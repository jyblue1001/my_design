magic
tech sky130A
magscale 1 2
timestamp 1751881932
<< error_p >>
rect 49250 -3550 49282 -3490
rect 49250 -4540 49268 -3550
<< nwell >>
rect 5930 6520 6950 7190
rect 7210 6520 9110 7190
rect 9370 6530 10390 7190
rect 5290 5400 6100 6060
rect 6360 5190 9960 6260
rect 10220 5400 11020 6060
rect 5260 4220 8020 4880
rect 8300 4220 11060 4880
rect 35930 3520 36950 4190
rect 37210 3520 39110 4190
rect 39370 3530 40390 4190
rect 35290 2400 36100 3060
rect 36360 2190 39960 3260
rect 40220 2400 41020 3060
rect 35260 1220 38020 1880
rect 38300 1220 41060 1880
<< pwell >>
rect 40 6840 2480 7330
rect 40 6310 2420 6800
rect 430 5890 2050 6270
rect 2610 6090 5020 7060
rect 430 5470 2050 5850
rect 2940 5680 4610 6050
rect 6150 3600 7650 4190
rect 8670 3600 10170 4190
rect -90 3370 260 3450
rect 5670 2650 8130 3540
rect 8190 2650 10650 3540
rect 5870 2100 10440 2610
rect 8440 2060 8852 2062
rect 6230 1460 7410 2060
rect 7460 1460 8860 2060
rect 8910 1460 10090 2060
rect 36150 600 37650 1190
rect 38670 600 40170 1190
rect 35670 -350 38130 540
rect 38190 -350 40650 540
rect 35870 -900 40440 -390
rect 38440 -940 38852 -938
rect 36230 -1540 37410 -940
rect 37460 -1540 38860 -940
rect 38910 -1540 40090 -940
rect 44040 -3160 46480 -2670
rect 44040 -3690 46420 -3200
rect 44430 -4110 46050 -3730
rect 46610 -3910 49020 -2940
rect 33590 -4373 34930 -4220
rect 33590 -5407 33743 -4373
rect 34777 -5407 34930 -4373
rect 33590 -5560 34930 -5407
rect 34950 -4373 36290 -4220
rect 34950 -5407 35103 -4373
rect 36137 -5407 36290 -4373
rect 34950 -5560 36290 -5407
rect 36310 -4373 37650 -4220
rect 36310 -5407 36463 -4373
rect 37497 -5407 37650 -4373
rect 44430 -4530 46050 -4150
rect 46940 -4320 48610 -3950
rect 36310 -5560 37650 -5407
rect 37640 -5580 37650 -5560
rect 33590 -5733 34930 -5580
rect 33590 -6767 33743 -5733
rect 34777 -6767 34930 -5733
rect 33590 -6920 34930 -6767
rect 34950 -5733 36290 -5580
rect 34950 -6767 35103 -5733
rect 36137 -6767 36290 -5733
rect 34950 -6920 36290 -6767
rect 36310 -5733 37650 -5580
rect 36310 -6767 36463 -5733
rect 37497 -6767 37650 -5733
rect 36310 -6920 37650 -6767
rect 37640 -6940 37650 -6920
rect 33590 -7093 34930 -6940
rect 33590 -8127 33743 -7093
rect 34777 -8127 34930 -7093
rect 33590 -8280 34930 -8127
rect 34950 -7093 36290 -6940
rect 34950 -8127 35103 -7093
rect 36137 -8127 36290 -7093
rect 34950 -8280 36290 -8127
rect 36310 -7093 37650 -6940
rect 36310 -8127 36463 -7093
rect 37497 -8127 37650 -7093
rect 36310 -8280 37650 -8127
rect 35560 -8600 35640 -8280
<< nbase >>
rect 33743 -5407 34777 -4373
rect 35103 -5407 36137 -4373
rect 36463 -5407 37497 -4373
rect 33743 -6767 34777 -5733
rect 35103 -6767 36137 -5733
rect 36463 -6767 37497 -5733
rect 33743 -8127 34777 -7093
rect 35103 -8127 36137 -7093
rect 36463 -8127 37497 -7093
<< nmos >>
rect 6340 3800 6380 3900
rect 6460 3800 6500 3900
rect 6580 3800 6620 3900
rect 6700 3800 6740 3900
rect 6820 3800 6860 3900
rect 6940 3800 6980 3900
rect 7060 3800 7100 3900
rect 7180 3800 7220 3900
rect 7300 3800 7340 3900
rect 7420 3800 7460 3900
rect 8860 3800 8900 3900
rect 8980 3800 9020 3900
rect 9100 3800 9140 3900
rect 9220 3800 9260 3900
rect 9340 3800 9380 3900
rect 9460 3800 9500 3900
rect 9580 3800 9620 3900
rect 9700 3800 9740 3900
rect 9820 3800 9860 3900
rect 9940 3800 9980 3900
rect 5860 2850 6860 3350
rect 6940 2850 7940 3350
rect 8380 2850 9380 3350
rect 9460 2850 10460 3350
rect 6120 2210 8120 2410
rect 8200 2210 10200 2410
rect 6420 1660 6450 1860
rect 6530 1660 6560 1860
rect 6640 1660 6670 1860
rect 6750 1660 6780 1860
rect 6860 1660 6890 1860
rect 6970 1660 7000 1860
rect 7080 1660 7110 1860
rect 7190 1660 7220 1860
rect 7650 1660 7680 1860
rect 7760 1660 7790 1860
rect 7870 1660 7900 1860
rect 7980 1660 8010 1860
rect 8090 1660 8120 1860
rect 8200 1660 8230 1860
rect 8310 1660 8340 1860
rect 8420 1660 8450 1860
rect 8530 1660 8560 1860
rect 8640 1660 8670 1860
rect 9100 1660 9130 1860
rect 9210 1660 9240 1860
rect 9320 1660 9350 1860
rect 9430 1660 9460 1860
rect 9540 1660 9570 1860
rect 9650 1660 9680 1860
rect 9760 1660 9790 1860
rect 9870 1660 9900 1860
rect 36340 800 36380 900
rect 36460 800 36500 900
rect 36580 800 36620 900
rect 36700 800 36740 900
rect 36820 800 36860 900
rect 36940 800 36980 900
rect 37060 800 37100 900
rect 37180 800 37220 900
rect 37300 800 37340 900
rect 37420 800 37460 900
rect 38860 800 38900 900
rect 38980 800 39020 900
rect 39100 800 39140 900
rect 39220 800 39260 900
rect 39340 800 39380 900
rect 39460 800 39500 900
rect 39580 800 39620 900
rect 39700 800 39740 900
rect 39820 800 39860 900
rect 39940 800 39980 900
rect 35860 -150 36860 350
rect 36940 -150 37940 350
rect 38380 -150 39380 350
rect 39460 -150 40460 350
rect 36120 -790 38120 -590
rect 38200 -790 40200 -590
rect 36420 -1340 36450 -1140
rect 36530 -1340 36560 -1140
rect 36640 -1340 36670 -1140
rect 36750 -1340 36780 -1140
rect 36860 -1340 36890 -1140
rect 36970 -1340 37000 -1140
rect 37080 -1340 37110 -1140
rect 37190 -1340 37220 -1140
rect 37650 -1340 37680 -1140
rect 37760 -1340 37790 -1140
rect 37870 -1340 37900 -1140
rect 37980 -1340 38010 -1140
rect 38090 -1340 38120 -1140
rect 38200 -1340 38230 -1140
rect 38310 -1340 38340 -1140
rect 38420 -1340 38450 -1140
rect 38530 -1340 38560 -1140
rect 38640 -1340 38670 -1140
rect 39100 -1340 39130 -1140
rect 39210 -1340 39240 -1140
rect 39320 -1340 39350 -1140
rect 39430 -1340 39460 -1140
rect 39540 -1340 39570 -1140
rect 39650 -1340 39680 -1140
rect 39760 -1340 39790 -1140
rect 39870 -1340 39900 -1140
<< pmos >>
rect 6150 6760 6180 6960
rect 6260 6760 6290 6960
rect 6370 6760 6400 6960
rect 6480 6760 6510 6960
rect 6590 6760 6620 6960
rect 6700 6760 6730 6960
rect 7430 6760 7460 6960
rect 7540 6760 7570 6960
rect 7650 6760 7680 6960
rect 7760 6760 7790 6960
rect 7870 6760 7900 6960
rect 7980 6760 8010 6960
rect 8090 6760 8120 6960
rect 8200 6760 8230 6960
rect 8310 6760 8340 6960
rect 8420 6760 8450 6960
rect 8530 6760 8560 6960
rect 8640 6760 8670 6960
rect 9590 6760 9620 6960
rect 9700 6760 9730 6960
rect 9810 6760 9840 6960
rect 9920 6760 9950 6960
rect 10030 6760 10060 6960
rect 10140 6760 10170 6960
rect 5510 5630 5540 5830
rect 5620 5630 5650 5830
rect 5730 5630 5760 5830
rect 5840 5630 5870 5830
rect 6580 5430 6680 6030
rect 6760 5430 6860 6030
rect 6940 5430 7040 6030
rect 7120 5430 7220 6030
rect 7300 5430 7400 6030
rect 7480 5430 7580 6030
rect 7660 5430 7760 6030
rect 7840 5430 7940 6030
rect 8020 5430 8120 6030
rect 8200 5430 8300 6030
rect 8380 5430 8480 6030
rect 8560 5430 8660 6030
rect 8740 5430 8840 6030
rect 8920 5430 9020 6030
rect 9100 5430 9200 6030
rect 9280 5430 9380 6030
rect 9460 5430 9560 6030
rect 9640 5430 9740 6030
rect 10440 5630 10470 5830
rect 10550 5630 10580 5830
rect 10660 5630 10690 5830
rect 10770 5630 10800 5830
rect 5480 4450 5520 4650
rect 5600 4450 5640 4650
rect 5720 4450 5760 4650
rect 5840 4450 5880 4650
rect 5960 4450 6000 4650
rect 6080 4450 6120 4650
rect 6200 4450 6240 4650
rect 6320 4450 6360 4650
rect 6440 4450 6480 4650
rect 6560 4450 6600 4650
rect 6680 4450 6720 4650
rect 6800 4450 6840 4650
rect 6920 4450 6960 4650
rect 7040 4450 7080 4650
rect 7160 4450 7200 4650
rect 7280 4450 7320 4650
rect 7400 4450 7440 4650
rect 7520 4450 7560 4650
rect 7640 4450 7680 4650
rect 7760 4450 7800 4650
rect 8520 4450 8560 4650
rect 8640 4450 8680 4650
rect 8760 4450 8800 4650
rect 8880 4450 8920 4650
rect 9000 4450 9040 4650
rect 9120 4450 9160 4650
rect 9240 4450 9280 4650
rect 9360 4450 9400 4650
rect 9480 4450 9520 4650
rect 9600 4450 9640 4650
rect 9720 4450 9760 4650
rect 9840 4450 9880 4650
rect 9960 4450 10000 4650
rect 10080 4450 10120 4650
rect 10200 4450 10240 4650
rect 10320 4450 10360 4650
rect 10440 4450 10480 4650
rect 10560 4450 10600 4650
rect 10680 4450 10720 4650
rect 10800 4450 10840 4650
rect 36150 3760 36180 3960
rect 36260 3760 36290 3960
rect 36370 3760 36400 3960
rect 36480 3760 36510 3960
rect 36590 3760 36620 3960
rect 36700 3760 36730 3960
rect 37430 3760 37460 3960
rect 37540 3760 37570 3960
rect 37650 3760 37680 3960
rect 37760 3760 37790 3960
rect 37870 3760 37900 3960
rect 37980 3760 38010 3960
rect 38090 3760 38120 3960
rect 38200 3760 38230 3960
rect 38310 3760 38340 3960
rect 38420 3760 38450 3960
rect 38530 3760 38560 3960
rect 38640 3760 38670 3960
rect 39590 3760 39620 3960
rect 39700 3760 39730 3960
rect 39810 3760 39840 3960
rect 39920 3760 39950 3960
rect 40030 3760 40060 3960
rect 40140 3760 40170 3960
rect 35510 2630 35540 2830
rect 35620 2630 35650 2830
rect 35730 2630 35760 2830
rect 35840 2630 35870 2830
rect 36580 2430 36680 3030
rect 36760 2430 36860 3030
rect 36940 2430 37040 3030
rect 37120 2430 37220 3030
rect 37300 2430 37400 3030
rect 37480 2430 37580 3030
rect 37660 2430 37760 3030
rect 37840 2430 37940 3030
rect 38020 2430 38120 3030
rect 38200 2430 38300 3030
rect 38380 2430 38480 3030
rect 38560 2430 38660 3030
rect 38740 2430 38840 3030
rect 38920 2430 39020 3030
rect 39100 2430 39200 3030
rect 39280 2430 39380 3030
rect 39460 2430 39560 3030
rect 39640 2430 39740 3030
rect 40440 2630 40470 2830
rect 40550 2630 40580 2830
rect 40660 2630 40690 2830
rect 40770 2630 40800 2830
rect 35480 1450 35520 1650
rect 35600 1450 35640 1650
rect 35720 1450 35760 1650
rect 35840 1450 35880 1650
rect 35960 1450 36000 1650
rect 36080 1450 36120 1650
rect 36200 1450 36240 1650
rect 36320 1450 36360 1650
rect 36440 1450 36480 1650
rect 36560 1450 36600 1650
rect 36680 1450 36720 1650
rect 36800 1450 36840 1650
rect 36920 1450 36960 1650
rect 37040 1450 37080 1650
rect 37160 1450 37200 1650
rect 37280 1450 37320 1650
rect 37400 1450 37440 1650
rect 37520 1450 37560 1650
rect 37640 1450 37680 1650
rect 37760 1450 37800 1650
rect 38520 1450 38560 1650
rect 38640 1450 38680 1650
rect 38760 1450 38800 1650
rect 38880 1450 38920 1650
rect 39000 1450 39040 1650
rect 39120 1450 39160 1650
rect 39240 1450 39280 1650
rect 39360 1450 39400 1650
rect 39480 1450 39520 1650
rect 39600 1450 39640 1650
rect 39720 1450 39760 1650
rect 39840 1450 39880 1650
rect 39960 1450 40000 1650
rect 40080 1450 40120 1650
rect 40200 1450 40240 1650
rect 40320 1450 40360 1650
rect 40440 1450 40480 1650
rect 40560 1450 40600 1650
rect 40680 1450 40720 1650
rect 40800 1450 40840 1650
<< ndiff >>
rect 6260 3870 6340 3900
rect 6260 3830 6280 3870
rect 6320 3830 6340 3870
rect 6260 3800 6340 3830
rect 6380 3870 6460 3900
rect 6380 3830 6400 3870
rect 6440 3830 6460 3870
rect 6380 3800 6460 3830
rect 6500 3870 6580 3900
rect 6500 3830 6520 3870
rect 6560 3830 6580 3870
rect 6500 3800 6580 3830
rect 6620 3870 6700 3900
rect 6620 3830 6640 3870
rect 6680 3830 6700 3870
rect 6620 3800 6700 3830
rect 6740 3870 6820 3900
rect 6740 3830 6760 3870
rect 6800 3830 6820 3870
rect 6740 3800 6820 3830
rect 6860 3870 6940 3900
rect 6860 3830 6880 3870
rect 6920 3830 6940 3870
rect 6860 3800 6940 3830
rect 6980 3870 7060 3900
rect 6980 3830 7000 3870
rect 7040 3830 7060 3870
rect 6980 3800 7060 3830
rect 7100 3870 7180 3900
rect 7100 3830 7120 3870
rect 7160 3830 7180 3870
rect 7100 3800 7180 3830
rect 7220 3870 7300 3900
rect 7220 3830 7240 3870
rect 7280 3830 7300 3870
rect 7220 3800 7300 3830
rect 7340 3870 7420 3900
rect 7340 3830 7360 3870
rect 7400 3830 7420 3870
rect 7340 3800 7420 3830
rect 7460 3870 7540 3900
rect 7460 3830 7480 3870
rect 7520 3830 7540 3870
rect 7460 3800 7540 3830
rect 8780 3870 8860 3900
rect 8780 3830 8800 3870
rect 8840 3830 8860 3870
rect 8780 3800 8860 3830
rect 8900 3870 8980 3900
rect 8900 3830 8920 3870
rect 8960 3830 8980 3870
rect 8900 3800 8980 3830
rect 9020 3870 9100 3900
rect 9020 3830 9040 3870
rect 9080 3830 9100 3870
rect 9020 3800 9100 3830
rect 9140 3870 9220 3900
rect 9140 3830 9160 3870
rect 9200 3830 9220 3870
rect 9140 3800 9220 3830
rect 9260 3870 9340 3900
rect 9260 3830 9280 3870
rect 9320 3830 9340 3870
rect 9260 3800 9340 3830
rect 9380 3870 9460 3900
rect 9380 3830 9400 3870
rect 9440 3830 9460 3870
rect 9380 3800 9460 3830
rect 9500 3870 9580 3900
rect 9500 3830 9520 3870
rect 9560 3830 9580 3870
rect 9500 3800 9580 3830
rect 9620 3870 9700 3900
rect 9620 3830 9640 3870
rect 9680 3830 9700 3870
rect 9620 3800 9700 3830
rect 9740 3870 9820 3900
rect 9740 3830 9760 3870
rect 9800 3830 9820 3870
rect 9740 3800 9820 3830
rect 9860 3870 9940 3900
rect 9860 3830 9880 3870
rect 9920 3830 9940 3870
rect 9860 3800 9940 3830
rect 9980 3870 10060 3900
rect 9980 3830 10000 3870
rect 10040 3830 10060 3870
rect 9980 3800 10060 3830
rect 5780 3320 5860 3350
rect 5780 3280 5800 3320
rect 5840 3280 5860 3320
rect 5780 3220 5860 3280
rect 5780 3180 5800 3220
rect 5840 3180 5860 3220
rect 5780 3120 5860 3180
rect 5780 3080 5800 3120
rect 5840 3080 5860 3120
rect 5780 3020 5860 3080
rect 5780 2980 5800 3020
rect 5840 2980 5860 3020
rect 5780 2920 5860 2980
rect 5780 2880 5800 2920
rect 5840 2880 5860 2920
rect 5780 2850 5860 2880
rect 6860 3320 6940 3350
rect 6860 3280 6880 3320
rect 6920 3280 6940 3320
rect 6860 3220 6940 3280
rect 6860 3180 6880 3220
rect 6920 3180 6940 3220
rect 6860 3120 6940 3180
rect 6860 3080 6880 3120
rect 6920 3080 6940 3120
rect 6860 3020 6940 3080
rect 6860 2980 6880 3020
rect 6920 2980 6940 3020
rect 6860 2920 6940 2980
rect 6860 2880 6880 2920
rect 6920 2880 6940 2920
rect 6860 2850 6940 2880
rect 7940 3320 8020 3350
rect 7940 3280 7960 3320
rect 8000 3280 8020 3320
rect 7940 3220 8020 3280
rect 7940 3180 7960 3220
rect 8000 3180 8020 3220
rect 7940 3120 8020 3180
rect 7940 3080 7960 3120
rect 8000 3080 8020 3120
rect 7940 3020 8020 3080
rect 7940 2980 7960 3020
rect 8000 2980 8020 3020
rect 7940 2920 8020 2980
rect 7940 2880 7960 2920
rect 8000 2880 8020 2920
rect 7940 2850 8020 2880
rect 8300 3320 8380 3350
rect 8300 3280 8320 3320
rect 8360 3280 8380 3320
rect 8300 3220 8380 3280
rect 8300 3180 8320 3220
rect 8360 3180 8380 3220
rect 8300 3120 8380 3180
rect 8300 3080 8320 3120
rect 8360 3080 8380 3120
rect 8300 3020 8380 3080
rect 8300 2980 8320 3020
rect 8360 2980 8380 3020
rect 8300 2920 8380 2980
rect 8300 2880 8320 2920
rect 8360 2880 8380 2920
rect 8300 2850 8380 2880
rect 9380 3320 9460 3350
rect 9380 3280 9400 3320
rect 9440 3280 9460 3320
rect 9380 3220 9460 3280
rect 9380 3180 9400 3220
rect 9440 3180 9460 3220
rect 9380 3120 9460 3180
rect 9380 3080 9400 3120
rect 9440 3080 9460 3120
rect 9380 3020 9460 3080
rect 9380 2980 9400 3020
rect 9440 2980 9460 3020
rect 9380 2920 9460 2980
rect 9380 2880 9400 2920
rect 9440 2880 9460 2920
rect 9380 2850 9460 2880
rect 10460 3320 10540 3350
rect 10460 3280 10480 3320
rect 10520 3280 10540 3320
rect 10460 3220 10540 3280
rect 10460 3180 10480 3220
rect 10520 3180 10540 3220
rect 10460 3120 10540 3180
rect 10460 3080 10480 3120
rect 10520 3080 10540 3120
rect 10460 3020 10540 3080
rect 10460 2980 10480 3020
rect 10520 2980 10540 3020
rect 10460 2920 10540 2980
rect 10460 2880 10480 2920
rect 10520 2880 10540 2920
rect 10460 2850 10540 2880
rect 6040 2380 6120 2410
rect 6040 2340 6060 2380
rect 6100 2340 6120 2380
rect 6040 2280 6120 2340
rect 6040 2240 6060 2280
rect 6100 2240 6120 2280
rect 6040 2210 6120 2240
rect 8120 2380 8200 2410
rect 8120 2340 8140 2380
rect 8180 2340 8200 2380
rect 8120 2280 8200 2340
rect 8120 2240 8140 2280
rect 8180 2240 8200 2280
rect 8120 2210 8200 2240
rect 10200 2380 10280 2410
rect 10200 2340 10220 2380
rect 10260 2340 10280 2380
rect 10200 2280 10280 2340
rect 10200 2240 10220 2280
rect 10260 2240 10280 2280
rect 10200 2210 10280 2240
rect 6340 1830 6420 1860
rect 6340 1790 6360 1830
rect 6400 1790 6420 1830
rect 6340 1730 6420 1790
rect 6340 1690 6360 1730
rect 6400 1690 6420 1730
rect 6340 1660 6420 1690
rect 6450 1830 6530 1860
rect 6450 1790 6470 1830
rect 6510 1790 6530 1830
rect 6450 1730 6530 1790
rect 6450 1690 6470 1730
rect 6510 1690 6530 1730
rect 6450 1660 6530 1690
rect 6560 1830 6640 1860
rect 6560 1790 6580 1830
rect 6620 1790 6640 1830
rect 6560 1730 6640 1790
rect 6560 1690 6580 1730
rect 6620 1690 6640 1730
rect 6560 1660 6640 1690
rect 6670 1830 6750 1860
rect 6670 1790 6690 1830
rect 6730 1790 6750 1830
rect 6670 1730 6750 1790
rect 6670 1690 6690 1730
rect 6730 1690 6750 1730
rect 6670 1660 6750 1690
rect 6780 1830 6860 1860
rect 6780 1790 6800 1830
rect 6840 1790 6860 1830
rect 6780 1730 6860 1790
rect 6780 1690 6800 1730
rect 6840 1690 6860 1730
rect 6780 1660 6860 1690
rect 6890 1830 6970 1860
rect 6890 1790 6910 1830
rect 6950 1790 6970 1830
rect 6890 1730 6970 1790
rect 6890 1690 6910 1730
rect 6950 1690 6970 1730
rect 6890 1660 6970 1690
rect 7000 1830 7080 1860
rect 7000 1790 7020 1830
rect 7060 1790 7080 1830
rect 7000 1730 7080 1790
rect 7000 1690 7020 1730
rect 7060 1690 7080 1730
rect 7000 1660 7080 1690
rect 7110 1830 7190 1860
rect 7110 1790 7130 1830
rect 7170 1790 7190 1830
rect 7110 1730 7190 1790
rect 7110 1690 7130 1730
rect 7170 1690 7190 1730
rect 7110 1660 7190 1690
rect 7220 1830 7300 1860
rect 7220 1790 7240 1830
rect 7280 1790 7300 1830
rect 7220 1730 7300 1790
rect 7220 1690 7240 1730
rect 7280 1690 7300 1730
rect 7220 1660 7300 1690
rect 7570 1830 7650 1860
rect 7570 1790 7590 1830
rect 7630 1790 7650 1830
rect 7570 1730 7650 1790
rect 7570 1690 7590 1730
rect 7630 1690 7650 1730
rect 7570 1660 7650 1690
rect 7680 1830 7760 1860
rect 7680 1790 7700 1830
rect 7740 1790 7760 1830
rect 7680 1730 7760 1790
rect 7680 1690 7700 1730
rect 7740 1690 7760 1730
rect 7680 1660 7760 1690
rect 7790 1830 7870 1860
rect 7790 1790 7810 1830
rect 7850 1790 7870 1830
rect 7790 1730 7870 1790
rect 7790 1690 7810 1730
rect 7850 1690 7870 1730
rect 7790 1660 7870 1690
rect 7900 1830 7980 1860
rect 7900 1790 7920 1830
rect 7960 1790 7980 1830
rect 7900 1730 7980 1790
rect 7900 1690 7920 1730
rect 7960 1690 7980 1730
rect 7900 1660 7980 1690
rect 8010 1830 8090 1860
rect 8010 1790 8030 1830
rect 8070 1790 8090 1830
rect 8010 1730 8090 1790
rect 8010 1690 8030 1730
rect 8070 1690 8090 1730
rect 8010 1660 8090 1690
rect 8120 1830 8200 1860
rect 8120 1790 8140 1830
rect 8180 1790 8200 1830
rect 8120 1730 8200 1790
rect 8120 1690 8140 1730
rect 8180 1690 8200 1730
rect 8120 1660 8200 1690
rect 8230 1830 8310 1860
rect 8230 1790 8250 1830
rect 8290 1790 8310 1830
rect 8230 1730 8310 1790
rect 8230 1690 8250 1730
rect 8290 1690 8310 1730
rect 8230 1660 8310 1690
rect 8340 1830 8420 1860
rect 8340 1790 8360 1830
rect 8400 1790 8420 1830
rect 8340 1730 8420 1790
rect 8340 1690 8360 1730
rect 8400 1690 8420 1730
rect 8340 1660 8420 1690
rect 8450 1830 8530 1860
rect 8450 1790 8470 1830
rect 8510 1790 8530 1830
rect 8450 1730 8530 1790
rect 8450 1690 8470 1730
rect 8510 1690 8530 1730
rect 8450 1660 8530 1690
rect 8560 1830 8640 1860
rect 8560 1790 8580 1830
rect 8620 1790 8640 1830
rect 8560 1730 8640 1790
rect 8560 1690 8580 1730
rect 8620 1690 8640 1730
rect 8560 1660 8640 1690
rect 8670 1830 8750 1860
rect 8670 1790 8690 1830
rect 8730 1790 8750 1830
rect 8670 1730 8750 1790
rect 8670 1690 8690 1730
rect 8730 1690 8750 1730
rect 8670 1660 8750 1690
rect 9020 1830 9100 1860
rect 9020 1790 9040 1830
rect 9080 1790 9100 1830
rect 9020 1730 9100 1790
rect 9020 1690 9040 1730
rect 9080 1690 9100 1730
rect 9020 1660 9100 1690
rect 9130 1830 9210 1860
rect 9130 1790 9150 1830
rect 9190 1790 9210 1830
rect 9130 1730 9210 1790
rect 9130 1690 9150 1730
rect 9190 1690 9210 1730
rect 9130 1660 9210 1690
rect 9240 1830 9320 1860
rect 9240 1790 9260 1830
rect 9300 1790 9320 1830
rect 9240 1730 9320 1790
rect 9240 1690 9260 1730
rect 9300 1690 9320 1730
rect 9240 1660 9320 1690
rect 9350 1830 9430 1860
rect 9350 1790 9370 1830
rect 9410 1790 9430 1830
rect 9350 1730 9430 1790
rect 9350 1690 9370 1730
rect 9410 1690 9430 1730
rect 9350 1660 9430 1690
rect 9460 1830 9540 1860
rect 9460 1790 9480 1830
rect 9520 1790 9540 1830
rect 9460 1730 9540 1790
rect 9460 1690 9480 1730
rect 9520 1690 9540 1730
rect 9460 1660 9540 1690
rect 9570 1830 9650 1860
rect 9570 1790 9590 1830
rect 9630 1790 9650 1830
rect 9570 1730 9650 1790
rect 9570 1690 9590 1730
rect 9630 1690 9650 1730
rect 9570 1660 9650 1690
rect 9680 1830 9760 1860
rect 9680 1790 9700 1830
rect 9740 1790 9760 1830
rect 9680 1730 9760 1790
rect 9680 1690 9700 1730
rect 9740 1690 9760 1730
rect 9680 1660 9760 1690
rect 9790 1830 9870 1860
rect 9790 1790 9810 1830
rect 9850 1790 9870 1830
rect 9790 1730 9870 1790
rect 9790 1690 9810 1730
rect 9850 1690 9870 1730
rect 9790 1660 9870 1690
rect 9900 1830 9980 1860
rect 9900 1790 9920 1830
rect 9960 1790 9980 1830
rect 9900 1730 9980 1790
rect 9900 1690 9920 1730
rect 9960 1690 9980 1730
rect 9900 1660 9980 1690
rect 36260 870 36340 900
rect 36260 830 36280 870
rect 36320 830 36340 870
rect 36260 800 36340 830
rect 36380 870 36460 900
rect 36380 830 36400 870
rect 36440 830 36460 870
rect 36380 800 36460 830
rect 36500 870 36580 900
rect 36500 830 36520 870
rect 36560 830 36580 870
rect 36500 800 36580 830
rect 36620 870 36700 900
rect 36620 830 36640 870
rect 36680 830 36700 870
rect 36620 800 36700 830
rect 36740 870 36820 900
rect 36740 830 36760 870
rect 36800 830 36820 870
rect 36740 800 36820 830
rect 36860 870 36940 900
rect 36860 830 36880 870
rect 36920 830 36940 870
rect 36860 800 36940 830
rect 36980 870 37060 900
rect 36980 830 37000 870
rect 37040 830 37060 870
rect 36980 800 37060 830
rect 37100 870 37180 900
rect 37100 830 37120 870
rect 37160 830 37180 870
rect 37100 800 37180 830
rect 37220 870 37300 900
rect 37220 830 37240 870
rect 37280 830 37300 870
rect 37220 800 37300 830
rect 37340 870 37420 900
rect 37340 830 37360 870
rect 37400 830 37420 870
rect 37340 800 37420 830
rect 37460 870 37540 900
rect 37460 830 37480 870
rect 37520 830 37540 870
rect 37460 800 37540 830
rect 38780 870 38860 900
rect 38780 830 38800 870
rect 38840 830 38860 870
rect 38780 800 38860 830
rect 38900 870 38980 900
rect 38900 830 38920 870
rect 38960 830 38980 870
rect 38900 800 38980 830
rect 39020 870 39100 900
rect 39020 830 39040 870
rect 39080 830 39100 870
rect 39020 800 39100 830
rect 39140 870 39220 900
rect 39140 830 39160 870
rect 39200 830 39220 870
rect 39140 800 39220 830
rect 39260 870 39340 900
rect 39260 830 39280 870
rect 39320 830 39340 870
rect 39260 800 39340 830
rect 39380 870 39460 900
rect 39380 830 39400 870
rect 39440 830 39460 870
rect 39380 800 39460 830
rect 39500 870 39580 900
rect 39500 830 39520 870
rect 39560 830 39580 870
rect 39500 800 39580 830
rect 39620 870 39700 900
rect 39620 830 39640 870
rect 39680 830 39700 870
rect 39620 800 39700 830
rect 39740 870 39820 900
rect 39740 830 39760 870
rect 39800 830 39820 870
rect 39740 800 39820 830
rect 39860 870 39940 900
rect 39860 830 39880 870
rect 39920 830 39940 870
rect 39860 800 39940 830
rect 39980 870 40060 900
rect 39980 830 40000 870
rect 40040 830 40060 870
rect 39980 800 40060 830
rect 35780 320 35860 350
rect 35780 280 35800 320
rect 35840 280 35860 320
rect 35780 220 35860 280
rect 35780 180 35800 220
rect 35840 180 35860 220
rect 35780 120 35860 180
rect 35780 80 35800 120
rect 35840 80 35860 120
rect 35780 20 35860 80
rect 35780 -20 35800 20
rect 35840 -20 35860 20
rect 35780 -80 35860 -20
rect 35780 -120 35800 -80
rect 35840 -120 35860 -80
rect 35780 -150 35860 -120
rect 36860 320 36940 350
rect 36860 280 36880 320
rect 36920 280 36940 320
rect 36860 220 36940 280
rect 36860 180 36880 220
rect 36920 180 36940 220
rect 36860 120 36940 180
rect 36860 80 36880 120
rect 36920 80 36940 120
rect 36860 20 36940 80
rect 36860 -20 36880 20
rect 36920 -20 36940 20
rect 36860 -80 36940 -20
rect 36860 -120 36880 -80
rect 36920 -120 36940 -80
rect 36860 -150 36940 -120
rect 37940 320 38020 350
rect 37940 280 37960 320
rect 38000 280 38020 320
rect 37940 220 38020 280
rect 37940 180 37960 220
rect 38000 180 38020 220
rect 37940 120 38020 180
rect 37940 80 37960 120
rect 38000 80 38020 120
rect 37940 20 38020 80
rect 37940 -20 37960 20
rect 38000 -20 38020 20
rect 37940 -80 38020 -20
rect 37940 -120 37960 -80
rect 38000 -120 38020 -80
rect 37940 -150 38020 -120
rect 38300 320 38380 350
rect 38300 280 38320 320
rect 38360 280 38380 320
rect 38300 220 38380 280
rect 38300 180 38320 220
rect 38360 180 38380 220
rect 38300 120 38380 180
rect 38300 80 38320 120
rect 38360 80 38380 120
rect 38300 20 38380 80
rect 38300 -20 38320 20
rect 38360 -20 38380 20
rect 38300 -80 38380 -20
rect 38300 -120 38320 -80
rect 38360 -120 38380 -80
rect 38300 -150 38380 -120
rect 39380 320 39460 350
rect 39380 280 39400 320
rect 39440 280 39460 320
rect 39380 220 39460 280
rect 39380 180 39400 220
rect 39440 180 39460 220
rect 39380 120 39460 180
rect 39380 80 39400 120
rect 39440 80 39460 120
rect 39380 20 39460 80
rect 39380 -20 39400 20
rect 39440 -20 39460 20
rect 39380 -80 39460 -20
rect 39380 -120 39400 -80
rect 39440 -120 39460 -80
rect 39380 -150 39460 -120
rect 40460 320 40540 350
rect 40460 280 40480 320
rect 40520 280 40540 320
rect 40460 220 40540 280
rect 40460 180 40480 220
rect 40520 180 40540 220
rect 40460 120 40540 180
rect 40460 80 40480 120
rect 40520 80 40540 120
rect 40460 20 40540 80
rect 40460 -20 40480 20
rect 40520 -20 40540 20
rect 40460 -80 40540 -20
rect 40460 -120 40480 -80
rect 40520 -120 40540 -80
rect 40460 -150 40540 -120
rect 36040 -620 36120 -590
rect 36040 -660 36060 -620
rect 36100 -660 36120 -620
rect 36040 -720 36120 -660
rect 36040 -760 36060 -720
rect 36100 -760 36120 -720
rect 36040 -790 36120 -760
rect 38120 -620 38200 -590
rect 38120 -660 38140 -620
rect 38180 -660 38200 -620
rect 38120 -720 38200 -660
rect 38120 -760 38140 -720
rect 38180 -760 38200 -720
rect 38120 -790 38200 -760
rect 40200 -620 40280 -590
rect 40200 -660 40220 -620
rect 40260 -660 40280 -620
rect 40200 -720 40280 -660
rect 40200 -760 40220 -720
rect 40260 -760 40280 -720
rect 40200 -790 40280 -760
rect 36340 -1170 36420 -1140
rect 36340 -1210 36360 -1170
rect 36400 -1210 36420 -1170
rect 36340 -1270 36420 -1210
rect 36340 -1310 36360 -1270
rect 36400 -1310 36420 -1270
rect 36340 -1340 36420 -1310
rect 36450 -1170 36530 -1140
rect 36450 -1210 36470 -1170
rect 36510 -1210 36530 -1170
rect 36450 -1270 36530 -1210
rect 36450 -1310 36470 -1270
rect 36510 -1310 36530 -1270
rect 36450 -1340 36530 -1310
rect 36560 -1170 36640 -1140
rect 36560 -1210 36580 -1170
rect 36620 -1210 36640 -1170
rect 36560 -1270 36640 -1210
rect 36560 -1310 36580 -1270
rect 36620 -1310 36640 -1270
rect 36560 -1340 36640 -1310
rect 36670 -1170 36750 -1140
rect 36670 -1210 36690 -1170
rect 36730 -1210 36750 -1170
rect 36670 -1270 36750 -1210
rect 36670 -1310 36690 -1270
rect 36730 -1310 36750 -1270
rect 36670 -1340 36750 -1310
rect 36780 -1170 36860 -1140
rect 36780 -1210 36800 -1170
rect 36840 -1210 36860 -1170
rect 36780 -1270 36860 -1210
rect 36780 -1310 36800 -1270
rect 36840 -1310 36860 -1270
rect 36780 -1340 36860 -1310
rect 36890 -1170 36970 -1140
rect 36890 -1210 36910 -1170
rect 36950 -1210 36970 -1170
rect 36890 -1270 36970 -1210
rect 36890 -1310 36910 -1270
rect 36950 -1310 36970 -1270
rect 36890 -1340 36970 -1310
rect 37000 -1170 37080 -1140
rect 37000 -1210 37020 -1170
rect 37060 -1210 37080 -1170
rect 37000 -1270 37080 -1210
rect 37000 -1310 37020 -1270
rect 37060 -1310 37080 -1270
rect 37000 -1340 37080 -1310
rect 37110 -1170 37190 -1140
rect 37110 -1210 37130 -1170
rect 37170 -1210 37190 -1170
rect 37110 -1270 37190 -1210
rect 37110 -1310 37130 -1270
rect 37170 -1310 37190 -1270
rect 37110 -1340 37190 -1310
rect 37220 -1170 37300 -1140
rect 37220 -1210 37240 -1170
rect 37280 -1210 37300 -1170
rect 37220 -1270 37300 -1210
rect 37220 -1310 37240 -1270
rect 37280 -1310 37300 -1270
rect 37220 -1340 37300 -1310
rect 37570 -1170 37650 -1140
rect 37570 -1210 37590 -1170
rect 37630 -1210 37650 -1170
rect 37570 -1270 37650 -1210
rect 37570 -1310 37590 -1270
rect 37630 -1310 37650 -1270
rect 37570 -1340 37650 -1310
rect 37680 -1170 37760 -1140
rect 37680 -1210 37700 -1170
rect 37740 -1210 37760 -1170
rect 37680 -1270 37760 -1210
rect 37680 -1310 37700 -1270
rect 37740 -1310 37760 -1270
rect 37680 -1340 37760 -1310
rect 37790 -1170 37870 -1140
rect 37790 -1210 37810 -1170
rect 37850 -1210 37870 -1170
rect 37790 -1270 37870 -1210
rect 37790 -1310 37810 -1270
rect 37850 -1310 37870 -1270
rect 37790 -1340 37870 -1310
rect 37900 -1170 37980 -1140
rect 37900 -1210 37920 -1170
rect 37960 -1210 37980 -1170
rect 37900 -1270 37980 -1210
rect 37900 -1310 37920 -1270
rect 37960 -1310 37980 -1270
rect 37900 -1340 37980 -1310
rect 38010 -1170 38090 -1140
rect 38010 -1210 38030 -1170
rect 38070 -1210 38090 -1170
rect 38010 -1270 38090 -1210
rect 38010 -1310 38030 -1270
rect 38070 -1310 38090 -1270
rect 38010 -1340 38090 -1310
rect 38120 -1170 38200 -1140
rect 38120 -1210 38140 -1170
rect 38180 -1210 38200 -1170
rect 38120 -1270 38200 -1210
rect 38120 -1310 38140 -1270
rect 38180 -1310 38200 -1270
rect 38120 -1340 38200 -1310
rect 38230 -1170 38310 -1140
rect 38230 -1210 38250 -1170
rect 38290 -1210 38310 -1170
rect 38230 -1270 38310 -1210
rect 38230 -1310 38250 -1270
rect 38290 -1310 38310 -1270
rect 38230 -1340 38310 -1310
rect 38340 -1170 38420 -1140
rect 38340 -1210 38360 -1170
rect 38400 -1210 38420 -1170
rect 38340 -1270 38420 -1210
rect 38340 -1310 38360 -1270
rect 38400 -1310 38420 -1270
rect 38340 -1340 38420 -1310
rect 38450 -1170 38530 -1140
rect 38450 -1210 38470 -1170
rect 38510 -1210 38530 -1170
rect 38450 -1270 38530 -1210
rect 38450 -1310 38470 -1270
rect 38510 -1310 38530 -1270
rect 38450 -1340 38530 -1310
rect 38560 -1170 38640 -1140
rect 38560 -1210 38580 -1170
rect 38620 -1210 38640 -1170
rect 38560 -1270 38640 -1210
rect 38560 -1310 38580 -1270
rect 38620 -1310 38640 -1270
rect 38560 -1340 38640 -1310
rect 38670 -1170 38750 -1140
rect 38670 -1210 38690 -1170
rect 38730 -1210 38750 -1170
rect 38670 -1270 38750 -1210
rect 38670 -1310 38690 -1270
rect 38730 -1310 38750 -1270
rect 38670 -1340 38750 -1310
rect 39020 -1170 39100 -1140
rect 39020 -1210 39040 -1170
rect 39080 -1210 39100 -1170
rect 39020 -1270 39100 -1210
rect 39020 -1310 39040 -1270
rect 39080 -1310 39100 -1270
rect 39020 -1340 39100 -1310
rect 39130 -1170 39210 -1140
rect 39130 -1210 39150 -1170
rect 39190 -1210 39210 -1170
rect 39130 -1270 39210 -1210
rect 39130 -1310 39150 -1270
rect 39190 -1310 39210 -1270
rect 39130 -1340 39210 -1310
rect 39240 -1170 39320 -1140
rect 39240 -1210 39260 -1170
rect 39300 -1210 39320 -1170
rect 39240 -1270 39320 -1210
rect 39240 -1310 39260 -1270
rect 39300 -1310 39320 -1270
rect 39240 -1340 39320 -1310
rect 39350 -1170 39430 -1140
rect 39350 -1210 39370 -1170
rect 39410 -1210 39430 -1170
rect 39350 -1270 39430 -1210
rect 39350 -1310 39370 -1270
rect 39410 -1310 39430 -1270
rect 39350 -1340 39430 -1310
rect 39460 -1170 39540 -1140
rect 39460 -1210 39480 -1170
rect 39520 -1210 39540 -1170
rect 39460 -1270 39540 -1210
rect 39460 -1310 39480 -1270
rect 39520 -1310 39540 -1270
rect 39460 -1340 39540 -1310
rect 39570 -1170 39650 -1140
rect 39570 -1210 39590 -1170
rect 39630 -1210 39650 -1170
rect 39570 -1270 39650 -1210
rect 39570 -1310 39590 -1270
rect 39630 -1310 39650 -1270
rect 39570 -1340 39650 -1310
rect 39680 -1170 39760 -1140
rect 39680 -1210 39700 -1170
rect 39740 -1210 39760 -1170
rect 39680 -1270 39760 -1210
rect 39680 -1310 39700 -1270
rect 39740 -1310 39760 -1270
rect 39680 -1340 39760 -1310
rect 39790 -1170 39870 -1140
rect 39790 -1210 39810 -1170
rect 39850 -1210 39870 -1170
rect 39790 -1270 39870 -1210
rect 39790 -1310 39810 -1270
rect 39850 -1310 39870 -1270
rect 39790 -1340 39870 -1310
rect 39900 -1170 39980 -1140
rect 39900 -1210 39920 -1170
rect 39960 -1210 39980 -1170
rect 39900 -1270 39980 -1210
rect 39900 -1310 39920 -1270
rect 39960 -1310 39980 -1270
rect 39900 -1340 39980 -1310
<< pdiff >>
rect 6070 6930 6150 6960
rect 6070 6786 6090 6930
rect 6130 6786 6150 6930
rect 6070 6760 6150 6786
rect 6180 6930 6260 6960
rect 6180 6786 6200 6930
rect 6240 6786 6260 6930
rect 6180 6760 6260 6786
rect 6290 6930 6370 6960
rect 6290 6786 6310 6930
rect 6350 6786 6370 6930
rect 6290 6760 6370 6786
rect 6400 6930 6480 6960
rect 6400 6786 6420 6930
rect 6460 6786 6480 6930
rect 6400 6760 6480 6786
rect 6510 6930 6590 6960
rect 6510 6786 6530 6930
rect 6570 6786 6590 6930
rect 6510 6760 6590 6786
rect 6620 6930 6700 6960
rect 6620 6786 6640 6930
rect 6680 6786 6700 6930
rect 6620 6760 6700 6786
rect 6730 6930 6810 6960
rect 6730 6786 6750 6930
rect 6790 6786 6810 6930
rect 6730 6760 6810 6786
rect 7350 6930 7430 6960
rect 7350 6890 7370 6930
rect 7410 6890 7430 6930
rect 7350 6830 7430 6890
rect 7350 6790 7370 6830
rect 7410 6790 7430 6830
rect 7350 6760 7430 6790
rect 7460 6930 7540 6960
rect 7460 6890 7480 6930
rect 7520 6890 7540 6930
rect 7460 6830 7540 6890
rect 7460 6790 7480 6830
rect 7520 6790 7540 6830
rect 7460 6760 7540 6790
rect 7570 6930 7650 6960
rect 7570 6890 7590 6930
rect 7630 6890 7650 6930
rect 7570 6830 7650 6890
rect 7570 6790 7590 6830
rect 7630 6790 7650 6830
rect 7570 6760 7650 6790
rect 7680 6930 7760 6960
rect 7680 6890 7700 6930
rect 7740 6890 7760 6930
rect 7680 6830 7760 6890
rect 7680 6790 7700 6830
rect 7740 6790 7760 6830
rect 7680 6760 7760 6790
rect 7790 6930 7870 6960
rect 7790 6890 7810 6930
rect 7850 6890 7870 6930
rect 7790 6830 7870 6890
rect 7790 6790 7810 6830
rect 7850 6790 7870 6830
rect 7790 6760 7870 6790
rect 7900 6930 7980 6960
rect 7900 6890 7920 6930
rect 7960 6890 7980 6930
rect 7900 6830 7980 6890
rect 7900 6790 7920 6830
rect 7960 6790 7980 6830
rect 7900 6760 7980 6790
rect 8010 6930 8090 6960
rect 8010 6890 8030 6930
rect 8070 6890 8090 6930
rect 8010 6830 8090 6890
rect 8010 6790 8030 6830
rect 8070 6790 8090 6830
rect 8010 6760 8090 6790
rect 8120 6930 8200 6960
rect 8120 6890 8140 6930
rect 8180 6890 8200 6930
rect 8120 6830 8200 6890
rect 8120 6790 8140 6830
rect 8180 6790 8200 6830
rect 8120 6760 8200 6790
rect 8230 6930 8310 6960
rect 8230 6890 8250 6930
rect 8290 6890 8310 6930
rect 8230 6830 8310 6890
rect 8230 6790 8250 6830
rect 8290 6790 8310 6830
rect 8230 6760 8310 6790
rect 8340 6930 8420 6960
rect 8340 6890 8360 6930
rect 8400 6890 8420 6930
rect 8340 6830 8420 6890
rect 8340 6790 8360 6830
rect 8400 6790 8420 6830
rect 8340 6760 8420 6790
rect 8450 6930 8530 6960
rect 8450 6890 8470 6930
rect 8510 6890 8530 6930
rect 8450 6830 8530 6890
rect 8450 6790 8470 6830
rect 8510 6790 8530 6830
rect 8450 6760 8530 6790
rect 8560 6930 8640 6960
rect 8560 6890 8580 6930
rect 8620 6890 8640 6930
rect 8560 6830 8640 6890
rect 8560 6790 8580 6830
rect 8620 6790 8640 6830
rect 8560 6760 8640 6790
rect 8670 6930 8750 6960
rect 8670 6890 8690 6930
rect 8730 6890 8750 6930
rect 8670 6830 8750 6890
rect 8670 6790 8690 6830
rect 8730 6790 8750 6830
rect 8670 6760 8750 6790
rect 9510 6930 9590 6960
rect 9510 6790 9530 6930
rect 9570 6790 9590 6930
rect 9510 6760 9590 6790
rect 9620 6930 9700 6960
rect 9620 6790 9640 6930
rect 9680 6790 9700 6930
rect 9620 6760 9700 6790
rect 9730 6930 9810 6960
rect 9730 6790 9750 6930
rect 9790 6790 9810 6930
rect 9730 6760 9810 6790
rect 9840 6930 9920 6960
rect 9840 6790 9860 6930
rect 9900 6790 9920 6930
rect 9840 6760 9920 6790
rect 9950 6930 10030 6960
rect 9950 6790 9970 6930
rect 10010 6790 10030 6930
rect 9950 6760 10030 6790
rect 10060 6930 10140 6960
rect 10060 6790 10080 6930
rect 10120 6790 10140 6930
rect 10060 6760 10140 6790
rect 10170 6930 10250 6960
rect 10170 6790 10190 6930
rect 10230 6790 10250 6930
rect 10170 6760 10250 6790
rect 5430 5800 5510 5830
rect 5430 5760 5450 5800
rect 5490 5760 5510 5800
rect 5430 5700 5510 5760
rect 5430 5660 5450 5700
rect 5490 5660 5510 5700
rect 5430 5630 5510 5660
rect 5540 5800 5620 5830
rect 5540 5760 5560 5800
rect 5600 5760 5620 5800
rect 5540 5700 5620 5760
rect 5540 5660 5560 5700
rect 5600 5660 5620 5700
rect 5540 5630 5620 5660
rect 5650 5800 5730 5830
rect 5650 5760 5670 5800
rect 5710 5760 5730 5800
rect 5650 5700 5730 5760
rect 5650 5660 5670 5700
rect 5710 5660 5730 5700
rect 5650 5630 5730 5660
rect 5760 5800 5840 5830
rect 5760 5760 5780 5800
rect 5820 5760 5840 5800
rect 5760 5700 5840 5760
rect 5760 5660 5780 5700
rect 5820 5660 5840 5700
rect 5760 5630 5840 5660
rect 5870 5800 5950 5830
rect 5870 5760 5890 5800
rect 5930 5760 5950 5800
rect 5870 5700 5950 5760
rect 5870 5660 5890 5700
rect 5930 5660 5950 5700
rect 5870 5630 5950 5660
rect 6500 6000 6580 6030
rect 6500 5960 6520 6000
rect 6560 5960 6580 6000
rect 6500 5900 6580 5960
rect 6500 5860 6520 5900
rect 6560 5860 6580 5900
rect 6500 5800 6580 5860
rect 6500 5760 6520 5800
rect 6560 5760 6580 5800
rect 6500 5700 6580 5760
rect 6500 5660 6520 5700
rect 6560 5660 6580 5700
rect 6500 5600 6580 5660
rect 6500 5560 6520 5600
rect 6560 5560 6580 5600
rect 6500 5500 6580 5560
rect 6500 5460 6520 5500
rect 6560 5460 6580 5500
rect 6500 5430 6580 5460
rect 6680 6000 6760 6030
rect 6680 5960 6700 6000
rect 6740 5960 6760 6000
rect 6680 5900 6760 5960
rect 6680 5860 6700 5900
rect 6740 5860 6760 5900
rect 6680 5800 6760 5860
rect 6680 5760 6700 5800
rect 6740 5760 6760 5800
rect 6680 5700 6760 5760
rect 6680 5660 6700 5700
rect 6740 5660 6760 5700
rect 6680 5600 6760 5660
rect 6680 5560 6700 5600
rect 6740 5560 6760 5600
rect 6680 5500 6760 5560
rect 6680 5460 6700 5500
rect 6740 5460 6760 5500
rect 6680 5430 6760 5460
rect 6860 6000 6940 6030
rect 6860 5960 6880 6000
rect 6920 5960 6940 6000
rect 6860 5900 6940 5960
rect 6860 5860 6880 5900
rect 6920 5860 6940 5900
rect 6860 5800 6940 5860
rect 6860 5760 6880 5800
rect 6920 5760 6940 5800
rect 6860 5700 6940 5760
rect 6860 5660 6880 5700
rect 6920 5660 6940 5700
rect 6860 5600 6940 5660
rect 6860 5560 6880 5600
rect 6920 5560 6940 5600
rect 6860 5500 6940 5560
rect 6860 5460 6880 5500
rect 6920 5460 6940 5500
rect 6860 5430 6940 5460
rect 7040 6000 7120 6030
rect 7040 5960 7060 6000
rect 7100 5960 7120 6000
rect 7040 5900 7120 5960
rect 7040 5860 7060 5900
rect 7100 5860 7120 5900
rect 7040 5800 7120 5860
rect 7040 5760 7060 5800
rect 7100 5760 7120 5800
rect 7040 5700 7120 5760
rect 7040 5660 7060 5700
rect 7100 5660 7120 5700
rect 7040 5600 7120 5660
rect 7040 5560 7060 5600
rect 7100 5560 7120 5600
rect 7040 5500 7120 5560
rect 7040 5460 7060 5500
rect 7100 5460 7120 5500
rect 7040 5430 7120 5460
rect 7220 6000 7300 6030
rect 7220 5960 7240 6000
rect 7280 5960 7300 6000
rect 7220 5900 7300 5960
rect 7220 5860 7240 5900
rect 7280 5860 7300 5900
rect 7220 5800 7300 5860
rect 7220 5760 7240 5800
rect 7280 5760 7300 5800
rect 7220 5700 7300 5760
rect 7220 5660 7240 5700
rect 7280 5660 7300 5700
rect 7220 5600 7300 5660
rect 7220 5560 7240 5600
rect 7280 5560 7300 5600
rect 7220 5500 7300 5560
rect 7220 5460 7240 5500
rect 7280 5460 7300 5500
rect 7220 5430 7300 5460
rect 7400 6000 7480 6030
rect 7400 5960 7420 6000
rect 7460 5960 7480 6000
rect 7400 5900 7480 5960
rect 7400 5860 7420 5900
rect 7460 5860 7480 5900
rect 7400 5800 7480 5860
rect 7400 5760 7420 5800
rect 7460 5760 7480 5800
rect 7400 5700 7480 5760
rect 7400 5660 7420 5700
rect 7460 5660 7480 5700
rect 7400 5600 7480 5660
rect 7400 5560 7420 5600
rect 7460 5560 7480 5600
rect 7400 5500 7480 5560
rect 7400 5460 7420 5500
rect 7460 5460 7480 5500
rect 7400 5430 7480 5460
rect 7580 6000 7660 6030
rect 7580 5960 7600 6000
rect 7640 5960 7660 6000
rect 7580 5900 7660 5960
rect 7580 5860 7600 5900
rect 7640 5860 7660 5900
rect 7580 5800 7660 5860
rect 7580 5760 7600 5800
rect 7640 5760 7660 5800
rect 7580 5700 7660 5760
rect 7580 5660 7600 5700
rect 7640 5660 7660 5700
rect 7580 5600 7660 5660
rect 7580 5560 7600 5600
rect 7640 5560 7660 5600
rect 7580 5500 7660 5560
rect 7580 5460 7600 5500
rect 7640 5460 7660 5500
rect 7580 5430 7660 5460
rect 7760 6000 7840 6030
rect 7760 5960 7780 6000
rect 7820 5960 7840 6000
rect 7760 5900 7840 5960
rect 7760 5860 7780 5900
rect 7820 5860 7840 5900
rect 7760 5800 7840 5860
rect 7760 5760 7780 5800
rect 7820 5760 7840 5800
rect 7760 5700 7840 5760
rect 7760 5660 7780 5700
rect 7820 5660 7840 5700
rect 7760 5600 7840 5660
rect 7760 5560 7780 5600
rect 7820 5560 7840 5600
rect 7760 5500 7840 5560
rect 7760 5460 7780 5500
rect 7820 5460 7840 5500
rect 7760 5430 7840 5460
rect 7940 6000 8020 6030
rect 7940 5960 7960 6000
rect 8000 5960 8020 6000
rect 7940 5900 8020 5960
rect 7940 5860 7960 5900
rect 8000 5860 8020 5900
rect 7940 5800 8020 5860
rect 7940 5760 7960 5800
rect 8000 5760 8020 5800
rect 7940 5700 8020 5760
rect 7940 5660 7960 5700
rect 8000 5660 8020 5700
rect 7940 5600 8020 5660
rect 7940 5560 7960 5600
rect 8000 5560 8020 5600
rect 7940 5500 8020 5560
rect 7940 5460 7960 5500
rect 8000 5460 8020 5500
rect 7940 5430 8020 5460
rect 8120 6000 8200 6030
rect 8120 5960 8140 6000
rect 8180 5960 8200 6000
rect 8120 5900 8200 5960
rect 8120 5860 8140 5900
rect 8180 5860 8200 5900
rect 8120 5800 8200 5860
rect 8120 5760 8140 5800
rect 8180 5760 8200 5800
rect 8120 5700 8200 5760
rect 8120 5660 8140 5700
rect 8180 5660 8200 5700
rect 8120 5600 8200 5660
rect 8120 5560 8140 5600
rect 8180 5560 8200 5600
rect 8120 5500 8200 5560
rect 8120 5460 8140 5500
rect 8180 5460 8200 5500
rect 8120 5430 8200 5460
rect 8300 6000 8380 6030
rect 8300 5960 8320 6000
rect 8360 5960 8380 6000
rect 8300 5900 8380 5960
rect 8300 5860 8320 5900
rect 8360 5860 8380 5900
rect 8300 5800 8380 5860
rect 8300 5760 8320 5800
rect 8360 5760 8380 5800
rect 8300 5700 8380 5760
rect 8300 5660 8320 5700
rect 8360 5660 8380 5700
rect 8300 5600 8380 5660
rect 8300 5560 8320 5600
rect 8360 5560 8380 5600
rect 8300 5500 8380 5560
rect 8300 5460 8320 5500
rect 8360 5460 8380 5500
rect 8300 5430 8380 5460
rect 8480 6000 8560 6030
rect 8480 5960 8500 6000
rect 8540 5960 8560 6000
rect 8480 5900 8560 5960
rect 8480 5860 8500 5900
rect 8540 5860 8560 5900
rect 8480 5800 8560 5860
rect 8480 5760 8500 5800
rect 8540 5760 8560 5800
rect 8480 5700 8560 5760
rect 8480 5660 8500 5700
rect 8540 5660 8560 5700
rect 8480 5600 8560 5660
rect 8480 5560 8500 5600
rect 8540 5560 8560 5600
rect 8480 5500 8560 5560
rect 8480 5460 8500 5500
rect 8540 5460 8560 5500
rect 8480 5430 8560 5460
rect 8660 6000 8740 6030
rect 8660 5960 8680 6000
rect 8720 5960 8740 6000
rect 8660 5900 8740 5960
rect 8660 5860 8680 5900
rect 8720 5860 8740 5900
rect 8660 5800 8740 5860
rect 8660 5760 8680 5800
rect 8720 5760 8740 5800
rect 8660 5700 8740 5760
rect 8660 5660 8680 5700
rect 8720 5660 8740 5700
rect 8660 5600 8740 5660
rect 8660 5560 8680 5600
rect 8720 5560 8740 5600
rect 8660 5500 8740 5560
rect 8660 5460 8680 5500
rect 8720 5460 8740 5500
rect 8660 5430 8740 5460
rect 8840 6000 8920 6030
rect 8840 5960 8860 6000
rect 8900 5960 8920 6000
rect 8840 5900 8920 5960
rect 8840 5860 8860 5900
rect 8900 5860 8920 5900
rect 8840 5800 8920 5860
rect 8840 5760 8860 5800
rect 8900 5760 8920 5800
rect 8840 5700 8920 5760
rect 8840 5660 8860 5700
rect 8900 5660 8920 5700
rect 8840 5600 8920 5660
rect 8840 5560 8860 5600
rect 8900 5560 8920 5600
rect 8840 5500 8920 5560
rect 8840 5460 8860 5500
rect 8900 5460 8920 5500
rect 8840 5430 8920 5460
rect 9020 6000 9100 6030
rect 9020 5960 9040 6000
rect 9080 5960 9100 6000
rect 9020 5900 9100 5960
rect 9020 5860 9040 5900
rect 9080 5860 9100 5900
rect 9020 5800 9100 5860
rect 9020 5760 9040 5800
rect 9080 5760 9100 5800
rect 9020 5700 9100 5760
rect 9020 5660 9040 5700
rect 9080 5660 9100 5700
rect 9020 5600 9100 5660
rect 9020 5560 9040 5600
rect 9080 5560 9100 5600
rect 9020 5500 9100 5560
rect 9020 5460 9040 5500
rect 9080 5460 9100 5500
rect 9020 5430 9100 5460
rect 9200 6000 9280 6030
rect 9200 5960 9220 6000
rect 9260 5960 9280 6000
rect 9200 5900 9280 5960
rect 9200 5860 9220 5900
rect 9260 5860 9280 5900
rect 9200 5800 9280 5860
rect 9200 5760 9220 5800
rect 9260 5760 9280 5800
rect 9200 5700 9280 5760
rect 9200 5660 9220 5700
rect 9260 5660 9280 5700
rect 9200 5600 9280 5660
rect 9200 5560 9220 5600
rect 9260 5560 9280 5600
rect 9200 5500 9280 5560
rect 9200 5460 9220 5500
rect 9260 5460 9280 5500
rect 9200 5430 9280 5460
rect 9380 6000 9460 6030
rect 9380 5960 9400 6000
rect 9440 5960 9460 6000
rect 9380 5900 9460 5960
rect 9380 5860 9400 5900
rect 9440 5860 9460 5900
rect 9380 5800 9460 5860
rect 9380 5760 9400 5800
rect 9440 5760 9460 5800
rect 9380 5700 9460 5760
rect 9380 5660 9400 5700
rect 9440 5660 9460 5700
rect 9380 5600 9460 5660
rect 9380 5560 9400 5600
rect 9440 5560 9460 5600
rect 9380 5500 9460 5560
rect 9380 5460 9400 5500
rect 9440 5460 9460 5500
rect 9380 5430 9460 5460
rect 9560 6000 9640 6030
rect 9560 5960 9580 6000
rect 9620 5960 9640 6000
rect 9560 5900 9640 5960
rect 9560 5860 9580 5900
rect 9620 5860 9640 5900
rect 9560 5800 9640 5860
rect 9560 5760 9580 5800
rect 9620 5760 9640 5800
rect 9560 5700 9640 5760
rect 9560 5660 9580 5700
rect 9620 5660 9640 5700
rect 9560 5600 9640 5660
rect 9560 5560 9580 5600
rect 9620 5560 9640 5600
rect 9560 5500 9640 5560
rect 9560 5460 9580 5500
rect 9620 5460 9640 5500
rect 9560 5430 9640 5460
rect 9740 6000 9820 6030
rect 9740 5960 9760 6000
rect 9800 5960 9820 6000
rect 9740 5900 9820 5960
rect 9740 5860 9760 5900
rect 9800 5860 9820 5900
rect 9740 5800 9820 5860
rect 9740 5760 9760 5800
rect 9800 5760 9820 5800
rect 9740 5700 9820 5760
rect 9740 5660 9760 5700
rect 9800 5660 9820 5700
rect 9740 5600 9820 5660
rect 9740 5560 9760 5600
rect 9800 5560 9820 5600
rect 9740 5500 9820 5560
rect 9740 5460 9760 5500
rect 9800 5460 9820 5500
rect 9740 5430 9820 5460
rect 10360 5800 10440 5830
rect 10360 5760 10380 5800
rect 10420 5760 10440 5800
rect 10360 5700 10440 5760
rect 10360 5660 10380 5700
rect 10420 5660 10440 5700
rect 10360 5630 10440 5660
rect 10470 5800 10550 5830
rect 10470 5760 10490 5800
rect 10530 5760 10550 5800
rect 10470 5700 10550 5760
rect 10470 5660 10490 5700
rect 10530 5660 10550 5700
rect 10470 5630 10550 5660
rect 10580 5800 10660 5830
rect 10580 5760 10600 5800
rect 10640 5760 10660 5800
rect 10580 5700 10660 5760
rect 10580 5660 10600 5700
rect 10640 5660 10660 5700
rect 10580 5630 10660 5660
rect 10690 5800 10770 5830
rect 10690 5760 10710 5800
rect 10750 5760 10770 5800
rect 10690 5700 10770 5760
rect 10690 5660 10710 5700
rect 10750 5660 10770 5700
rect 10690 5630 10770 5660
rect 10800 5800 10880 5830
rect 10800 5760 10820 5800
rect 10860 5760 10880 5800
rect 10800 5700 10880 5760
rect 10800 5660 10820 5700
rect 10860 5660 10880 5700
rect 10800 5630 10880 5660
rect 5400 4620 5480 4650
rect 5400 4580 5420 4620
rect 5460 4580 5480 4620
rect 5400 4520 5480 4580
rect 5400 4480 5420 4520
rect 5460 4480 5480 4520
rect 5400 4450 5480 4480
rect 5520 4620 5600 4650
rect 5520 4580 5540 4620
rect 5580 4580 5600 4620
rect 5520 4520 5600 4580
rect 5520 4480 5540 4520
rect 5580 4480 5600 4520
rect 5520 4450 5600 4480
rect 5640 4620 5720 4650
rect 5640 4580 5660 4620
rect 5700 4580 5720 4620
rect 5640 4520 5720 4580
rect 5640 4480 5660 4520
rect 5700 4480 5720 4520
rect 5640 4450 5720 4480
rect 5760 4620 5840 4650
rect 5760 4580 5780 4620
rect 5820 4580 5840 4620
rect 5760 4520 5840 4580
rect 5760 4480 5780 4520
rect 5820 4480 5840 4520
rect 5760 4450 5840 4480
rect 5880 4620 5960 4650
rect 5880 4580 5900 4620
rect 5940 4580 5960 4620
rect 5880 4520 5960 4580
rect 5880 4480 5900 4520
rect 5940 4480 5960 4520
rect 5880 4450 5960 4480
rect 6000 4620 6080 4650
rect 6000 4580 6020 4620
rect 6060 4580 6080 4620
rect 6000 4520 6080 4580
rect 6000 4480 6020 4520
rect 6060 4480 6080 4520
rect 6000 4450 6080 4480
rect 6120 4620 6200 4650
rect 6120 4580 6140 4620
rect 6180 4580 6200 4620
rect 6120 4520 6200 4580
rect 6120 4480 6140 4520
rect 6180 4480 6200 4520
rect 6120 4450 6200 4480
rect 6240 4620 6320 4650
rect 6240 4580 6260 4620
rect 6300 4580 6320 4620
rect 6240 4520 6320 4580
rect 6240 4480 6260 4520
rect 6300 4480 6320 4520
rect 6240 4450 6320 4480
rect 6360 4620 6440 4650
rect 6360 4580 6380 4620
rect 6420 4580 6440 4620
rect 6360 4520 6440 4580
rect 6360 4480 6380 4520
rect 6420 4480 6440 4520
rect 6360 4450 6440 4480
rect 6480 4620 6560 4650
rect 6480 4580 6500 4620
rect 6540 4580 6560 4620
rect 6480 4520 6560 4580
rect 6480 4480 6500 4520
rect 6540 4480 6560 4520
rect 6480 4450 6560 4480
rect 6600 4620 6680 4650
rect 6600 4580 6620 4620
rect 6660 4580 6680 4620
rect 6600 4520 6680 4580
rect 6600 4480 6620 4520
rect 6660 4480 6680 4520
rect 6600 4450 6680 4480
rect 6720 4620 6800 4650
rect 6720 4580 6740 4620
rect 6780 4580 6800 4620
rect 6720 4520 6800 4580
rect 6720 4480 6740 4520
rect 6780 4480 6800 4520
rect 6720 4450 6800 4480
rect 6840 4620 6920 4650
rect 6840 4580 6860 4620
rect 6900 4580 6920 4620
rect 6840 4520 6920 4580
rect 6840 4480 6860 4520
rect 6900 4480 6920 4520
rect 6840 4450 6920 4480
rect 6960 4620 7040 4650
rect 6960 4580 6980 4620
rect 7020 4580 7040 4620
rect 6960 4520 7040 4580
rect 6960 4480 6980 4520
rect 7020 4480 7040 4520
rect 6960 4450 7040 4480
rect 7080 4620 7160 4650
rect 7080 4580 7100 4620
rect 7140 4580 7160 4620
rect 7080 4520 7160 4580
rect 7080 4480 7100 4520
rect 7140 4480 7160 4520
rect 7080 4450 7160 4480
rect 7200 4620 7280 4650
rect 7200 4580 7220 4620
rect 7260 4580 7280 4620
rect 7200 4520 7280 4580
rect 7200 4480 7220 4520
rect 7260 4480 7280 4520
rect 7200 4450 7280 4480
rect 7320 4620 7400 4650
rect 7320 4580 7340 4620
rect 7380 4580 7400 4620
rect 7320 4520 7400 4580
rect 7320 4480 7340 4520
rect 7380 4480 7400 4520
rect 7320 4450 7400 4480
rect 7440 4620 7520 4650
rect 7440 4580 7460 4620
rect 7500 4580 7520 4620
rect 7440 4520 7520 4580
rect 7440 4480 7460 4520
rect 7500 4480 7520 4520
rect 7440 4450 7520 4480
rect 7560 4620 7640 4650
rect 7560 4580 7580 4620
rect 7620 4580 7640 4620
rect 7560 4520 7640 4580
rect 7560 4480 7580 4520
rect 7620 4480 7640 4520
rect 7560 4450 7640 4480
rect 7680 4620 7760 4650
rect 7680 4580 7700 4620
rect 7740 4580 7760 4620
rect 7680 4520 7760 4580
rect 7680 4480 7700 4520
rect 7740 4480 7760 4520
rect 7680 4450 7760 4480
rect 7800 4620 7880 4650
rect 7800 4580 7820 4620
rect 7860 4580 7880 4620
rect 7800 4520 7880 4580
rect 7800 4480 7820 4520
rect 7860 4480 7880 4520
rect 7800 4450 7880 4480
rect 8440 4620 8520 4650
rect 8440 4580 8460 4620
rect 8500 4580 8520 4620
rect 8440 4520 8520 4580
rect 8440 4480 8460 4520
rect 8500 4480 8520 4520
rect 8440 4450 8520 4480
rect 8560 4620 8640 4650
rect 8560 4580 8580 4620
rect 8620 4580 8640 4620
rect 8560 4520 8640 4580
rect 8560 4480 8580 4520
rect 8620 4480 8640 4520
rect 8560 4450 8640 4480
rect 8680 4620 8760 4650
rect 8680 4580 8700 4620
rect 8740 4580 8760 4620
rect 8680 4520 8760 4580
rect 8680 4480 8700 4520
rect 8740 4480 8760 4520
rect 8680 4450 8760 4480
rect 8800 4620 8880 4650
rect 8800 4580 8820 4620
rect 8860 4580 8880 4620
rect 8800 4520 8880 4580
rect 8800 4480 8820 4520
rect 8860 4480 8880 4520
rect 8800 4450 8880 4480
rect 8920 4620 9000 4650
rect 8920 4580 8940 4620
rect 8980 4580 9000 4620
rect 8920 4520 9000 4580
rect 8920 4480 8940 4520
rect 8980 4480 9000 4520
rect 8920 4450 9000 4480
rect 9040 4620 9120 4650
rect 9040 4580 9060 4620
rect 9100 4580 9120 4620
rect 9040 4520 9120 4580
rect 9040 4480 9060 4520
rect 9100 4480 9120 4520
rect 9040 4450 9120 4480
rect 9160 4620 9240 4650
rect 9160 4580 9180 4620
rect 9220 4580 9240 4620
rect 9160 4520 9240 4580
rect 9160 4480 9180 4520
rect 9220 4480 9240 4520
rect 9160 4450 9240 4480
rect 9280 4620 9360 4650
rect 9280 4580 9300 4620
rect 9340 4580 9360 4620
rect 9280 4520 9360 4580
rect 9280 4480 9300 4520
rect 9340 4480 9360 4520
rect 9280 4450 9360 4480
rect 9400 4620 9480 4650
rect 9400 4580 9420 4620
rect 9460 4580 9480 4620
rect 9400 4520 9480 4580
rect 9400 4480 9420 4520
rect 9460 4480 9480 4520
rect 9400 4450 9480 4480
rect 9520 4620 9600 4650
rect 9520 4580 9540 4620
rect 9580 4580 9600 4620
rect 9520 4520 9600 4580
rect 9520 4480 9540 4520
rect 9580 4480 9600 4520
rect 9520 4450 9600 4480
rect 9640 4620 9720 4650
rect 9640 4580 9660 4620
rect 9700 4580 9720 4620
rect 9640 4520 9720 4580
rect 9640 4480 9660 4520
rect 9700 4480 9720 4520
rect 9640 4450 9720 4480
rect 9760 4620 9840 4650
rect 9760 4580 9780 4620
rect 9820 4580 9840 4620
rect 9760 4520 9840 4580
rect 9760 4480 9780 4520
rect 9820 4480 9840 4520
rect 9760 4450 9840 4480
rect 9880 4620 9960 4650
rect 9880 4580 9900 4620
rect 9940 4580 9960 4620
rect 9880 4520 9960 4580
rect 9880 4480 9900 4520
rect 9940 4480 9960 4520
rect 9880 4450 9960 4480
rect 10000 4620 10080 4650
rect 10000 4580 10020 4620
rect 10060 4580 10080 4620
rect 10000 4520 10080 4580
rect 10000 4480 10020 4520
rect 10060 4480 10080 4520
rect 10000 4450 10080 4480
rect 10120 4620 10200 4650
rect 10120 4580 10140 4620
rect 10180 4580 10200 4620
rect 10120 4520 10200 4580
rect 10120 4480 10140 4520
rect 10180 4480 10200 4520
rect 10120 4450 10200 4480
rect 10240 4620 10320 4650
rect 10240 4580 10260 4620
rect 10300 4580 10320 4620
rect 10240 4520 10320 4580
rect 10240 4480 10260 4520
rect 10300 4480 10320 4520
rect 10240 4450 10320 4480
rect 10360 4620 10440 4650
rect 10360 4580 10380 4620
rect 10420 4580 10440 4620
rect 10360 4520 10440 4580
rect 10360 4480 10380 4520
rect 10420 4480 10440 4520
rect 10360 4450 10440 4480
rect 10480 4620 10560 4650
rect 10480 4580 10500 4620
rect 10540 4580 10560 4620
rect 10480 4520 10560 4580
rect 10480 4480 10500 4520
rect 10540 4480 10560 4520
rect 10480 4450 10560 4480
rect 10600 4620 10680 4650
rect 10600 4580 10620 4620
rect 10660 4580 10680 4620
rect 10600 4520 10680 4580
rect 10600 4480 10620 4520
rect 10660 4480 10680 4520
rect 10600 4450 10680 4480
rect 10720 4620 10800 4650
rect 10720 4580 10740 4620
rect 10780 4580 10800 4620
rect 10720 4520 10800 4580
rect 10720 4480 10740 4520
rect 10780 4480 10800 4520
rect 10720 4450 10800 4480
rect 10840 4620 10920 4650
rect 10840 4580 10860 4620
rect 10900 4580 10920 4620
rect 10840 4520 10920 4580
rect 10840 4480 10860 4520
rect 10900 4480 10920 4520
rect 10840 4450 10920 4480
rect 36070 3930 36150 3960
rect 36070 3786 36090 3930
rect 36130 3786 36150 3930
rect 36070 3760 36150 3786
rect 36180 3930 36260 3960
rect 36180 3786 36200 3930
rect 36240 3786 36260 3930
rect 36180 3760 36260 3786
rect 36290 3930 36370 3960
rect 36290 3786 36310 3930
rect 36350 3786 36370 3930
rect 36290 3760 36370 3786
rect 36400 3930 36480 3960
rect 36400 3786 36420 3930
rect 36460 3786 36480 3930
rect 36400 3760 36480 3786
rect 36510 3930 36590 3960
rect 36510 3786 36530 3930
rect 36570 3786 36590 3930
rect 36510 3760 36590 3786
rect 36620 3930 36700 3960
rect 36620 3786 36640 3930
rect 36680 3786 36700 3930
rect 36620 3760 36700 3786
rect 36730 3930 36810 3960
rect 36730 3786 36750 3930
rect 36790 3786 36810 3930
rect 36730 3760 36810 3786
rect 37350 3930 37430 3960
rect 37350 3890 37370 3930
rect 37410 3890 37430 3930
rect 37350 3830 37430 3890
rect 37350 3790 37370 3830
rect 37410 3790 37430 3830
rect 37350 3760 37430 3790
rect 37460 3930 37540 3960
rect 37460 3890 37480 3930
rect 37520 3890 37540 3930
rect 37460 3830 37540 3890
rect 37460 3790 37480 3830
rect 37520 3790 37540 3830
rect 37460 3760 37540 3790
rect 37570 3930 37650 3960
rect 37570 3890 37590 3930
rect 37630 3890 37650 3930
rect 37570 3830 37650 3890
rect 37570 3790 37590 3830
rect 37630 3790 37650 3830
rect 37570 3760 37650 3790
rect 37680 3930 37760 3960
rect 37680 3890 37700 3930
rect 37740 3890 37760 3930
rect 37680 3830 37760 3890
rect 37680 3790 37700 3830
rect 37740 3790 37760 3830
rect 37680 3760 37760 3790
rect 37790 3930 37870 3960
rect 37790 3890 37810 3930
rect 37850 3890 37870 3930
rect 37790 3830 37870 3890
rect 37790 3790 37810 3830
rect 37850 3790 37870 3830
rect 37790 3760 37870 3790
rect 37900 3930 37980 3960
rect 37900 3890 37920 3930
rect 37960 3890 37980 3930
rect 37900 3830 37980 3890
rect 37900 3790 37920 3830
rect 37960 3790 37980 3830
rect 37900 3760 37980 3790
rect 38010 3930 38090 3960
rect 38010 3890 38030 3930
rect 38070 3890 38090 3930
rect 38010 3830 38090 3890
rect 38010 3790 38030 3830
rect 38070 3790 38090 3830
rect 38010 3760 38090 3790
rect 38120 3930 38200 3960
rect 38120 3890 38140 3930
rect 38180 3890 38200 3930
rect 38120 3830 38200 3890
rect 38120 3790 38140 3830
rect 38180 3790 38200 3830
rect 38120 3760 38200 3790
rect 38230 3930 38310 3960
rect 38230 3890 38250 3930
rect 38290 3890 38310 3930
rect 38230 3830 38310 3890
rect 38230 3790 38250 3830
rect 38290 3790 38310 3830
rect 38230 3760 38310 3790
rect 38340 3930 38420 3960
rect 38340 3890 38360 3930
rect 38400 3890 38420 3930
rect 38340 3830 38420 3890
rect 38340 3790 38360 3830
rect 38400 3790 38420 3830
rect 38340 3760 38420 3790
rect 38450 3930 38530 3960
rect 38450 3890 38470 3930
rect 38510 3890 38530 3930
rect 38450 3830 38530 3890
rect 38450 3790 38470 3830
rect 38510 3790 38530 3830
rect 38450 3760 38530 3790
rect 38560 3930 38640 3960
rect 38560 3890 38580 3930
rect 38620 3890 38640 3930
rect 38560 3830 38640 3890
rect 38560 3790 38580 3830
rect 38620 3790 38640 3830
rect 38560 3760 38640 3790
rect 38670 3930 38750 3960
rect 38670 3890 38690 3930
rect 38730 3890 38750 3930
rect 38670 3830 38750 3890
rect 38670 3790 38690 3830
rect 38730 3790 38750 3830
rect 38670 3760 38750 3790
rect 39510 3930 39590 3960
rect 39510 3790 39530 3930
rect 39570 3790 39590 3930
rect 39510 3760 39590 3790
rect 39620 3930 39700 3960
rect 39620 3790 39640 3930
rect 39680 3790 39700 3930
rect 39620 3760 39700 3790
rect 39730 3930 39810 3960
rect 39730 3790 39750 3930
rect 39790 3790 39810 3930
rect 39730 3760 39810 3790
rect 39840 3930 39920 3960
rect 39840 3790 39860 3930
rect 39900 3790 39920 3930
rect 39840 3760 39920 3790
rect 39950 3930 40030 3960
rect 39950 3790 39970 3930
rect 40010 3790 40030 3930
rect 39950 3760 40030 3790
rect 40060 3930 40140 3960
rect 40060 3790 40080 3930
rect 40120 3790 40140 3930
rect 40060 3760 40140 3790
rect 40170 3930 40250 3960
rect 40170 3790 40190 3930
rect 40230 3790 40250 3930
rect 40170 3760 40250 3790
rect 35430 2800 35510 2830
rect 35430 2760 35450 2800
rect 35490 2760 35510 2800
rect 35430 2700 35510 2760
rect 35430 2660 35450 2700
rect 35490 2660 35510 2700
rect 35430 2630 35510 2660
rect 35540 2800 35620 2830
rect 35540 2760 35560 2800
rect 35600 2760 35620 2800
rect 35540 2700 35620 2760
rect 35540 2660 35560 2700
rect 35600 2660 35620 2700
rect 35540 2630 35620 2660
rect 35650 2800 35730 2830
rect 35650 2760 35670 2800
rect 35710 2760 35730 2800
rect 35650 2700 35730 2760
rect 35650 2660 35670 2700
rect 35710 2660 35730 2700
rect 35650 2630 35730 2660
rect 35760 2800 35840 2830
rect 35760 2760 35780 2800
rect 35820 2760 35840 2800
rect 35760 2700 35840 2760
rect 35760 2660 35780 2700
rect 35820 2660 35840 2700
rect 35760 2630 35840 2660
rect 35870 2800 35950 2830
rect 35870 2760 35890 2800
rect 35930 2760 35950 2800
rect 35870 2700 35950 2760
rect 35870 2660 35890 2700
rect 35930 2660 35950 2700
rect 35870 2630 35950 2660
rect 36500 3000 36580 3030
rect 36500 2960 36520 3000
rect 36560 2960 36580 3000
rect 36500 2900 36580 2960
rect 36500 2860 36520 2900
rect 36560 2860 36580 2900
rect 36500 2800 36580 2860
rect 36500 2760 36520 2800
rect 36560 2760 36580 2800
rect 36500 2700 36580 2760
rect 36500 2660 36520 2700
rect 36560 2660 36580 2700
rect 36500 2600 36580 2660
rect 36500 2560 36520 2600
rect 36560 2560 36580 2600
rect 36500 2500 36580 2560
rect 36500 2460 36520 2500
rect 36560 2460 36580 2500
rect 36500 2430 36580 2460
rect 36680 3000 36760 3030
rect 36680 2960 36700 3000
rect 36740 2960 36760 3000
rect 36680 2900 36760 2960
rect 36680 2860 36700 2900
rect 36740 2860 36760 2900
rect 36680 2800 36760 2860
rect 36680 2760 36700 2800
rect 36740 2760 36760 2800
rect 36680 2700 36760 2760
rect 36680 2660 36700 2700
rect 36740 2660 36760 2700
rect 36680 2600 36760 2660
rect 36680 2560 36700 2600
rect 36740 2560 36760 2600
rect 36680 2500 36760 2560
rect 36680 2460 36700 2500
rect 36740 2460 36760 2500
rect 36680 2430 36760 2460
rect 36860 3000 36940 3030
rect 36860 2960 36880 3000
rect 36920 2960 36940 3000
rect 36860 2900 36940 2960
rect 36860 2860 36880 2900
rect 36920 2860 36940 2900
rect 36860 2800 36940 2860
rect 36860 2760 36880 2800
rect 36920 2760 36940 2800
rect 36860 2700 36940 2760
rect 36860 2660 36880 2700
rect 36920 2660 36940 2700
rect 36860 2600 36940 2660
rect 36860 2560 36880 2600
rect 36920 2560 36940 2600
rect 36860 2500 36940 2560
rect 36860 2460 36880 2500
rect 36920 2460 36940 2500
rect 36860 2430 36940 2460
rect 37040 3000 37120 3030
rect 37040 2960 37060 3000
rect 37100 2960 37120 3000
rect 37040 2900 37120 2960
rect 37040 2860 37060 2900
rect 37100 2860 37120 2900
rect 37040 2800 37120 2860
rect 37040 2760 37060 2800
rect 37100 2760 37120 2800
rect 37040 2700 37120 2760
rect 37040 2660 37060 2700
rect 37100 2660 37120 2700
rect 37040 2600 37120 2660
rect 37040 2560 37060 2600
rect 37100 2560 37120 2600
rect 37040 2500 37120 2560
rect 37040 2460 37060 2500
rect 37100 2460 37120 2500
rect 37040 2430 37120 2460
rect 37220 3000 37300 3030
rect 37220 2960 37240 3000
rect 37280 2960 37300 3000
rect 37220 2900 37300 2960
rect 37220 2860 37240 2900
rect 37280 2860 37300 2900
rect 37220 2800 37300 2860
rect 37220 2760 37240 2800
rect 37280 2760 37300 2800
rect 37220 2700 37300 2760
rect 37220 2660 37240 2700
rect 37280 2660 37300 2700
rect 37220 2600 37300 2660
rect 37220 2560 37240 2600
rect 37280 2560 37300 2600
rect 37220 2500 37300 2560
rect 37220 2460 37240 2500
rect 37280 2460 37300 2500
rect 37220 2430 37300 2460
rect 37400 3000 37480 3030
rect 37400 2960 37420 3000
rect 37460 2960 37480 3000
rect 37400 2900 37480 2960
rect 37400 2860 37420 2900
rect 37460 2860 37480 2900
rect 37400 2800 37480 2860
rect 37400 2760 37420 2800
rect 37460 2760 37480 2800
rect 37400 2700 37480 2760
rect 37400 2660 37420 2700
rect 37460 2660 37480 2700
rect 37400 2600 37480 2660
rect 37400 2560 37420 2600
rect 37460 2560 37480 2600
rect 37400 2500 37480 2560
rect 37400 2460 37420 2500
rect 37460 2460 37480 2500
rect 37400 2430 37480 2460
rect 37580 3000 37660 3030
rect 37580 2960 37600 3000
rect 37640 2960 37660 3000
rect 37580 2900 37660 2960
rect 37580 2860 37600 2900
rect 37640 2860 37660 2900
rect 37580 2800 37660 2860
rect 37580 2760 37600 2800
rect 37640 2760 37660 2800
rect 37580 2700 37660 2760
rect 37580 2660 37600 2700
rect 37640 2660 37660 2700
rect 37580 2600 37660 2660
rect 37580 2560 37600 2600
rect 37640 2560 37660 2600
rect 37580 2500 37660 2560
rect 37580 2460 37600 2500
rect 37640 2460 37660 2500
rect 37580 2430 37660 2460
rect 37760 3000 37840 3030
rect 37760 2960 37780 3000
rect 37820 2960 37840 3000
rect 37760 2900 37840 2960
rect 37760 2860 37780 2900
rect 37820 2860 37840 2900
rect 37760 2800 37840 2860
rect 37760 2760 37780 2800
rect 37820 2760 37840 2800
rect 37760 2700 37840 2760
rect 37760 2660 37780 2700
rect 37820 2660 37840 2700
rect 37760 2600 37840 2660
rect 37760 2560 37780 2600
rect 37820 2560 37840 2600
rect 37760 2500 37840 2560
rect 37760 2460 37780 2500
rect 37820 2460 37840 2500
rect 37760 2430 37840 2460
rect 37940 3000 38020 3030
rect 37940 2960 37960 3000
rect 38000 2960 38020 3000
rect 37940 2900 38020 2960
rect 37940 2860 37960 2900
rect 38000 2860 38020 2900
rect 37940 2800 38020 2860
rect 37940 2760 37960 2800
rect 38000 2760 38020 2800
rect 37940 2700 38020 2760
rect 37940 2660 37960 2700
rect 38000 2660 38020 2700
rect 37940 2600 38020 2660
rect 37940 2560 37960 2600
rect 38000 2560 38020 2600
rect 37940 2500 38020 2560
rect 37940 2460 37960 2500
rect 38000 2460 38020 2500
rect 37940 2430 38020 2460
rect 38120 3000 38200 3030
rect 38120 2960 38140 3000
rect 38180 2960 38200 3000
rect 38120 2900 38200 2960
rect 38120 2860 38140 2900
rect 38180 2860 38200 2900
rect 38120 2800 38200 2860
rect 38120 2760 38140 2800
rect 38180 2760 38200 2800
rect 38120 2700 38200 2760
rect 38120 2660 38140 2700
rect 38180 2660 38200 2700
rect 38120 2600 38200 2660
rect 38120 2560 38140 2600
rect 38180 2560 38200 2600
rect 38120 2500 38200 2560
rect 38120 2460 38140 2500
rect 38180 2460 38200 2500
rect 38120 2430 38200 2460
rect 38300 3000 38380 3030
rect 38300 2960 38320 3000
rect 38360 2960 38380 3000
rect 38300 2900 38380 2960
rect 38300 2860 38320 2900
rect 38360 2860 38380 2900
rect 38300 2800 38380 2860
rect 38300 2760 38320 2800
rect 38360 2760 38380 2800
rect 38300 2700 38380 2760
rect 38300 2660 38320 2700
rect 38360 2660 38380 2700
rect 38300 2600 38380 2660
rect 38300 2560 38320 2600
rect 38360 2560 38380 2600
rect 38300 2500 38380 2560
rect 38300 2460 38320 2500
rect 38360 2460 38380 2500
rect 38300 2430 38380 2460
rect 38480 3000 38560 3030
rect 38480 2960 38500 3000
rect 38540 2960 38560 3000
rect 38480 2900 38560 2960
rect 38480 2860 38500 2900
rect 38540 2860 38560 2900
rect 38480 2800 38560 2860
rect 38480 2760 38500 2800
rect 38540 2760 38560 2800
rect 38480 2700 38560 2760
rect 38480 2660 38500 2700
rect 38540 2660 38560 2700
rect 38480 2600 38560 2660
rect 38480 2560 38500 2600
rect 38540 2560 38560 2600
rect 38480 2500 38560 2560
rect 38480 2460 38500 2500
rect 38540 2460 38560 2500
rect 38480 2430 38560 2460
rect 38660 3000 38740 3030
rect 38660 2960 38680 3000
rect 38720 2960 38740 3000
rect 38660 2900 38740 2960
rect 38660 2860 38680 2900
rect 38720 2860 38740 2900
rect 38660 2800 38740 2860
rect 38660 2760 38680 2800
rect 38720 2760 38740 2800
rect 38660 2700 38740 2760
rect 38660 2660 38680 2700
rect 38720 2660 38740 2700
rect 38660 2600 38740 2660
rect 38660 2560 38680 2600
rect 38720 2560 38740 2600
rect 38660 2500 38740 2560
rect 38660 2460 38680 2500
rect 38720 2460 38740 2500
rect 38660 2430 38740 2460
rect 38840 3000 38920 3030
rect 38840 2960 38860 3000
rect 38900 2960 38920 3000
rect 38840 2900 38920 2960
rect 38840 2860 38860 2900
rect 38900 2860 38920 2900
rect 38840 2800 38920 2860
rect 38840 2760 38860 2800
rect 38900 2760 38920 2800
rect 38840 2700 38920 2760
rect 38840 2660 38860 2700
rect 38900 2660 38920 2700
rect 38840 2600 38920 2660
rect 38840 2560 38860 2600
rect 38900 2560 38920 2600
rect 38840 2500 38920 2560
rect 38840 2460 38860 2500
rect 38900 2460 38920 2500
rect 38840 2430 38920 2460
rect 39020 3000 39100 3030
rect 39020 2960 39040 3000
rect 39080 2960 39100 3000
rect 39020 2900 39100 2960
rect 39020 2860 39040 2900
rect 39080 2860 39100 2900
rect 39020 2800 39100 2860
rect 39020 2760 39040 2800
rect 39080 2760 39100 2800
rect 39020 2700 39100 2760
rect 39020 2660 39040 2700
rect 39080 2660 39100 2700
rect 39020 2600 39100 2660
rect 39020 2560 39040 2600
rect 39080 2560 39100 2600
rect 39020 2500 39100 2560
rect 39020 2460 39040 2500
rect 39080 2460 39100 2500
rect 39020 2430 39100 2460
rect 39200 3000 39280 3030
rect 39200 2960 39220 3000
rect 39260 2960 39280 3000
rect 39200 2900 39280 2960
rect 39200 2860 39220 2900
rect 39260 2860 39280 2900
rect 39200 2800 39280 2860
rect 39200 2760 39220 2800
rect 39260 2760 39280 2800
rect 39200 2700 39280 2760
rect 39200 2660 39220 2700
rect 39260 2660 39280 2700
rect 39200 2600 39280 2660
rect 39200 2560 39220 2600
rect 39260 2560 39280 2600
rect 39200 2500 39280 2560
rect 39200 2460 39220 2500
rect 39260 2460 39280 2500
rect 39200 2430 39280 2460
rect 39380 3000 39460 3030
rect 39380 2960 39400 3000
rect 39440 2960 39460 3000
rect 39380 2900 39460 2960
rect 39380 2860 39400 2900
rect 39440 2860 39460 2900
rect 39380 2800 39460 2860
rect 39380 2760 39400 2800
rect 39440 2760 39460 2800
rect 39380 2700 39460 2760
rect 39380 2660 39400 2700
rect 39440 2660 39460 2700
rect 39380 2600 39460 2660
rect 39380 2560 39400 2600
rect 39440 2560 39460 2600
rect 39380 2500 39460 2560
rect 39380 2460 39400 2500
rect 39440 2460 39460 2500
rect 39380 2430 39460 2460
rect 39560 3000 39640 3030
rect 39560 2960 39580 3000
rect 39620 2960 39640 3000
rect 39560 2900 39640 2960
rect 39560 2860 39580 2900
rect 39620 2860 39640 2900
rect 39560 2800 39640 2860
rect 39560 2760 39580 2800
rect 39620 2760 39640 2800
rect 39560 2700 39640 2760
rect 39560 2660 39580 2700
rect 39620 2660 39640 2700
rect 39560 2600 39640 2660
rect 39560 2560 39580 2600
rect 39620 2560 39640 2600
rect 39560 2500 39640 2560
rect 39560 2460 39580 2500
rect 39620 2460 39640 2500
rect 39560 2430 39640 2460
rect 39740 3000 39820 3030
rect 39740 2960 39760 3000
rect 39800 2960 39820 3000
rect 39740 2900 39820 2960
rect 39740 2860 39760 2900
rect 39800 2860 39820 2900
rect 39740 2800 39820 2860
rect 39740 2760 39760 2800
rect 39800 2760 39820 2800
rect 39740 2700 39820 2760
rect 39740 2660 39760 2700
rect 39800 2660 39820 2700
rect 39740 2600 39820 2660
rect 39740 2560 39760 2600
rect 39800 2560 39820 2600
rect 39740 2500 39820 2560
rect 39740 2460 39760 2500
rect 39800 2460 39820 2500
rect 39740 2430 39820 2460
rect 40360 2800 40440 2830
rect 40360 2760 40380 2800
rect 40420 2760 40440 2800
rect 40360 2700 40440 2760
rect 40360 2660 40380 2700
rect 40420 2660 40440 2700
rect 40360 2630 40440 2660
rect 40470 2800 40550 2830
rect 40470 2760 40490 2800
rect 40530 2760 40550 2800
rect 40470 2700 40550 2760
rect 40470 2660 40490 2700
rect 40530 2660 40550 2700
rect 40470 2630 40550 2660
rect 40580 2800 40660 2830
rect 40580 2760 40600 2800
rect 40640 2760 40660 2800
rect 40580 2700 40660 2760
rect 40580 2660 40600 2700
rect 40640 2660 40660 2700
rect 40580 2630 40660 2660
rect 40690 2800 40770 2830
rect 40690 2760 40710 2800
rect 40750 2760 40770 2800
rect 40690 2700 40770 2760
rect 40690 2660 40710 2700
rect 40750 2660 40770 2700
rect 40690 2630 40770 2660
rect 40800 2800 40880 2830
rect 40800 2760 40820 2800
rect 40860 2760 40880 2800
rect 40800 2700 40880 2760
rect 40800 2660 40820 2700
rect 40860 2660 40880 2700
rect 40800 2630 40880 2660
rect 35400 1620 35480 1650
rect 35400 1580 35420 1620
rect 35460 1580 35480 1620
rect 35400 1520 35480 1580
rect 35400 1480 35420 1520
rect 35460 1480 35480 1520
rect 35400 1450 35480 1480
rect 35520 1620 35600 1650
rect 35520 1580 35540 1620
rect 35580 1580 35600 1620
rect 35520 1520 35600 1580
rect 35520 1480 35540 1520
rect 35580 1480 35600 1520
rect 35520 1450 35600 1480
rect 35640 1620 35720 1650
rect 35640 1580 35660 1620
rect 35700 1580 35720 1620
rect 35640 1520 35720 1580
rect 35640 1480 35660 1520
rect 35700 1480 35720 1520
rect 35640 1450 35720 1480
rect 35760 1620 35840 1650
rect 35760 1580 35780 1620
rect 35820 1580 35840 1620
rect 35760 1520 35840 1580
rect 35760 1480 35780 1520
rect 35820 1480 35840 1520
rect 35760 1450 35840 1480
rect 35880 1620 35960 1650
rect 35880 1580 35900 1620
rect 35940 1580 35960 1620
rect 35880 1520 35960 1580
rect 35880 1480 35900 1520
rect 35940 1480 35960 1520
rect 35880 1450 35960 1480
rect 36000 1620 36080 1650
rect 36000 1580 36020 1620
rect 36060 1580 36080 1620
rect 36000 1520 36080 1580
rect 36000 1480 36020 1520
rect 36060 1480 36080 1520
rect 36000 1450 36080 1480
rect 36120 1620 36200 1650
rect 36120 1580 36140 1620
rect 36180 1580 36200 1620
rect 36120 1520 36200 1580
rect 36120 1480 36140 1520
rect 36180 1480 36200 1520
rect 36120 1450 36200 1480
rect 36240 1620 36320 1650
rect 36240 1580 36260 1620
rect 36300 1580 36320 1620
rect 36240 1520 36320 1580
rect 36240 1480 36260 1520
rect 36300 1480 36320 1520
rect 36240 1450 36320 1480
rect 36360 1620 36440 1650
rect 36360 1580 36380 1620
rect 36420 1580 36440 1620
rect 36360 1520 36440 1580
rect 36360 1480 36380 1520
rect 36420 1480 36440 1520
rect 36360 1450 36440 1480
rect 36480 1620 36560 1650
rect 36480 1580 36500 1620
rect 36540 1580 36560 1620
rect 36480 1520 36560 1580
rect 36480 1480 36500 1520
rect 36540 1480 36560 1520
rect 36480 1450 36560 1480
rect 36600 1620 36680 1650
rect 36600 1580 36620 1620
rect 36660 1580 36680 1620
rect 36600 1520 36680 1580
rect 36600 1480 36620 1520
rect 36660 1480 36680 1520
rect 36600 1450 36680 1480
rect 36720 1620 36800 1650
rect 36720 1580 36740 1620
rect 36780 1580 36800 1620
rect 36720 1520 36800 1580
rect 36720 1480 36740 1520
rect 36780 1480 36800 1520
rect 36720 1450 36800 1480
rect 36840 1620 36920 1650
rect 36840 1580 36860 1620
rect 36900 1580 36920 1620
rect 36840 1520 36920 1580
rect 36840 1480 36860 1520
rect 36900 1480 36920 1520
rect 36840 1450 36920 1480
rect 36960 1620 37040 1650
rect 36960 1580 36980 1620
rect 37020 1580 37040 1620
rect 36960 1520 37040 1580
rect 36960 1480 36980 1520
rect 37020 1480 37040 1520
rect 36960 1450 37040 1480
rect 37080 1620 37160 1650
rect 37080 1580 37100 1620
rect 37140 1580 37160 1620
rect 37080 1520 37160 1580
rect 37080 1480 37100 1520
rect 37140 1480 37160 1520
rect 37080 1450 37160 1480
rect 37200 1620 37280 1650
rect 37200 1580 37220 1620
rect 37260 1580 37280 1620
rect 37200 1520 37280 1580
rect 37200 1480 37220 1520
rect 37260 1480 37280 1520
rect 37200 1450 37280 1480
rect 37320 1620 37400 1650
rect 37320 1580 37340 1620
rect 37380 1580 37400 1620
rect 37320 1520 37400 1580
rect 37320 1480 37340 1520
rect 37380 1480 37400 1520
rect 37320 1450 37400 1480
rect 37440 1620 37520 1650
rect 37440 1580 37460 1620
rect 37500 1580 37520 1620
rect 37440 1520 37520 1580
rect 37440 1480 37460 1520
rect 37500 1480 37520 1520
rect 37440 1450 37520 1480
rect 37560 1620 37640 1650
rect 37560 1580 37580 1620
rect 37620 1580 37640 1620
rect 37560 1520 37640 1580
rect 37560 1480 37580 1520
rect 37620 1480 37640 1520
rect 37560 1450 37640 1480
rect 37680 1620 37760 1650
rect 37680 1580 37700 1620
rect 37740 1580 37760 1620
rect 37680 1520 37760 1580
rect 37680 1480 37700 1520
rect 37740 1480 37760 1520
rect 37680 1450 37760 1480
rect 37800 1620 37880 1650
rect 37800 1580 37820 1620
rect 37860 1580 37880 1620
rect 37800 1520 37880 1580
rect 37800 1480 37820 1520
rect 37860 1480 37880 1520
rect 37800 1450 37880 1480
rect 38440 1620 38520 1650
rect 38440 1580 38460 1620
rect 38500 1580 38520 1620
rect 38440 1520 38520 1580
rect 38440 1480 38460 1520
rect 38500 1480 38520 1520
rect 38440 1450 38520 1480
rect 38560 1620 38640 1650
rect 38560 1580 38580 1620
rect 38620 1580 38640 1620
rect 38560 1520 38640 1580
rect 38560 1480 38580 1520
rect 38620 1480 38640 1520
rect 38560 1450 38640 1480
rect 38680 1620 38760 1650
rect 38680 1580 38700 1620
rect 38740 1580 38760 1620
rect 38680 1520 38760 1580
rect 38680 1480 38700 1520
rect 38740 1480 38760 1520
rect 38680 1450 38760 1480
rect 38800 1620 38880 1650
rect 38800 1580 38820 1620
rect 38860 1580 38880 1620
rect 38800 1520 38880 1580
rect 38800 1480 38820 1520
rect 38860 1480 38880 1520
rect 38800 1450 38880 1480
rect 38920 1620 39000 1650
rect 38920 1580 38940 1620
rect 38980 1580 39000 1620
rect 38920 1520 39000 1580
rect 38920 1480 38940 1520
rect 38980 1480 39000 1520
rect 38920 1450 39000 1480
rect 39040 1620 39120 1650
rect 39040 1580 39060 1620
rect 39100 1580 39120 1620
rect 39040 1520 39120 1580
rect 39040 1480 39060 1520
rect 39100 1480 39120 1520
rect 39040 1450 39120 1480
rect 39160 1620 39240 1650
rect 39160 1580 39180 1620
rect 39220 1580 39240 1620
rect 39160 1520 39240 1580
rect 39160 1480 39180 1520
rect 39220 1480 39240 1520
rect 39160 1450 39240 1480
rect 39280 1620 39360 1650
rect 39280 1580 39300 1620
rect 39340 1580 39360 1620
rect 39280 1520 39360 1580
rect 39280 1480 39300 1520
rect 39340 1480 39360 1520
rect 39280 1450 39360 1480
rect 39400 1620 39480 1650
rect 39400 1580 39420 1620
rect 39460 1580 39480 1620
rect 39400 1520 39480 1580
rect 39400 1480 39420 1520
rect 39460 1480 39480 1520
rect 39400 1450 39480 1480
rect 39520 1620 39600 1650
rect 39520 1580 39540 1620
rect 39580 1580 39600 1620
rect 39520 1520 39600 1580
rect 39520 1480 39540 1520
rect 39580 1480 39600 1520
rect 39520 1450 39600 1480
rect 39640 1620 39720 1650
rect 39640 1580 39660 1620
rect 39700 1580 39720 1620
rect 39640 1520 39720 1580
rect 39640 1480 39660 1520
rect 39700 1480 39720 1520
rect 39640 1450 39720 1480
rect 39760 1620 39840 1650
rect 39760 1580 39780 1620
rect 39820 1580 39840 1620
rect 39760 1520 39840 1580
rect 39760 1480 39780 1520
rect 39820 1480 39840 1520
rect 39760 1450 39840 1480
rect 39880 1620 39960 1650
rect 39880 1580 39900 1620
rect 39940 1580 39960 1620
rect 39880 1520 39960 1580
rect 39880 1480 39900 1520
rect 39940 1480 39960 1520
rect 39880 1450 39960 1480
rect 40000 1620 40080 1650
rect 40000 1580 40020 1620
rect 40060 1580 40080 1620
rect 40000 1520 40080 1580
rect 40000 1480 40020 1520
rect 40060 1480 40080 1520
rect 40000 1450 40080 1480
rect 40120 1620 40200 1650
rect 40120 1580 40140 1620
rect 40180 1580 40200 1620
rect 40120 1520 40200 1580
rect 40120 1480 40140 1520
rect 40180 1480 40200 1520
rect 40120 1450 40200 1480
rect 40240 1620 40320 1650
rect 40240 1580 40260 1620
rect 40300 1580 40320 1620
rect 40240 1520 40320 1580
rect 40240 1480 40260 1520
rect 40300 1480 40320 1520
rect 40240 1450 40320 1480
rect 40360 1620 40440 1650
rect 40360 1580 40380 1620
rect 40420 1580 40440 1620
rect 40360 1520 40440 1580
rect 40360 1480 40380 1520
rect 40420 1480 40440 1520
rect 40360 1450 40440 1480
rect 40480 1620 40560 1650
rect 40480 1580 40500 1620
rect 40540 1580 40560 1620
rect 40480 1520 40560 1580
rect 40480 1480 40500 1520
rect 40540 1480 40560 1520
rect 40480 1450 40560 1480
rect 40600 1620 40680 1650
rect 40600 1580 40620 1620
rect 40660 1580 40680 1620
rect 40600 1520 40680 1580
rect 40600 1480 40620 1520
rect 40660 1480 40680 1520
rect 40600 1450 40680 1480
rect 40720 1620 40800 1650
rect 40720 1580 40740 1620
rect 40780 1580 40800 1620
rect 40720 1520 40800 1580
rect 40720 1480 40740 1520
rect 40780 1480 40800 1520
rect 40720 1450 40800 1480
rect 40840 1620 40920 1650
rect 40840 1580 40860 1620
rect 40900 1580 40920 1620
rect 40840 1520 40920 1580
rect 40840 1480 40860 1520
rect 40900 1480 40920 1520
rect 40840 1450 40920 1480
rect 33920 -4602 34600 -4550
rect 33920 -4636 33972 -4602
rect 34006 -4636 34062 -4602
rect 34096 -4636 34152 -4602
rect 34186 -4636 34242 -4602
rect 34276 -4636 34332 -4602
rect 34366 -4636 34422 -4602
rect 34456 -4636 34512 -4602
rect 34546 -4636 34600 -4602
rect 33920 -4692 34600 -4636
rect 33920 -4726 33972 -4692
rect 34006 -4726 34062 -4692
rect 34096 -4726 34152 -4692
rect 34186 -4726 34242 -4692
rect 34276 -4726 34332 -4692
rect 34366 -4726 34422 -4692
rect 34456 -4726 34512 -4692
rect 34546 -4726 34600 -4692
rect 33920 -4782 34600 -4726
rect 33920 -4816 33972 -4782
rect 34006 -4816 34062 -4782
rect 34096 -4816 34152 -4782
rect 34186 -4816 34242 -4782
rect 34276 -4816 34332 -4782
rect 34366 -4816 34422 -4782
rect 34456 -4816 34512 -4782
rect 34546 -4816 34600 -4782
rect 33920 -4872 34600 -4816
rect 33920 -4906 33972 -4872
rect 34006 -4906 34062 -4872
rect 34096 -4906 34152 -4872
rect 34186 -4906 34242 -4872
rect 34276 -4906 34332 -4872
rect 34366 -4906 34422 -4872
rect 34456 -4906 34512 -4872
rect 34546 -4906 34600 -4872
rect 33920 -4962 34600 -4906
rect 33920 -4996 33972 -4962
rect 34006 -4996 34062 -4962
rect 34096 -4996 34152 -4962
rect 34186 -4996 34242 -4962
rect 34276 -4996 34332 -4962
rect 34366 -4996 34422 -4962
rect 34456 -4996 34512 -4962
rect 34546 -4996 34600 -4962
rect 33920 -5052 34600 -4996
rect 33920 -5086 33972 -5052
rect 34006 -5086 34062 -5052
rect 34096 -5086 34152 -5052
rect 34186 -5086 34242 -5052
rect 34276 -5086 34332 -5052
rect 34366 -5086 34422 -5052
rect 34456 -5086 34512 -5052
rect 34546 -5086 34600 -5052
rect 33920 -5142 34600 -5086
rect 33920 -5176 33972 -5142
rect 34006 -5176 34062 -5142
rect 34096 -5176 34152 -5142
rect 34186 -5176 34242 -5142
rect 34276 -5176 34332 -5142
rect 34366 -5176 34422 -5142
rect 34456 -5176 34512 -5142
rect 34546 -5176 34600 -5142
rect 33920 -5230 34600 -5176
rect 35280 -4602 35960 -4550
rect 35280 -4636 35332 -4602
rect 35366 -4636 35422 -4602
rect 35456 -4636 35512 -4602
rect 35546 -4636 35602 -4602
rect 35636 -4636 35692 -4602
rect 35726 -4636 35782 -4602
rect 35816 -4636 35872 -4602
rect 35906 -4636 35960 -4602
rect 35280 -4692 35960 -4636
rect 35280 -4726 35332 -4692
rect 35366 -4726 35422 -4692
rect 35456 -4726 35512 -4692
rect 35546 -4726 35602 -4692
rect 35636 -4726 35692 -4692
rect 35726 -4726 35782 -4692
rect 35816 -4726 35872 -4692
rect 35906 -4726 35960 -4692
rect 35280 -4782 35960 -4726
rect 35280 -4816 35332 -4782
rect 35366 -4816 35422 -4782
rect 35456 -4816 35512 -4782
rect 35546 -4816 35602 -4782
rect 35636 -4816 35692 -4782
rect 35726 -4816 35782 -4782
rect 35816 -4816 35872 -4782
rect 35906 -4816 35960 -4782
rect 35280 -4872 35960 -4816
rect 35280 -4906 35332 -4872
rect 35366 -4906 35422 -4872
rect 35456 -4906 35512 -4872
rect 35546 -4906 35602 -4872
rect 35636 -4906 35692 -4872
rect 35726 -4906 35782 -4872
rect 35816 -4906 35872 -4872
rect 35906 -4906 35960 -4872
rect 35280 -4962 35960 -4906
rect 35280 -4996 35332 -4962
rect 35366 -4996 35422 -4962
rect 35456 -4996 35512 -4962
rect 35546 -4996 35602 -4962
rect 35636 -4996 35692 -4962
rect 35726 -4996 35782 -4962
rect 35816 -4996 35872 -4962
rect 35906 -4996 35960 -4962
rect 35280 -5052 35960 -4996
rect 35280 -5086 35332 -5052
rect 35366 -5086 35422 -5052
rect 35456 -5086 35512 -5052
rect 35546 -5086 35602 -5052
rect 35636 -5086 35692 -5052
rect 35726 -5086 35782 -5052
rect 35816 -5086 35872 -5052
rect 35906 -5086 35960 -5052
rect 35280 -5142 35960 -5086
rect 35280 -5176 35332 -5142
rect 35366 -5176 35422 -5142
rect 35456 -5176 35512 -5142
rect 35546 -5176 35602 -5142
rect 35636 -5176 35692 -5142
rect 35726 -5176 35782 -5142
rect 35816 -5176 35872 -5142
rect 35906 -5176 35960 -5142
rect 35280 -5230 35960 -5176
rect 36640 -4602 37320 -4550
rect 36640 -4636 36692 -4602
rect 36726 -4636 36782 -4602
rect 36816 -4636 36872 -4602
rect 36906 -4636 36962 -4602
rect 36996 -4636 37052 -4602
rect 37086 -4636 37142 -4602
rect 37176 -4636 37232 -4602
rect 37266 -4636 37320 -4602
rect 36640 -4692 37320 -4636
rect 36640 -4726 36692 -4692
rect 36726 -4726 36782 -4692
rect 36816 -4726 36872 -4692
rect 36906 -4726 36962 -4692
rect 36996 -4726 37052 -4692
rect 37086 -4726 37142 -4692
rect 37176 -4726 37232 -4692
rect 37266 -4726 37320 -4692
rect 36640 -4782 37320 -4726
rect 36640 -4816 36692 -4782
rect 36726 -4816 36782 -4782
rect 36816 -4816 36872 -4782
rect 36906 -4816 36962 -4782
rect 36996 -4816 37052 -4782
rect 37086 -4816 37142 -4782
rect 37176 -4816 37232 -4782
rect 37266 -4816 37320 -4782
rect 36640 -4872 37320 -4816
rect 36640 -4906 36692 -4872
rect 36726 -4906 36782 -4872
rect 36816 -4906 36872 -4872
rect 36906 -4906 36962 -4872
rect 36996 -4906 37052 -4872
rect 37086 -4906 37142 -4872
rect 37176 -4906 37232 -4872
rect 37266 -4906 37320 -4872
rect 36640 -4962 37320 -4906
rect 36640 -4996 36692 -4962
rect 36726 -4996 36782 -4962
rect 36816 -4996 36872 -4962
rect 36906 -4996 36962 -4962
rect 36996 -4996 37052 -4962
rect 37086 -4996 37142 -4962
rect 37176 -4996 37232 -4962
rect 37266 -4996 37320 -4962
rect 36640 -5052 37320 -4996
rect 36640 -5086 36692 -5052
rect 36726 -5086 36782 -5052
rect 36816 -5086 36872 -5052
rect 36906 -5086 36962 -5052
rect 36996 -5086 37052 -5052
rect 37086 -5086 37142 -5052
rect 37176 -5086 37232 -5052
rect 37266 -5086 37320 -5052
rect 36640 -5142 37320 -5086
rect 36640 -5176 36692 -5142
rect 36726 -5176 36782 -5142
rect 36816 -5176 36872 -5142
rect 36906 -5176 36962 -5142
rect 36996 -5176 37052 -5142
rect 37086 -5176 37142 -5142
rect 37176 -5176 37232 -5142
rect 37266 -5176 37320 -5142
rect 36640 -5230 37320 -5176
rect 33920 -5962 34600 -5910
rect 33920 -5996 33972 -5962
rect 34006 -5996 34062 -5962
rect 34096 -5996 34152 -5962
rect 34186 -5996 34242 -5962
rect 34276 -5996 34332 -5962
rect 34366 -5996 34422 -5962
rect 34456 -5996 34512 -5962
rect 34546 -5996 34600 -5962
rect 33920 -6052 34600 -5996
rect 33920 -6086 33972 -6052
rect 34006 -6086 34062 -6052
rect 34096 -6086 34152 -6052
rect 34186 -6086 34242 -6052
rect 34276 -6086 34332 -6052
rect 34366 -6086 34422 -6052
rect 34456 -6086 34512 -6052
rect 34546 -6086 34600 -6052
rect 33920 -6142 34600 -6086
rect 33920 -6176 33972 -6142
rect 34006 -6176 34062 -6142
rect 34096 -6176 34152 -6142
rect 34186 -6176 34242 -6142
rect 34276 -6176 34332 -6142
rect 34366 -6176 34422 -6142
rect 34456 -6176 34512 -6142
rect 34546 -6176 34600 -6142
rect 33920 -6232 34600 -6176
rect 33920 -6266 33972 -6232
rect 34006 -6266 34062 -6232
rect 34096 -6266 34152 -6232
rect 34186 -6266 34242 -6232
rect 34276 -6266 34332 -6232
rect 34366 -6266 34422 -6232
rect 34456 -6266 34512 -6232
rect 34546 -6266 34600 -6232
rect 33920 -6322 34600 -6266
rect 33920 -6356 33972 -6322
rect 34006 -6356 34062 -6322
rect 34096 -6356 34152 -6322
rect 34186 -6356 34242 -6322
rect 34276 -6356 34332 -6322
rect 34366 -6356 34422 -6322
rect 34456 -6356 34512 -6322
rect 34546 -6356 34600 -6322
rect 33920 -6412 34600 -6356
rect 33920 -6446 33972 -6412
rect 34006 -6446 34062 -6412
rect 34096 -6446 34152 -6412
rect 34186 -6446 34242 -6412
rect 34276 -6446 34332 -6412
rect 34366 -6446 34422 -6412
rect 34456 -6446 34512 -6412
rect 34546 -6446 34600 -6412
rect 33920 -6502 34600 -6446
rect 33920 -6536 33972 -6502
rect 34006 -6536 34062 -6502
rect 34096 -6536 34152 -6502
rect 34186 -6536 34242 -6502
rect 34276 -6536 34332 -6502
rect 34366 -6536 34422 -6502
rect 34456 -6536 34512 -6502
rect 34546 -6536 34600 -6502
rect 33920 -6590 34600 -6536
rect 35280 -5962 35960 -5910
rect 35280 -5996 35332 -5962
rect 35366 -5996 35422 -5962
rect 35456 -5996 35512 -5962
rect 35546 -5996 35602 -5962
rect 35636 -5996 35692 -5962
rect 35726 -5996 35782 -5962
rect 35816 -5996 35872 -5962
rect 35906 -5996 35960 -5962
rect 35280 -6052 35960 -5996
rect 35280 -6086 35332 -6052
rect 35366 -6086 35422 -6052
rect 35456 -6086 35512 -6052
rect 35546 -6086 35602 -6052
rect 35636 -6086 35692 -6052
rect 35726 -6086 35782 -6052
rect 35816 -6086 35872 -6052
rect 35906 -6086 35960 -6052
rect 35280 -6142 35960 -6086
rect 35280 -6176 35332 -6142
rect 35366 -6176 35422 -6142
rect 35456 -6176 35512 -6142
rect 35546 -6176 35602 -6142
rect 35636 -6176 35692 -6142
rect 35726 -6176 35782 -6142
rect 35816 -6176 35872 -6142
rect 35906 -6176 35960 -6142
rect 35280 -6232 35960 -6176
rect 35280 -6266 35332 -6232
rect 35366 -6266 35422 -6232
rect 35456 -6266 35512 -6232
rect 35546 -6266 35602 -6232
rect 35636 -6266 35692 -6232
rect 35726 -6266 35782 -6232
rect 35816 -6266 35872 -6232
rect 35906 -6266 35960 -6232
rect 35280 -6322 35960 -6266
rect 35280 -6356 35332 -6322
rect 35366 -6356 35422 -6322
rect 35456 -6356 35512 -6322
rect 35546 -6356 35602 -6322
rect 35636 -6356 35692 -6322
rect 35726 -6356 35782 -6322
rect 35816 -6356 35872 -6322
rect 35906 -6356 35960 -6322
rect 35280 -6412 35960 -6356
rect 35280 -6446 35332 -6412
rect 35366 -6446 35422 -6412
rect 35456 -6446 35512 -6412
rect 35546 -6446 35602 -6412
rect 35636 -6446 35692 -6412
rect 35726 -6446 35782 -6412
rect 35816 -6446 35872 -6412
rect 35906 -6446 35960 -6412
rect 35280 -6502 35960 -6446
rect 35280 -6536 35332 -6502
rect 35366 -6536 35422 -6502
rect 35456 -6536 35512 -6502
rect 35546 -6536 35602 -6502
rect 35636 -6536 35692 -6502
rect 35726 -6536 35782 -6502
rect 35816 -6536 35872 -6502
rect 35906 -6536 35960 -6502
rect 35280 -6590 35960 -6536
rect 36640 -5962 37320 -5910
rect 36640 -5996 36692 -5962
rect 36726 -5996 36782 -5962
rect 36816 -5996 36872 -5962
rect 36906 -5996 36962 -5962
rect 36996 -5996 37052 -5962
rect 37086 -5996 37142 -5962
rect 37176 -5996 37232 -5962
rect 37266 -5996 37320 -5962
rect 36640 -6052 37320 -5996
rect 36640 -6086 36692 -6052
rect 36726 -6086 36782 -6052
rect 36816 -6086 36872 -6052
rect 36906 -6086 36962 -6052
rect 36996 -6086 37052 -6052
rect 37086 -6086 37142 -6052
rect 37176 -6086 37232 -6052
rect 37266 -6086 37320 -6052
rect 36640 -6142 37320 -6086
rect 36640 -6176 36692 -6142
rect 36726 -6176 36782 -6142
rect 36816 -6176 36872 -6142
rect 36906 -6176 36962 -6142
rect 36996 -6176 37052 -6142
rect 37086 -6176 37142 -6142
rect 37176 -6176 37232 -6142
rect 37266 -6176 37320 -6142
rect 36640 -6232 37320 -6176
rect 36640 -6266 36692 -6232
rect 36726 -6266 36782 -6232
rect 36816 -6266 36872 -6232
rect 36906 -6266 36962 -6232
rect 36996 -6266 37052 -6232
rect 37086 -6266 37142 -6232
rect 37176 -6266 37232 -6232
rect 37266 -6266 37320 -6232
rect 36640 -6322 37320 -6266
rect 36640 -6356 36692 -6322
rect 36726 -6356 36782 -6322
rect 36816 -6356 36872 -6322
rect 36906 -6356 36962 -6322
rect 36996 -6356 37052 -6322
rect 37086 -6356 37142 -6322
rect 37176 -6356 37232 -6322
rect 37266 -6356 37320 -6322
rect 36640 -6412 37320 -6356
rect 36640 -6446 36692 -6412
rect 36726 -6446 36782 -6412
rect 36816 -6446 36872 -6412
rect 36906 -6446 36962 -6412
rect 36996 -6446 37052 -6412
rect 37086 -6446 37142 -6412
rect 37176 -6446 37232 -6412
rect 37266 -6446 37320 -6412
rect 36640 -6502 37320 -6446
rect 36640 -6536 36692 -6502
rect 36726 -6536 36782 -6502
rect 36816 -6536 36872 -6502
rect 36906 -6536 36962 -6502
rect 36996 -6536 37052 -6502
rect 37086 -6536 37142 -6502
rect 37176 -6536 37232 -6502
rect 37266 -6536 37320 -6502
rect 36640 -6590 37320 -6536
rect 33920 -7322 34600 -7270
rect 33920 -7356 33972 -7322
rect 34006 -7356 34062 -7322
rect 34096 -7356 34152 -7322
rect 34186 -7356 34242 -7322
rect 34276 -7356 34332 -7322
rect 34366 -7356 34422 -7322
rect 34456 -7356 34512 -7322
rect 34546 -7356 34600 -7322
rect 33920 -7412 34600 -7356
rect 33920 -7446 33972 -7412
rect 34006 -7446 34062 -7412
rect 34096 -7446 34152 -7412
rect 34186 -7446 34242 -7412
rect 34276 -7446 34332 -7412
rect 34366 -7446 34422 -7412
rect 34456 -7446 34512 -7412
rect 34546 -7446 34600 -7412
rect 33920 -7502 34600 -7446
rect 33920 -7536 33972 -7502
rect 34006 -7536 34062 -7502
rect 34096 -7536 34152 -7502
rect 34186 -7536 34242 -7502
rect 34276 -7536 34332 -7502
rect 34366 -7536 34422 -7502
rect 34456 -7536 34512 -7502
rect 34546 -7536 34600 -7502
rect 33920 -7592 34600 -7536
rect 33920 -7626 33972 -7592
rect 34006 -7626 34062 -7592
rect 34096 -7626 34152 -7592
rect 34186 -7626 34242 -7592
rect 34276 -7626 34332 -7592
rect 34366 -7626 34422 -7592
rect 34456 -7626 34512 -7592
rect 34546 -7626 34600 -7592
rect 33920 -7682 34600 -7626
rect 33920 -7716 33972 -7682
rect 34006 -7716 34062 -7682
rect 34096 -7716 34152 -7682
rect 34186 -7716 34242 -7682
rect 34276 -7716 34332 -7682
rect 34366 -7716 34422 -7682
rect 34456 -7716 34512 -7682
rect 34546 -7716 34600 -7682
rect 33920 -7772 34600 -7716
rect 33920 -7806 33972 -7772
rect 34006 -7806 34062 -7772
rect 34096 -7806 34152 -7772
rect 34186 -7806 34242 -7772
rect 34276 -7806 34332 -7772
rect 34366 -7806 34422 -7772
rect 34456 -7806 34512 -7772
rect 34546 -7806 34600 -7772
rect 33920 -7862 34600 -7806
rect 33920 -7896 33972 -7862
rect 34006 -7896 34062 -7862
rect 34096 -7896 34152 -7862
rect 34186 -7896 34242 -7862
rect 34276 -7896 34332 -7862
rect 34366 -7896 34422 -7862
rect 34456 -7896 34512 -7862
rect 34546 -7896 34600 -7862
rect 33920 -7950 34600 -7896
rect 35280 -7322 35960 -7270
rect 35280 -7356 35332 -7322
rect 35366 -7356 35422 -7322
rect 35456 -7356 35512 -7322
rect 35546 -7356 35602 -7322
rect 35636 -7356 35692 -7322
rect 35726 -7356 35782 -7322
rect 35816 -7356 35872 -7322
rect 35906 -7356 35960 -7322
rect 35280 -7412 35960 -7356
rect 35280 -7446 35332 -7412
rect 35366 -7446 35422 -7412
rect 35456 -7446 35512 -7412
rect 35546 -7446 35602 -7412
rect 35636 -7446 35692 -7412
rect 35726 -7446 35782 -7412
rect 35816 -7446 35872 -7412
rect 35906 -7446 35960 -7412
rect 35280 -7502 35960 -7446
rect 35280 -7536 35332 -7502
rect 35366 -7536 35422 -7502
rect 35456 -7536 35512 -7502
rect 35546 -7536 35602 -7502
rect 35636 -7536 35692 -7502
rect 35726 -7536 35782 -7502
rect 35816 -7536 35872 -7502
rect 35906 -7536 35960 -7502
rect 35280 -7592 35960 -7536
rect 35280 -7626 35332 -7592
rect 35366 -7626 35422 -7592
rect 35456 -7626 35512 -7592
rect 35546 -7626 35602 -7592
rect 35636 -7626 35692 -7592
rect 35726 -7626 35782 -7592
rect 35816 -7626 35872 -7592
rect 35906 -7626 35960 -7592
rect 35280 -7682 35960 -7626
rect 35280 -7716 35332 -7682
rect 35366 -7716 35422 -7682
rect 35456 -7716 35512 -7682
rect 35546 -7716 35602 -7682
rect 35636 -7716 35692 -7682
rect 35726 -7716 35782 -7682
rect 35816 -7716 35872 -7682
rect 35906 -7716 35960 -7682
rect 35280 -7772 35960 -7716
rect 35280 -7806 35332 -7772
rect 35366 -7806 35422 -7772
rect 35456 -7806 35512 -7772
rect 35546 -7806 35602 -7772
rect 35636 -7806 35692 -7772
rect 35726 -7806 35782 -7772
rect 35816 -7806 35872 -7772
rect 35906 -7806 35960 -7772
rect 35280 -7862 35960 -7806
rect 35280 -7896 35332 -7862
rect 35366 -7896 35422 -7862
rect 35456 -7896 35512 -7862
rect 35546 -7896 35602 -7862
rect 35636 -7896 35692 -7862
rect 35726 -7896 35782 -7862
rect 35816 -7896 35872 -7862
rect 35906 -7896 35960 -7862
rect 35280 -7950 35960 -7896
rect 36640 -7322 37320 -7270
rect 36640 -7356 36692 -7322
rect 36726 -7356 36782 -7322
rect 36816 -7356 36872 -7322
rect 36906 -7356 36962 -7322
rect 36996 -7356 37052 -7322
rect 37086 -7356 37142 -7322
rect 37176 -7356 37232 -7322
rect 37266 -7356 37320 -7322
rect 36640 -7412 37320 -7356
rect 36640 -7446 36692 -7412
rect 36726 -7446 36782 -7412
rect 36816 -7446 36872 -7412
rect 36906 -7446 36962 -7412
rect 36996 -7446 37052 -7412
rect 37086 -7446 37142 -7412
rect 37176 -7446 37232 -7412
rect 37266 -7446 37320 -7412
rect 36640 -7502 37320 -7446
rect 36640 -7536 36692 -7502
rect 36726 -7536 36782 -7502
rect 36816 -7536 36872 -7502
rect 36906 -7536 36962 -7502
rect 36996 -7536 37052 -7502
rect 37086 -7536 37142 -7502
rect 37176 -7536 37232 -7502
rect 37266 -7536 37320 -7502
rect 36640 -7592 37320 -7536
rect 36640 -7626 36692 -7592
rect 36726 -7626 36782 -7592
rect 36816 -7626 36872 -7592
rect 36906 -7626 36962 -7592
rect 36996 -7626 37052 -7592
rect 37086 -7626 37142 -7592
rect 37176 -7626 37232 -7592
rect 37266 -7626 37320 -7592
rect 36640 -7682 37320 -7626
rect 36640 -7716 36692 -7682
rect 36726 -7716 36782 -7682
rect 36816 -7716 36872 -7682
rect 36906 -7716 36962 -7682
rect 36996 -7716 37052 -7682
rect 37086 -7716 37142 -7682
rect 37176 -7716 37232 -7682
rect 37266 -7716 37320 -7682
rect 36640 -7772 37320 -7716
rect 36640 -7806 36692 -7772
rect 36726 -7806 36782 -7772
rect 36816 -7806 36872 -7772
rect 36906 -7806 36962 -7772
rect 36996 -7806 37052 -7772
rect 37086 -7806 37142 -7772
rect 37176 -7806 37232 -7772
rect 37266 -7806 37320 -7772
rect 36640 -7862 37320 -7806
rect 36640 -7896 36692 -7862
rect 36726 -7896 36782 -7862
rect 36816 -7896 36872 -7862
rect 36906 -7896 36962 -7862
rect 36996 -7896 37052 -7862
rect 37086 -7896 37142 -7862
rect 37176 -7896 37232 -7862
rect 37266 -7896 37320 -7862
rect 36640 -7950 37320 -7896
<< ndiffc >>
rect 6280 3830 6320 3870
rect 6400 3830 6440 3870
rect 6520 3830 6560 3870
rect 6640 3830 6680 3870
rect 6760 3830 6800 3870
rect 6880 3830 6920 3870
rect 7000 3830 7040 3870
rect 7120 3830 7160 3870
rect 7240 3830 7280 3870
rect 7360 3830 7400 3870
rect 7480 3830 7520 3870
rect 8800 3830 8840 3870
rect 8920 3830 8960 3870
rect 9040 3830 9080 3870
rect 9160 3830 9200 3870
rect 9280 3830 9320 3870
rect 9400 3830 9440 3870
rect 9520 3830 9560 3870
rect 9640 3830 9680 3870
rect 9760 3830 9800 3870
rect 9880 3830 9920 3870
rect 10000 3830 10040 3870
rect 5800 3280 5840 3320
rect 5800 3180 5840 3220
rect 5800 3080 5840 3120
rect 5800 2980 5840 3020
rect 5800 2880 5840 2920
rect 6880 3280 6920 3320
rect 6880 3180 6920 3220
rect 6880 3080 6920 3120
rect 6880 2980 6920 3020
rect 6880 2880 6920 2920
rect 7960 3280 8000 3320
rect 7960 3180 8000 3220
rect 7960 3080 8000 3120
rect 7960 2980 8000 3020
rect 7960 2880 8000 2920
rect 8320 3280 8360 3320
rect 8320 3180 8360 3220
rect 8320 3080 8360 3120
rect 8320 2980 8360 3020
rect 8320 2880 8360 2920
rect 9400 3280 9440 3320
rect 9400 3180 9440 3220
rect 9400 3080 9440 3120
rect 9400 2980 9440 3020
rect 9400 2880 9440 2920
rect 10480 3280 10520 3320
rect 10480 3180 10520 3220
rect 10480 3080 10520 3120
rect 10480 2980 10520 3020
rect 10480 2880 10520 2920
rect 6060 2340 6100 2380
rect 6060 2240 6100 2280
rect 8140 2340 8180 2380
rect 8140 2240 8180 2280
rect 10220 2340 10260 2380
rect 10220 2240 10260 2280
rect 6360 1790 6400 1830
rect 6360 1690 6400 1730
rect 6470 1790 6510 1830
rect 6470 1690 6510 1730
rect 6580 1790 6620 1830
rect 6580 1690 6620 1730
rect 6690 1790 6730 1830
rect 6690 1690 6730 1730
rect 6800 1790 6840 1830
rect 6800 1690 6840 1730
rect 6910 1790 6950 1830
rect 6910 1690 6950 1730
rect 7020 1790 7060 1830
rect 7020 1690 7060 1730
rect 7130 1790 7170 1830
rect 7130 1690 7170 1730
rect 7240 1790 7280 1830
rect 7240 1690 7280 1730
rect 7590 1790 7630 1830
rect 7590 1690 7630 1730
rect 7700 1790 7740 1830
rect 7700 1690 7740 1730
rect 7810 1790 7850 1830
rect 7810 1690 7850 1730
rect 7920 1790 7960 1830
rect 7920 1690 7960 1730
rect 8030 1790 8070 1830
rect 8030 1690 8070 1730
rect 8140 1790 8180 1830
rect 8140 1690 8180 1730
rect 8250 1790 8290 1830
rect 8250 1690 8290 1730
rect 8360 1790 8400 1830
rect 8360 1690 8400 1730
rect 8470 1790 8510 1830
rect 8470 1690 8510 1730
rect 8580 1790 8620 1830
rect 8580 1690 8620 1730
rect 8690 1790 8730 1830
rect 8690 1690 8730 1730
rect 9040 1790 9080 1830
rect 9040 1690 9080 1730
rect 9150 1790 9190 1830
rect 9150 1690 9190 1730
rect 9260 1790 9300 1830
rect 9260 1690 9300 1730
rect 9370 1790 9410 1830
rect 9370 1690 9410 1730
rect 9480 1790 9520 1830
rect 9480 1690 9520 1730
rect 9590 1790 9630 1830
rect 9590 1690 9630 1730
rect 9700 1790 9740 1830
rect 9700 1690 9740 1730
rect 9810 1790 9850 1830
rect 9810 1690 9850 1730
rect 9920 1790 9960 1830
rect 9920 1690 9960 1730
rect 36280 830 36320 870
rect 36400 830 36440 870
rect 36520 830 36560 870
rect 36640 830 36680 870
rect 36760 830 36800 870
rect 36880 830 36920 870
rect 37000 830 37040 870
rect 37120 830 37160 870
rect 37240 830 37280 870
rect 37360 830 37400 870
rect 37480 830 37520 870
rect 38800 830 38840 870
rect 38920 830 38960 870
rect 39040 830 39080 870
rect 39160 830 39200 870
rect 39280 830 39320 870
rect 39400 830 39440 870
rect 39520 830 39560 870
rect 39640 830 39680 870
rect 39760 830 39800 870
rect 39880 830 39920 870
rect 40000 830 40040 870
rect 35800 280 35840 320
rect 35800 180 35840 220
rect 35800 80 35840 120
rect 35800 -20 35840 20
rect 35800 -120 35840 -80
rect 36880 280 36920 320
rect 36880 180 36920 220
rect 36880 80 36920 120
rect 36880 -20 36920 20
rect 36880 -120 36920 -80
rect 37960 280 38000 320
rect 37960 180 38000 220
rect 37960 80 38000 120
rect 37960 -20 38000 20
rect 37960 -120 38000 -80
rect 38320 280 38360 320
rect 38320 180 38360 220
rect 38320 80 38360 120
rect 38320 -20 38360 20
rect 38320 -120 38360 -80
rect 39400 280 39440 320
rect 39400 180 39440 220
rect 39400 80 39440 120
rect 39400 -20 39440 20
rect 39400 -120 39440 -80
rect 40480 280 40520 320
rect 40480 180 40520 220
rect 40480 80 40520 120
rect 40480 -20 40520 20
rect 40480 -120 40520 -80
rect 36060 -660 36100 -620
rect 36060 -760 36100 -720
rect 38140 -660 38180 -620
rect 38140 -760 38180 -720
rect 40220 -660 40260 -620
rect 40220 -760 40260 -720
rect 36360 -1210 36400 -1170
rect 36360 -1310 36400 -1270
rect 36470 -1210 36510 -1170
rect 36470 -1310 36510 -1270
rect 36580 -1210 36620 -1170
rect 36580 -1310 36620 -1270
rect 36690 -1210 36730 -1170
rect 36690 -1310 36730 -1270
rect 36800 -1210 36840 -1170
rect 36800 -1310 36840 -1270
rect 36910 -1210 36950 -1170
rect 36910 -1310 36950 -1270
rect 37020 -1210 37060 -1170
rect 37020 -1310 37060 -1270
rect 37130 -1210 37170 -1170
rect 37130 -1310 37170 -1270
rect 37240 -1210 37280 -1170
rect 37240 -1310 37280 -1270
rect 37590 -1210 37630 -1170
rect 37590 -1310 37630 -1270
rect 37700 -1210 37740 -1170
rect 37700 -1310 37740 -1270
rect 37810 -1210 37850 -1170
rect 37810 -1310 37850 -1270
rect 37920 -1210 37960 -1170
rect 37920 -1310 37960 -1270
rect 38030 -1210 38070 -1170
rect 38030 -1310 38070 -1270
rect 38140 -1210 38180 -1170
rect 38140 -1310 38180 -1270
rect 38250 -1210 38290 -1170
rect 38250 -1310 38290 -1270
rect 38360 -1210 38400 -1170
rect 38360 -1310 38400 -1270
rect 38470 -1210 38510 -1170
rect 38470 -1310 38510 -1270
rect 38580 -1210 38620 -1170
rect 38580 -1310 38620 -1270
rect 38690 -1210 38730 -1170
rect 38690 -1310 38730 -1270
rect 39040 -1210 39080 -1170
rect 39040 -1310 39080 -1270
rect 39150 -1210 39190 -1170
rect 39150 -1310 39190 -1270
rect 39260 -1210 39300 -1170
rect 39260 -1310 39300 -1270
rect 39370 -1210 39410 -1170
rect 39370 -1310 39410 -1270
rect 39480 -1210 39520 -1170
rect 39480 -1310 39520 -1270
rect 39590 -1210 39630 -1170
rect 39590 -1310 39630 -1270
rect 39700 -1210 39740 -1170
rect 39700 -1310 39740 -1270
rect 39810 -1210 39850 -1170
rect 39810 -1310 39850 -1270
rect 39920 -1210 39960 -1170
rect 39920 -1310 39960 -1270
<< pdiffc >>
rect 6090 6786 6130 6930
rect 6200 6786 6240 6930
rect 6310 6786 6350 6930
rect 6420 6786 6460 6930
rect 6530 6786 6570 6930
rect 6640 6786 6680 6930
rect 6750 6786 6790 6930
rect 7370 6890 7410 6930
rect 7370 6790 7410 6830
rect 7480 6890 7520 6930
rect 7480 6790 7520 6830
rect 7590 6890 7630 6930
rect 7590 6790 7630 6830
rect 7700 6890 7740 6930
rect 7700 6790 7740 6830
rect 7810 6890 7850 6930
rect 7810 6790 7850 6830
rect 7920 6890 7960 6930
rect 7920 6790 7960 6830
rect 8030 6890 8070 6930
rect 8030 6790 8070 6830
rect 8140 6890 8180 6930
rect 8140 6790 8180 6830
rect 8250 6890 8290 6930
rect 8250 6790 8290 6830
rect 8360 6890 8400 6930
rect 8360 6790 8400 6830
rect 8470 6890 8510 6930
rect 8470 6790 8510 6830
rect 8580 6890 8620 6930
rect 8580 6790 8620 6830
rect 8690 6890 8730 6930
rect 8690 6790 8730 6830
rect 9530 6790 9570 6930
rect 9640 6790 9680 6930
rect 9750 6790 9790 6930
rect 9860 6790 9900 6930
rect 9970 6790 10010 6930
rect 10080 6790 10120 6930
rect 10190 6790 10230 6930
rect 5450 5760 5490 5800
rect 5450 5660 5490 5700
rect 5560 5760 5600 5800
rect 5560 5660 5600 5700
rect 5670 5760 5710 5800
rect 5670 5660 5710 5700
rect 5780 5760 5820 5800
rect 5780 5660 5820 5700
rect 5890 5760 5930 5800
rect 5890 5660 5930 5700
rect 6520 5960 6560 6000
rect 6520 5860 6560 5900
rect 6520 5760 6560 5800
rect 6520 5660 6560 5700
rect 6520 5560 6560 5600
rect 6520 5460 6560 5500
rect 6700 5960 6740 6000
rect 6700 5860 6740 5900
rect 6700 5760 6740 5800
rect 6700 5660 6740 5700
rect 6700 5560 6740 5600
rect 6700 5460 6740 5500
rect 6880 5960 6920 6000
rect 6880 5860 6920 5900
rect 6880 5760 6920 5800
rect 6880 5660 6920 5700
rect 6880 5560 6920 5600
rect 6880 5460 6920 5500
rect 7060 5960 7100 6000
rect 7060 5860 7100 5900
rect 7060 5760 7100 5800
rect 7060 5660 7100 5700
rect 7060 5560 7100 5600
rect 7060 5460 7100 5500
rect 7240 5960 7280 6000
rect 7240 5860 7280 5900
rect 7240 5760 7280 5800
rect 7240 5660 7280 5700
rect 7240 5560 7280 5600
rect 7240 5460 7280 5500
rect 7420 5960 7460 6000
rect 7420 5860 7460 5900
rect 7420 5760 7460 5800
rect 7420 5660 7460 5700
rect 7420 5560 7460 5600
rect 7420 5460 7460 5500
rect 7600 5960 7640 6000
rect 7600 5860 7640 5900
rect 7600 5760 7640 5800
rect 7600 5660 7640 5700
rect 7600 5560 7640 5600
rect 7600 5460 7640 5500
rect 7780 5960 7820 6000
rect 7780 5860 7820 5900
rect 7780 5760 7820 5800
rect 7780 5660 7820 5700
rect 7780 5560 7820 5600
rect 7780 5460 7820 5500
rect 7960 5960 8000 6000
rect 7960 5860 8000 5900
rect 7960 5760 8000 5800
rect 7960 5660 8000 5700
rect 7960 5560 8000 5600
rect 7960 5460 8000 5500
rect 8140 5960 8180 6000
rect 8140 5860 8180 5900
rect 8140 5760 8180 5800
rect 8140 5660 8180 5700
rect 8140 5560 8180 5600
rect 8140 5460 8180 5500
rect 8320 5960 8360 6000
rect 8320 5860 8360 5900
rect 8320 5760 8360 5800
rect 8320 5660 8360 5700
rect 8320 5560 8360 5600
rect 8320 5460 8360 5500
rect 8500 5960 8540 6000
rect 8500 5860 8540 5900
rect 8500 5760 8540 5800
rect 8500 5660 8540 5700
rect 8500 5560 8540 5600
rect 8500 5460 8540 5500
rect 8680 5960 8720 6000
rect 8680 5860 8720 5900
rect 8680 5760 8720 5800
rect 8680 5660 8720 5700
rect 8680 5560 8720 5600
rect 8680 5460 8720 5500
rect 8860 5960 8900 6000
rect 8860 5860 8900 5900
rect 8860 5760 8900 5800
rect 8860 5660 8900 5700
rect 8860 5560 8900 5600
rect 8860 5460 8900 5500
rect 9040 5960 9080 6000
rect 9040 5860 9080 5900
rect 9040 5760 9080 5800
rect 9040 5660 9080 5700
rect 9040 5560 9080 5600
rect 9040 5460 9080 5500
rect 9220 5960 9260 6000
rect 9220 5860 9260 5900
rect 9220 5760 9260 5800
rect 9220 5660 9260 5700
rect 9220 5560 9260 5600
rect 9220 5460 9260 5500
rect 9400 5960 9440 6000
rect 9400 5860 9440 5900
rect 9400 5760 9440 5800
rect 9400 5660 9440 5700
rect 9400 5560 9440 5600
rect 9400 5460 9440 5500
rect 9580 5960 9620 6000
rect 9580 5860 9620 5900
rect 9580 5760 9620 5800
rect 9580 5660 9620 5700
rect 9580 5560 9620 5600
rect 9580 5460 9620 5500
rect 9760 5960 9800 6000
rect 9760 5860 9800 5900
rect 9760 5760 9800 5800
rect 9760 5660 9800 5700
rect 9760 5560 9800 5600
rect 9760 5460 9800 5500
rect 10380 5760 10420 5800
rect 10380 5660 10420 5700
rect 10490 5760 10530 5800
rect 10490 5660 10530 5700
rect 10600 5760 10640 5800
rect 10600 5660 10640 5700
rect 10710 5760 10750 5800
rect 10710 5660 10750 5700
rect 10820 5760 10860 5800
rect 10820 5660 10860 5700
rect 5420 4580 5460 4620
rect 5420 4480 5460 4520
rect 5540 4580 5580 4620
rect 5540 4480 5580 4520
rect 5660 4580 5700 4620
rect 5660 4480 5700 4520
rect 5780 4580 5820 4620
rect 5780 4480 5820 4520
rect 5900 4580 5940 4620
rect 5900 4480 5940 4520
rect 6020 4580 6060 4620
rect 6020 4480 6060 4520
rect 6140 4580 6180 4620
rect 6140 4480 6180 4520
rect 6260 4580 6300 4620
rect 6260 4480 6300 4520
rect 6380 4580 6420 4620
rect 6380 4480 6420 4520
rect 6500 4580 6540 4620
rect 6500 4480 6540 4520
rect 6620 4580 6660 4620
rect 6620 4480 6660 4520
rect 6740 4580 6780 4620
rect 6740 4480 6780 4520
rect 6860 4580 6900 4620
rect 6860 4480 6900 4520
rect 6980 4580 7020 4620
rect 6980 4480 7020 4520
rect 7100 4580 7140 4620
rect 7100 4480 7140 4520
rect 7220 4580 7260 4620
rect 7220 4480 7260 4520
rect 7340 4580 7380 4620
rect 7340 4480 7380 4520
rect 7460 4580 7500 4620
rect 7460 4480 7500 4520
rect 7580 4580 7620 4620
rect 7580 4480 7620 4520
rect 7700 4580 7740 4620
rect 7700 4480 7740 4520
rect 7820 4580 7860 4620
rect 7820 4480 7860 4520
rect 8460 4580 8500 4620
rect 8460 4480 8500 4520
rect 8580 4580 8620 4620
rect 8580 4480 8620 4520
rect 8700 4580 8740 4620
rect 8700 4480 8740 4520
rect 8820 4580 8860 4620
rect 8820 4480 8860 4520
rect 8940 4580 8980 4620
rect 8940 4480 8980 4520
rect 9060 4580 9100 4620
rect 9060 4480 9100 4520
rect 9180 4580 9220 4620
rect 9180 4480 9220 4520
rect 9300 4580 9340 4620
rect 9300 4480 9340 4520
rect 9420 4580 9460 4620
rect 9420 4480 9460 4520
rect 9540 4580 9580 4620
rect 9540 4480 9580 4520
rect 9660 4580 9700 4620
rect 9660 4480 9700 4520
rect 9780 4580 9820 4620
rect 9780 4480 9820 4520
rect 9900 4580 9940 4620
rect 9900 4480 9940 4520
rect 10020 4580 10060 4620
rect 10020 4480 10060 4520
rect 10140 4580 10180 4620
rect 10140 4480 10180 4520
rect 10260 4580 10300 4620
rect 10260 4480 10300 4520
rect 10380 4580 10420 4620
rect 10380 4480 10420 4520
rect 10500 4580 10540 4620
rect 10500 4480 10540 4520
rect 10620 4580 10660 4620
rect 10620 4480 10660 4520
rect 10740 4580 10780 4620
rect 10740 4480 10780 4520
rect 10860 4580 10900 4620
rect 10860 4480 10900 4520
rect 36090 3786 36130 3930
rect 36200 3786 36240 3930
rect 36310 3786 36350 3930
rect 36420 3786 36460 3930
rect 36530 3786 36570 3930
rect 36640 3786 36680 3930
rect 36750 3786 36790 3930
rect 37370 3890 37410 3930
rect 37370 3790 37410 3830
rect 37480 3890 37520 3930
rect 37480 3790 37520 3830
rect 37590 3890 37630 3930
rect 37590 3790 37630 3830
rect 37700 3890 37740 3930
rect 37700 3790 37740 3830
rect 37810 3890 37850 3930
rect 37810 3790 37850 3830
rect 37920 3890 37960 3930
rect 37920 3790 37960 3830
rect 38030 3890 38070 3930
rect 38030 3790 38070 3830
rect 38140 3890 38180 3930
rect 38140 3790 38180 3830
rect 38250 3890 38290 3930
rect 38250 3790 38290 3830
rect 38360 3890 38400 3930
rect 38360 3790 38400 3830
rect 38470 3890 38510 3930
rect 38470 3790 38510 3830
rect 38580 3890 38620 3930
rect 38580 3790 38620 3830
rect 38690 3890 38730 3930
rect 38690 3790 38730 3830
rect 39530 3790 39570 3930
rect 39640 3790 39680 3930
rect 39750 3790 39790 3930
rect 39860 3790 39900 3930
rect 39970 3790 40010 3930
rect 40080 3790 40120 3930
rect 40190 3790 40230 3930
rect 35450 2760 35490 2800
rect 35450 2660 35490 2700
rect 35560 2760 35600 2800
rect 35560 2660 35600 2700
rect 35670 2760 35710 2800
rect 35670 2660 35710 2700
rect 35780 2760 35820 2800
rect 35780 2660 35820 2700
rect 35890 2760 35930 2800
rect 35890 2660 35930 2700
rect 36520 2960 36560 3000
rect 36520 2860 36560 2900
rect 36520 2760 36560 2800
rect 36520 2660 36560 2700
rect 36520 2560 36560 2600
rect 36520 2460 36560 2500
rect 36700 2960 36740 3000
rect 36700 2860 36740 2900
rect 36700 2760 36740 2800
rect 36700 2660 36740 2700
rect 36700 2560 36740 2600
rect 36700 2460 36740 2500
rect 36880 2960 36920 3000
rect 36880 2860 36920 2900
rect 36880 2760 36920 2800
rect 36880 2660 36920 2700
rect 36880 2560 36920 2600
rect 36880 2460 36920 2500
rect 37060 2960 37100 3000
rect 37060 2860 37100 2900
rect 37060 2760 37100 2800
rect 37060 2660 37100 2700
rect 37060 2560 37100 2600
rect 37060 2460 37100 2500
rect 37240 2960 37280 3000
rect 37240 2860 37280 2900
rect 37240 2760 37280 2800
rect 37240 2660 37280 2700
rect 37240 2560 37280 2600
rect 37240 2460 37280 2500
rect 37420 2960 37460 3000
rect 37420 2860 37460 2900
rect 37420 2760 37460 2800
rect 37420 2660 37460 2700
rect 37420 2560 37460 2600
rect 37420 2460 37460 2500
rect 37600 2960 37640 3000
rect 37600 2860 37640 2900
rect 37600 2760 37640 2800
rect 37600 2660 37640 2700
rect 37600 2560 37640 2600
rect 37600 2460 37640 2500
rect 37780 2960 37820 3000
rect 37780 2860 37820 2900
rect 37780 2760 37820 2800
rect 37780 2660 37820 2700
rect 37780 2560 37820 2600
rect 37780 2460 37820 2500
rect 37960 2960 38000 3000
rect 37960 2860 38000 2900
rect 37960 2760 38000 2800
rect 37960 2660 38000 2700
rect 37960 2560 38000 2600
rect 37960 2460 38000 2500
rect 38140 2960 38180 3000
rect 38140 2860 38180 2900
rect 38140 2760 38180 2800
rect 38140 2660 38180 2700
rect 38140 2560 38180 2600
rect 38140 2460 38180 2500
rect 38320 2960 38360 3000
rect 38320 2860 38360 2900
rect 38320 2760 38360 2800
rect 38320 2660 38360 2700
rect 38320 2560 38360 2600
rect 38320 2460 38360 2500
rect 38500 2960 38540 3000
rect 38500 2860 38540 2900
rect 38500 2760 38540 2800
rect 38500 2660 38540 2700
rect 38500 2560 38540 2600
rect 38500 2460 38540 2500
rect 38680 2960 38720 3000
rect 38680 2860 38720 2900
rect 38680 2760 38720 2800
rect 38680 2660 38720 2700
rect 38680 2560 38720 2600
rect 38680 2460 38720 2500
rect 38860 2960 38900 3000
rect 38860 2860 38900 2900
rect 38860 2760 38900 2800
rect 38860 2660 38900 2700
rect 38860 2560 38900 2600
rect 38860 2460 38900 2500
rect 39040 2960 39080 3000
rect 39040 2860 39080 2900
rect 39040 2760 39080 2800
rect 39040 2660 39080 2700
rect 39040 2560 39080 2600
rect 39040 2460 39080 2500
rect 39220 2960 39260 3000
rect 39220 2860 39260 2900
rect 39220 2760 39260 2800
rect 39220 2660 39260 2700
rect 39220 2560 39260 2600
rect 39220 2460 39260 2500
rect 39400 2960 39440 3000
rect 39400 2860 39440 2900
rect 39400 2760 39440 2800
rect 39400 2660 39440 2700
rect 39400 2560 39440 2600
rect 39400 2460 39440 2500
rect 39580 2960 39620 3000
rect 39580 2860 39620 2900
rect 39580 2760 39620 2800
rect 39580 2660 39620 2700
rect 39580 2560 39620 2600
rect 39580 2460 39620 2500
rect 39760 2960 39800 3000
rect 39760 2860 39800 2900
rect 39760 2760 39800 2800
rect 39760 2660 39800 2700
rect 39760 2560 39800 2600
rect 39760 2460 39800 2500
rect 40380 2760 40420 2800
rect 40380 2660 40420 2700
rect 40490 2760 40530 2800
rect 40490 2660 40530 2700
rect 40600 2760 40640 2800
rect 40600 2660 40640 2700
rect 40710 2760 40750 2800
rect 40710 2660 40750 2700
rect 40820 2760 40860 2800
rect 40820 2660 40860 2700
rect 35420 1580 35460 1620
rect 35420 1480 35460 1520
rect 35540 1580 35580 1620
rect 35540 1480 35580 1520
rect 35660 1580 35700 1620
rect 35660 1480 35700 1520
rect 35780 1580 35820 1620
rect 35780 1480 35820 1520
rect 35900 1580 35940 1620
rect 35900 1480 35940 1520
rect 36020 1580 36060 1620
rect 36020 1480 36060 1520
rect 36140 1580 36180 1620
rect 36140 1480 36180 1520
rect 36260 1580 36300 1620
rect 36260 1480 36300 1520
rect 36380 1580 36420 1620
rect 36380 1480 36420 1520
rect 36500 1580 36540 1620
rect 36500 1480 36540 1520
rect 36620 1580 36660 1620
rect 36620 1480 36660 1520
rect 36740 1580 36780 1620
rect 36740 1480 36780 1520
rect 36860 1580 36900 1620
rect 36860 1480 36900 1520
rect 36980 1580 37020 1620
rect 36980 1480 37020 1520
rect 37100 1580 37140 1620
rect 37100 1480 37140 1520
rect 37220 1580 37260 1620
rect 37220 1480 37260 1520
rect 37340 1580 37380 1620
rect 37340 1480 37380 1520
rect 37460 1580 37500 1620
rect 37460 1480 37500 1520
rect 37580 1580 37620 1620
rect 37580 1480 37620 1520
rect 37700 1580 37740 1620
rect 37700 1480 37740 1520
rect 37820 1580 37860 1620
rect 37820 1480 37860 1520
rect 38460 1580 38500 1620
rect 38460 1480 38500 1520
rect 38580 1580 38620 1620
rect 38580 1480 38620 1520
rect 38700 1580 38740 1620
rect 38700 1480 38740 1520
rect 38820 1580 38860 1620
rect 38820 1480 38860 1520
rect 38940 1580 38980 1620
rect 38940 1480 38980 1520
rect 39060 1580 39100 1620
rect 39060 1480 39100 1520
rect 39180 1580 39220 1620
rect 39180 1480 39220 1520
rect 39300 1580 39340 1620
rect 39300 1480 39340 1520
rect 39420 1580 39460 1620
rect 39420 1480 39460 1520
rect 39540 1580 39580 1620
rect 39540 1480 39580 1520
rect 39660 1580 39700 1620
rect 39660 1480 39700 1520
rect 39780 1580 39820 1620
rect 39780 1480 39820 1520
rect 39900 1580 39940 1620
rect 39900 1480 39940 1520
rect 40020 1580 40060 1620
rect 40020 1480 40060 1520
rect 40140 1580 40180 1620
rect 40140 1480 40180 1520
rect 40260 1580 40300 1620
rect 40260 1480 40300 1520
rect 40380 1580 40420 1620
rect 40380 1480 40420 1520
rect 40500 1580 40540 1620
rect 40500 1480 40540 1520
rect 40620 1580 40660 1620
rect 40620 1480 40660 1520
rect 40740 1580 40780 1620
rect 40740 1480 40780 1520
rect 40860 1580 40900 1620
rect 40860 1480 40900 1520
rect 33972 -4636 34006 -4602
rect 34062 -4636 34096 -4602
rect 34152 -4636 34186 -4602
rect 34242 -4636 34276 -4602
rect 34332 -4636 34366 -4602
rect 34422 -4636 34456 -4602
rect 34512 -4636 34546 -4602
rect 33972 -4726 34006 -4692
rect 34062 -4726 34096 -4692
rect 34152 -4726 34186 -4692
rect 34242 -4726 34276 -4692
rect 34332 -4726 34366 -4692
rect 34422 -4726 34456 -4692
rect 34512 -4726 34546 -4692
rect 33972 -4816 34006 -4782
rect 34062 -4816 34096 -4782
rect 34152 -4816 34186 -4782
rect 34242 -4816 34276 -4782
rect 34332 -4816 34366 -4782
rect 34422 -4816 34456 -4782
rect 34512 -4816 34546 -4782
rect 33972 -4906 34006 -4872
rect 34062 -4906 34096 -4872
rect 34152 -4906 34186 -4872
rect 34242 -4906 34276 -4872
rect 34332 -4906 34366 -4872
rect 34422 -4906 34456 -4872
rect 34512 -4906 34546 -4872
rect 33972 -4996 34006 -4962
rect 34062 -4996 34096 -4962
rect 34152 -4996 34186 -4962
rect 34242 -4996 34276 -4962
rect 34332 -4996 34366 -4962
rect 34422 -4996 34456 -4962
rect 34512 -4996 34546 -4962
rect 33972 -5086 34006 -5052
rect 34062 -5086 34096 -5052
rect 34152 -5086 34186 -5052
rect 34242 -5086 34276 -5052
rect 34332 -5086 34366 -5052
rect 34422 -5086 34456 -5052
rect 34512 -5086 34546 -5052
rect 33972 -5176 34006 -5142
rect 34062 -5176 34096 -5142
rect 34152 -5176 34186 -5142
rect 34242 -5176 34276 -5142
rect 34332 -5176 34366 -5142
rect 34422 -5176 34456 -5142
rect 34512 -5176 34546 -5142
rect 35332 -4636 35366 -4602
rect 35422 -4636 35456 -4602
rect 35512 -4636 35546 -4602
rect 35602 -4636 35636 -4602
rect 35692 -4636 35726 -4602
rect 35782 -4636 35816 -4602
rect 35872 -4636 35906 -4602
rect 35332 -4726 35366 -4692
rect 35422 -4726 35456 -4692
rect 35512 -4726 35546 -4692
rect 35602 -4726 35636 -4692
rect 35692 -4726 35726 -4692
rect 35782 -4726 35816 -4692
rect 35872 -4726 35906 -4692
rect 35332 -4816 35366 -4782
rect 35422 -4816 35456 -4782
rect 35512 -4816 35546 -4782
rect 35602 -4816 35636 -4782
rect 35692 -4816 35726 -4782
rect 35782 -4816 35816 -4782
rect 35872 -4816 35906 -4782
rect 35332 -4906 35366 -4872
rect 35422 -4906 35456 -4872
rect 35512 -4906 35546 -4872
rect 35602 -4906 35636 -4872
rect 35692 -4906 35726 -4872
rect 35782 -4906 35816 -4872
rect 35872 -4906 35906 -4872
rect 35332 -4996 35366 -4962
rect 35422 -4996 35456 -4962
rect 35512 -4996 35546 -4962
rect 35602 -4996 35636 -4962
rect 35692 -4996 35726 -4962
rect 35782 -4996 35816 -4962
rect 35872 -4996 35906 -4962
rect 35332 -5086 35366 -5052
rect 35422 -5086 35456 -5052
rect 35512 -5086 35546 -5052
rect 35602 -5086 35636 -5052
rect 35692 -5086 35726 -5052
rect 35782 -5086 35816 -5052
rect 35872 -5086 35906 -5052
rect 35332 -5176 35366 -5142
rect 35422 -5176 35456 -5142
rect 35512 -5176 35546 -5142
rect 35602 -5176 35636 -5142
rect 35692 -5176 35726 -5142
rect 35782 -5176 35816 -5142
rect 35872 -5176 35906 -5142
rect 36692 -4636 36726 -4602
rect 36782 -4636 36816 -4602
rect 36872 -4636 36906 -4602
rect 36962 -4636 36996 -4602
rect 37052 -4636 37086 -4602
rect 37142 -4636 37176 -4602
rect 37232 -4636 37266 -4602
rect 36692 -4726 36726 -4692
rect 36782 -4726 36816 -4692
rect 36872 -4726 36906 -4692
rect 36962 -4726 36996 -4692
rect 37052 -4726 37086 -4692
rect 37142 -4726 37176 -4692
rect 37232 -4726 37266 -4692
rect 36692 -4816 36726 -4782
rect 36782 -4816 36816 -4782
rect 36872 -4816 36906 -4782
rect 36962 -4816 36996 -4782
rect 37052 -4816 37086 -4782
rect 37142 -4816 37176 -4782
rect 37232 -4816 37266 -4782
rect 36692 -4906 36726 -4872
rect 36782 -4906 36816 -4872
rect 36872 -4906 36906 -4872
rect 36962 -4906 36996 -4872
rect 37052 -4906 37086 -4872
rect 37142 -4906 37176 -4872
rect 37232 -4906 37266 -4872
rect 36692 -4996 36726 -4962
rect 36782 -4996 36816 -4962
rect 36872 -4996 36906 -4962
rect 36962 -4996 36996 -4962
rect 37052 -4996 37086 -4962
rect 37142 -4996 37176 -4962
rect 37232 -4996 37266 -4962
rect 36692 -5086 36726 -5052
rect 36782 -5086 36816 -5052
rect 36872 -5086 36906 -5052
rect 36962 -5086 36996 -5052
rect 37052 -5086 37086 -5052
rect 37142 -5086 37176 -5052
rect 37232 -5086 37266 -5052
rect 36692 -5176 36726 -5142
rect 36782 -5176 36816 -5142
rect 36872 -5176 36906 -5142
rect 36962 -5176 36996 -5142
rect 37052 -5176 37086 -5142
rect 37142 -5176 37176 -5142
rect 37232 -5176 37266 -5142
rect 33972 -5996 34006 -5962
rect 34062 -5996 34096 -5962
rect 34152 -5996 34186 -5962
rect 34242 -5996 34276 -5962
rect 34332 -5996 34366 -5962
rect 34422 -5996 34456 -5962
rect 34512 -5996 34546 -5962
rect 33972 -6086 34006 -6052
rect 34062 -6086 34096 -6052
rect 34152 -6086 34186 -6052
rect 34242 -6086 34276 -6052
rect 34332 -6086 34366 -6052
rect 34422 -6086 34456 -6052
rect 34512 -6086 34546 -6052
rect 33972 -6176 34006 -6142
rect 34062 -6176 34096 -6142
rect 34152 -6176 34186 -6142
rect 34242 -6176 34276 -6142
rect 34332 -6176 34366 -6142
rect 34422 -6176 34456 -6142
rect 34512 -6176 34546 -6142
rect 33972 -6266 34006 -6232
rect 34062 -6266 34096 -6232
rect 34152 -6266 34186 -6232
rect 34242 -6266 34276 -6232
rect 34332 -6266 34366 -6232
rect 34422 -6266 34456 -6232
rect 34512 -6266 34546 -6232
rect 33972 -6356 34006 -6322
rect 34062 -6356 34096 -6322
rect 34152 -6356 34186 -6322
rect 34242 -6356 34276 -6322
rect 34332 -6356 34366 -6322
rect 34422 -6356 34456 -6322
rect 34512 -6356 34546 -6322
rect 33972 -6446 34006 -6412
rect 34062 -6446 34096 -6412
rect 34152 -6446 34186 -6412
rect 34242 -6446 34276 -6412
rect 34332 -6446 34366 -6412
rect 34422 -6446 34456 -6412
rect 34512 -6446 34546 -6412
rect 33972 -6536 34006 -6502
rect 34062 -6536 34096 -6502
rect 34152 -6536 34186 -6502
rect 34242 -6536 34276 -6502
rect 34332 -6536 34366 -6502
rect 34422 -6536 34456 -6502
rect 34512 -6536 34546 -6502
rect 35332 -5996 35366 -5962
rect 35422 -5996 35456 -5962
rect 35512 -5996 35546 -5962
rect 35602 -5996 35636 -5962
rect 35692 -5996 35726 -5962
rect 35782 -5996 35816 -5962
rect 35872 -5996 35906 -5962
rect 35332 -6086 35366 -6052
rect 35422 -6086 35456 -6052
rect 35512 -6086 35546 -6052
rect 35602 -6086 35636 -6052
rect 35692 -6086 35726 -6052
rect 35782 -6086 35816 -6052
rect 35872 -6086 35906 -6052
rect 35332 -6176 35366 -6142
rect 35422 -6176 35456 -6142
rect 35512 -6176 35546 -6142
rect 35602 -6176 35636 -6142
rect 35692 -6176 35726 -6142
rect 35782 -6176 35816 -6142
rect 35872 -6176 35906 -6142
rect 35332 -6266 35366 -6232
rect 35422 -6266 35456 -6232
rect 35512 -6266 35546 -6232
rect 35602 -6266 35636 -6232
rect 35692 -6266 35726 -6232
rect 35782 -6266 35816 -6232
rect 35872 -6266 35906 -6232
rect 35332 -6356 35366 -6322
rect 35422 -6356 35456 -6322
rect 35512 -6356 35546 -6322
rect 35602 -6356 35636 -6322
rect 35692 -6356 35726 -6322
rect 35782 -6356 35816 -6322
rect 35872 -6356 35906 -6322
rect 35332 -6446 35366 -6412
rect 35422 -6446 35456 -6412
rect 35512 -6446 35546 -6412
rect 35602 -6446 35636 -6412
rect 35692 -6446 35726 -6412
rect 35782 -6446 35816 -6412
rect 35872 -6446 35906 -6412
rect 35332 -6536 35366 -6502
rect 35422 -6536 35456 -6502
rect 35512 -6536 35546 -6502
rect 35602 -6536 35636 -6502
rect 35692 -6536 35726 -6502
rect 35782 -6536 35816 -6502
rect 35872 -6536 35906 -6502
rect 36692 -5996 36726 -5962
rect 36782 -5996 36816 -5962
rect 36872 -5996 36906 -5962
rect 36962 -5996 36996 -5962
rect 37052 -5996 37086 -5962
rect 37142 -5996 37176 -5962
rect 37232 -5996 37266 -5962
rect 36692 -6086 36726 -6052
rect 36782 -6086 36816 -6052
rect 36872 -6086 36906 -6052
rect 36962 -6086 36996 -6052
rect 37052 -6086 37086 -6052
rect 37142 -6086 37176 -6052
rect 37232 -6086 37266 -6052
rect 36692 -6176 36726 -6142
rect 36782 -6176 36816 -6142
rect 36872 -6176 36906 -6142
rect 36962 -6176 36996 -6142
rect 37052 -6176 37086 -6142
rect 37142 -6176 37176 -6142
rect 37232 -6176 37266 -6142
rect 36692 -6266 36726 -6232
rect 36782 -6266 36816 -6232
rect 36872 -6266 36906 -6232
rect 36962 -6266 36996 -6232
rect 37052 -6266 37086 -6232
rect 37142 -6266 37176 -6232
rect 37232 -6266 37266 -6232
rect 36692 -6356 36726 -6322
rect 36782 -6356 36816 -6322
rect 36872 -6356 36906 -6322
rect 36962 -6356 36996 -6322
rect 37052 -6356 37086 -6322
rect 37142 -6356 37176 -6322
rect 37232 -6356 37266 -6322
rect 36692 -6446 36726 -6412
rect 36782 -6446 36816 -6412
rect 36872 -6446 36906 -6412
rect 36962 -6446 36996 -6412
rect 37052 -6446 37086 -6412
rect 37142 -6446 37176 -6412
rect 37232 -6446 37266 -6412
rect 36692 -6536 36726 -6502
rect 36782 -6536 36816 -6502
rect 36872 -6536 36906 -6502
rect 36962 -6536 36996 -6502
rect 37052 -6536 37086 -6502
rect 37142 -6536 37176 -6502
rect 37232 -6536 37266 -6502
rect 33972 -7356 34006 -7322
rect 34062 -7356 34096 -7322
rect 34152 -7356 34186 -7322
rect 34242 -7356 34276 -7322
rect 34332 -7356 34366 -7322
rect 34422 -7356 34456 -7322
rect 34512 -7356 34546 -7322
rect 33972 -7446 34006 -7412
rect 34062 -7446 34096 -7412
rect 34152 -7446 34186 -7412
rect 34242 -7446 34276 -7412
rect 34332 -7446 34366 -7412
rect 34422 -7446 34456 -7412
rect 34512 -7446 34546 -7412
rect 33972 -7536 34006 -7502
rect 34062 -7536 34096 -7502
rect 34152 -7536 34186 -7502
rect 34242 -7536 34276 -7502
rect 34332 -7536 34366 -7502
rect 34422 -7536 34456 -7502
rect 34512 -7536 34546 -7502
rect 33972 -7626 34006 -7592
rect 34062 -7626 34096 -7592
rect 34152 -7626 34186 -7592
rect 34242 -7626 34276 -7592
rect 34332 -7626 34366 -7592
rect 34422 -7626 34456 -7592
rect 34512 -7626 34546 -7592
rect 33972 -7716 34006 -7682
rect 34062 -7716 34096 -7682
rect 34152 -7716 34186 -7682
rect 34242 -7716 34276 -7682
rect 34332 -7716 34366 -7682
rect 34422 -7716 34456 -7682
rect 34512 -7716 34546 -7682
rect 33972 -7806 34006 -7772
rect 34062 -7806 34096 -7772
rect 34152 -7806 34186 -7772
rect 34242 -7806 34276 -7772
rect 34332 -7806 34366 -7772
rect 34422 -7806 34456 -7772
rect 34512 -7806 34546 -7772
rect 33972 -7896 34006 -7862
rect 34062 -7896 34096 -7862
rect 34152 -7896 34186 -7862
rect 34242 -7896 34276 -7862
rect 34332 -7896 34366 -7862
rect 34422 -7896 34456 -7862
rect 34512 -7896 34546 -7862
rect 35332 -7356 35366 -7322
rect 35422 -7356 35456 -7322
rect 35512 -7356 35546 -7322
rect 35602 -7356 35636 -7322
rect 35692 -7356 35726 -7322
rect 35782 -7356 35816 -7322
rect 35872 -7356 35906 -7322
rect 35332 -7446 35366 -7412
rect 35422 -7446 35456 -7412
rect 35512 -7446 35546 -7412
rect 35602 -7446 35636 -7412
rect 35692 -7446 35726 -7412
rect 35782 -7446 35816 -7412
rect 35872 -7446 35906 -7412
rect 35332 -7536 35366 -7502
rect 35422 -7536 35456 -7502
rect 35512 -7536 35546 -7502
rect 35602 -7536 35636 -7502
rect 35692 -7536 35726 -7502
rect 35782 -7536 35816 -7502
rect 35872 -7536 35906 -7502
rect 35332 -7626 35366 -7592
rect 35422 -7626 35456 -7592
rect 35512 -7626 35546 -7592
rect 35602 -7626 35636 -7592
rect 35692 -7626 35726 -7592
rect 35782 -7626 35816 -7592
rect 35872 -7626 35906 -7592
rect 35332 -7716 35366 -7682
rect 35422 -7716 35456 -7682
rect 35512 -7716 35546 -7682
rect 35602 -7716 35636 -7682
rect 35692 -7716 35726 -7682
rect 35782 -7716 35816 -7682
rect 35872 -7716 35906 -7682
rect 35332 -7806 35366 -7772
rect 35422 -7806 35456 -7772
rect 35512 -7806 35546 -7772
rect 35602 -7806 35636 -7772
rect 35692 -7806 35726 -7772
rect 35782 -7806 35816 -7772
rect 35872 -7806 35906 -7772
rect 35332 -7896 35366 -7862
rect 35422 -7896 35456 -7862
rect 35512 -7896 35546 -7862
rect 35602 -7896 35636 -7862
rect 35692 -7896 35726 -7862
rect 35782 -7896 35816 -7862
rect 35872 -7896 35906 -7862
rect 36692 -7356 36726 -7322
rect 36782 -7356 36816 -7322
rect 36872 -7356 36906 -7322
rect 36962 -7356 36996 -7322
rect 37052 -7356 37086 -7322
rect 37142 -7356 37176 -7322
rect 37232 -7356 37266 -7322
rect 36692 -7446 36726 -7412
rect 36782 -7446 36816 -7412
rect 36872 -7446 36906 -7412
rect 36962 -7446 36996 -7412
rect 37052 -7446 37086 -7412
rect 37142 -7446 37176 -7412
rect 37232 -7446 37266 -7412
rect 36692 -7536 36726 -7502
rect 36782 -7536 36816 -7502
rect 36872 -7536 36906 -7502
rect 36962 -7536 36996 -7502
rect 37052 -7536 37086 -7502
rect 37142 -7536 37176 -7502
rect 37232 -7536 37266 -7502
rect 36692 -7626 36726 -7592
rect 36782 -7626 36816 -7592
rect 36872 -7626 36906 -7592
rect 36962 -7626 36996 -7592
rect 37052 -7626 37086 -7592
rect 37142 -7626 37176 -7592
rect 37232 -7626 37266 -7592
rect 36692 -7716 36726 -7682
rect 36782 -7716 36816 -7682
rect 36872 -7716 36906 -7682
rect 36962 -7716 36996 -7682
rect 37052 -7716 37086 -7682
rect 37142 -7716 37176 -7682
rect 37232 -7716 37266 -7682
rect 36692 -7806 36726 -7772
rect 36782 -7806 36816 -7772
rect 36872 -7806 36906 -7772
rect 36962 -7806 36996 -7772
rect 37052 -7806 37086 -7772
rect 37142 -7806 37176 -7772
rect 37232 -7806 37266 -7772
rect 36692 -7896 36726 -7862
rect 36782 -7896 36816 -7862
rect 36872 -7896 36906 -7862
rect 36962 -7896 36996 -7862
rect 37052 -7896 37086 -7862
rect 37142 -7896 37176 -7862
rect 37232 -7896 37266 -7862
<< psubdiff >>
rect 50 7280 1180 7320
rect 1340 7280 2470 7320
rect 50 7160 90 7280
rect 2430 7160 2470 7280
rect 50 6890 90 7000
rect 2430 6890 2470 7000
rect 50 6850 1180 6890
rect 1340 6850 2470 6890
rect 2620 7010 3690 7050
rect 3850 7010 5010 7050
rect 50 6750 1150 6790
rect 1310 6750 2410 6790
rect 50 6630 90 6750
rect 2370 6630 2410 6750
rect 50 6360 90 6470
rect 2370 6360 2410 6470
rect 50 6320 1150 6360
rect 1310 6320 2410 6360
rect 2620 6650 2660 7010
rect 4970 6650 5010 7010
rect 440 6220 1150 6260
rect 1310 6220 2040 6260
rect 440 6160 480 6220
rect 2000 6160 2040 6220
rect 440 5940 480 6000
rect 2620 6140 2660 6490
rect 4970 6140 5010 6490
rect 2620 6100 3690 6140
rect 3850 6100 5010 6140
rect 2000 5940 2040 6000
rect 440 5900 1150 5940
rect 1310 5900 2040 5940
rect 2950 6000 3690 6040
rect 3850 6000 4600 6040
rect 2950 5940 2990 6000
rect 440 5800 1150 5840
rect 1310 5800 2040 5840
rect 440 5740 480 5800
rect 2000 5740 2040 5800
rect 440 5520 480 5580
rect 4560 5940 4600 6000
rect 2950 5730 2990 5780
rect 4560 5730 4600 5780
rect 2950 5690 3690 5730
rect 3850 5690 4600 5730
rect 2000 5520 2040 5580
rect 440 5480 1150 5520
rect 1310 5480 2040 5520
rect 6160 4140 6820 4180
rect 6980 4140 7640 4180
rect 6160 3930 6200 4140
rect 7600 3930 7640 4140
rect 6160 3650 6200 3770
rect 7600 3650 7640 3770
rect 6160 3610 6820 3650
rect 6980 3610 7640 3650
rect 8680 4140 9340 4180
rect 9500 4140 10160 4180
rect 8680 3930 8720 4140
rect 10120 3930 10160 4140
rect 8680 3650 8720 3770
rect 10120 3650 10160 3770
rect 8680 3610 10160 3650
rect 5680 3490 6820 3530
rect 6980 3490 8120 3530
rect -100 3430 200 3460
rect -100 3390 -70 3430
rect -30 3390 30 3430
rect 70 3390 130 3430
rect 170 3390 200 3430
rect -100 3360 200 3390
rect 5680 3180 5720 3490
rect 5680 2700 5720 3020
rect 8080 3180 8120 3490
rect 8080 2700 8120 3020
rect 5680 2660 6820 2700
rect 6980 2660 8120 2700
rect 8200 3490 9340 3530
rect 9500 3490 10640 3530
rect 8200 3180 8240 3490
rect 8200 2700 8240 3020
rect 10600 3180 10640 3490
rect 10600 2700 10640 3020
rect 8200 2660 9340 2700
rect 9500 2660 10640 2700
rect 5880 2560 8080 2600
rect 8240 2560 10430 2600
rect 5880 2390 5920 2560
rect 5880 2150 5920 2230
rect 10390 2390 10430 2560
rect 10390 2150 10430 2230
rect 5880 2110 8080 2150
rect 8240 2110 10430 2150
rect 6240 2010 6800 2050
rect 6960 2010 7400 2050
rect 6240 1840 6280 2010
rect 6240 1510 6280 1680
rect 7360 1840 7400 2010
rect 7360 1510 7400 1680
rect 6240 1470 7400 1510
rect 7470 2010 8080 2050
rect 8240 2010 8850 2050
rect 7470 1840 7510 2010
rect 7470 1510 7510 1680
rect 8810 1840 8850 2010
rect 8810 1510 8850 1680
rect 7470 1470 8080 1510
rect 8240 1470 8850 1510
rect 8920 2010 9360 2050
rect 9520 2010 10080 2050
rect 8920 1840 8960 2010
rect 8920 1510 8960 1680
rect 10040 1840 10080 2010
rect 10040 1510 10080 1680
rect 8920 1470 10080 1510
rect 36160 1140 36820 1180
rect 36980 1140 37640 1180
rect 36160 930 36200 1140
rect 37600 930 37640 1140
rect 36160 650 36200 770
rect 37600 650 37640 770
rect 36160 610 36820 650
rect 36980 610 37640 650
rect 38680 1140 39340 1180
rect 39500 1140 40160 1180
rect 38680 930 38720 1140
rect 40120 930 40160 1140
rect 38680 650 38720 770
rect 40120 650 40160 770
rect 38680 610 40160 650
rect 35680 490 36820 530
rect 36980 490 38120 530
rect 35680 180 35720 490
rect 35680 -300 35720 20
rect 38080 180 38120 490
rect 38080 -300 38120 20
rect 35680 -340 36820 -300
rect 36980 -340 38120 -300
rect 38200 490 39340 530
rect 39500 490 40640 530
rect 38200 180 38240 490
rect 38200 -300 38240 20
rect 40600 180 40640 490
rect 40600 -300 40640 20
rect 38200 -340 39340 -300
rect 39500 -340 40640 -300
rect 35880 -440 38080 -400
rect 38240 -440 40430 -400
rect 35880 -610 35920 -440
rect 35880 -850 35920 -770
rect 40390 -610 40430 -440
rect 40390 -850 40430 -770
rect 35880 -890 38080 -850
rect 38240 -890 40430 -850
rect 36240 -990 36800 -950
rect 36960 -990 37400 -950
rect 36240 -1160 36280 -990
rect 36240 -1490 36280 -1320
rect 37360 -1160 37400 -990
rect 37360 -1490 37400 -1320
rect 36240 -1530 37400 -1490
rect 37470 -990 38080 -950
rect 38240 -990 38850 -950
rect 37470 -1160 37510 -990
rect 37470 -1490 37510 -1320
rect 38810 -1160 38850 -990
rect 38810 -1490 38850 -1320
rect 37470 -1530 38080 -1490
rect 38240 -1530 38850 -1490
rect 38920 -990 39360 -950
rect 39520 -990 40080 -950
rect 38920 -1160 38960 -990
rect 38920 -1490 38960 -1320
rect 40040 -1160 40080 -990
rect 40040 -1490 40080 -1320
rect 38920 -1530 40080 -1490
rect 44050 -2720 45180 -2680
rect 45340 -2720 46470 -2680
rect 44050 -2840 44090 -2720
rect 46430 -2840 46470 -2720
rect 44050 -3110 44090 -3000
rect 46430 -3110 46470 -3000
rect 44050 -3150 45180 -3110
rect 45340 -3150 46470 -3110
rect 46620 -2990 47690 -2950
rect 47850 -2990 49010 -2950
rect 44050 -3250 45150 -3210
rect 45310 -3250 46410 -3210
rect 44050 -3370 44090 -3250
rect 46370 -3370 46410 -3250
rect 44050 -3640 44090 -3530
rect 46370 -3640 46410 -3530
rect 44050 -3680 45150 -3640
rect 45310 -3680 46410 -3640
rect 46620 -3350 46660 -2990
rect 48970 -3350 49010 -2990
rect 44440 -3780 45150 -3740
rect 45310 -3780 46040 -3740
rect 44440 -3840 44480 -3780
rect 46000 -3840 46040 -3780
rect 44440 -4060 44480 -4000
rect 46620 -3860 46660 -3510
rect 48970 -3860 49010 -3510
rect 46620 -3900 47690 -3860
rect 47850 -3900 49010 -3860
rect 46000 -4060 46040 -4000
rect 44440 -4100 45150 -4060
rect 45310 -4100 46040 -4060
rect 46950 -4000 47690 -3960
rect 47850 -4000 48600 -3960
rect 46950 -4060 46990 -4000
rect 44440 -4200 45150 -4160
rect 45310 -4200 46040 -4160
rect 33616 -4279 34904 -4246
rect 33616 -4313 33674 -4279
rect 33708 -4313 33764 -4279
rect 33798 -4313 33854 -4279
rect 33888 -4313 33944 -4279
rect 33978 -4313 34034 -4279
rect 34068 -4313 34124 -4279
rect 34158 -4313 34214 -4279
rect 34248 -4313 34304 -4279
rect 34338 -4313 34394 -4279
rect 34428 -4313 34484 -4279
rect 34518 -4313 34574 -4279
rect 34608 -4313 34664 -4279
rect 34698 -4313 34754 -4279
rect 34788 -4313 34904 -4279
rect 33616 -4347 34904 -4313
rect 33616 -4380 33717 -4347
rect 33616 -4414 33651 -4380
rect 33685 -4414 33717 -4380
rect 34803 -4380 34904 -4347
rect 33616 -4470 33717 -4414
rect 33616 -4504 33651 -4470
rect 33685 -4504 33717 -4470
rect 33616 -4560 33717 -4504
rect 33616 -4594 33651 -4560
rect 33685 -4594 33717 -4560
rect 33616 -4650 33717 -4594
rect 33616 -4684 33651 -4650
rect 33685 -4684 33717 -4650
rect 33616 -4740 33717 -4684
rect 33616 -4774 33651 -4740
rect 33685 -4774 33717 -4740
rect 33616 -4830 33717 -4774
rect 33616 -4864 33651 -4830
rect 33685 -4864 33717 -4830
rect 33616 -4920 33717 -4864
rect 33616 -4954 33651 -4920
rect 33685 -4954 33717 -4920
rect 33616 -5010 33717 -4954
rect 33616 -5044 33651 -5010
rect 33685 -5044 33717 -5010
rect 33616 -5100 33717 -5044
rect 33616 -5134 33651 -5100
rect 33685 -5134 33717 -5100
rect 33616 -5190 33717 -5134
rect 33616 -5224 33651 -5190
rect 33685 -5224 33717 -5190
rect 33616 -5280 33717 -5224
rect 33616 -5314 33651 -5280
rect 33685 -5314 33717 -5280
rect 33616 -5370 33717 -5314
rect 33616 -5404 33651 -5370
rect 33685 -5404 33717 -5370
rect 34803 -4414 34838 -4380
rect 34872 -4414 34904 -4380
rect 34803 -4470 34904 -4414
rect 34803 -4504 34838 -4470
rect 34872 -4504 34904 -4470
rect 34803 -4560 34904 -4504
rect 34803 -4594 34838 -4560
rect 34872 -4594 34904 -4560
rect 34803 -4650 34904 -4594
rect 34803 -4684 34838 -4650
rect 34872 -4684 34904 -4650
rect 34803 -4740 34904 -4684
rect 34803 -4774 34838 -4740
rect 34872 -4774 34904 -4740
rect 34803 -4830 34904 -4774
rect 34803 -4864 34838 -4830
rect 34872 -4864 34904 -4830
rect 34803 -4920 34904 -4864
rect 34803 -4954 34838 -4920
rect 34872 -4954 34904 -4920
rect 34803 -5010 34904 -4954
rect 34803 -5044 34838 -5010
rect 34872 -5044 34904 -5010
rect 34803 -5100 34904 -5044
rect 34803 -5134 34838 -5100
rect 34872 -5134 34904 -5100
rect 34803 -5190 34904 -5134
rect 34803 -5224 34838 -5190
rect 34872 -5224 34904 -5190
rect 34803 -5280 34904 -5224
rect 34803 -5314 34838 -5280
rect 34872 -5314 34904 -5280
rect 34803 -5370 34904 -5314
rect 33616 -5433 33717 -5404
rect 34803 -5404 34838 -5370
rect 34872 -5404 34904 -5370
rect 34803 -5433 34904 -5404
rect 33616 -5466 34904 -5433
rect 33616 -5500 33674 -5466
rect 33708 -5500 33764 -5466
rect 33798 -5500 33854 -5466
rect 33888 -5500 33944 -5466
rect 33978 -5500 34034 -5466
rect 34068 -5500 34124 -5466
rect 34158 -5500 34214 -5466
rect 34248 -5500 34304 -5466
rect 34338 -5500 34394 -5466
rect 34428 -5500 34484 -5466
rect 34518 -5500 34574 -5466
rect 34608 -5500 34664 -5466
rect 34698 -5500 34754 -5466
rect 34788 -5500 34904 -5466
rect 33616 -5534 34904 -5500
rect 34976 -4279 36264 -4246
rect 34976 -4313 35034 -4279
rect 35068 -4313 35124 -4279
rect 35158 -4313 35214 -4279
rect 35248 -4313 35304 -4279
rect 35338 -4313 35394 -4279
rect 35428 -4313 35484 -4279
rect 35518 -4313 35574 -4279
rect 35608 -4313 35664 -4279
rect 35698 -4313 35754 -4279
rect 35788 -4313 35844 -4279
rect 35878 -4313 35934 -4279
rect 35968 -4313 36024 -4279
rect 36058 -4313 36114 -4279
rect 36148 -4313 36264 -4279
rect 34976 -4347 36264 -4313
rect 34976 -4380 35077 -4347
rect 34976 -4414 35011 -4380
rect 35045 -4414 35077 -4380
rect 36163 -4380 36264 -4347
rect 34976 -4470 35077 -4414
rect 34976 -4504 35011 -4470
rect 35045 -4504 35077 -4470
rect 34976 -4560 35077 -4504
rect 34976 -4594 35011 -4560
rect 35045 -4594 35077 -4560
rect 34976 -4650 35077 -4594
rect 34976 -4684 35011 -4650
rect 35045 -4684 35077 -4650
rect 34976 -4740 35077 -4684
rect 34976 -4774 35011 -4740
rect 35045 -4774 35077 -4740
rect 34976 -4830 35077 -4774
rect 34976 -4864 35011 -4830
rect 35045 -4864 35077 -4830
rect 34976 -4920 35077 -4864
rect 34976 -4954 35011 -4920
rect 35045 -4954 35077 -4920
rect 34976 -5010 35077 -4954
rect 34976 -5044 35011 -5010
rect 35045 -5044 35077 -5010
rect 34976 -5100 35077 -5044
rect 34976 -5134 35011 -5100
rect 35045 -5134 35077 -5100
rect 34976 -5190 35077 -5134
rect 34976 -5224 35011 -5190
rect 35045 -5224 35077 -5190
rect 34976 -5280 35077 -5224
rect 34976 -5314 35011 -5280
rect 35045 -5314 35077 -5280
rect 34976 -5370 35077 -5314
rect 34976 -5404 35011 -5370
rect 35045 -5404 35077 -5370
rect 36163 -4414 36198 -4380
rect 36232 -4414 36264 -4380
rect 36163 -4470 36264 -4414
rect 36163 -4504 36198 -4470
rect 36232 -4504 36264 -4470
rect 36163 -4560 36264 -4504
rect 36163 -4594 36198 -4560
rect 36232 -4594 36264 -4560
rect 36163 -4650 36264 -4594
rect 36163 -4684 36198 -4650
rect 36232 -4684 36264 -4650
rect 36163 -4740 36264 -4684
rect 36163 -4774 36198 -4740
rect 36232 -4774 36264 -4740
rect 36163 -4830 36264 -4774
rect 36163 -4864 36198 -4830
rect 36232 -4864 36264 -4830
rect 36163 -4920 36264 -4864
rect 36163 -4954 36198 -4920
rect 36232 -4954 36264 -4920
rect 36163 -5010 36264 -4954
rect 36163 -5044 36198 -5010
rect 36232 -5044 36264 -5010
rect 36163 -5100 36264 -5044
rect 36163 -5134 36198 -5100
rect 36232 -5134 36264 -5100
rect 36163 -5190 36264 -5134
rect 36163 -5224 36198 -5190
rect 36232 -5224 36264 -5190
rect 36163 -5280 36264 -5224
rect 36163 -5314 36198 -5280
rect 36232 -5314 36264 -5280
rect 36163 -5370 36264 -5314
rect 34976 -5433 35077 -5404
rect 36163 -5404 36198 -5370
rect 36232 -5404 36264 -5370
rect 36163 -5433 36264 -5404
rect 34976 -5466 36264 -5433
rect 34976 -5500 35034 -5466
rect 35068 -5500 35124 -5466
rect 35158 -5500 35214 -5466
rect 35248 -5500 35304 -5466
rect 35338 -5500 35394 -5466
rect 35428 -5500 35484 -5466
rect 35518 -5500 35574 -5466
rect 35608 -5500 35664 -5466
rect 35698 -5500 35754 -5466
rect 35788 -5500 35844 -5466
rect 35878 -5500 35934 -5466
rect 35968 -5500 36024 -5466
rect 36058 -5500 36114 -5466
rect 36148 -5500 36264 -5466
rect 34976 -5534 36264 -5500
rect 36336 -4279 37624 -4246
rect 36336 -4313 36394 -4279
rect 36428 -4313 36484 -4279
rect 36518 -4313 36574 -4279
rect 36608 -4313 36664 -4279
rect 36698 -4313 36754 -4279
rect 36788 -4313 36844 -4279
rect 36878 -4313 36934 -4279
rect 36968 -4313 37024 -4279
rect 37058 -4313 37114 -4279
rect 37148 -4313 37204 -4279
rect 37238 -4313 37294 -4279
rect 37328 -4313 37384 -4279
rect 37418 -4313 37474 -4279
rect 37508 -4313 37624 -4279
rect 36336 -4347 37624 -4313
rect 36336 -4380 36437 -4347
rect 36336 -4414 36371 -4380
rect 36405 -4414 36437 -4380
rect 37523 -4380 37624 -4347
rect 36336 -4470 36437 -4414
rect 36336 -4504 36371 -4470
rect 36405 -4504 36437 -4470
rect 36336 -4560 36437 -4504
rect 36336 -4594 36371 -4560
rect 36405 -4594 36437 -4560
rect 36336 -4650 36437 -4594
rect 36336 -4684 36371 -4650
rect 36405 -4684 36437 -4650
rect 36336 -4740 36437 -4684
rect 36336 -4774 36371 -4740
rect 36405 -4774 36437 -4740
rect 36336 -4830 36437 -4774
rect 36336 -4864 36371 -4830
rect 36405 -4864 36437 -4830
rect 36336 -4920 36437 -4864
rect 36336 -4954 36371 -4920
rect 36405 -4954 36437 -4920
rect 36336 -5010 36437 -4954
rect 36336 -5044 36371 -5010
rect 36405 -5044 36437 -5010
rect 36336 -5100 36437 -5044
rect 36336 -5134 36371 -5100
rect 36405 -5134 36437 -5100
rect 36336 -5190 36437 -5134
rect 36336 -5224 36371 -5190
rect 36405 -5224 36437 -5190
rect 36336 -5280 36437 -5224
rect 36336 -5314 36371 -5280
rect 36405 -5314 36437 -5280
rect 36336 -5370 36437 -5314
rect 36336 -5404 36371 -5370
rect 36405 -5404 36437 -5370
rect 37523 -4414 37558 -4380
rect 37592 -4414 37624 -4380
rect 37523 -4470 37624 -4414
rect 37523 -4504 37558 -4470
rect 37592 -4504 37624 -4470
rect 37523 -4560 37624 -4504
rect 44440 -4260 44480 -4200
rect 46000 -4260 46040 -4200
rect 44440 -4480 44480 -4420
rect 48560 -4060 48600 -4000
rect 46950 -4270 46990 -4220
rect 48560 -4270 48600 -4220
rect 46950 -4310 47690 -4270
rect 47850 -4310 48600 -4270
rect 46000 -4480 46040 -4420
rect 44440 -4520 45150 -4480
rect 45310 -4520 46040 -4480
rect 37523 -4594 37558 -4560
rect 37592 -4594 37624 -4560
rect 37523 -4650 37624 -4594
rect 37523 -4684 37558 -4650
rect 37592 -4684 37624 -4650
rect 37523 -4740 37624 -4684
rect 37523 -4774 37558 -4740
rect 37592 -4774 37624 -4740
rect 37523 -4830 37624 -4774
rect 37523 -4864 37558 -4830
rect 37592 -4864 37624 -4830
rect 37523 -4920 37624 -4864
rect 37523 -4954 37558 -4920
rect 37592 -4954 37624 -4920
rect 37523 -5010 37624 -4954
rect 37523 -5044 37558 -5010
rect 37592 -5044 37624 -5010
rect 37523 -5100 37624 -5044
rect 37523 -5134 37558 -5100
rect 37592 -5134 37624 -5100
rect 37523 -5190 37624 -5134
rect 37523 -5224 37558 -5190
rect 37592 -5224 37624 -5190
rect 37523 -5280 37624 -5224
rect 37523 -5314 37558 -5280
rect 37592 -5314 37624 -5280
rect 37523 -5370 37624 -5314
rect 36336 -5433 36437 -5404
rect 37523 -5404 37558 -5370
rect 37592 -5404 37624 -5370
rect 37523 -5433 37624 -5404
rect 36336 -5466 37624 -5433
rect 36336 -5500 36394 -5466
rect 36428 -5500 36484 -5466
rect 36518 -5500 36574 -5466
rect 36608 -5500 36664 -5466
rect 36698 -5500 36754 -5466
rect 36788 -5500 36844 -5466
rect 36878 -5500 36934 -5466
rect 36968 -5500 37024 -5466
rect 37058 -5500 37114 -5466
rect 37148 -5500 37204 -5466
rect 37238 -5500 37294 -5466
rect 37328 -5500 37384 -5466
rect 37418 -5500 37474 -5466
rect 37508 -5500 37624 -5466
rect 36336 -5534 37624 -5500
rect 33616 -5639 34904 -5606
rect 33616 -5673 33674 -5639
rect 33708 -5673 33764 -5639
rect 33798 -5673 33854 -5639
rect 33888 -5673 33944 -5639
rect 33978 -5673 34034 -5639
rect 34068 -5673 34124 -5639
rect 34158 -5673 34214 -5639
rect 34248 -5673 34304 -5639
rect 34338 -5673 34394 -5639
rect 34428 -5673 34484 -5639
rect 34518 -5673 34574 -5639
rect 34608 -5673 34664 -5639
rect 34698 -5673 34754 -5639
rect 34788 -5673 34904 -5639
rect 33616 -5707 34904 -5673
rect 33616 -5740 33717 -5707
rect 33616 -5774 33651 -5740
rect 33685 -5774 33717 -5740
rect 34803 -5740 34904 -5707
rect 33616 -5830 33717 -5774
rect 33616 -5864 33651 -5830
rect 33685 -5864 33717 -5830
rect 33616 -5920 33717 -5864
rect 33616 -5954 33651 -5920
rect 33685 -5954 33717 -5920
rect 33616 -6010 33717 -5954
rect 33616 -6044 33651 -6010
rect 33685 -6044 33717 -6010
rect 33616 -6100 33717 -6044
rect 33616 -6134 33651 -6100
rect 33685 -6134 33717 -6100
rect 33616 -6190 33717 -6134
rect 33616 -6224 33651 -6190
rect 33685 -6224 33717 -6190
rect 33616 -6280 33717 -6224
rect 33616 -6314 33651 -6280
rect 33685 -6314 33717 -6280
rect 33616 -6370 33717 -6314
rect 33616 -6404 33651 -6370
rect 33685 -6404 33717 -6370
rect 33616 -6460 33717 -6404
rect 33616 -6494 33651 -6460
rect 33685 -6494 33717 -6460
rect 33616 -6550 33717 -6494
rect 33616 -6584 33651 -6550
rect 33685 -6584 33717 -6550
rect 33616 -6640 33717 -6584
rect 33616 -6674 33651 -6640
rect 33685 -6674 33717 -6640
rect 33616 -6730 33717 -6674
rect 33616 -6764 33651 -6730
rect 33685 -6764 33717 -6730
rect 34803 -5774 34838 -5740
rect 34872 -5774 34904 -5740
rect 34803 -5830 34904 -5774
rect 34803 -5864 34838 -5830
rect 34872 -5864 34904 -5830
rect 34803 -5920 34904 -5864
rect 34803 -5954 34838 -5920
rect 34872 -5954 34904 -5920
rect 34803 -6010 34904 -5954
rect 34803 -6044 34838 -6010
rect 34872 -6044 34904 -6010
rect 34803 -6100 34904 -6044
rect 34803 -6134 34838 -6100
rect 34872 -6134 34904 -6100
rect 34803 -6190 34904 -6134
rect 34803 -6224 34838 -6190
rect 34872 -6224 34904 -6190
rect 34803 -6280 34904 -6224
rect 34803 -6314 34838 -6280
rect 34872 -6314 34904 -6280
rect 34803 -6370 34904 -6314
rect 34803 -6404 34838 -6370
rect 34872 -6404 34904 -6370
rect 34803 -6460 34904 -6404
rect 34803 -6494 34838 -6460
rect 34872 -6494 34904 -6460
rect 34803 -6550 34904 -6494
rect 34803 -6584 34838 -6550
rect 34872 -6584 34904 -6550
rect 34803 -6640 34904 -6584
rect 34803 -6674 34838 -6640
rect 34872 -6674 34904 -6640
rect 34803 -6730 34904 -6674
rect 33616 -6793 33717 -6764
rect 34803 -6764 34838 -6730
rect 34872 -6764 34904 -6730
rect 34803 -6793 34904 -6764
rect 33616 -6826 34904 -6793
rect 33616 -6860 33674 -6826
rect 33708 -6860 33764 -6826
rect 33798 -6860 33854 -6826
rect 33888 -6860 33944 -6826
rect 33978 -6860 34034 -6826
rect 34068 -6860 34124 -6826
rect 34158 -6860 34214 -6826
rect 34248 -6860 34304 -6826
rect 34338 -6860 34394 -6826
rect 34428 -6860 34484 -6826
rect 34518 -6860 34574 -6826
rect 34608 -6860 34664 -6826
rect 34698 -6860 34754 -6826
rect 34788 -6860 34904 -6826
rect 33616 -6894 34904 -6860
rect 34976 -5639 36264 -5606
rect 34976 -5673 35034 -5639
rect 35068 -5673 35124 -5639
rect 35158 -5673 35214 -5639
rect 35248 -5673 35304 -5639
rect 35338 -5673 35394 -5639
rect 35428 -5673 35484 -5639
rect 35518 -5673 35574 -5639
rect 35608 -5673 35664 -5639
rect 35698 -5673 35754 -5639
rect 35788 -5673 35844 -5639
rect 35878 -5673 35934 -5639
rect 35968 -5673 36024 -5639
rect 36058 -5673 36114 -5639
rect 36148 -5673 36264 -5639
rect 34976 -5707 36264 -5673
rect 34976 -5740 35077 -5707
rect 34976 -5774 35011 -5740
rect 35045 -5774 35077 -5740
rect 36163 -5740 36264 -5707
rect 34976 -5830 35077 -5774
rect 34976 -5864 35011 -5830
rect 35045 -5864 35077 -5830
rect 34976 -5920 35077 -5864
rect 34976 -5954 35011 -5920
rect 35045 -5954 35077 -5920
rect 34976 -6010 35077 -5954
rect 34976 -6044 35011 -6010
rect 35045 -6044 35077 -6010
rect 34976 -6100 35077 -6044
rect 34976 -6134 35011 -6100
rect 35045 -6134 35077 -6100
rect 34976 -6190 35077 -6134
rect 34976 -6224 35011 -6190
rect 35045 -6224 35077 -6190
rect 34976 -6280 35077 -6224
rect 34976 -6314 35011 -6280
rect 35045 -6314 35077 -6280
rect 34976 -6370 35077 -6314
rect 34976 -6404 35011 -6370
rect 35045 -6404 35077 -6370
rect 34976 -6460 35077 -6404
rect 34976 -6494 35011 -6460
rect 35045 -6494 35077 -6460
rect 34976 -6550 35077 -6494
rect 34976 -6584 35011 -6550
rect 35045 -6584 35077 -6550
rect 34976 -6640 35077 -6584
rect 34976 -6674 35011 -6640
rect 35045 -6674 35077 -6640
rect 34976 -6730 35077 -6674
rect 34976 -6764 35011 -6730
rect 35045 -6764 35077 -6730
rect 36163 -5774 36198 -5740
rect 36232 -5774 36264 -5740
rect 36163 -5830 36264 -5774
rect 36163 -5864 36198 -5830
rect 36232 -5864 36264 -5830
rect 36163 -5920 36264 -5864
rect 36163 -5954 36198 -5920
rect 36232 -5954 36264 -5920
rect 36163 -6010 36264 -5954
rect 36163 -6044 36198 -6010
rect 36232 -6044 36264 -6010
rect 36163 -6100 36264 -6044
rect 36163 -6134 36198 -6100
rect 36232 -6134 36264 -6100
rect 36163 -6190 36264 -6134
rect 36163 -6224 36198 -6190
rect 36232 -6224 36264 -6190
rect 36163 -6280 36264 -6224
rect 36163 -6314 36198 -6280
rect 36232 -6314 36264 -6280
rect 36163 -6370 36264 -6314
rect 36163 -6404 36198 -6370
rect 36232 -6404 36264 -6370
rect 36163 -6460 36264 -6404
rect 36163 -6494 36198 -6460
rect 36232 -6494 36264 -6460
rect 36163 -6550 36264 -6494
rect 36163 -6584 36198 -6550
rect 36232 -6584 36264 -6550
rect 36163 -6640 36264 -6584
rect 36163 -6674 36198 -6640
rect 36232 -6674 36264 -6640
rect 36163 -6730 36264 -6674
rect 34976 -6793 35077 -6764
rect 36163 -6764 36198 -6730
rect 36232 -6764 36264 -6730
rect 36163 -6793 36264 -6764
rect 34976 -6826 36264 -6793
rect 34976 -6860 35034 -6826
rect 35068 -6860 35124 -6826
rect 35158 -6860 35214 -6826
rect 35248 -6860 35304 -6826
rect 35338 -6860 35394 -6826
rect 35428 -6860 35484 -6826
rect 35518 -6860 35574 -6826
rect 35608 -6860 35664 -6826
rect 35698 -6860 35754 -6826
rect 35788 -6860 35844 -6826
rect 35878 -6860 35934 -6826
rect 35968 -6860 36024 -6826
rect 36058 -6860 36114 -6826
rect 36148 -6860 36264 -6826
rect 34976 -6894 36264 -6860
rect 36336 -5639 37624 -5606
rect 36336 -5673 36394 -5639
rect 36428 -5673 36484 -5639
rect 36518 -5673 36574 -5639
rect 36608 -5673 36664 -5639
rect 36698 -5673 36754 -5639
rect 36788 -5673 36844 -5639
rect 36878 -5673 36934 -5639
rect 36968 -5673 37024 -5639
rect 37058 -5673 37114 -5639
rect 37148 -5673 37204 -5639
rect 37238 -5673 37294 -5639
rect 37328 -5673 37384 -5639
rect 37418 -5673 37474 -5639
rect 37508 -5673 37624 -5639
rect 36336 -5707 37624 -5673
rect 36336 -5740 36437 -5707
rect 36336 -5774 36371 -5740
rect 36405 -5774 36437 -5740
rect 37523 -5740 37624 -5707
rect 36336 -5830 36437 -5774
rect 36336 -5864 36371 -5830
rect 36405 -5864 36437 -5830
rect 36336 -5920 36437 -5864
rect 36336 -5954 36371 -5920
rect 36405 -5954 36437 -5920
rect 36336 -6010 36437 -5954
rect 36336 -6044 36371 -6010
rect 36405 -6044 36437 -6010
rect 36336 -6100 36437 -6044
rect 36336 -6134 36371 -6100
rect 36405 -6134 36437 -6100
rect 36336 -6190 36437 -6134
rect 36336 -6224 36371 -6190
rect 36405 -6224 36437 -6190
rect 36336 -6280 36437 -6224
rect 36336 -6314 36371 -6280
rect 36405 -6314 36437 -6280
rect 36336 -6370 36437 -6314
rect 36336 -6404 36371 -6370
rect 36405 -6404 36437 -6370
rect 36336 -6460 36437 -6404
rect 36336 -6494 36371 -6460
rect 36405 -6494 36437 -6460
rect 36336 -6550 36437 -6494
rect 36336 -6584 36371 -6550
rect 36405 -6584 36437 -6550
rect 36336 -6640 36437 -6584
rect 36336 -6674 36371 -6640
rect 36405 -6674 36437 -6640
rect 36336 -6730 36437 -6674
rect 36336 -6764 36371 -6730
rect 36405 -6764 36437 -6730
rect 37523 -5774 37558 -5740
rect 37592 -5774 37624 -5740
rect 37523 -5830 37624 -5774
rect 37523 -5864 37558 -5830
rect 37592 -5864 37624 -5830
rect 37523 -5920 37624 -5864
rect 37523 -5954 37558 -5920
rect 37592 -5954 37624 -5920
rect 37523 -6010 37624 -5954
rect 37523 -6044 37558 -6010
rect 37592 -6044 37624 -6010
rect 37523 -6100 37624 -6044
rect 37523 -6134 37558 -6100
rect 37592 -6134 37624 -6100
rect 37523 -6190 37624 -6134
rect 37523 -6224 37558 -6190
rect 37592 -6224 37624 -6190
rect 37523 -6280 37624 -6224
rect 37523 -6314 37558 -6280
rect 37592 -6314 37624 -6280
rect 37523 -6370 37624 -6314
rect 37523 -6404 37558 -6370
rect 37592 -6404 37624 -6370
rect 37523 -6460 37624 -6404
rect 37523 -6494 37558 -6460
rect 37592 -6494 37624 -6460
rect 37523 -6550 37624 -6494
rect 37523 -6584 37558 -6550
rect 37592 -6584 37624 -6550
rect 37523 -6640 37624 -6584
rect 37523 -6674 37558 -6640
rect 37592 -6674 37624 -6640
rect 37523 -6730 37624 -6674
rect 36336 -6793 36437 -6764
rect 37523 -6764 37558 -6730
rect 37592 -6764 37624 -6730
rect 37523 -6793 37624 -6764
rect 36336 -6826 37624 -6793
rect 36336 -6860 36394 -6826
rect 36428 -6860 36484 -6826
rect 36518 -6860 36574 -6826
rect 36608 -6860 36664 -6826
rect 36698 -6860 36754 -6826
rect 36788 -6860 36844 -6826
rect 36878 -6860 36934 -6826
rect 36968 -6860 37024 -6826
rect 37058 -6860 37114 -6826
rect 37148 -6860 37204 -6826
rect 37238 -6860 37294 -6826
rect 37328 -6860 37384 -6826
rect 37418 -6860 37474 -6826
rect 37508 -6860 37624 -6826
rect 36336 -6894 37624 -6860
rect 33616 -6999 34904 -6966
rect 33616 -7033 33674 -6999
rect 33708 -7033 33764 -6999
rect 33798 -7033 33854 -6999
rect 33888 -7033 33944 -6999
rect 33978 -7033 34034 -6999
rect 34068 -7033 34124 -6999
rect 34158 -7033 34214 -6999
rect 34248 -7033 34304 -6999
rect 34338 -7033 34394 -6999
rect 34428 -7033 34484 -6999
rect 34518 -7033 34574 -6999
rect 34608 -7033 34664 -6999
rect 34698 -7033 34754 -6999
rect 34788 -7033 34904 -6999
rect 33616 -7067 34904 -7033
rect 33616 -7100 33717 -7067
rect 33616 -7134 33651 -7100
rect 33685 -7134 33717 -7100
rect 34803 -7100 34904 -7067
rect 33616 -7190 33717 -7134
rect 33616 -7224 33651 -7190
rect 33685 -7224 33717 -7190
rect 33616 -7280 33717 -7224
rect 33616 -7314 33651 -7280
rect 33685 -7314 33717 -7280
rect 33616 -7370 33717 -7314
rect 33616 -7404 33651 -7370
rect 33685 -7404 33717 -7370
rect 33616 -7460 33717 -7404
rect 33616 -7494 33651 -7460
rect 33685 -7494 33717 -7460
rect 33616 -7550 33717 -7494
rect 33616 -7584 33651 -7550
rect 33685 -7584 33717 -7550
rect 33616 -7640 33717 -7584
rect 33616 -7674 33651 -7640
rect 33685 -7674 33717 -7640
rect 33616 -7730 33717 -7674
rect 33616 -7764 33651 -7730
rect 33685 -7764 33717 -7730
rect 33616 -7820 33717 -7764
rect 33616 -7854 33651 -7820
rect 33685 -7854 33717 -7820
rect 33616 -7910 33717 -7854
rect 33616 -7944 33651 -7910
rect 33685 -7944 33717 -7910
rect 33616 -8000 33717 -7944
rect 33616 -8034 33651 -8000
rect 33685 -8034 33717 -8000
rect 33616 -8090 33717 -8034
rect 33616 -8124 33651 -8090
rect 33685 -8124 33717 -8090
rect 34803 -7134 34838 -7100
rect 34872 -7134 34904 -7100
rect 34803 -7190 34904 -7134
rect 34803 -7224 34838 -7190
rect 34872 -7224 34904 -7190
rect 34803 -7280 34904 -7224
rect 34803 -7314 34838 -7280
rect 34872 -7314 34904 -7280
rect 34803 -7370 34904 -7314
rect 34803 -7404 34838 -7370
rect 34872 -7404 34904 -7370
rect 34803 -7460 34904 -7404
rect 34803 -7494 34838 -7460
rect 34872 -7494 34904 -7460
rect 34803 -7550 34904 -7494
rect 34803 -7584 34838 -7550
rect 34872 -7584 34904 -7550
rect 34803 -7640 34904 -7584
rect 34803 -7674 34838 -7640
rect 34872 -7674 34904 -7640
rect 34803 -7730 34904 -7674
rect 34803 -7764 34838 -7730
rect 34872 -7764 34904 -7730
rect 34803 -7820 34904 -7764
rect 34803 -7854 34838 -7820
rect 34872 -7854 34904 -7820
rect 34803 -7910 34904 -7854
rect 34803 -7944 34838 -7910
rect 34872 -7944 34904 -7910
rect 34803 -8000 34904 -7944
rect 34803 -8034 34838 -8000
rect 34872 -8034 34904 -8000
rect 34803 -8090 34904 -8034
rect 33616 -8153 33717 -8124
rect 34803 -8124 34838 -8090
rect 34872 -8124 34904 -8090
rect 34803 -8153 34904 -8124
rect 33616 -8186 34904 -8153
rect 33616 -8220 33674 -8186
rect 33708 -8220 33764 -8186
rect 33798 -8220 33854 -8186
rect 33888 -8220 33944 -8186
rect 33978 -8220 34034 -8186
rect 34068 -8220 34124 -8186
rect 34158 -8220 34214 -8186
rect 34248 -8220 34304 -8186
rect 34338 -8220 34394 -8186
rect 34428 -8220 34484 -8186
rect 34518 -8220 34574 -8186
rect 34608 -8220 34664 -8186
rect 34698 -8220 34754 -8186
rect 34788 -8220 34904 -8186
rect 33616 -8254 34904 -8220
rect 34976 -6999 36264 -6966
rect 34976 -7033 35034 -6999
rect 35068 -7033 35124 -6999
rect 35158 -7033 35214 -6999
rect 35248 -7033 35304 -6999
rect 35338 -7033 35394 -6999
rect 35428 -7033 35484 -6999
rect 35518 -7033 35574 -6999
rect 35608 -7033 35664 -6999
rect 35698 -7033 35754 -6999
rect 35788 -7033 35844 -6999
rect 35878 -7033 35934 -6999
rect 35968 -7033 36024 -6999
rect 36058 -7033 36114 -6999
rect 36148 -7033 36264 -6999
rect 34976 -7067 36264 -7033
rect 34976 -7100 35077 -7067
rect 34976 -7134 35011 -7100
rect 35045 -7134 35077 -7100
rect 36163 -7100 36264 -7067
rect 34976 -7190 35077 -7134
rect 34976 -7224 35011 -7190
rect 35045 -7224 35077 -7190
rect 34976 -7280 35077 -7224
rect 34976 -7314 35011 -7280
rect 35045 -7314 35077 -7280
rect 34976 -7370 35077 -7314
rect 34976 -7404 35011 -7370
rect 35045 -7404 35077 -7370
rect 34976 -7460 35077 -7404
rect 34976 -7494 35011 -7460
rect 35045 -7494 35077 -7460
rect 34976 -7550 35077 -7494
rect 34976 -7584 35011 -7550
rect 35045 -7584 35077 -7550
rect 34976 -7640 35077 -7584
rect 34976 -7674 35011 -7640
rect 35045 -7674 35077 -7640
rect 34976 -7730 35077 -7674
rect 34976 -7764 35011 -7730
rect 35045 -7764 35077 -7730
rect 34976 -7820 35077 -7764
rect 34976 -7854 35011 -7820
rect 35045 -7854 35077 -7820
rect 34976 -7910 35077 -7854
rect 34976 -7944 35011 -7910
rect 35045 -7944 35077 -7910
rect 34976 -8000 35077 -7944
rect 34976 -8034 35011 -8000
rect 35045 -8034 35077 -8000
rect 34976 -8090 35077 -8034
rect 34976 -8124 35011 -8090
rect 35045 -8124 35077 -8090
rect 36163 -7134 36198 -7100
rect 36232 -7134 36264 -7100
rect 36163 -7190 36264 -7134
rect 36163 -7224 36198 -7190
rect 36232 -7224 36264 -7190
rect 36163 -7280 36264 -7224
rect 36163 -7314 36198 -7280
rect 36232 -7314 36264 -7280
rect 36163 -7370 36264 -7314
rect 36163 -7404 36198 -7370
rect 36232 -7404 36264 -7370
rect 36163 -7460 36264 -7404
rect 36163 -7494 36198 -7460
rect 36232 -7494 36264 -7460
rect 36163 -7550 36264 -7494
rect 36163 -7584 36198 -7550
rect 36232 -7584 36264 -7550
rect 36163 -7640 36264 -7584
rect 36163 -7674 36198 -7640
rect 36232 -7674 36264 -7640
rect 36163 -7730 36264 -7674
rect 36163 -7764 36198 -7730
rect 36232 -7764 36264 -7730
rect 36163 -7820 36264 -7764
rect 36163 -7854 36198 -7820
rect 36232 -7854 36264 -7820
rect 36163 -7910 36264 -7854
rect 36163 -7944 36198 -7910
rect 36232 -7944 36264 -7910
rect 36163 -8000 36264 -7944
rect 36163 -8034 36198 -8000
rect 36232 -8034 36264 -8000
rect 36163 -8090 36264 -8034
rect 34976 -8153 35077 -8124
rect 36163 -8124 36198 -8090
rect 36232 -8124 36264 -8090
rect 36163 -8153 36264 -8124
rect 34976 -8186 36264 -8153
rect 34976 -8220 35034 -8186
rect 35068 -8220 35124 -8186
rect 35158 -8220 35214 -8186
rect 35248 -8220 35304 -8186
rect 35338 -8220 35394 -8186
rect 35428 -8220 35484 -8186
rect 35518 -8220 35574 -8186
rect 35608 -8220 35664 -8186
rect 35698 -8220 35754 -8186
rect 35788 -8220 35844 -8186
rect 35878 -8220 35934 -8186
rect 35968 -8220 36024 -8186
rect 36058 -8220 36114 -8186
rect 36148 -8220 36264 -8186
rect 34976 -8254 36264 -8220
rect 36336 -6999 37624 -6966
rect 36336 -7033 36394 -6999
rect 36428 -7033 36484 -6999
rect 36518 -7033 36574 -6999
rect 36608 -7033 36664 -6999
rect 36698 -7033 36754 -6999
rect 36788 -7033 36844 -6999
rect 36878 -7033 36934 -6999
rect 36968 -7033 37024 -6999
rect 37058 -7033 37114 -6999
rect 37148 -7033 37204 -6999
rect 37238 -7033 37294 -6999
rect 37328 -7033 37384 -6999
rect 37418 -7033 37474 -6999
rect 37508 -7033 37624 -6999
rect 36336 -7067 37624 -7033
rect 36336 -7100 36437 -7067
rect 36336 -7134 36371 -7100
rect 36405 -7134 36437 -7100
rect 37523 -7100 37624 -7067
rect 36336 -7190 36437 -7134
rect 36336 -7224 36371 -7190
rect 36405 -7224 36437 -7190
rect 36336 -7280 36437 -7224
rect 36336 -7314 36371 -7280
rect 36405 -7314 36437 -7280
rect 36336 -7370 36437 -7314
rect 36336 -7404 36371 -7370
rect 36405 -7404 36437 -7370
rect 36336 -7460 36437 -7404
rect 36336 -7494 36371 -7460
rect 36405 -7494 36437 -7460
rect 36336 -7550 36437 -7494
rect 36336 -7584 36371 -7550
rect 36405 -7584 36437 -7550
rect 36336 -7640 36437 -7584
rect 36336 -7674 36371 -7640
rect 36405 -7674 36437 -7640
rect 36336 -7730 36437 -7674
rect 36336 -7764 36371 -7730
rect 36405 -7764 36437 -7730
rect 36336 -7820 36437 -7764
rect 36336 -7854 36371 -7820
rect 36405 -7854 36437 -7820
rect 36336 -7910 36437 -7854
rect 36336 -7944 36371 -7910
rect 36405 -7944 36437 -7910
rect 36336 -8000 36437 -7944
rect 36336 -8034 36371 -8000
rect 36405 -8034 36437 -8000
rect 36336 -8090 36437 -8034
rect 36336 -8124 36371 -8090
rect 36405 -8124 36437 -8090
rect 37523 -7134 37558 -7100
rect 37592 -7134 37624 -7100
rect 37523 -7190 37624 -7134
rect 37523 -7224 37558 -7190
rect 37592 -7224 37624 -7190
rect 37523 -7280 37624 -7224
rect 37523 -7314 37558 -7280
rect 37592 -7314 37624 -7280
rect 37523 -7370 37624 -7314
rect 37523 -7404 37558 -7370
rect 37592 -7404 37624 -7370
rect 37523 -7460 37624 -7404
rect 37523 -7494 37558 -7460
rect 37592 -7494 37624 -7460
rect 37523 -7550 37624 -7494
rect 37523 -7584 37558 -7550
rect 37592 -7584 37624 -7550
rect 37523 -7640 37624 -7584
rect 37523 -7674 37558 -7640
rect 37592 -7674 37624 -7640
rect 37523 -7730 37624 -7674
rect 37523 -7764 37558 -7730
rect 37592 -7764 37624 -7730
rect 37523 -7820 37624 -7764
rect 37523 -7854 37558 -7820
rect 37592 -7854 37624 -7820
rect 37523 -7910 37624 -7854
rect 37523 -7944 37558 -7910
rect 37592 -7944 37624 -7910
rect 37523 -8000 37624 -7944
rect 37523 -8034 37558 -8000
rect 37592 -8034 37624 -8000
rect 37523 -8090 37624 -8034
rect 36336 -8153 36437 -8124
rect 37523 -8124 37558 -8090
rect 37592 -8124 37624 -8090
rect 37523 -8153 37624 -8124
rect 36336 -8186 37624 -8153
rect 36336 -8220 36394 -8186
rect 36428 -8220 36484 -8186
rect 36518 -8220 36574 -8186
rect 36608 -8220 36664 -8186
rect 36698 -8220 36754 -8186
rect 36788 -8220 36844 -8186
rect 36878 -8220 36934 -8186
rect 36968 -8220 37024 -8186
rect 37058 -8220 37114 -8186
rect 37148 -8220 37204 -8186
rect 37238 -8220 37294 -8186
rect 37328 -8220 37384 -8186
rect 37418 -8220 37474 -8186
rect 37508 -8220 37624 -8186
rect 36336 -8254 37624 -8220
rect 35550 -8340 35650 -8310
rect 35550 -8380 35580 -8340
rect 35620 -8380 35650 -8340
rect 35550 -8440 35650 -8380
rect 35550 -8480 35580 -8440
rect 35620 -8480 35650 -8440
rect 35550 -8540 35650 -8480
rect 35550 -8580 35580 -8540
rect 35620 -8580 35650 -8540
rect 35550 -8610 35650 -8580
<< nsubdiff >>
rect 5970 7110 6360 7150
rect 6520 7110 6910 7150
rect 5970 6940 6010 7110
rect 5970 6610 6010 6780
rect 6870 6940 6910 7110
rect 6870 6610 6910 6780
rect 5970 6570 6360 6610
rect 6520 6570 6910 6610
rect 7250 7110 8080 7150
rect 8240 7110 9070 7150
rect 7250 6940 7290 7110
rect 7250 6610 7290 6780
rect 9030 6940 9070 7110
rect 9030 6610 9070 6780
rect 7250 6570 8080 6610
rect 8240 6570 9070 6610
rect 9410 7110 9800 7150
rect 9960 7110 10350 7150
rect 9410 6940 9450 7110
rect 9410 6610 9450 6780
rect 10310 6940 10350 7110
rect 10310 6610 10350 6780
rect 9410 6570 9800 6610
rect 9930 6570 10350 6610
rect 6400 6180 8080 6220
rect 8240 6180 9920 6220
rect 5330 5980 5610 6020
rect 5770 5980 6050 6020
rect 5330 5810 5370 5980
rect 5330 5480 5370 5650
rect 6010 5810 6050 5980
rect 6010 5480 6050 5650
rect 5330 5440 5610 5480
rect 5770 5440 6050 5480
rect 6400 5810 6440 6180
rect 6400 5270 6440 5650
rect 9880 5810 9920 6180
rect 9880 5270 9920 5650
rect 10260 5980 10540 6020
rect 10700 5980 10980 6020
rect 10260 5810 10300 5980
rect 10260 5480 10300 5650
rect 10940 5810 10980 5980
rect 10940 5480 10980 5650
rect 10260 5440 10540 5480
rect 10700 5440 10980 5480
rect 6400 5230 8080 5270
rect 8240 5230 9920 5270
rect 5300 4800 6560 4840
rect 6720 4800 7980 4840
rect 5300 4630 5340 4800
rect 5300 4300 5340 4470
rect 7940 4630 7980 4800
rect 7940 4300 7980 4470
rect 5300 4260 6560 4300
rect 6720 4260 7980 4300
rect 8340 4800 9600 4840
rect 9760 4800 11020 4840
rect 8340 4630 8380 4800
rect 8340 4300 8380 4470
rect 10980 4630 11020 4800
rect 10980 4300 11020 4470
rect 8340 4260 9600 4300
rect 9760 4260 11020 4300
rect 35970 4110 36360 4150
rect 36520 4110 36910 4150
rect 35970 3940 36010 4110
rect 35970 3610 36010 3780
rect 36870 3940 36910 4110
rect 36870 3610 36910 3780
rect 35970 3570 36360 3610
rect 36520 3570 36910 3610
rect 37250 4110 38080 4150
rect 38240 4110 39070 4150
rect 37250 3940 37290 4110
rect 37250 3610 37290 3780
rect 39030 3940 39070 4110
rect 39030 3610 39070 3780
rect 37250 3570 38080 3610
rect 38240 3570 39070 3610
rect 39410 4110 39800 4150
rect 39960 4110 40350 4150
rect 39410 3940 39450 4110
rect 39410 3610 39450 3780
rect 40310 3940 40350 4110
rect 40310 3610 40350 3780
rect 39410 3570 39800 3610
rect 39930 3570 40350 3610
rect 36400 3180 38080 3220
rect 38240 3180 39920 3220
rect 35330 2980 35610 3020
rect 35770 2980 36050 3020
rect 35330 2810 35370 2980
rect 35330 2480 35370 2650
rect 36010 2810 36050 2980
rect 36010 2480 36050 2650
rect 35330 2440 35610 2480
rect 35770 2440 36050 2480
rect 36400 2810 36440 3180
rect 36400 2270 36440 2650
rect 39880 2810 39920 3180
rect 39880 2270 39920 2650
rect 40260 2980 40540 3020
rect 40700 2980 40980 3020
rect 40260 2810 40300 2980
rect 40260 2480 40300 2650
rect 40940 2810 40980 2980
rect 40940 2480 40980 2650
rect 40260 2440 40540 2480
rect 40700 2440 40980 2480
rect 36400 2230 38080 2270
rect 38240 2230 39920 2270
rect 35300 1800 36560 1840
rect 36720 1800 37980 1840
rect 35300 1630 35340 1800
rect 35300 1300 35340 1470
rect 37940 1630 37980 1800
rect 37940 1300 37980 1470
rect 35300 1260 36560 1300
rect 36720 1260 37980 1300
rect 38340 1800 39600 1840
rect 39760 1800 41020 1840
rect 38340 1630 38380 1800
rect 38340 1300 38380 1470
rect 40980 1630 41020 1800
rect 40980 1300 41020 1470
rect 38340 1260 39600 1300
rect 39760 1260 41020 1300
rect 33779 -4428 34741 -4409
rect 33779 -4462 33874 -4428
rect 33908 -4462 33964 -4428
rect 33998 -4462 34054 -4428
rect 34088 -4462 34144 -4428
rect 34178 -4462 34234 -4428
rect 34268 -4462 34324 -4428
rect 34358 -4462 34414 -4428
rect 34448 -4462 34504 -4428
rect 34538 -4462 34594 -4428
rect 34628 -4462 34741 -4428
rect 33779 -4481 34741 -4462
rect 33779 -4486 33851 -4481
rect 33779 -4520 33798 -4486
rect 33832 -4520 33851 -4486
rect 33779 -4576 33851 -4520
rect 34669 -4520 34741 -4481
rect 33779 -4610 33798 -4576
rect 33832 -4610 33851 -4576
rect 33779 -4666 33851 -4610
rect 33779 -4700 33798 -4666
rect 33832 -4700 33851 -4666
rect 33779 -4756 33851 -4700
rect 33779 -4790 33798 -4756
rect 33832 -4790 33851 -4756
rect 33779 -4846 33851 -4790
rect 33779 -4880 33798 -4846
rect 33832 -4880 33851 -4846
rect 33779 -4936 33851 -4880
rect 33779 -4970 33798 -4936
rect 33832 -4970 33851 -4936
rect 33779 -5026 33851 -4970
rect 33779 -5060 33798 -5026
rect 33832 -5060 33851 -5026
rect 33779 -5116 33851 -5060
rect 33779 -5150 33798 -5116
rect 33832 -5150 33851 -5116
rect 33779 -5206 33851 -5150
rect 33779 -5240 33798 -5206
rect 33832 -5240 33851 -5206
rect 34669 -4554 34688 -4520
rect 34722 -4554 34741 -4520
rect 34669 -4610 34741 -4554
rect 34669 -4644 34688 -4610
rect 34722 -4644 34741 -4610
rect 34669 -4700 34741 -4644
rect 34669 -4734 34688 -4700
rect 34722 -4734 34741 -4700
rect 34669 -4790 34741 -4734
rect 34669 -4824 34688 -4790
rect 34722 -4824 34741 -4790
rect 34669 -4880 34741 -4824
rect 34669 -4914 34688 -4880
rect 34722 -4914 34741 -4880
rect 34669 -4970 34741 -4914
rect 34669 -5004 34688 -4970
rect 34722 -5004 34741 -4970
rect 34669 -5060 34741 -5004
rect 34669 -5094 34688 -5060
rect 34722 -5094 34741 -5060
rect 34669 -5150 34741 -5094
rect 34669 -5184 34688 -5150
rect 34722 -5184 34741 -5150
rect 33779 -5299 33851 -5240
rect 34669 -5240 34741 -5184
rect 34669 -5274 34688 -5240
rect 34722 -5274 34741 -5240
rect 34669 -5299 34741 -5274
rect 33779 -5318 34741 -5299
rect 33779 -5352 33855 -5318
rect 33889 -5352 33945 -5318
rect 33979 -5352 34035 -5318
rect 34069 -5352 34125 -5318
rect 34159 -5352 34215 -5318
rect 34249 -5352 34305 -5318
rect 34339 -5352 34395 -5318
rect 34429 -5352 34485 -5318
rect 34519 -5352 34575 -5318
rect 34609 -5352 34741 -5318
rect 33779 -5371 34741 -5352
rect 35139 -4428 36101 -4409
rect 35139 -4462 35234 -4428
rect 35268 -4462 35324 -4428
rect 35358 -4462 35414 -4428
rect 35448 -4462 35504 -4428
rect 35538 -4462 35594 -4428
rect 35628 -4462 35684 -4428
rect 35718 -4462 35774 -4428
rect 35808 -4462 35864 -4428
rect 35898 -4462 35954 -4428
rect 35988 -4462 36101 -4428
rect 35139 -4481 36101 -4462
rect 35139 -4486 35211 -4481
rect 35139 -4520 35158 -4486
rect 35192 -4520 35211 -4486
rect 35139 -4576 35211 -4520
rect 36029 -4520 36101 -4481
rect 35139 -4610 35158 -4576
rect 35192 -4610 35211 -4576
rect 35139 -4666 35211 -4610
rect 35139 -4700 35158 -4666
rect 35192 -4700 35211 -4666
rect 35139 -4756 35211 -4700
rect 35139 -4790 35158 -4756
rect 35192 -4790 35211 -4756
rect 35139 -4846 35211 -4790
rect 35139 -4880 35158 -4846
rect 35192 -4880 35211 -4846
rect 35139 -4936 35211 -4880
rect 35139 -4970 35158 -4936
rect 35192 -4970 35211 -4936
rect 35139 -5026 35211 -4970
rect 35139 -5060 35158 -5026
rect 35192 -5060 35211 -5026
rect 35139 -5116 35211 -5060
rect 35139 -5150 35158 -5116
rect 35192 -5150 35211 -5116
rect 35139 -5206 35211 -5150
rect 35139 -5240 35158 -5206
rect 35192 -5240 35211 -5206
rect 36029 -4554 36048 -4520
rect 36082 -4554 36101 -4520
rect 36029 -4610 36101 -4554
rect 36029 -4644 36048 -4610
rect 36082 -4644 36101 -4610
rect 36029 -4700 36101 -4644
rect 36029 -4734 36048 -4700
rect 36082 -4734 36101 -4700
rect 36029 -4790 36101 -4734
rect 36029 -4824 36048 -4790
rect 36082 -4824 36101 -4790
rect 36029 -4880 36101 -4824
rect 36029 -4914 36048 -4880
rect 36082 -4914 36101 -4880
rect 36029 -4970 36101 -4914
rect 36029 -5004 36048 -4970
rect 36082 -5004 36101 -4970
rect 36029 -5060 36101 -5004
rect 36029 -5094 36048 -5060
rect 36082 -5094 36101 -5060
rect 36029 -5150 36101 -5094
rect 36029 -5184 36048 -5150
rect 36082 -5184 36101 -5150
rect 35139 -5299 35211 -5240
rect 36029 -5240 36101 -5184
rect 36029 -5274 36048 -5240
rect 36082 -5274 36101 -5240
rect 36029 -5299 36101 -5274
rect 35139 -5318 36101 -5299
rect 35139 -5352 35215 -5318
rect 35249 -5352 35305 -5318
rect 35339 -5352 35395 -5318
rect 35429 -5352 35485 -5318
rect 35519 -5352 35575 -5318
rect 35609 -5352 35665 -5318
rect 35699 -5352 35755 -5318
rect 35789 -5352 35845 -5318
rect 35879 -5352 35935 -5318
rect 35969 -5352 36101 -5318
rect 35139 -5371 36101 -5352
rect 36499 -4428 37461 -4409
rect 36499 -4462 36594 -4428
rect 36628 -4462 36684 -4428
rect 36718 -4462 36774 -4428
rect 36808 -4462 36864 -4428
rect 36898 -4462 36954 -4428
rect 36988 -4462 37044 -4428
rect 37078 -4462 37134 -4428
rect 37168 -4462 37224 -4428
rect 37258 -4462 37314 -4428
rect 37348 -4462 37461 -4428
rect 36499 -4481 37461 -4462
rect 36499 -4486 36571 -4481
rect 36499 -4520 36518 -4486
rect 36552 -4520 36571 -4486
rect 36499 -4576 36571 -4520
rect 37389 -4520 37461 -4481
rect 36499 -4610 36518 -4576
rect 36552 -4610 36571 -4576
rect 36499 -4666 36571 -4610
rect 36499 -4700 36518 -4666
rect 36552 -4700 36571 -4666
rect 36499 -4756 36571 -4700
rect 36499 -4790 36518 -4756
rect 36552 -4790 36571 -4756
rect 36499 -4846 36571 -4790
rect 36499 -4880 36518 -4846
rect 36552 -4880 36571 -4846
rect 36499 -4936 36571 -4880
rect 36499 -4970 36518 -4936
rect 36552 -4970 36571 -4936
rect 36499 -5026 36571 -4970
rect 36499 -5060 36518 -5026
rect 36552 -5060 36571 -5026
rect 36499 -5116 36571 -5060
rect 36499 -5150 36518 -5116
rect 36552 -5150 36571 -5116
rect 36499 -5206 36571 -5150
rect 36499 -5240 36518 -5206
rect 36552 -5240 36571 -5206
rect 37389 -4554 37408 -4520
rect 37442 -4554 37461 -4520
rect 37389 -4610 37461 -4554
rect 37389 -4644 37408 -4610
rect 37442 -4644 37461 -4610
rect 37389 -4700 37461 -4644
rect 37389 -4734 37408 -4700
rect 37442 -4734 37461 -4700
rect 37389 -4790 37461 -4734
rect 37389 -4824 37408 -4790
rect 37442 -4824 37461 -4790
rect 37389 -4880 37461 -4824
rect 37389 -4914 37408 -4880
rect 37442 -4914 37461 -4880
rect 37389 -4970 37461 -4914
rect 37389 -5004 37408 -4970
rect 37442 -5004 37461 -4970
rect 37389 -5060 37461 -5004
rect 37389 -5094 37408 -5060
rect 37442 -5094 37461 -5060
rect 37389 -5150 37461 -5094
rect 37389 -5184 37408 -5150
rect 37442 -5184 37461 -5150
rect 36499 -5299 36571 -5240
rect 37389 -5240 37461 -5184
rect 37389 -5274 37408 -5240
rect 37442 -5274 37461 -5240
rect 37389 -5299 37461 -5274
rect 36499 -5318 37461 -5299
rect 36499 -5352 36575 -5318
rect 36609 -5352 36665 -5318
rect 36699 -5352 36755 -5318
rect 36789 -5352 36845 -5318
rect 36879 -5352 36935 -5318
rect 36969 -5352 37025 -5318
rect 37059 -5352 37115 -5318
rect 37149 -5352 37205 -5318
rect 37239 -5352 37295 -5318
rect 37329 -5352 37461 -5318
rect 36499 -5371 37461 -5352
rect 33779 -5788 34741 -5769
rect 33779 -5822 33874 -5788
rect 33908 -5822 33964 -5788
rect 33998 -5822 34054 -5788
rect 34088 -5822 34144 -5788
rect 34178 -5822 34234 -5788
rect 34268 -5822 34324 -5788
rect 34358 -5822 34414 -5788
rect 34448 -5822 34504 -5788
rect 34538 -5822 34594 -5788
rect 34628 -5822 34741 -5788
rect 33779 -5841 34741 -5822
rect 33779 -5846 33851 -5841
rect 33779 -5880 33798 -5846
rect 33832 -5880 33851 -5846
rect 33779 -5936 33851 -5880
rect 34669 -5880 34741 -5841
rect 33779 -5970 33798 -5936
rect 33832 -5970 33851 -5936
rect 33779 -6026 33851 -5970
rect 33779 -6060 33798 -6026
rect 33832 -6060 33851 -6026
rect 33779 -6116 33851 -6060
rect 33779 -6150 33798 -6116
rect 33832 -6150 33851 -6116
rect 33779 -6206 33851 -6150
rect 33779 -6240 33798 -6206
rect 33832 -6240 33851 -6206
rect 33779 -6296 33851 -6240
rect 33779 -6330 33798 -6296
rect 33832 -6330 33851 -6296
rect 33779 -6386 33851 -6330
rect 33779 -6420 33798 -6386
rect 33832 -6420 33851 -6386
rect 33779 -6476 33851 -6420
rect 33779 -6510 33798 -6476
rect 33832 -6510 33851 -6476
rect 33779 -6566 33851 -6510
rect 33779 -6600 33798 -6566
rect 33832 -6600 33851 -6566
rect 34669 -5914 34688 -5880
rect 34722 -5914 34741 -5880
rect 34669 -5970 34741 -5914
rect 34669 -6004 34688 -5970
rect 34722 -6004 34741 -5970
rect 34669 -6060 34741 -6004
rect 34669 -6094 34688 -6060
rect 34722 -6094 34741 -6060
rect 34669 -6150 34741 -6094
rect 34669 -6184 34688 -6150
rect 34722 -6184 34741 -6150
rect 34669 -6240 34741 -6184
rect 34669 -6274 34688 -6240
rect 34722 -6274 34741 -6240
rect 34669 -6330 34741 -6274
rect 34669 -6364 34688 -6330
rect 34722 -6364 34741 -6330
rect 34669 -6420 34741 -6364
rect 34669 -6454 34688 -6420
rect 34722 -6454 34741 -6420
rect 34669 -6510 34741 -6454
rect 34669 -6544 34688 -6510
rect 34722 -6544 34741 -6510
rect 33779 -6659 33851 -6600
rect 34669 -6600 34741 -6544
rect 34669 -6634 34688 -6600
rect 34722 -6634 34741 -6600
rect 34669 -6659 34741 -6634
rect 33779 -6678 34741 -6659
rect 33779 -6712 33855 -6678
rect 33889 -6712 33945 -6678
rect 33979 -6712 34035 -6678
rect 34069 -6712 34125 -6678
rect 34159 -6712 34215 -6678
rect 34249 -6712 34305 -6678
rect 34339 -6712 34395 -6678
rect 34429 -6712 34485 -6678
rect 34519 -6712 34575 -6678
rect 34609 -6712 34741 -6678
rect 33779 -6731 34741 -6712
rect 35139 -5788 36101 -5769
rect 35139 -5822 35234 -5788
rect 35268 -5822 35324 -5788
rect 35358 -5822 35414 -5788
rect 35448 -5822 35504 -5788
rect 35538 -5822 35594 -5788
rect 35628 -5822 35684 -5788
rect 35718 -5822 35774 -5788
rect 35808 -5822 35864 -5788
rect 35898 -5822 35954 -5788
rect 35988 -5822 36101 -5788
rect 35139 -5841 36101 -5822
rect 35139 -5846 35211 -5841
rect 35139 -5880 35158 -5846
rect 35192 -5880 35211 -5846
rect 35139 -5936 35211 -5880
rect 36029 -5880 36101 -5841
rect 35139 -5970 35158 -5936
rect 35192 -5970 35211 -5936
rect 35139 -6026 35211 -5970
rect 35139 -6060 35158 -6026
rect 35192 -6060 35211 -6026
rect 35139 -6116 35211 -6060
rect 35139 -6150 35158 -6116
rect 35192 -6150 35211 -6116
rect 35139 -6206 35211 -6150
rect 35139 -6240 35158 -6206
rect 35192 -6240 35211 -6206
rect 35139 -6296 35211 -6240
rect 35139 -6330 35158 -6296
rect 35192 -6330 35211 -6296
rect 35139 -6386 35211 -6330
rect 35139 -6420 35158 -6386
rect 35192 -6420 35211 -6386
rect 35139 -6476 35211 -6420
rect 35139 -6510 35158 -6476
rect 35192 -6510 35211 -6476
rect 35139 -6566 35211 -6510
rect 35139 -6600 35158 -6566
rect 35192 -6600 35211 -6566
rect 36029 -5914 36048 -5880
rect 36082 -5914 36101 -5880
rect 36029 -5970 36101 -5914
rect 36029 -6004 36048 -5970
rect 36082 -6004 36101 -5970
rect 36029 -6060 36101 -6004
rect 36029 -6094 36048 -6060
rect 36082 -6094 36101 -6060
rect 36029 -6150 36101 -6094
rect 36029 -6184 36048 -6150
rect 36082 -6184 36101 -6150
rect 36029 -6240 36101 -6184
rect 36029 -6274 36048 -6240
rect 36082 -6274 36101 -6240
rect 36029 -6330 36101 -6274
rect 36029 -6364 36048 -6330
rect 36082 -6364 36101 -6330
rect 36029 -6420 36101 -6364
rect 36029 -6454 36048 -6420
rect 36082 -6454 36101 -6420
rect 36029 -6510 36101 -6454
rect 36029 -6544 36048 -6510
rect 36082 -6544 36101 -6510
rect 35139 -6659 35211 -6600
rect 36029 -6600 36101 -6544
rect 36029 -6634 36048 -6600
rect 36082 -6634 36101 -6600
rect 36029 -6659 36101 -6634
rect 35139 -6678 36101 -6659
rect 35139 -6712 35215 -6678
rect 35249 -6712 35305 -6678
rect 35339 -6712 35395 -6678
rect 35429 -6712 35485 -6678
rect 35519 -6712 35575 -6678
rect 35609 -6712 35665 -6678
rect 35699 -6712 35755 -6678
rect 35789 -6712 35845 -6678
rect 35879 -6712 35935 -6678
rect 35969 -6712 36101 -6678
rect 35139 -6731 36101 -6712
rect 36499 -5788 37461 -5769
rect 36499 -5822 36594 -5788
rect 36628 -5822 36684 -5788
rect 36718 -5822 36774 -5788
rect 36808 -5822 36864 -5788
rect 36898 -5822 36954 -5788
rect 36988 -5822 37044 -5788
rect 37078 -5822 37134 -5788
rect 37168 -5822 37224 -5788
rect 37258 -5822 37314 -5788
rect 37348 -5822 37461 -5788
rect 36499 -5841 37461 -5822
rect 36499 -5846 36571 -5841
rect 36499 -5880 36518 -5846
rect 36552 -5880 36571 -5846
rect 36499 -5936 36571 -5880
rect 37389 -5880 37461 -5841
rect 36499 -5970 36518 -5936
rect 36552 -5970 36571 -5936
rect 36499 -6026 36571 -5970
rect 36499 -6060 36518 -6026
rect 36552 -6060 36571 -6026
rect 36499 -6116 36571 -6060
rect 36499 -6150 36518 -6116
rect 36552 -6150 36571 -6116
rect 36499 -6206 36571 -6150
rect 36499 -6240 36518 -6206
rect 36552 -6240 36571 -6206
rect 36499 -6296 36571 -6240
rect 36499 -6330 36518 -6296
rect 36552 -6330 36571 -6296
rect 36499 -6386 36571 -6330
rect 36499 -6420 36518 -6386
rect 36552 -6420 36571 -6386
rect 36499 -6476 36571 -6420
rect 36499 -6510 36518 -6476
rect 36552 -6510 36571 -6476
rect 36499 -6566 36571 -6510
rect 36499 -6600 36518 -6566
rect 36552 -6600 36571 -6566
rect 37389 -5914 37408 -5880
rect 37442 -5914 37461 -5880
rect 37389 -5970 37461 -5914
rect 37389 -6004 37408 -5970
rect 37442 -6004 37461 -5970
rect 37389 -6060 37461 -6004
rect 37389 -6094 37408 -6060
rect 37442 -6094 37461 -6060
rect 37389 -6150 37461 -6094
rect 37389 -6184 37408 -6150
rect 37442 -6184 37461 -6150
rect 37389 -6240 37461 -6184
rect 37389 -6274 37408 -6240
rect 37442 -6274 37461 -6240
rect 37389 -6330 37461 -6274
rect 37389 -6364 37408 -6330
rect 37442 -6364 37461 -6330
rect 37389 -6420 37461 -6364
rect 37389 -6454 37408 -6420
rect 37442 -6454 37461 -6420
rect 37389 -6510 37461 -6454
rect 37389 -6544 37408 -6510
rect 37442 -6544 37461 -6510
rect 36499 -6659 36571 -6600
rect 37389 -6600 37461 -6544
rect 37389 -6634 37408 -6600
rect 37442 -6634 37461 -6600
rect 37389 -6659 37461 -6634
rect 36499 -6678 37461 -6659
rect 36499 -6712 36575 -6678
rect 36609 -6712 36665 -6678
rect 36699 -6712 36755 -6678
rect 36789 -6712 36845 -6678
rect 36879 -6712 36935 -6678
rect 36969 -6712 37025 -6678
rect 37059 -6712 37115 -6678
rect 37149 -6712 37205 -6678
rect 37239 -6712 37295 -6678
rect 37329 -6712 37461 -6678
rect 36499 -6731 37461 -6712
rect 33779 -7148 34741 -7129
rect 33779 -7182 33874 -7148
rect 33908 -7182 33964 -7148
rect 33998 -7182 34054 -7148
rect 34088 -7182 34144 -7148
rect 34178 -7182 34234 -7148
rect 34268 -7182 34324 -7148
rect 34358 -7182 34414 -7148
rect 34448 -7182 34504 -7148
rect 34538 -7182 34594 -7148
rect 34628 -7182 34741 -7148
rect 33779 -7201 34741 -7182
rect 33779 -7206 33851 -7201
rect 33779 -7240 33798 -7206
rect 33832 -7240 33851 -7206
rect 33779 -7296 33851 -7240
rect 34669 -7240 34741 -7201
rect 33779 -7330 33798 -7296
rect 33832 -7330 33851 -7296
rect 33779 -7386 33851 -7330
rect 33779 -7420 33798 -7386
rect 33832 -7420 33851 -7386
rect 33779 -7476 33851 -7420
rect 33779 -7510 33798 -7476
rect 33832 -7510 33851 -7476
rect 33779 -7566 33851 -7510
rect 33779 -7600 33798 -7566
rect 33832 -7600 33851 -7566
rect 33779 -7656 33851 -7600
rect 33779 -7690 33798 -7656
rect 33832 -7690 33851 -7656
rect 33779 -7746 33851 -7690
rect 33779 -7780 33798 -7746
rect 33832 -7780 33851 -7746
rect 33779 -7836 33851 -7780
rect 33779 -7870 33798 -7836
rect 33832 -7870 33851 -7836
rect 33779 -7926 33851 -7870
rect 33779 -7960 33798 -7926
rect 33832 -7960 33851 -7926
rect 34669 -7274 34688 -7240
rect 34722 -7274 34741 -7240
rect 34669 -7330 34741 -7274
rect 34669 -7364 34688 -7330
rect 34722 -7364 34741 -7330
rect 34669 -7420 34741 -7364
rect 34669 -7454 34688 -7420
rect 34722 -7454 34741 -7420
rect 34669 -7510 34741 -7454
rect 34669 -7544 34688 -7510
rect 34722 -7544 34741 -7510
rect 34669 -7600 34741 -7544
rect 34669 -7634 34688 -7600
rect 34722 -7634 34741 -7600
rect 34669 -7690 34741 -7634
rect 34669 -7724 34688 -7690
rect 34722 -7724 34741 -7690
rect 34669 -7780 34741 -7724
rect 34669 -7814 34688 -7780
rect 34722 -7814 34741 -7780
rect 34669 -7870 34741 -7814
rect 34669 -7904 34688 -7870
rect 34722 -7904 34741 -7870
rect 33779 -8019 33851 -7960
rect 34669 -7960 34741 -7904
rect 34669 -7994 34688 -7960
rect 34722 -7994 34741 -7960
rect 34669 -8019 34741 -7994
rect 33779 -8038 34741 -8019
rect 33779 -8072 33855 -8038
rect 33889 -8072 33945 -8038
rect 33979 -8072 34035 -8038
rect 34069 -8072 34125 -8038
rect 34159 -8072 34215 -8038
rect 34249 -8072 34305 -8038
rect 34339 -8072 34395 -8038
rect 34429 -8072 34485 -8038
rect 34519 -8072 34575 -8038
rect 34609 -8072 34741 -8038
rect 33779 -8091 34741 -8072
rect 35139 -7148 36101 -7129
rect 35139 -7182 35234 -7148
rect 35268 -7182 35324 -7148
rect 35358 -7182 35414 -7148
rect 35448 -7182 35504 -7148
rect 35538 -7182 35594 -7148
rect 35628 -7182 35684 -7148
rect 35718 -7182 35774 -7148
rect 35808 -7182 35864 -7148
rect 35898 -7182 35954 -7148
rect 35988 -7182 36101 -7148
rect 35139 -7201 36101 -7182
rect 35139 -7206 35211 -7201
rect 35139 -7240 35158 -7206
rect 35192 -7240 35211 -7206
rect 35139 -7296 35211 -7240
rect 36029 -7240 36101 -7201
rect 35139 -7330 35158 -7296
rect 35192 -7330 35211 -7296
rect 35139 -7386 35211 -7330
rect 35139 -7420 35158 -7386
rect 35192 -7420 35211 -7386
rect 35139 -7476 35211 -7420
rect 35139 -7510 35158 -7476
rect 35192 -7510 35211 -7476
rect 35139 -7566 35211 -7510
rect 35139 -7600 35158 -7566
rect 35192 -7600 35211 -7566
rect 35139 -7656 35211 -7600
rect 35139 -7690 35158 -7656
rect 35192 -7690 35211 -7656
rect 35139 -7746 35211 -7690
rect 35139 -7780 35158 -7746
rect 35192 -7780 35211 -7746
rect 35139 -7836 35211 -7780
rect 35139 -7870 35158 -7836
rect 35192 -7870 35211 -7836
rect 35139 -7926 35211 -7870
rect 35139 -7960 35158 -7926
rect 35192 -7960 35211 -7926
rect 36029 -7274 36048 -7240
rect 36082 -7274 36101 -7240
rect 36029 -7330 36101 -7274
rect 36029 -7364 36048 -7330
rect 36082 -7364 36101 -7330
rect 36029 -7420 36101 -7364
rect 36029 -7454 36048 -7420
rect 36082 -7454 36101 -7420
rect 36029 -7510 36101 -7454
rect 36029 -7544 36048 -7510
rect 36082 -7544 36101 -7510
rect 36029 -7600 36101 -7544
rect 36029 -7634 36048 -7600
rect 36082 -7634 36101 -7600
rect 36029 -7690 36101 -7634
rect 36029 -7724 36048 -7690
rect 36082 -7724 36101 -7690
rect 36029 -7780 36101 -7724
rect 36029 -7814 36048 -7780
rect 36082 -7814 36101 -7780
rect 36029 -7870 36101 -7814
rect 36029 -7904 36048 -7870
rect 36082 -7904 36101 -7870
rect 35139 -8019 35211 -7960
rect 36029 -7960 36101 -7904
rect 36029 -7994 36048 -7960
rect 36082 -7994 36101 -7960
rect 36029 -8019 36101 -7994
rect 35139 -8038 36101 -8019
rect 35139 -8072 35215 -8038
rect 35249 -8072 35305 -8038
rect 35339 -8072 35395 -8038
rect 35429 -8072 35485 -8038
rect 35519 -8072 35575 -8038
rect 35609 -8072 35665 -8038
rect 35699 -8072 35755 -8038
rect 35789 -8072 35845 -8038
rect 35879 -8072 35935 -8038
rect 35969 -8072 36101 -8038
rect 35139 -8091 36101 -8072
rect 36499 -7148 37461 -7129
rect 36499 -7182 36594 -7148
rect 36628 -7182 36684 -7148
rect 36718 -7182 36774 -7148
rect 36808 -7182 36864 -7148
rect 36898 -7182 36954 -7148
rect 36988 -7182 37044 -7148
rect 37078 -7182 37134 -7148
rect 37168 -7182 37224 -7148
rect 37258 -7182 37314 -7148
rect 37348 -7182 37461 -7148
rect 36499 -7201 37461 -7182
rect 36499 -7206 36571 -7201
rect 36499 -7240 36518 -7206
rect 36552 -7240 36571 -7206
rect 36499 -7296 36571 -7240
rect 37389 -7240 37461 -7201
rect 36499 -7330 36518 -7296
rect 36552 -7330 36571 -7296
rect 36499 -7386 36571 -7330
rect 36499 -7420 36518 -7386
rect 36552 -7420 36571 -7386
rect 36499 -7476 36571 -7420
rect 36499 -7510 36518 -7476
rect 36552 -7510 36571 -7476
rect 36499 -7566 36571 -7510
rect 36499 -7600 36518 -7566
rect 36552 -7600 36571 -7566
rect 36499 -7656 36571 -7600
rect 36499 -7690 36518 -7656
rect 36552 -7690 36571 -7656
rect 36499 -7746 36571 -7690
rect 36499 -7780 36518 -7746
rect 36552 -7780 36571 -7746
rect 36499 -7836 36571 -7780
rect 36499 -7870 36518 -7836
rect 36552 -7870 36571 -7836
rect 36499 -7926 36571 -7870
rect 36499 -7960 36518 -7926
rect 36552 -7960 36571 -7926
rect 37389 -7274 37408 -7240
rect 37442 -7274 37461 -7240
rect 37389 -7330 37461 -7274
rect 37389 -7364 37408 -7330
rect 37442 -7364 37461 -7330
rect 37389 -7420 37461 -7364
rect 37389 -7454 37408 -7420
rect 37442 -7454 37461 -7420
rect 37389 -7510 37461 -7454
rect 37389 -7544 37408 -7510
rect 37442 -7544 37461 -7510
rect 37389 -7600 37461 -7544
rect 37389 -7634 37408 -7600
rect 37442 -7634 37461 -7600
rect 37389 -7690 37461 -7634
rect 37389 -7724 37408 -7690
rect 37442 -7724 37461 -7690
rect 37389 -7780 37461 -7724
rect 37389 -7814 37408 -7780
rect 37442 -7814 37461 -7780
rect 37389 -7870 37461 -7814
rect 37389 -7904 37408 -7870
rect 37442 -7904 37461 -7870
rect 36499 -8019 36571 -7960
rect 37389 -7960 37461 -7904
rect 37389 -7994 37408 -7960
rect 37442 -7994 37461 -7960
rect 37389 -8019 37461 -7994
rect 36499 -8038 37461 -8019
rect 36499 -8072 36575 -8038
rect 36609 -8072 36665 -8038
rect 36699 -8072 36755 -8038
rect 36789 -8072 36845 -8038
rect 36879 -8072 36935 -8038
rect 36969 -8072 37025 -8038
rect 37059 -8072 37115 -8038
rect 37149 -8072 37205 -8038
rect 37239 -8072 37295 -8038
rect 37329 -8072 37461 -8038
rect 36499 -8091 37461 -8072
<< psubdiffcont >>
rect 1180 7280 1340 7320
rect 50 7000 90 7160
rect 2430 7000 2470 7160
rect 1180 6850 1340 6890
rect 3690 7010 3850 7050
rect 1150 6750 1310 6790
rect 50 6470 90 6630
rect 2370 6470 2410 6630
rect 1150 6320 1310 6360
rect 2620 6490 2660 6650
rect 1150 6220 1310 6260
rect 440 6000 480 6160
rect 2000 6000 2040 6160
rect 4970 6490 5010 6650
rect 3690 6100 3850 6140
rect 1150 5900 1310 5940
rect 3690 6000 3850 6040
rect 1150 5800 1310 5840
rect 440 5580 480 5740
rect 2000 5580 2040 5740
rect 2950 5780 2990 5940
rect 4560 5780 4600 5940
rect 3690 5690 3850 5730
rect 1150 5480 1310 5520
rect 6820 4140 6980 4180
rect 6160 3770 6200 3930
rect 7600 3770 7640 3930
rect 6820 3610 6980 3650
rect 9340 4140 9500 4180
rect 8680 3770 8720 3930
rect 10120 3770 10160 3930
rect 6820 3490 6980 3530
rect -70 3390 -30 3430
rect 30 3390 70 3430
rect 130 3390 170 3430
rect 5680 3020 5720 3180
rect 8080 3020 8120 3180
rect 6820 2660 6980 2700
rect 9340 3490 9500 3530
rect 8200 3020 8240 3180
rect 10600 3020 10640 3180
rect 9340 2660 9500 2700
rect 8080 2560 8240 2600
rect 5880 2230 5920 2390
rect 10390 2230 10430 2390
rect 8080 2110 8240 2150
rect 6800 2010 6960 2050
rect 6240 1680 6280 1840
rect 7360 1680 7400 1840
rect 8080 2010 8240 2050
rect 7470 1680 7510 1840
rect 8810 1680 8850 1840
rect 8080 1470 8240 1510
rect 9360 2010 9520 2050
rect 8920 1680 8960 1840
rect 10040 1680 10080 1840
rect 36820 1140 36980 1180
rect 36160 770 36200 930
rect 37600 770 37640 930
rect 36820 610 36980 650
rect 39340 1140 39500 1180
rect 38680 770 38720 930
rect 40120 770 40160 930
rect 36820 490 36980 530
rect 35680 20 35720 180
rect 38080 20 38120 180
rect 36820 -340 36980 -300
rect 39340 490 39500 530
rect 38200 20 38240 180
rect 40600 20 40640 180
rect 39340 -340 39500 -300
rect 38080 -440 38240 -400
rect 35880 -770 35920 -610
rect 40390 -770 40430 -610
rect 38080 -890 38240 -850
rect 36800 -990 36960 -950
rect 36240 -1320 36280 -1160
rect 37360 -1320 37400 -1160
rect 38080 -990 38240 -950
rect 37470 -1320 37510 -1160
rect 38810 -1320 38850 -1160
rect 38080 -1530 38240 -1490
rect 39360 -990 39520 -950
rect 38920 -1320 38960 -1160
rect 40040 -1320 40080 -1160
rect 45180 -2720 45340 -2680
rect 44050 -3000 44090 -2840
rect 46430 -3000 46470 -2840
rect 45180 -3150 45340 -3110
rect 47690 -2990 47850 -2950
rect 45150 -3250 45310 -3210
rect 44050 -3530 44090 -3370
rect 46370 -3530 46410 -3370
rect 45150 -3680 45310 -3640
rect 46620 -3510 46660 -3350
rect 45150 -3780 45310 -3740
rect 44440 -4000 44480 -3840
rect 46000 -4000 46040 -3840
rect 48970 -3510 49010 -3350
rect 47690 -3900 47850 -3860
rect 45150 -4100 45310 -4060
rect 47690 -4000 47850 -3960
rect 45150 -4200 45310 -4160
rect 33674 -4313 33708 -4279
rect 33764 -4313 33798 -4279
rect 33854 -4313 33888 -4279
rect 33944 -4313 33978 -4279
rect 34034 -4313 34068 -4279
rect 34124 -4313 34158 -4279
rect 34214 -4313 34248 -4279
rect 34304 -4313 34338 -4279
rect 34394 -4313 34428 -4279
rect 34484 -4313 34518 -4279
rect 34574 -4313 34608 -4279
rect 34664 -4313 34698 -4279
rect 34754 -4313 34788 -4279
rect 33651 -4414 33685 -4380
rect 33651 -4504 33685 -4470
rect 33651 -4594 33685 -4560
rect 33651 -4684 33685 -4650
rect 33651 -4774 33685 -4740
rect 33651 -4864 33685 -4830
rect 33651 -4954 33685 -4920
rect 33651 -5044 33685 -5010
rect 33651 -5134 33685 -5100
rect 33651 -5224 33685 -5190
rect 33651 -5314 33685 -5280
rect 33651 -5404 33685 -5370
rect 34838 -4414 34872 -4380
rect 34838 -4504 34872 -4470
rect 34838 -4594 34872 -4560
rect 34838 -4684 34872 -4650
rect 34838 -4774 34872 -4740
rect 34838 -4864 34872 -4830
rect 34838 -4954 34872 -4920
rect 34838 -5044 34872 -5010
rect 34838 -5134 34872 -5100
rect 34838 -5224 34872 -5190
rect 34838 -5314 34872 -5280
rect 34838 -5404 34872 -5370
rect 33674 -5500 33708 -5466
rect 33764 -5500 33798 -5466
rect 33854 -5500 33888 -5466
rect 33944 -5500 33978 -5466
rect 34034 -5500 34068 -5466
rect 34124 -5500 34158 -5466
rect 34214 -5500 34248 -5466
rect 34304 -5500 34338 -5466
rect 34394 -5500 34428 -5466
rect 34484 -5500 34518 -5466
rect 34574 -5500 34608 -5466
rect 34664 -5500 34698 -5466
rect 34754 -5500 34788 -5466
rect 35034 -4313 35068 -4279
rect 35124 -4313 35158 -4279
rect 35214 -4313 35248 -4279
rect 35304 -4313 35338 -4279
rect 35394 -4313 35428 -4279
rect 35484 -4313 35518 -4279
rect 35574 -4313 35608 -4279
rect 35664 -4313 35698 -4279
rect 35754 -4313 35788 -4279
rect 35844 -4313 35878 -4279
rect 35934 -4313 35968 -4279
rect 36024 -4313 36058 -4279
rect 36114 -4313 36148 -4279
rect 35011 -4414 35045 -4380
rect 35011 -4504 35045 -4470
rect 35011 -4594 35045 -4560
rect 35011 -4684 35045 -4650
rect 35011 -4774 35045 -4740
rect 35011 -4864 35045 -4830
rect 35011 -4954 35045 -4920
rect 35011 -5044 35045 -5010
rect 35011 -5134 35045 -5100
rect 35011 -5224 35045 -5190
rect 35011 -5314 35045 -5280
rect 35011 -5404 35045 -5370
rect 36198 -4414 36232 -4380
rect 36198 -4504 36232 -4470
rect 36198 -4594 36232 -4560
rect 36198 -4684 36232 -4650
rect 36198 -4774 36232 -4740
rect 36198 -4864 36232 -4830
rect 36198 -4954 36232 -4920
rect 36198 -5044 36232 -5010
rect 36198 -5134 36232 -5100
rect 36198 -5224 36232 -5190
rect 36198 -5314 36232 -5280
rect 36198 -5404 36232 -5370
rect 35034 -5500 35068 -5466
rect 35124 -5500 35158 -5466
rect 35214 -5500 35248 -5466
rect 35304 -5500 35338 -5466
rect 35394 -5500 35428 -5466
rect 35484 -5500 35518 -5466
rect 35574 -5500 35608 -5466
rect 35664 -5500 35698 -5466
rect 35754 -5500 35788 -5466
rect 35844 -5500 35878 -5466
rect 35934 -5500 35968 -5466
rect 36024 -5500 36058 -5466
rect 36114 -5500 36148 -5466
rect 36394 -4313 36428 -4279
rect 36484 -4313 36518 -4279
rect 36574 -4313 36608 -4279
rect 36664 -4313 36698 -4279
rect 36754 -4313 36788 -4279
rect 36844 -4313 36878 -4279
rect 36934 -4313 36968 -4279
rect 37024 -4313 37058 -4279
rect 37114 -4313 37148 -4279
rect 37204 -4313 37238 -4279
rect 37294 -4313 37328 -4279
rect 37384 -4313 37418 -4279
rect 37474 -4313 37508 -4279
rect 36371 -4414 36405 -4380
rect 36371 -4504 36405 -4470
rect 36371 -4594 36405 -4560
rect 36371 -4684 36405 -4650
rect 36371 -4774 36405 -4740
rect 36371 -4864 36405 -4830
rect 36371 -4954 36405 -4920
rect 36371 -5044 36405 -5010
rect 36371 -5134 36405 -5100
rect 36371 -5224 36405 -5190
rect 36371 -5314 36405 -5280
rect 36371 -5404 36405 -5370
rect 37558 -4414 37592 -4380
rect 37558 -4504 37592 -4470
rect 44440 -4420 44480 -4260
rect 46000 -4420 46040 -4260
rect 46950 -4220 46990 -4060
rect 48560 -4220 48600 -4060
rect 47690 -4310 47850 -4270
rect 45150 -4520 45310 -4480
rect 37558 -4594 37592 -4560
rect 37558 -4684 37592 -4650
rect 37558 -4774 37592 -4740
rect 37558 -4864 37592 -4830
rect 37558 -4954 37592 -4920
rect 37558 -5044 37592 -5010
rect 37558 -5134 37592 -5100
rect 37558 -5224 37592 -5190
rect 37558 -5314 37592 -5280
rect 37558 -5404 37592 -5370
rect 36394 -5500 36428 -5466
rect 36484 -5500 36518 -5466
rect 36574 -5500 36608 -5466
rect 36664 -5500 36698 -5466
rect 36754 -5500 36788 -5466
rect 36844 -5500 36878 -5466
rect 36934 -5500 36968 -5466
rect 37024 -5500 37058 -5466
rect 37114 -5500 37148 -5466
rect 37204 -5500 37238 -5466
rect 37294 -5500 37328 -5466
rect 37384 -5500 37418 -5466
rect 37474 -5500 37508 -5466
rect 33674 -5673 33708 -5639
rect 33764 -5673 33798 -5639
rect 33854 -5673 33888 -5639
rect 33944 -5673 33978 -5639
rect 34034 -5673 34068 -5639
rect 34124 -5673 34158 -5639
rect 34214 -5673 34248 -5639
rect 34304 -5673 34338 -5639
rect 34394 -5673 34428 -5639
rect 34484 -5673 34518 -5639
rect 34574 -5673 34608 -5639
rect 34664 -5673 34698 -5639
rect 34754 -5673 34788 -5639
rect 33651 -5774 33685 -5740
rect 33651 -5864 33685 -5830
rect 33651 -5954 33685 -5920
rect 33651 -6044 33685 -6010
rect 33651 -6134 33685 -6100
rect 33651 -6224 33685 -6190
rect 33651 -6314 33685 -6280
rect 33651 -6404 33685 -6370
rect 33651 -6494 33685 -6460
rect 33651 -6584 33685 -6550
rect 33651 -6674 33685 -6640
rect 33651 -6764 33685 -6730
rect 34838 -5774 34872 -5740
rect 34838 -5864 34872 -5830
rect 34838 -5954 34872 -5920
rect 34838 -6044 34872 -6010
rect 34838 -6134 34872 -6100
rect 34838 -6224 34872 -6190
rect 34838 -6314 34872 -6280
rect 34838 -6404 34872 -6370
rect 34838 -6494 34872 -6460
rect 34838 -6584 34872 -6550
rect 34838 -6674 34872 -6640
rect 34838 -6764 34872 -6730
rect 33674 -6860 33708 -6826
rect 33764 -6860 33798 -6826
rect 33854 -6860 33888 -6826
rect 33944 -6860 33978 -6826
rect 34034 -6860 34068 -6826
rect 34124 -6860 34158 -6826
rect 34214 -6860 34248 -6826
rect 34304 -6860 34338 -6826
rect 34394 -6860 34428 -6826
rect 34484 -6860 34518 -6826
rect 34574 -6860 34608 -6826
rect 34664 -6860 34698 -6826
rect 34754 -6860 34788 -6826
rect 35034 -5673 35068 -5639
rect 35124 -5673 35158 -5639
rect 35214 -5673 35248 -5639
rect 35304 -5673 35338 -5639
rect 35394 -5673 35428 -5639
rect 35484 -5673 35518 -5639
rect 35574 -5673 35608 -5639
rect 35664 -5673 35698 -5639
rect 35754 -5673 35788 -5639
rect 35844 -5673 35878 -5639
rect 35934 -5673 35968 -5639
rect 36024 -5673 36058 -5639
rect 36114 -5673 36148 -5639
rect 35011 -5774 35045 -5740
rect 35011 -5864 35045 -5830
rect 35011 -5954 35045 -5920
rect 35011 -6044 35045 -6010
rect 35011 -6134 35045 -6100
rect 35011 -6224 35045 -6190
rect 35011 -6314 35045 -6280
rect 35011 -6404 35045 -6370
rect 35011 -6494 35045 -6460
rect 35011 -6584 35045 -6550
rect 35011 -6674 35045 -6640
rect 35011 -6764 35045 -6730
rect 36198 -5774 36232 -5740
rect 36198 -5864 36232 -5830
rect 36198 -5954 36232 -5920
rect 36198 -6044 36232 -6010
rect 36198 -6134 36232 -6100
rect 36198 -6224 36232 -6190
rect 36198 -6314 36232 -6280
rect 36198 -6404 36232 -6370
rect 36198 -6494 36232 -6460
rect 36198 -6584 36232 -6550
rect 36198 -6674 36232 -6640
rect 36198 -6764 36232 -6730
rect 35034 -6860 35068 -6826
rect 35124 -6860 35158 -6826
rect 35214 -6860 35248 -6826
rect 35304 -6860 35338 -6826
rect 35394 -6860 35428 -6826
rect 35484 -6860 35518 -6826
rect 35574 -6860 35608 -6826
rect 35664 -6860 35698 -6826
rect 35754 -6860 35788 -6826
rect 35844 -6860 35878 -6826
rect 35934 -6860 35968 -6826
rect 36024 -6860 36058 -6826
rect 36114 -6860 36148 -6826
rect 36394 -5673 36428 -5639
rect 36484 -5673 36518 -5639
rect 36574 -5673 36608 -5639
rect 36664 -5673 36698 -5639
rect 36754 -5673 36788 -5639
rect 36844 -5673 36878 -5639
rect 36934 -5673 36968 -5639
rect 37024 -5673 37058 -5639
rect 37114 -5673 37148 -5639
rect 37204 -5673 37238 -5639
rect 37294 -5673 37328 -5639
rect 37384 -5673 37418 -5639
rect 37474 -5673 37508 -5639
rect 36371 -5774 36405 -5740
rect 36371 -5864 36405 -5830
rect 36371 -5954 36405 -5920
rect 36371 -6044 36405 -6010
rect 36371 -6134 36405 -6100
rect 36371 -6224 36405 -6190
rect 36371 -6314 36405 -6280
rect 36371 -6404 36405 -6370
rect 36371 -6494 36405 -6460
rect 36371 -6584 36405 -6550
rect 36371 -6674 36405 -6640
rect 36371 -6764 36405 -6730
rect 37558 -5774 37592 -5740
rect 37558 -5864 37592 -5830
rect 37558 -5954 37592 -5920
rect 37558 -6044 37592 -6010
rect 37558 -6134 37592 -6100
rect 37558 -6224 37592 -6190
rect 37558 -6314 37592 -6280
rect 37558 -6404 37592 -6370
rect 37558 -6494 37592 -6460
rect 37558 -6584 37592 -6550
rect 37558 -6674 37592 -6640
rect 37558 -6764 37592 -6730
rect 36394 -6860 36428 -6826
rect 36484 -6860 36518 -6826
rect 36574 -6860 36608 -6826
rect 36664 -6860 36698 -6826
rect 36754 -6860 36788 -6826
rect 36844 -6860 36878 -6826
rect 36934 -6860 36968 -6826
rect 37024 -6860 37058 -6826
rect 37114 -6860 37148 -6826
rect 37204 -6860 37238 -6826
rect 37294 -6860 37328 -6826
rect 37384 -6860 37418 -6826
rect 37474 -6860 37508 -6826
rect 33674 -7033 33708 -6999
rect 33764 -7033 33798 -6999
rect 33854 -7033 33888 -6999
rect 33944 -7033 33978 -6999
rect 34034 -7033 34068 -6999
rect 34124 -7033 34158 -6999
rect 34214 -7033 34248 -6999
rect 34304 -7033 34338 -6999
rect 34394 -7033 34428 -6999
rect 34484 -7033 34518 -6999
rect 34574 -7033 34608 -6999
rect 34664 -7033 34698 -6999
rect 34754 -7033 34788 -6999
rect 33651 -7134 33685 -7100
rect 33651 -7224 33685 -7190
rect 33651 -7314 33685 -7280
rect 33651 -7404 33685 -7370
rect 33651 -7494 33685 -7460
rect 33651 -7584 33685 -7550
rect 33651 -7674 33685 -7640
rect 33651 -7764 33685 -7730
rect 33651 -7854 33685 -7820
rect 33651 -7944 33685 -7910
rect 33651 -8034 33685 -8000
rect 33651 -8124 33685 -8090
rect 34838 -7134 34872 -7100
rect 34838 -7224 34872 -7190
rect 34838 -7314 34872 -7280
rect 34838 -7404 34872 -7370
rect 34838 -7494 34872 -7460
rect 34838 -7584 34872 -7550
rect 34838 -7674 34872 -7640
rect 34838 -7764 34872 -7730
rect 34838 -7854 34872 -7820
rect 34838 -7944 34872 -7910
rect 34838 -8034 34872 -8000
rect 34838 -8124 34872 -8090
rect 33674 -8220 33708 -8186
rect 33764 -8220 33798 -8186
rect 33854 -8220 33888 -8186
rect 33944 -8220 33978 -8186
rect 34034 -8220 34068 -8186
rect 34124 -8220 34158 -8186
rect 34214 -8220 34248 -8186
rect 34304 -8220 34338 -8186
rect 34394 -8220 34428 -8186
rect 34484 -8220 34518 -8186
rect 34574 -8220 34608 -8186
rect 34664 -8220 34698 -8186
rect 34754 -8220 34788 -8186
rect 35034 -7033 35068 -6999
rect 35124 -7033 35158 -6999
rect 35214 -7033 35248 -6999
rect 35304 -7033 35338 -6999
rect 35394 -7033 35428 -6999
rect 35484 -7033 35518 -6999
rect 35574 -7033 35608 -6999
rect 35664 -7033 35698 -6999
rect 35754 -7033 35788 -6999
rect 35844 -7033 35878 -6999
rect 35934 -7033 35968 -6999
rect 36024 -7033 36058 -6999
rect 36114 -7033 36148 -6999
rect 35011 -7134 35045 -7100
rect 35011 -7224 35045 -7190
rect 35011 -7314 35045 -7280
rect 35011 -7404 35045 -7370
rect 35011 -7494 35045 -7460
rect 35011 -7584 35045 -7550
rect 35011 -7674 35045 -7640
rect 35011 -7764 35045 -7730
rect 35011 -7854 35045 -7820
rect 35011 -7944 35045 -7910
rect 35011 -8034 35045 -8000
rect 35011 -8124 35045 -8090
rect 36198 -7134 36232 -7100
rect 36198 -7224 36232 -7190
rect 36198 -7314 36232 -7280
rect 36198 -7404 36232 -7370
rect 36198 -7494 36232 -7460
rect 36198 -7584 36232 -7550
rect 36198 -7674 36232 -7640
rect 36198 -7764 36232 -7730
rect 36198 -7854 36232 -7820
rect 36198 -7944 36232 -7910
rect 36198 -8034 36232 -8000
rect 36198 -8124 36232 -8090
rect 35034 -8220 35068 -8186
rect 35124 -8220 35158 -8186
rect 35214 -8220 35248 -8186
rect 35304 -8220 35338 -8186
rect 35394 -8220 35428 -8186
rect 35484 -8220 35518 -8186
rect 35574 -8220 35608 -8186
rect 35664 -8220 35698 -8186
rect 35754 -8220 35788 -8186
rect 35844 -8220 35878 -8186
rect 35934 -8220 35968 -8186
rect 36024 -8220 36058 -8186
rect 36114 -8220 36148 -8186
rect 36394 -7033 36428 -6999
rect 36484 -7033 36518 -6999
rect 36574 -7033 36608 -6999
rect 36664 -7033 36698 -6999
rect 36754 -7033 36788 -6999
rect 36844 -7033 36878 -6999
rect 36934 -7033 36968 -6999
rect 37024 -7033 37058 -6999
rect 37114 -7033 37148 -6999
rect 37204 -7033 37238 -6999
rect 37294 -7033 37328 -6999
rect 37384 -7033 37418 -6999
rect 37474 -7033 37508 -6999
rect 36371 -7134 36405 -7100
rect 36371 -7224 36405 -7190
rect 36371 -7314 36405 -7280
rect 36371 -7404 36405 -7370
rect 36371 -7494 36405 -7460
rect 36371 -7584 36405 -7550
rect 36371 -7674 36405 -7640
rect 36371 -7764 36405 -7730
rect 36371 -7854 36405 -7820
rect 36371 -7944 36405 -7910
rect 36371 -8034 36405 -8000
rect 36371 -8124 36405 -8090
rect 37558 -7134 37592 -7100
rect 37558 -7224 37592 -7190
rect 37558 -7314 37592 -7280
rect 37558 -7404 37592 -7370
rect 37558 -7494 37592 -7460
rect 37558 -7584 37592 -7550
rect 37558 -7674 37592 -7640
rect 37558 -7764 37592 -7730
rect 37558 -7854 37592 -7820
rect 37558 -7944 37592 -7910
rect 37558 -8034 37592 -8000
rect 37558 -8124 37592 -8090
rect 36394 -8220 36428 -8186
rect 36484 -8220 36518 -8186
rect 36574 -8220 36608 -8186
rect 36664 -8220 36698 -8186
rect 36754 -8220 36788 -8186
rect 36844 -8220 36878 -8186
rect 36934 -8220 36968 -8186
rect 37024 -8220 37058 -8186
rect 37114 -8220 37148 -8186
rect 37204 -8220 37238 -8186
rect 37294 -8220 37328 -8186
rect 37384 -8220 37418 -8186
rect 37474 -8220 37508 -8186
rect 35580 -8380 35620 -8340
rect 35580 -8480 35620 -8440
rect 35580 -8580 35620 -8540
<< nsubdiffcont >>
rect 6360 7110 6520 7150
rect 5970 6780 6010 6940
rect 6870 6780 6910 6940
rect 6360 6570 6520 6610
rect 8080 7110 8240 7150
rect 7250 6780 7290 6940
rect 9030 6780 9070 6940
rect 8080 6570 8240 6610
rect 9800 7110 9960 7150
rect 9410 6780 9450 6940
rect 10310 6780 10350 6940
rect 9800 6570 9930 6610
rect 8080 6180 8240 6220
rect 5610 5980 5770 6020
rect 5330 5650 5370 5810
rect 6010 5650 6050 5810
rect 5610 5440 5770 5480
rect 6400 5650 6440 5810
rect 9880 5650 9920 5810
rect 10540 5980 10700 6020
rect 10260 5650 10300 5810
rect 10940 5650 10980 5810
rect 10540 5440 10700 5480
rect 8080 5230 8240 5270
rect 6560 4800 6720 4840
rect 5300 4470 5340 4630
rect 7940 4470 7980 4630
rect 6560 4260 6720 4300
rect 9600 4800 9760 4840
rect 8340 4470 8380 4630
rect 10980 4470 11020 4630
rect 9600 4260 9760 4300
rect 36360 4110 36520 4150
rect 35970 3780 36010 3940
rect 36870 3780 36910 3940
rect 36360 3570 36520 3610
rect 38080 4110 38240 4150
rect 37250 3780 37290 3940
rect 39030 3780 39070 3940
rect 38080 3570 38240 3610
rect 39800 4110 39960 4150
rect 39410 3780 39450 3940
rect 40310 3780 40350 3940
rect 39800 3570 39930 3610
rect 38080 3180 38240 3220
rect 35610 2980 35770 3020
rect 35330 2650 35370 2810
rect 36010 2650 36050 2810
rect 35610 2440 35770 2480
rect 36400 2650 36440 2810
rect 39880 2650 39920 2810
rect 40540 2980 40700 3020
rect 40260 2650 40300 2810
rect 40940 2650 40980 2810
rect 40540 2440 40700 2480
rect 38080 2230 38240 2270
rect 36560 1800 36720 1840
rect 35300 1470 35340 1630
rect 37940 1470 37980 1630
rect 36560 1260 36720 1300
rect 39600 1800 39760 1840
rect 38340 1470 38380 1630
rect 40980 1470 41020 1630
rect 39600 1260 39760 1300
rect 33874 -4462 33908 -4428
rect 33964 -4462 33998 -4428
rect 34054 -4462 34088 -4428
rect 34144 -4462 34178 -4428
rect 34234 -4462 34268 -4428
rect 34324 -4462 34358 -4428
rect 34414 -4462 34448 -4428
rect 34504 -4462 34538 -4428
rect 34594 -4462 34628 -4428
rect 33798 -4520 33832 -4486
rect 33798 -4610 33832 -4576
rect 33798 -4700 33832 -4666
rect 33798 -4790 33832 -4756
rect 33798 -4880 33832 -4846
rect 33798 -4970 33832 -4936
rect 33798 -5060 33832 -5026
rect 33798 -5150 33832 -5116
rect 33798 -5240 33832 -5206
rect 34688 -4554 34722 -4520
rect 34688 -4644 34722 -4610
rect 34688 -4734 34722 -4700
rect 34688 -4824 34722 -4790
rect 34688 -4914 34722 -4880
rect 34688 -5004 34722 -4970
rect 34688 -5094 34722 -5060
rect 34688 -5184 34722 -5150
rect 34688 -5274 34722 -5240
rect 33855 -5352 33889 -5318
rect 33945 -5352 33979 -5318
rect 34035 -5352 34069 -5318
rect 34125 -5352 34159 -5318
rect 34215 -5352 34249 -5318
rect 34305 -5352 34339 -5318
rect 34395 -5352 34429 -5318
rect 34485 -5352 34519 -5318
rect 34575 -5352 34609 -5318
rect 35234 -4462 35268 -4428
rect 35324 -4462 35358 -4428
rect 35414 -4462 35448 -4428
rect 35504 -4462 35538 -4428
rect 35594 -4462 35628 -4428
rect 35684 -4462 35718 -4428
rect 35774 -4462 35808 -4428
rect 35864 -4462 35898 -4428
rect 35954 -4462 35988 -4428
rect 35158 -4520 35192 -4486
rect 35158 -4610 35192 -4576
rect 35158 -4700 35192 -4666
rect 35158 -4790 35192 -4756
rect 35158 -4880 35192 -4846
rect 35158 -4970 35192 -4936
rect 35158 -5060 35192 -5026
rect 35158 -5150 35192 -5116
rect 35158 -5240 35192 -5206
rect 36048 -4554 36082 -4520
rect 36048 -4644 36082 -4610
rect 36048 -4734 36082 -4700
rect 36048 -4824 36082 -4790
rect 36048 -4914 36082 -4880
rect 36048 -5004 36082 -4970
rect 36048 -5094 36082 -5060
rect 36048 -5184 36082 -5150
rect 36048 -5274 36082 -5240
rect 35215 -5352 35249 -5318
rect 35305 -5352 35339 -5318
rect 35395 -5352 35429 -5318
rect 35485 -5352 35519 -5318
rect 35575 -5352 35609 -5318
rect 35665 -5352 35699 -5318
rect 35755 -5352 35789 -5318
rect 35845 -5352 35879 -5318
rect 35935 -5352 35969 -5318
rect 36594 -4462 36628 -4428
rect 36684 -4462 36718 -4428
rect 36774 -4462 36808 -4428
rect 36864 -4462 36898 -4428
rect 36954 -4462 36988 -4428
rect 37044 -4462 37078 -4428
rect 37134 -4462 37168 -4428
rect 37224 -4462 37258 -4428
rect 37314 -4462 37348 -4428
rect 36518 -4520 36552 -4486
rect 36518 -4610 36552 -4576
rect 36518 -4700 36552 -4666
rect 36518 -4790 36552 -4756
rect 36518 -4880 36552 -4846
rect 36518 -4970 36552 -4936
rect 36518 -5060 36552 -5026
rect 36518 -5150 36552 -5116
rect 36518 -5240 36552 -5206
rect 37408 -4554 37442 -4520
rect 37408 -4644 37442 -4610
rect 37408 -4734 37442 -4700
rect 37408 -4824 37442 -4790
rect 37408 -4914 37442 -4880
rect 37408 -5004 37442 -4970
rect 37408 -5094 37442 -5060
rect 37408 -5184 37442 -5150
rect 37408 -5274 37442 -5240
rect 36575 -5352 36609 -5318
rect 36665 -5352 36699 -5318
rect 36755 -5352 36789 -5318
rect 36845 -5352 36879 -5318
rect 36935 -5352 36969 -5318
rect 37025 -5352 37059 -5318
rect 37115 -5352 37149 -5318
rect 37205 -5352 37239 -5318
rect 37295 -5352 37329 -5318
rect 33874 -5822 33908 -5788
rect 33964 -5822 33998 -5788
rect 34054 -5822 34088 -5788
rect 34144 -5822 34178 -5788
rect 34234 -5822 34268 -5788
rect 34324 -5822 34358 -5788
rect 34414 -5822 34448 -5788
rect 34504 -5822 34538 -5788
rect 34594 -5822 34628 -5788
rect 33798 -5880 33832 -5846
rect 33798 -5970 33832 -5936
rect 33798 -6060 33832 -6026
rect 33798 -6150 33832 -6116
rect 33798 -6240 33832 -6206
rect 33798 -6330 33832 -6296
rect 33798 -6420 33832 -6386
rect 33798 -6510 33832 -6476
rect 33798 -6600 33832 -6566
rect 34688 -5914 34722 -5880
rect 34688 -6004 34722 -5970
rect 34688 -6094 34722 -6060
rect 34688 -6184 34722 -6150
rect 34688 -6274 34722 -6240
rect 34688 -6364 34722 -6330
rect 34688 -6454 34722 -6420
rect 34688 -6544 34722 -6510
rect 34688 -6634 34722 -6600
rect 33855 -6712 33889 -6678
rect 33945 -6712 33979 -6678
rect 34035 -6712 34069 -6678
rect 34125 -6712 34159 -6678
rect 34215 -6712 34249 -6678
rect 34305 -6712 34339 -6678
rect 34395 -6712 34429 -6678
rect 34485 -6712 34519 -6678
rect 34575 -6712 34609 -6678
rect 35234 -5822 35268 -5788
rect 35324 -5822 35358 -5788
rect 35414 -5822 35448 -5788
rect 35504 -5822 35538 -5788
rect 35594 -5822 35628 -5788
rect 35684 -5822 35718 -5788
rect 35774 -5822 35808 -5788
rect 35864 -5822 35898 -5788
rect 35954 -5822 35988 -5788
rect 35158 -5880 35192 -5846
rect 35158 -5970 35192 -5936
rect 35158 -6060 35192 -6026
rect 35158 -6150 35192 -6116
rect 35158 -6240 35192 -6206
rect 35158 -6330 35192 -6296
rect 35158 -6420 35192 -6386
rect 35158 -6510 35192 -6476
rect 35158 -6600 35192 -6566
rect 36048 -5914 36082 -5880
rect 36048 -6004 36082 -5970
rect 36048 -6094 36082 -6060
rect 36048 -6184 36082 -6150
rect 36048 -6274 36082 -6240
rect 36048 -6364 36082 -6330
rect 36048 -6454 36082 -6420
rect 36048 -6544 36082 -6510
rect 36048 -6634 36082 -6600
rect 35215 -6712 35249 -6678
rect 35305 -6712 35339 -6678
rect 35395 -6712 35429 -6678
rect 35485 -6712 35519 -6678
rect 35575 -6712 35609 -6678
rect 35665 -6712 35699 -6678
rect 35755 -6712 35789 -6678
rect 35845 -6712 35879 -6678
rect 35935 -6712 35969 -6678
rect 36594 -5822 36628 -5788
rect 36684 -5822 36718 -5788
rect 36774 -5822 36808 -5788
rect 36864 -5822 36898 -5788
rect 36954 -5822 36988 -5788
rect 37044 -5822 37078 -5788
rect 37134 -5822 37168 -5788
rect 37224 -5822 37258 -5788
rect 37314 -5822 37348 -5788
rect 36518 -5880 36552 -5846
rect 36518 -5970 36552 -5936
rect 36518 -6060 36552 -6026
rect 36518 -6150 36552 -6116
rect 36518 -6240 36552 -6206
rect 36518 -6330 36552 -6296
rect 36518 -6420 36552 -6386
rect 36518 -6510 36552 -6476
rect 36518 -6600 36552 -6566
rect 37408 -5914 37442 -5880
rect 37408 -6004 37442 -5970
rect 37408 -6094 37442 -6060
rect 37408 -6184 37442 -6150
rect 37408 -6274 37442 -6240
rect 37408 -6364 37442 -6330
rect 37408 -6454 37442 -6420
rect 37408 -6544 37442 -6510
rect 37408 -6634 37442 -6600
rect 36575 -6712 36609 -6678
rect 36665 -6712 36699 -6678
rect 36755 -6712 36789 -6678
rect 36845 -6712 36879 -6678
rect 36935 -6712 36969 -6678
rect 37025 -6712 37059 -6678
rect 37115 -6712 37149 -6678
rect 37205 -6712 37239 -6678
rect 37295 -6712 37329 -6678
rect 33874 -7182 33908 -7148
rect 33964 -7182 33998 -7148
rect 34054 -7182 34088 -7148
rect 34144 -7182 34178 -7148
rect 34234 -7182 34268 -7148
rect 34324 -7182 34358 -7148
rect 34414 -7182 34448 -7148
rect 34504 -7182 34538 -7148
rect 34594 -7182 34628 -7148
rect 33798 -7240 33832 -7206
rect 33798 -7330 33832 -7296
rect 33798 -7420 33832 -7386
rect 33798 -7510 33832 -7476
rect 33798 -7600 33832 -7566
rect 33798 -7690 33832 -7656
rect 33798 -7780 33832 -7746
rect 33798 -7870 33832 -7836
rect 33798 -7960 33832 -7926
rect 34688 -7274 34722 -7240
rect 34688 -7364 34722 -7330
rect 34688 -7454 34722 -7420
rect 34688 -7544 34722 -7510
rect 34688 -7634 34722 -7600
rect 34688 -7724 34722 -7690
rect 34688 -7814 34722 -7780
rect 34688 -7904 34722 -7870
rect 34688 -7994 34722 -7960
rect 33855 -8072 33889 -8038
rect 33945 -8072 33979 -8038
rect 34035 -8072 34069 -8038
rect 34125 -8072 34159 -8038
rect 34215 -8072 34249 -8038
rect 34305 -8072 34339 -8038
rect 34395 -8072 34429 -8038
rect 34485 -8072 34519 -8038
rect 34575 -8072 34609 -8038
rect 35234 -7182 35268 -7148
rect 35324 -7182 35358 -7148
rect 35414 -7182 35448 -7148
rect 35504 -7182 35538 -7148
rect 35594 -7182 35628 -7148
rect 35684 -7182 35718 -7148
rect 35774 -7182 35808 -7148
rect 35864 -7182 35898 -7148
rect 35954 -7182 35988 -7148
rect 35158 -7240 35192 -7206
rect 35158 -7330 35192 -7296
rect 35158 -7420 35192 -7386
rect 35158 -7510 35192 -7476
rect 35158 -7600 35192 -7566
rect 35158 -7690 35192 -7656
rect 35158 -7780 35192 -7746
rect 35158 -7870 35192 -7836
rect 35158 -7960 35192 -7926
rect 36048 -7274 36082 -7240
rect 36048 -7364 36082 -7330
rect 36048 -7454 36082 -7420
rect 36048 -7544 36082 -7510
rect 36048 -7634 36082 -7600
rect 36048 -7724 36082 -7690
rect 36048 -7814 36082 -7780
rect 36048 -7904 36082 -7870
rect 36048 -7994 36082 -7960
rect 35215 -8072 35249 -8038
rect 35305 -8072 35339 -8038
rect 35395 -8072 35429 -8038
rect 35485 -8072 35519 -8038
rect 35575 -8072 35609 -8038
rect 35665 -8072 35699 -8038
rect 35755 -8072 35789 -8038
rect 35845 -8072 35879 -8038
rect 35935 -8072 35969 -8038
rect 36594 -7182 36628 -7148
rect 36684 -7182 36718 -7148
rect 36774 -7182 36808 -7148
rect 36864 -7182 36898 -7148
rect 36954 -7182 36988 -7148
rect 37044 -7182 37078 -7148
rect 37134 -7182 37168 -7148
rect 37224 -7182 37258 -7148
rect 37314 -7182 37348 -7148
rect 36518 -7240 36552 -7206
rect 36518 -7330 36552 -7296
rect 36518 -7420 36552 -7386
rect 36518 -7510 36552 -7476
rect 36518 -7600 36552 -7566
rect 36518 -7690 36552 -7656
rect 36518 -7780 36552 -7746
rect 36518 -7870 36552 -7836
rect 36518 -7960 36552 -7926
rect 37408 -7274 37442 -7240
rect 37408 -7364 37442 -7330
rect 37408 -7454 37442 -7420
rect 37408 -7544 37442 -7510
rect 37408 -7634 37442 -7600
rect 37408 -7724 37442 -7690
rect 37408 -7814 37442 -7780
rect 37408 -7904 37442 -7870
rect 37408 -7994 37442 -7960
rect 36575 -8072 36609 -8038
rect 36665 -8072 36699 -8038
rect 36755 -8072 36789 -8038
rect 36845 -8072 36879 -8038
rect 36935 -8072 36969 -8038
rect 37025 -8072 37059 -8038
rect 37115 -8072 37149 -8038
rect 37205 -8072 37239 -8038
rect 37295 -8072 37329 -8038
<< poly >>
rect 6070 7050 6150 7070
rect 6070 7010 6090 7050
rect 6130 7020 6150 7050
rect 6410 7050 6470 7070
rect 6130 7010 6180 7020
rect 6410 7010 6420 7050
rect 6460 7010 6470 7050
rect 6730 7050 6810 7070
rect 6730 7010 6750 7050
rect 6790 7010 6810 7050
rect 6070 6990 6180 7010
rect 6150 6960 6180 6990
rect 6260 6980 6620 7010
rect 6260 6960 6290 6980
rect 6370 6960 6400 6980
rect 6480 6960 6510 6980
rect 6590 6960 6620 6980
rect 6700 6980 6810 7010
rect 6700 6960 6730 6980
rect 6150 6730 6180 6760
rect 6260 6730 6290 6760
rect 6370 6730 6400 6760
rect 6480 6730 6510 6760
rect 6590 6730 6620 6760
rect 6700 6730 6730 6760
rect 7350 7050 7430 7070
rect 7350 7010 7370 7050
rect 7410 7020 7430 7050
rect 8130 7050 8190 7070
rect 7410 7010 7460 7020
rect 8130 7010 8140 7050
rect 8180 7010 8190 7050
rect 8670 7050 8750 7070
rect 8670 7020 8690 7050
rect 8640 7010 8690 7020
rect 8730 7010 8750 7050
rect 7350 6990 7460 7010
rect 7430 6960 7460 6990
rect 7540 6980 8560 7010
rect 7540 6960 7570 6980
rect 7650 6960 7680 6980
rect 7760 6960 7790 6980
rect 7870 6960 7900 6980
rect 7980 6960 8010 6980
rect 8090 6960 8120 6980
rect 8200 6960 8230 6980
rect 8310 6960 8340 6980
rect 8420 6960 8450 6980
rect 8530 6960 8560 6980
rect 8640 6990 8750 7010
rect 8640 6960 8670 6990
rect 7430 6730 7460 6760
rect 7540 6730 7570 6760
rect 7650 6730 7680 6760
rect 7760 6730 7790 6760
rect 7870 6730 7900 6760
rect 7980 6730 8010 6760
rect 8090 6730 8120 6760
rect 8200 6730 8230 6760
rect 8310 6730 8340 6760
rect 8420 6730 8450 6760
rect 8530 6730 8560 6760
rect 8640 6730 8670 6760
rect 9510 7050 9590 7070
rect 9510 7010 9530 7050
rect 9570 7020 9590 7050
rect 9850 7050 9910 7070
rect 9570 7010 9620 7020
rect 9850 7010 9860 7050
rect 9900 7010 9910 7050
rect 10170 7050 10250 7070
rect 10170 7020 10190 7050
rect 10140 7010 10190 7020
rect 10230 7010 10250 7050
rect 9510 6990 9620 7010
rect 9590 6960 9620 6990
rect 9700 6980 10060 7010
rect 9700 6960 9730 6980
rect 9810 6960 9840 6980
rect 9920 6960 9950 6980
rect 10030 6960 10060 6980
rect 10140 6990 10250 7010
rect 10140 6960 10170 6990
rect 9590 6730 9620 6760
rect 9700 6730 9730 6760
rect 9810 6730 9840 6760
rect 9920 6730 9950 6760
rect 10030 6730 10060 6760
rect 10140 6730 10170 6760
rect 5440 5920 5500 5940
rect 5440 5880 5450 5920
rect 5490 5880 5500 5920
rect 5880 5920 5940 5940
rect 5880 5880 5890 5920
rect 5930 5880 5940 5920
rect 5440 5850 5540 5880
rect 5510 5830 5540 5850
rect 5620 5830 5650 5860
rect 5730 5830 5760 5860
rect 5840 5850 5940 5880
rect 5840 5830 5870 5850
rect 5510 5600 5540 5630
rect 5620 5610 5650 5630
rect 5730 5610 5760 5630
rect 5620 5580 5760 5610
rect 5840 5600 5870 5630
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 6500 6120 6580 6140
rect 6500 6080 6520 6120
rect 6560 6090 6580 6120
rect 9740 6120 9820 6140
rect 9740 6090 9760 6120
rect 6560 6080 6680 6090
rect 6500 6060 6680 6080
rect 9640 6080 9760 6090
rect 9800 6080 9820 6120
rect 9640 6060 9820 6080
rect 6580 6030 6680 6060
rect 6760 6030 6860 6060
rect 6940 6030 7040 6060
rect 7120 6030 7220 6060
rect 7300 6030 7400 6060
rect 7480 6030 7580 6060
rect 7660 6030 7760 6060
rect 7840 6030 7940 6060
rect 8020 6030 8120 6060
rect 8200 6030 8300 6060
rect 8380 6030 8480 6060
rect 8560 6030 8660 6060
rect 8740 6030 8840 6060
rect 8920 6030 9020 6060
rect 9100 6030 9200 6060
rect 9280 6030 9380 6060
rect 9460 6030 9560 6060
rect 9640 6030 9740 6060
rect 6580 5400 6680 5430
rect 6760 5410 6860 5430
rect 6940 5410 7040 5430
rect 7120 5410 7220 5430
rect 7300 5410 7400 5430
rect 7480 5410 7580 5430
rect 7660 5410 7760 5430
rect 7840 5410 7940 5430
rect 8020 5410 8120 5430
rect 8200 5410 8300 5430
rect 8380 5410 8480 5430
rect 8560 5410 8660 5430
rect 8740 5410 8840 5430
rect 8920 5410 9020 5430
rect 9100 5410 9200 5430
rect 9280 5410 9380 5430
rect 9460 5410 9560 5430
rect 6760 5380 9560 5410
rect 9640 5400 9740 5430
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 10370 5920 10430 5940
rect 10370 5880 10380 5920
rect 10420 5890 10430 5920
rect 10810 5920 10870 5940
rect 10810 5890 10820 5920
rect 10420 5880 10470 5890
rect 10370 5860 10470 5880
rect 10770 5880 10820 5890
rect 10860 5880 10870 5920
rect 10770 5860 10870 5880
rect 10440 5830 10470 5860
rect 10550 5830 10580 5860
rect 10660 5830 10690 5860
rect 10770 5830 10800 5860
rect 10440 5600 10470 5630
rect 10550 5610 10580 5630
rect 10660 5610 10690 5630
rect 10550 5580 10690 5610
rect 10770 5600 10800 5630
rect 10580 5540 10600 5580
rect 10640 5540 10660 5580
rect 10580 5520 10660 5540
rect 5480 4650 5520 4680
rect 5600 4650 5640 4680
rect 5720 4650 5760 4680
rect 5840 4650 5880 4680
rect 5960 4650 6000 4680
rect 6080 4650 6120 4680
rect 6200 4650 6240 4680
rect 6320 4650 6360 4680
rect 6440 4650 6480 4680
rect 6560 4650 6600 4680
rect 6680 4650 6720 4680
rect 6800 4650 6840 4680
rect 6920 4650 6960 4680
rect 7040 4650 7080 4680
rect 7160 4650 7200 4680
rect 7280 4650 7320 4680
rect 7400 4650 7440 4680
rect 7520 4650 7560 4680
rect 7640 4650 7680 4680
rect 7760 4650 7800 4680
rect 5480 4430 5520 4450
rect 5410 4400 5520 4430
rect 5600 4420 5640 4450
rect 5720 4430 5760 4450
rect 5840 4430 5880 4450
rect 5960 4430 6000 4450
rect 6080 4430 6120 4450
rect 5580 4400 5660 4420
rect 5720 4400 6120 4430
rect 6200 4430 6240 4450
rect 6320 4430 6360 4450
rect 6200 4400 6360 4430
rect 6440 4430 6480 4450
rect 6560 4430 6600 4450
rect 6680 4430 6720 4450
rect 6800 4430 6840 4450
rect 6440 4400 6840 4430
rect 6920 4430 6960 4450
rect 7040 4430 7080 4450
rect 6920 4400 7080 4430
rect 7160 4430 7200 4450
rect 7280 4430 7320 4450
rect 7400 4430 7440 4450
rect 7520 4430 7560 4450
rect 7160 4400 7560 4430
rect 7640 4420 7680 4450
rect 7760 4430 7800 4450
rect 7630 4400 7690 4420
rect 7760 4400 7870 4430
rect 5410 4360 5420 4400
rect 5460 4360 5470 4400
rect 5410 4340 5470 4360
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4360 5780 4400
rect 5820 4360 5840 4400
rect 5760 4340 5840 4360
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4360 6500 4400
rect 6540 4360 6560 4400
rect 6480 4340 6560 4360
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4360 7220 4400
rect 7260 4360 7280 4400
rect 7200 4340 7280 4360
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 7810 4360 7820 4400
rect 7860 4360 7870 4400
rect 7810 4340 7870 4360
rect 8520 4650 8560 4680
rect 8640 4650 8680 4680
rect 8760 4650 8800 4680
rect 8880 4650 8920 4680
rect 9000 4650 9040 4680
rect 9120 4650 9160 4680
rect 9240 4650 9280 4680
rect 9360 4650 9400 4680
rect 9480 4650 9520 4680
rect 9600 4650 9640 4680
rect 9720 4650 9760 4680
rect 9840 4650 9880 4680
rect 9960 4650 10000 4680
rect 10080 4650 10120 4680
rect 10200 4650 10240 4680
rect 10320 4650 10360 4680
rect 10440 4650 10480 4680
rect 10560 4650 10600 4680
rect 10680 4650 10720 4680
rect 10800 4650 10840 4680
rect 8520 4430 8560 4450
rect 8450 4400 8560 4430
rect 8640 4420 8680 4450
rect 8760 4430 8800 4450
rect 8880 4430 8920 4450
rect 9000 4430 9040 4450
rect 9120 4430 9160 4450
rect 8630 4400 8690 4420
rect 8760 4400 9160 4430
rect 9240 4430 9280 4450
rect 9360 4430 9400 4450
rect 9240 4400 9400 4430
rect 9480 4430 9520 4450
rect 9600 4430 9640 4450
rect 9720 4430 9760 4450
rect 9840 4430 9880 4450
rect 9480 4400 9880 4430
rect 9960 4430 10000 4450
rect 10080 4430 10120 4450
rect 9960 4400 10120 4430
rect 10200 4430 10240 4450
rect 10320 4430 10360 4450
rect 10440 4430 10480 4450
rect 10560 4430 10600 4450
rect 10200 4400 10600 4430
rect 10680 4420 10720 4450
rect 10800 4430 10840 4450
rect 10660 4400 10740 4420
rect 10800 4400 10910 4430
rect 8450 4360 8460 4400
rect 8500 4360 8510 4400
rect 8450 4340 8510 4360
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 9040 4360 9060 4400
rect 9100 4360 9120 4400
rect 9040 4340 9120 4360
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9760 4360 9780 4400
rect 9820 4360 9840 4400
rect 9760 4340 9840 4360
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10480 4360 10500 4400
rect 10540 4360 10560 4400
rect 10480 4340 10560 4360
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 10850 4360 10860 4400
rect 10900 4360 10910 4400
rect 10850 4340 10910 4360
rect 6380 4080 6460 4100
rect 6380 4040 6400 4080
rect 6440 4040 6460 4080
rect 6380 4010 6460 4040
rect 6380 3980 7460 4010
rect 6340 3900 6380 3930
rect 6460 3900 6500 3980
rect 6580 3900 6620 3980
rect 6700 3900 6740 3930
rect 6820 3900 6860 3930
rect 6940 3900 6980 3980
rect 7060 3900 7100 3980
rect 7180 3900 7220 3930
rect 7300 3900 7340 3930
rect 7420 3900 7460 3980
rect 6340 3770 6380 3800
rect 6460 3770 6500 3800
rect 6580 3770 6620 3800
rect 6260 3750 6380 3770
rect 6260 3710 6280 3750
rect 6320 3720 6380 3750
rect 6700 3720 6740 3800
rect 6820 3720 6860 3800
rect 6940 3770 6980 3800
rect 7060 3770 7100 3800
rect 7180 3720 7220 3800
rect 7300 3720 7340 3800
rect 7420 3770 7460 3800
rect 6320 3710 7340 3720
rect 6260 3690 7340 3710
rect 9860 4080 9940 4100
rect 9860 4040 9880 4080
rect 9920 4040 9940 4080
rect 9860 4010 9940 4040
rect 8860 3980 9940 4010
rect 8860 3900 8900 3980
rect 8980 3900 9020 3930
rect 9100 3900 9140 3930
rect 9220 3900 9260 3980
rect 9340 3900 9380 3980
rect 9460 3900 9500 3930
rect 9580 3900 9620 3930
rect 9700 3900 9740 3980
rect 9820 3900 9860 3980
rect 9940 3900 9980 3930
rect 8860 3770 8900 3800
rect 8980 3720 9020 3800
rect 9100 3720 9140 3800
rect 9220 3770 9260 3800
rect 9340 3770 9380 3800
rect 9460 3720 9500 3800
rect 9580 3720 9620 3800
rect 9700 3770 9740 3800
rect 9820 3770 9860 3800
rect 9940 3770 9980 3800
rect 9940 3750 10060 3770
rect 9940 3720 10000 3750
rect 8980 3710 10000 3720
rect 10040 3710 10060 3750
rect 8980 3690 10060 3710
rect 36070 4050 36150 4070
rect 36070 4010 36090 4050
rect 36130 4020 36150 4050
rect 36410 4050 36470 4070
rect 36130 4010 36180 4020
rect 36410 4010 36420 4050
rect 36460 4010 36470 4050
rect 36730 4050 36810 4070
rect 36730 4010 36750 4050
rect 36790 4010 36810 4050
rect 36070 3990 36180 4010
rect 36150 3960 36180 3990
rect 36260 3980 36620 4010
rect 36260 3960 36290 3980
rect 36370 3960 36400 3980
rect 36480 3960 36510 3980
rect 36590 3960 36620 3980
rect 36700 3980 36810 4010
rect 36700 3960 36730 3980
rect 36150 3730 36180 3760
rect 36260 3730 36290 3760
rect 36370 3730 36400 3760
rect 36480 3730 36510 3760
rect 36590 3730 36620 3760
rect 36700 3730 36730 3760
rect 37350 4050 37430 4070
rect 37350 4010 37370 4050
rect 37410 4020 37430 4050
rect 38130 4050 38190 4070
rect 37410 4010 37460 4020
rect 38130 4010 38140 4050
rect 38180 4010 38190 4050
rect 38670 4050 38750 4070
rect 38670 4020 38690 4050
rect 38640 4010 38690 4020
rect 38730 4010 38750 4050
rect 37350 3990 37460 4010
rect 37430 3960 37460 3990
rect 37540 3980 38560 4010
rect 37540 3960 37570 3980
rect 37650 3960 37680 3980
rect 37760 3960 37790 3980
rect 37870 3960 37900 3980
rect 37980 3960 38010 3980
rect 38090 3960 38120 3980
rect 38200 3960 38230 3980
rect 38310 3960 38340 3980
rect 38420 3960 38450 3980
rect 38530 3960 38560 3980
rect 38640 3990 38750 4010
rect 38640 3960 38670 3990
rect 37430 3730 37460 3760
rect 37540 3730 37570 3760
rect 37650 3730 37680 3760
rect 37760 3730 37790 3760
rect 37870 3730 37900 3760
rect 37980 3730 38010 3760
rect 38090 3730 38120 3760
rect 38200 3730 38230 3760
rect 38310 3730 38340 3760
rect 38420 3730 38450 3760
rect 38530 3730 38560 3760
rect 38640 3730 38670 3760
rect 39510 4050 39590 4070
rect 39510 4010 39530 4050
rect 39570 4020 39590 4050
rect 39850 4050 39910 4070
rect 39570 4010 39620 4020
rect 39850 4010 39860 4050
rect 39900 4010 39910 4050
rect 40170 4050 40250 4070
rect 40170 4020 40190 4050
rect 40140 4010 40190 4020
rect 40230 4010 40250 4050
rect 39510 3990 39620 4010
rect 39590 3960 39620 3990
rect 39700 3980 40060 4010
rect 39700 3960 39730 3980
rect 39810 3960 39840 3980
rect 39920 3960 39950 3980
rect 40030 3960 40060 3980
rect 40140 3990 40250 4010
rect 40140 3960 40170 3990
rect 39590 3730 39620 3760
rect 39700 3730 39730 3760
rect 39810 3730 39840 3760
rect 39920 3730 39950 3760
rect 40030 3730 40060 3760
rect 40140 3730 40170 3760
rect 5960 3430 6040 3450
rect 5960 3390 5980 3430
rect 6020 3390 6040 3430
rect 5960 3380 6040 3390
rect 6200 3430 6280 3450
rect 6200 3390 6220 3430
rect 6260 3390 6280 3430
rect 6200 3380 6280 3390
rect 6440 3430 6520 3450
rect 6440 3390 6460 3430
rect 6500 3390 6520 3430
rect 6440 3380 6520 3390
rect 6680 3430 6760 3450
rect 6680 3390 6700 3430
rect 6740 3390 6760 3430
rect 6680 3380 6760 3390
rect 7160 3430 7240 3450
rect 7160 3390 7180 3430
rect 7220 3390 7240 3430
rect 7160 3380 7240 3390
rect 7400 3430 7480 3450
rect 7400 3390 7420 3430
rect 7460 3390 7480 3430
rect 7400 3380 7480 3390
rect 7640 3430 7720 3450
rect 7640 3390 7660 3430
rect 7700 3390 7720 3430
rect 7640 3380 7720 3390
rect 5860 3350 6860 3380
rect 6940 3350 7940 3380
rect 5860 2820 6860 2850
rect 6940 2820 7940 2850
rect 8600 3430 8680 3450
rect 8600 3390 8620 3430
rect 8660 3390 8680 3430
rect 8600 3380 8680 3390
rect 8840 3430 8920 3450
rect 8840 3390 8860 3430
rect 8900 3390 8920 3430
rect 8840 3380 8920 3390
rect 9080 3430 9160 3450
rect 9080 3390 9100 3430
rect 9140 3390 9160 3430
rect 9080 3380 9160 3390
rect 9560 3430 9640 3450
rect 9560 3390 9580 3430
rect 9620 3390 9640 3430
rect 9560 3380 9640 3390
rect 9800 3430 9880 3450
rect 9800 3390 9820 3430
rect 9860 3390 9880 3430
rect 9800 3380 9880 3390
rect 10040 3430 10120 3450
rect 10040 3390 10060 3430
rect 10100 3390 10120 3430
rect 10040 3380 10120 3390
rect 10280 3430 10360 3450
rect 10280 3390 10300 3430
rect 10340 3390 10360 3430
rect 10280 3380 10360 3390
rect 8380 3350 9380 3380
rect 9460 3350 10460 3380
rect 8380 2820 9380 2850
rect 9460 2820 10460 2850
rect 35440 2920 35500 2940
rect 35440 2880 35450 2920
rect 35490 2880 35500 2920
rect 35880 2920 35940 2940
rect 35880 2880 35890 2920
rect 35930 2880 35940 2920
rect 35440 2850 35540 2880
rect 35510 2830 35540 2850
rect 35620 2830 35650 2860
rect 35730 2830 35760 2860
rect 35840 2850 35940 2880
rect 35840 2830 35870 2850
rect 6200 2500 6280 2520
rect 6200 2460 6220 2500
rect 6260 2460 6280 2500
rect 6200 2440 6280 2460
rect 6360 2500 6440 2520
rect 6360 2460 6380 2500
rect 6420 2460 6440 2500
rect 6360 2440 6440 2460
rect 6520 2500 6600 2520
rect 6520 2460 6540 2500
rect 6580 2460 6600 2500
rect 6520 2440 6600 2460
rect 6680 2500 6760 2520
rect 6680 2460 6700 2500
rect 6740 2460 6760 2500
rect 6680 2440 6760 2460
rect 6840 2500 6920 2520
rect 6840 2460 6860 2500
rect 6900 2460 6920 2500
rect 6840 2440 6920 2460
rect 7000 2500 7080 2520
rect 7000 2460 7020 2500
rect 7060 2460 7080 2500
rect 7000 2440 7080 2460
rect 7160 2500 7240 2520
rect 7160 2460 7180 2500
rect 7220 2460 7240 2500
rect 7160 2440 7240 2460
rect 7320 2500 7400 2520
rect 7320 2460 7340 2500
rect 7380 2460 7400 2500
rect 7320 2440 7400 2460
rect 7480 2500 7560 2520
rect 7480 2460 7500 2500
rect 7540 2460 7560 2500
rect 7480 2440 7560 2460
rect 7640 2500 7720 2520
rect 7640 2460 7660 2500
rect 7700 2460 7720 2500
rect 7640 2440 7720 2460
rect 7800 2500 7880 2520
rect 7800 2460 7820 2500
rect 7860 2460 7880 2500
rect 7800 2440 7880 2460
rect 7960 2500 8040 2520
rect 7960 2460 7980 2500
rect 8020 2460 8040 2500
rect 7960 2440 8040 2460
rect 8280 2500 8360 2520
rect 8280 2460 8300 2500
rect 8340 2460 8360 2500
rect 8280 2440 8360 2460
rect 8440 2500 8520 2520
rect 8440 2460 8460 2500
rect 8500 2460 8520 2500
rect 8440 2440 8520 2460
rect 8600 2500 8680 2520
rect 8600 2460 8620 2500
rect 8660 2460 8680 2500
rect 8600 2440 8680 2460
rect 8760 2500 8840 2520
rect 8760 2460 8780 2500
rect 8820 2460 8840 2500
rect 8760 2440 8840 2460
rect 8920 2500 9000 2520
rect 8920 2460 8940 2500
rect 8980 2460 9000 2500
rect 8920 2440 9000 2460
rect 9080 2500 9160 2520
rect 9080 2460 9100 2500
rect 9140 2460 9160 2500
rect 9080 2440 9160 2460
rect 9240 2500 9320 2520
rect 9240 2460 9260 2500
rect 9300 2460 9320 2500
rect 9240 2440 9320 2460
rect 9400 2500 9480 2520
rect 9400 2460 9420 2500
rect 9460 2460 9480 2500
rect 9400 2440 9480 2460
rect 9560 2500 9640 2520
rect 9560 2460 9580 2500
rect 9620 2460 9640 2500
rect 9560 2440 9640 2460
rect 9720 2500 9800 2520
rect 9720 2460 9740 2500
rect 9780 2460 9800 2500
rect 9720 2440 9800 2460
rect 9880 2500 9960 2520
rect 9880 2460 9900 2500
rect 9940 2460 9960 2500
rect 9880 2440 9960 2460
rect 10040 2500 10120 2520
rect 10040 2460 10060 2500
rect 10100 2460 10120 2500
rect 10040 2440 10120 2460
rect 6120 2410 8120 2440
rect 8200 2410 10200 2440
rect 35510 2600 35540 2630
rect 35620 2610 35650 2630
rect 35730 2610 35760 2630
rect 35620 2580 35760 2610
rect 35840 2600 35870 2630
rect 35650 2540 35670 2580
rect 35710 2540 35730 2580
rect 35650 2520 35730 2540
rect 36500 3120 36580 3140
rect 36500 3080 36520 3120
rect 36560 3090 36580 3120
rect 39740 3120 39820 3140
rect 39740 3090 39760 3120
rect 36560 3080 36680 3090
rect 36500 3060 36680 3080
rect 39640 3080 39760 3090
rect 39800 3080 39820 3120
rect 39640 3060 39820 3080
rect 36580 3030 36680 3060
rect 36760 3030 36860 3060
rect 36940 3030 37040 3060
rect 37120 3030 37220 3060
rect 37300 3030 37400 3060
rect 37480 3030 37580 3060
rect 37660 3030 37760 3060
rect 37840 3030 37940 3060
rect 38020 3030 38120 3060
rect 38200 3030 38300 3060
rect 38380 3030 38480 3060
rect 38560 3030 38660 3060
rect 38740 3030 38840 3060
rect 38920 3030 39020 3060
rect 39100 3030 39200 3060
rect 39280 3030 39380 3060
rect 39460 3030 39560 3060
rect 39640 3030 39740 3060
rect 36580 2400 36680 2430
rect 36760 2410 36860 2430
rect 36940 2410 37040 2430
rect 37120 2410 37220 2430
rect 37300 2410 37400 2430
rect 37480 2410 37580 2430
rect 37660 2410 37760 2430
rect 37840 2410 37940 2430
rect 38020 2410 38120 2430
rect 38200 2410 38300 2430
rect 38380 2410 38480 2430
rect 38560 2410 38660 2430
rect 38740 2410 38840 2430
rect 38920 2410 39020 2430
rect 39100 2410 39200 2430
rect 39280 2410 39380 2430
rect 39460 2410 39560 2430
rect 36760 2380 39560 2410
rect 39640 2400 39740 2430
rect 37940 2340 37960 2380
rect 38000 2340 38020 2380
rect 37940 2320 38020 2340
rect 39380 2340 39400 2380
rect 39440 2340 39460 2380
rect 39380 2320 39460 2340
rect 40370 2920 40430 2940
rect 40370 2880 40380 2920
rect 40420 2890 40430 2920
rect 40810 2920 40870 2940
rect 40810 2890 40820 2920
rect 40420 2880 40470 2890
rect 40370 2860 40470 2880
rect 40770 2880 40820 2890
rect 40860 2880 40870 2920
rect 40770 2860 40870 2880
rect 40440 2830 40470 2860
rect 40550 2830 40580 2860
rect 40660 2830 40690 2860
rect 40770 2830 40800 2860
rect 40440 2600 40470 2630
rect 40550 2610 40580 2630
rect 40660 2610 40690 2630
rect 40550 2580 40690 2610
rect 40770 2600 40800 2630
rect 40580 2540 40600 2580
rect 40640 2540 40660 2580
rect 40580 2520 40660 2540
rect 6120 2180 8120 2210
rect 8200 2180 10200 2210
rect 6900 1950 6960 1970
rect 6900 1910 6910 1950
rect 6950 1910 6960 1950
rect 6420 1860 6450 1890
rect 6530 1880 7110 1910
rect 6530 1860 6560 1880
rect 6640 1860 6670 1880
rect 6750 1860 6780 1880
rect 6860 1860 6890 1880
rect 6970 1860 7000 1880
rect 7080 1860 7110 1880
rect 7190 1860 7220 1890
rect 6420 1640 6450 1660
rect 6350 1610 6450 1640
rect 6530 1630 6560 1660
rect 6640 1630 6670 1660
rect 6750 1630 6780 1660
rect 6860 1630 6890 1660
rect 6970 1630 7000 1660
rect 7080 1630 7110 1660
rect 7190 1640 7220 1660
rect 7190 1610 7290 1640
rect 6350 1570 6360 1610
rect 6400 1570 6410 1610
rect 6350 1550 6410 1570
rect 7230 1570 7240 1610
rect 7280 1570 7290 1610
rect 7230 1550 7290 1570
rect 8130 1950 8190 1970
rect 8130 1910 8140 1950
rect 8180 1910 8190 1950
rect 7650 1860 7680 1890
rect 7760 1880 8560 1910
rect 7760 1860 7790 1880
rect 7870 1860 7900 1880
rect 7980 1860 8010 1880
rect 8090 1860 8120 1880
rect 8200 1860 8230 1880
rect 8310 1860 8340 1880
rect 8420 1860 8450 1880
rect 8530 1860 8560 1880
rect 8640 1860 8670 1890
rect 7650 1640 7680 1660
rect 7580 1610 7680 1640
rect 7760 1630 7790 1660
rect 7870 1630 7900 1660
rect 7980 1630 8010 1660
rect 8090 1630 8120 1660
rect 8200 1630 8230 1660
rect 8310 1630 8340 1660
rect 8420 1630 8450 1660
rect 8530 1630 8560 1660
rect 8640 1640 8670 1660
rect 7730 1610 7810 1630
rect 8640 1610 8740 1640
rect 7580 1570 7590 1610
rect 7630 1570 7640 1610
rect 7580 1550 7640 1570
rect 7730 1570 7750 1610
rect 7790 1570 7810 1610
rect 7730 1550 7810 1570
rect 8680 1570 8690 1610
rect 8730 1570 8740 1610
rect 8680 1550 8740 1570
rect 9360 1950 9420 1970
rect 9360 1910 9370 1950
rect 9410 1910 9420 1950
rect 9100 1860 9130 1890
rect 9210 1880 9790 1910
rect 9210 1860 9240 1880
rect 9320 1860 9350 1880
rect 9430 1860 9460 1880
rect 9540 1860 9570 1880
rect 9650 1860 9680 1880
rect 9760 1860 9790 1880
rect 9870 1860 9900 1890
rect 9100 1640 9130 1660
rect 9030 1610 9130 1640
rect 9210 1630 9240 1660
rect 9320 1630 9350 1660
rect 9430 1630 9460 1660
rect 9540 1630 9570 1660
rect 9650 1630 9680 1660
rect 9760 1630 9790 1660
rect 9870 1640 9900 1660
rect 9870 1610 9970 1640
rect 9030 1570 9040 1610
rect 9080 1570 9090 1610
rect 9030 1550 9090 1570
rect 9910 1570 9920 1610
rect 9960 1570 9970 1610
rect 9910 1550 9970 1570
rect 35480 1650 35520 1680
rect 35600 1650 35640 1680
rect 35720 1650 35760 1680
rect 35840 1650 35880 1680
rect 35960 1650 36000 1680
rect 36080 1650 36120 1680
rect 36200 1650 36240 1680
rect 36320 1650 36360 1680
rect 36440 1650 36480 1680
rect 36560 1650 36600 1680
rect 36680 1650 36720 1680
rect 36800 1650 36840 1680
rect 36920 1650 36960 1680
rect 37040 1650 37080 1680
rect 37160 1650 37200 1680
rect 37280 1650 37320 1680
rect 37400 1650 37440 1680
rect 37520 1650 37560 1680
rect 37640 1650 37680 1680
rect 37760 1650 37800 1680
rect 35480 1430 35520 1450
rect 35410 1400 35520 1430
rect 35600 1420 35640 1450
rect 35720 1430 35760 1450
rect 35840 1430 35880 1450
rect 35960 1430 36000 1450
rect 36080 1430 36120 1450
rect 35580 1400 35660 1420
rect 35720 1400 36120 1430
rect 36200 1430 36240 1450
rect 36320 1430 36360 1450
rect 36200 1400 36360 1430
rect 36440 1430 36480 1450
rect 36560 1430 36600 1450
rect 36680 1430 36720 1450
rect 36800 1430 36840 1450
rect 36440 1400 36840 1430
rect 36920 1430 36960 1450
rect 37040 1430 37080 1450
rect 36920 1400 37080 1430
rect 37160 1430 37200 1450
rect 37280 1430 37320 1450
rect 37400 1430 37440 1450
rect 37520 1430 37560 1450
rect 37160 1400 37560 1430
rect 37640 1420 37680 1450
rect 37760 1430 37800 1450
rect 37630 1400 37690 1420
rect 37760 1400 37870 1430
rect 35410 1360 35420 1400
rect 35460 1360 35470 1400
rect 35410 1340 35470 1360
rect 35580 1360 35600 1400
rect 35640 1360 35660 1400
rect 35580 1340 35660 1360
rect 35760 1360 35780 1400
rect 35820 1360 35840 1400
rect 35760 1340 35840 1360
rect 36240 1360 36260 1400
rect 36300 1360 36320 1400
rect 36240 1340 36320 1360
rect 36480 1360 36500 1400
rect 36540 1360 36560 1400
rect 36480 1340 36560 1360
rect 36960 1360 36980 1400
rect 37020 1360 37040 1400
rect 36960 1340 37040 1360
rect 37200 1360 37220 1400
rect 37260 1360 37280 1400
rect 37200 1340 37280 1360
rect 37630 1360 37640 1400
rect 37680 1360 37690 1400
rect 37630 1340 37690 1360
rect 37810 1360 37820 1400
rect 37860 1360 37870 1400
rect 37810 1340 37870 1360
rect 38520 1650 38560 1680
rect 38640 1650 38680 1680
rect 38760 1650 38800 1680
rect 38880 1650 38920 1680
rect 39000 1650 39040 1680
rect 39120 1650 39160 1680
rect 39240 1650 39280 1680
rect 39360 1650 39400 1680
rect 39480 1650 39520 1680
rect 39600 1650 39640 1680
rect 39720 1650 39760 1680
rect 39840 1650 39880 1680
rect 39960 1650 40000 1680
rect 40080 1650 40120 1680
rect 40200 1650 40240 1680
rect 40320 1650 40360 1680
rect 40440 1650 40480 1680
rect 40560 1650 40600 1680
rect 40680 1650 40720 1680
rect 40800 1650 40840 1680
rect 38520 1430 38560 1450
rect 38450 1400 38560 1430
rect 38640 1420 38680 1450
rect 38760 1430 38800 1450
rect 38880 1430 38920 1450
rect 39000 1430 39040 1450
rect 39120 1430 39160 1450
rect 38630 1400 38690 1420
rect 38760 1400 39160 1430
rect 39240 1430 39280 1450
rect 39360 1430 39400 1450
rect 39240 1400 39400 1430
rect 39480 1430 39520 1450
rect 39600 1430 39640 1450
rect 39720 1430 39760 1450
rect 39840 1430 39880 1450
rect 39480 1400 39880 1430
rect 39960 1430 40000 1450
rect 40080 1430 40120 1450
rect 39960 1400 40120 1430
rect 40200 1430 40240 1450
rect 40320 1430 40360 1450
rect 40440 1430 40480 1450
rect 40560 1430 40600 1450
rect 40200 1400 40600 1430
rect 40680 1420 40720 1450
rect 40800 1430 40840 1450
rect 40660 1400 40740 1420
rect 40800 1400 40910 1430
rect 38450 1360 38460 1400
rect 38500 1360 38510 1400
rect 38450 1340 38510 1360
rect 38630 1360 38640 1400
rect 38680 1360 38690 1400
rect 38630 1340 38690 1360
rect 39040 1360 39060 1400
rect 39100 1360 39120 1400
rect 39040 1340 39120 1360
rect 39280 1360 39300 1400
rect 39340 1360 39360 1400
rect 39280 1340 39360 1360
rect 39760 1360 39780 1400
rect 39820 1360 39840 1400
rect 39760 1340 39840 1360
rect 40000 1360 40020 1400
rect 40060 1360 40080 1400
rect 40000 1340 40080 1360
rect 40480 1360 40500 1400
rect 40540 1360 40560 1400
rect 40480 1340 40560 1360
rect 40660 1360 40680 1400
rect 40720 1360 40740 1400
rect 40660 1340 40740 1360
rect 40850 1360 40860 1400
rect 40900 1360 40910 1400
rect 40850 1340 40910 1360
rect 36380 1080 36460 1100
rect 36380 1040 36400 1080
rect 36440 1040 36460 1080
rect 36380 1010 36460 1040
rect 36380 980 37460 1010
rect 36340 900 36380 930
rect 36460 900 36500 980
rect 36580 900 36620 980
rect 36700 900 36740 930
rect 36820 900 36860 930
rect 36940 900 36980 980
rect 37060 900 37100 980
rect 37180 900 37220 930
rect 37300 900 37340 930
rect 37420 900 37460 980
rect 36340 770 36380 800
rect 36460 770 36500 800
rect 36580 770 36620 800
rect 36260 750 36380 770
rect 36260 710 36280 750
rect 36320 720 36380 750
rect 36700 720 36740 800
rect 36820 720 36860 800
rect 36940 770 36980 800
rect 37060 770 37100 800
rect 37180 720 37220 800
rect 37300 720 37340 800
rect 37420 770 37460 800
rect 36320 710 37340 720
rect 36260 690 37340 710
rect 39860 1080 39940 1100
rect 39860 1040 39880 1080
rect 39920 1040 39940 1080
rect 39860 1010 39940 1040
rect 38860 980 39940 1010
rect 38860 900 38900 980
rect 38980 900 39020 930
rect 39100 900 39140 930
rect 39220 900 39260 980
rect 39340 900 39380 980
rect 39460 900 39500 930
rect 39580 900 39620 930
rect 39700 900 39740 980
rect 39820 900 39860 980
rect 39940 900 39980 930
rect 38860 770 38900 800
rect 38980 720 39020 800
rect 39100 720 39140 800
rect 39220 770 39260 800
rect 39340 770 39380 800
rect 39460 720 39500 800
rect 39580 720 39620 800
rect 39700 770 39740 800
rect 39820 770 39860 800
rect 39940 770 39980 800
rect 39940 750 40060 770
rect 39940 720 40000 750
rect 38980 710 40000 720
rect 40040 710 40060 750
rect 38980 690 40060 710
rect 35960 430 36040 450
rect 35960 390 35980 430
rect 36020 390 36040 430
rect 35960 380 36040 390
rect 36200 430 36280 450
rect 36200 390 36220 430
rect 36260 390 36280 430
rect 36200 380 36280 390
rect 36440 430 36520 450
rect 36440 390 36460 430
rect 36500 390 36520 430
rect 36440 380 36520 390
rect 36680 430 36760 450
rect 36680 390 36700 430
rect 36740 390 36760 430
rect 36680 380 36760 390
rect 37160 430 37240 450
rect 37160 390 37180 430
rect 37220 390 37240 430
rect 37160 380 37240 390
rect 37400 430 37480 450
rect 37400 390 37420 430
rect 37460 390 37480 430
rect 37400 380 37480 390
rect 37640 430 37720 450
rect 37640 390 37660 430
rect 37700 390 37720 430
rect 37640 380 37720 390
rect 35860 350 36860 380
rect 36940 350 37940 380
rect 35860 -180 36860 -150
rect 36940 -180 37940 -150
rect 38600 430 38680 450
rect 38600 390 38620 430
rect 38660 390 38680 430
rect 38600 380 38680 390
rect 38840 430 38920 450
rect 38840 390 38860 430
rect 38900 390 38920 430
rect 38840 380 38920 390
rect 39080 430 39160 450
rect 39080 390 39100 430
rect 39140 390 39160 430
rect 39080 380 39160 390
rect 39560 430 39640 450
rect 39560 390 39580 430
rect 39620 390 39640 430
rect 39560 380 39640 390
rect 39800 430 39880 450
rect 39800 390 39820 430
rect 39860 390 39880 430
rect 39800 380 39880 390
rect 40040 430 40120 450
rect 40040 390 40060 430
rect 40100 390 40120 430
rect 40040 380 40120 390
rect 40280 430 40360 450
rect 40280 390 40300 430
rect 40340 390 40360 430
rect 40280 380 40360 390
rect 38380 350 39380 380
rect 39460 350 40460 380
rect 38380 -180 39380 -150
rect 39460 -180 40460 -150
rect 36200 -500 36280 -480
rect 36200 -540 36220 -500
rect 36260 -540 36280 -500
rect 36200 -560 36280 -540
rect 36360 -500 36440 -480
rect 36360 -540 36380 -500
rect 36420 -540 36440 -500
rect 36360 -560 36440 -540
rect 36520 -500 36600 -480
rect 36520 -540 36540 -500
rect 36580 -540 36600 -500
rect 36520 -560 36600 -540
rect 36680 -500 36760 -480
rect 36680 -540 36700 -500
rect 36740 -540 36760 -500
rect 36680 -560 36760 -540
rect 36840 -500 36920 -480
rect 36840 -540 36860 -500
rect 36900 -540 36920 -500
rect 36840 -560 36920 -540
rect 37000 -500 37080 -480
rect 37000 -540 37020 -500
rect 37060 -540 37080 -500
rect 37000 -560 37080 -540
rect 37160 -500 37240 -480
rect 37160 -540 37180 -500
rect 37220 -540 37240 -500
rect 37160 -560 37240 -540
rect 37320 -500 37400 -480
rect 37320 -540 37340 -500
rect 37380 -540 37400 -500
rect 37320 -560 37400 -540
rect 37480 -500 37560 -480
rect 37480 -540 37500 -500
rect 37540 -540 37560 -500
rect 37480 -560 37560 -540
rect 37640 -500 37720 -480
rect 37640 -540 37660 -500
rect 37700 -540 37720 -500
rect 37640 -560 37720 -540
rect 37800 -500 37880 -480
rect 37800 -540 37820 -500
rect 37860 -540 37880 -500
rect 37800 -560 37880 -540
rect 37960 -500 38040 -480
rect 37960 -540 37980 -500
rect 38020 -540 38040 -500
rect 37960 -560 38040 -540
rect 38280 -500 38360 -480
rect 38280 -540 38300 -500
rect 38340 -540 38360 -500
rect 38280 -560 38360 -540
rect 38440 -500 38520 -480
rect 38440 -540 38460 -500
rect 38500 -540 38520 -500
rect 38440 -560 38520 -540
rect 38600 -500 38680 -480
rect 38600 -540 38620 -500
rect 38660 -540 38680 -500
rect 38600 -560 38680 -540
rect 38760 -500 38840 -480
rect 38760 -540 38780 -500
rect 38820 -540 38840 -500
rect 38760 -560 38840 -540
rect 38920 -500 39000 -480
rect 38920 -540 38940 -500
rect 38980 -540 39000 -500
rect 38920 -560 39000 -540
rect 39080 -500 39160 -480
rect 39080 -540 39100 -500
rect 39140 -540 39160 -500
rect 39080 -560 39160 -540
rect 39240 -500 39320 -480
rect 39240 -540 39260 -500
rect 39300 -540 39320 -500
rect 39240 -560 39320 -540
rect 39400 -500 39480 -480
rect 39400 -540 39420 -500
rect 39460 -540 39480 -500
rect 39400 -560 39480 -540
rect 39560 -500 39640 -480
rect 39560 -540 39580 -500
rect 39620 -540 39640 -500
rect 39560 -560 39640 -540
rect 39720 -500 39800 -480
rect 39720 -540 39740 -500
rect 39780 -540 39800 -500
rect 39720 -560 39800 -540
rect 39880 -500 39960 -480
rect 39880 -540 39900 -500
rect 39940 -540 39960 -500
rect 39880 -560 39960 -540
rect 40040 -500 40120 -480
rect 40040 -540 40060 -500
rect 40100 -540 40120 -500
rect 40040 -560 40120 -540
rect 36120 -590 38120 -560
rect 38200 -590 40200 -560
rect 36120 -820 38120 -790
rect 38200 -820 40200 -790
rect 36900 -1050 36960 -1030
rect 36900 -1090 36910 -1050
rect 36950 -1090 36960 -1050
rect 36420 -1140 36450 -1110
rect 36530 -1120 37110 -1090
rect 36530 -1140 36560 -1120
rect 36640 -1140 36670 -1120
rect 36750 -1140 36780 -1120
rect 36860 -1140 36890 -1120
rect 36970 -1140 37000 -1120
rect 37080 -1140 37110 -1120
rect 37190 -1140 37220 -1110
rect 36420 -1360 36450 -1340
rect 36350 -1390 36450 -1360
rect 36530 -1370 36560 -1340
rect 36640 -1370 36670 -1340
rect 36750 -1370 36780 -1340
rect 36860 -1370 36890 -1340
rect 36970 -1370 37000 -1340
rect 37080 -1370 37110 -1340
rect 37190 -1360 37220 -1340
rect 37190 -1390 37290 -1360
rect 36350 -1430 36360 -1390
rect 36400 -1430 36410 -1390
rect 36350 -1450 36410 -1430
rect 37230 -1430 37240 -1390
rect 37280 -1430 37290 -1390
rect 37230 -1450 37290 -1430
rect 38130 -1050 38190 -1030
rect 38130 -1090 38140 -1050
rect 38180 -1090 38190 -1050
rect 37650 -1140 37680 -1110
rect 37760 -1120 38560 -1090
rect 37760 -1140 37790 -1120
rect 37870 -1140 37900 -1120
rect 37980 -1140 38010 -1120
rect 38090 -1140 38120 -1120
rect 38200 -1140 38230 -1120
rect 38310 -1140 38340 -1120
rect 38420 -1140 38450 -1120
rect 38530 -1140 38560 -1120
rect 38640 -1140 38670 -1110
rect 37650 -1360 37680 -1340
rect 37580 -1390 37680 -1360
rect 37760 -1370 37790 -1340
rect 37870 -1370 37900 -1340
rect 37980 -1370 38010 -1340
rect 38090 -1370 38120 -1340
rect 38200 -1370 38230 -1340
rect 38310 -1370 38340 -1340
rect 38420 -1370 38450 -1340
rect 38530 -1370 38560 -1340
rect 38640 -1360 38670 -1340
rect 37730 -1390 37810 -1370
rect 38640 -1390 38740 -1360
rect 37580 -1430 37590 -1390
rect 37630 -1430 37640 -1390
rect 37580 -1450 37640 -1430
rect 37730 -1430 37750 -1390
rect 37790 -1430 37810 -1390
rect 37730 -1450 37810 -1430
rect 38680 -1430 38690 -1390
rect 38730 -1430 38740 -1390
rect 38680 -1450 38740 -1430
rect 39360 -1050 39420 -1030
rect 39360 -1090 39370 -1050
rect 39410 -1090 39420 -1050
rect 39100 -1140 39130 -1110
rect 39210 -1120 39790 -1090
rect 39210 -1140 39240 -1120
rect 39320 -1140 39350 -1120
rect 39430 -1140 39460 -1120
rect 39540 -1140 39570 -1120
rect 39650 -1140 39680 -1120
rect 39760 -1140 39790 -1120
rect 39870 -1140 39900 -1110
rect 39100 -1360 39130 -1340
rect 39030 -1390 39130 -1360
rect 39210 -1370 39240 -1340
rect 39320 -1370 39350 -1340
rect 39430 -1370 39460 -1340
rect 39540 -1370 39570 -1340
rect 39650 -1370 39680 -1340
rect 39760 -1370 39790 -1340
rect 39870 -1360 39900 -1340
rect 39870 -1390 39970 -1360
rect 39030 -1430 39040 -1390
rect 39080 -1430 39090 -1390
rect 39030 -1450 39090 -1430
rect 39910 -1430 39920 -1390
rect 39960 -1430 39970 -1390
rect 39910 -1450 39970 -1430
<< polycont >>
rect 6090 7010 6130 7050
rect 6420 7010 6460 7050
rect 6750 7010 6790 7050
rect 7370 7010 7410 7050
rect 8140 7010 8180 7050
rect 8690 7010 8730 7050
rect 9530 7010 9570 7050
rect 9860 7010 9900 7050
rect 10190 7010 10230 7050
rect 5450 5880 5490 5920
rect 5890 5880 5930 5920
rect 5670 5540 5710 5580
rect 6520 6080 6560 6120
rect 9760 6080 9800 6120
rect 7960 5340 8000 5380
rect 9400 5340 9440 5380
rect 10380 5880 10420 5920
rect 10820 5880 10860 5920
rect 10600 5540 10640 5580
rect 5420 4360 5460 4400
rect 5600 4360 5640 4400
rect 5780 4360 5820 4400
rect 6260 4360 6300 4400
rect 6500 4360 6540 4400
rect 6980 4360 7020 4400
rect 7220 4360 7260 4400
rect 7640 4360 7680 4400
rect 7820 4360 7860 4400
rect 8460 4360 8500 4400
rect 8640 4360 8680 4400
rect 9060 4360 9100 4400
rect 9300 4360 9340 4400
rect 9780 4360 9820 4400
rect 10020 4360 10060 4400
rect 10500 4360 10540 4400
rect 10680 4360 10720 4400
rect 10860 4360 10900 4400
rect 6400 4040 6440 4080
rect 6280 3710 6320 3750
rect 9880 4040 9920 4080
rect 10000 3710 10040 3750
rect 36090 4010 36130 4050
rect 36420 4010 36460 4050
rect 36750 4010 36790 4050
rect 37370 4010 37410 4050
rect 38140 4010 38180 4050
rect 38690 4010 38730 4050
rect 39530 4010 39570 4050
rect 39860 4010 39900 4050
rect 40190 4010 40230 4050
rect 5980 3390 6020 3430
rect 6220 3390 6260 3430
rect 6460 3390 6500 3430
rect 6700 3390 6740 3430
rect 7180 3390 7220 3430
rect 7420 3390 7460 3430
rect 7660 3390 7700 3430
rect 8620 3390 8660 3430
rect 8860 3390 8900 3430
rect 9100 3390 9140 3430
rect 9580 3390 9620 3430
rect 9820 3390 9860 3430
rect 10060 3390 10100 3430
rect 10300 3390 10340 3430
rect 35450 2880 35490 2920
rect 35890 2880 35930 2920
rect 6220 2460 6260 2500
rect 6380 2460 6420 2500
rect 6540 2460 6580 2500
rect 6700 2460 6740 2500
rect 6860 2460 6900 2500
rect 7020 2460 7060 2500
rect 7180 2460 7220 2500
rect 7340 2460 7380 2500
rect 7500 2460 7540 2500
rect 7660 2460 7700 2500
rect 7820 2460 7860 2500
rect 7980 2460 8020 2500
rect 8300 2460 8340 2500
rect 8460 2460 8500 2500
rect 8620 2460 8660 2500
rect 8780 2460 8820 2500
rect 8940 2460 8980 2500
rect 9100 2460 9140 2500
rect 9260 2460 9300 2500
rect 9420 2460 9460 2500
rect 9580 2460 9620 2500
rect 9740 2460 9780 2500
rect 9900 2460 9940 2500
rect 10060 2460 10100 2500
rect 35670 2540 35710 2580
rect 36520 3080 36560 3120
rect 39760 3080 39800 3120
rect 37960 2340 38000 2380
rect 39400 2340 39440 2380
rect 40380 2880 40420 2920
rect 40820 2880 40860 2920
rect 40600 2540 40640 2580
rect 6910 1910 6950 1950
rect 6360 1570 6400 1610
rect 7240 1570 7280 1610
rect 8140 1910 8180 1950
rect 7590 1570 7630 1610
rect 7750 1570 7790 1610
rect 8690 1570 8730 1610
rect 9370 1910 9410 1950
rect 9040 1570 9080 1610
rect 9920 1570 9960 1610
rect 35420 1360 35460 1400
rect 35600 1360 35640 1400
rect 35780 1360 35820 1400
rect 36260 1360 36300 1400
rect 36500 1360 36540 1400
rect 36980 1360 37020 1400
rect 37220 1360 37260 1400
rect 37640 1360 37680 1400
rect 37820 1360 37860 1400
rect 38460 1360 38500 1400
rect 38640 1360 38680 1400
rect 39060 1360 39100 1400
rect 39300 1360 39340 1400
rect 39780 1360 39820 1400
rect 40020 1360 40060 1400
rect 40500 1360 40540 1400
rect 40680 1360 40720 1400
rect 40860 1360 40900 1400
rect 36400 1040 36440 1080
rect 36280 710 36320 750
rect 39880 1040 39920 1080
rect 40000 710 40040 750
rect 35980 390 36020 430
rect 36220 390 36260 430
rect 36460 390 36500 430
rect 36700 390 36740 430
rect 37180 390 37220 430
rect 37420 390 37460 430
rect 37660 390 37700 430
rect 38620 390 38660 430
rect 38860 390 38900 430
rect 39100 390 39140 430
rect 39580 390 39620 430
rect 39820 390 39860 430
rect 40060 390 40100 430
rect 40300 390 40340 430
rect 36220 -540 36260 -500
rect 36380 -540 36420 -500
rect 36540 -540 36580 -500
rect 36700 -540 36740 -500
rect 36860 -540 36900 -500
rect 37020 -540 37060 -500
rect 37180 -540 37220 -500
rect 37340 -540 37380 -500
rect 37500 -540 37540 -500
rect 37660 -540 37700 -500
rect 37820 -540 37860 -500
rect 37980 -540 38020 -500
rect 38300 -540 38340 -500
rect 38460 -540 38500 -500
rect 38620 -540 38660 -500
rect 38780 -540 38820 -500
rect 38940 -540 38980 -500
rect 39100 -540 39140 -500
rect 39260 -540 39300 -500
rect 39420 -540 39460 -500
rect 39580 -540 39620 -500
rect 39740 -540 39780 -500
rect 39900 -540 39940 -500
rect 40060 -540 40100 -500
rect 36910 -1090 36950 -1050
rect 36360 -1430 36400 -1390
rect 37240 -1430 37280 -1390
rect 38140 -1090 38180 -1050
rect 37590 -1430 37630 -1390
rect 37750 -1430 37790 -1390
rect 38690 -1430 38730 -1390
rect 39370 -1090 39410 -1050
rect 39040 -1430 39080 -1390
rect 39920 -1430 39960 -1390
<< xpolycontact >>
rect 222 7110 662 7180
rect 1890 7110 2330 7180
rect 222 6990 662 7060
rect 1890 6990 2330 7060
rect 222 6580 662 6650
rect 1830 6580 2270 6650
rect 222 6460 662 6530
rect 1830 6460 2270 6530
rect 2792 6840 3232 6910
rect 4400 6840 4840 6910
rect 2792 6720 3232 6790
rect 4400 6720 4840 6790
rect 2792 6600 3232 6670
rect 4400 6600 4840 6670
rect 612 6050 1050 6120
rect 1428 6050 1868 6120
rect 2792 6480 3232 6550
rect 4400 6480 4840 6550
rect 2792 6360 3232 6430
rect 4400 6360 4840 6430
rect 2792 6240 3232 6310
rect 4400 6240 4840 6310
rect 612 5630 1050 5700
rect 1428 5630 1868 5700
rect 3122 5830 3562 5900
rect 3990 5830 4430 5900
rect 44222 -2890 44662 -2820
rect 45890 -2890 46330 -2820
rect 44222 -3010 44662 -2940
rect 45890 -3010 46330 -2940
rect 44222 -3420 44662 -3350
rect 45830 -3420 46270 -3350
rect 44222 -3540 44662 -3470
rect 45830 -3540 46270 -3470
rect 46792 -3160 47232 -3090
rect 48400 -3160 48840 -3090
rect 46792 -3280 47232 -3210
rect 48400 -3280 48840 -3210
rect 46792 -3400 47232 -3330
rect 48400 -3400 48840 -3330
rect 44612 -3950 45050 -3880
rect 45428 -3950 45868 -3880
rect 46792 -3520 47232 -3450
rect 48400 -3520 48840 -3450
rect 46792 -3640 47232 -3570
rect 48400 -3640 48840 -3570
rect 46792 -3760 47232 -3690
rect 48400 -3760 48840 -3690
rect 44612 -4370 45050 -4300
rect 45428 -4370 45868 -4300
rect 47122 -4170 47562 -4100
rect 47990 -4170 48430 -4100
<< ppolyres >>
rect 1050 6050 1428 6120
rect 1050 5630 1428 5700
rect 45050 -3950 45428 -3880
rect 45050 -4370 45428 -4300
<< xpolyres >>
rect 662 7110 1890 7180
rect 662 6990 1890 7060
rect 662 6580 1830 6650
rect 662 6460 1830 6530
rect 3232 6840 4400 6910
rect 3232 6720 4400 6790
rect 3232 6600 4400 6670
rect 3232 6480 4400 6550
rect 3232 6360 4400 6430
rect 3232 6240 4400 6310
rect 3562 5830 3990 5900
rect 44662 -2890 45890 -2820
rect 44662 -3010 45890 -2940
rect 44662 -3420 45830 -3350
rect 44662 -3540 45830 -3470
rect 47232 -3160 48400 -3090
rect 47232 -3280 48400 -3210
rect 47232 -3400 48400 -3330
rect 47232 -3520 48400 -3450
rect 47232 -3640 48400 -3570
rect 47232 -3760 48400 -3690
rect 47562 -4170 47990 -4100
<< locali >>
rect 50 7280 1180 7320
rect 1340 7280 2470 7320
rect 50 7160 90 7280
rect 132 7170 222 7180
rect 132 7120 152 7170
rect 202 7120 222 7170
rect 132 7110 222 7120
rect 2260 7060 2330 7110
rect 50 6890 90 7000
rect 132 7050 222 7060
rect 132 7000 152 7050
rect 202 7000 222 7050
rect 132 6990 222 7000
rect 2430 7160 2470 7280
rect 5970 7110 6360 7150
rect 6520 7110 6910 7150
rect 2430 6890 2470 7000
rect 50 6850 1180 6890
rect 1340 6850 2470 6890
rect 2620 7010 3690 7050
rect 3850 7010 5010 7050
rect 1230 6790 1270 6850
rect 50 6750 1150 6790
rect 1310 6750 2410 6790
rect 50 6630 90 6750
rect 132 6640 222 6650
rect 132 6590 152 6640
rect 202 6590 222 6640
rect 132 6580 222 6590
rect 2200 6530 2270 6580
rect 50 6360 90 6470
rect 132 6520 222 6530
rect 132 6470 152 6520
rect 202 6470 222 6520
rect 132 6460 222 6470
rect 2370 6630 2410 6750
rect 2620 6650 2660 7010
rect 2702 6900 2792 6910
rect 2702 6850 2722 6900
rect 2772 6850 2792 6900
rect 2702 6840 2792 6850
rect 4840 6840 4920 6910
rect 2702 6780 2792 6790
rect 2702 6730 2722 6780
rect 2772 6730 2792 6780
rect 2702 6720 2792 6730
rect 4770 6670 4840 6720
rect 2410 6570 2450 6590
rect 2430 6530 2450 6570
rect 2410 6510 2450 6530
rect 2580 6570 2620 6590
rect 2580 6530 2600 6570
rect 2580 6510 2620 6530
rect 1190 6380 1270 6400
rect 1190 6360 1210 6380
rect 1250 6360 1270 6380
rect 2370 6360 2410 6470
rect 50 6320 1150 6360
rect 1310 6320 2410 6360
rect 1210 6260 1250 6320
rect 440 6220 1150 6260
rect 1310 6220 2040 6260
rect 440 6160 480 6220
rect 2000 6160 2040 6220
rect 522 6110 612 6120
rect 522 6060 542 6110
rect 592 6060 612 6110
rect 522 6050 612 6060
rect 1868 6110 1958 6120
rect 1868 6060 1888 6110
rect 1938 6060 1958 6110
rect 1868 6050 1958 6060
rect 440 5940 480 6000
rect 2620 6140 2660 6490
rect 2712 6600 2792 6670
rect 2712 6310 2752 6600
rect 4880 6550 4920 6840
rect 4840 6480 4920 6550
rect 4970 6650 5010 7010
rect 5970 6940 6010 7110
rect 6090 7070 6130 7110
rect 6750 7070 6790 7110
rect 6070 7050 6150 7070
rect 6070 7010 6090 7050
rect 6130 7010 6150 7050
rect 6070 6990 6150 7010
rect 6290 7050 6370 7070
rect 6290 7010 6310 7050
rect 6350 7010 6370 7050
rect 6290 6990 6370 7010
rect 6410 7050 6470 7070
rect 6410 7010 6420 7050
rect 6460 7010 6470 7050
rect 6410 6990 6470 7010
rect 6510 7050 6590 7070
rect 6510 7010 6530 7050
rect 6570 7010 6590 7050
rect 6510 6990 6590 7010
rect 6630 7050 6690 7070
rect 6630 7010 6640 7050
rect 6680 7010 6690 7050
rect 6630 6990 6690 7010
rect 6730 7050 6810 7070
rect 6730 7010 6750 7050
rect 6790 7010 6810 7050
rect 6730 6990 6810 7010
rect 6090 6950 6130 6990
rect 6310 6950 6350 6990
rect 6530 6950 6570 6990
rect 6640 6950 6680 6990
rect 6750 6950 6790 6990
rect 5970 6610 6010 6780
rect 6080 6930 6140 6950
rect 6080 6786 6090 6930
rect 6130 6786 6140 6930
rect 6080 6770 6140 6786
rect 6190 6930 6250 6950
rect 6190 6786 6200 6930
rect 6240 6786 6250 6930
rect 6190 6770 6250 6786
rect 6300 6930 6360 6950
rect 6300 6786 6310 6930
rect 6350 6786 6360 6930
rect 6300 6770 6360 6786
rect 6410 6930 6470 6950
rect 6410 6786 6420 6930
rect 6460 6786 6470 6930
rect 6410 6770 6470 6786
rect 6520 6930 6580 6950
rect 6520 6786 6530 6930
rect 6570 6786 6580 6930
rect 6520 6770 6580 6786
rect 6630 6930 6690 6950
rect 6630 6786 6640 6930
rect 6680 6786 6690 6930
rect 6630 6770 6690 6786
rect 6740 6930 6800 6950
rect 6740 6786 6750 6930
rect 6790 6786 6800 6930
rect 6740 6770 6800 6786
rect 6870 6940 6910 7110
rect 6200 6730 6240 6770
rect 6420 6730 6460 6770
rect 6640 6730 6680 6770
rect 6180 6710 6260 6730
rect 6180 6670 6200 6710
rect 6240 6670 6260 6710
rect 6180 6650 6260 6670
rect 6400 6710 6480 6730
rect 6400 6670 6420 6710
rect 6460 6670 6480 6710
rect 6400 6650 6480 6670
rect 6620 6710 6700 6730
rect 6620 6670 6640 6710
rect 6680 6670 6700 6710
rect 6620 6650 6700 6670
rect 6870 6610 6910 6780
rect 5970 6570 6360 6610
rect 6520 6570 6910 6610
rect 7250 7110 8080 7150
rect 8240 7110 9070 7150
rect 7250 6940 7290 7110
rect 7370 7070 7410 7110
rect 8690 7070 8730 7110
rect 7350 7050 7430 7070
rect 7350 7010 7370 7050
rect 7410 7010 7430 7050
rect 7350 6990 7430 7010
rect 7570 7050 7650 7070
rect 7570 7010 7590 7050
rect 7630 7010 7650 7050
rect 7570 6990 7650 7010
rect 7790 7050 7870 7070
rect 7790 7010 7810 7050
rect 7850 7010 7870 7050
rect 7790 6990 7870 7010
rect 8010 7050 8090 7070
rect 8010 7010 8030 7050
rect 8070 7010 8090 7050
rect 8010 6990 8090 7010
rect 8130 7050 8190 7070
rect 8130 7010 8140 7050
rect 8180 7010 8190 7050
rect 8130 6990 8190 7010
rect 8230 7050 8310 7070
rect 8230 7010 8250 7050
rect 8290 7010 8310 7050
rect 8230 6990 8310 7010
rect 8450 7050 8530 7070
rect 8450 7010 8470 7050
rect 8510 7010 8530 7050
rect 8450 6990 8530 7010
rect 8570 7050 8630 7070
rect 8570 7010 8580 7050
rect 8620 7010 8630 7050
rect 8570 6990 8630 7010
rect 8670 7050 8750 7070
rect 8670 7010 8690 7050
rect 8730 7010 8750 7050
rect 8670 6990 8750 7010
rect 7370 6950 7410 6990
rect 7590 6950 7630 6990
rect 7810 6950 7850 6990
rect 8030 6950 8070 6990
rect 8250 6950 8290 6990
rect 8470 6950 8510 6990
rect 8580 6950 8620 6990
rect 8690 6950 8730 6990
rect 7250 6610 7290 6780
rect 7360 6930 7420 6950
rect 7360 6890 7370 6930
rect 7410 6890 7420 6930
rect 7360 6830 7420 6890
rect 7360 6790 7370 6830
rect 7410 6790 7420 6830
rect 7360 6770 7420 6790
rect 7470 6930 7530 6950
rect 7470 6890 7480 6930
rect 7520 6890 7530 6930
rect 7470 6830 7530 6890
rect 7470 6790 7480 6830
rect 7520 6790 7530 6830
rect 7470 6770 7530 6790
rect 7580 6930 7640 6950
rect 7580 6890 7590 6930
rect 7630 6890 7640 6930
rect 7580 6830 7640 6890
rect 7580 6790 7590 6830
rect 7630 6790 7640 6830
rect 7580 6770 7640 6790
rect 7690 6930 7750 6950
rect 7690 6890 7700 6930
rect 7740 6890 7750 6930
rect 7690 6830 7750 6890
rect 7690 6790 7700 6830
rect 7740 6790 7750 6830
rect 7690 6770 7750 6790
rect 7800 6930 7860 6950
rect 7800 6890 7810 6930
rect 7850 6890 7860 6930
rect 7800 6830 7860 6890
rect 7800 6790 7810 6830
rect 7850 6790 7860 6830
rect 7800 6770 7860 6790
rect 7910 6930 7970 6950
rect 7910 6890 7920 6930
rect 7960 6890 7970 6930
rect 7910 6830 7970 6890
rect 7910 6790 7920 6830
rect 7960 6790 7970 6830
rect 7910 6770 7970 6790
rect 8020 6930 8080 6950
rect 8020 6890 8030 6930
rect 8070 6890 8080 6930
rect 8020 6830 8080 6890
rect 8020 6790 8030 6830
rect 8070 6790 8080 6830
rect 8020 6770 8080 6790
rect 8130 6930 8190 6950
rect 8130 6890 8140 6930
rect 8180 6890 8190 6930
rect 8130 6830 8190 6890
rect 8130 6790 8140 6830
rect 8180 6790 8190 6830
rect 8130 6770 8190 6790
rect 8240 6930 8300 6950
rect 8240 6890 8250 6930
rect 8290 6890 8300 6930
rect 8240 6830 8300 6890
rect 8240 6790 8250 6830
rect 8290 6790 8300 6830
rect 8240 6770 8300 6790
rect 8350 6930 8410 6950
rect 8350 6890 8360 6930
rect 8400 6890 8410 6930
rect 8350 6830 8410 6890
rect 8350 6790 8360 6830
rect 8400 6790 8410 6830
rect 8350 6770 8410 6790
rect 8460 6930 8520 6950
rect 8460 6890 8470 6930
rect 8510 6890 8520 6930
rect 8460 6830 8520 6890
rect 8460 6790 8470 6830
rect 8510 6790 8520 6830
rect 8460 6770 8520 6790
rect 8570 6930 8630 6950
rect 8570 6890 8580 6930
rect 8620 6890 8630 6930
rect 8570 6830 8630 6890
rect 8570 6790 8580 6830
rect 8620 6790 8630 6830
rect 8570 6770 8630 6790
rect 8680 6930 8740 6950
rect 8680 6890 8690 6930
rect 8730 6890 8740 6930
rect 8680 6830 8740 6890
rect 8680 6790 8690 6830
rect 8730 6790 8740 6830
rect 8680 6770 8740 6790
rect 9030 6940 9070 7110
rect 7480 6730 7520 6770
rect 7700 6730 7740 6770
rect 7920 6730 7960 6770
rect 8140 6730 8180 6770
rect 8360 6730 8400 6770
rect 8580 6730 8620 6770
rect 7460 6710 7540 6730
rect 7460 6670 7480 6710
rect 7520 6670 7540 6710
rect 7460 6650 7540 6670
rect 7680 6710 7760 6730
rect 7680 6670 7700 6710
rect 7740 6670 7760 6710
rect 7680 6650 7760 6670
rect 7900 6710 7980 6730
rect 7900 6670 7920 6710
rect 7960 6670 7980 6710
rect 7900 6650 7980 6670
rect 8120 6710 8200 6730
rect 8120 6670 8140 6710
rect 8180 6670 8200 6710
rect 8120 6650 8200 6670
rect 8340 6710 8420 6730
rect 8340 6670 8360 6710
rect 8400 6670 8420 6710
rect 8340 6650 8420 6670
rect 8560 6710 8640 6730
rect 8560 6670 8580 6710
rect 8620 6670 8640 6710
rect 8560 6650 8640 6670
rect 9030 6610 9070 6780
rect 7250 6570 8080 6610
rect 8240 6570 9070 6610
rect 9410 7110 9800 7150
rect 9960 7110 10350 7150
rect 9410 6940 9450 7110
rect 9530 7070 9570 7110
rect 10190 7070 10230 7110
rect 9510 7050 9590 7070
rect 9510 7010 9530 7050
rect 9570 7010 9590 7050
rect 9510 6990 9590 7010
rect 9730 7050 9810 7070
rect 9730 7010 9750 7050
rect 9790 7010 9810 7050
rect 9730 6990 9810 7010
rect 9850 7050 9910 7070
rect 9850 7010 9860 7050
rect 9900 7010 9910 7050
rect 9850 6990 9910 7010
rect 9950 7050 10030 7070
rect 9950 7010 9970 7050
rect 10010 7010 10030 7050
rect 9950 6990 10030 7010
rect 10170 7050 10250 7070
rect 10170 7010 10190 7050
rect 10230 7010 10250 7050
rect 10170 6990 10250 7010
rect 9530 6950 9570 6990
rect 9750 6950 9790 6990
rect 9970 6950 10010 6990
rect 10190 6950 10230 6990
rect 9410 6610 9450 6780
rect 9520 6930 9580 6950
rect 9520 6790 9530 6930
rect 9570 6790 9580 6930
rect 9520 6770 9580 6790
rect 9630 6930 9690 6950
rect 9630 6790 9640 6930
rect 9680 6790 9690 6930
rect 9630 6770 9690 6790
rect 9740 6930 9800 6950
rect 9740 6790 9750 6930
rect 9790 6790 9800 6930
rect 9740 6770 9800 6790
rect 9850 6930 9910 6950
rect 9850 6790 9860 6930
rect 9900 6790 9910 6930
rect 9850 6770 9910 6790
rect 9960 6930 10020 6950
rect 9960 6790 9970 6930
rect 10010 6790 10020 6930
rect 9960 6770 10020 6790
rect 10070 6930 10130 6950
rect 10070 6790 10080 6930
rect 10120 6790 10130 6930
rect 10070 6770 10130 6790
rect 10180 6930 10240 6950
rect 10180 6790 10190 6930
rect 10230 6790 10240 6930
rect 10180 6770 10240 6790
rect 10310 6940 10350 7110
rect 9640 6730 9680 6770
rect 9860 6730 9900 6770
rect 10080 6730 10120 6770
rect 9620 6710 9700 6730
rect 9620 6670 9640 6710
rect 9680 6670 9700 6710
rect 9620 6650 9700 6670
rect 9840 6710 9920 6730
rect 9840 6670 9860 6710
rect 9900 6670 9920 6710
rect 9840 6650 9920 6670
rect 10060 6710 10140 6730
rect 10060 6670 10080 6710
rect 10120 6670 10140 6710
rect 10060 6650 10140 6670
rect 10310 6610 10350 6780
rect 9410 6570 9800 6610
rect 9930 6570 10350 6610
rect 2792 6430 2862 6480
rect 4840 6420 4930 6430
rect 4840 6370 4860 6420
rect 4910 6370 4930 6420
rect 4840 6360 4930 6370
rect 2712 6240 2792 6310
rect 4840 6300 4930 6320
rect 4840 6250 4860 6300
rect 4910 6250 4930 6300
rect 4840 6230 4930 6250
rect 4970 6140 5010 6490
rect 2620 6100 3690 6140
rect 3850 6100 5010 6140
rect 6400 6180 8080 6220
rect 8240 6180 9920 6220
rect 3750 6040 3790 6100
rect 5650 6040 5730 6060
rect 2000 5940 2040 6000
rect 440 5900 1150 5940
rect 1310 5900 2040 5940
rect 2950 6000 3690 6040
rect 3850 6000 4600 6040
rect 5650 6020 5670 6040
rect 5710 6020 5730 6040
rect 2950 5940 2990 6000
rect 1210 5840 1250 5900
rect 440 5800 1150 5840
rect 1310 5800 2040 5840
rect 440 5740 480 5800
rect 2000 5740 2040 5800
rect 522 5690 612 5700
rect 522 5640 542 5690
rect 592 5640 612 5690
rect 522 5630 612 5640
rect 1868 5690 1958 5700
rect 1868 5640 1888 5690
rect 1938 5640 1958 5690
rect 1868 5630 1958 5640
rect 440 5520 480 5580
rect 4560 5940 4600 6000
rect 3032 5890 3122 5900
rect 3032 5840 3052 5890
rect 3102 5840 3122 5890
rect 3032 5830 3122 5840
rect 4430 5890 4520 5900
rect 4430 5840 4450 5890
rect 4500 5840 4520 5890
rect 4430 5830 4520 5840
rect 2950 5730 2990 5780
rect 4560 5730 4600 5780
rect 2950 5690 3690 5730
rect 3850 5690 4600 5730
rect 5330 5980 5610 6020
rect 5770 5980 6050 6020
rect 5330 5810 5370 5980
rect 5450 5940 5490 5980
rect 5890 5940 5930 5980
rect 2000 5520 2040 5580
rect 440 5480 1150 5520
rect 1310 5480 2040 5520
rect 5330 5480 5370 5650
rect 5440 5920 5500 5940
rect 5440 5880 5450 5920
rect 5490 5880 5500 5920
rect 5440 5800 5500 5880
rect 5650 5920 5730 5940
rect 5650 5880 5670 5920
rect 5710 5880 5730 5920
rect 5650 5860 5730 5880
rect 5880 5920 5940 5940
rect 5880 5880 5890 5920
rect 5930 5880 5940 5920
rect 5670 5820 5710 5860
rect 5440 5760 5450 5800
rect 5490 5760 5500 5800
rect 5440 5700 5500 5760
rect 5440 5660 5450 5700
rect 5490 5660 5500 5700
rect 5440 5640 5500 5660
rect 5550 5800 5610 5820
rect 5550 5760 5560 5800
rect 5600 5760 5610 5800
rect 5550 5700 5610 5760
rect 5550 5660 5560 5700
rect 5600 5660 5610 5700
rect 5550 5640 5610 5660
rect 5660 5800 5720 5820
rect 5660 5760 5670 5800
rect 5710 5760 5720 5800
rect 5660 5700 5720 5760
rect 5660 5660 5670 5700
rect 5710 5660 5720 5700
rect 5660 5640 5720 5660
rect 5770 5800 5830 5820
rect 5770 5760 5780 5800
rect 5820 5760 5830 5800
rect 5770 5700 5830 5760
rect 5770 5660 5780 5700
rect 5820 5660 5830 5700
rect 5770 5640 5830 5660
rect 5880 5800 5940 5880
rect 5880 5760 5890 5800
rect 5930 5760 5940 5800
rect 5880 5700 5940 5760
rect 5880 5660 5890 5700
rect 5930 5660 5940 5700
rect 5880 5640 5940 5660
rect 6010 5810 6050 5980
rect 5560 5600 5600 5640
rect 5780 5600 5820 5640
rect 5520 5580 5600 5600
rect 5520 5540 5540 5580
rect 5580 5540 5600 5580
rect 5520 5520 5600 5540
rect 5650 5580 5730 5600
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 5780 5580 5860 5600
rect 5780 5540 5800 5580
rect 5840 5540 5860 5580
rect 5780 5520 5860 5540
rect 6010 5480 6050 5650
rect 5330 5440 5610 5480
rect 5770 5440 6050 5480
rect 6400 5810 6440 6180
rect 6520 6140 6560 6180
rect 9760 6140 9800 6180
rect 6500 6120 6580 6140
rect 6500 6080 6520 6120
rect 6560 6080 6580 6120
rect 6500 6060 6580 6080
rect 6860 6120 6940 6140
rect 6860 6080 6880 6120
rect 6920 6080 6940 6120
rect 6860 6060 6940 6080
rect 7220 6120 7300 6140
rect 7220 6080 7240 6120
rect 7280 6080 7300 6120
rect 7220 6060 7300 6080
rect 7580 6120 7660 6140
rect 7580 6080 7600 6120
rect 7640 6080 7660 6120
rect 7580 6060 7660 6080
rect 7940 6120 8020 6140
rect 7940 6080 7960 6120
rect 8000 6080 8020 6120
rect 7940 6060 8020 6080
rect 8300 6120 8380 6140
rect 8300 6080 8320 6120
rect 8360 6080 8380 6120
rect 8300 6060 8380 6080
rect 8660 6120 8740 6140
rect 8660 6080 8680 6120
rect 8720 6080 8740 6120
rect 8660 6060 8740 6080
rect 9020 6120 9100 6140
rect 9020 6080 9040 6120
rect 9080 6080 9100 6120
rect 9020 6060 9100 6080
rect 9380 6120 9460 6140
rect 9380 6080 9400 6120
rect 9440 6080 9460 6120
rect 9380 6060 9460 6080
rect 9740 6120 9820 6140
rect 9740 6080 9760 6120
rect 9800 6080 9820 6120
rect 9740 6060 9820 6080
rect 6520 6020 6560 6060
rect 6880 6020 6920 6060
rect 7240 6020 7280 6060
rect 7600 6020 7640 6060
rect 7960 6020 8000 6060
rect 8320 6020 8360 6060
rect 8680 6020 8720 6060
rect 9040 6020 9080 6060
rect 9400 6020 9440 6060
rect 9760 6020 9800 6060
rect 1300 4110 1550 5400
rect 2660 4110 2910 5400
rect 4020 4110 4270 5400
rect 6400 5270 6440 5650
rect 6510 6000 6570 6020
rect 6510 5960 6520 6000
rect 6560 5960 6570 6000
rect 6510 5900 6570 5960
rect 6510 5860 6520 5900
rect 6560 5860 6570 5900
rect 6510 5800 6570 5860
rect 6510 5760 6520 5800
rect 6560 5760 6570 5800
rect 6510 5700 6570 5760
rect 6510 5660 6520 5700
rect 6560 5660 6570 5700
rect 6510 5600 6570 5660
rect 6510 5560 6520 5600
rect 6560 5560 6570 5600
rect 6510 5500 6570 5560
rect 6510 5460 6520 5500
rect 6560 5460 6570 5500
rect 6510 5440 6570 5460
rect 6690 6000 6750 6020
rect 6690 5960 6700 6000
rect 6740 5960 6750 6000
rect 6690 5900 6750 5960
rect 6690 5860 6700 5900
rect 6740 5860 6750 5900
rect 6690 5800 6750 5860
rect 6690 5760 6700 5800
rect 6740 5760 6750 5800
rect 6690 5700 6750 5760
rect 6690 5660 6700 5700
rect 6740 5660 6750 5700
rect 6690 5600 6750 5660
rect 6690 5560 6700 5600
rect 6740 5560 6750 5600
rect 6690 5500 6750 5560
rect 6690 5460 6700 5500
rect 6740 5460 6750 5500
rect 6690 5440 6750 5460
rect 6870 6000 6930 6020
rect 6870 5960 6880 6000
rect 6920 5960 6930 6000
rect 6870 5900 6930 5960
rect 6870 5860 6880 5900
rect 6920 5860 6930 5900
rect 6870 5800 6930 5860
rect 6870 5760 6880 5800
rect 6920 5760 6930 5800
rect 6870 5700 6930 5760
rect 6870 5660 6880 5700
rect 6920 5660 6930 5700
rect 6870 5600 6930 5660
rect 6870 5560 6880 5600
rect 6920 5560 6930 5600
rect 6870 5500 6930 5560
rect 6870 5460 6880 5500
rect 6920 5460 6930 5500
rect 6870 5440 6930 5460
rect 7050 6000 7110 6020
rect 7050 5960 7060 6000
rect 7100 5960 7110 6000
rect 7050 5900 7110 5960
rect 7050 5860 7060 5900
rect 7100 5860 7110 5900
rect 7050 5800 7110 5860
rect 7050 5760 7060 5800
rect 7100 5760 7110 5800
rect 7050 5700 7110 5760
rect 7050 5660 7060 5700
rect 7100 5660 7110 5700
rect 7050 5600 7110 5660
rect 7050 5560 7060 5600
rect 7100 5560 7110 5600
rect 7050 5500 7110 5560
rect 7050 5460 7060 5500
rect 7100 5460 7110 5500
rect 7050 5440 7110 5460
rect 7230 6000 7290 6020
rect 7230 5960 7240 6000
rect 7280 5960 7290 6000
rect 7230 5900 7290 5960
rect 7230 5860 7240 5900
rect 7280 5860 7290 5900
rect 7230 5800 7290 5860
rect 7230 5760 7240 5800
rect 7280 5760 7290 5800
rect 7230 5700 7290 5760
rect 7230 5660 7240 5700
rect 7280 5660 7290 5700
rect 7230 5600 7290 5660
rect 7230 5560 7240 5600
rect 7280 5560 7290 5600
rect 7230 5500 7290 5560
rect 7230 5460 7240 5500
rect 7280 5460 7290 5500
rect 7230 5440 7290 5460
rect 7410 6000 7470 6020
rect 7410 5960 7420 6000
rect 7460 5960 7470 6000
rect 7410 5900 7470 5960
rect 7410 5860 7420 5900
rect 7460 5860 7470 5900
rect 7410 5800 7470 5860
rect 7410 5760 7420 5800
rect 7460 5760 7470 5800
rect 7410 5700 7470 5760
rect 7410 5660 7420 5700
rect 7460 5660 7470 5700
rect 7410 5600 7470 5660
rect 7410 5560 7420 5600
rect 7460 5560 7470 5600
rect 7410 5500 7470 5560
rect 7410 5460 7420 5500
rect 7460 5460 7470 5500
rect 7410 5440 7470 5460
rect 7590 6000 7650 6020
rect 7590 5960 7600 6000
rect 7640 5960 7650 6000
rect 7590 5900 7650 5960
rect 7590 5860 7600 5900
rect 7640 5860 7650 5900
rect 7590 5800 7650 5860
rect 7590 5760 7600 5800
rect 7640 5760 7650 5800
rect 7590 5700 7650 5760
rect 7590 5660 7600 5700
rect 7640 5660 7650 5700
rect 7590 5600 7650 5660
rect 7590 5560 7600 5600
rect 7640 5560 7650 5600
rect 7590 5500 7650 5560
rect 7590 5460 7600 5500
rect 7640 5460 7650 5500
rect 7590 5440 7650 5460
rect 7770 6000 7830 6020
rect 7770 5960 7780 6000
rect 7820 5960 7830 6000
rect 7770 5900 7830 5960
rect 7770 5860 7780 5900
rect 7820 5860 7830 5900
rect 7770 5800 7830 5860
rect 7770 5760 7780 5800
rect 7820 5760 7830 5800
rect 7770 5700 7830 5760
rect 7770 5660 7780 5700
rect 7820 5660 7830 5700
rect 7770 5600 7830 5660
rect 7770 5560 7780 5600
rect 7820 5560 7830 5600
rect 7770 5500 7830 5560
rect 7770 5460 7780 5500
rect 7820 5460 7830 5500
rect 7770 5440 7830 5460
rect 7950 6000 8010 6020
rect 7950 5960 7960 6000
rect 8000 5960 8010 6000
rect 7950 5900 8010 5960
rect 7950 5860 7960 5900
rect 8000 5860 8010 5900
rect 7950 5800 8010 5860
rect 7950 5760 7960 5800
rect 8000 5760 8010 5800
rect 7950 5700 8010 5760
rect 7950 5660 7960 5700
rect 8000 5660 8010 5700
rect 7950 5600 8010 5660
rect 7950 5560 7960 5600
rect 8000 5560 8010 5600
rect 7950 5500 8010 5560
rect 7950 5460 7960 5500
rect 8000 5460 8010 5500
rect 7950 5440 8010 5460
rect 8130 6000 8190 6020
rect 8130 5960 8140 6000
rect 8180 5960 8190 6000
rect 8130 5900 8190 5960
rect 8130 5860 8140 5900
rect 8180 5860 8190 5900
rect 8130 5800 8190 5860
rect 8130 5760 8140 5800
rect 8180 5760 8190 5800
rect 8130 5700 8190 5760
rect 8130 5660 8140 5700
rect 8180 5660 8190 5700
rect 8130 5600 8190 5660
rect 8130 5560 8140 5600
rect 8180 5560 8190 5600
rect 8130 5500 8190 5560
rect 8130 5460 8140 5500
rect 8180 5460 8190 5500
rect 8130 5440 8190 5460
rect 8310 6000 8370 6020
rect 8310 5960 8320 6000
rect 8360 5960 8370 6000
rect 8310 5900 8370 5960
rect 8310 5860 8320 5900
rect 8360 5860 8370 5900
rect 8310 5800 8370 5860
rect 8310 5760 8320 5800
rect 8360 5760 8370 5800
rect 8310 5700 8370 5760
rect 8310 5660 8320 5700
rect 8360 5660 8370 5700
rect 8310 5600 8370 5660
rect 8310 5560 8320 5600
rect 8360 5560 8370 5600
rect 8310 5500 8370 5560
rect 8310 5460 8320 5500
rect 8360 5460 8370 5500
rect 8310 5440 8370 5460
rect 8490 6000 8550 6020
rect 8490 5960 8500 6000
rect 8540 5960 8550 6000
rect 8490 5900 8550 5960
rect 8490 5860 8500 5900
rect 8540 5860 8550 5900
rect 8490 5800 8550 5860
rect 8490 5760 8500 5800
rect 8540 5760 8550 5800
rect 8490 5700 8550 5760
rect 8490 5660 8500 5700
rect 8540 5660 8550 5700
rect 8490 5600 8550 5660
rect 8490 5560 8500 5600
rect 8540 5560 8550 5600
rect 8490 5500 8550 5560
rect 8490 5460 8500 5500
rect 8540 5460 8550 5500
rect 8490 5440 8550 5460
rect 8670 6000 8730 6020
rect 8670 5960 8680 6000
rect 8720 5960 8730 6000
rect 8670 5900 8730 5960
rect 8670 5860 8680 5900
rect 8720 5860 8730 5900
rect 8670 5800 8730 5860
rect 8670 5760 8680 5800
rect 8720 5760 8730 5800
rect 8670 5700 8730 5760
rect 8670 5660 8680 5700
rect 8720 5660 8730 5700
rect 8670 5600 8730 5660
rect 8670 5560 8680 5600
rect 8720 5560 8730 5600
rect 8670 5500 8730 5560
rect 8670 5460 8680 5500
rect 8720 5460 8730 5500
rect 8670 5440 8730 5460
rect 8850 6000 8910 6020
rect 8850 5960 8860 6000
rect 8900 5960 8910 6000
rect 8850 5900 8910 5960
rect 8850 5860 8860 5900
rect 8900 5860 8910 5900
rect 8850 5800 8910 5860
rect 8850 5760 8860 5800
rect 8900 5760 8910 5800
rect 8850 5700 8910 5760
rect 8850 5660 8860 5700
rect 8900 5660 8910 5700
rect 8850 5600 8910 5660
rect 8850 5560 8860 5600
rect 8900 5560 8910 5600
rect 8850 5500 8910 5560
rect 8850 5460 8860 5500
rect 8900 5460 8910 5500
rect 8850 5440 8910 5460
rect 9030 6000 9090 6020
rect 9030 5960 9040 6000
rect 9080 5960 9090 6000
rect 9030 5900 9090 5960
rect 9030 5860 9040 5900
rect 9080 5860 9090 5900
rect 9030 5800 9090 5860
rect 9030 5760 9040 5800
rect 9080 5760 9090 5800
rect 9030 5700 9090 5760
rect 9030 5660 9040 5700
rect 9080 5660 9090 5700
rect 9030 5600 9090 5660
rect 9030 5560 9040 5600
rect 9080 5560 9090 5600
rect 9030 5500 9090 5560
rect 9030 5460 9040 5500
rect 9080 5460 9090 5500
rect 9030 5440 9090 5460
rect 9210 6000 9270 6020
rect 9210 5960 9220 6000
rect 9260 5960 9270 6000
rect 9210 5900 9270 5960
rect 9210 5860 9220 5900
rect 9260 5860 9270 5900
rect 9210 5800 9270 5860
rect 9210 5760 9220 5800
rect 9260 5760 9270 5800
rect 9210 5700 9270 5760
rect 9210 5660 9220 5700
rect 9260 5660 9270 5700
rect 9210 5600 9270 5660
rect 9210 5560 9220 5600
rect 9260 5560 9270 5600
rect 9210 5500 9270 5560
rect 9210 5460 9220 5500
rect 9260 5460 9270 5500
rect 9210 5440 9270 5460
rect 9390 6000 9450 6020
rect 9390 5960 9400 6000
rect 9440 5960 9450 6000
rect 9390 5900 9450 5960
rect 9390 5860 9400 5900
rect 9440 5860 9450 5900
rect 9390 5800 9450 5860
rect 9390 5760 9400 5800
rect 9440 5760 9450 5800
rect 9390 5700 9450 5760
rect 9390 5660 9400 5700
rect 9440 5660 9450 5700
rect 9390 5600 9450 5660
rect 9390 5560 9400 5600
rect 9440 5560 9450 5600
rect 9390 5500 9450 5560
rect 9390 5460 9400 5500
rect 9440 5460 9450 5500
rect 9390 5440 9450 5460
rect 9570 6000 9630 6020
rect 9570 5960 9580 6000
rect 9620 5960 9630 6000
rect 9570 5900 9630 5960
rect 9570 5860 9580 5900
rect 9620 5860 9630 5900
rect 9570 5800 9630 5860
rect 9570 5760 9580 5800
rect 9620 5760 9630 5800
rect 9570 5700 9630 5760
rect 9570 5660 9580 5700
rect 9620 5660 9630 5700
rect 9570 5600 9630 5660
rect 9570 5560 9580 5600
rect 9620 5560 9630 5600
rect 9570 5500 9630 5560
rect 9570 5460 9580 5500
rect 9620 5460 9630 5500
rect 9570 5440 9630 5460
rect 9750 6000 9810 6020
rect 9750 5960 9760 6000
rect 9800 5960 9810 6000
rect 9750 5900 9810 5960
rect 9750 5860 9760 5900
rect 9800 5860 9810 5900
rect 9750 5800 9810 5860
rect 9750 5760 9760 5800
rect 9800 5760 9810 5800
rect 9750 5700 9810 5760
rect 9750 5660 9760 5700
rect 9800 5660 9810 5700
rect 9750 5600 9810 5660
rect 9750 5560 9760 5600
rect 9800 5560 9810 5600
rect 9750 5500 9810 5560
rect 9750 5460 9760 5500
rect 9800 5460 9810 5500
rect 9750 5440 9810 5460
rect 9880 5810 9920 6180
rect 10580 6040 10660 6080
rect 10580 6020 10600 6040
rect 10640 6020 10660 6040
rect 6700 5400 6740 5440
rect 7060 5400 7100 5440
rect 7420 5400 7460 5440
rect 7780 5400 7820 5440
rect 8140 5400 8180 5440
rect 8500 5400 8540 5440
rect 8860 5400 8900 5440
rect 9220 5400 9260 5440
rect 9580 5400 9620 5440
rect 6680 5380 6760 5400
rect 6680 5340 6700 5380
rect 6740 5340 6760 5380
rect 6680 5320 6760 5340
rect 7040 5380 7120 5400
rect 7040 5340 7060 5380
rect 7100 5340 7120 5380
rect 7040 5320 7120 5340
rect 7400 5380 7480 5400
rect 7400 5340 7420 5380
rect 7460 5340 7480 5380
rect 7400 5320 7480 5340
rect 7760 5380 7840 5400
rect 7760 5340 7780 5380
rect 7820 5340 7840 5380
rect 7760 5320 7840 5340
rect 7940 5380 8020 5400
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 8120 5380 8200 5400
rect 8120 5340 8140 5380
rect 8180 5340 8200 5380
rect 8120 5320 8200 5340
rect 8480 5380 8560 5400
rect 8480 5340 8500 5380
rect 8540 5340 8560 5380
rect 8480 5320 8560 5340
rect 8840 5380 8920 5400
rect 8840 5340 8860 5380
rect 8900 5340 8920 5380
rect 8840 5320 8920 5340
rect 9200 5380 9280 5400
rect 9200 5340 9220 5380
rect 9260 5340 9280 5380
rect 9200 5320 9280 5340
rect 9380 5380 9460 5400
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 9560 5380 9640 5400
rect 9560 5340 9580 5380
rect 9620 5340 9640 5380
rect 9560 5320 9640 5340
rect 9880 5270 9920 5650
rect 10260 5980 10540 6020
rect 10700 5980 10980 6020
rect 10260 5810 10300 5980
rect 10380 5940 10420 5980
rect 10820 5940 10860 5980
rect 10370 5920 10430 5940
rect 10370 5880 10380 5920
rect 10420 5880 10430 5920
rect 10370 5860 10430 5880
rect 10580 5920 10660 5940
rect 10580 5880 10600 5920
rect 10640 5880 10660 5920
rect 10580 5860 10660 5880
rect 10810 5920 10870 5940
rect 10810 5880 10820 5920
rect 10860 5880 10870 5920
rect 10810 5860 10870 5880
rect 10380 5820 10420 5860
rect 10600 5820 10640 5860
rect 10820 5820 10860 5860
rect 10260 5480 10300 5650
rect 10370 5800 10430 5820
rect 10370 5760 10380 5800
rect 10420 5760 10430 5800
rect 10370 5700 10430 5760
rect 10370 5660 10380 5700
rect 10420 5660 10430 5700
rect 10370 5640 10430 5660
rect 10480 5800 10540 5820
rect 10480 5760 10490 5800
rect 10530 5760 10540 5800
rect 10480 5700 10540 5760
rect 10480 5660 10490 5700
rect 10530 5660 10540 5700
rect 10480 5640 10540 5660
rect 10590 5800 10650 5820
rect 10590 5760 10600 5800
rect 10640 5760 10650 5800
rect 10590 5700 10650 5760
rect 10590 5660 10600 5700
rect 10640 5660 10650 5700
rect 10590 5640 10650 5660
rect 10700 5800 10760 5820
rect 10700 5760 10710 5800
rect 10750 5760 10760 5800
rect 10700 5700 10760 5760
rect 10700 5660 10710 5700
rect 10750 5660 10760 5700
rect 10700 5640 10760 5660
rect 10810 5800 10870 5820
rect 10810 5760 10820 5800
rect 10860 5760 10870 5800
rect 10810 5700 10870 5760
rect 10810 5660 10820 5700
rect 10860 5660 10870 5700
rect 10810 5640 10870 5660
rect 10940 5810 10980 5980
rect 10490 5600 10530 5640
rect 10710 5600 10750 5640
rect 10450 5580 10530 5600
rect 10450 5540 10470 5580
rect 10510 5540 10530 5580
rect 10450 5520 10530 5540
rect 10580 5580 10660 5600
rect 10580 5540 10600 5580
rect 10640 5540 10660 5580
rect 10580 5520 10660 5540
rect 10710 5580 10790 5600
rect 10710 5540 10730 5580
rect 10770 5540 10790 5580
rect 10710 5520 10790 5540
rect 10940 5480 10980 5650
rect 10260 5440 10540 5480
rect 10700 5440 10980 5480
rect 6400 5230 8080 5270
rect 8240 5230 9920 5270
rect 6600 4860 6680 4880
rect 6600 4840 6620 4860
rect 6660 4840 6680 4860
rect 8680 4860 8760 4880
rect 8680 4840 8700 4860
rect 5300 4800 6560 4840
rect 6720 4800 7980 4840
rect 5300 4630 5340 4800
rect 5520 4740 5600 4760
rect 5520 4700 5540 4740
rect 5580 4700 5600 4740
rect 5520 4680 5600 4700
rect 5650 4740 5710 4760
rect 5650 4700 5660 4740
rect 5700 4700 5710 4740
rect 5650 4680 5710 4700
rect 5890 4740 5950 4760
rect 5890 4700 5900 4740
rect 5940 4700 5950 4740
rect 5890 4680 5950 4700
rect 6130 4740 6190 4760
rect 6130 4700 6140 4740
rect 6180 4700 6190 4740
rect 6130 4680 6190 4700
rect 6240 4740 6320 4760
rect 6240 4700 6260 4740
rect 6300 4700 6320 4740
rect 6240 4680 6320 4700
rect 6370 4740 6430 4760
rect 6370 4700 6380 4740
rect 6420 4700 6430 4740
rect 6370 4680 6430 4700
rect 6610 4740 6670 4760
rect 6610 4700 6620 4740
rect 6660 4700 6670 4740
rect 6610 4680 6670 4700
rect 6850 4740 6910 4760
rect 6850 4700 6860 4740
rect 6900 4700 6910 4740
rect 6850 4680 6910 4700
rect 6960 4740 7040 4760
rect 6960 4700 6980 4740
rect 7020 4700 7040 4740
rect 6960 4680 7040 4700
rect 7090 4740 7150 4760
rect 7090 4700 7100 4740
rect 7140 4700 7150 4740
rect 7090 4680 7150 4700
rect 7330 4740 7390 4760
rect 7330 4700 7340 4740
rect 7380 4700 7390 4740
rect 7330 4680 7390 4700
rect 7570 4740 7630 4760
rect 7570 4700 7580 4740
rect 7620 4700 7630 4740
rect 7570 4680 7630 4700
rect 7680 4740 7760 4760
rect 7680 4700 7700 4740
rect 7740 4700 7760 4740
rect 7680 4680 7760 4700
rect 5540 4640 5580 4680
rect 5660 4640 5700 4680
rect 5900 4640 5940 4680
rect 6140 4640 6180 4680
rect 6260 4640 6300 4680
rect 6380 4640 6420 4680
rect 6620 4640 6660 4680
rect 6860 4640 6900 4680
rect 6980 4640 7020 4680
rect 7100 4640 7140 4680
rect 7340 4640 7380 4680
rect 7580 4640 7620 4680
rect 7700 4640 7740 4680
rect 5300 4300 5340 4470
rect 5410 4620 5470 4640
rect 5410 4580 5420 4620
rect 5460 4580 5470 4620
rect 5410 4520 5470 4580
rect 5410 4480 5420 4520
rect 5460 4480 5470 4520
rect 5410 4400 5470 4480
rect 5530 4620 5590 4640
rect 5530 4580 5540 4620
rect 5580 4580 5590 4620
rect 5530 4520 5590 4580
rect 5530 4480 5540 4520
rect 5580 4480 5590 4520
rect 5530 4460 5590 4480
rect 5650 4620 5710 4640
rect 5650 4580 5660 4620
rect 5700 4580 5710 4620
rect 5650 4520 5710 4580
rect 5650 4480 5660 4520
rect 5700 4480 5710 4520
rect 5650 4460 5710 4480
rect 5770 4620 5830 4640
rect 5770 4580 5780 4620
rect 5820 4580 5830 4620
rect 5770 4520 5830 4580
rect 5770 4480 5780 4520
rect 5820 4480 5830 4520
rect 5770 4460 5830 4480
rect 5890 4620 5950 4640
rect 5890 4580 5900 4620
rect 5940 4580 5950 4620
rect 5890 4520 5950 4580
rect 5890 4480 5900 4520
rect 5940 4480 5950 4520
rect 5890 4460 5950 4480
rect 6010 4620 6070 4640
rect 6010 4580 6020 4620
rect 6060 4580 6070 4620
rect 6010 4520 6070 4580
rect 6010 4480 6020 4520
rect 6060 4480 6070 4520
rect 6010 4460 6070 4480
rect 6130 4620 6190 4640
rect 6130 4580 6140 4620
rect 6180 4580 6190 4620
rect 6130 4520 6190 4580
rect 6130 4480 6140 4520
rect 6180 4480 6190 4520
rect 6130 4460 6190 4480
rect 6250 4620 6310 4640
rect 6250 4580 6260 4620
rect 6300 4580 6310 4620
rect 6250 4520 6310 4580
rect 6250 4480 6260 4520
rect 6300 4480 6310 4520
rect 6250 4460 6310 4480
rect 6370 4620 6430 4640
rect 6370 4580 6380 4620
rect 6420 4580 6430 4620
rect 6370 4520 6430 4580
rect 6370 4480 6380 4520
rect 6420 4480 6430 4520
rect 6370 4460 6430 4480
rect 6490 4620 6550 4640
rect 6490 4580 6500 4620
rect 6540 4580 6550 4620
rect 6490 4520 6550 4580
rect 6490 4480 6500 4520
rect 6540 4480 6550 4520
rect 6490 4460 6550 4480
rect 6610 4620 6670 4640
rect 6610 4580 6620 4620
rect 6660 4580 6670 4620
rect 6610 4520 6670 4580
rect 6610 4480 6620 4520
rect 6660 4480 6670 4520
rect 6610 4460 6670 4480
rect 6730 4620 6790 4640
rect 6730 4580 6740 4620
rect 6780 4580 6790 4620
rect 6730 4520 6790 4580
rect 6730 4480 6740 4520
rect 6780 4480 6790 4520
rect 6730 4460 6790 4480
rect 6850 4620 6910 4640
rect 6850 4580 6860 4620
rect 6900 4580 6910 4620
rect 6850 4520 6910 4580
rect 6850 4480 6860 4520
rect 6900 4480 6910 4520
rect 6850 4460 6910 4480
rect 6970 4620 7030 4640
rect 6970 4580 6980 4620
rect 7020 4580 7030 4620
rect 6970 4520 7030 4580
rect 6970 4480 6980 4520
rect 7020 4480 7030 4520
rect 6970 4460 7030 4480
rect 7090 4620 7150 4640
rect 7090 4580 7100 4620
rect 7140 4580 7150 4620
rect 7090 4520 7150 4580
rect 7090 4480 7100 4520
rect 7140 4480 7150 4520
rect 7090 4460 7150 4480
rect 7210 4620 7270 4640
rect 7210 4580 7220 4620
rect 7260 4580 7270 4620
rect 7210 4520 7270 4580
rect 7210 4480 7220 4520
rect 7260 4480 7270 4520
rect 7210 4460 7270 4480
rect 7330 4620 7390 4640
rect 7330 4580 7340 4620
rect 7380 4580 7390 4620
rect 7330 4520 7390 4580
rect 7330 4480 7340 4520
rect 7380 4480 7390 4520
rect 7330 4460 7390 4480
rect 7450 4620 7510 4640
rect 7450 4580 7460 4620
rect 7500 4580 7510 4620
rect 7450 4520 7510 4580
rect 7450 4480 7460 4520
rect 7500 4480 7510 4520
rect 7450 4460 7510 4480
rect 7570 4620 7630 4640
rect 7570 4580 7580 4620
rect 7620 4580 7630 4620
rect 7570 4520 7630 4580
rect 7570 4480 7580 4520
rect 7620 4480 7630 4520
rect 7570 4460 7630 4480
rect 7690 4620 7750 4640
rect 7690 4580 7700 4620
rect 7740 4580 7750 4620
rect 7690 4520 7750 4580
rect 7690 4480 7700 4520
rect 7740 4480 7750 4520
rect 7690 4460 7750 4480
rect 7810 4620 7870 4640
rect 7810 4580 7820 4620
rect 7860 4580 7870 4620
rect 7810 4520 7870 4580
rect 7810 4480 7820 4520
rect 7860 4480 7870 4520
rect 5780 4420 5820 4460
rect 6020 4420 6060 4460
rect 6500 4420 6540 4460
rect 6740 4420 6780 4460
rect 7220 4420 7260 4460
rect 7460 4420 7500 4460
rect 5410 4360 5420 4400
rect 5460 4360 5470 4400
rect 5410 4340 5470 4360
rect 5580 4400 5660 4420
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4400 5840 4420
rect 5760 4360 5780 4400
rect 5820 4360 5840 4400
rect 5760 4340 5840 4360
rect 6000 4400 6080 4420
rect 6000 4360 6020 4400
rect 6060 4360 6080 4400
rect 6000 4340 6080 4360
rect 6240 4400 6320 4420
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4400 6560 4420
rect 6480 4360 6500 4400
rect 6540 4360 6560 4400
rect 6480 4340 6560 4360
rect 6720 4400 6800 4420
rect 6720 4360 6740 4400
rect 6780 4360 6800 4400
rect 6720 4340 6800 4360
rect 6960 4400 7040 4420
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4400 7280 4420
rect 7200 4360 7220 4400
rect 7260 4360 7280 4400
rect 7200 4340 7280 4360
rect 7440 4400 7520 4420
rect 7440 4360 7460 4400
rect 7500 4360 7520 4400
rect 7440 4340 7520 4360
rect 7630 4400 7690 4420
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 7810 4400 7870 4480
rect 7810 4360 7820 4400
rect 7860 4360 7870 4400
rect 7810 4340 7870 4360
rect 7940 4630 7980 4800
rect 5420 4300 5460 4340
rect 7820 4300 7860 4340
rect 7940 4300 7980 4470
rect 5300 4260 6560 4300
rect 6720 4260 7980 4300
rect 8340 4820 8700 4840
rect 8740 4840 8760 4860
rect 8920 4860 9000 4880
rect 8920 4840 8940 4860
rect 8740 4820 8940 4840
rect 8980 4840 9000 4860
rect 9160 4860 9240 4880
rect 9160 4840 9180 4860
rect 8980 4820 9180 4840
rect 9220 4840 9240 4860
rect 9400 4860 9480 4880
rect 9400 4840 9420 4860
rect 9220 4820 9420 4840
rect 9460 4840 9480 4860
rect 9640 4860 9720 4880
rect 9640 4840 9660 4860
rect 9700 4840 9720 4860
rect 9880 4860 9960 4880
rect 9880 4840 9900 4860
rect 9460 4820 9600 4840
rect 9760 4820 9900 4840
rect 9940 4840 9960 4860
rect 10120 4860 10200 4880
rect 10120 4840 10140 4860
rect 9940 4820 10140 4840
rect 10180 4840 10200 4860
rect 10360 4860 10440 4880
rect 10360 4840 10380 4860
rect 10180 4820 10380 4840
rect 10420 4840 10440 4860
rect 10600 4860 10680 4880
rect 10600 4840 10620 4860
rect 10420 4820 10620 4840
rect 10660 4840 10680 4860
rect 10660 4820 11020 4840
rect 8340 4800 9600 4820
rect 9760 4800 11020 4820
rect 8340 4630 8380 4800
rect 8560 4740 8640 4760
rect 8560 4700 8580 4740
rect 8620 4700 8640 4740
rect 8560 4680 8640 4700
rect 8690 4740 8750 4760
rect 8690 4700 8700 4740
rect 8740 4700 8750 4740
rect 8690 4680 8750 4700
rect 8930 4740 8990 4760
rect 8930 4700 8940 4740
rect 8980 4700 8990 4740
rect 8930 4680 8990 4700
rect 9170 4740 9230 4760
rect 9170 4700 9180 4740
rect 9220 4700 9230 4740
rect 9170 4680 9230 4700
rect 9280 4740 9360 4760
rect 9280 4700 9300 4740
rect 9340 4700 9360 4740
rect 9280 4680 9360 4700
rect 9410 4740 9470 4760
rect 9410 4700 9420 4740
rect 9460 4700 9470 4740
rect 9410 4680 9470 4700
rect 9650 4740 9710 4760
rect 9650 4700 9660 4740
rect 9700 4700 9710 4740
rect 9650 4680 9710 4700
rect 9890 4740 9950 4760
rect 9890 4700 9900 4740
rect 9940 4700 9950 4740
rect 9890 4680 9950 4700
rect 10000 4740 10080 4760
rect 10000 4700 10020 4740
rect 10060 4700 10080 4740
rect 10000 4680 10080 4700
rect 10130 4740 10190 4760
rect 10130 4700 10140 4740
rect 10180 4700 10190 4740
rect 10130 4680 10190 4700
rect 10370 4740 10430 4760
rect 10370 4700 10380 4740
rect 10420 4700 10430 4740
rect 10370 4680 10430 4700
rect 10610 4740 10670 4760
rect 10610 4700 10620 4740
rect 10660 4700 10670 4740
rect 10610 4680 10670 4700
rect 10720 4740 10800 4760
rect 10720 4700 10740 4740
rect 10780 4700 10800 4740
rect 10720 4680 10800 4700
rect 8580 4640 8620 4680
rect 8700 4640 8740 4680
rect 8940 4640 8980 4680
rect 9180 4640 9220 4680
rect 9300 4640 9340 4680
rect 9420 4640 9460 4680
rect 9660 4640 9700 4680
rect 9900 4640 9940 4680
rect 10020 4640 10060 4680
rect 10140 4640 10180 4680
rect 10380 4640 10420 4680
rect 10620 4640 10660 4680
rect 10740 4640 10780 4680
rect 8340 4300 8380 4470
rect 8450 4620 8510 4640
rect 8450 4580 8460 4620
rect 8500 4580 8510 4620
rect 8450 4520 8510 4580
rect 8450 4480 8460 4520
rect 8500 4480 8510 4520
rect 8450 4400 8510 4480
rect 8570 4620 8630 4640
rect 8570 4580 8580 4620
rect 8620 4580 8630 4620
rect 8570 4520 8630 4580
rect 8570 4480 8580 4520
rect 8620 4480 8630 4520
rect 8570 4460 8630 4480
rect 8690 4620 8750 4640
rect 8690 4580 8700 4620
rect 8740 4580 8750 4620
rect 8690 4520 8750 4580
rect 8690 4480 8700 4520
rect 8740 4480 8750 4520
rect 8690 4460 8750 4480
rect 8810 4620 8870 4640
rect 8810 4580 8820 4620
rect 8860 4580 8870 4620
rect 8810 4520 8870 4580
rect 8810 4480 8820 4520
rect 8860 4480 8870 4520
rect 8810 4460 8870 4480
rect 8930 4620 8990 4640
rect 8930 4580 8940 4620
rect 8980 4580 8990 4620
rect 8930 4520 8990 4580
rect 8930 4480 8940 4520
rect 8980 4480 8990 4520
rect 8930 4460 8990 4480
rect 9050 4620 9110 4640
rect 9050 4580 9060 4620
rect 9100 4580 9110 4620
rect 9050 4520 9110 4580
rect 9050 4480 9060 4520
rect 9100 4480 9110 4520
rect 9050 4460 9110 4480
rect 9170 4620 9230 4640
rect 9170 4580 9180 4620
rect 9220 4580 9230 4620
rect 9170 4520 9230 4580
rect 9170 4480 9180 4520
rect 9220 4480 9230 4520
rect 9170 4460 9230 4480
rect 9290 4620 9350 4640
rect 9290 4580 9300 4620
rect 9340 4580 9350 4620
rect 9290 4520 9350 4580
rect 9290 4480 9300 4520
rect 9340 4480 9350 4520
rect 9290 4460 9350 4480
rect 9410 4620 9470 4640
rect 9410 4580 9420 4620
rect 9460 4580 9470 4620
rect 9410 4520 9470 4580
rect 9410 4480 9420 4520
rect 9460 4480 9470 4520
rect 9410 4460 9470 4480
rect 9530 4620 9590 4640
rect 9530 4580 9540 4620
rect 9580 4580 9590 4620
rect 9530 4520 9590 4580
rect 9530 4480 9540 4520
rect 9580 4480 9590 4520
rect 9530 4460 9590 4480
rect 9650 4620 9710 4640
rect 9650 4580 9660 4620
rect 9700 4580 9710 4620
rect 9650 4520 9710 4580
rect 9650 4480 9660 4520
rect 9700 4480 9710 4520
rect 9650 4460 9710 4480
rect 9770 4620 9830 4640
rect 9770 4580 9780 4620
rect 9820 4580 9830 4620
rect 9770 4520 9830 4580
rect 9770 4480 9780 4520
rect 9820 4480 9830 4520
rect 9770 4460 9830 4480
rect 9890 4620 9950 4640
rect 9890 4580 9900 4620
rect 9940 4580 9950 4620
rect 9890 4520 9950 4580
rect 9890 4480 9900 4520
rect 9940 4480 9950 4520
rect 9890 4460 9950 4480
rect 10010 4620 10070 4640
rect 10010 4580 10020 4620
rect 10060 4580 10070 4620
rect 10010 4520 10070 4580
rect 10010 4480 10020 4520
rect 10060 4480 10070 4520
rect 10010 4460 10070 4480
rect 10130 4620 10190 4640
rect 10130 4580 10140 4620
rect 10180 4580 10190 4620
rect 10130 4520 10190 4580
rect 10130 4480 10140 4520
rect 10180 4480 10190 4520
rect 10130 4460 10190 4480
rect 10250 4620 10310 4640
rect 10250 4580 10260 4620
rect 10300 4580 10310 4620
rect 10250 4520 10310 4580
rect 10250 4480 10260 4520
rect 10300 4480 10310 4520
rect 10250 4460 10310 4480
rect 10370 4620 10430 4640
rect 10370 4580 10380 4620
rect 10420 4580 10430 4620
rect 10370 4520 10430 4580
rect 10370 4480 10380 4520
rect 10420 4480 10430 4520
rect 10370 4460 10430 4480
rect 10490 4620 10550 4640
rect 10490 4580 10500 4620
rect 10540 4580 10550 4620
rect 10490 4520 10550 4580
rect 10490 4480 10500 4520
rect 10540 4480 10550 4520
rect 10490 4460 10550 4480
rect 10610 4620 10670 4640
rect 10610 4580 10620 4620
rect 10660 4580 10670 4620
rect 10610 4520 10670 4580
rect 10610 4480 10620 4520
rect 10660 4480 10670 4520
rect 10610 4460 10670 4480
rect 10730 4620 10790 4640
rect 10730 4580 10740 4620
rect 10780 4580 10790 4620
rect 10730 4520 10790 4580
rect 10730 4480 10740 4520
rect 10780 4480 10790 4520
rect 10730 4460 10790 4480
rect 10850 4620 10910 4640
rect 10850 4580 10860 4620
rect 10900 4580 10910 4620
rect 10850 4520 10910 4580
rect 10850 4480 10860 4520
rect 10900 4480 10910 4520
rect 8820 4420 8860 4460
rect 9060 4420 9100 4460
rect 9540 4420 9580 4460
rect 9780 4420 9820 4460
rect 10260 4420 10300 4460
rect 10500 4420 10540 4460
rect 8450 4360 8460 4400
rect 8500 4360 8510 4400
rect 8450 4340 8510 4360
rect 8630 4400 8690 4420
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 8800 4400 8880 4420
rect 8800 4360 8820 4400
rect 8860 4360 8880 4400
rect 8800 4340 8880 4360
rect 9040 4400 9120 4420
rect 9040 4360 9060 4400
rect 9100 4360 9120 4400
rect 9040 4340 9120 4360
rect 9280 4400 9360 4420
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9520 4400 9600 4420
rect 9520 4360 9540 4400
rect 9580 4360 9600 4400
rect 9520 4340 9600 4360
rect 9760 4400 9840 4420
rect 9760 4360 9780 4400
rect 9820 4360 9840 4400
rect 9760 4340 9840 4360
rect 10000 4400 10080 4420
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10240 4400 10320 4420
rect 10240 4360 10260 4400
rect 10300 4360 10320 4400
rect 10240 4340 10320 4360
rect 10480 4400 10560 4420
rect 10480 4360 10500 4400
rect 10540 4360 10560 4400
rect 10480 4340 10560 4360
rect 10660 4400 10740 4420
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 10850 4400 10910 4480
rect 10850 4360 10860 4400
rect 10900 4360 10910 4400
rect 10850 4340 10910 4360
rect 10980 4630 11020 4800
rect 8460 4300 8500 4340
rect 10860 4300 10900 4340
rect 10980 4300 11020 4470
rect 8340 4260 9600 4300
rect 9760 4260 11020 4300
rect 250 4030 4270 4110
rect -90 3430 260 3450
rect -90 3390 -70 3430
rect -30 3390 30 3430
rect 70 3390 130 3430
rect 170 3390 260 3430
rect -90 3370 260 3390
rect 1300 2750 1550 4030
rect 2660 2750 2910 4030
rect 4020 2750 4270 4030
rect 6160 4140 6820 4180
rect 6980 4140 7640 4180
rect 6160 3930 6200 4140
rect 6380 4080 6460 4100
rect 6380 4040 6400 4080
rect 6440 4040 6460 4080
rect 6380 4020 6460 4040
rect 6260 3990 6340 4010
rect 6260 3950 6280 3990
rect 6320 3950 6340 3990
rect 6260 3930 6340 3950
rect 6510 3990 6570 4010
rect 6510 3950 6520 3990
rect 6560 3950 6570 3990
rect 6510 3930 6570 3950
rect 6740 3990 6820 4010
rect 6740 3950 6760 3990
rect 6800 3950 6820 3990
rect 6740 3930 6820 3950
rect 6990 3990 7050 4010
rect 6990 3950 7000 3990
rect 7040 3950 7050 3990
rect 6990 3930 7050 3950
rect 7220 3990 7300 4010
rect 7220 3950 7240 3990
rect 7280 3950 7300 3990
rect 7220 3930 7300 3950
rect 7470 3990 7530 4010
rect 7470 3950 7480 3990
rect 7520 3950 7530 3990
rect 7470 3930 7530 3950
rect 7600 3930 7640 4140
rect 6280 3890 6320 3930
rect 6520 3890 6560 3930
rect 6760 3890 6800 3930
rect 7000 3890 7040 3930
rect 7240 3890 7280 3930
rect 7480 3890 7520 3930
rect 6270 3870 6330 3890
rect 6270 3830 6280 3870
rect 6320 3830 6330 3870
rect 6270 3810 6330 3830
rect 6390 3870 6450 3890
rect 6390 3830 6400 3870
rect 6440 3830 6450 3870
rect 6390 3810 6450 3830
rect 6510 3870 6570 3890
rect 6510 3830 6520 3870
rect 6560 3830 6570 3870
rect 6510 3810 6570 3830
rect 6630 3870 6690 3890
rect 6630 3830 6640 3870
rect 6680 3830 6690 3870
rect 6630 3810 6690 3830
rect 6750 3870 6810 3890
rect 6750 3830 6760 3870
rect 6800 3830 6810 3870
rect 6750 3810 6810 3830
rect 6870 3870 6930 3890
rect 6870 3830 6880 3870
rect 6920 3830 6930 3870
rect 6870 3810 6930 3830
rect 6990 3870 7050 3890
rect 6990 3830 7000 3870
rect 7040 3830 7050 3870
rect 6990 3810 7050 3830
rect 7110 3870 7170 3890
rect 7110 3830 7120 3870
rect 7160 3830 7170 3870
rect 7110 3810 7170 3830
rect 7230 3870 7290 3890
rect 7230 3830 7240 3870
rect 7280 3830 7290 3870
rect 7230 3810 7290 3830
rect 7350 3870 7410 3890
rect 7350 3830 7360 3870
rect 7400 3830 7410 3870
rect 7350 3810 7410 3830
rect 7470 3870 7530 3890
rect 7470 3830 7480 3870
rect 7520 3830 7530 3870
rect 7470 3810 7530 3830
rect 7580 3810 7600 3890
rect 8680 4140 9340 4180
rect 9500 4140 10160 4180
rect 8680 3930 8720 4140
rect 9860 4080 9940 4100
rect 9860 4040 9880 4080
rect 9920 4040 9940 4080
rect 9860 4020 9940 4040
rect 8790 3990 8850 4010
rect 8790 3950 8800 3990
rect 8840 3950 8850 3990
rect 8790 3930 8850 3950
rect 9020 3990 9100 4010
rect 9020 3950 9040 3990
rect 9080 3950 9100 3990
rect 9020 3930 9100 3950
rect 9270 3990 9330 4010
rect 9270 3950 9280 3990
rect 9320 3950 9330 3990
rect 9270 3930 9330 3950
rect 9500 3990 9580 4010
rect 9500 3950 9520 3990
rect 9560 3950 9580 3990
rect 9500 3930 9580 3950
rect 9750 3990 9810 4010
rect 9750 3950 9760 3990
rect 9800 3950 9810 3990
rect 9750 3930 9810 3950
rect 9980 3990 10060 4010
rect 9980 3950 10000 3990
rect 10040 3950 10060 3990
rect 9980 3930 10060 3950
rect 10120 3930 10160 4140
rect 6400 3770 6440 3810
rect 6640 3770 6680 3810
rect 6880 3770 6920 3810
rect 7120 3770 7160 3810
rect 7360 3770 7400 3810
rect 7640 3810 7660 3890
rect 8660 3810 8680 3890
rect 8800 3890 8840 3930
rect 9040 3890 9080 3930
rect 9280 3890 9320 3930
rect 9520 3890 9560 3930
rect 9760 3890 9800 3930
rect 10000 3890 10040 3930
rect 6160 3650 6200 3770
rect 6260 3750 6340 3770
rect 6260 3710 6280 3750
rect 6320 3710 6340 3750
rect 6260 3690 6340 3710
rect 6390 3750 6450 3770
rect 6390 3710 6400 3750
rect 6440 3710 6450 3750
rect 6390 3690 6450 3710
rect 6630 3750 6690 3770
rect 6630 3710 6640 3750
rect 6680 3710 6690 3750
rect 6630 3690 6690 3710
rect 6870 3750 6930 3770
rect 6870 3710 6880 3750
rect 6920 3710 6930 3750
rect 6870 3690 6930 3710
rect 7110 3750 7170 3770
rect 7110 3710 7120 3750
rect 7160 3710 7170 3750
rect 7110 3690 7170 3710
rect 7350 3750 7410 3770
rect 7350 3710 7360 3750
rect 7400 3710 7410 3750
rect 7350 3690 7410 3710
rect 7600 3650 7640 3770
rect 6160 3610 6820 3650
rect 6980 3610 7640 3650
rect 8720 3810 8740 3890
rect 8790 3870 8850 3890
rect 8790 3830 8800 3870
rect 8840 3830 8850 3870
rect 8790 3810 8850 3830
rect 8910 3870 8970 3890
rect 8910 3830 8920 3870
rect 8960 3830 8970 3870
rect 8910 3810 8970 3830
rect 9030 3870 9090 3890
rect 9030 3830 9040 3870
rect 9080 3830 9090 3870
rect 9030 3810 9090 3830
rect 9150 3870 9210 3890
rect 9150 3830 9160 3870
rect 9200 3830 9210 3870
rect 9150 3810 9210 3830
rect 9270 3870 9330 3890
rect 9270 3830 9280 3870
rect 9320 3830 9330 3870
rect 9270 3810 9330 3830
rect 9390 3870 9450 3890
rect 9390 3830 9400 3870
rect 9440 3830 9450 3870
rect 9390 3810 9450 3830
rect 9510 3870 9570 3890
rect 9510 3830 9520 3870
rect 9560 3830 9570 3870
rect 9510 3810 9570 3830
rect 9630 3870 9690 3890
rect 9630 3830 9640 3870
rect 9680 3830 9690 3870
rect 9630 3810 9690 3830
rect 9750 3870 9810 3890
rect 9750 3830 9760 3870
rect 9800 3830 9810 3870
rect 9750 3810 9810 3830
rect 9870 3870 9930 3890
rect 9870 3830 9880 3870
rect 9920 3830 9930 3870
rect 9870 3810 9930 3830
rect 9990 3870 10050 3890
rect 9990 3830 10000 3870
rect 10040 3830 10050 3870
rect 9990 3810 10050 3830
rect 8920 3770 8960 3810
rect 9160 3770 9200 3810
rect 9400 3770 9440 3810
rect 9640 3770 9680 3810
rect 9880 3770 9920 3810
rect 8680 3650 8720 3770
rect 8910 3750 8970 3770
rect 8910 3710 8920 3750
rect 8960 3710 8970 3750
rect 8910 3690 8970 3710
rect 9150 3750 9210 3770
rect 9150 3710 9160 3750
rect 9200 3710 9210 3750
rect 9150 3690 9210 3710
rect 9390 3750 9450 3770
rect 9390 3710 9400 3750
rect 9440 3710 9450 3750
rect 9390 3690 9450 3710
rect 9630 3750 9690 3770
rect 9630 3710 9640 3750
rect 9680 3710 9690 3750
rect 9630 3690 9690 3710
rect 9870 3750 9930 3770
rect 9870 3710 9880 3750
rect 9920 3710 9930 3750
rect 9870 3690 9930 3710
rect 9980 3750 10060 3770
rect 9980 3710 10000 3750
rect 10040 3710 10060 3750
rect 9980 3690 10060 3710
rect 10120 3650 10160 3770
rect 8680 3610 10160 3650
rect 35970 4110 36360 4150
rect 36520 4110 36910 4150
rect 35970 3940 36010 4110
rect 36090 4070 36130 4110
rect 36750 4070 36790 4110
rect 36070 4050 36150 4070
rect 36070 4010 36090 4050
rect 36130 4010 36150 4050
rect 36070 3990 36150 4010
rect 36290 4050 36370 4070
rect 36290 4010 36310 4050
rect 36350 4010 36370 4050
rect 36290 3990 36370 4010
rect 36410 4050 36470 4070
rect 36410 4010 36420 4050
rect 36460 4010 36470 4050
rect 36410 3990 36470 4010
rect 36510 4050 36590 4070
rect 36510 4010 36530 4050
rect 36570 4010 36590 4050
rect 36510 3990 36590 4010
rect 36630 4050 36690 4070
rect 36630 4010 36640 4050
rect 36680 4010 36690 4050
rect 36630 3990 36690 4010
rect 36730 4050 36810 4070
rect 36730 4010 36750 4050
rect 36790 4010 36810 4050
rect 36730 3990 36810 4010
rect 36090 3950 36130 3990
rect 36310 3950 36350 3990
rect 36530 3950 36570 3990
rect 36640 3950 36680 3990
rect 36750 3950 36790 3990
rect 35970 3610 36010 3780
rect 36080 3930 36140 3950
rect 36080 3786 36090 3930
rect 36130 3786 36140 3930
rect 36080 3770 36140 3786
rect 36190 3930 36250 3950
rect 36190 3786 36200 3930
rect 36240 3786 36250 3930
rect 36190 3770 36250 3786
rect 36300 3930 36360 3950
rect 36300 3786 36310 3930
rect 36350 3786 36360 3930
rect 36300 3770 36360 3786
rect 36410 3930 36470 3950
rect 36410 3786 36420 3930
rect 36460 3786 36470 3930
rect 36410 3770 36470 3786
rect 36520 3930 36580 3950
rect 36520 3786 36530 3930
rect 36570 3786 36580 3930
rect 36520 3770 36580 3786
rect 36630 3930 36690 3950
rect 36630 3786 36640 3930
rect 36680 3786 36690 3930
rect 36630 3770 36690 3786
rect 36740 3930 36800 3950
rect 36740 3786 36750 3930
rect 36790 3786 36800 3930
rect 36740 3770 36800 3786
rect 36870 3940 36910 4110
rect 36200 3730 36240 3770
rect 36420 3730 36460 3770
rect 36640 3730 36680 3770
rect 36180 3710 36260 3730
rect 36180 3670 36200 3710
rect 36240 3670 36260 3710
rect 36180 3650 36260 3670
rect 36400 3710 36480 3730
rect 36400 3670 36420 3710
rect 36460 3670 36480 3710
rect 36400 3650 36480 3670
rect 36620 3710 36700 3730
rect 36620 3670 36640 3710
rect 36680 3670 36700 3710
rect 36620 3650 36700 3670
rect 36870 3610 36910 3780
rect 9860 3570 9940 3610
rect 35970 3570 36360 3610
rect 36520 3570 36910 3610
rect 37250 4110 38080 4150
rect 38240 4110 39070 4150
rect 37250 3940 37290 4110
rect 37370 4070 37410 4110
rect 38690 4070 38730 4110
rect 37350 4050 37430 4070
rect 37350 4010 37370 4050
rect 37410 4010 37430 4050
rect 37350 3990 37430 4010
rect 37570 4050 37650 4070
rect 37570 4010 37590 4050
rect 37630 4010 37650 4050
rect 37570 3990 37650 4010
rect 37790 4050 37870 4070
rect 37790 4010 37810 4050
rect 37850 4010 37870 4050
rect 37790 3990 37870 4010
rect 38010 4050 38090 4070
rect 38010 4010 38030 4050
rect 38070 4010 38090 4050
rect 38010 3990 38090 4010
rect 38130 4050 38190 4070
rect 38130 4010 38140 4050
rect 38180 4010 38190 4050
rect 38130 3990 38190 4010
rect 38230 4050 38310 4070
rect 38230 4010 38250 4050
rect 38290 4010 38310 4050
rect 38230 3990 38310 4010
rect 38450 4050 38530 4070
rect 38450 4010 38470 4050
rect 38510 4010 38530 4050
rect 38450 3990 38530 4010
rect 38570 4050 38630 4070
rect 38570 4010 38580 4050
rect 38620 4010 38630 4050
rect 38570 3990 38630 4010
rect 38670 4050 38750 4070
rect 38670 4010 38690 4050
rect 38730 4010 38750 4050
rect 38670 3990 38750 4010
rect 37370 3950 37410 3990
rect 37590 3950 37630 3990
rect 37810 3950 37850 3990
rect 38030 3950 38070 3990
rect 38250 3950 38290 3990
rect 38470 3950 38510 3990
rect 38580 3950 38620 3990
rect 38690 3950 38730 3990
rect 37250 3610 37290 3780
rect 37360 3930 37420 3950
rect 37360 3890 37370 3930
rect 37410 3890 37420 3930
rect 37360 3830 37420 3890
rect 37360 3790 37370 3830
rect 37410 3790 37420 3830
rect 37360 3770 37420 3790
rect 37470 3930 37530 3950
rect 37470 3890 37480 3930
rect 37520 3890 37530 3930
rect 37470 3830 37530 3890
rect 37470 3790 37480 3830
rect 37520 3790 37530 3830
rect 37470 3770 37530 3790
rect 37580 3930 37640 3950
rect 37580 3890 37590 3930
rect 37630 3890 37640 3930
rect 37580 3830 37640 3890
rect 37580 3790 37590 3830
rect 37630 3790 37640 3830
rect 37580 3770 37640 3790
rect 37690 3930 37750 3950
rect 37690 3890 37700 3930
rect 37740 3890 37750 3930
rect 37690 3830 37750 3890
rect 37690 3790 37700 3830
rect 37740 3790 37750 3830
rect 37690 3770 37750 3790
rect 37800 3930 37860 3950
rect 37800 3890 37810 3930
rect 37850 3890 37860 3930
rect 37800 3830 37860 3890
rect 37800 3790 37810 3830
rect 37850 3790 37860 3830
rect 37800 3770 37860 3790
rect 37910 3930 37970 3950
rect 37910 3890 37920 3930
rect 37960 3890 37970 3930
rect 37910 3830 37970 3890
rect 37910 3790 37920 3830
rect 37960 3790 37970 3830
rect 37910 3770 37970 3790
rect 38020 3930 38080 3950
rect 38020 3890 38030 3930
rect 38070 3890 38080 3930
rect 38020 3830 38080 3890
rect 38020 3790 38030 3830
rect 38070 3790 38080 3830
rect 38020 3770 38080 3790
rect 38130 3930 38190 3950
rect 38130 3890 38140 3930
rect 38180 3890 38190 3930
rect 38130 3830 38190 3890
rect 38130 3790 38140 3830
rect 38180 3790 38190 3830
rect 38130 3770 38190 3790
rect 38240 3930 38300 3950
rect 38240 3890 38250 3930
rect 38290 3890 38300 3930
rect 38240 3830 38300 3890
rect 38240 3790 38250 3830
rect 38290 3790 38300 3830
rect 38240 3770 38300 3790
rect 38350 3930 38410 3950
rect 38350 3890 38360 3930
rect 38400 3890 38410 3930
rect 38350 3830 38410 3890
rect 38350 3790 38360 3830
rect 38400 3790 38410 3830
rect 38350 3770 38410 3790
rect 38460 3930 38520 3950
rect 38460 3890 38470 3930
rect 38510 3890 38520 3930
rect 38460 3830 38520 3890
rect 38460 3790 38470 3830
rect 38510 3790 38520 3830
rect 38460 3770 38520 3790
rect 38570 3930 38630 3950
rect 38570 3890 38580 3930
rect 38620 3890 38630 3930
rect 38570 3830 38630 3890
rect 38570 3790 38580 3830
rect 38620 3790 38630 3830
rect 38570 3770 38630 3790
rect 38680 3930 38740 3950
rect 38680 3890 38690 3930
rect 38730 3890 38740 3930
rect 38680 3830 38740 3890
rect 38680 3790 38690 3830
rect 38730 3790 38740 3830
rect 38680 3770 38740 3790
rect 39030 3940 39070 4110
rect 37480 3730 37520 3770
rect 37700 3730 37740 3770
rect 37920 3730 37960 3770
rect 38140 3730 38180 3770
rect 38360 3730 38400 3770
rect 38580 3730 38620 3770
rect 37460 3710 37540 3730
rect 37460 3670 37480 3710
rect 37520 3670 37540 3710
rect 37460 3650 37540 3670
rect 37680 3710 37760 3730
rect 37680 3670 37700 3710
rect 37740 3670 37760 3710
rect 37680 3650 37760 3670
rect 37900 3710 37980 3730
rect 37900 3670 37920 3710
rect 37960 3670 37980 3710
rect 37900 3650 37980 3670
rect 38120 3710 38200 3730
rect 38120 3670 38140 3710
rect 38180 3670 38200 3710
rect 38120 3650 38200 3670
rect 38340 3710 38420 3730
rect 38340 3670 38360 3710
rect 38400 3670 38420 3710
rect 38340 3650 38420 3670
rect 38560 3710 38640 3730
rect 38560 3670 38580 3710
rect 38620 3670 38640 3710
rect 38560 3650 38640 3670
rect 39030 3610 39070 3780
rect 37250 3570 38080 3610
rect 38240 3570 39070 3610
rect 39410 4110 39800 4150
rect 39960 4110 40350 4150
rect 39410 3940 39450 4110
rect 39530 4070 39570 4110
rect 40190 4070 40230 4110
rect 39510 4050 39590 4070
rect 39510 4010 39530 4050
rect 39570 4010 39590 4050
rect 39510 3990 39590 4010
rect 39730 4050 39810 4070
rect 39730 4010 39750 4050
rect 39790 4010 39810 4050
rect 39730 3990 39810 4010
rect 39850 4050 39910 4070
rect 39850 4010 39860 4050
rect 39900 4010 39910 4050
rect 39850 3990 39910 4010
rect 39950 4050 40030 4070
rect 39950 4010 39970 4050
rect 40010 4010 40030 4050
rect 39950 3990 40030 4010
rect 40170 4050 40250 4070
rect 40170 4010 40190 4050
rect 40230 4010 40250 4050
rect 40170 3990 40250 4010
rect 39530 3950 39570 3990
rect 39750 3950 39790 3990
rect 39970 3950 40010 3990
rect 40190 3950 40230 3990
rect 39410 3610 39450 3780
rect 39520 3930 39580 3950
rect 39520 3790 39530 3930
rect 39570 3790 39580 3930
rect 39520 3770 39580 3790
rect 39630 3930 39690 3950
rect 39630 3790 39640 3930
rect 39680 3790 39690 3930
rect 39630 3770 39690 3790
rect 39740 3930 39800 3950
rect 39740 3790 39750 3930
rect 39790 3790 39800 3930
rect 39740 3770 39800 3790
rect 39850 3930 39910 3950
rect 39850 3790 39860 3930
rect 39900 3790 39910 3930
rect 39850 3770 39910 3790
rect 39960 3930 40020 3950
rect 39960 3790 39970 3930
rect 40010 3790 40020 3930
rect 39960 3770 40020 3790
rect 40070 3930 40130 3950
rect 40070 3790 40080 3930
rect 40120 3790 40130 3930
rect 40070 3770 40130 3790
rect 40180 3930 40240 3950
rect 40180 3790 40190 3930
rect 40230 3790 40240 3930
rect 40180 3770 40240 3790
rect 40310 3940 40350 4110
rect 39640 3730 39680 3770
rect 39860 3730 39900 3770
rect 40080 3730 40120 3770
rect 39620 3710 39700 3730
rect 39620 3670 39640 3710
rect 39680 3670 39700 3710
rect 39620 3650 39700 3670
rect 39840 3710 39920 3730
rect 39840 3670 39860 3710
rect 39900 3670 39920 3710
rect 39840 3650 39920 3670
rect 40060 3710 40140 3730
rect 40060 3670 40080 3710
rect 40120 3670 40140 3710
rect 40060 3650 40140 3670
rect 40310 3610 40350 3780
rect 39410 3570 39800 3610
rect 39930 3570 40350 3610
rect 250 2670 4270 2750
rect 1300 1380 1550 2670
rect 2660 1380 2910 2670
rect 4020 1390 4270 2670
rect 5680 3490 6820 3530
rect 6980 3490 8120 3530
rect 5680 3180 5720 3490
rect 5960 3430 6040 3450
rect 5780 3400 5860 3420
rect 5780 3360 5800 3400
rect 5840 3360 5860 3400
rect 5960 3390 5980 3430
rect 6020 3390 6040 3430
rect 5960 3370 6040 3390
rect 6200 3430 6280 3450
rect 6200 3390 6220 3430
rect 6260 3390 6280 3430
rect 6200 3370 6280 3390
rect 6440 3430 6520 3450
rect 6440 3390 6460 3430
rect 6500 3390 6520 3430
rect 6440 3370 6520 3390
rect 6680 3430 6760 3450
rect 6680 3390 6700 3430
rect 6740 3390 6760 3430
rect 6680 3370 6760 3390
rect 7160 3430 7240 3450
rect 7160 3390 7180 3430
rect 7220 3390 7240 3430
rect 7160 3370 7240 3390
rect 7400 3430 7480 3450
rect 7400 3390 7420 3430
rect 7460 3390 7480 3430
rect 7400 3370 7480 3390
rect 7640 3430 7720 3450
rect 7640 3390 7660 3430
rect 7700 3390 7720 3430
rect 7640 3370 7720 3390
rect 7940 3400 8020 3420
rect 5780 3340 5860 3360
rect 7940 3360 7960 3400
rect 8000 3360 8020 3400
rect 7940 3340 8020 3360
rect 5680 2700 5720 3020
rect 5790 3320 5850 3340
rect 5790 3280 5800 3320
rect 5840 3280 5850 3320
rect 5790 3220 5850 3280
rect 5790 3180 5800 3220
rect 5840 3180 5850 3220
rect 5790 3120 5850 3180
rect 5790 3080 5800 3120
rect 5840 3080 5850 3120
rect 5790 3020 5850 3080
rect 5790 2980 5800 3020
rect 5840 2980 5850 3020
rect 5790 2920 5850 2980
rect 5790 2880 5800 2920
rect 5840 2880 5850 2920
rect 5790 2860 5850 2880
rect 6870 3320 6930 3340
rect 6870 3280 6880 3320
rect 6920 3280 6930 3320
rect 6870 3220 6930 3280
rect 6870 3180 6880 3220
rect 6920 3180 6930 3220
rect 6870 3120 6930 3180
rect 6870 3080 6880 3120
rect 6920 3080 6930 3120
rect 6870 3020 6930 3080
rect 6870 2980 6880 3020
rect 6920 2980 6930 3020
rect 6870 2920 6930 2980
rect 6870 2880 6880 2920
rect 6920 2880 6930 2920
rect 6870 2860 6930 2880
rect 7950 3320 8010 3340
rect 7950 3280 7960 3320
rect 8000 3280 8010 3320
rect 7950 3220 8010 3280
rect 7950 3180 7960 3220
rect 8000 3180 8010 3220
rect 7950 3120 8010 3180
rect 7950 3080 7960 3120
rect 8000 3080 8010 3120
rect 7950 3020 8010 3080
rect 7950 2980 7960 3020
rect 8000 2980 8010 3020
rect 7950 2920 8010 2980
rect 7950 2880 7960 2920
rect 8000 2880 8010 2920
rect 7950 2860 8010 2880
rect 8080 3180 8120 3490
rect 6880 2820 6920 2860
rect 6860 2800 6940 2820
rect 6860 2760 6880 2800
rect 6920 2760 6940 2800
rect 6860 2740 6940 2760
rect 6880 2700 6920 2740
rect 8080 2700 8120 3020
rect 5680 2660 6820 2700
rect 6980 2660 8120 2700
rect 8200 3490 9340 3530
rect 9500 3490 10640 3530
rect 8200 3180 8240 3490
rect 8600 3430 8680 3450
rect 8300 3400 8380 3420
rect 8300 3360 8320 3400
rect 8360 3360 8380 3400
rect 8600 3390 8620 3430
rect 8660 3390 8680 3430
rect 8600 3370 8680 3390
rect 8840 3430 8920 3450
rect 8840 3390 8860 3430
rect 8900 3390 8920 3430
rect 8840 3370 8920 3390
rect 9080 3430 9160 3450
rect 9080 3390 9100 3430
rect 9140 3390 9160 3430
rect 9080 3370 9160 3390
rect 9560 3430 9640 3450
rect 9560 3390 9580 3430
rect 9620 3390 9640 3430
rect 9560 3370 9640 3390
rect 9800 3430 9880 3450
rect 9800 3390 9820 3430
rect 9860 3390 9880 3430
rect 9800 3370 9880 3390
rect 10040 3430 10120 3450
rect 10040 3390 10060 3430
rect 10100 3390 10120 3430
rect 10040 3370 10120 3390
rect 10280 3430 10360 3450
rect 10280 3390 10300 3430
rect 10340 3390 10360 3430
rect 10280 3370 10360 3390
rect 10460 3400 10540 3420
rect 8300 3340 8380 3360
rect 10460 3360 10480 3400
rect 10520 3360 10540 3400
rect 10460 3340 10540 3360
rect 8200 2700 8240 3020
rect 8310 3320 8370 3340
rect 8310 3280 8320 3320
rect 8360 3280 8370 3320
rect 8310 3220 8370 3280
rect 8310 3180 8320 3220
rect 8360 3180 8370 3220
rect 8310 3120 8370 3180
rect 8310 3080 8320 3120
rect 8360 3080 8370 3120
rect 8310 3020 8370 3080
rect 8310 2980 8320 3020
rect 8360 2980 8370 3020
rect 8310 2920 8370 2980
rect 8310 2880 8320 2920
rect 8360 2880 8370 2920
rect 8310 2860 8370 2880
rect 9390 3320 9450 3340
rect 9390 3280 9400 3320
rect 9440 3280 9450 3320
rect 9390 3220 9450 3280
rect 9390 3180 9400 3220
rect 9440 3180 9450 3220
rect 9390 3120 9450 3180
rect 9390 3080 9400 3120
rect 9440 3080 9450 3120
rect 9390 3020 9450 3080
rect 9390 2980 9400 3020
rect 9440 2980 9450 3020
rect 9390 2920 9450 2980
rect 9390 2880 9400 2920
rect 9440 2880 9450 2920
rect 9390 2860 9450 2880
rect 10470 3320 10530 3340
rect 10470 3280 10480 3320
rect 10520 3280 10530 3320
rect 10470 3220 10530 3280
rect 10470 3180 10480 3220
rect 10520 3180 10530 3220
rect 10470 3120 10530 3180
rect 10470 3080 10480 3120
rect 10520 3080 10530 3120
rect 10470 3020 10530 3080
rect 10470 2980 10480 3020
rect 10520 2980 10530 3020
rect 10470 2920 10530 2980
rect 10470 2880 10480 2920
rect 10520 2880 10530 2920
rect 10470 2860 10530 2880
rect 10600 3180 10640 3490
rect 36400 3180 38080 3220
rect 38240 3180 39920 3220
rect 35650 3040 35730 3060
rect 35650 3020 35670 3040
rect 35710 3020 35730 3040
rect 9400 2820 9440 2860
rect 9380 2800 9460 2820
rect 9380 2760 9400 2800
rect 9440 2760 9460 2800
rect 9380 2740 9460 2760
rect 9400 2700 9440 2740
rect 10600 2700 10640 3020
rect 8200 2660 9340 2700
rect 9500 2660 10640 2700
rect 35330 2980 35610 3020
rect 35770 2980 36050 3020
rect 35330 2810 35370 2980
rect 35450 2940 35490 2980
rect 35890 2940 35930 2980
rect 5880 2560 8080 2600
rect 8240 2560 10430 2600
rect 5880 2390 5920 2560
rect 6040 2500 6120 2520
rect 6040 2460 6060 2500
rect 6100 2460 6120 2500
rect 6040 2440 6120 2460
rect 6200 2500 6280 2520
rect 6200 2460 6220 2500
rect 6260 2460 6280 2500
rect 6200 2440 6280 2460
rect 6360 2500 6440 2520
rect 6360 2460 6380 2500
rect 6420 2460 6440 2500
rect 6360 2440 6440 2460
rect 6520 2500 6600 2520
rect 6520 2460 6540 2500
rect 6580 2460 6600 2500
rect 6520 2440 6600 2460
rect 6680 2500 6760 2520
rect 6680 2460 6700 2500
rect 6740 2460 6760 2500
rect 6680 2440 6760 2460
rect 6840 2500 6920 2520
rect 6840 2460 6860 2500
rect 6900 2460 6920 2500
rect 6840 2440 6920 2460
rect 7000 2500 7080 2520
rect 7000 2460 7020 2500
rect 7060 2460 7080 2500
rect 7000 2440 7080 2460
rect 7160 2500 7240 2520
rect 7160 2460 7180 2500
rect 7220 2460 7240 2500
rect 7160 2440 7240 2460
rect 7320 2500 7400 2520
rect 7320 2460 7340 2500
rect 7380 2460 7400 2500
rect 7320 2440 7400 2460
rect 7480 2500 7560 2520
rect 7480 2460 7500 2500
rect 7540 2460 7560 2500
rect 7480 2440 7560 2460
rect 7640 2500 7720 2520
rect 7640 2460 7660 2500
rect 7700 2460 7720 2500
rect 7640 2440 7720 2460
rect 7800 2500 7880 2520
rect 7800 2460 7820 2500
rect 7860 2460 7880 2500
rect 7800 2440 7880 2460
rect 7960 2500 8040 2520
rect 7960 2460 7980 2500
rect 8020 2460 8040 2500
rect 7960 2440 8040 2460
rect 8120 2500 8200 2520
rect 8120 2460 8140 2500
rect 8180 2460 8200 2500
rect 8120 2440 8200 2460
rect 8280 2500 8360 2520
rect 8280 2460 8300 2500
rect 8340 2460 8360 2500
rect 8280 2440 8360 2460
rect 8440 2500 8520 2520
rect 8440 2460 8460 2500
rect 8500 2460 8520 2500
rect 8440 2440 8520 2460
rect 8600 2500 8680 2520
rect 8600 2460 8620 2500
rect 8660 2460 8680 2500
rect 8600 2440 8680 2460
rect 8760 2500 8840 2520
rect 8760 2460 8780 2500
rect 8820 2460 8840 2500
rect 8760 2440 8840 2460
rect 8920 2500 9000 2520
rect 8920 2460 8940 2500
rect 8980 2460 9000 2500
rect 8920 2440 9000 2460
rect 9080 2500 9160 2520
rect 9080 2460 9100 2500
rect 9140 2460 9160 2500
rect 9080 2440 9160 2460
rect 9240 2500 9320 2520
rect 9240 2460 9260 2500
rect 9300 2460 9320 2500
rect 9240 2440 9320 2460
rect 9400 2500 9480 2520
rect 9400 2460 9420 2500
rect 9460 2460 9480 2500
rect 9400 2440 9480 2460
rect 9560 2500 9640 2520
rect 9560 2460 9580 2500
rect 9620 2460 9640 2500
rect 9560 2440 9640 2460
rect 9720 2500 9800 2520
rect 9720 2460 9740 2500
rect 9780 2460 9800 2500
rect 9720 2440 9800 2460
rect 9880 2500 9960 2520
rect 9880 2460 9900 2500
rect 9940 2460 9960 2500
rect 9880 2440 9960 2460
rect 10040 2500 10120 2520
rect 10040 2460 10060 2500
rect 10100 2460 10120 2500
rect 10040 2440 10120 2460
rect 6060 2400 6100 2440
rect 8140 2400 8180 2440
rect 6050 2380 6110 2400
rect 6050 2350 6060 2380
rect 5960 2340 6060 2350
rect 6100 2340 6110 2380
rect 5960 2330 6110 2340
rect 5960 2290 5980 2330
rect 6020 2290 6110 2330
rect 5960 2280 6110 2290
rect 5960 2270 6060 2280
rect 5880 2150 5920 2230
rect 6050 2240 6060 2270
rect 6100 2240 6110 2280
rect 6050 2220 6110 2240
rect 8130 2380 8190 2400
rect 8130 2340 8140 2380
rect 8180 2340 8190 2380
rect 8130 2280 8190 2340
rect 8130 2240 8140 2280
rect 8180 2240 8190 2280
rect 8130 2220 8190 2240
rect 10210 2380 10270 2400
rect 10210 2340 10220 2380
rect 10260 2350 10270 2380
rect 10390 2390 10430 2560
rect 35330 2480 35370 2650
rect 35440 2920 35500 2940
rect 35440 2880 35450 2920
rect 35490 2880 35500 2920
rect 35440 2800 35500 2880
rect 35650 2920 35730 2940
rect 35650 2880 35670 2920
rect 35710 2880 35730 2920
rect 35650 2860 35730 2880
rect 35880 2920 35940 2940
rect 35880 2880 35890 2920
rect 35930 2880 35940 2920
rect 35670 2820 35710 2860
rect 35440 2760 35450 2800
rect 35490 2760 35500 2800
rect 35440 2700 35500 2760
rect 35440 2660 35450 2700
rect 35490 2660 35500 2700
rect 35440 2640 35500 2660
rect 35550 2800 35610 2820
rect 35550 2760 35560 2800
rect 35600 2760 35610 2800
rect 35550 2700 35610 2760
rect 35550 2660 35560 2700
rect 35600 2660 35610 2700
rect 35550 2640 35610 2660
rect 35660 2800 35720 2820
rect 35660 2760 35670 2800
rect 35710 2760 35720 2800
rect 35660 2700 35720 2760
rect 35660 2660 35670 2700
rect 35710 2660 35720 2700
rect 35660 2640 35720 2660
rect 35770 2800 35830 2820
rect 35770 2760 35780 2800
rect 35820 2760 35830 2800
rect 35770 2700 35830 2760
rect 35770 2660 35780 2700
rect 35820 2660 35830 2700
rect 35770 2640 35830 2660
rect 35880 2800 35940 2880
rect 35880 2760 35890 2800
rect 35930 2760 35940 2800
rect 35880 2700 35940 2760
rect 35880 2660 35890 2700
rect 35930 2660 35940 2700
rect 35880 2640 35940 2660
rect 36010 2810 36050 2980
rect 35560 2600 35600 2640
rect 35780 2600 35820 2640
rect 35520 2580 35600 2600
rect 35520 2540 35540 2580
rect 35580 2540 35600 2580
rect 35520 2520 35600 2540
rect 35650 2580 35730 2600
rect 35650 2540 35670 2580
rect 35710 2540 35730 2580
rect 35650 2520 35730 2540
rect 35780 2580 35860 2600
rect 35780 2540 35800 2580
rect 35840 2540 35860 2580
rect 35780 2520 35860 2540
rect 36010 2480 36050 2650
rect 35330 2440 35610 2480
rect 35770 2440 36050 2480
rect 36400 2810 36440 3180
rect 36520 3140 36560 3180
rect 39760 3140 39800 3180
rect 36500 3120 36580 3140
rect 36500 3080 36520 3120
rect 36560 3080 36580 3120
rect 36500 3060 36580 3080
rect 36860 3120 36940 3140
rect 36860 3080 36880 3120
rect 36920 3080 36940 3120
rect 36860 3060 36940 3080
rect 37220 3120 37300 3140
rect 37220 3080 37240 3120
rect 37280 3080 37300 3120
rect 37220 3060 37300 3080
rect 37580 3120 37660 3140
rect 37580 3080 37600 3120
rect 37640 3080 37660 3120
rect 37580 3060 37660 3080
rect 37940 3120 38020 3140
rect 37940 3080 37960 3120
rect 38000 3080 38020 3120
rect 37940 3060 38020 3080
rect 38300 3120 38380 3140
rect 38300 3080 38320 3120
rect 38360 3080 38380 3120
rect 38300 3060 38380 3080
rect 38660 3120 38740 3140
rect 38660 3080 38680 3120
rect 38720 3080 38740 3120
rect 38660 3060 38740 3080
rect 39020 3120 39100 3140
rect 39020 3080 39040 3120
rect 39080 3080 39100 3120
rect 39020 3060 39100 3080
rect 39380 3120 39460 3140
rect 39380 3080 39400 3120
rect 39440 3080 39460 3120
rect 39380 3060 39460 3080
rect 39740 3120 39820 3140
rect 39740 3080 39760 3120
rect 39800 3080 39820 3120
rect 39740 3060 39820 3080
rect 36520 3020 36560 3060
rect 36880 3020 36920 3060
rect 37240 3020 37280 3060
rect 37600 3020 37640 3060
rect 37960 3020 38000 3060
rect 38320 3020 38360 3060
rect 38680 3020 38720 3060
rect 39040 3020 39080 3060
rect 39400 3020 39440 3060
rect 39760 3020 39800 3060
rect 10260 2340 10350 2350
rect 10210 2330 10350 2340
rect 10210 2290 10290 2330
rect 10330 2290 10350 2330
rect 10210 2280 10350 2290
rect 10210 2240 10220 2280
rect 10260 2270 10350 2280
rect 10260 2240 10270 2270
rect 10210 2220 10270 2240
rect 36400 2270 36440 2650
rect 36510 3000 36570 3020
rect 36510 2960 36520 3000
rect 36560 2960 36570 3000
rect 36510 2900 36570 2960
rect 36510 2860 36520 2900
rect 36560 2860 36570 2900
rect 36510 2800 36570 2860
rect 36510 2760 36520 2800
rect 36560 2760 36570 2800
rect 36510 2700 36570 2760
rect 36510 2660 36520 2700
rect 36560 2660 36570 2700
rect 36510 2600 36570 2660
rect 36510 2560 36520 2600
rect 36560 2560 36570 2600
rect 36510 2500 36570 2560
rect 36510 2460 36520 2500
rect 36560 2460 36570 2500
rect 36510 2440 36570 2460
rect 36690 3000 36750 3020
rect 36690 2960 36700 3000
rect 36740 2960 36750 3000
rect 36690 2900 36750 2960
rect 36690 2860 36700 2900
rect 36740 2860 36750 2900
rect 36690 2800 36750 2860
rect 36690 2760 36700 2800
rect 36740 2760 36750 2800
rect 36690 2700 36750 2760
rect 36690 2660 36700 2700
rect 36740 2660 36750 2700
rect 36690 2600 36750 2660
rect 36690 2560 36700 2600
rect 36740 2560 36750 2600
rect 36690 2500 36750 2560
rect 36690 2460 36700 2500
rect 36740 2460 36750 2500
rect 36690 2440 36750 2460
rect 36870 3000 36930 3020
rect 36870 2960 36880 3000
rect 36920 2960 36930 3000
rect 36870 2900 36930 2960
rect 36870 2860 36880 2900
rect 36920 2860 36930 2900
rect 36870 2800 36930 2860
rect 36870 2760 36880 2800
rect 36920 2760 36930 2800
rect 36870 2700 36930 2760
rect 36870 2660 36880 2700
rect 36920 2660 36930 2700
rect 36870 2600 36930 2660
rect 36870 2560 36880 2600
rect 36920 2560 36930 2600
rect 36870 2500 36930 2560
rect 36870 2460 36880 2500
rect 36920 2460 36930 2500
rect 36870 2440 36930 2460
rect 37050 3000 37110 3020
rect 37050 2960 37060 3000
rect 37100 2960 37110 3000
rect 37050 2900 37110 2960
rect 37050 2860 37060 2900
rect 37100 2860 37110 2900
rect 37050 2800 37110 2860
rect 37050 2760 37060 2800
rect 37100 2760 37110 2800
rect 37050 2700 37110 2760
rect 37050 2660 37060 2700
rect 37100 2660 37110 2700
rect 37050 2600 37110 2660
rect 37050 2560 37060 2600
rect 37100 2560 37110 2600
rect 37050 2500 37110 2560
rect 37050 2460 37060 2500
rect 37100 2460 37110 2500
rect 37050 2440 37110 2460
rect 37230 3000 37290 3020
rect 37230 2960 37240 3000
rect 37280 2960 37290 3000
rect 37230 2900 37290 2960
rect 37230 2860 37240 2900
rect 37280 2860 37290 2900
rect 37230 2800 37290 2860
rect 37230 2760 37240 2800
rect 37280 2760 37290 2800
rect 37230 2700 37290 2760
rect 37230 2660 37240 2700
rect 37280 2660 37290 2700
rect 37230 2600 37290 2660
rect 37230 2560 37240 2600
rect 37280 2560 37290 2600
rect 37230 2500 37290 2560
rect 37230 2460 37240 2500
rect 37280 2460 37290 2500
rect 37230 2440 37290 2460
rect 37410 3000 37470 3020
rect 37410 2960 37420 3000
rect 37460 2960 37470 3000
rect 37410 2900 37470 2960
rect 37410 2860 37420 2900
rect 37460 2860 37470 2900
rect 37410 2800 37470 2860
rect 37410 2760 37420 2800
rect 37460 2760 37470 2800
rect 37410 2700 37470 2760
rect 37410 2660 37420 2700
rect 37460 2660 37470 2700
rect 37410 2600 37470 2660
rect 37410 2560 37420 2600
rect 37460 2560 37470 2600
rect 37410 2500 37470 2560
rect 37410 2460 37420 2500
rect 37460 2460 37470 2500
rect 37410 2440 37470 2460
rect 37590 3000 37650 3020
rect 37590 2960 37600 3000
rect 37640 2960 37650 3000
rect 37590 2900 37650 2960
rect 37590 2860 37600 2900
rect 37640 2860 37650 2900
rect 37590 2800 37650 2860
rect 37590 2760 37600 2800
rect 37640 2760 37650 2800
rect 37590 2700 37650 2760
rect 37590 2660 37600 2700
rect 37640 2660 37650 2700
rect 37590 2600 37650 2660
rect 37590 2560 37600 2600
rect 37640 2560 37650 2600
rect 37590 2500 37650 2560
rect 37590 2460 37600 2500
rect 37640 2460 37650 2500
rect 37590 2440 37650 2460
rect 37770 3000 37830 3020
rect 37770 2960 37780 3000
rect 37820 2960 37830 3000
rect 37770 2900 37830 2960
rect 37770 2860 37780 2900
rect 37820 2860 37830 2900
rect 37770 2800 37830 2860
rect 37770 2760 37780 2800
rect 37820 2760 37830 2800
rect 37770 2700 37830 2760
rect 37770 2660 37780 2700
rect 37820 2660 37830 2700
rect 37770 2600 37830 2660
rect 37770 2560 37780 2600
rect 37820 2560 37830 2600
rect 37770 2500 37830 2560
rect 37770 2460 37780 2500
rect 37820 2460 37830 2500
rect 37770 2440 37830 2460
rect 37950 3000 38010 3020
rect 37950 2960 37960 3000
rect 38000 2960 38010 3000
rect 37950 2900 38010 2960
rect 37950 2860 37960 2900
rect 38000 2860 38010 2900
rect 37950 2800 38010 2860
rect 37950 2760 37960 2800
rect 38000 2760 38010 2800
rect 37950 2700 38010 2760
rect 37950 2660 37960 2700
rect 38000 2660 38010 2700
rect 37950 2600 38010 2660
rect 37950 2560 37960 2600
rect 38000 2560 38010 2600
rect 37950 2500 38010 2560
rect 37950 2460 37960 2500
rect 38000 2460 38010 2500
rect 37950 2440 38010 2460
rect 38130 3000 38190 3020
rect 38130 2960 38140 3000
rect 38180 2960 38190 3000
rect 38130 2900 38190 2960
rect 38130 2860 38140 2900
rect 38180 2860 38190 2900
rect 38130 2800 38190 2860
rect 38130 2760 38140 2800
rect 38180 2760 38190 2800
rect 38130 2700 38190 2760
rect 38130 2660 38140 2700
rect 38180 2660 38190 2700
rect 38130 2600 38190 2660
rect 38130 2560 38140 2600
rect 38180 2560 38190 2600
rect 38130 2500 38190 2560
rect 38130 2460 38140 2500
rect 38180 2460 38190 2500
rect 38130 2440 38190 2460
rect 38310 3000 38370 3020
rect 38310 2960 38320 3000
rect 38360 2960 38370 3000
rect 38310 2900 38370 2960
rect 38310 2860 38320 2900
rect 38360 2860 38370 2900
rect 38310 2800 38370 2860
rect 38310 2760 38320 2800
rect 38360 2760 38370 2800
rect 38310 2700 38370 2760
rect 38310 2660 38320 2700
rect 38360 2660 38370 2700
rect 38310 2600 38370 2660
rect 38310 2560 38320 2600
rect 38360 2560 38370 2600
rect 38310 2500 38370 2560
rect 38310 2460 38320 2500
rect 38360 2460 38370 2500
rect 38310 2440 38370 2460
rect 38490 3000 38550 3020
rect 38490 2960 38500 3000
rect 38540 2960 38550 3000
rect 38490 2900 38550 2960
rect 38490 2860 38500 2900
rect 38540 2860 38550 2900
rect 38490 2800 38550 2860
rect 38490 2760 38500 2800
rect 38540 2760 38550 2800
rect 38490 2700 38550 2760
rect 38490 2660 38500 2700
rect 38540 2660 38550 2700
rect 38490 2600 38550 2660
rect 38490 2560 38500 2600
rect 38540 2560 38550 2600
rect 38490 2500 38550 2560
rect 38490 2460 38500 2500
rect 38540 2460 38550 2500
rect 38490 2440 38550 2460
rect 38670 3000 38730 3020
rect 38670 2960 38680 3000
rect 38720 2960 38730 3000
rect 38670 2900 38730 2960
rect 38670 2860 38680 2900
rect 38720 2860 38730 2900
rect 38670 2800 38730 2860
rect 38670 2760 38680 2800
rect 38720 2760 38730 2800
rect 38670 2700 38730 2760
rect 38670 2660 38680 2700
rect 38720 2660 38730 2700
rect 38670 2600 38730 2660
rect 38670 2560 38680 2600
rect 38720 2560 38730 2600
rect 38670 2500 38730 2560
rect 38670 2460 38680 2500
rect 38720 2460 38730 2500
rect 38670 2440 38730 2460
rect 38850 3000 38910 3020
rect 38850 2960 38860 3000
rect 38900 2960 38910 3000
rect 38850 2900 38910 2960
rect 38850 2860 38860 2900
rect 38900 2860 38910 2900
rect 38850 2800 38910 2860
rect 38850 2760 38860 2800
rect 38900 2760 38910 2800
rect 38850 2700 38910 2760
rect 38850 2660 38860 2700
rect 38900 2660 38910 2700
rect 38850 2600 38910 2660
rect 38850 2560 38860 2600
rect 38900 2560 38910 2600
rect 38850 2500 38910 2560
rect 38850 2460 38860 2500
rect 38900 2460 38910 2500
rect 38850 2440 38910 2460
rect 39030 3000 39090 3020
rect 39030 2960 39040 3000
rect 39080 2960 39090 3000
rect 39030 2900 39090 2960
rect 39030 2860 39040 2900
rect 39080 2860 39090 2900
rect 39030 2800 39090 2860
rect 39030 2760 39040 2800
rect 39080 2760 39090 2800
rect 39030 2700 39090 2760
rect 39030 2660 39040 2700
rect 39080 2660 39090 2700
rect 39030 2600 39090 2660
rect 39030 2560 39040 2600
rect 39080 2560 39090 2600
rect 39030 2500 39090 2560
rect 39030 2460 39040 2500
rect 39080 2460 39090 2500
rect 39030 2440 39090 2460
rect 39210 3000 39270 3020
rect 39210 2960 39220 3000
rect 39260 2960 39270 3000
rect 39210 2900 39270 2960
rect 39210 2860 39220 2900
rect 39260 2860 39270 2900
rect 39210 2800 39270 2860
rect 39210 2760 39220 2800
rect 39260 2760 39270 2800
rect 39210 2700 39270 2760
rect 39210 2660 39220 2700
rect 39260 2660 39270 2700
rect 39210 2600 39270 2660
rect 39210 2560 39220 2600
rect 39260 2560 39270 2600
rect 39210 2500 39270 2560
rect 39210 2460 39220 2500
rect 39260 2460 39270 2500
rect 39210 2440 39270 2460
rect 39390 3000 39450 3020
rect 39390 2960 39400 3000
rect 39440 2960 39450 3000
rect 39390 2900 39450 2960
rect 39390 2860 39400 2900
rect 39440 2860 39450 2900
rect 39390 2800 39450 2860
rect 39390 2760 39400 2800
rect 39440 2760 39450 2800
rect 39390 2700 39450 2760
rect 39390 2660 39400 2700
rect 39440 2660 39450 2700
rect 39390 2600 39450 2660
rect 39390 2560 39400 2600
rect 39440 2560 39450 2600
rect 39390 2500 39450 2560
rect 39390 2460 39400 2500
rect 39440 2460 39450 2500
rect 39390 2440 39450 2460
rect 39570 3000 39630 3020
rect 39570 2960 39580 3000
rect 39620 2960 39630 3000
rect 39570 2900 39630 2960
rect 39570 2860 39580 2900
rect 39620 2860 39630 2900
rect 39570 2800 39630 2860
rect 39570 2760 39580 2800
rect 39620 2760 39630 2800
rect 39570 2700 39630 2760
rect 39570 2660 39580 2700
rect 39620 2660 39630 2700
rect 39570 2600 39630 2660
rect 39570 2560 39580 2600
rect 39620 2560 39630 2600
rect 39570 2500 39630 2560
rect 39570 2460 39580 2500
rect 39620 2460 39630 2500
rect 39570 2440 39630 2460
rect 39750 3000 39810 3020
rect 39750 2960 39760 3000
rect 39800 2960 39810 3000
rect 39750 2900 39810 2960
rect 39750 2860 39760 2900
rect 39800 2860 39810 2900
rect 39750 2800 39810 2860
rect 39750 2760 39760 2800
rect 39800 2760 39810 2800
rect 39750 2700 39810 2760
rect 39750 2660 39760 2700
rect 39800 2660 39810 2700
rect 39750 2600 39810 2660
rect 39750 2560 39760 2600
rect 39800 2560 39810 2600
rect 39750 2500 39810 2560
rect 39750 2460 39760 2500
rect 39800 2460 39810 2500
rect 39750 2440 39810 2460
rect 39880 2810 39920 3180
rect 40580 3040 40660 3080
rect 40580 3020 40600 3040
rect 40640 3020 40660 3040
rect 36700 2400 36740 2440
rect 37060 2400 37100 2440
rect 37420 2400 37460 2440
rect 37780 2400 37820 2440
rect 38140 2400 38180 2440
rect 38500 2400 38540 2440
rect 38860 2400 38900 2440
rect 39220 2400 39260 2440
rect 39580 2400 39620 2440
rect 36680 2380 36760 2400
rect 36680 2340 36700 2380
rect 36740 2340 36760 2380
rect 36680 2320 36760 2340
rect 37040 2380 37120 2400
rect 37040 2340 37060 2380
rect 37100 2340 37120 2380
rect 37040 2320 37120 2340
rect 37400 2380 37480 2400
rect 37400 2340 37420 2380
rect 37460 2340 37480 2380
rect 37400 2320 37480 2340
rect 37760 2380 37840 2400
rect 37760 2340 37780 2380
rect 37820 2340 37840 2380
rect 37760 2320 37840 2340
rect 37940 2380 38020 2400
rect 37940 2340 37960 2380
rect 38000 2340 38020 2380
rect 37940 2320 38020 2340
rect 38120 2380 38200 2400
rect 38120 2340 38140 2380
rect 38180 2340 38200 2380
rect 38120 2320 38200 2340
rect 38480 2380 38560 2400
rect 38480 2340 38500 2380
rect 38540 2340 38560 2380
rect 38480 2320 38560 2340
rect 38840 2380 38920 2400
rect 38840 2340 38860 2380
rect 38900 2340 38920 2380
rect 38840 2320 38920 2340
rect 39200 2380 39280 2400
rect 39200 2340 39220 2380
rect 39260 2340 39280 2380
rect 39200 2320 39280 2340
rect 39380 2380 39460 2400
rect 39380 2340 39400 2380
rect 39440 2340 39460 2380
rect 39380 2320 39460 2340
rect 39560 2380 39640 2400
rect 39560 2340 39580 2380
rect 39620 2340 39640 2380
rect 39560 2320 39640 2340
rect 39880 2270 39920 2650
rect 40260 2980 40540 3020
rect 40700 2980 40980 3020
rect 40260 2810 40300 2980
rect 40380 2940 40420 2980
rect 40820 2940 40860 2980
rect 40370 2920 40430 2940
rect 40370 2880 40380 2920
rect 40420 2880 40430 2920
rect 40370 2860 40430 2880
rect 40580 2920 40660 2940
rect 40580 2880 40600 2920
rect 40640 2880 40660 2920
rect 40580 2860 40660 2880
rect 40810 2920 40870 2940
rect 40810 2880 40820 2920
rect 40860 2880 40870 2920
rect 40810 2860 40870 2880
rect 40380 2820 40420 2860
rect 40600 2820 40640 2860
rect 40820 2820 40860 2860
rect 40260 2480 40300 2650
rect 40370 2800 40430 2820
rect 40370 2760 40380 2800
rect 40420 2760 40430 2800
rect 40370 2700 40430 2760
rect 40370 2660 40380 2700
rect 40420 2660 40430 2700
rect 40370 2640 40430 2660
rect 40480 2800 40540 2820
rect 40480 2760 40490 2800
rect 40530 2760 40540 2800
rect 40480 2700 40540 2760
rect 40480 2660 40490 2700
rect 40530 2660 40540 2700
rect 40480 2640 40540 2660
rect 40590 2800 40650 2820
rect 40590 2760 40600 2800
rect 40640 2760 40650 2800
rect 40590 2700 40650 2760
rect 40590 2660 40600 2700
rect 40640 2660 40650 2700
rect 40590 2640 40650 2660
rect 40700 2800 40760 2820
rect 40700 2760 40710 2800
rect 40750 2760 40760 2800
rect 40700 2700 40760 2760
rect 40700 2660 40710 2700
rect 40750 2660 40760 2700
rect 40700 2640 40760 2660
rect 40810 2800 40870 2820
rect 40810 2760 40820 2800
rect 40860 2760 40870 2800
rect 40810 2700 40870 2760
rect 40810 2660 40820 2700
rect 40860 2660 40870 2700
rect 40810 2640 40870 2660
rect 40940 2810 40980 2980
rect 40490 2600 40530 2640
rect 40710 2600 40750 2640
rect 40450 2580 40530 2600
rect 40450 2540 40470 2580
rect 40510 2540 40530 2580
rect 40450 2520 40530 2540
rect 40580 2580 40660 2600
rect 40580 2540 40600 2580
rect 40640 2540 40660 2580
rect 40580 2520 40660 2540
rect 40710 2580 40790 2600
rect 40710 2540 40730 2580
rect 40770 2540 40790 2580
rect 40710 2520 40790 2540
rect 40940 2480 40980 2650
rect 40260 2440 40540 2480
rect 40700 2440 40980 2480
rect 36400 2230 38080 2270
rect 38240 2230 39920 2270
rect 10390 2150 10430 2230
rect 5880 2110 8080 2150
rect 8240 2110 10430 2150
rect 6240 2010 6800 2050
rect 6960 2010 7400 2050
rect 6240 1840 6280 2010
rect 6560 1950 6640 1970
rect 6560 1910 6580 1950
rect 6620 1910 6640 1950
rect 6560 1890 6640 1910
rect 6780 1950 6860 1970
rect 6780 1910 6800 1950
rect 6840 1910 6860 1950
rect 6780 1890 6860 1910
rect 6900 1950 6960 1970
rect 6900 1910 6910 1950
rect 6950 1910 6960 1950
rect 6900 1890 6960 1910
rect 7000 1950 7080 1970
rect 7000 1910 7020 1950
rect 7060 1910 7080 1950
rect 7000 1890 7080 1910
rect 6580 1850 6620 1890
rect 6800 1850 6840 1890
rect 7020 1850 7060 1890
rect 6240 1510 6280 1680
rect 6350 1830 6410 1850
rect 6350 1790 6360 1830
rect 6400 1790 6410 1830
rect 6350 1730 6410 1790
rect 6350 1690 6360 1730
rect 6400 1690 6410 1730
rect 6350 1610 6410 1690
rect 6460 1830 6520 1850
rect 6460 1790 6470 1830
rect 6510 1790 6520 1830
rect 6460 1730 6520 1790
rect 6460 1690 6470 1730
rect 6510 1690 6520 1730
rect 6460 1670 6520 1690
rect 6570 1830 6630 1850
rect 6570 1790 6580 1830
rect 6620 1790 6630 1830
rect 6570 1730 6630 1790
rect 6570 1690 6580 1730
rect 6620 1690 6630 1730
rect 6570 1670 6630 1690
rect 6680 1830 6740 1850
rect 6680 1790 6690 1830
rect 6730 1790 6740 1830
rect 6680 1730 6740 1790
rect 6680 1690 6690 1730
rect 6730 1690 6740 1730
rect 6680 1670 6740 1690
rect 6790 1830 6850 1850
rect 6790 1790 6800 1830
rect 6840 1790 6850 1830
rect 6790 1730 6850 1790
rect 6790 1690 6800 1730
rect 6840 1690 6850 1730
rect 6790 1670 6850 1690
rect 6900 1830 6960 1850
rect 6900 1790 6910 1830
rect 6950 1790 6960 1830
rect 6900 1730 6960 1790
rect 6900 1690 6910 1730
rect 6950 1690 6960 1730
rect 6900 1670 6960 1690
rect 7010 1830 7070 1850
rect 7010 1790 7020 1830
rect 7060 1790 7070 1830
rect 7010 1730 7070 1790
rect 7010 1690 7020 1730
rect 7060 1690 7070 1730
rect 7010 1670 7070 1690
rect 7120 1830 7180 1850
rect 7120 1790 7130 1830
rect 7170 1790 7180 1830
rect 7120 1730 7180 1790
rect 7120 1690 7130 1730
rect 7170 1690 7180 1730
rect 7120 1670 7180 1690
rect 7230 1830 7290 1850
rect 7230 1790 7240 1830
rect 7280 1790 7290 1830
rect 7230 1730 7290 1790
rect 7230 1690 7240 1730
rect 7280 1690 7290 1730
rect 6470 1630 6510 1670
rect 6690 1630 6730 1670
rect 6910 1630 6950 1670
rect 7130 1630 7170 1670
rect 6350 1570 6360 1610
rect 6400 1570 6410 1610
rect 6350 1550 6410 1570
rect 6450 1610 6530 1630
rect 6450 1570 6470 1610
rect 6510 1570 6530 1610
rect 6450 1550 6530 1570
rect 6670 1610 6750 1630
rect 6670 1570 6690 1610
rect 6730 1570 6750 1610
rect 6670 1550 6750 1570
rect 6890 1610 6970 1630
rect 6890 1570 6910 1610
rect 6950 1570 6970 1610
rect 6890 1550 6970 1570
rect 7110 1610 7190 1630
rect 7110 1570 7130 1610
rect 7170 1570 7190 1610
rect 7110 1550 7190 1570
rect 7230 1610 7290 1690
rect 7230 1570 7240 1610
rect 7280 1570 7290 1610
rect 7230 1550 7290 1570
rect 7360 1840 7400 2010
rect 6360 1510 6400 1550
rect 7240 1510 7280 1550
rect 7360 1510 7400 1680
rect 6240 1470 7400 1510
rect 7470 2010 8080 2050
rect 8240 2010 8850 2050
rect 7470 1840 7510 2010
rect 7790 1950 7870 1970
rect 7790 1910 7810 1950
rect 7850 1910 7870 1950
rect 7790 1890 7870 1910
rect 8010 1950 8090 1970
rect 8010 1910 8030 1950
rect 8070 1910 8090 1950
rect 8010 1890 8090 1910
rect 8130 1950 8190 1970
rect 8130 1910 8140 1950
rect 8180 1910 8190 1950
rect 8130 1890 8190 1910
rect 8230 1950 8310 1970
rect 8230 1910 8250 1950
rect 8290 1910 8310 1950
rect 8230 1890 8310 1910
rect 8450 1950 8530 1970
rect 8450 1910 8470 1950
rect 8510 1910 8530 1950
rect 8450 1890 8530 1910
rect 7810 1850 7850 1890
rect 8030 1850 8070 1890
rect 8250 1850 8290 1890
rect 8470 1850 8510 1890
rect 7470 1510 7510 1680
rect 7580 1830 7640 1850
rect 7580 1790 7590 1830
rect 7630 1790 7640 1830
rect 7580 1730 7640 1790
rect 7580 1690 7590 1730
rect 7630 1690 7640 1730
rect 7580 1610 7640 1690
rect 7690 1830 7750 1850
rect 7690 1790 7700 1830
rect 7740 1790 7750 1830
rect 7690 1730 7750 1790
rect 7690 1690 7700 1730
rect 7740 1690 7750 1730
rect 7690 1670 7750 1690
rect 7800 1830 7860 1850
rect 7800 1790 7810 1830
rect 7850 1790 7860 1830
rect 7800 1730 7860 1790
rect 7800 1690 7810 1730
rect 7850 1690 7860 1730
rect 7800 1670 7860 1690
rect 7910 1830 7970 1850
rect 7910 1790 7920 1830
rect 7960 1790 7970 1830
rect 7910 1730 7970 1790
rect 7910 1690 7920 1730
rect 7960 1690 7970 1730
rect 7910 1670 7970 1690
rect 8020 1830 8080 1850
rect 8020 1790 8030 1830
rect 8070 1790 8080 1830
rect 8020 1730 8080 1790
rect 8020 1690 8030 1730
rect 8070 1690 8080 1730
rect 8020 1670 8080 1690
rect 8130 1830 8190 1850
rect 8130 1790 8140 1830
rect 8180 1790 8190 1830
rect 8130 1730 8190 1790
rect 8130 1690 8140 1730
rect 8180 1690 8190 1730
rect 8130 1670 8190 1690
rect 8240 1830 8300 1850
rect 8240 1790 8250 1830
rect 8290 1790 8300 1830
rect 8240 1730 8300 1790
rect 8240 1690 8250 1730
rect 8290 1690 8300 1730
rect 8240 1670 8300 1690
rect 8350 1830 8410 1850
rect 8350 1790 8360 1830
rect 8400 1790 8410 1830
rect 8350 1730 8410 1790
rect 8350 1690 8360 1730
rect 8400 1690 8410 1730
rect 8350 1670 8410 1690
rect 8460 1830 8520 1850
rect 8460 1790 8470 1830
rect 8510 1790 8520 1830
rect 8460 1730 8520 1790
rect 8460 1690 8470 1730
rect 8510 1690 8520 1730
rect 8460 1670 8520 1690
rect 8570 1830 8630 1850
rect 8570 1790 8580 1830
rect 8620 1790 8630 1830
rect 8570 1730 8630 1790
rect 8570 1690 8580 1730
rect 8620 1690 8630 1730
rect 8570 1670 8630 1690
rect 8680 1830 8740 1850
rect 8680 1790 8690 1830
rect 8730 1790 8740 1830
rect 8680 1730 8740 1790
rect 8680 1690 8690 1730
rect 8730 1690 8740 1730
rect 7580 1570 7590 1610
rect 7630 1570 7640 1610
rect 7580 1550 7640 1570
rect 7700 1630 7740 1670
rect 7920 1630 7960 1670
rect 8140 1630 8180 1670
rect 8360 1630 8400 1670
rect 8580 1630 8620 1670
rect 7700 1610 7810 1630
rect 7700 1570 7750 1610
rect 7790 1570 7810 1610
rect 7700 1550 7810 1570
rect 7900 1610 7980 1630
rect 7900 1570 7920 1610
rect 7960 1570 7980 1610
rect 7900 1550 7980 1570
rect 8120 1610 8200 1630
rect 8120 1570 8140 1610
rect 8180 1570 8200 1610
rect 8120 1550 8200 1570
rect 8340 1610 8420 1630
rect 8340 1570 8360 1610
rect 8400 1570 8420 1610
rect 8340 1550 8420 1570
rect 8560 1610 8640 1630
rect 8560 1570 8580 1610
rect 8620 1570 8640 1610
rect 8560 1550 8640 1570
rect 8680 1610 8740 1690
rect 8680 1570 8690 1610
rect 8730 1570 8740 1610
rect 8680 1550 8740 1570
rect 8810 1840 8850 2010
rect 7590 1510 7630 1550
rect 8690 1510 8730 1550
rect 8810 1510 8850 1680
rect 7470 1470 8080 1510
rect 8240 1470 8850 1510
rect 8920 2010 9360 2050
rect 9520 2010 10080 2050
rect 8920 1840 8960 2010
rect 9240 1950 9320 1970
rect 9240 1910 9260 1950
rect 9300 1910 9320 1950
rect 9240 1890 9320 1910
rect 9360 1950 9420 1970
rect 9360 1910 9370 1950
rect 9410 1910 9420 1950
rect 9360 1890 9420 1910
rect 9460 1950 9540 1970
rect 9460 1910 9480 1950
rect 9520 1910 9540 1950
rect 9460 1890 9540 1910
rect 9680 1950 9760 1970
rect 9680 1910 9700 1950
rect 9740 1910 9760 1950
rect 9680 1890 9760 1910
rect 9260 1850 9300 1890
rect 9480 1850 9520 1890
rect 9700 1850 9740 1890
rect 8920 1510 8960 1680
rect 9030 1830 9090 1850
rect 9030 1790 9040 1830
rect 9080 1790 9090 1830
rect 9030 1730 9090 1790
rect 9030 1690 9040 1730
rect 9080 1690 9090 1730
rect 9030 1610 9090 1690
rect 9140 1830 9200 1850
rect 9140 1790 9150 1830
rect 9190 1790 9200 1830
rect 9140 1730 9200 1790
rect 9140 1690 9150 1730
rect 9190 1690 9200 1730
rect 9140 1670 9200 1690
rect 9250 1830 9310 1850
rect 9250 1790 9260 1830
rect 9300 1790 9310 1830
rect 9250 1730 9310 1790
rect 9250 1690 9260 1730
rect 9300 1690 9310 1730
rect 9250 1670 9310 1690
rect 9360 1830 9420 1850
rect 9360 1790 9370 1830
rect 9410 1790 9420 1830
rect 9360 1730 9420 1790
rect 9360 1690 9370 1730
rect 9410 1690 9420 1730
rect 9360 1670 9420 1690
rect 9470 1830 9530 1850
rect 9470 1790 9480 1830
rect 9520 1790 9530 1830
rect 9470 1730 9530 1790
rect 9470 1690 9480 1730
rect 9520 1690 9530 1730
rect 9470 1670 9530 1690
rect 9580 1830 9640 1850
rect 9580 1790 9590 1830
rect 9630 1790 9640 1830
rect 9580 1730 9640 1790
rect 9580 1690 9590 1730
rect 9630 1690 9640 1730
rect 9580 1670 9640 1690
rect 9690 1830 9750 1850
rect 9690 1790 9700 1830
rect 9740 1790 9750 1830
rect 9690 1730 9750 1790
rect 9690 1690 9700 1730
rect 9740 1690 9750 1730
rect 9690 1670 9750 1690
rect 9800 1830 9860 1850
rect 9800 1790 9810 1830
rect 9850 1790 9860 1830
rect 9800 1730 9860 1790
rect 9800 1690 9810 1730
rect 9850 1690 9860 1730
rect 9800 1670 9860 1690
rect 9910 1830 9970 1850
rect 9910 1790 9920 1830
rect 9960 1790 9970 1830
rect 9910 1730 9970 1790
rect 9910 1690 9920 1730
rect 9960 1690 9970 1730
rect 9150 1630 9190 1670
rect 9370 1630 9410 1670
rect 9590 1630 9630 1670
rect 9810 1630 9850 1670
rect 9030 1570 9040 1610
rect 9080 1570 9090 1610
rect 9030 1550 9090 1570
rect 9130 1610 9210 1630
rect 9130 1570 9150 1610
rect 9190 1570 9210 1610
rect 9130 1550 9210 1570
rect 9350 1610 9430 1630
rect 9350 1570 9370 1610
rect 9410 1570 9430 1610
rect 9350 1550 9430 1570
rect 9570 1610 9650 1630
rect 9570 1570 9590 1610
rect 9630 1570 9650 1610
rect 9570 1550 9650 1570
rect 9790 1610 9870 1630
rect 9790 1570 9810 1610
rect 9850 1570 9870 1610
rect 9790 1550 9870 1570
rect 9910 1610 9970 1690
rect 9910 1570 9920 1610
rect 9960 1570 9970 1610
rect 9910 1550 9970 1570
rect 10040 1840 10080 2010
rect 36600 1860 36680 1880
rect 36600 1840 36620 1860
rect 36660 1840 36680 1860
rect 38680 1860 38760 1880
rect 38680 1840 38700 1860
rect 9040 1510 9080 1550
rect 9920 1510 9960 1550
rect 10040 1510 10080 1680
rect 8920 1470 10080 1510
rect 35300 1800 36560 1840
rect 36720 1800 37980 1840
rect 35300 1630 35340 1800
rect 35520 1740 35600 1760
rect 35520 1700 35540 1740
rect 35580 1700 35600 1740
rect 35520 1680 35600 1700
rect 35650 1740 35710 1760
rect 35650 1700 35660 1740
rect 35700 1700 35710 1740
rect 35650 1680 35710 1700
rect 35890 1740 35950 1760
rect 35890 1700 35900 1740
rect 35940 1700 35950 1740
rect 35890 1680 35950 1700
rect 36130 1740 36190 1760
rect 36130 1700 36140 1740
rect 36180 1700 36190 1740
rect 36130 1680 36190 1700
rect 36240 1740 36320 1760
rect 36240 1700 36260 1740
rect 36300 1700 36320 1740
rect 36240 1680 36320 1700
rect 36370 1740 36430 1760
rect 36370 1700 36380 1740
rect 36420 1700 36430 1740
rect 36370 1680 36430 1700
rect 36610 1740 36670 1760
rect 36610 1700 36620 1740
rect 36660 1700 36670 1740
rect 36610 1680 36670 1700
rect 36850 1740 36910 1760
rect 36850 1700 36860 1740
rect 36900 1700 36910 1740
rect 36850 1680 36910 1700
rect 36960 1740 37040 1760
rect 36960 1700 36980 1740
rect 37020 1700 37040 1740
rect 36960 1680 37040 1700
rect 37090 1740 37150 1760
rect 37090 1700 37100 1740
rect 37140 1700 37150 1740
rect 37090 1680 37150 1700
rect 37330 1740 37390 1760
rect 37330 1700 37340 1740
rect 37380 1700 37390 1740
rect 37330 1680 37390 1700
rect 37570 1740 37630 1760
rect 37570 1700 37580 1740
rect 37620 1700 37630 1740
rect 37570 1680 37630 1700
rect 37680 1740 37760 1760
rect 37680 1700 37700 1740
rect 37740 1700 37760 1740
rect 37680 1680 37760 1700
rect 35540 1640 35580 1680
rect 35660 1640 35700 1680
rect 35900 1640 35940 1680
rect 36140 1640 36180 1680
rect 36260 1640 36300 1680
rect 36380 1640 36420 1680
rect 36620 1640 36660 1680
rect 36860 1640 36900 1680
rect 36980 1640 37020 1680
rect 37100 1640 37140 1680
rect 37340 1640 37380 1680
rect 37580 1640 37620 1680
rect 37700 1640 37740 1680
rect 35300 1300 35340 1470
rect 35410 1620 35470 1640
rect 35410 1580 35420 1620
rect 35460 1580 35470 1620
rect 35410 1520 35470 1580
rect 35410 1480 35420 1520
rect 35460 1480 35470 1520
rect 35410 1400 35470 1480
rect 35530 1620 35590 1640
rect 35530 1580 35540 1620
rect 35580 1580 35590 1620
rect 35530 1520 35590 1580
rect 35530 1480 35540 1520
rect 35580 1480 35590 1520
rect 35530 1460 35590 1480
rect 35650 1620 35710 1640
rect 35650 1580 35660 1620
rect 35700 1580 35710 1620
rect 35650 1520 35710 1580
rect 35650 1480 35660 1520
rect 35700 1480 35710 1520
rect 35650 1460 35710 1480
rect 35770 1620 35830 1640
rect 35770 1580 35780 1620
rect 35820 1580 35830 1620
rect 35770 1520 35830 1580
rect 35770 1480 35780 1520
rect 35820 1480 35830 1520
rect 35770 1460 35830 1480
rect 35890 1620 35950 1640
rect 35890 1580 35900 1620
rect 35940 1580 35950 1620
rect 35890 1520 35950 1580
rect 35890 1480 35900 1520
rect 35940 1480 35950 1520
rect 35890 1460 35950 1480
rect 36010 1620 36070 1640
rect 36010 1580 36020 1620
rect 36060 1580 36070 1620
rect 36010 1520 36070 1580
rect 36010 1480 36020 1520
rect 36060 1480 36070 1520
rect 36010 1460 36070 1480
rect 36130 1620 36190 1640
rect 36130 1580 36140 1620
rect 36180 1580 36190 1620
rect 36130 1520 36190 1580
rect 36130 1480 36140 1520
rect 36180 1480 36190 1520
rect 36130 1460 36190 1480
rect 36250 1620 36310 1640
rect 36250 1580 36260 1620
rect 36300 1580 36310 1620
rect 36250 1520 36310 1580
rect 36250 1480 36260 1520
rect 36300 1480 36310 1520
rect 36250 1460 36310 1480
rect 36370 1620 36430 1640
rect 36370 1580 36380 1620
rect 36420 1580 36430 1620
rect 36370 1520 36430 1580
rect 36370 1480 36380 1520
rect 36420 1480 36430 1520
rect 36370 1460 36430 1480
rect 36490 1620 36550 1640
rect 36490 1580 36500 1620
rect 36540 1580 36550 1620
rect 36490 1520 36550 1580
rect 36490 1480 36500 1520
rect 36540 1480 36550 1520
rect 36490 1460 36550 1480
rect 36610 1620 36670 1640
rect 36610 1580 36620 1620
rect 36660 1580 36670 1620
rect 36610 1520 36670 1580
rect 36610 1480 36620 1520
rect 36660 1480 36670 1520
rect 36610 1460 36670 1480
rect 36730 1620 36790 1640
rect 36730 1580 36740 1620
rect 36780 1580 36790 1620
rect 36730 1520 36790 1580
rect 36730 1480 36740 1520
rect 36780 1480 36790 1520
rect 36730 1460 36790 1480
rect 36850 1620 36910 1640
rect 36850 1580 36860 1620
rect 36900 1580 36910 1620
rect 36850 1520 36910 1580
rect 36850 1480 36860 1520
rect 36900 1480 36910 1520
rect 36850 1460 36910 1480
rect 36970 1620 37030 1640
rect 36970 1580 36980 1620
rect 37020 1580 37030 1620
rect 36970 1520 37030 1580
rect 36970 1480 36980 1520
rect 37020 1480 37030 1520
rect 36970 1460 37030 1480
rect 37090 1620 37150 1640
rect 37090 1580 37100 1620
rect 37140 1580 37150 1620
rect 37090 1520 37150 1580
rect 37090 1480 37100 1520
rect 37140 1480 37150 1520
rect 37090 1460 37150 1480
rect 37210 1620 37270 1640
rect 37210 1580 37220 1620
rect 37260 1580 37270 1620
rect 37210 1520 37270 1580
rect 37210 1480 37220 1520
rect 37260 1480 37270 1520
rect 37210 1460 37270 1480
rect 37330 1620 37390 1640
rect 37330 1580 37340 1620
rect 37380 1580 37390 1620
rect 37330 1520 37390 1580
rect 37330 1480 37340 1520
rect 37380 1480 37390 1520
rect 37330 1460 37390 1480
rect 37450 1620 37510 1640
rect 37450 1580 37460 1620
rect 37500 1580 37510 1620
rect 37450 1520 37510 1580
rect 37450 1480 37460 1520
rect 37500 1480 37510 1520
rect 37450 1460 37510 1480
rect 37570 1620 37630 1640
rect 37570 1580 37580 1620
rect 37620 1580 37630 1620
rect 37570 1520 37630 1580
rect 37570 1480 37580 1520
rect 37620 1480 37630 1520
rect 37570 1460 37630 1480
rect 37690 1620 37750 1640
rect 37690 1580 37700 1620
rect 37740 1580 37750 1620
rect 37690 1520 37750 1580
rect 37690 1480 37700 1520
rect 37740 1480 37750 1520
rect 37690 1460 37750 1480
rect 37810 1620 37870 1640
rect 37810 1580 37820 1620
rect 37860 1580 37870 1620
rect 37810 1520 37870 1580
rect 37810 1480 37820 1520
rect 37860 1480 37870 1520
rect 35780 1420 35820 1460
rect 36020 1420 36060 1460
rect 36500 1420 36540 1460
rect 36740 1420 36780 1460
rect 37220 1420 37260 1460
rect 37460 1420 37500 1460
rect 35410 1360 35420 1400
rect 35460 1360 35470 1400
rect 35410 1340 35470 1360
rect 35580 1400 35660 1420
rect 35580 1360 35600 1400
rect 35640 1360 35660 1400
rect 35580 1340 35660 1360
rect 35760 1400 35840 1420
rect 35760 1360 35780 1400
rect 35820 1360 35840 1400
rect 35760 1340 35840 1360
rect 36000 1400 36080 1420
rect 36000 1360 36020 1400
rect 36060 1360 36080 1400
rect 36000 1340 36080 1360
rect 36240 1400 36320 1420
rect 36240 1360 36260 1400
rect 36300 1360 36320 1400
rect 36240 1340 36320 1360
rect 36480 1400 36560 1420
rect 36480 1360 36500 1400
rect 36540 1360 36560 1400
rect 36480 1340 36560 1360
rect 36720 1400 36800 1420
rect 36720 1360 36740 1400
rect 36780 1360 36800 1400
rect 36720 1340 36800 1360
rect 36960 1400 37040 1420
rect 36960 1360 36980 1400
rect 37020 1360 37040 1400
rect 36960 1340 37040 1360
rect 37200 1400 37280 1420
rect 37200 1360 37220 1400
rect 37260 1360 37280 1400
rect 37200 1340 37280 1360
rect 37440 1400 37520 1420
rect 37440 1360 37460 1400
rect 37500 1360 37520 1400
rect 37440 1340 37520 1360
rect 37630 1400 37690 1420
rect 37630 1360 37640 1400
rect 37680 1360 37690 1400
rect 37630 1340 37690 1360
rect 37810 1400 37870 1480
rect 37810 1360 37820 1400
rect 37860 1360 37870 1400
rect 37810 1340 37870 1360
rect 37940 1630 37980 1800
rect 35420 1300 35460 1340
rect 37820 1300 37860 1340
rect 37940 1300 37980 1470
rect 35300 1260 36560 1300
rect 36720 1260 37980 1300
rect 38340 1820 38700 1840
rect 38740 1840 38760 1860
rect 38920 1860 39000 1880
rect 38920 1840 38940 1860
rect 38740 1820 38940 1840
rect 38980 1840 39000 1860
rect 39160 1860 39240 1880
rect 39160 1840 39180 1860
rect 38980 1820 39180 1840
rect 39220 1840 39240 1860
rect 39400 1860 39480 1880
rect 39400 1840 39420 1860
rect 39220 1820 39420 1840
rect 39460 1840 39480 1860
rect 39640 1860 39720 1880
rect 39640 1840 39660 1860
rect 39700 1840 39720 1860
rect 39880 1860 39960 1880
rect 39880 1840 39900 1860
rect 39460 1820 39600 1840
rect 39760 1820 39900 1840
rect 39940 1840 39960 1860
rect 40120 1860 40200 1880
rect 40120 1840 40140 1860
rect 39940 1820 40140 1840
rect 40180 1840 40200 1860
rect 40360 1860 40440 1880
rect 40360 1840 40380 1860
rect 40180 1820 40380 1840
rect 40420 1840 40440 1860
rect 40600 1860 40680 1880
rect 40600 1840 40620 1860
rect 40420 1820 40620 1840
rect 40660 1840 40680 1860
rect 40660 1820 41020 1840
rect 38340 1800 39600 1820
rect 39760 1800 41020 1820
rect 38340 1630 38380 1800
rect 38560 1740 38640 1760
rect 38560 1700 38580 1740
rect 38620 1700 38640 1740
rect 38560 1680 38640 1700
rect 38690 1740 38750 1760
rect 38690 1700 38700 1740
rect 38740 1700 38750 1740
rect 38690 1680 38750 1700
rect 38930 1740 38990 1760
rect 38930 1700 38940 1740
rect 38980 1700 38990 1740
rect 38930 1680 38990 1700
rect 39170 1740 39230 1760
rect 39170 1700 39180 1740
rect 39220 1700 39230 1740
rect 39170 1680 39230 1700
rect 39280 1740 39360 1760
rect 39280 1700 39300 1740
rect 39340 1700 39360 1740
rect 39280 1680 39360 1700
rect 39410 1740 39470 1760
rect 39410 1700 39420 1740
rect 39460 1700 39470 1740
rect 39410 1680 39470 1700
rect 39650 1740 39710 1760
rect 39650 1700 39660 1740
rect 39700 1700 39710 1740
rect 39650 1680 39710 1700
rect 39890 1740 39950 1760
rect 39890 1700 39900 1740
rect 39940 1700 39950 1740
rect 39890 1680 39950 1700
rect 40000 1740 40080 1760
rect 40000 1700 40020 1740
rect 40060 1700 40080 1740
rect 40000 1680 40080 1700
rect 40130 1740 40190 1760
rect 40130 1700 40140 1740
rect 40180 1700 40190 1740
rect 40130 1680 40190 1700
rect 40370 1740 40430 1760
rect 40370 1700 40380 1740
rect 40420 1700 40430 1740
rect 40370 1680 40430 1700
rect 40610 1740 40670 1760
rect 40610 1700 40620 1740
rect 40660 1700 40670 1740
rect 40610 1680 40670 1700
rect 40720 1740 40800 1760
rect 40720 1700 40740 1740
rect 40780 1700 40800 1740
rect 40720 1680 40800 1700
rect 38580 1640 38620 1680
rect 38700 1640 38740 1680
rect 38940 1640 38980 1680
rect 39180 1640 39220 1680
rect 39300 1640 39340 1680
rect 39420 1640 39460 1680
rect 39660 1640 39700 1680
rect 39900 1640 39940 1680
rect 40020 1640 40060 1680
rect 40140 1640 40180 1680
rect 40380 1640 40420 1680
rect 40620 1640 40660 1680
rect 40740 1640 40780 1680
rect 38340 1300 38380 1470
rect 38450 1620 38510 1640
rect 38450 1580 38460 1620
rect 38500 1580 38510 1620
rect 38450 1520 38510 1580
rect 38450 1480 38460 1520
rect 38500 1480 38510 1520
rect 38450 1400 38510 1480
rect 38570 1620 38630 1640
rect 38570 1580 38580 1620
rect 38620 1580 38630 1620
rect 38570 1520 38630 1580
rect 38570 1480 38580 1520
rect 38620 1480 38630 1520
rect 38570 1460 38630 1480
rect 38690 1620 38750 1640
rect 38690 1580 38700 1620
rect 38740 1580 38750 1620
rect 38690 1520 38750 1580
rect 38690 1480 38700 1520
rect 38740 1480 38750 1520
rect 38690 1460 38750 1480
rect 38810 1620 38870 1640
rect 38810 1580 38820 1620
rect 38860 1580 38870 1620
rect 38810 1520 38870 1580
rect 38810 1480 38820 1520
rect 38860 1480 38870 1520
rect 38810 1460 38870 1480
rect 38930 1620 38990 1640
rect 38930 1580 38940 1620
rect 38980 1580 38990 1620
rect 38930 1520 38990 1580
rect 38930 1480 38940 1520
rect 38980 1480 38990 1520
rect 38930 1460 38990 1480
rect 39050 1620 39110 1640
rect 39050 1580 39060 1620
rect 39100 1580 39110 1620
rect 39050 1520 39110 1580
rect 39050 1480 39060 1520
rect 39100 1480 39110 1520
rect 39050 1460 39110 1480
rect 39170 1620 39230 1640
rect 39170 1580 39180 1620
rect 39220 1580 39230 1620
rect 39170 1520 39230 1580
rect 39170 1480 39180 1520
rect 39220 1480 39230 1520
rect 39170 1460 39230 1480
rect 39290 1620 39350 1640
rect 39290 1580 39300 1620
rect 39340 1580 39350 1620
rect 39290 1520 39350 1580
rect 39290 1480 39300 1520
rect 39340 1480 39350 1520
rect 39290 1460 39350 1480
rect 39410 1620 39470 1640
rect 39410 1580 39420 1620
rect 39460 1580 39470 1620
rect 39410 1520 39470 1580
rect 39410 1480 39420 1520
rect 39460 1480 39470 1520
rect 39410 1460 39470 1480
rect 39530 1620 39590 1640
rect 39530 1580 39540 1620
rect 39580 1580 39590 1620
rect 39530 1520 39590 1580
rect 39530 1480 39540 1520
rect 39580 1480 39590 1520
rect 39530 1460 39590 1480
rect 39650 1620 39710 1640
rect 39650 1580 39660 1620
rect 39700 1580 39710 1620
rect 39650 1520 39710 1580
rect 39650 1480 39660 1520
rect 39700 1480 39710 1520
rect 39650 1460 39710 1480
rect 39770 1620 39830 1640
rect 39770 1580 39780 1620
rect 39820 1580 39830 1620
rect 39770 1520 39830 1580
rect 39770 1480 39780 1520
rect 39820 1480 39830 1520
rect 39770 1460 39830 1480
rect 39890 1620 39950 1640
rect 39890 1580 39900 1620
rect 39940 1580 39950 1620
rect 39890 1520 39950 1580
rect 39890 1480 39900 1520
rect 39940 1480 39950 1520
rect 39890 1460 39950 1480
rect 40010 1620 40070 1640
rect 40010 1580 40020 1620
rect 40060 1580 40070 1620
rect 40010 1520 40070 1580
rect 40010 1480 40020 1520
rect 40060 1480 40070 1520
rect 40010 1460 40070 1480
rect 40130 1620 40190 1640
rect 40130 1580 40140 1620
rect 40180 1580 40190 1620
rect 40130 1520 40190 1580
rect 40130 1480 40140 1520
rect 40180 1480 40190 1520
rect 40130 1460 40190 1480
rect 40250 1620 40310 1640
rect 40250 1580 40260 1620
rect 40300 1580 40310 1620
rect 40250 1520 40310 1580
rect 40250 1480 40260 1520
rect 40300 1480 40310 1520
rect 40250 1460 40310 1480
rect 40370 1620 40430 1640
rect 40370 1580 40380 1620
rect 40420 1580 40430 1620
rect 40370 1520 40430 1580
rect 40370 1480 40380 1520
rect 40420 1480 40430 1520
rect 40370 1460 40430 1480
rect 40490 1620 40550 1640
rect 40490 1580 40500 1620
rect 40540 1580 40550 1620
rect 40490 1520 40550 1580
rect 40490 1480 40500 1520
rect 40540 1480 40550 1520
rect 40490 1460 40550 1480
rect 40610 1620 40670 1640
rect 40610 1580 40620 1620
rect 40660 1580 40670 1620
rect 40610 1520 40670 1580
rect 40610 1480 40620 1520
rect 40660 1480 40670 1520
rect 40610 1460 40670 1480
rect 40730 1620 40790 1640
rect 40730 1580 40740 1620
rect 40780 1580 40790 1620
rect 40730 1520 40790 1580
rect 40730 1480 40740 1520
rect 40780 1480 40790 1520
rect 40730 1460 40790 1480
rect 40850 1620 40910 1640
rect 40850 1580 40860 1620
rect 40900 1580 40910 1620
rect 40850 1520 40910 1580
rect 40850 1480 40860 1520
rect 40900 1480 40910 1520
rect 38820 1420 38860 1460
rect 39060 1420 39100 1460
rect 39540 1420 39580 1460
rect 39780 1420 39820 1460
rect 40260 1420 40300 1460
rect 40500 1420 40540 1460
rect 38450 1360 38460 1400
rect 38500 1360 38510 1400
rect 38450 1340 38510 1360
rect 38630 1400 38690 1420
rect 38630 1360 38640 1400
rect 38680 1360 38690 1400
rect 38630 1340 38690 1360
rect 38800 1400 38880 1420
rect 38800 1360 38820 1400
rect 38860 1360 38880 1400
rect 38800 1340 38880 1360
rect 39040 1400 39120 1420
rect 39040 1360 39060 1400
rect 39100 1360 39120 1400
rect 39040 1340 39120 1360
rect 39280 1400 39360 1420
rect 39280 1360 39300 1400
rect 39340 1360 39360 1400
rect 39280 1340 39360 1360
rect 39520 1400 39600 1420
rect 39520 1360 39540 1400
rect 39580 1360 39600 1400
rect 39520 1340 39600 1360
rect 39760 1400 39840 1420
rect 39760 1360 39780 1400
rect 39820 1360 39840 1400
rect 39760 1340 39840 1360
rect 40000 1400 40080 1420
rect 40000 1360 40020 1400
rect 40060 1360 40080 1400
rect 40000 1340 40080 1360
rect 40240 1400 40320 1420
rect 40240 1360 40260 1400
rect 40300 1360 40320 1400
rect 40240 1340 40320 1360
rect 40480 1400 40560 1420
rect 40480 1360 40500 1400
rect 40540 1360 40560 1400
rect 40480 1340 40560 1360
rect 40660 1400 40740 1420
rect 40660 1360 40680 1400
rect 40720 1360 40740 1400
rect 40660 1340 40740 1360
rect 40850 1400 40910 1480
rect 40850 1360 40860 1400
rect 40900 1360 40910 1400
rect 40850 1340 40910 1360
rect 40980 1630 41020 1800
rect 38460 1300 38500 1340
rect 40860 1300 40900 1340
rect 40980 1300 41020 1470
rect 38340 1260 39600 1300
rect 39760 1260 41020 1300
rect 36160 1140 36820 1180
rect 36980 1140 37640 1180
rect 36160 930 36200 1140
rect 36380 1080 36460 1100
rect 36380 1040 36400 1080
rect 36440 1040 36460 1080
rect 36380 1020 36460 1040
rect 36260 990 36340 1010
rect 36260 950 36280 990
rect 36320 950 36340 990
rect 36260 930 36340 950
rect 36510 990 36570 1010
rect 36510 950 36520 990
rect 36560 950 36570 990
rect 36510 930 36570 950
rect 36740 990 36820 1010
rect 36740 950 36760 990
rect 36800 950 36820 990
rect 36740 930 36820 950
rect 36990 990 37050 1010
rect 36990 950 37000 990
rect 37040 950 37050 990
rect 36990 930 37050 950
rect 37220 990 37300 1010
rect 37220 950 37240 990
rect 37280 950 37300 990
rect 37220 930 37300 950
rect 37470 990 37530 1010
rect 37470 950 37480 990
rect 37520 950 37530 990
rect 37470 930 37530 950
rect 37600 930 37640 1140
rect 36280 890 36320 930
rect 36520 890 36560 930
rect 36760 890 36800 930
rect 37000 890 37040 930
rect 37240 890 37280 930
rect 37480 890 37520 930
rect 36270 870 36330 890
rect 36270 830 36280 870
rect 36320 830 36330 870
rect 36270 810 36330 830
rect 36390 870 36450 890
rect 36390 830 36400 870
rect 36440 830 36450 870
rect 36390 810 36450 830
rect 36510 870 36570 890
rect 36510 830 36520 870
rect 36560 830 36570 870
rect 36510 810 36570 830
rect 36630 870 36690 890
rect 36630 830 36640 870
rect 36680 830 36690 870
rect 36630 810 36690 830
rect 36750 870 36810 890
rect 36750 830 36760 870
rect 36800 830 36810 870
rect 36750 810 36810 830
rect 36870 870 36930 890
rect 36870 830 36880 870
rect 36920 830 36930 870
rect 36870 810 36930 830
rect 36990 870 37050 890
rect 36990 830 37000 870
rect 37040 830 37050 870
rect 36990 810 37050 830
rect 37110 870 37170 890
rect 37110 830 37120 870
rect 37160 830 37170 870
rect 37110 810 37170 830
rect 37230 870 37290 890
rect 37230 830 37240 870
rect 37280 830 37290 870
rect 37230 810 37290 830
rect 37350 870 37410 890
rect 37350 830 37360 870
rect 37400 830 37410 870
rect 37350 810 37410 830
rect 37470 870 37530 890
rect 37470 830 37480 870
rect 37520 830 37530 870
rect 37470 810 37530 830
rect 37580 810 37600 890
rect 38680 1140 39340 1180
rect 39500 1140 40160 1180
rect 38680 930 38720 1140
rect 39860 1080 39940 1100
rect 39860 1040 39880 1080
rect 39920 1040 39940 1080
rect 39860 1020 39940 1040
rect 38790 990 38850 1010
rect 38790 950 38800 990
rect 38840 950 38850 990
rect 38790 930 38850 950
rect 39020 990 39100 1010
rect 39020 950 39040 990
rect 39080 950 39100 990
rect 39020 930 39100 950
rect 39270 990 39330 1010
rect 39270 950 39280 990
rect 39320 950 39330 990
rect 39270 930 39330 950
rect 39500 990 39580 1010
rect 39500 950 39520 990
rect 39560 950 39580 990
rect 39500 930 39580 950
rect 39750 990 39810 1010
rect 39750 950 39760 990
rect 39800 950 39810 990
rect 39750 930 39810 950
rect 39980 990 40060 1010
rect 39980 950 40000 990
rect 40040 950 40060 990
rect 39980 930 40060 950
rect 40120 930 40160 1140
rect 36400 770 36440 810
rect 36640 770 36680 810
rect 36880 770 36920 810
rect 37120 770 37160 810
rect 37360 770 37400 810
rect 37640 810 37660 890
rect 38660 810 38680 890
rect 38800 890 38840 930
rect 39040 890 39080 930
rect 39280 890 39320 930
rect 39520 890 39560 930
rect 39760 890 39800 930
rect 40000 890 40040 930
rect 36160 650 36200 770
rect 36260 750 36340 770
rect 36260 710 36280 750
rect 36320 710 36340 750
rect 36260 690 36340 710
rect 36390 750 36450 770
rect 36390 710 36400 750
rect 36440 710 36450 750
rect 36390 690 36450 710
rect 36630 750 36690 770
rect 36630 710 36640 750
rect 36680 710 36690 750
rect 36630 690 36690 710
rect 36870 750 36930 770
rect 36870 710 36880 750
rect 36920 710 36930 750
rect 36870 690 36930 710
rect 37110 750 37170 770
rect 37110 710 37120 750
rect 37160 710 37170 750
rect 37110 690 37170 710
rect 37350 750 37410 770
rect 37350 710 37360 750
rect 37400 710 37410 750
rect 37350 690 37410 710
rect 37600 650 37640 770
rect 36160 610 36820 650
rect 36980 610 37640 650
rect 38720 810 38740 890
rect 38790 870 38850 890
rect 38790 830 38800 870
rect 38840 830 38850 870
rect 38790 810 38850 830
rect 38910 870 38970 890
rect 38910 830 38920 870
rect 38960 830 38970 870
rect 38910 810 38970 830
rect 39030 870 39090 890
rect 39030 830 39040 870
rect 39080 830 39090 870
rect 39030 810 39090 830
rect 39150 870 39210 890
rect 39150 830 39160 870
rect 39200 830 39210 870
rect 39150 810 39210 830
rect 39270 870 39330 890
rect 39270 830 39280 870
rect 39320 830 39330 870
rect 39270 810 39330 830
rect 39390 870 39450 890
rect 39390 830 39400 870
rect 39440 830 39450 870
rect 39390 810 39450 830
rect 39510 870 39570 890
rect 39510 830 39520 870
rect 39560 830 39570 870
rect 39510 810 39570 830
rect 39630 870 39690 890
rect 39630 830 39640 870
rect 39680 830 39690 870
rect 39630 810 39690 830
rect 39750 870 39810 890
rect 39750 830 39760 870
rect 39800 830 39810 870
rect 39750 810 39810 830
rect 39870 870 39930 890
rect 39870 830 39880 870
rect 39920 830 39930 870
rect 39870 810 39930 830
rect 39990 870 40050 890
rect 39990 830 40000 870
rect 40040 830 40050 870
rect 39990 810 40050 830
rect 38920 770 38960 810
rect 39160 770 39200 810
rect 39400 770 39440 810
rect 39640 770 39680 810
rect 39880 770 39920 810
rect 38680 650 38720 770
rect 38910 750 38970 770
rect 38910 710 38920 750
rect 38960 710 38970 750
rect 38910 690 38970 710
rect 39150 750 39210 770
rect 39150 710 39160 750
rect 39200 710 39210 750
rect 39150 690 39210 710
rect 39390 750 39450 770
rect 39390 710 39400 750
rect 39440 710 39450 750
rect 39390 690 39450 710
rect 39630 750 39690 770
rect 39630 710 39640 750
rect 39680 710 39690 750
rect 39630 690 39690 710
rect 39870 750 39930 770
rect 39870 710 39880 750
rect 39920 710 39930 750
rect 39870 690 39930 710
rect 39980 750 40060 770
rect 39980 710 40000 750
rect 40040 710 40060 750
rect 39980 690 40060 710
rect 40120 650 40160 770
rect 38680 610 40160 650
rect 39860 570 39940 610
rect 35680 490 36820 530
rect 36980 490 38120 530
rect 35680 180 35720 490
rect 35960 430 36040 450
rect 35780 400 35860 420
rect 35780 360 35800 400
rect 35840 360 35860 400
rect 35960 390 35980 430
rect 36020 390 36040 430
rect 35960 370 36040 390
rect 36200 430 36280 450
rect 36200 390 36220 430
rect 36260 390 36280 430
rect 36200 370 36280 390
rect 36440 430 36520 450
rect 36440 390 36460 430
rect 36500 390 36520 430
rect 36440 370 36520 390
rect 36680 430 36760 450
rect 36680 390 36700 430
rect 36740 390 36760 430
rect 36680 370 36760 390
rect 37160 430 37240 450
rect 37160 390 37180 430
rect 37220 390 37240 430
rect 37160 370 37240 390
rect 37400 430 37480 450
rect 37400 390 37420 430
rect 37460 390 37480 430
rect 37400 370 37480 390
rect 37640 430 37720 450
rect 37640 390 37660 430
rect 37700 390 37720 430
rect 37640 370 37720 390
rect 37940 400 38020 420
rect 35780 340 35860 360
rect 37940 360 37960 400
rect 38000 360 38020 400
rect 37940 340 38020 360
rect 35680 -300 35720 20
rect 35790 320 35850 340
rect 35790 280 35800 320
rect 35840 280 35850 320
rect 35790 220 35850 280
rect 35790 180 35800 220
rect 35840 180 35850 220
rect 35790 120 35850 180
rect 35790 80 35800 120
rect 35840 80 35850 120
rect 35790 20 35850 80
rect 35790 -20 35800 20
rect 35840 -20 35850 20
rect 35790 -80 35850 -20
rect 35790 -120 35800 -80
rect 35840 -120 35850 -80
rect 35790 -140 35850 -120
rect 36870 320 36930 340
rect 36870 280 36880 320
rect 36920 280 36930 320
rect 36870 220 36930 280
rect 36870 180 36880 220
rect 36920 180 36930 220
rect 36870 120 36930 180
rect 36870 80 36880 120
rect 36920 80 36930 120
rect 36870 20 36930 80
rect 36870 -20 36880 20
rect 36920 -20 36930 20
rect 36870 -80 36930 -20
rect 36870 -120 36880 -80
rect 36920 -120 36930 -80
rect 36870 -140 36930 -120
rect 37950 320 38010 340
rect 37950 280 37960 320
rect 38000 280 38010 320
rect 37950 220 38010 280
rect 37950 180 37960 220
rect 38000 180 38010 220
rect 37950 120 38010 180
rect 37950 80 37960 120
rect 38000 80 38010 120
rect 37950 20 38010 80
rect 37950 -20 37960 20
rect 38000 -20 38010 20
rect 37950 -80 38010 -20
rect 37950 -120 37960 -80
rect 38000 -120 38010 -80
rect 37950 -140 38010 -120
rect 38080 180 38120 490
rect 36880 -180 36920 -140
rect 36860 -200 36940 -180
rect 36860 -240 36880 -200
rect 36920 -240 36940 -200
rect 36860 -260 36940 -240
rect 36880 -300 36920 -260
rect 38080 -300 38120 20
rect 35680 -340 36820 -300
rect 36980 -340 38120 -300
rect 38200 490 39340 530
rect 39500 490 40640 530
rect 38200 180 38240 490
rect 38600 430 38680 450
rect 38300 400 38380 420
rect 38300 360 38320 400
rect 38360 360 38380 400
rect 38600 390 38620 430
rect 38660 390 38680 430
rect 38600 370 38680 390
rect 38840 430 38920 450
rect 38840 390 38860 430
rect 38900 390 38920 430
rect 38840 370 38920 390
rect 39080 430 39160 450
rect 39080 390 39100 430
rect 39140 390 39160 430
rect 39080 370 39160 390
rect 39560 430 39640 450
rect 39560 390 39580 430
rect 39620 390 39640 430
rect 39560 370 39640 390
rect 39800 430 39880 450
rect 39800 390 39820 430
rect 39860 390 39880 430
rect 39800 370 39880 390
rect 40040 430 40120 450
rect 40040 390 40060 430
rect 40100 390 40120 430
rect 40040 370 40120 390
rect 40280 430 40360 450
rect 40280 390 40300 430
rect 40340 390 40360 430
rect 40280 370 40360 390
rect 40460 400 40540 420
rect 38300 340 38380 360
rect 40460 360 40480 400
rect 40520 360 40540 400
rect 40460 340 40540 360
rect 38200 -300 38240 20
rect 38310 320 38370 340
rect 38310 280 38320 320
rect 38360 280 38370 320
rect 38310 220 38370 280
rect 38310 180 38320 220
rect 38360 180 38370 220
rect 38310 120 38370 180
rect 38310 80 38320 120
rect 38360 80 38370 120
rect 38310 20 38370 80
rect 38310 -20 38320 20
rect 38360 -20 38370 20
rect 38310 -80 38370 -20
rect 38310 -120 38320 -80
rect 38360 -120 38370 -80
rect 38310 -140 38370 -120
rect 39390 320 39450 340
rect 39390 280 39400 320
rect 39440 280 39450 320
rect 39390 220 39450 280
rect 39390 180 39400 220
rect 39440 180 39450 220
rect 39390 120 39450 180
rect 39390 80 39400 120
rect 39440 80 39450 120
rect 39390 20 39450 80
rect 39390 -20 39400 20
rect 39440 -20 39450 20
rect 39390 -80 39450 -20
rect 39390 -120 39400 -80
rect 39440 -120 39450 -80
rect 39390 -140 39450 -120
rect 40470 320 40530 340
rect 40470 280 40480 320
rect 40520 280 40530 320
rect 40470 220 40530 280
rect 40470 180 40480 220
rect 40520 180 40530 220
rect 40470 120 40530 180
rect 40470 80 40480 120
rect 40520 80 40530 120
rect 40470 20 40530 80
rect 40470 -20 40480 20
rect 40520 -20 40530 20
rect 40470 -80 40530 -20
rect 40470 -120 40480 -80
rect 40520 -120 40530 -80
rect 40470 -140 40530 -120
rect 40600 180 40640 490
rect 39400 -180 39440 -140
rect 39380 -200 39460 -180
rect 39380 -240 39400 -200
rect 39440 -240 39460 -200
rect 39380 -260 39460 -240
rect 39400 -300 39440 -260
rect 40600 -300 40640 20
rect 38200 -340 39340 -300
rect 39500 -340 40640 -300
rect 35880 -440 38080 -400
rect 38240 -440 40430 -400
rect 35880 -610 35920 -440
rect 36040 -500 36120 -480
rect 36040 -540 36060 -500
rect 36100 -540 36120 -500
rect 36040 -560 36120 -540
rect 36200 -500 36280 -480
rect 36200 -540 36220 -500
rect 36260 -540 36280 -500
rect 36200 -560 36280 -540
rect 36360 -500 36440 -480
rect 36360 -540 36380 -500
rect 36420 -540 36440 -500
rect 36360 -560 36440 -540
rect 36520 -500 36600 -480
rect 36520 -540 36540 -500
rect 36580 -540 36600 -500
rect 36520 -560 36600 -540
rect 36680 -500 36760 -480
rect 36680 -540 36700 -500
rect 36740 -540 36760 -500
rect 36680 -560 36760 -540
rect 36840 -500 36920 -480
rect 36840 -540 36860 -500
rect 36900 -540 36920 -500
rect 36840 -560 36920 -540
rect 37000 -500 37080 -480
rect 37000 -540 37020 -500
rect 37060 -540 37080 -500
rect 37000 -560 37080 -540
rect 37160 -500 37240 -480
rect 37160 -540 37180 -500
rect 37220 -540 37240 -500
rect 37160 -560 37240 -540
rect 37320 -500 37400 -480
rect 37320 -540 37340 -500
rect 37380 -540 37400 -500
rect 37320 -560 37400 -540
rect 37480 -500 37560 -480
rect 37480 -540 37500 -500
rect 37540 -540 37560 -500
rect 37480 -560 37560 -540
rect 37640 -500 37720 -480
rect 37640 -540 37660 -500
rect 37700 -540 37720 -500
rect 37640 -560 37720 -540
rect 37800 -500 37880 -480
rect 37800 -540 37820 -500
rect 37860 -540 37880 -500
rect 37800 -560 37880 -540
rect 37960 -500 38040 -480
rect 37960 -540 37980 -500
rect 38020 -540 38040 -500
rect 37960 -560 38040 -540
rect 38120 -500 38200 -480
rect 38120 -540 38140 -500
rect 38180 -540 38200 -500
rect 38120 -560 38200 -540
rect 38280 -500 38360 -480
rect 38280 -540 38300 -500
rect 38340 -540 38360 -500
rect 38280 -560 38360 -540
rect 38440 -500 38520 -480
rect 38440 -540 38460 -500
rect 38500 -540 38520 -500
rect 38440 -560 38520 -540
rect 38600 -500 38680 -480
rect 38600 -540 38620 -500
rect 38660 -540 38680 -500
rect 38600 -560 38680 -540
rect 38760 -500 38840 -480
rect 38760 -540 38780 -500
rect 38820 -540 38840 -500
rect 38760 -560 38840 -540
rect 38920 -500 39000 -480
rect 38920 -540 38940 -500
rect 38980 -540 39000 -500
rect 38920 -560 39000 -540
rect 39080 -500 39160 -480
rect 39080 -540 39100 -500
rect 39140 -540 39160 -500
rect 39080 -560 39160 -540
rect 39240 -500 39320 -480
rect 39240 -540 39260 -500
rect 39300 -540 39320 -500
rect 39240 -560 39320 -540
rect 39400 -500 39480 -480
rect 39400 -540 39420 -500
rect 39460 -540 39480 -500
rect 39400 -560 39480 -540
rect 39560 -500 39640 -480
rect 39560 -540 39580 -500
rect 39620 -540 39640 -500
rect 39560 -560 39640 -540
rect 39720 -500 39800 -480
rect 39720 -540 39740 -500
rect 39780 -540 39800 -500
rect 39720 -560 39800 -540
rect 39880 -500 39960 -480
rect 39880 -540 39900 -500
rect 39940 -540 39960 -500
rect 39880 -560 39960 -540
rect 40040 -500 40120 -480
rect 40040 -540 40060 -500
rect 40100 -540 40120 -500
rect 40040 -560 40120 -540
rect 36060 -600 36100 -560
rect 38140 -600 38180 -560
rect 36050 -620 36110 -600
rect 36050 -650 36060 -620
rect 35960 -660 36060 -650
rect 36100 -660 36110 -620
rect 35960 -670 36110 -660
rect 35960 -710 35980 -670
rect 36020 -710 36110 -670
rect 35960 -720 36110 -710
rect 35960 -730 36060 -720
rect 35880 -850 35920 -770
rect 36050 -760 36060 -730
rect 36100 -760 36110 -720
rect 36050 -780 36110 -760
rect 38130 -620 38190 -600
rect 38130 -660 38140 -620
rect 38180 -660 38190 -620
rect 38130 -720 38190 -660
rect 38130 -760 38140 -720
rect 38180 -760 38190 -720
rect 38130 -780 38190 -760
rect 40210 -620 40270 -600
rect 40210 -660 40220 -620
rect 40260 -650 40270 -620
rect 40390 -610 40430 -440
rect 40260 -660 40350 -650
rect 40210 -670 40350 -660
rect 40210 -710 40290 -670
rect 40330 -710 40350 -670
rect 40210 -720 40350 -710
rect 40210 -760 40220 -720
rect 40260 -730 40350 -720
rect 40260 -760 40270 -730
rect 40210 -780 40270 -760
rect 40390 -850 40430 -770
rect 35880 -890 38080 -850
rect 38240 -890 40430 -850
rect 36240 -990 36800 -950
rect 36960 -990 37400 -950
rect 36240 -1160 36280 -990
rect 36560 -1050 36640 -1030
rect 36560 -1090 36580 -1050
rect 36620 -1090 36640 -1050
rect 36560 -1110 36640 -1090
rect 36780 -1050 36860 -1030
rect 36780 -1090 36800 -1050
rect 36840 -1090 36860 -1050
rect 36780 -1110 36860 -1090
rect 36900 -1050 36960 -1030
rect 36900 -1090 36910 -1050
rect 36950 -1090 36960 -1050
rect 36900 -1110 36960 -1090
rect 37000 -1050 37080 -1030
rect 37000 -1090 37020 -1050
rect 37060 -1090 37080 -1050
rect 37000 -1110 37080 -1090
rect 36580 -1150 36620 -1110
rect 36800 -1150 36840 -1110
rect 37020 -1150 37060 -1110
rect 36240 -1490 36280 -1320
rect 36350 -1170 36410 -1150
rect 36350 -1210 36360 -1170
rect 36400 -1210 36410 -1170
rect 36350 -1270 36410 -1210
rect 36350 -1310 36360 -1270
rect 36400 -1310 36410 -1270
rect 36350 -1390 36410 -1310
rect 36460 -1170 36520 -1150
rect 36460 -1210 36470 -1170
rect 36510 -1210 36520 -1170
rect 36460 -1270 36520 -1210
rect 36460 -1310 36470 -1270
rect 36510 -1310 36520 -1270
rect 36460 -1330 36520 -1310
rect 36570 -1170 36630 -1150
rect 36570 -1210 36580 -1170
rect 36620 -1210 36630 -1170
rect 36570 -1270 36630 -1210
rect 36570 -1310 36580 -1270
rect 36620 -1310 36630 -1270
rect 36570 -1330 36630 -1310
rect 36680 -1170 36740 -1150
rect 36680 -1210 36690 -1170
rect 36730 -1210 36740 -1170
rect 36680 -1270 36740 -1210
rect 36680 -1310 36690 -1270
rect 36730 -1310 36740 -1270
rect 36680 -1330 36740 -1310
rect 36790 -1170 36850 -1150
rect 36790 -1210 36800 -1170
rect 36840 -1210 36850 -1170
rect 36790 -1270 36850 -1210
rect 36790 -1310 36800 -1270
rect 36840 -1310 36850 -1270
rect 36790 -1330 36850 -1310
rect 36900 -1170 36960 -1150
rect 36900 -1210 36910 -1170
rect 36950 -1210 36960 -1170
rect 36900 -1270 36960 -1210
rect 36900 -1310 36910 -1270
rect 36950 -1310 36960 -1270
rect 36900 -1330 36960 -1310
rect 37010 -1170 37070 -1150
rect 37010 -1210 37020 -1170
rect 37060 -1210 37070 -1170
rect 37010 -1270 37070 -1210
rect 37010 -1310 37020 -1270
rect 37060 -1310 37070 -1270
rect 37010 -1330 37070 -1310
rect 37120 -1170 37180 -1150
rect 37120 -1210 37130 -1170
rect 37170 -1210 37180 -1170
rect 37120 -1270 37180 -1210
rect 37120 -1310 37130 -1270
rect 37170 -1310 37180 -1270
rect 37120 -1330 37180 -1310
rect 37230 -1170 37290 -1150
rect 37230 -1210 37240 -1170
rect 37280 -1210 37290 -1170
rect 37230 -1270 37290 -1210
rect 37230 -1310 37240 -1270
rect 37280 -1310 37290 -1270
rect 36470 -1370 36510 -1330
rect 36690 -1370 36730 -1330
rect 36910 -1370 36950 -1330
rect 37130 -1370 37170 -1330
rect 36350 -1430 36360 -1390
rect 36400 -1430 36410 -1390
rect 36350 -1450 36410 -1430
rect 36450 -1390 36530 -1370
rect 36450 -1430 36470 -1390
rect 36510 -1430 36530 -1390
rect 36450 -1450 36530 -1430
rect 36670 -1390 36750 -1370
rect 36670 -1430 36690 -1390
rect 36730 -1430 36750 -1390
rect 36670 -1450 36750 -1430
rect 36890 -1390 36970 -1370
rect 36890 -1430 36910 -1390
rect 36950 -1430 36970 -1390
rect 36890 -1450 36970 -1430
rect 37110 -1390 37190 -1370
rect 37110 -1430 37130 -1390
rect 37170 -1430 37190 -1390
rect 37110 -1450 37190 -1430
rect 37230 -1390 37290 -1310
rect 37230 -1430 37240 -1390
rect 37280 -1430 37290 -1390
rect 37230 -1450 37290 -1430
rect 37360 -1160 37400 -990
rect 36360 -1490 36400 -1450
rect 37240 -1490 37280 -1450
rect 37360 -1490 37400 -1320
rect 36240 -1530 37400 -1490
rect 37470 -990 38080 -950
rect 38240 -990 38850 -950
rect 37470 -1160 37510 -990
rect 37790 -1050 37870 -1030
rect 37790 -1090 37810 -1050
rect 37850 -1090 37870 -1050
rect 37790 -1110 37870 -1090
rect 38010 -1050 38090 -1030
rect 38010 -1090 38030 -1050
rect 38070 -1090 38090 -1050
rect 38010 -1110 38090 -1090
rect 38130 -1050 38190 -1030
rect 38130 -1090 38140 -1050
rect 38180 -1090 38190 -1050
rect 38130 -1110 38190 -1090
rect 38230 -1050 38310 -1030
rect 38230 -1090 38250 -1050
rect 38290 -1090 38310 -1050
rect 38230 -1110 38310 -1090
rect 38450 -1050 38530 -1030
rect 38450 -1090 38470 -1050
rect 38510 -1090 38530 -1050
rect 38450 -1110 38530 -1090
rect 37810 -1150 37850 -1110
rect 38030 -1150 38070 -1110
rect 38250 -1150 38290 -1110
rect 38470 -1150 38510 -1110
rect 37470 -1490 37510 -1320
rect 37580 -1170 37640 -1150
rect 37580 -1210 37590 -1170
rect 37630 -1210 37640 -1170
rect 37580 -1270 37640 -1210
rect 37580 -1310 37590 -1270
rect 37630 -1310 37640 -1270
rect 37580 -1390 37640 -1310
rect 37690 -1170 37750 -1150
rect 37690 -1210 37700 -1170
rect 37740 -1210 37750 -1170
rect 37690 -1270 37750 -1210
rect 37690 -1310 37700 -1270
rect 37740 -1310 37750 -1270
rect 37690 -1330 37750 -1310
rect 37800 -1170 37860 -1150
rect 37800 -1210 37810 -1170
rect 37850 -1210 37860 -1170
rect 37800 -1270 37860 -1210
rect 37800 -1310 37810 -1270
rect 37850 -1310 37860 -1270
rect 37800 -1330 37860 -1310
rect 37910 -1170 37970 -1150
rect 37910 -1210 37920 -1170
rect 37960 -1210 37970 -1170
rect 37910 -1270 37970 -1210
rect 37910 -1310 37920 -1270
rect 37960 -1310 37970 -1270
rect 37910 -1330 37970 -1310
rect 38020 -1170 38080 -1150
rect 38020 -1210 38030 -1170
rect 38070 -1210 38080 -1170
rect 38020 -1270 38080 -1210
rect 38020 -1310 38030 -1270
rect 38070 -1310 38080 -1270
rect 38020 -1330 38080 -1310
rect 38130 -1170 38190 -1150
rect 38130 -1210 38140 -1170
rect 38180 -1210 38190 -1170
rect 38130 -1270 38190 -1210
rect 38130 -1310 38140 -1270
rect 38180 -1310 38190 -1270
rect 38130 -1330 38190 -1310
rect 38240 -1170 38300 -1150
rect 38240 -1210 38250 -1170
rect 38290 -1210 38300 -1170
rect 38240 -1270 38300 -1210
rect 38240 -1310 38250 -1270
rect 38290 -1310 38300 -1270
rect 38240 -1330 38300 -1310
rect 38350 -1170 38410 -1150
rect 38350 -1210 38360 -1170
rect 38400 -1210 38410 -1170
rect 38350 -1270 38410 -1210
rect 38350 -1310 38360 -1270
rect 38400 -1310 38410 -1270
rect 38350 -1330 38410 -1310
rect 38460 -1170 38520 -1150
rect 38460 -1210 38470 -1170
rect 38510 -1210 38520 -1170
rect 38460 -1270 38520 -1210
rect 38460 -1310 38470 -1270
rect 38510 -1310 38520 -1270
rect 38460 -1330 38520 -1310
rect 38570 -1170 38630 -1150
rect 38570 -1210 38580 -1170
rect 38620 -1210 38630 -1170
rect 38570 -1270 38630 -1210
rect 38570 -1310 38580 -1270
rect 38620 -1310 38630 -1270
rect 38570 -1330 38630 -1310
rect 38680 -1170 38740 -1150
rect 38680 -1210 38690 -1170
rect 38730 -1210 38740 -1170
rect 38680 -1270 38740 -1210
rect 38680 -1310 38690 -1270
rect 38730 -1310 38740 -1270
rect 37580 -1430 37590 -1390
rect 37630 -1430 37640 -1390
rect 37580 -1450 37640 -1430
rect 37700 -1370 37740 -1330
rect 37920 -1370 37960 -1330
rect 38140 -1370 38180 -1330
rect 38360 -1370 38400 -1330
rect 38580 -1370 38620 -1330
rect 37700 -1390 37810 -1370
rect 37700 -1430 37750 -1390
rect 37790 -1430 37810 -1390
rect 37700 -1450 37810 -1430
rect 37900 -1390 37980 -1370
rect 37900 -1430 37920 -1390
rect 37960 -1430 37980 -1390
rect 37900 -1450 37980 -1430
rect 38120 -1390 38200 -1370
rect 38120 -1430 38140 -1390
rect 38180 -1430 38200 -1390
rect 38120 -1450 38200 -1430
rect 38340 -1390 38420 -1370
rect 38340 -1430 38360 -1390
rect 38400 -1430 38420 -1390
rect 38340 -1450 38420 -1430
rect 38560 -1390 38640 -1370
rect 38560 -1430 38580 -1390
rect 38620 -1430 38640 -1390
rect 38560 -1450 38640 -1430
rect 38680 -1390 38740 -1310
rect 38680 -1430 38690 -1390
rect 38730 -1430 38740 -1390
rect 38680 -1450 38740 -1430
rect 38810 -1160 38850 -990
rect 37590 -1490 37630 -1450
rect 38690 -1490 38730 -1450
rect 38810 -1490 38850 -1320
rect 37470 -1530 38080 -1490
rect 38240 -1530 38850 -1490
rect 38920 -990 39360 -950
rect 39520 -990 40080 -950
rect 38920 -1160 38960 -990
rect 39240 -1050 39320 -1030
rect 39240 -1090 39260 -1050
rect 39300 -1090 39320 -1050
rect 39240 -1110 39320 -1090
rect 39360 -1050 39420 -1030
rect 39360 -1090 39370 -1050
rect 39410 -1090 39420 -1050
rect 39360 -1110 39420 -1090
rect 39460 -1050 39540 -1030
rect 39460 -1090 39480 -1050
rect 39520 -1090 39540 -1050
rect 39460 -1110 39540 -1090
rect 39680 -1050 39760 -1030
rect 39680 -1090 39700 -1050
rect 39740 -1090 39760 -1050
rect 39680 -1110 39760 -1090
rect 39260 -1150 39300 -1110
rect 39480 -1150 39520 -1110
rect 39700 -1150 39740 -1110
rect 38920 -1490 38960 -1320
rect 39030 -1170 39090 -1150
rect 39030 -1210 39040 -1170
rect 39080 -1210 39090 -1170
rect 39030 -1270 39090 -1210
rect 39030 -1310 39040 -1270
rect 39080 -1310 39090 -1270
rect 39030 -1390 39090 -1310
rect 39140 -1170 39200 -1150
rect 39140 -1210 39150 -1170
rect 39190 -1210 39200 -1170
rect 39140 -1270 39200 -1210
rect 39140 -1310 39150 -1270
rect 39190 -1310 39200 -1270
rect 39140 -1330 39200 -1310
rect 39250 -1170 39310 -1150
rect 39250 -1210 39260 -1170
rect 39300 -1210 39310 -1170
rect 39250 -1270 39310 -1210
rect 39250 -1310 39260 -1270
rect 39300 -1310 39310 -1270
rect 39250 -1330 39310 -1310
rect 39360 -1170 39420 -1150
rect 39360 -1210 39370 -1170
rect 39410 -1210 39420 -1170
rect 39360 -1270 39420 -1210
rect 39360 -1310 39370 -1270
rect 39410 -1310 39420 -1270
rect 39360 -1330 39420 -1310
rect 39470 -1170 39530 -1150
rect 39470 -1210 39480 -1170
rect 39520 -1210 39530 -1170
rect 39470 -1270 39530 -1210
rect 39470 -1310 39480 -1270
rect 39520 -1310 39530 -1270
rect 39470 -1330 39530 -1310
rect 39580 -1170 39640 -1150
rect 39580 -1210 39590 -1170
rect 39630 -1210 39640 -1170
rect 39580 -1270 39640 -1210
rect 39580 -1310 39590 -1270
rect 39630 -1310 39640 -1270
rect 39580 -1330 39640 -1310
rect 39690 -1170 39750 -1150
rect 39690 -1210 39700 -1170
rect 39740 -1210 39750 -1170
rect 39690 -1270 39750 -1210
rect 39690 -1310 39700 -1270
rect 39740 -1310 39750 -1270
rect 39690 -1330 39750 -1310
rect 39800 -1170 39860 -1150
rect 39800 -1210 39810 -1170
rect 39850 -1210 39860 -1170
rect 39800 -1270 39860 -1210
rect 39800 -1310 39810 -1270
rect 39850 -1310 39860 -1270
rect 39800 -1330 39860 -1310
rect 39910 -1170 39970 -1150
rect 39910 -1210 39920 -1170
rect 39960 -1210 39970 -1170
rect 39910 -1270 39970 -1210
rect 39910 -1310 39920 -1270
rect 39960 -1310 39970 -1270
rect 39150 -1370 39190 -1330
rect 39370 -1370 39410 -1330
rect 39590 -1370 39630 -1330
rect 39810 -1370 39850 -1330
rect 39030 -1430 39040 -1390
rect 39080 -1430 39090 -1390
rect 39030 -1450 39090 -1430
rect 39130 -1390 39210 -1370
rect 39130 -1430 39150 -1390
rect 39190 -1430 39210 -1390
rect 39130 -1450 39210 -1430
rect 39350 -1390 39430 -1370
rect 39350 -1430 39370 -1390
rect 39410 -1430 39430 -1390
rect 39350 -1450 39430 -1430
rect 39570 -1390 39650 -1370
rect 39570 -1430 39590 -1390
rect 39630 -1430 39650 -1390
rect 39570 -1450 39650 -1430
rect 39790 -1390 39870 -1370
rect 39790 -1430 39810 -1390
rect 39850 -1430 39870 -1390
rect 39790 -1450 39870 -1430
rect 39910 -1390 39970 -1310
rect 39910 -1430 39920 -1390
rect 39960 -1430 39970 -1390
rect 39910 -1450 39970 -1430
rect 40040 -1160 40080 -990
rect 39040 -1490 39080 -1450
rect 39920 -1490 39960 -1450
rect 40040 -1490 40080 -1320
rect 38920 -1530 40080 -1490
rect 44050 -2720 45180 -2680
rect 45340 -2720 46470 -2680
rect 44050 -2840 44090 -2720
rect 44132 -2830 44222 -2820
rect 44132 -2880 44152 -2830
rect 44202 -2880 44222 -2830
rect 44132 -2890 44222 -2880
rect 46260 -2940 46330 -2890
rect 44050 -3110 44090 -3000
rect 44132 -2950 44222 -2940
rect 44132 -3000 44152 -2950
rect 44202 -3000 44222 -2950
rect 44132 -3010 44222 -3000
rect 46430 -2840 46470 -2720
rect 46430 -3110 46470 -3000
rect 44050 -3150 45180 -3110
rect 45340 -3150 46470 -3110
rect 46620 -2990 47690 -2950
rect 47850 -2990 49010 -2950
rect 45230 -3210 45270 -3150
rect 44050 -3250 45150 -3210
rect 45310 -3250 46410 -3210
rect 44050 -3370 44090 -3250
rect 44132 -3360 44222 -3350
rect 44132 -3410 44152 -3360
rect 44202 -3410 44222 -3360
rect 44132 -3420 44222 -3410
rect 46200 -3470 46270 -3420
rect 44050 -3640 44090 -3530
rect 44132 -3480 44222 -3470
rect 44132 -3530 44152 -3480
rect 44202 -3530 44222 -3480
rect 44132 -3540 44222 -3530
rect 46370 -3370 46410 -3250
rect 46620 -3350 46660 -2990
rect 46702 -3100 46792 -3090
rect 46702 -3150 46722 -3100
rect 46772 -3150 46792 -3100
rect 46702 -3160 46792 -3150
rect 48840 -3160 48920 -3090
rect 46702 -3220 46792 -3210
rect 46702 -3270 46722 -3220
rect 46772 -3270 46792 -3220
rect 46702 -3280 46792 -3270
rect 48770 -3330 48840 -3280
rect 46410 -3430 46450 -3410
rect 46430 -3470 46450 -3430
rect 46410 -3490 46450 -3470
rect 46580 -3430 46620 -3410
rect 46580 -3470 46600 -3430
rect 46580 -3490 46620 -3470
rect 45190 -3620 45270 -3600
rect 45190 -3640 45210 -3620
rect 45250 -3640 45270 -3620
rect 46370 -3640 46410 -3530
rect 44050 -3680 45150 -3640
rect 45310 -3680 46410 -3640
rect 45210 -3740 45250 -3680
rect 44440 -3780 45150 -3740
rect 45310 -3780 46040 -3740
rect 44440 -3840 44480 -3780
rect 46000 -3840 46040 -3780
rect 44522 -3890 44612 -3880
rect 44522 -3940 44542 -3890
rect 44592 -3940 44612 -3890
rect 44522 -3950 44612 -3940
rect 45868 -3890 45958 -3880
rect 45868 -3940 45888 -3890
rect 45938 -3940 45958 -3890
rect 45868 -3950 45958 -3940
rect 44440 -4060 44480 -4000
rect 46620 -3860 46660 -3510
rect 46712 -3400 46792 -3330
rect 46712 -3690 46752 -3400
rect 48880 -3450 48920 -3160
rect 48840 -3520 48920 -3450
rect 48970 -3350 49010 -2990
rect 46792 -3570 46862 -3520
rect 48840 -3580 48930 -3570
rect 48840 -3630 48860 -3580
rect 48910 -3630 48930 -3580
rect 48840 -3640 48930 -3630
rect 46712 -3760 46792 -3690
rect 48840 -3700 48930 -3680
rect 48840 -3750 48860 -3700
rect 48910 -3750 48930 -3700
rect 48840 -3770 48930 -3750
rect 48970 -3860 49010 -3510
rect 46620 -3900 47690 -3860
rect 47850 -3900 49010 -3860
rect 47750 -3960 47790 -3900
rect 46000 -4060 46040 -4000
rect 44440 -4100 45150 -4060
rect 45310 -4100 46040 -4060
rect 46950 -4000 47690 -3960
rect 47850 -4000 48600 -3960
rect 46950 -4060 46990 -4000
rect 45210 -4160 45250 -4100
rect 44440 -4200 45150 -4160
rect 45310 -4200 46040 -4160
rect 33610 -4246 37620 -4240
rect 33610 -4279 37624 -4246
rect 33610 -4313 33674 -4279
rect 33708 -4313 33764 -4279
rect 33798 -4313 33854 -4279
rect 33888 -4313 33944 -4279
rect 33978 -4313 34034 -4279
rect 34068 -4313 34124 -4279
rect 34158 -4313 34214 -4279
rect 34248 -4313 34304 -4279
rect 34338 -4313 34394 -4279
rect 34428 -4313 34484 -4279
rect 34518 -4313 34574 -4279
rect 34608 -4313 34664 -4279
rect 34698 -4313 34754 -4279
rect 34788 -4313 35034 -4279
rect 35068 -4313 35124 -4279
rect 35158 -4313 35214 -4279
rect 35248 -4313 35304 -4279
rect 35338 -4313 35394 -4279
rect 35428 -4313 35484 -4279
rect 35518 -4313 35574 -4279
rect 35608 -4313 35664 -4279
rect 35698 -4313 35754 -4279
rect 35788 -4313 35844 -4279
rect 35878 -4313 35934 -4279
rect 35968 -4313 36024 -4279
rect 36058 -4313 36114 -4279
rect 36148 -4313 36394 -4279
rect 36428 -4313 36484 -4279
rect 36518 -4313 36574 -4279
rect 36608 -4313 36664 -4279
rect 36698 -4313 36754 -4279
rect 36788 -4313 36844 -4279
rect 36878 -4313 36934 -4279
rect 36968 -4313 37024 -4279
rect 37058 -4313 37114 -4279
rect 37148 -4313 37204 -4279
rect 37238 -4313 37294 -4279
rect 37328 -4313 37384 -4279
rect 37418 -4313 37474 -4279
rect 37508 -4313 37624 -4279
rect 33610 -4380 37624 -4313
rect 33610 -4414 33651 -4380
rect 33685 -4414 34838 -4380
rect 34872 -4414 35011 -4380
rect 35045 -4414 36198 -4380
rect 36232 -4414 36371 -4380
rect 36405 -4414 37558 -4380
rect 37592 -4414 37624 -4380
rect 33610 -4428 37624 -4414
rect 33610 -4462 33874 -4428
rect 33908 -4462 33964 -4428
rect 33998 -4462 34054 -4428
rect 34088 -4462 34144 -4428
rect 34178 -4462 34234 -4428
rect 34268 -4462 34324 -4428
rect 34358 -4462 34414 -4428
rect 34448 -4462 34504 -4428
rect 34538 -4462 34594 -4428
rect 34628 -4462 35234 -4428
rect 35268 -4462 35324 -4428
rect 35358 -4462 35414 -4428
rect 35448 -4462 35504 -4428
rect 35538 -4462 35594 -4428
rect 35628 -4462 35684 -4428
rect 35718 -4462 35774 -4428
rect 35808 -4462 35864 -4428
rect 35898 -4462 35954 -4428
rect 35988 -4462 36594 -4428
rect 36628 -4462 36684 -4428
rect 36718 -4462 36774 -4428
rect 36808 -4462 36864 -4428
rect 36898 -4462 36954 -4428
rect 36988 -4462 37044 -4428
rect 37078 -4462 37134 -4428
rect 37168 -4462 37224 -4428
rect 37258 -4462 37314 -4428
rect 37348 -4462 37624 -4428
rect 33610 -4470 37624 -4462
rect 33610 -4490 33651 -4470
rect 33616 -4504 33651 -4490
rect 33685 -4486 34838 -4470
rect 33685 -4490 33798 -4486
rect 33685 -4504 33715 -4490
rect 33616 -4560 33715 -4504
rect 33616 -4594 33651 -4560
rect 33685 -4594 33715 -4560
rect 33616 -4650 33715 -4594
rect 33616 -4684 33651 -4650
rect 33685 -4684 33715 -4650
rect 33616 -4740 33715 -4684
rect 33616 -4774 33651 -4740
rect 33685 -4774 33715 -4740
rect 33616 -4830 33715 -4774
rect 33616 -4864 33651 -4830
rect 33685 -4864 33715 -4830
rect 33616 -4920 33715 -4864
rect 33616 -4954 33651 -4920
rect 33685 -4954 33715 -4920
rect 33616 -5010 33715 -4954
rect 33616 -5044 33651 -5010
rect 33685 -5044 33715 -5010
rect 33616 -5100 33715 -5044
rect 33616 -5134 33651 -5100
rect 33685 -5134 33715 -5100
rect 33616 -5190 33715 -5134
rect 33616 -5224 33651 -5190
rect 33685 -5224 33715 -5190
rect 33616 -5280 33715 -5224
rect 33616 -5314 33651 -5280
rect 33685 -5314 33715 -5280
rect 33616 -5370 33715 -5314
rect 33616 -5404 33651 -5370
rect 33685 -5404 33715 -5370
rect 33779 -4520 33798 -4490
rect 33832 -4490 34838 -4486
rect 33832 -4520 33851 -4490
rect 33779 -4576 33851 -4520
rect 34669 -4520 34741 -4490
rect 33779 -4610 33798 -4576
rect 33832 -4610 33851 -4576
rect 33779 -4666 33851 -4610
rect 33779 -4700 33798 -4666
rect 33832 -4700 33851 -4666
rect 33779 -4756 33851 -4700
rect 33779 -4790 33798 -4756
rect 33832 -4790 33851 -4756
rect 33779 -4846 33851 -4790
rect 33779 -4880 33798 -4846
rect 33832 -4880 33851 -4846
rect 33779 -4936 33851 -4880
rect 33779 -4970 33798 -4936
rect 33832 -4970 33851 -4936
rect 33779 -5026 33851 -4970
rect 33779 -5060 33798 -5026
rect 33832 -5060 33851 -5026
rect 33779 -5116 33851 -5060
rect 33779 -5150 33798 -5116
rect 33832 -5150 33851 -5116
rect 33779 -5206 33851 -5150
rect 33779 -5240 33798 -5206
rect 33832 -5240 33851 -5206
rect 33913 -4602 34607 -4543
rect 33913 -4636 33972 -4602
rect 34006 -4630 34062 -4602
rect 34034 -4636 34062 -4630
rect 34096 -4630 34152 -4602
rect 34096 -4636 34100 -4630
rect 33913 -4664 34000 -4636
rect 34034 -4664 34100 -4636
rect 34134 -4636 34152 -4630
rect 34186 -4630 34242 -4602
rect 34186 -4636 34200 -4630
rect 34134 -4664 34200 -4636
rect 34234 -4636 34242 -4630
rect 34276 -4630 34332 -4602
rect 34366 -4630 34422 -4602
rect 34456 -4630 34512 -4602
rect 34276 -4636 34300 -4630
rect 34366 -4636 34400 -4630
rect 34456 -4636 34500 -4630
rect 34546 -4636 34607 -4602
rect 34234 -4664 34300 -4636
rect 34334 -4664 34400 -4636
rect 34434 -4664 34500 -4636
rect 34534 -4664 34607 -4636
rect 33913 -4692 34607 -4664
rect 33913 -4726 33972 -4692
rect 34006 -4726 34062 -4692
rect 34096 -4726 34152 -4692
rect 34186 -4726 34242 -4692
rect 34276 -4726 34332 -4692
rect 34366 -4726 34422 -4692
rect 34456 -4726 34512 -4692
rect 34546 -4726 34607 -4692
rect 33913 -4730 34607 -4726
rect 33913 -4764 34000 -4730
rect 34034 -4764 34100 -4730
rect 34134 -4764 34200 -4730
rect 34234 -4764 34300 -4730
rect 34334 -4764 34400 -4730
rect 34434 -4764 34500 -4730
rect 34534 -4764 34607 -4730
rect 33913 -4782 34607 -4764
rect 33913 -4816 33972 -4782
rect 34006 -4816 34062 -4782
rect 34096 -4816 34152 -4782
rect 34186 -4816 34242 -4782
rect 34276 -4816 34332 -4782
rect 34366 -4816 34422 -4782
rect 34456 -4816 34512 -4782
rect 34546 -4816 34607 -4782
rect 33913 -4830 34607 -4816
rect 33913 -4864 34000 -4830
rect 34034 -4864 34100 -4830
rect 34134 -4864 34200 -4830
rect 34234 -4864 34300 -4830
rect 34334 -4864 34400 -4830
rect 34434 -4864 34500 -4830
rect 34534 -4864 34607 -4830
rect 33913 -4872 34607 -4864
rect 33913 -4906 33972 -4872
rect 34006 -4906 34062 -4872
rect 34096 -4906 34152 -4872
rect 34186 -4906 34242 -4872
rect 34276 -4906 34332 -4872
rect 34366 -4906 34422 -4872
rect 34456 -4906 34512 -4872
rect 34546 -4906 34607 -4872
rect 33913 -4930 34607 -4906
rect 33913 -4962 34000 -4930
rect 34034 -4962 34100 -4930
rect 33913 -4996 33972 -4962
rect 34034 -4964 34062 -4962
rect 34006 -4996 34062 -4964
rect 34096 -4964 34100 -4962
rect 34134 -4962 34200 -4930
rect 34134 -4964 34152 -4962
rect 34096 -4996 34152 -4964
rect 34186 -4964 34200 -4962
rect 34234 -4962 34300 -4930
rect 34334 -4962 34400 -4930
rect 34434 -4962 34500 -4930
rect 34534 -4962 34607 -4930
rect 34234 -4964 34242 -4962
rect 34186 -4996 34242 -4964
rect 34276 -4964 34300 -4962
rect 34366 -4964 34400 -4962
rect 34456 -4964 34500 -4962
rect 34276 -4996 34332 -4964
rect 34366 -4996 34422 -4964
rect 34456 -4996 34512 -4964
rect 34546 -4996 34607 -4962
rect 33913 -5030 34607 -4996
rect 33913 -5052 34000 -5030
rect 34034 -5052 34100 -5030
rect 33913 -5086 33972 -5052
rect 34034 -5064 34062 -5052
rect 34006 -5086 34062 -5064
rect 34096 -5064 34100 -5052
rect 34134 -5052 34200 -5030
rect 34134 -5064 34152 -5052
rect 34096 -5086 34152 -5064
rect 34186 -5064 34200 -5052
rect 34234 -5052 34300 -5030
rect 34334 -5052 34400 -5030
rect 34434 -5052 34500 -5030
rect 34534 -5052 34607 -5030
rect 34234 -5064 34242 -5052
rect 34186 -5086 34242 -5064
rect 34276 -5064 34300 -5052
rect 34366 -5064 34400 -5052
rect 34456 -5064 34500 -5052
rect 34276 -5086 34332 -5064
rect 34366 -5086 34422 -5064
rect 34456 -5086 34512 -5064
rect 34546 -5086 34607 -5052
rect 33913 -5130 34607 -5086
rect 33913 -5142 34000 -5130
rect 34034 -5142 34100 -5130
rect 33913 -5176 33972 -5142
rect 34034 -5164 34062 -5142
rect 34006 -5176 34062 -5164
rect 34096 -5164 34100 -5142
rect 34134 -5142 34200 -5130
rect 34134 -5164 34152 -5142
rect 34096 -5176 34152 -5164
rect 34186 -5164 34200 -5142
rect 34234 -5142 34300 -5130
rect 34334 -5142 34400 -5130
rect 34434 -5142 34500 -5130
rect 34534 -5142 34607 -5130
rect 34234 -5164 34242 -5142
rect 34186 -5176 34242 -5164
rect 34276 -5164 34300 -5142
rect 34366 -5164 34400 -5142
rect 34456 -5164 34500 -5142
rect 34276 -5176 34332 -5164
rect 34366 -5176 34422 -5164
rect 34456 -5176 34512 -5164
rect 34546 -5176 34607 -5142
rect 33913 -5237 34607 -5176
rect 34669 -4554 34688 -4520
rect 34722 -4554 34741 -4520
rect 34669 -4610 34741 -4554
rect 34669 -4644 34688 -4610
rect 34722 -4644 34741 -4610
rect 34669 -4700 34741 -4644
rect 34669 -4734 34688 -4700
rect 34722 -4734 34741 -4700
rect 34669 -4790 34741 -4734
rect 34669 -4824 34688 -4790
rect 34722 -4824 34741 -4790
rect 34669 -4880 34741 -4824
rect 34669 -4914 34688 -4880
rect 34722 -4914 34741 -4880
rect 34669 -4970 34741 -4914
rect 34669 -5004 34688 -4970
rect 34722 -5004 34741 -4970
rect 34669 -5060 34741 -5004
rect 34669 -5094 34688 -5060
rect 34722 -5094 34741 -5060
rect 34669 -5150 34741 -5094
rect 34669 -5184 34688 -5150
rect 34722 -5184 34741 -5150
rect 33779 -5299 33851 -5240
rect 34669 -5240 34741 -5184
rect 34669 -5274 34688 -5240
rect 34722 -5274 34741 -5240
rect 34669 -5299 34741 -5274
rect 33779 -5318 34741 -5299
rect 33779 -5352 33855 -5318
rect 33889 -5352 33945 -5318
rect 33979 -5352 34035 -5318
rect 34069 -5352 34125 -5318
rect 34159 -5352 34215 -5318
rect 34249 -5352 34305 -5318
rect 34339 -5352 34395 -5318
rect 34429 -5352 34485 -5318
rect 34519 -5352 34575 -5318
rect 34609 -5352 34741 -5318
rect 33779 -5371 34741 -5352
rect 34805 -4504 34838 -4490
rect 34872 -4504 35011 -4470
rect 35045 -4486 36198 -4470
rect 35045 -4490 35158 -4486
rect 35045 -4504 35075 -4490
rect 34805 -4560 35075 -4504
rect 34805 -4594 34838 -4560
rect 34872 -4594 35011 -4560
rect 35045 -4594 35075 -4560
rect 34805 -4650 35075 -4594
rect 34805 -4684 34838 -4650
rect 34872 -4684 35011 -4650
rect 35045 -4684 35075 -4650
rect 34805 -4740 35075 -4684
rect 34805 -4774 34838 -4740
rect 34872 -4774 35011 -4740
rect 35045 -4774 35075 -4740
rect 34805 -4830 35075 -4774
rect 34805 -4864 34838 -4830
rect 34872 -4864 35011 -4830
rect 35045 -4864 35075 -4830
rect 34805 -4920 35075 -4864
rect 34805 -4954 34838 -4920
rect 34872 -4954 35011 -4920
rect 35045 -4954 35075 -4920
rect 34805 -5010 35075 -4954
rect 34805 -5044 34838 -5010
rect 34872 -5044 35011 -5010
rect 35045 -5044 35075 -5010
rect 34805 -5100 35075 -5044
rect 34805 -5134 34838 -5100
rect 34872 -5134 35011 -5100
rect 35045 -5134 35075 -5100
rect 34805 -5190 35075 -5134
rect 34805 -5224 34838 -5190
rect 34872 -5224 35011 -5190
rect 35045 -5224 35075 -5190
rect 34805 -5280 35075 -5224
rect 34805 -5314 34838 -5280
rect 34872 -5314 35011 -5280
rect 35045 -5314 35075 -5280
rect 34805 -5370 35075 -5314
rect 33616 -5435 33715 -5404
rect 34805 -5404 34838 -5370
rect 34872 -5404 35011 -5370
rect 35045 -5404 35075 -5370
rect 35139 -4520 35158 -4490
rect 35192 -4490 36198 -4486
rect 35192 -4520 35211 -4490
rect 35139 -4576 35211 -4520
rect 36029 -4520 36101 -4490
rect 35139 -4610 35158 -4576
rect 35192 -4610 35211 -4576
rect 35139 -4666 35211 -4610
rect 35139 -4700 35158 -4666
rect 35192 -4700 35211 -4666
rect 35139 -4756 35211 -4700
rect 35139 -4790 35158 -4756
rect 35192 -4790 35211 -4756
rect 35139 -4846 35211 -4790
rect 35139 -4880 35158 -4846
rect 35192 -4880 35211 -4846
rect 35139 -4936 35211 -4880
rect 35139 -4970 35158 -4936
rect 35192 -4970 35211 -4936
rect 35139 -5026 35211 -4970
rect 35139 -5060 35158 -5026
rect 35192 -5060 35211 -5026
rect 35139 -5116 35211 -5060
rect 35139 -5150 35158 -5116
rect 35192 -5150 35211 -5116
rect 35139 -5206 35211 -5150
rect 35139 -5240 35158 -5206
rect 35192 -5240 35211 -5206
rect 35273 -4602 35967 -4543
rect 35273 -4636 35332 -4602
rect 35366 -4630 35422 -4602
rect 35394 -4636 35422 -4630
rect 35456 -4630 35512 -4602
rect 35456 -4636 35460 -4630
rect 35273 -4664 35360 -4636
rect 35394 -4664 35460 -4636
rect 35494 -4636 35512 -4630
rect 35546 -4630 35602 -4602
rect 35546 -4636 35560 -4630
rect 35494 -4664 35560 -4636
rect 35594 -4636 35602 -4630
rect 35636 -4630 35692 -4602
rect 35726 -4630 35782 -4602
rect 35816 -4630 35872 -4602
rect 35636 -4636 35660 -4630
rect 35726 -4636 35760 -4630
rect 35816 -4636 35860 -4630
rect 35906 -4636 35967 -4602
rect 35594 -4664 35660 -4636
rect 35694 -4664 35760 -4636
rect 35794 -4664 35860 -4636
rect 35894 -4664 35967 -4636
rect 35273 -4692 35967 -4664
rect 35273 -4726 35332 -4692
rect 35366 -4726 35422 -4692
rect 35456 -4726 35512 -4692
rect 35546 -4726 35602 -4692
rect 35636 -4726 35692 -4692
rect 35726 -4726 35782 -4692
rect 35816 -4726 35872 -4692
rect 35906 -4726 35967 -4692
rect 35273 -4730 35967 -4726
rect 35273 -4764 35360 -4730
rect 35394 -4764 35460 -4730
rect 35494 -4764 35560 -4730
rect 35594 -4764 35660 -4730
rect 35694 -4764 35760 -4730
rect 35794 -4764 35860 -4730
rect 35894 -4764 35967 -4730
rect 35273 -4782 35967 -4764
rect 35273 -4816 35332 -4782
rect 35366 -4816 35422 -4782
rect 35456 -4816 35512 -4782
rect 35546 -4816 35602 -4782
rect 35636 -4816 35692 -4782
rect 35726 -4816 35782 -4782
rect 35816 -4816 35872 -4782
rect 35906 -4816 35967 -4782
rect 35273 -4830 35967 -4816
rect 35273 -4864 35360 -4830
rect 35394 -4864 35460 -4830
rect 35494 -4864 35560 -4830
rect 35594 -4864 35660 -4830
rect 35694 -4864 35760 -4830
rect 35794 -4864 35860 -4830
rect 35894 -4864 35967 -4830
rect 35273 -4872 35967 -4864
rect 35273 -4906 35332 -4872
rect 35366 -4906 35422 -4872
rect 35456 -4906 35512 -4872
rect 35546 -4906 35602 -4872
rect 35636 -4906 35692 -4872
rect 35726 -4906 35782 -4872
rect 35816 -4906 35872 -4872
rect 35906 -4906 35967 -4872
rect 35273 -4930 35967 -4906
rect 35273 -4962 35360 -4930
rect 35394 -4962 35460 -4930
rect 35273 -4996 35332 -4962
rect 35394 -4964 35422 -4962
rect 35366 -4996 35422 -4964
rect 35456 -4964 35460 -4962
rect 35494 -4962 35560 -4930
rect 35494 -4964 35512 -4962
rect 35456 -4996 35512 -4964
rect 35546 -4964 35560 -4962
rect 35594 -4962 35660 -4930
rect 35694 -4962 35760 -4930
rect 35794 -4962 35860 -4930
rect 35894 -4962 35967 -4930
rect 35594 -4964 35602 -4962
rect 35546 -4996 35602 -4964
rect 35636 -4964 35660 -4962
rect 35726 -4964 35760 -4962
rect 35816 -4964 35860 -4962
rect 35636 -4996 35692 -4964
rect 35726 -4996 35782 -4964
rect 35816 -4996 35872 -4964
rect 35906 -4996 35967 -4962
rect 35273 -5030 35967 -4996
rect 35273 -5052 35360 -5030
rect 35394 -5052 35460 -5030
rect 35273 -5086 35332 -5052
rect 35394 -5064 35422 -5052
rect 35366 -5086 35422 -5064
rect 35456 -5064 35460 -5052
rect 35494 -5052 35560 -5030
rect 35494 -5064 35512 -5052
rect 35456 -5086 35512 -5064
rect 35546 -5064 35560 -5052
rect 35594 -5052 35660 -5030
rect 35694 -5052 35760 -5030
rect 35794 -5052 35860 -5030
rect 35894 -5052 35967 -5030
rect 35594 -5064 35602 -5052
rect 35546 -5086 35602 -5064
rect 35636 -5064 35660 -5052
rect 35726 -5064 35760 -5052
rect 35816 -5064 35860 -5052
rect 35636 -5086 35692 -5064
rect 35726 -5086 35782 -5064
rect 35816 -5086 35872 -5064
rect 35906 -5086 35967 -5052
rect 35273 -5130 35967 -5086
rect 35273 -5142 35360 -5130
rect 35394 -5142 35460 -5130
rect 35273 -5176 35332 -5142
rect 35394 -5164 35422 -5142
rect 35366 -5176 35422 -5164
rect 35456 -5164 35460 -5142
rect 35494 -5142 35560 -5130
rect 35494 -5164 35512 -5142
rect 35456 -5176 35512 -5164
rect 35546 -5164 35560 -5142
rect 35594 -5142 35660 -5130
rect 35694 -5142 35760 -5130
rect 35794 -5142 35860 -5130
rect 35894 -5142 35967 -5130
rect 35594 -5164 35602 -5142
rect 35546 -5176 35602 -5164
rect 35636 -5164 35660 -5142
rect 35726 -5164 35760 -5142
rect 35816 -5164 35860 -5142
rect 35636 -5176 35692 -5164
rect 35726 -5176 35782 -5164
rect 35816 -5176 35872 -5164
rect 35906 -5176 35967 -5142
rect 35273 -5237 35967 -5176
rect 36029 -4554 36048 -4520
rect 36082 -4554 36101 -4520
rect 36029 -4610 36101 -4554
rect 36029 -4644 36048 -4610
rect 36082 -4644 36101 -4610
rect 36029 -4700 36101 -4644
rect 36029 -4734 36048 -4700
rect 36082 -4734 36101 -4700
rect 36029 -4790 36101 -4734
rect 36029 -4824 36048 -4790
rect 36082 -4824 36101 -4790
rect 36029 -4880 36101 -4824
rect 36029 -4914 36048 -4880
rect 36082 -4914 36101 -4880
rect 36029 -4970 36101 -4914
rect 36029 -5004 36048 -4970
rect 36082 -5004 36101 -4970
rect 36029 -5060 36101 -5004
rect 36029 -5094 36048 -5060
rect 36082 -5094 36101 -5060
rect 36029 -5150 36101 -5094
rect 36029 -5184 36048 -5150
rect 36082 -5184 36101 -5150
rect 35139 -5299 35211 -5240
rect 36029 -5240 36101 -5184
rect 36029 -5274 36048 -5240
rect 36082 -5274 36101 -5240
rect 36029 -5299 36101 -5274
rect 35139 -5318 36101 -5299
rect 35139 -5352 35215 -5318
rect 35249 -5352 35305 -5318
rect 35339 -5352 35395 -5318
rect 35429 -5352 35485 -5318
rect 35519 -5352 35575 -5318
rect 35609 -5352 35665 -5318
rect 35699 -5352 35755 -5318
rect 35789 -5352 35845 -5318
rect 35879 -5352 35935 -5318
rect 35969 -5352 36101 -5318
rect 35139 -5371 36101 -5352
rect 36165 -4504 36198 -4490
rect 36232 -4504 36371 -4470
rect 36405 -4486 37558 -4470
rect 36405 -4490 36518 -4486
rect 36405 -4504 36435 -4490
rect 36165 -4560 36435 -4504
rect 36165 -4594 36198 -4560
rect 36232 -4594 36371 -4560
rect 36405 -4594 36435 -4560
rect 36165 -4650 36435 -4594
rect 36165 -4684 36198 -4650
rect 36232 -4684 36371 -4650
rect 36405 -4684 36435 -4650
rect 36165 -4740 36435 -4684
rect 36165 -4774 36198 -4740
rect 36232 -4774 36371 -4740
rect 36405 -4774 36435 -4740
rect 36165 -4830 36435 -4774
rect 36165 -4864 36198 -4830
rect 36232 -4864 36371 -4830
rect 36405 -4864 36435 -4830
rect 36165 -4920 36435 -4864
rect 36165 -4954 36198 -4920
rect 36232 -4954 36371 -4920
rect 36405 -4954 36435 -4920
rect 36165 -5010 36435 -4954
rect 36165 -5044 36198 -5010
rect 36232 -5044 36371 -5010
rect 36405 -5044 36435 -5010
rect 36165 -5100 36435 -5044
rect 36165 -5134 36198 -5100
rect 36232 -5134 36371 -5100
rect 36405 -5134 36435 -5100
rect 36165 -5190 36435 -5134
rect 36165 -5224 36198 -5190
rect 36232 -5224 36371 -5190
rect 36405 -5224 36435 -5190
rect 36165 -5280 36435 -5224
rect 36165 -5314 36198 -5280
rect 36232 -5314 36371 -5280
rect 36405 -5314 36435 -5280
rect 36165 -5370 36435 -5314
rect 34805 -5435 35075 -5404
rect 36165 -5404 36198 -5370
rect 36232 -5404 36371 -5370
rect 36405 -5404 36435 -5370
rect 36499 -4520 36518 -4490
rect 36552 -4490 37558 -4486
rect 36552 -4520 36571 -4490
rect 36499 -4576 36571 -4520
rect 37389 -4520 37461 -4490
rect 36499 -4610 36518 -4576
rect 36552 -4610 36571 -4576
rect 36499 -4666 36571 -4610
rect 36499 -4700 36518 -4666
rect 36552 -4700 36571 -4666
rect 36499 -4756 36571 -4700
rect 36499 -4790 36518 -4756
rect 36552 -4790 36571 -4756
rect 36499 -4846 36571 -4790
rect 36499 -4880 36518 -4846
rect 36552 -4880 36571 -4846
rect 36499 -4936 36571 -4880
rect 36499 -4970 36518 -4936
rect 36552 -4970 36571 -4936
rect 36499 -5026 36571 -4970
rect 36499 -5060 36518 -5026
rect 36552 -5060 36571 -5026
rect 36499 -5116 36571 -5060
rect 36499 -5150 36518 -5116
rect 36552 -5150 36571 -5116
rect 36499 -5206 36571 -5150
rect 36499 -5240 36518 -5206
rect 36552 -5240 36571 -5206
rect 36633 -4602 37327 -4543
rect 36633 -4636 36692 -4602
rect 36726 -4630 36782 -4602
rect 36754 -4636 36782 -4630
rect 36816 -4630 36872 -4602
rect 36816 -4636 36820 -4630
rect 36633 -4664 36720 -4636
rect 36754 -4664 36820 -4636
rect 36854 -4636 36872 -4630
rect 36906 -4630 36962 -4602
rect 36906 -4636 36920 -4630
rect 36854 -4664 36920 -4636
rect 36954 -4636 36962 -4630
rect 36996 -4630 37052 -4602
rect 37086 -4630 37142 -4602
rect 37176 -4630 37232 -4602
rect 36996 -4636 37020 -4630
rect 37086 -4636 37120 -4630
rect 37176 -4636 37220 -4630
rect 37266 -4636 37327 -4602
rect 36954 -4664 37020 -4636
rect 37054 -4664 37120 -4636
rect 37154 -4664 37220 -4636
rect 37254 -4664 37327 -4636
rect 36633 -4692 37327 -4664
rect 36633 -4726 36692 -4692
rect 36726 -4726 36782 -4692
rect 36816 -4726 36872 -4692
rect 36906 -4726 36962 -4692
rect 36996 -4726 37052 -4692
rect 37086 -4726 37142 -4692
rect 37176 -4726 37232 -4692
rect 37266 -4726 37327 -4692
rect 36633 -4730 37327 -4726
rect 36633 -4764 36720 -4730
rect 36754 -4764 36820 -4730
rect 36854 -4764 36920 -4730
rect 36954 -4764 37020 -4730
rect 37054 -4764 37120 -4730
rect 37154 -4764 37220 -4730
rect 37254 -4764 37327 -4730
rect 36633 -4782 37327 -4764
rect 36633 -4816 36692 -4782
rect 36726 -4816 36782 -4782
rect 36816 -4816 36872 -4782
rect 36906 -4816 36962 -4782
rect 36996 -4816 37052 -4782
rect 37086 -4816 37142 -4782
rect 37176 -4816 37232 -4782
rect 37266 -4816 37327 -4782
rect 36633 -4830 37327 -4816
rect 36633 -4864 36720 -4830
rect 36754 -4864 36820 -4830
rect 36854 -4864 36920 -4830
rect 36954 -4864 37020 -4830
rect 37054 -4864 37120 -4830
rect 37154 -4864 37220 -4830
rect 37254 -4864 37327 -4830
rect 36633 -4872 37327 -4864
rect 36633 -4906 36692 -4872
rect 36726 -4906 36782 -4872
rect 36816 -4906 36872 -4872
rect 36906 -4906 36962 -4872
rect 36996 -4906 37052 -4872
rect 37086 -4906 37142 -4872
rect 37176 -4906 37232 -4872
rect 37266 -4906 37327 -4872
rect 36633 -4930 37327 -4906
rect 36633 -4962 36720 -4930
rect 36754 -4962 36820 -4930
rect 36633 -4996 36692 -4962
rect 36754 -4964 36782 -4962
rect 36726 -4996 36782 -4964
rect 36816 -4964 36820 -4962
rect 36854 -4962 36920 -4930
rect 36854 -4964 36872 -4962
rect 36816 -4996 36872 -4964
rect 36906 -4964 36920 -4962
rect 36954 -4962 37020 -4930
rect 37054 -4962 37120 -4930
rect 37154 -4962 37220 -4930
rect 37254 -4962 37327 -4930
rect 36954 -4964 36962 -4962
rect 36906 -4996 36962 -4964
rect 36996 -4964 37020 -4962
rect 37086 -4964 37120 -4962
rect 37176 -4964 37220 -4962
rect 36996 -4996 37052 -4964
rect 37086 -4996 37142 -4964
rect 37176 -4996 37232 -4964
rect 37266 -4996 37327 -4962
rect 36633 -5030 37327 -4996
rect 36633 -5052 36720 -5030
rect 36754 -5052 36820 -5030
rect 36633 -5086 36692 -5052
rect 36754 -5064 36782 -5052
rect 36726 -5086 36782 -5064
rect 36816 -5064 36820 -5052
rect 36854 -5052 36920 -5030
rect 36854 -5064 36872 -5052
rect 36816 -5086 36872 -5064
rect 36906 -5064 36920 -5052
rect 36954 -5052 37020 -5030
rect 37054 -5052 37120 -5030
rect 37154 -5052 37220 -5030
rect 37254 -5052 37327 -5030
rect 36954 -5064 36962 -5052
rect 36906 -5086 36962 -5064
rect 36996 -5064 37020 -5052
rect 37086 -5064 37120 -5052
rect 37176 -5064 37220 -5052
rect 36996 -5086 37052 -5064
rect 37086 -5086 37142 -5064
rect 37176 -5086 37232 -5064
rect 37266 -5086 37327 -5052
rect 36633 -5130 37327 -5086
rect 36633 -5142 36720 -5130
rect 36754 -5142 36820 -5130
rect 36633 -5176 36692 -5142
rect 36754 -5164 36782 -5142
rect 36726 -5176 36782 -5164
rect 36816 -5164 36820 -5142
rect 36854 -5142 36920 -5130
rect 36854 -5164 36872 -5142
rect 36816 -5176 36872 -5164
rect 36906 -5164 36920 -5142
rect 36954 -5142 37020 -5130
rect 37054 -5142 37120 -5130
rect 37154 -5142 37220 -5130
rect 37254 -5142 37327 -5130
rect 36954 -5164 36962 -5142
rect 36906 -5176 36962 -5164
rect 36996 -5164 37020 -5142
rect 37086 -5164 37120 -5142
rect 37176 -5164 37220 -5142
rect 36996 -5176 37052 -5164
rect 37086 -5176 37142 -5164
rect 37176 -5176 37232 -5164
rect 37266 -5176 37327 -5142
rect 36633 -5237 37327 -5176
rect 37389 -4554 37408 -4520
rect 37442 -4554 37461 -4520
rect 37389 -4610 37461 -4554
rect 37389 -4644 37408 -4610
rect 37442 -4644 37461 -4610
rect 37389 -4700 37461 -4644
rect 37389 -4734 37408 -4700
rect 37442 -4734 37461 -4700
rect 37389 -4790 37461 -4734
rect 37389 -4824 37408 -4790
rect 37442 -4824 37461 -4790
rect 37389 -4880 37461 -4824
rect 37389 -4914 37408 -4880
rect 37442 -4914 37461 -4880
rect 37389 -4970 37461 -4914
rect 37389 -5004 37408 -4970
rect 37442 -5004 37461 -4970
rect 37389 -5060 37461 -5004
rect 37389 -5094 37408 -5060
rect 37442 -5094 37461 -5060
rect 37389 -5150 37461 -5094
rect 37389 -5184 37408 -5150
rect 37442 -5184 37461 -5150
rect 36499 -5299 36571 -5240
rect 37389 -5240 37461 -5184
rect 37389 -5274 37408 -5240
rect 37442 -5274 37461 -5240
rect 37389 -5299 37461 -5274
rect 36499 -5318 37461 -5299
rect 36499 -5352 36575 -5318
rect 36609 -5352 36665 -5318
rect 36699 -5352 36755 -5318
rect 36789 -5352 36845 -5318
rect 36879 -5352 36935 -5318
rect 36969 -5352 37025 -5318
rect 37059 -5352 37115 -5318
rect 37149 -5352 37205 -5318
rect 37239 -5352 37295 -5318
rect 37329 -5352 37461 -5318
rect 36499 -5371 37461 -5352
rect 37525 -4504 37558 -4490
rect 37592 -4504 37624 -4470
rect 37525 -4560 37624 -4504
rect 44440 -4260 44480 -4200
rect 46000 -4260 46040 -4200
rect 44522 -4310 44612 -4300
rect 44522 -4360 44542 -4310
rect 44592 -4360 44612 -4310
rect 44522 -4370 44612 -4360
rect 45868 -4310 45958 -4300
rect 45868 -4360 45888 -4310
rect 45938 -4360 45958 -4310
rect 45868 -4370 45958 -4360
rect 44440 -4480 44480 -4420
rect 48560 -4060 48600 -4000
rect 47032 -4110 47122 -4100
rect 47032 -4160 47052 -4110
rect 47102 -4160 47122 -4110
rect 47032 -4170 47122 -4160
rect 48430 -4110 48520 -4100
rect 48430 -4160 48450 -4110
rect 48500 -4160 48520 -4110
rect 48430 -4170 48520 -4160
rect 46950 -4270 46990 -4220
rect 48560 -4270 48600 -4220
rect 46950 -4310 47690 -4270
rect 47850 -4310 48600 -4270
rect 46000 -4480 46040 -4420
rect 44440 -4520 45150 -4480
rect 45310 -4520 46040 -4480
rect 37525 -4594 37558 -4560
rect 37592 -4594 37624 -4560
rect 37525 -4650 37624 -4594
rect 37525 -4684 37558 -4650
rect 37592 -4684 37624 -4650
rect 37525 -4740 37624 -4684
rect 37525 -4774 37558 -4740
rect 37592 -4774 37624 -4740
rect 37525 -4830 37624 -4774
rect 37525 -4864 37558 -4830
rect 37592 -4864 37624 -4830
rect 37525 -4920 37624 -4864
rect 37525 -4954 37558 -4920
rect 37592 -4954 37624 -4920
rect 37525 -5010 37624 -4954
rect 37525 -5044 37558 -5010
rect 37592 -5044 37624 -5010
rect 37525 -5100 37624 -5044
rect 37525 -5134 37558 -5100
rect 37592 -5134 37624 -5100
rect 37525 -5190 37624 -5134
rect 37525 -5224 37558 -5190
rect 37592 -5224 37624 -5190
rect 37525 -5280 37624 -5224
rect 37525 -5314 37558 -5280
rect 37592 -5314 37624 -5280
rect 37525 -5370 37624 -5314
rect 36165 -5435 36435 -5404
rect 37525 -5404 37558 -5370
rect 37592 -5404 37624 -5370
rect 37525 -5435 37624 -5404
rect 33616 -5466 37624 -5435
rect 33616 -5500 33674 -5466
rect 33708 -5500 33764 -5466
rect 33798 -5500 33854 -5466
rect 33888 -5500 33944 -5466
rect 33978 -5500 34034 -5466
rect 34068 -5500 34124 -5466
rect 34158 -5500 34214 -5466
rect 34248 -5500 34304 -5466
rect 34338 -5500 34394 -5466
rect 34428 -5500 34484 -5466
rect 34518 -5500 34574 -5466
rect 34608 -5500 34664 -5466
rect 34698 -5500 34754 -5466
rect 34788 -5500 35034 -5466
rect 35068 -5500 35124 -5466
rect 35158 -5500 35214 -5466
rect 35248 -5500 35304 -5466
rect 35338 -5500 35394 -5466
rect 35428 -5500 35484 -5466
rect 35518 -5500 35574 -5466
rect 35608 -5500 35664 -5466
rect 35698 -5500 35754 -5466
rect 35788 -5500 35844 -5466
rect 35878 -5500 35934 -5466
rect 35968 -5500 36024 -5466
rect 36058 -5500 36114 -5466
rect 36148 -5500 36394 -5466
rect 36428 -5500 36484 -5466
rect 36518 -5500 36574 -5466
rect 36608 -5500 36664 -5466
rect 36698 -5500 36754 -5466
rect 36788 -5500 36844 -5466
rect 36878 -5500 36934 -5466
rect 36968 -5500 37024 -5466
rect 37058 -5500 37114 -5466
rect 37148 -5500 37204 -5466
rect 37238 -5500 37294 -5466
rect 37328 -5500 37384 -5466
rect 37418 -5500 37474 -5466
rect 37508 -5500 37624 -5466
rect 33616 -5534 37624 -5500
rect 34900 -5600 34980 -5534
rect 36260 -5600 36340 -5534
rect 33610 -5639 37630 -5600
rect 33610 -5673 33674 -5639
rect 33708 -5673 33764 -5639
rect 33798 -5673 33854 -5639
rect 33888 -5673 33944 -5639
rect 33978 -5673 34034 -5639
rect 34068 -5673 34124 -5639
rect 34158 -5673 34214 -5639
rect 34248 -5673 34304 -5639
rect 34338 -5673 34394 -5639
rect 34428 -5673 34484 -5639
rect 34518 -5673 34574 -5639
rect 34608 -5673 34664 -5639
rect 34698 -5673 34754 -5639
rect 34788 -5673 35034 -5639
rect 35068 -5673 35124 -5639
rect 35158 -5673 35214 -5639
rect 35248 -5673 35304 -5639
rect 35338 -5673 35394 -5639
rect 35428 -5673 35484 -5639
rect 35518 -5673 35574 -5639
rect 35608 -5673 35664 -5639
rect 35698 -5673 35754 -5639
rect 35788 -5673 35844 -5639
rect 35878 -5673 35934 -5639
rect 35968 -5673 36024 -5639
rect 36058 -5673 36114 -5639
rect 36148 -5673 36394 -5639
rect 36428 -5673 36484 -5639
rect 36518 -5673 36574 -5639
rect 36608 -5673 36664 -5639
rect 36698 -5673 36754 -5639
rect 36788 -5673 36844 -5639
rect 36878 -5673 36934 -5639
rect 36968 -5673 37024 -5639
rect 37058 -5673 37114 -5639
rect 37148 -5673 37204 -5639
rect 37238 -5673 37294 -5639
rect 37328 -5673 37384 -5639
rect 37418 -5673 37474 -5639
rect 37508 -5673 37630 -5639
rect 33610 -5740 37630 -5673
rect 33610 -5774 33651 -5740
rect 33685 -5774 34838 -5740
rect 34872 -5774 35011 -5740
rect 35045 -5774 36198 -5740
rect 36232 -5774 36371 -5740
rect 36405 -5774 37558 -5740
rect 37592 -5774 37630 -5740
rect 33610 -5788 37630 -5774
rect 33610 -5822 33874 -5788
rect 33908 -5822 33964 -5788
rect 33998 -5822 34054 -5788
rect 34088 -5822 34144 -5788
rect 34178 -5822 34234 -5788
rect 34268 -5822 34324 -5788
rect 34358 -5822 34414 -5788
rect 34448 -5822 34504 -5788
rect 34538 -5822 34594 -5788
rect 34628 -5822 35234 -5788
rect 35268 -5822 35324 -5788
rect 35358 -5822 35414 -5788
rect 35448 -5822 35504 -5788
rect 35538 -5822 35594 -5788
rect 35628 -5822 35684 -5788
rect 35718 -5822 35774 -5788
rect 35808 -5822 35864 -5788
rect 35898 -5822 35954 -5788
rect 35988 -5822 36594 -5788
rect 36628 -5822 36684 -5788
rect 36718 -5822 36774 -5788
rect 36808 -5822 36864 -5788
rect 36898 -5822 36954 -5788
rect 36988 -5822 37044 -5788
rect 37078 -5822 37134 -5788
rect 37168 -5822 37224 -5788
rect 37258 -5822 37314 -5788
rect 37348 -5822 37630 -5788
rect 33610 -5830 37630 -5822
rect 33610 -5850 33651 -5830
rect 33616 -5864 33651 -5850
rect 33685 -5846 34838 -5830
rect 33685 -5850 33798 -5846
rect 33685 -5864 33715 -5850
rect 33616 -5920 33715 -5864
rect 33616 -5954 33651 -5920
rect 33685 -5954 33715 -5920
rect 33616 -6010 33715 -5954
rect 33616 -6044 33651 -6010
rect 33685 -6044 33715 -6010
rect 33616 -6100 33715 -6044
rect 33616 -6134 33651 -6100
rect 33685 -6134 33715 -6100
rect 33616 -6190 33715 -6134
rect 33616 -6224 33651 -6190
rect 33685 -6224 33715 -6190
rect 33616 -6280 33715 -6224
rect 33616 -6314 33651 -6280
rect 33685 -6314 33715 -6280
rect 33616 -6370 33715 -6314
rect 33616 -6404 33651 -6370
rect 33685 -6404 33715 -6370
rect 33616 -6460 33715 -6404
rect 33616 -6494 33651 -6460
rect 33685 -6494 33715 -6460
rect 33616 -6550 33715 -6494
rect 33616 -6584 33651 -6550
rect 33685 -6584 33715 -6550
rect 33616 -6640 33715 -6584
rect 33616 -6674 33651 -6640
rect 33685 -6674 33715 -6640
rect 33616 -6730 33715 -6674
rect 33616 -6764 33651 -6730
rect 33685 -6764 33715 -6730
rect 33779 -5880 33798 -5850
rect 33832 -5850 34838 -5846
rect 33832 -5880 33851 -5850
rect 33779 -5936 33851 -5880
rect 34669 -5880 34741 -5850
rect 33779 -5970 33798 -5936
rect 33832 -5970 33851 -5936
rect 33779 -6026 33851 -5970
rect 33779 -6060 33798 -6026
rect 33832 -6060 33851 -6026
rect 33779 -6116 33851 -6060
rect 33779 -6150 33798 -6116
rect 33832 -6150 33851 -6116
rect 33779 -6206 33851 -6150
rect 33779 -6240 33798 -6206
rect 33832 -6240 33851 -6206
rect 33779 -6296 33851 -6240
rect 33779 -6330 33798 -6296
rect 33832 -6330 33851 -6296
rect 33779 -6386 33851 -6330
rect 33779 -6420 33798 -6386
rect 33832 -6420 33851 -6386
rect 33779 -6476 33851 -6420
rect 33779 -6510 33798 -6476
rect 33832 -6510 33851 -6476
rect 33779 -6566 33851 -6510
rect 33779 -6600 33798 -6566
rect 33832 -6600 33851 -6566
rect 33913 -5962 34607 -5903
rect 33913 -5996 33972 -5962
rect 34006 -5990 34062 -5962
rect 34034 -5996 34062 -5990
rect 34096 -5990 34152 -5962
rect 34096 -5996 34100 -5990
rect 33913 -6024 34000 -5996
rect 34034 -6024 34100 -5996
rect 34134 -5996 34152 -5990
rect 34186 -5990 34242 -5962
rect 34186 -5996 34200 -5990
rect 34134 -6024 34200 -5996
rect 34234 -5996 34242 -5990
rect 34276 -5990 34332 -5962
rect 34366 -5990 34422 -5962
rect 34456 -5990 34512 -5962
rect 34276 -5996 34300 -5990
rect 34366 -5996 34400 -5990
rect 34456 -5996 34500 -5990
rect 34546 -5996 34607 -5962
rect 34234 -6024 34300 -5996
rect 34334 -6024 34400 -5996
rect 34434 -6024 34500 -5996
rect 34534 -6024 34607 -5996
rect 33913 -6052 34607 -6024
rect 33913 -6086 33972 -6052
rect 34006 -6086 34062 -6052
rect 34096 -6086 34152 -6052
rect 34186 -6086 34242 -6052
rect 34276 -6086 34332 -6052
rect 34366 -6086 34422 -6052
rect 34456 -6086 34512 -6052
rect 34546 -6086 34607 -6052
rect 33913 -6090 34607 -6086
rect 33913 -6124 34000 -6090
rect 34034 -6124 34100 -6090
rect 34134 -6124 34200 -6090
rect 34234 -6124 34300 -6090
rect 34334 -6124 34400 -6090
rect 34434 -6124 34500 -6090
rect 34534 -6124 34607 -6090
rect 33913 -6142 34607 -6124
rect 33913 -6176 33972 -6142
rect 34006 -6176 34062 -6142
rect 34096 -6176 34152 -6142
rect 34186 -6176 34242 -6142
rect 34276 -6176 34332 -6142
rect 34366 -6176 34422 -6142
rect 34456 -6176 34512 -6142
rect 34546 -6176 34607 -6142
rect 33913 -6190 34607 -6176
rect 33913 -6224 34000 -6190
rect 34034 -6224 34100 -6190
rect 34134 -6224 34200 -6190
rect 34234 -6224 34300 -6190
rect 34334 -6224 34400 -6190
rect 34434 -6224 34500 -6190
rect 34534 -6224 34607 -6190
rect 33913 -6232 34607 -6224
rect 33913 -6266 33972 -6232
rect 34006 -6266 34062 -6232
rect 34096 -6266 34152 -6232
rect 34186 -6266 34242 -6232
rect 34276 -6266 34332 -6232
rect 34366 -6266 34422 -6232
rect 34456 -6266 34512 -6232
rect 34546 -6266 34607 -6232
rect 33913 -6290 34607 -6266
rect 33913 -6322 34000 -6290
rect 34034 -6322 34100 -6290
rect 33913 -6356 33972 -6322
rect 34034 -6324 34062 -6322
rect 34006 -6356 34062 -6324
rect 34096 -6324 34100 -6322
rect 34134 -6322 34200 -6290
rect 34134 -6324 34152 -6322
rect 34096 -6356 34152 -6324
rect 34186 -6324 34200 -6322
rect 34234 -6322 34300 -6290
rect 34334 -6322 34400 -6290
rect 34434 -6322 34500 -6290
rect 34534 -6322 34607 -6290
rect 34234 -6324 34242 -6322
rect 34186 -6356 34242 -6324
rect 34276 -6324 34300 -6322
rect 34366 -6324 34400 -6322
rect 34456 -6324 34500 -6322
rect 34276 -6356 34332 -6324
rect 34366 -6356 34422 -6324
rect 34456 -6356 34512 -6324
rect 34546 -6356 34607 -6322
rect 33913 -6390 34607 -6356
rect 33913 -6412 34000 -6390
rect 34034 -6412 34100 -6390
rect 33913 -6446 33972 -6412
rect 34034 -6424 34062 -6412
rect 34006 -6446 34062 -6424
rect 34096 -6424 34100 -6412
rect 34134 -6412 34200 -6390
rect 34134 -6424 34152 -6412
rect 34096 -6446 34152 -6424
rect 34186 -6424 34200 -6412
rect 34234 -6412 34300 -6390
rect 34334 -6412 34400 -6390
rect 34434 -6412 34500 -6390
rect 34534 -6412 34607 -6390
rect 34234 -6424 34242 -6412
rect 34186 -6446 34242 -6424
rect 34276 -6424 34300 -6412
rect 34366 -6424 34400 -6412
rect 34456 -6424 34500 -6412
rect 34276 -6446 34332 -6424
rect 34366 -6446 34422 -6424
rect 34456 -6446 34512 -6424
rect 34546 -6446 34607 -6412
rect 33913 -6490 34607 -6446
rect 33913 -6502 34000 -6490
rect 34034 -6502 34100 -6490
rect 33913 -6536 33972 -6502
rect 34034 -6524 34062 -6502
rect 34006 -6536 34062 -6524
rect 34096 -6524 34100 -6502
rect 34134 -6502 34200 -6490
rect 34134 -6524 34152 -6502
rect 34096 -6536 34152 -6524
rect 34186 -6524 34200 -6502
rect 34234 -6502 34300 -6490
rect 34334 -6502 34400 -6490
rect 34434 -6502 34500 -6490
rect 34534 -6502 34607 -6490
rect 34234 -6524 34242 -6502
rect 34186 -6536 34242 -6524
rect 34276 -6524 34300 -6502
rect 34366 -6524 34400 -6502
rect 34456 -6524 34500 -6502
rect 34276 -6536 34332 -6524
rect 34366 -6536 34422 -6524
rect 34456 -6536 34512 -6524
rect 34546 -6536 34607 -6502
rect 33913 -6597 34607 -6536
rect 34669 -5914 34688 -5880
rect 34722 -5914 34741 -5880
rect 34669 -5970 34741 -5914
rect 34669 -6004 34688 -5970
rect 34722 -6004 34741 -5970
rect 34669 -6060 34741 -6004
rect 34669 -6094 34688 -6060
rect 34722 -6094 34741 -6060
rect 34669 -6150 34741 -6094
rect 34669 -6184 34688 -6150
rect 34722 -6184 34741 -6150
rect 34669 -6240 34741 -6184
rect 34669 -6274 34688 -6240
rect 34722 -6274 34741 -6240
rect 34669 -6330 34741 -6274
rect 34669 -6364 34688 -6330
rect 34722 -6364 34741 -6330
rect 34669 -6420 34741 -6364
rect 34669 -6454 34688 -6420
rect 34722 -6454 34741 -6420
rect 34669 -6510 34741 -6454
rect 34669 -6544 34688 -6510
rect 34722 -6544 34741 -6510
rect 33779 -6659 33851 -6600
rect 34669 -6600 34741 -6544
rect 34669 -6634 34688 -6600
rect 34722 -6634 34741 -6600
rect 34669 -6659 34741 -6634
rect 33779 -6678 34741 -6659
rect 33779 -6712 33855 -6678
rect 33889 -6712 33945 -6678
rect 33979 -6712 34035 -6678
rect 34069 -6712 34125 -6678
rect 34159 -6712 34215 -6678
rect 34249 -6712 34305 -6678
rect 34339 -6712 34395 -6678
rect 34429 -6712 34485 -6678
rect 34519 -6712 34575 -6678
rect 34609 -6712 34741 -6678
rect 33779 -6731 34741 -6712
rect 34805 -5864 34838 -5850
rect 34872 -5864 35011 -5830
rect 35045 -5846 36198 -5830
rect 35045 -5850 35158 -5846
rect 35045 -5864 35075 -5850
rect 34805 -5920 35075 -5864
rect 34805 -5954 34838 -5920
rect 34872 -5954 35011 -5920
rect 35045 -5954 35075 -5920
rect 34805 -6010 35075 -5954
rect 34805 -6044 34838 -6010
rect 34872 -6044 35011 -6010
rect 35045 -6044 35075 -6010
rect 34805 -6100 35075 -6044
rect 34805 -6134 34838 -6100
rect 34872 -6134 35011 -6100
rect 35045 -6134 35075 -6100
rect 34805 -6190 35075 -6134
rect 34805 -6224 34838 -6190
rect 34872 -6224 35011 -6190
rect 35045 -6224 35075 -6190
rect 34805 -6280 35075 -6224
rect 34805 -6314 34838 -6280
rect 34872 -6314 35011 -6280
rect 35045 -6314 35075 -6280
rect 34805 -6370 35075 -6314
rect 34805 -6404 34838 -6370
rect 34872 -6404 35011 -6370
rect 35045 -6404 35075 -6370
rect 34805 -6460 35075 -6404
rect 34805 -6494 34838 -6460
rect 34872 -6494 35011 -6460
rect 35045 -6494 35075 -6460
rect 34805 -6550 35075 -6494
rect 34805 -6584 34838 -6550
rect 34872 -6584 35011 -6550
rect 35045 -6584 35075 -6550
rect 34805 -6640 35075 -6584
rect 34805 -6674 34838 -6640
rect 34872 -6674 35011 -6640
rect 35045 -6674 35075 -6640
rect 34805 -6730 35075 -6674
rect 33616 -6795 33715 -6764
rect 34805 -6764 34838 -6730
rect 34872 -6764 35011 -6730
rect 35045 -6764 35075 -6730
rect 35139 -5880 35158 -5850
rect 35192 -5850 36198 -5846
rect 35192 -5880 35211 -5850
rect 35139 -5936 35211 -5880
rect 36029 -5880 36101 -5850
rect 35139 -5970 35158 -5936
rect 35192 -5970 35211 -5936
rect 35139 -6026 35211 -5970
rect 35139 -6060 35158 -6026
rect 35192 -6060 35211 -6026
rect 35139 -6116 35211 -6060
rect 35139 -6150 35158 -6116
rect 35192 -6150 35211 -6116
rect 35139 -6206 35211 -6150
rect 35139 -6240 35158 -6206
rect 35192 -6240 35211 -6206
rect 35139 -6296 35211 -6240
rect 35139 -6330 35158 -6296
rect 35192 -6330 35211 -6296
rect 35139 -6386 35211 -6330
rect 35139 -6420 35158 -6386
rect 35192 -6420 35211 -6386
rect 35139 -6476 35211 -6420
rect 35139 -6510 35158 -6476
rect 35192 -6510 35211 -6476
rect 35139 -6566 35211 -6510
rect 35139 -6600 35158 -6566
rect 35192 -6600 35211 -6566
rect 35273 -5962 35967 -5903
rect 35273 -5996 35332 -5962
rect 35366 -5990 35422 -5962
rect 35394 -5996 35422 -5990
rect 35456 -5990 35512 -5962
rect 35456 -5996 35460 -5990
rect 35273 -6024 35360 -5996
rect 35394 -6024 35460 -5996
rect 35494 -5996 35512 -5990
rect 35546 -5990 35602 -5962
rect 35546 -5996 35560 -5990
rect 35494 -6024 35560 -5996
rect 35594 -5996 35602 -5990
rect 35636 -5990 35692 -5962
rect 35726 -5990 35782 -5962
rect 35816 -5990 35872 -5962
rect 35636 -5996 35660 -5990
rect 35726 -5996 35760 -5990
rect 35816 -5996 35860 -5990
rect 35906 -5996 35967 -5962
rect 35594 -6024 35660 -5996
rect 35694 -6024 35760 -5996
rect 35794 -6024 35860 -5996
rect 35894 -6024 35967 -5996
rect 35273 -6052 35967 -6024
rect 35273 -6086 35332 -6052
rect 35366 -6086 35422 -6052
rect 35456 -6086 35512 -6052
rect 35546 -6086 35602 -6052
rect 35636 -6086 35692 -6052
rect 35726 -6086 35782 -6052
rect 35816 -6086 35872 -6052
rect 35906 -6086 35967 -6052
rect 35273 -6090 35967 -6086
rect 35273 -6124 35360 -6090
rect 35394 -6124 35460 -6090
rect 35494 -6124 35560 -6090
rect 35594 -6124 35660 -6090
rect 35694 -6124 35760 -6090
rect 35794 -6124 35860 -6090
rect 35894 -6124 35967 -6090
rect 35273 -6142 35967 -6124
rect 35273 -6176 35332 -6142
rect 35366 -6176 35422 -6142
rect 35456 -6176 35512 -6142
rect 35546 -6176 35602 -6142
rect 35636 -6176 35692 -6142
rect 35726 -6176 35782 -6142
rect 35816 -6176 35872 -6142
rect 35906 -6176 35967 -6142
rect 35273 -6190 35967 -6176
rect 35273 -6224 35360 -6190
rect 35394 -6224 35460 -6190
rect 35494 -6224 35560 -6190
rect 35594 -6224 35660 -6190
rect 35694 -6224 35760 -6190
rect 35794 -6224 35860 -6190
rect 35894 -6224 35967 -6190
rect 35273 -6232 35967 -6224
rect 35273 -6266 35332 -6232
rect 35366 -6266 35422 -6232
rect 35456 -6266 35512 -6232
rect 35546 -6266 35602 -6232
rect 35636 -6266 35692 -6232
rect 35726 -6266 35782 -6232
rect 35816 -6266 35872 -6232
rect 35906 -6266 35967 -6232
rect 35273 -6290 35967 -6266
rect 35273 -6322 35360 -6290
rect 35394 -6322 35460 -6290
rect 35273 -6356 35332 -6322
rect 35394 -6324 35422 -6322
rect 35366 -6356 35422 -6324
rect 35456 -6324 35460 -6322
rect 35494 -6322 35560 -6290
rect 35494 -6324 35512 -6322
rect 35456 -6356 35512 -6324
rect 35546 -6324 35560 -6322
rect 35594 -6322 35660 -6290
rect 35694 -6322 35760 -6290
rect 35794 -6322 35860 -6290
rect 35894 -6322 35967 -6290
rect 35594 -6324 35602 -6322
rect 35546 -6356 35602 -6324
rect 35636 -6324 35660 -6322
rect 35726 -6324 35760 -6322
rect 35816 -6324 35860 -6322
rect 35636 -6356 35692 -6324
rect 35726 -6356 35782 -6324
rect 35816 -6356 35872 -6324
rect 35906 -6356 35967 -6322
rect 35273 -6390 35967 -6356
rect 35273 -6412 35360 -6390
rect 35394 -6412 35460 -6390
rect 35273 -6446 35332 -6412
rect 35394 -6424 35422 -6412
rect 35366 -6446 35422 -6424
rect 35456 -6424 35460 -6412
rect 35494 -6412 35560 -6390
rect 35494 -6424 35512 -6412
rect 35456 -6446 35512 -6424
rect 35546 -6424 35560 -6412
rect 35594 -6412 35660 -6390
rect 35694 -6412 35760 -6390
rect 35794 -6412 35860 -6390
rect 35894 -6412 35967 -6390
rect 35594 -6424 35602 -6412
rect 35546 -6446 35602 -6424
rect 35636 -6424 35660 -6412
rect 35726 -6424 35760 -6412
rect 35816 -6424 35860 -6412
rect 35636 -6446 35692 -6424
rect 35726 -6446 35782 -6424
rect 35816 -6446 35872 -6424
rect 35906 -6446 35967 -6412
rect 35273 -6490 35967 -6446
rect 35273 -6502 35360 -6490
rect 35394 -6502 35460 -6490
rect 35273 -6536 35332 -6502
rect 35394 -6524 35422 -6502
rect 35366 -6536 35422 -6524
rect 35456 -6524 35460 -6502
rect 35494 -6502 35560 -6490
rect 35494 -6524 35512 -6502
rect 35456 -6536 35512 -6524
rect 35546 -6524 35560 -6502
rect 35594 -6502 35660 -6490
rect 35694 -6502 35760 -6490
rect 35794 -6502 35860 -6490
rect 35894 -6502 35967 -6490
rect 35594 -6524 35602 -6502
rect 35546 -6536 35602 -6524
rect 35636 -6524 35660 -6502
rect 35726 -6524 35760 -6502
rect 35816 -6524 35860 -6502
rect 35636 -6536 35692 -6524
rect 35726 -6536 35782 -6524
rect 35816 -6536 35872 -6524
rect 35906 -6536 35967 -6502
rect 35273 -6597 35967 -6536
rect 36029 -5914 36048 -5880
rect 36082 -5914 36101 -5880
rect 36029 -5970 36101 -5914
rect 36029 -6004 36048 -5970
rect 36082 -6004 36101 -5970
rect 36029 -6060 36101 -6004
rect 36029 -6094 36048 -6060
rect 36082 -6094 36101 -6060
rect 36029 -6150 36101 -6094
rect 36029 -6184 36048 -6150
rect 36082 -6184 36101 -6150
rect 36029 -6240 36101 -6184
rect 36029 -6274 36048 -6240
rect 36082 -6274 36101 -6240
rect 36029 -6330 36101 -6274
rect 36029 -6364 36048 -6330
rect 36082 -6364 36101 -6330
rect 36029 -6420 36101 -6364
rect 36029 -6454 36048 -6420
rect 36082 -6454 36101 -6420
rect 36029 -6510 36101 -6454
rect 36029 -6544 36048 -6510
rect 36082 -6544 36101 -6510
rect 35139 -6659 35211 -6600
rect 36029 -6600 36101 -6544
rect 36029 -6634 36048 -6600
rect 36082 -6634 36101 -6600
rect 36029 -6659 36101 -6634
rect 35139 -6678 36101 -6659
rect 35139 -6712 35215 -6678
rect 35249 -6712 35305 -6678
rect 35339 -6712 35395 -6678
rect 35429 -6712 35485 -6678
rect 35519 -6712 35575 -6678
rect 35609 -6712 35665 -6678
rect 35699 -6712 35755 -6678
rect 35789 -6712 35845 -6678
rect 35879 -6712 35935 -6678
rect 35969 -6712 36101 -6678
rect 35139 -6731 36101 -6712
rect 36165 -5864 36198 -5850
rect 36232 -5864 36371 -5830
rect 36405 -5846 37558 -5830
rect 36405 -5850 36518 -5846
rect 36405 -5864 36435 -5850
rect 36165 -5920 36435 -5864
rect 36165 -5954 36198 -5920
rect 36232 -5954 36371 -5920
rect 36405 -5954 36435 -5920
rect 36165 -6010 36435 -5954
rect 36165 -6044 36198 -6010
rect 36232 -6044 36371 -6010
rect 36405 -6044 36435 -6010
rect 36165 -6100 36435 -6044
rect 36165 -6134 36198 -6100
rect 36232 -6134 36371 -6100
rect 36405 -6134 36435 -6100
rect 36165 -6190 36435 -6134
rect 36165 -6224 36198 -6190
rect 36232 -6224 36371 -6190
rect 36405 -6224 36435 -6190
rect 36165 -6280 36435 -6224
rect 36165 -6314 36198 -6280
rect 36232 -6314 36371 -6280
rect 36405 -6314 36435 -6280
rect 36165 -6370 36435 -6314
rect 36165 -6404 36198 -6370
rect 36232 -6404 36371 -6370
rect 36405 -6404 36435 -6370
rect 36165 -6460 36435 -6404
rect 36165 -6494 36198 -6460
rect 36232 -6494 36371 -6460
rect 36405 -6494 36435 -6460
rect 36165 -6550 36435 -6494
rect 36165 -6584 36198 -6550
rect 36232 -6584 36371 -6550
rect 36405 -6584 36435 -6550
rect 36165 -6640 36435 -6584
rect 36165 -6674 36198 -6640
rect 36232 -6674 36371 -6640
rect 36405 -6674 36435 -6640
rect 36165 -6730 36435 -6674
rect 34805 -6795 35075 -6764
rect 36165 -6764 36198 -6730
rect 36232 -6764 36371 -6730
rect 36405 -6764 36435 -6730
rect 36499 -5880 36518 -5850
rect 36552 -5850 37558 -5846
rect 36552 -5880 36571 -5850
rect 36499 -5936 36571 -5880
rect 37389 -5880 37461 -5850
rect 36499 -5970 36518 -5936
rect 36552 -5970 36571 -5936
rect 36499 -6026 36571 -5970
rect 36499 -6060 36518 -6026
rect 36552 -6060 36571 -6026
rect 36499 -6116 36571 -6060
rect 36499 -6150 36518 -6116
rect 36552 -6150 36571 -6116
rect 36499 -6206 36571 -6150
rect 36499 -6240 36518 -6206
rect 36552 -6240 36571 -6206
rect 36499 -6296 36571 -6240
rect 36499 -6330 36518 -6296
rect 36552 -6330 36571 -6296
rect 36499 -6386 36571 -6330
rect 36499 -6420 36518 -6386
rect 36552 -6420 36571 -6386
rect 36499 -6476 36571 -6420
rect 36499 -6510 36518 -6476
rect 36552 -6510 36571 -6476
rect 36499 -6566 36571 -6510
rect 36499 -6600 36518 -6566
rect 36552 -6600 36571 -6566
rect 36633 -5962 37327 -5903
rect 36633 -5996 36692 -5962
rect 36726 -5990 36782 -5962
rect 36754 -5996 36782 -5990
rect 36816 -5990 36872 -5962
rect 36816 -5996 36820 -5990
rect 36633 -6024 36720 -5996
rect 36754 -6024 36820 -5996
rect 36854 -5996 36872 -5990
rect 36906 -5990 36962 -5962
rect 36906 -5996 36920 -5990
rect 36854 -6024 36920 -5996
rect 36954 -5996 36962 -5990
rect 36996 -5990 37052 -5962
rect 37086 -5990 37142 -5962
rect 37176 -5990 37232 -5962
rect 36996 -5996 37020 -5990
rect 37086 -5996 37120 -5990
rect 37176 -5996 37220 -5990
rect 37266 -5996 37327 -5962
rect 36954 -6024 37020 -5996
rect 37054 -6024 37120 -5996
rect 37154 -6024 37220 -5996
rect 37254 -6024 37327 -5996
rect 36633 -6052 37327 -6024
rect 36633 -6086 36692 -6052
rect 36726 -6086 36782 -6052
rect 36816 -6086 36872 -6052
rect 36906 -6086 36962 -6052
rect 36996 -6086 37052 -6052
rect 37086 -6086 37142 -6052
rect 37176 -6086 37232 -6052
rect 37266 -6086 37327 -6052
rect 36633 -6090 37327 -6086
rect 36633 -6124 36720 -6090
rect 36754 -6124 36820 -6090
rect 36854 -6124 36920 -6090
rect 36954 -6124 37020 -6090
rect 37054 -6124 37120 -6090
rect 37154 -6124 37220 -6090
rect 37254 -6124 37327 -6090
rect 36633 -6142 37327 -6124
rect 36633 -6176 36692 -6142
rect 36726 -6176 36782 -6142
rect 36816 -6176 36872 -6142
rect 36906 -6176 36962 -6142
rect 36996 -6176 37052 -6142
rect 37086 -6176 37142 -6142
rect 37176 -6176 37232 -6142
rect 37266 -6176 37327 -6142
rect 36633 -6190 37327 -6176
rect 36633 -6224 36720 -6190
rect 36754 -6224 36820 -6190
rect 36854 -6224 36920 -6190
rect 36954 -6224 37020 -6190
rect 37054 -6224 37120 -6190
rect 37154 -6224 37220 -6190
rect 37254 -6224 37327 -6190
rect 36633 -6232 37327 -6224
rect 36633 -6266 36692 -6232
rect 36726 -6266 36782 -6232
rect 36816 -6266 36872 -6232
rect 36906 -6266 36962 -6232
rect 36996 -6266 37052 -6232
rect 37086 -6266 37142 -6232
rect 37176 -6266 37232 -6232
rect 37266 -6266 37327 -6232
rect 36633 -6290 37327 -6266
rect 36633 -6322 36720 -6290
rect 36754 -6322 36820 -6290
rect 36633 -6356 36692 -6322
rect 36754 -6324 36782 -6322
rect 36726 -6356 36782 -6324
rect 36816 -6324 36820 -6322
rect 36854 -6322 36920 -6290
rect 36854 -6324 36872 -6322
rect 36816 -6356 36872 -6324
rect 36906 -6324 36920 -6322
rect 36954 -6322 37020 -6290
rect 37054 -6322 37120 -6290
rect 37154 -6322 37220 -6290
rect 37254 -6322 37327 -6290
rect 36954 -6324 36962 -6322
rect 36906 -6356 36962 -6324
rect 36996 -6324 37020 -6322
rect 37086 -6324 37120 -6322
rect 37176 -6324 37220 -6322
rect 36996 -6356 37052 -6324
rect 37086 -6356 37142 -6324
rect 37176 -6356 37232 -6324
rect 37266 -6356 37327 -6322
rect 36633 -6390 37327 -6356
rect 36633 -6412 36720 -6390
rect 36754 -6412 36820 -6390
rect 36633 -6446 36692 -6412
rect 36754 -6424 36782 -6412
rect 36726 -6446 36782 -6424
rect 36816 -6424 36820 -6412
rect 36854 -6412 36920 -6390
rect 36854 -6424 36872 -6412
rect 36816 -6446 36872 -6424
rect 36906 -6424 36920 -6412
rect 36954 -6412 37020 -6390
rect 37054 -6412 37120 -6390
rect 37154 -6412 37220 -6390
rect 37254 -6412 37327 -6390
rect 36954 -6424 36962 -6412
rect 36906 -6446 36962 -6424
rect 36996 -6424 37020 -6412
rect 37086 -6424 37120 -6412
rect 37176 -6424 37220 -6412
rect 36996 -6446 37052 -6424
rect 37086 -6446 37142 -6424
rect 37176 -6446 37232 -6424
rect 37266 -6446 37327 -6412
rect 36633 -6490 37327 -6446
rect 36633 -6502 36720 -6490
rect 36754 -6502 36820 -6490
rect 36633 -6536 36692 -6502
rect 36754 -6524 36782 -6502
rect 36726 -6536 36782 -6524
rect 36816 -6524 36820 -6502
rect 36854 -6502 36920 -6490
rect 36854 -6524 36872 -6502
rect 36816 -6536 36872 -6524
rect 36906 -6524 36920 -6502
rect 36954 -6502 37020 -6490
rect 37054 -6502 37120 -6490
rect 37154 -6502 37220 -6490
rect 37254 -6502 37327 -6490
rect 36954 -6524 36962 -6502
rect 36906 -6536 36962 -6524
rect 36996 -6524 37020 -6502
rect 37086 -6524 37120 -6502
rect 37176 -6524 37220 -6502
rect 36996 -6536 37052 -6524
rect 37086 -6536 37142 -6524
rect 37176 -6536 37232 -6524
rect 37266 -6536 37327 -6502
rect 36633 -6597 37327 -6536
rect 37389 -5914 37408 -5880
rect 37442 -5914 37461 -5880
rect 37389 -5970 37461 -5914
rect 37389 -6004 37408 -5970
rect 37442 -6004 37461 -5970
rect 37389 -6060 37461 -6004
rect 37389 -6094 37408 -6060
rect 37442 -6094 37461 -6060
rect 37389 -6150 37461 -6094
rect 37389 -6184 37408 -6150
rect 37442 -6184 37461 -6150
rect 37389 -6240 37461 -6184
rect 37389 -6274 37408 -6240
rect 37442 -6274 37461 -6240
rect 37389 -6330 37461 -6274
rect 37389 -6364 37408 -6330
rect 37442 -6364 37461 -6330
rect 37389 -6420 37461 -6364
rect 37389 -6454 37408 -6420
rect 37442 -6454 37461 -6420
rect 37389 -6510 37461 -6454
rect 37389 -6544 37408 -6510
rect 37442 -6544 37461 -6510
rect 36499 -6659 36571 -6600
rect 37389 -6600 37461 -6544
rect 37389 -6634 37408 -6600
rect 37442 -6634 37461 -6600
rect 37389 -6659 37461 -6634
rect 36499 -6678 37461 -6659
rect 36499 -6712 36575 -6678
rect 36609 -6712 36665 -6678
rect 36699 -6712 36755 -6678
rect 36789 -6712 36845 -6678
rect 36879 -6712 36935 -6678
rect 36969 -6712 37025 -6678
rect 37059 -6712 37115 -6678
rect 37149 -6712 37205 -6678
rect 37239 -6712 37295 -6678
rect 37329 -6712 37461 -6678
rect 36499 -6731 37461 -6712
rect 37525 -5864 37558 -5850
rect 37592 -5850 37630 -5830
rect 37592 -5864 37624 -5850
rect 37525 -5920 37624 -5864
rect 37525 -5954 37558 -5920
rect 37592 -5954 37624 -5920
rect 37525 -6010 37624 -5954
rect 37525 -6044 37558 -6010
rect 37592 -6044 37624 -6010
rect 37525 -6100 37624 -6044
rect 37525 -6134 37558 -6100
rect 37592 -6134 37624 -6100
rect 37525 -6190 37624 -6134
rect 37525 -6224 37558 -6190
rect 37592 -6224 37624 -6190
rect 37525 -6280 37624 -6224
rect 37525 -6314 37558 -6280
rect 37592 -6314 37624 -6280
rect 37525 -6370 37624 -6314
rect 37525 -6404 37558 -6370
rect 37592 -6404 37624 -6370
rect 37525 -6460 37624 -6404
rect 37525 -6494 37558 -6460
rect 37592 -6494 37624 -6460
rect 37525 -6550 37624 -6494
rect 37525 -6584 37558 -6550
rect 37592 -6584 37624 -6550
rect 37525 -6640 37624 -6584
rect 37525 -6674 37558 -6640
rect 37592 -6674 37624 -6640
rect 37525 -6730 37624 -6674
rect 36165 -6795 36435 -6764
rect 37525 -6764 37558 -6730
rect 37592 -6764 37624 -6730
rect 37525 -6795 37624 -6764
rect 33616 -6826 37624 -6795
rect 33616 -6860 33674 -6826
rect 33708 -6860 33764 -6826
rect 33798 -6860 33854 -6826
rect 33888 -6860 33944 -6826
rect 33978 -6860 34034 -6826
rect 34068 -6860 34124 -6826
rect 34158 -6860 34214 -6826
rect 34248 -6860 34304 -6826
rect 34338 -6860 34394 -6826
rect 34428 -6860 34484 -6826
rect 34518 -6860 34574 -6826
rect 34608 -6860 34664 -6826
rect 34698 -6860 34754 -6826
rect 34788 -6860 35034 -6826
rect 35068 -6860 35124 -6826
rect 35158 -6860 35214 -6826
rect 35248 -6860 35304 -6826
rect 35338 -6860 35394 -6826
rect 35428 -6860 35484 -6826
rect 35518 -6860 35574 -6826
rect 35608 -6860 35664 -6826
rect 35698 -6860 35754 -6826
rect 35788 -6860 35844 -6826
rect 35878 -6860 35934 -6826
rect 35968 -6860 36024 -6826
rect 36058 -6860 36114 -6826
rect 36148 -6860 36394 -6826
rect 36428 -6860 36484 -6826
rect 36518 -6860 36574 -6826
rect 36608 -6860 36664 -6826
rect 36698 -6860 36754 -6826
rect 36788 -6860 36844 -6826
rect 36878 -6860 36934 -6826
rect 36968 -6860 37024 -6826
rect 37058 -6860 37114 -6826
rect 37148 -6860 37204 -6826
rect 37238 -6860 37294 -6826
rect 37328 -6860 37384 -6826
rect 37418 -6860 37474 -6826
rect 37508 -6860 37624 -6826
rect 33616 -6894 37624 -6860
rect 34900 -6960 34980 -6894
rect 36260 -6960 36340 -6894
rect 33610 -6999 37630 -6960
rect 33610 -7033 33674 -6999
rect 33708 -7033 33764 -6999
rect 33798 -7033 33854 -6999
rect 33888 -7033 33944 -6999
rect 33978 -7033 34034 -6999
rect 34068 -7033 34124 -6999
rect 34158 -7033 34214 -6999
rect 34248 -7033 34304 -6999
rect 34338 -7033 34394 -6999
rect 34428 -7033 34484 -6999
rect 34518 -7033 34574 -6999
rect 34608 -7033 34664 -6999
rect 34698 -7033 34754 -6999
rect 34788 -7033 35034 -6999
rect 35068 -7033 35124 -6999
rect 35158 -7033 35214 -6999
rect 35248 -7033 35304 -6999
rect 35338 -7033 35394 -6999
rect 35428 -7033 35484 -6999
rect 35518 -7033 35574 -6999
rect 35608 -7033 35664 -6999
rect 35698 -7033 35754 -6999
rect 35788 -7033 35844 -6999
rect 35878 -7033 35934 -6999
rect 35968 -7033 36024 -6999
rect 36058 -7033 36114 -6999
rect 36148 -7033 36394 -6999
rect 36428 -7033 36484 -6999
rect 36518 -7033 36574 -6999
rect 36608 -7033 36664 -6999
rect 36698 -7033 36754 -6999
rect 36788 -7033 36844 -6999
rect 36878 -7033 36934 -6999
rect 36968 -7033 37024 -6999
rect 37058 -7033 37114 -6999
rect 37148 -7033 37204 -6999
rect 37238 -7033 37294 -6999
rect 37328 -7033 37384 -6999
rect 37418 -7033 37474 -6999
rect 37508 -7033 37630 -6999
rect 33610 -7100 37630 -7033
rect 33610 -7134 33651 -7100
rect 33685 -7134 34838 -7100
rect 34872 -7134 35011 -7100
rect 35045 -7134 36198 -7100
rect 36232 -7134 36371 -7100
rect 36405 -7134 37558 -7100
rect 37592 -7134 37630 -7100
rect 33610 -7148 37630 -7134
rect 33610 -7182 33874 -7148
rect 33908 -7182 33964 -7148
rect 33998 -7182 34054 -7148
rect 34088 -7182 34144 -7148
rect 34178 -7182 34234 -7148
rect 34268 -7182 34324 -7148
rect 34358 -7182 34414 -7148
rect 34448 -7182 34504 -7148
rect 34538 -7182 34594 -7148
rect 34628 -7182 35234 -7148
rect 35268 -7182 35324 -7148
rect 35358 -7182 35414 -7148
rect 35448 -7182 35504 -7148
rect 35538 -7182 35594 -7148
rect 35628 -7182 35684 -7148
rect 35718 -7182 35774 -7148
rect 35808 -7182 35864 -7148
rect 35898 -7182 35954 -7148
rect 35988 -7182 36594 -7148
rect 36628 -7182 36684 -7148
rect 36718 -7182 36774 -7148
rect 36808 -7182 36864 -7148
rect 36898 -7182 36954 -7148
rect 36988 -7182 37044 -7148
rect 37078 -7182 37134 -7148
rect 37168 -7182 37224 -7148
rect 37258 -7182 37314 -7148
rect 37348 -7182 37630 -7148
rect 33610 -7190 37630 -7182
rect 33610 -7210 33651 -7190
rect 33616 -7224 33651 -7210
rect 33685 -7206 34838 -7190
rect 33685 -7210 33798 -7206
rect 33685 -7224 33715 -7210
rect 33616 -7280 33715 -7224
rect 33616 -7314 33651 -7280
rect 33685 -7314 33715 -7280
rect 33616 -7370 33715 -7314
rect 33616 -7404 33651 -7370
rect 33685 -7404 33715 -7370
rect 33616 -7460 33715 -7404
rect 33616 -7494 33651 -7460
rect 33685 -7494 33715 -7460
rect 33616 -7550 33715 -7494
rect 33616 -7584 33651 -7550
rect 33685 -7584 33715 -7550
rect 33616 -7640 33715 -7584
rect 33616 -7674 33651 -7640
rect 33685 -7674 33715 -7640
rect 33616 -7730 33715 -7674
rect 33616 -7764 33651 -7730
rect 33685 -7764 33715 -7730
rect 33616 -7820 33715 -7764
rect 33616 -7854 33651 -7820
rect 33685 -7854 33715 -7820
rect 33616 -7910 33715 -7854
rect 33616 -7944 33651 -7910
rect 33685 -7944 33715 -7910
rect 33616 -8000 33715 -7944
rect 33616 -8034 33651 -8000
rect 33685 -8034 33715 -8000
rect 33616 -8090 33715 -8034
rect 33616 -8124 33651 -8090
rect 33685 -8124 33715 -8090
rect 33779 -7240 33798 -7210
rect 33832 -7210 34838 -7206
rect 33832 -7240 33851 -7210
rect 33779 -7296 33851 -7240
rect 34669 -7240 34741 -7210
rect 33779 -7330 33798 -7296
rect 33832 -7330 33851 -7296
rect 33779 -7386 33851 -7330
rect 33779 -7420 33798 -7386
rect 33832 -7420 33851 -7386
rect 33779 -7476 33851 -7420
rect 33779 -7510 33798 -7476
rect 33832 -7510 33851 -7476
rect 33779 -7566 33851 -7510
rect 33779 -7600 33798 -7566
rect 33832 -7600 33851 -7566
rect 33779 -7656 33851 -7600
rect 33779 -7690 33798 -7656
rect 33832 -7690 33851 -7656
rect 33779 -7746 33851 -7690
rect 33779 -7780 33798 -7746
rect 33832 -7780 33851 -7746
rect 33779 -7836 33851 -7780
rect 33779 -7870 33798 -7836
rect 33832 -7870 33851 -7836
rect 33779 -7926 33851 -7870
rect 33779 -7960 33798 -7926
rect 33832 -7960 33851 -7926
rect 33913 -7322 34607 -7263
rect 33913 -7356 33972 -7322
rect 34006 -7350 34062 -7322
rect 34034 -7356 34062 -7350
rect 34096 -7350 34152 -7322
rect 34096 -7356 34100 -7350
rect 33913 -7384 34000 -7356
rect 34034 -7384 34100 -7356
rect 34134 -7356 34152 -7350
rect 34186 -7350 34242 -7322
rect 34186 -7356 34200 -7350
rect 34134 -7384 34200 -7356
rect 34234 -7356 34242 -7350
rect 34276 -7350 34332 -7322
rect 34366 -7350 34422 -7322
rect 34456 -7350 34512 -7322
rect 34276 -7356 34300 -7350
rect 34366 -7356 34400 -7350
rect 34456 -7356 34500 -7350
rect 34546 -7356 34607 -7322
rect 34234 -7384 34300 -7356
rect 34334 -7384 34400 -7356
rect 34434 -7384 34500 -7356
rect 34534 -7384 34607 -7356
rect 33913 -7412 34607 -7384
rect 33913 -7446 33972 -7412
rect 34006 -7446 34062 -7412
rect 34096 -7446 34152 -7412
rect 34186 -7446 34242 -7412
rect 34276 -7446 34332 -7412
rect 34366 -7446 34422 -7412
rect 34456 -7446 34512 -7412
rect 34546 -7446 34607 -7412
rect 33913 -7450 34607 -7446
rect 33913 -7484 34000 -7450
rect 34034 -7484 34100 -7450
rect 34134 -7484 34200 -7450
rect 34234 -7484 34300 -7450
rect 34334 -7484 34400 -7450
rect 34434 -7484 34500 -7450
rect 34534 -7484 34607 -7450
rect 33913 -7502 34607 -7484
rect 33913 -7536 33972 -7502
rect 34006 -7536 34062 -7502
rect 34096 -7536 34152 -7502
rect 34186 -7536 34242 -7502
rect 34276 -7536 34332 -7502
rect 34366 -7536 34422 -7502
rect 34456 -7536 34512 -7502
rect 34546 -7536 34607 -7502
rect 33913 -7550 34607 -7536
rect 33913 -7584 34000 -7550
rect 34034 -7584 34100 -7550
rect 34134 -7584 34200 -7550
rect 34234 -7584 34300 -7550
rect 34334 -7584 34400 -7550
rect 34434 -7584 34500 -7550
rect 34534 -7584 34607 -7550
rect 33913 -7592 34607 -7584
rect 33913 -7626 33972 -7592
rect 34006 -7626 34062 -7592
rect 34096 -7626 34152 -7592
rect 34186 -7626 34242 -7592
rect 34276 -7626 34332 -7592
rect 34366 -7626 34422 -7592
rect 34456 -7626 34512 -7592
rect 34546 -7626 34607 -7592
rect 33913 -7650 34607 -7626
rect 33913 -7682 34000 -7650
rect 34034 -7682 34100 -7650
rect 33913 -7716 33972 -7682
rect 34034 -7684 34062 -7682
rect 34006 -7716 34062 -7684
rect 34096 -7684 34100 -7682
rect 34134 -7682 34200 -7650
rect 34134 -7684 34152 -7682
rect 34096 -7716 34152 -7684
rect 34186 -7684 34200 -7682
rect 34234 -7682 34300 -7650
rect 34334 -7682 34400 -7650
rect 34434 -7682 34500 -7650
rect 34534 -7682 34607 -7650
rect 34234 -7684 34242 -7682
rect 34186 -7716 34242 -7684
rect 34276 -7684 34300 -7682
rect 34366 -7684 34400 -7682
rect 34456 -7684 34500 -7682
rect 34276 -7716 34332 -7684
rect 34366 -7716 34422 -7684
rect 34456 -7716 34512 -7684
rect 34546 -7716 34607 -7682
rect 33913 -7750 34607 -7716
rect 33913 -7772 34000 -7750
rect 34034 -7772 34100 -7750
rect 33913 -7806 33972 -7772
rect 34034 -7784 34062 -7772
rect 34006 -7806 34062 -7784
rect 34096 -7784 34100 -7772
rect 34134 -7772 34200 -7750
rect 34134 -7784 34152 -7772
rect 34096 -7806 34152 -7784
rect 34186 -7784 34200 -7772
rect 34234 -7772 34300 -7750
rect 34334 -7772 34400 -7750
rect 34434 -7772 34500 -7750
rect 34534 -7772 34607 -7750
rect 34234 -7784 34242 -7772
rect 34186 -7806 34242 -7784
rect 34276 -7784 34300 -7772
rect 34366 -7784 34400 -7772
rect 34456 -7784 34500 -7772
rect 34276 -7806 34332 -7784
rect 34366 -7806 34422 -7784
rect 34456 -7806 34512 -7784
rect 34546 -7806 34607 -7772
rect 33913 -7850 34607 -7806
rect 33913 -7862 34000 -7850
rect 34034 -7862 34100 -7850
rect 33913 -7896 33972 -7862
rect 34034 -7884 34062 -7862
rect 34006 -7896 34062 -7884
rect 34096 -7884 34100 -7862
rect 34134 -7862 34200 -7850
rect 34134 -7884 34152 -7862
rect 34096 -7896 34152 -7884
rect 34186 -7884 34200 -7862
rect 34234 -7862 34300 -7850
rect 34334 -7862 34400 -7850
rect 34434 -7862 34500 -7850
rect 34534 -7862 34607 -7850
rect 34234 -7884 34242 -7862
rect 34186 -7896 34242 -7884
rect 34276 -7884 34300 -7862
rect 34366 -7884 34400 -7862
rect 34456 -7884 34500 -7862
rect 34276 -7896 34332 -7884
rect 34366 -7896 34422 -7884
rect 34456 -7896 34512 -7884
rect 34546 -7896 34607 -7862
rect 33913 -7957 34607 -7896
rect 34669 -7274 34688 -7240
rect 34722 -7274 34741 -7240
rect 34669 -7330 34741 -7274
rect 34669 -7364 34688 -7330
rect 34722 -7364 34741 -7330
rect 34669 -7420 34741 -7364
rect 34669 -7454 34688 -7420
rect 34722 -7454 34741 -7420
rect 34669 -7510 34741 -7454
rect 34669 -7544 34688 -7510
rect 34722 -7544 34741 -7510
rect 34669 -7600 34741 -7544
rect 34669 -7634 34688 -7600
rect 34722 -7634 34741 -7600
rect 34669 -7690 34741 -7634
rect 34669 -7724 34688 -7690
rect 34722 -7724 34741 -7690
rect 34669 -7780 34741 -7724
rect 34669 -7814 34688 -7780
rect 34722 -7814 34741 -7780
rect 34669 -7870 34741 -7814
rect 34669 -7904 34688 -7870
rect 34722 -7904 34741 -7870
rect 33779 -8019 33851 -7960
rect 34669 -7960 34741 -7904
rect 34669 -7994 34688 -7960
rect 34722 -7994 34741 -7960
rect 34669 -8019 34741 -7994
rect 33779 -8038 34741 -8019
rect 33779 -8072 33855 -8038
rect 33889 -8072 33945 -8038
rect 33979 -8072 34035 -8038
rect 34069 -8072 34125 -8038
rect 34159 -8072 34215 -8038
rect 34249 -8072 34305 -8038
rect 34339 -8072 34395 -8038
rect 34429 -8072 34485 -8038
rect 34519 -8072 34575 -8038
rect 34609 -8072 34741 -8038
rect 33779 -8091 34741 -8072
rect 34805 -7224 34838 -7210
rect 34872 -7224 35011 -7190
rect 35045 -7206 36198 -7190
rect 35045 -7210 35158 -7206
rect 35045 -7224 35075 -7210
rect 34805 -7280 35075 -7224
rect 34805 -7314 34838 -7280
rect 34872 -7314 35011 -7280
rect 35045 -7314 35075 -7280
rect 34805 -7370 35075 -7314
rect 34805 -7404 34838 -7370
rect 34872 -7404 35011 -7370
rect 35045 -7404 35075 -7370
rect 34805 -7460 35075 -7404
rect 34805 -7494 34838 -7460
rect 34872 -7494 35011 -7460
rect 35045 -7494 35075 -7460
rect 34805 -7550 35075 -7494
rect 34805 -7584 34838 -7550
rect 34872 -7584 35011 -7550
rect 35045 -7584 35075 -7550
rect 34805 -7640 35075 -7584
rect 34805 -7674 34838 -7640
rect 34872 -7674 35011 -7640
rect 35045 -7674 35075 -7640
rect 34805 -7730 35075 -7674
rect 34805 -7764 34838 -7730
rect 34872 -7764 35011 -7730
rect 35045 -7764 35075 -7730
rect 34805 -7820 35075 -7764
rect 34805 -7854 34838 -7820
rect 34872 -7854 35011 -7820
rect 35045 -7854 35075 -7820
rect 34805 -7910 35075 -7854
rect 34805 -7944 34838 -7910
rect 34872 -7944 35011 -7910
rect 35045 -7944 35075 -7910
rect 34805 -8000 35075 -7944
rect 34805 -8034 34838 -8000
rect 34872 -8034 35011 -8000
rect 35045 -8034 35075 -8000
rect 34805 -8090 35075 -8034
rect 33616 -8155 33715 -8124
rect 34805 -8124 34838 -8090
rect 34872 -8124 35011 -8090
rect 35045 -8124 35075 -8090
rect 35139 -7240 35158 -7210
rect 35192 -7210 36198 -7206
rect 35192 -7240 35211 -7210
rect 35139 -7296 35211 -7240
rect 36029 -7240 36101 -7210
rect 35139 -7330 35158 -7296
rect 35192 -7330 35211 -7296
rect 35139 -7386 35211 -7330
rect 35139 -7420 35158 -7386
rect 35192 -7420 35211 -7386
rect 35139 -7476 35211 -7420
rect 35139 -7510 35158 -7476
rect 35192 -7510 35211 -7476
rect 35139 -7566 35211 -7510
rect 35139 -7600 35158 -7566
rect 35192 -7600 35211 -7566
rect 35139 -7656 35211 -7600
rect 35139 -7690 35158 -7656
rect 35192 -7690 35211 -7656
rect 35139 -7746 35211 -7690
rect 35139 -7780 35158 -7746
rect 35192 -7780 35211 -7746
rect 35139 -7836 35211 -7780
rect 35139 -7870 35158 -7836
rect 35192 -7870 35211 -7836
rect 35139 -7926 35211 -7870
rect 35139 -7960 35158 -7926
rect 35192 -7960 35211 -7926
rect 35273 -7322 35967 -7263
rect 35273 -7356 35332 -7322
rect 35366 -7350 35422 -7322
rect 35394 -7356 35422 -7350
rect 35456 -7350 35512 -7322
rect 35456 -7356 35460 -7350
rect 35273 -7384 35360 -7356
rect 35394 -7384 35460 -7356
rect 35494 -7356 35512 -7350
rect 35546 -7350 35602 -7322
rect 35546 -7356 35560 -7350
rect 35494 -7384 35560 -7356
rect 35594 -7356 35602 -7350
rect 35636 -7350 35692 -7322
rect 35726 -7350 35782 -7322
rect 35816 -7350 35872 -7322
rect 35636 -7356 35660 -7350
rect 35726 -7356 35760 -7350
rect 35816 -7356 35860 -7350
rect 35906 -7356 35967 -7322
rect 35594 -7384 35660 -7356
rect 35694 -7384 35760 -7356
rect 35794 -7384 35860 -7356
rect 35894 -7384 35967 -7356
rect 35273 -7412 35967 -7384
rect 35273 -7446 35332 -7412
rect 35366 -7446 35422 -7412
rect 35456 -7446 35512 -7412
rect 35546 -7446 35602 -7412
rect 35636 -7446 35692 -7412
rect 35726 -7446 35782 -7412
rect 35816 -7446 35872 -7412
rect 35906 -7446 35967 -7412
rect 35273 -7450 35967 -7446
rect 35273 -7484 35360 -7450
rect 35394 -7484 35460 -7450
rect 35494 -7484 35560 -7450
rect 35594 -7484 35660 -7450
rect 35694 -7484 35760 -7450
rect 35794 -7484 35860 -7450
rect 35894 -7484 35967 -7450
rect 35273 -7502 35967 -7484
rect 35273 -7536 35332 -7502
rect 35366 -7536 35422 -7502
rect 35456 -7536 35512 -7502
rect 35546 -7536 35602 -7502
rect 35636 -7536 35692 -7502
rect 35726 -7536 35782 -7502
rect 35816 -7536 35872 -7502
rect 35906 -7536 35967 -7502
rect 35273 -7550 35967 -7536
rect 35273 -7584 35360 -7550
rect 35394 -7584 35460 -7550
rect 35494 -7584 35560 -7550
rect 35594 -7584 35660 -7550
rect 35694 -7584 35760 -7550
rect 35794 -7584 35860 -7550
rect 35894 -7584 35967 -7550
rect 35273 -7592 35967 -7584
rect 35273 -7626 35332 -7592
rect 35366 -7626 35422 -7592
rect 35456 -7626 35512 -7592
rect 35546 -7626 35602 -7592
rect 35636 -7626 35692 -7592
rect 35726 -7626 35782 -7592
rect 35816 -7626 35872 -7592
rect 35906 -7626 35967 -7592
rect 35273 -7650 35967 -7626
rect 35273 -7682 35360 -7650
rect 35394 -7682 35460 -7650
rect 35273 -7716 35332 -7682
rect 35394 -7684 35422 -7682
rect 35366 -7716 35422 -7684
rect 35456 -7684 35460 -7682
rect 35494 -7682 35560 -7650
rect 35494 -7684 35512 -7682
rect 35456 -7716 35512 -7684
rect 35546 -7684 35560 -7682
rect 35594 -7682 35660 -7650
rect 35694 -7682 35760 -7650
rect 35794 -7682 35860 -7650
rect 35894 -7682 35967 -7650
rect 35594 -7684 35602 -7682
rect 35546 -7716 35602 -7684
rect 35636 -7684 35660 -7682
rect 35726 -7684 35760 -7682
rect 35816 -7684 35860 -7682
rect 35636 -7716 35692 -7684
rect 35726 -7716 35782 -7684
rect 35816 -7716 35872 -7684
rect 35906 -7716 35967 -7682
rect 35273 -7750 35967 -7716
rect 35273 -7772 35360 -7750
rect 35394 -7772 35460 -7750
rect 35273 -7806 35332 -7772
rect 35394 -7784 35422 -7772
rect 35366 -7806 35422 -7784
rect 35456 -7784 35460 -7772
rect 35494 -7772 35560 -7750
rect 35494 -7784 35512 -7772
rect 35456 -7806 35512 -7784
rect 35546 -7784 35560 -7772
rect 35594 -7772 35660 -7750
rect 35694 -7772 35760 -7750
rect 35794 -7772 35860 -7750
rect 35894 -7772 35967 -7750
rect 35594 -7784 35602 -7772
rect 35546 -7806 35602 -7784
rect 35636 -7784 35660 -7772
rect 35726 -7784 35760 -7772
rect 35816 -7784 35860 -7772
rect 35636 -7806 35692 -7784
rect 35726 -7806 35782 -7784
rect 35816 -7806 35872 -7784
rect 35906 -7806 35967 -7772
rect 35273 -7850 35967 -7806
rect 35273 -7862 35360 -7850
rect 35394 -7862 35460 -7850
rect 35273 -7896 35332 -7862
rect 35394 -7884 35422 -7862
rect 35366 -7896 35422 -7884
rect 35456 -7884 35460 -7862
rect 35494 -7862 35560 -7850
rect 35494 -7884 35512 -7862
rect 35456 -7896 35512 -7884
rect 35546 -7884 35560 -7862
rect 35594 -7862 35660 -7850
rect 35694 -7862 35760 -7850
rect 35794 -7862 35860 -7850
rect 35894 -7862 35967 -7850
rect 35594 -7884 35602 -7862
rect 35546 -7896 35602 -7884
rect 35636 -7884 35660 -7862
rect 35726 -7884 35760 -7862
rect 35816 -7884 35860 -7862
rect 35636 -7896 35692 -7884
rect 35726 -7896 35782 -7884
rect 35816 -7896 35872 -7884
rect 35906 -7896 35967 -7862
rect 35273 -7957 35967 -7896
rect 36029 -7274 36048 -7240
rect 36082 -7274 36101 -7240
rect 36029 -7330 36101 -7274
rect 36029 -7364 36048 -7330
rect 36082 -7364 36101 -7330
rect 36029 -7420 36101 -7364
rect 36029 -7454 36048 -7420
rect 36082 -7454 36101 -7420
rect 36029 -7510 36101 -7454
rect 36029 -7544 36048 -7510
rect 36082 -7544 36101 -7510
rect 36029 -7600 36101 -7544
rect 36029 -7634 36048 -7600
rect 36082 -7634 36101 -7600
rect 36029 -7690 36101 -7634
rect 36029 -7724 36048 -7690
rect 36082 -7724 36101 -7690
rect 36029 -7780 36101 -7724
rect 36029 -7814 36048 -7780
rect 36082 -7814 36101 -7780
rect 36029 -7870 36101 -7814
rect 36029 -7904 36048 -7870
rect 36082 -7904 36101 -7870
rect 35139 -8019 35211 -7960
rect 36029 -7960 36101 -7904
rect 36029 -7994 36048 -7960
rect 36082 -7994 36101 -7960
rect 36029 -8019 36101 -7994
rect 35139 -8038 36101 -8019
rect 35139 -8072 35215 -8038
rect 35249 -8072 35305 -8038
rect 35339 -8072 35395 -8038
rect 35429 -8072 35485 -8038
rect 35519 -8072 35575 -8038
rect 35609 -8072 35665 -8038
rect 35699 -8072 35755 -8038
rect 35789 -8072 35845 -8038
rect 35879 -8072 35935 -8038
rect 35969 -8072 36101 -8038
rect 35139 -8091 36101 -8072
rect 36165 -7224 36198 -7210
rect 36232 -7224 36371 -7190
rect 36405 -7206 37558 -7190
rect 36405 -7210 36518 -7206
rect 36405 -7224 36435 -7210
rect 36165 -7280 36435 -7224
rect 36165 -7314 36198 -7280
rect 36232 -7314 36371 -7280
rect 36405 -7314 36435 -7280
rect 36165 -7370 36435 -7314
rect 36165 -7404 36198 -7370
rect 36232 -7404 36371 -7370
rect 36405 -7404 36435 -7370
rect 36165 -7460 36435 -7404
rect 36165 -7494 36198 -7460
rect 36232 -7494 36371 -7460
rect 36405 -7494 36435 -7460
rect 36165 -7550 36435 -7494
rect 36165 -7584 36198 -7550
rect 36232 -7584 36371 -7550
rect 36405 -7584 36435 -7550
rect 36165 -7640 36435 -7584
rect 36165 -7674 36198 -7640
rect 36232 -7674 36371 -7640
rect 36405 -7674 36435 -7640
rect 36165 -7730 36435 -7674
rect 36165 -7764 36198 -7730
rect 36232 -7764 36371 -7730
rect 36405 -7764 36435 -7730
rect 36165 -7820 36435 -7764
rect 36165 -7854 36198 -7820
rect 36232 -7854 36371 -7820
rect 36405 -7854 36435 -7820
rect 36165 -7910 36435 -7854
rect 36165 -7944 36198 -7910
rect 36232 -7944 36371 -7910
rect 36405 -7944 36435 -7910
rect 36165 -8000 36435 -7944
rect 36165 -8034 36198 -8000
rect 36232 -8034 36371 -8000
rect 36405 -8034 36435 -8000
rect 36165 -8090 36435 -8034
rect 34805 -8155 35075 -8124
rect 36165 -8124 36198 -8090
rect 36232 -8124 36371 -8090
rect 36405 -8124 36435 -8090
rect 36499 -7240 36518 -7210
rect 36552 -7210 37558 -7206
rect 36552 -7240 36571 -7210
rect 36499 -7296 36571 -7240
rect 37389 -7240 37461 -7210
rect 36499 -7330 36518 -7296
rect 36552 -7330 36571 -7296
rect 36499 -7386 36571 -7330
rect 36499 -7420 36518 -7386
rect 36552 -7420 36571 -7386
rect 36499 -7476 36571 -7420
rect 36499 -7510 36518 -7476
rect 36552 -7510 36571 -7476
rect 36499 -7566 36571 -7510
rect 36499 -7600 36518 -7566
rect 36552 -7600 36571 -7566
rect 36499 -7656 36571 -7600
rect 36499 -7690 36518 -7656
rect 36552 -7690 36571 -7656
rect 36499 -7746 36571 -7690
rect 36499 -7780 36518 -7746
rect 36552 -7780 36571 -7746
rect 36499 -7836 36571 -7780
rect 36499 -7870 36518 -7836
rect 36552 -7870 36571 -7836
rect 36499 -7926 36571 -7870
rect 36499 -7960 36518 -7926
rect 36552 -7960 36571 -7926
rect 36633 -7322 37327 -7263
rect 36633 -7356 36692 -7322
rect 36726 -7350 36782 -7322
rect 36754 -7356 36782 -7350
rect 36816 -7350 36872 -7322
rect 36816 -7356 36820 -7350
rect 36633 -7384 36720 -7356
rect 36754 -7384 36820 -7356
rect 36854 -7356 36872 -7350
rect 36906 -7350 36962 -7322
rect 36906 -7356 36920 -7350
rect 36854 -7384 36920 -7356
rect 36954 -7356 36962 -7350
rect 36996 -7350 37052 -7322
rect 37086 -7350 37142 -7322
rect 37176 -7350 37232 -7322
rect 36996 -7356 37020 -7350
rect 37086 -7356 37120 -7350
rect 37176 -7356 37220 -7350
rect 37266 -7356 37327 -7322
rect 36954 -7384 37020 -7356
rect 37054 -7384 37120 -7356
rect 37154 -7384 37220 -7356
rect 37254 -7384 37327 -7356
rect 36633 -7412 37327 -7384
rect 36633 -7446 36692 -7412
rect 36726 -7446 36782 -7412
rect 36816 -7446 36872 -7412
rect 36906 -7446 36962 -7412
rect 36996 -7446 37052 -7412
rect 37086 -7446 37142 -7412
rect 37176 -7446 37232 -7412
rect 37266 -7446 37327 -7412
rect 36633 -7450 37327 -7446
rect 36633 -7484 36720 -7450
rect 36754 -7484 36820 -7450
rect 36854 -7484 36920 -7450
rect 36954 -7484 37020 -7450
rect 37054 -7484 37120 -7450
rect 37154 -7484 37220 -7450
rect 37254 -7484 37327 -7450
rect 36633 -7502 37327 -7484
rect 36633 -7536 36692 -7502
rect 36726 -7536 36782 -7502
rect 36816 -7536 36872 -7502
rect 36906 -7536 36962 -7502
rect 36996 -7536 37052 -7502
rect 37086 -7536 37142 -7502
rect 37176 -7536 37232 -7502
rect 37266 -7536 37327 -7502
rect 36633 -7550 37327 -7536
rect 36633 -7584 36720 -7550
rect 36754 -7584 36820 -7550
rect 36854 -7584 36920 -7550
rect 36954 -7584 37020 -7550
rect 37054 -7584 37120 -7550
rect 37154 -7584 37220 -7550
rect 37254 -7584 37327 -7550
rect 36633 -7592 37327 -7584
rect 36633 -7626 36692 -7592
rect 36726 -7626 36782 -7592
rect 36816 -7626 36872 -7592
rect 36906 -7626 36962 -7592
rect 36996 -7626 37052 -7592
rect 37086 -7626 37142 -7592
rect 37176 -7626 37232 -7592
rect 37266 -7626 37327 -7592
rect 36633 -7650 37327 -7626
rect 36633 -7682 36720 -7650
rect 36754 -7682 36820 -7650
rect 36633 -7716 36692 -7682
rect 36754 -7684 36782 -7682
rect 36726 -7716 36782 -7684
rect 36816 -7684 36820 -7682
rect 36854 -7682 36920 -7650
rect 36854 -7684 36872 -7682
rect 36816 -7716 36872 -7684
rect 36906 -7684 36920 -7682
rect 36954 -7682 37020 -7650
rect 37054 -7682 37120 -7650
rect 37154 -7682 37220 -7650
rect 37254 -7682 37327 -7650
rect 36954 -7684 36962 -7682
rect 36906 -7716 36962 -7684
rect 36996 -7684 37020 -7682
rect 37086 -7684 37120 -7682
rect 37176 -7684 37220 -7682
rect 36996 -7716 37052 -7684
rect 37086 -7716 37142 -7684
rect 37176 -7716 37232 -7684
rect 37266 -7716 37327 -7682
rect 36633 -7750 37327 -7716
rect 36633 -7772 36720 -7750
rect 36754 -7772 36820 -7750
rect 36633 -7806 36692 -7772
rect 36754 -7784 36782 -7772
rect 36726 -7806 36782 -7784
rect 36816 -7784 36820 -7772
rect 36854 -7772 36920 -7750
rect 36854 -7784 36872 -7772
rect 36816 -7806 36872 -7784
rect 36906 -7784 36920 -7772
rect 36954 -7772 37020 -7750
rect 37054 -7772 37120 -7750
rect 37154 -7772 37220 -7750
rect 37254 -7772 37327 -7750
rect 36954 -7784 36962 -7772
rect 36906 -7806 36962 -7784
rect 36996 -7784 37020 -7772
rect 37086 -7784 37120 -7772
rect 37176 -7784 37220 -7772
rect 36996 -7806 37052 -7784
rect 37086 -7806 37142 -7784
rect 37176 -7806 37232 -7784
rect 37266 -7806 37327 -7772
rect 36633 -7850 37327 -7806
rect 36633 -7862 36720 -7850
rect 36754 -7862 36820 -7850
rect 36633 -7896 36692 -7862
rect 36754 -7884 36782 -7862
rect 36726 -7896 36782 -7884
rect 36816 -7884 36820 -7862
rect 36854 -7862 36920 -7850
rect 36854 -7884 36872 -7862
rect 36816 -7896 36872 -7884
rect 36906 -7884 36920 -7862
rect 36954 -7862 37020 -7850
rect 37054 -7862 37120 -7850
rect 37154 -7862 37220 -7850
rect 37254 -7862 37327 -7850
rect 36954 -7884 36962 -7862
rect 36906 -7896 36962 -7884
rect 36996 -7884 37020 -7862
rect 37086 -7884 37120 -7862
rect 37176 -7884 37220 -7862
rect 36996 -7896 37052 -7884
rect 37086 -7896 37142 -7884
rect 37176 -7896 37232 -7884
rect 37266 -7896 37327 -7862
rect 36633 -7957 37327 -7896
rect 37389 -7274 37408 -7240
rect 37442 -7274 37461 -7240
rect 37389 -7330 37461 -7274
rect 37389 -7364 37408 -7330
rect 37442 -7364 37461 -7330
rect 37389 -7420 37461 -7364
rect 37389 -7454 37408 -7420
rect 37442 -7454 37461 -7420
rect 37389 -7510 37461 -7454
rect 37389 -7544 37408 -7510
rect 37442 -7544 37461 -7510
rect 37389 -7600 37461 -7544
rect 37389 -7634 37408 -7600
rect 37442 -7634 37461 -7600
rect 37389 -7690 37461 -7634
rect 37389 -7724 37408 -7690
rect 37442 -7724 37461 -7690
rect 37389 -7780 37461 -7724
rect 37389 -7814 37408 -7780
rect 37442 -7814 37461 -7780
rect 37389 -7870 37461 -7814
rect 37389 -7904 37408 -7870
rect 37442 -7904 37461 -7870
rect 36499 -8019 36571 -7960
rect 37389 -7960 37461 -7904
rect 37389 -7994 37408 -7960
rect 37442 -7994 37461 -7960
rect 37389 -8019 37461 -7994
rect 36499 -8038 37461 -8019
rect 36499 -8072 36575 -8038
rect 36609 -8072 36665 -8038
rect 36699 -8072 36755 -8038
rect 36789 -8072 36845 -8038
rect 36879 -8072 36935 -8038
rect 36969 -8072 37025 -8038
rect 37059 -8072 37115 -8038
rect 37149 -8072 37205 -8038
rect 37239 -8072 37295 -8038
rect 37329 -8072 37461 -8038
rect 36499 -8091 37461 -8072
rect 37525 -7224 37558 -7210
rect 37592 -7210 37630 -7190
rect 37592 -7224 37624 -7210
rect 37525 -7280 37624 -7224
rect 37525 -7314 37558 -7280
rect 37592 -7314 37624 -7280
rect 37525 -7370 37624 -7314
rect 37525 -7404 37558 -7370
rect 37592 -7404 37624 -7370
rect 37525 -7460 37624 -7404
rect 37525 -7494 37558 -7460
rect 37592 -7494 37624 -7460
rect 37525 -7550 37624 -7494
rect 37525 -7584 37558 -7550
rect 37592 -7584 37624 -7550
rect 37525 -7640 37624 -7584
rect 37525 -7674 37558 -7640
rect 37592 -7674 37624 -7640
rect 37525 -7730 37624 -7674
rect 37525 -7764 37558 -7730
rect 37592 -7764 37624 -7730
rect 37525 -7820 37624 -7764
rect 37525 -7854 37558 -7820
rect 37592 -7854 37624 -7820
rect 37525 -7910 37624 -7854
rect 37525 -7944 37558 -7910
rect 37592 -7944 37624 -7910
rect 37525 -8000 37624 -7944
rect 37525 -8034 37558 -8000
rect 37592 -8034 37624 -8000
rect 37525 -8090 37624 -8034
rect 36165 -8155 36435 -8124
rect 37525 -8124 37558 -8090
rect 37592 -8124 37624 -8090
rect 37525 -8155 37624 -8124
rect 33616 -8186 37624 -8155
rect 33616 -8220 33674 -8186
rect 33708 -8220 33764 -8186
rect 33798 -8220 33854 -8186
rect 33888 -8220 33944 -8186
rect 33978 -8220 34034 -8186
rect 34068 -8220 34124 -8186
rect 34158 -8220 34214 -8186
rect 34248 -8220 34304 -8186
rect 34338 -8220 34394 -8186
rect 34428 -8220 34484 -8186
rect 34518 -8220 34574 -8186
rect 34608 -8220 34664 -8186
rect 34698 -8220 34754 -8186
rect 34788 -8220 35034 -8186
rect 35068 -8220 35124 -8186
rect 35158 -8220 35214 -8186
rect 35248 -8220 35304 -8186
rect 35338 -8220 35394 -8186
rect 35428 -8220 35484 -8186
rect 35518 -8220 35574 -8186
rect 35608 -8220 35664 -8186
rect 35698 -8220 35754 -8186
rect 35788 -8220 35844 -8186
rect 35878 -8220 35934 -8186
rect 35968 -8220 36024 -8186
rect 36058 -8220 36114 -8186
rect 36148 -8220 36394 -8186
rect 36428 -8220 36484 -8186
rect 36518 -8220 36574 -8186
rect 36608 -8220 36664 -8186
rect 36698 -8220 36754 -8186
rect 36788 -8220 36844 -8186
rect 36878 -8220 36934 -8186
rect 36968 -8220 37024 -8186
rect 37058 -8220 37114 -8186
rect 37148 -8220 37204 -8186
rect 37238 -8220 37294 -8186
rect 37328 -8220 37384 -8186
rect 37418 -8220 37474 -8186
rect 37508 -8220 37624 -8186
rect 33616 -8254 37624 -8220
rect 34900 -8260 34980 -8254
rect 35560 -8340 35640 -8254
rect 36260 -8260 36340 -8254
rect 35560 -8380 35580 -8340
rect 35620 -8380 35640 -8340
rect 35560 -8440 35640 -8380
rect 35560 -8480 35580 -8440
rect 35620 -8480 35640 -8440
rect 35560 -8540 35640 -8480
rect 35560 -8580 35580 -8540
rect 35620 -8580 35640 -8540
rect 35560 -8600 35640 -8580
<< viali >>
rect 152 7120 202 7170
rect 152 7000 202 7050
rect 152 6590 202 6640
rect 152 6470 202 6520
rect 2722 6850 2772 6900
rect 2722 6730 2772 6780
rect 2390 6530 2410 6570
rect 2410 6530 2430 6570
rect 2600 6530 2620 6570
rect 2620 6530 2640 6570
rect 1210 6360 1250 6380
rect 1210 6340 1250 6360
rect 542 6060 592 6110
rect 1888 6060 1938 6110
rect 6090 7010 6130 7050
rect 6310 7010 6350 7050
rect 6420 7010 6460 7050
rect 6530 7010 6570 7050
rect 6640 7010 6680 7050
rect 6750 7010 6790 7050
rect 6200 6670 6240 6710
rect 6420 6670 6460 6710
rect 6640 6670 6680 6710
rect 7370 7010 7410 7050
rect 7590 7010 7630 7050
rect 7810 7010 7850 7050
rect 8030 7010 8070 7050
rect 8140 7010 8180 7050
rect 8250 7010 8290 7050
rect 8470 7010 8510 7050
rect 8580 7010 8620 7050
rect 8690 7010 8730 7050
rect 7480 6670 7520 6710
rect 7700 6670 7740 6710
rect 7920 6670 7960 6710
rect 8140 6670 8180 6710
rect 8360 6670 8400 6710
rect 8580 6670 8620 6710
rect 9530 7010 9570 7050
rect 9750 7010 9790 7050
rect 9860 7010 9900 7050
rect 9970 7010 10010 7050
rect 10190 7010 10230 7050
rect 9640 6670 9680 6710
rect 9860 6670 9900 6710
rect 10080 6670 10120 6710
rect 4860 6370 4910 6420
rect 4860 6250 4910 6300
rect 5670 6020 5710 6040
rect 542 5640 592 5690
rect 1888 5640 1938 5690
rect 3052 5840 3102 5890
rect 4450 5840 4500 5890
rect 5670 6000 5710 6020
rect 5670 5880 5710 5920
rect 5540 5540 5580 5580
rect 5670 5540 5710 5580
rect 5800 5540 5840 5580
rect 6520 6080 6560 6120
rect 6880 6080 6920 6120
rect 7240 6080 7280 6120
rect 7600 6080 7640 6120
rect 7960 6080 8000 6120
rect 8320 6080 8360 6120
rect 8680 6080 8720 6120
rect 9040 6080 9080 6120
rect 9400 6080 9440 6120
rect 9760 6080 9800 6120
rect 10600 6020 10640 6040
rect 6700 5340 6740 5380
rect 7060 5340 7100 5380
rect 7420 5340 7460 5380
rect 7780 5340 7820 5380
rect 7960 5340 8000 5380
rect 8140 5340 8180 5380
rect 8500 5340 8540 5380
rect 8860 5340 8900 5380
rect 9220 5340 9260 5380
rect 9400 5340 9440 5380
rect 9580 5340 9620 5380
rect 10600 6000 10640 6020
rect 10600 5880 10640 5920
rect 10470 5540 10510 5580
rect 10600 5540 10640 5580
rect 10730 5540 10770 5580
rect 6620 4840 6660 4860
rect 6620 4820 6660 4840
rect 5540 4700 5580 4740
rect 5660 4700 5700 4740
rect 5900 4700 5940 4740
rect 6140 4700 6180 4740
rect 6260 4700 6300 4740
rect 6380 4700 6420 4740
rect 6620 4700 6660 4740
rect 6860 4700 6900 4740
rect 6980 4700 7020 4740
rect 7100 4700 7140 4740
rect 7340 4700 7380 4740
rect 7580 4700 7620 4740
rect 7700 4700 7740 4740
rect 5600 4360 5640 4400
rect 5780 4360 5820 4400
rect 6020 4360 6060 4400
rect 6260 4360 6300 4400
rect 6500 4360 6540 4400
rect 6740 4360 6780 4400
rect 6980 4360 7020 4400
rect 7220 4360 7260 4400
rect 7460 4360 7500 4400
rect 7640 4360 7680 4400
rect 8700 4820 8740 4860
rect 8940 4820 8980 4860
rect 9180 4820 9220 4860
rect 9420 4820 9460 4860
rect 9660 4840 9700 4860
rect 9660 4820 9700 4840
rect 9900 4820 9940 4860
rect 10140 4820 10180 4860
rect 10380 4820 10420 4860
rect 10620 4820 10660 4860
rect 8580 4700 8620 4740
rect 8700 4700 8740 4740
rect 8940 4700 8980 4740
rect 9180 4700 9220 4740
rect 9300 4700 9340 4740
rect 9420 4700 9460 4740
rect 9660 4700 9700 4740
rect 9900 4700 9940 4740
rect 10020 4700 10060 4740
rect 10140 4700 10180 4740
rect 10380 4700 10420 4740
rect 10620 4700 10660 4740
rect 10740 4700 10780 4740
rect 8640 4360 8680 4400
rect 8820 4360 8860 4400
rect 9060 4360 9100 4400
rect 9300 4360 9340 4400
rect 9540 4360 9580 4400
rect 9780 4360 9820 4400
rect 10020 4360 10060 4400
rect 10260 4360 10300 4400
rect 10500 4360 10540 4400
rect 10680 4360 10720 4400
rect -70 3390 -30 3430
rect 6400 4040 6440 4080
rect 6280 3950 6320 3990
rect 6520 3950 6560 3990
rect 6760 3950 6800 3990
rect 7000 3950 7040 3990
rect 7240 3950 7280 3990
rect 7480 3950 7520 3990
rect 9880 4040 9920 4080
rect 8800 3950 8840 3990
rect 9040 3950 9080 3990
rect 9280 3950 9320 3990
rect 9520 3950 9560 3990
rect 9760 3950 9800 3990
rect 10000 3950 10040 3990
rect 7600 3830 7640 3870
rect 8680 3830 8720 3870
rect 6280 3710 6320 3750
rect 6400 3710 6440 3750
rect 6640 3710 6680 3750
rect 6880 3710 6920 3750
rect 7120 3710 7160 3750
rect 7360 3710 7400 3750
rect 8920 3710 8960 3750
rect 9160 3710 9200 3750
rect 9400 3710 9440 3750
rect 9640 3710 9680 3750
rect 9880 3710 9920 3750
rect 10000 3710 10040 3750
rect 36090 4010 36130 4050
rect 36310 4010 36350 4050
rect 36420 4010 36460 4050
rect 36530 4010 36570 4050
rect 36640 4010 36680 4050
rect 36750 4010 36790 4050
rect 36200 3670 36240 3710
rect 36420 3670 36460 3710
rect 36640 3670 36680 3710
rect 37370 4010 37410 4050
rect 37590 4010 37630 4050
rect 37810 4010 37850 4050
rect 38030 4010 38070 4050
rect 38140 4010 38180 4050
rect 38250 4010 38290 4050
rect 38470 4010 38510 4050
rect 38580 4010 38620 4050
rect 38690 4010 38730 4050
rect 37480 3670 37520 3710
rect 37700 3670 37740 3710
rect 37920 3670 37960 3710
rect 38140 3670 38180 3710
rect 38360 3670 38400 3710
rect 38580 3670 38620 3710
rect 39530 4010 39570 4050
rect 39750 4010 39790 4050
rect 39860 4010 39900 4050
rect 39970 4010 40010 4050
rect 40190 4010 40230 4050
rect 39640 3670 39680 3710
rect 39860 3670 39900 3710
rect 40080 3670 40120 3710
rect 5800 3360 5840 3400
rect 5980 3390 6020 3430
rect 6220 3390 6260 3430
rect 6460 3390 6500 3430
rect 6700 3390 6740 3430
rect 7180 3390 7220 3430
rect 7420 3390 7460 3430
rect 7660 3390 7700 3430
rect 7960 3360 8000 3400
rect 6880 2760 6920 2800
rect 8320 3360 8360 3400
rect 8620 3390 8660 3430
rect 8860 3390 8900 3430
rect 9100 3390 9140 3430
rect 9580 3390 9620 3430
rect 9820 3390 9860 3430
rect 10060 3390 10100 3430
rect 10300 3390 10340 3430
rect 10480 3360 10520 3400
rect 35670 3020 35710 3040
rect 9400 2760 9440 2800
rect 35670 3000 35710 3020
rect 8140 2560 8180 2600
rect 6060 2460 6100 2500
rect 6220 2460 6260 2500
rect 6380 2460 6420 2500
rect 6540 2460 6580 2500
rect 6700 2460 6740 2500
rect 6860 2460 6900 2500
rect 7020 2460 7060 2500
rect 7180 2460 7220 2500
rect 7340 2460 7380 2500
rect 7500 2460 7540 2500
rect 7660 2460 7700 2500
rect 7820 2460 7860 2500
rect 7980 2460 8020 2500
rect 8140 2460 8180 2500
rect 8300 2460 8340 2500
rect 8460 2460 8500 2500
rect 8620 2460 8660 2500
rect 8780 2460 8820 2500
rect 8940 2460 8980 2500
rect 9100 2460 9140 2500
rect 9260 2460 9300 2500
rect 9420 2460 9460 2500
rect 9580 2460 9620 2500
rect 9740 2460 9780 2500
rect 9900 2460 9940 2500
rect 10060 2460 10100 2500
rect 5980 2290 6020 2330
rect 35670 2880 35710 2920
rect 35540 2540 35580 2580
rect 35670 2540 35710 2580
rect 35800 2540 35840 2580
rect 36520 3080 36560 3120
rect 36880 3080 36920 3120
rect 37240 3080 37280 3120
rect 37600 3080 37640 3120
rect 37960 3080 38000 3120
rect 38320 3080 38360 3120
rect 38680 3080 38720 3120
rect 39040 3080 39080 3120
rect 39400 3080 39440 3120
rect 39760 3080 39800 3120
rect 10290 2290 10330 2330
rect 40600 3020 40640 3040
rect 36700 2340 36740 2380
rect 37060 2340 37100 2380
rect 37420 2340 37460 2380
rect 37780 2340 37820 2380
rect 37960 2340 38000 2380
rect 38140 2340 38180 2380
rect 38500 2340 38540 2380
rect 38860 2340 38900 2380
rect 39220 2340 39260 2380
rect 39400 2340 39440 2380
rect 39580 2340 39620 2380
rect 40600 3000 40640 3020
rect 40600 2880 40640 2920
rect 40470 2540 40510 2580
rect 40600 2540 40640 2580
rect 40730 2540 40770 2580
rect 6580 1910 6620 1950
rect 6800 1910 6840 1950
rect 6910 1910 6950 1950
rect 7020 1910 7060 1950
rect 6470 1570 6510 1610
rect 6690 1570 6730 1610
rect 6910 1570 6950 1610
rect 7130 1570 7170 1610
rect 7360 1740 7400 1780
rect 7810 1910 7850 1950
rect 8030 1910 8070 1950
rect 8140 1910 8180 1950
rect 8250 1910 8290 1950
rect 8470 1910 8510 1950
rect 7470 1740 7510 1780
rect 7750 1570 7790 1610
rect 7920 1570 7960 1610
rect 8140 1570 8180 1610
rect 8360 1570 8400 1610
rect 8580 1570 8620 1610
rect 8810 1740 8850 1780
rect 9260 1910 9300 1950
rect 9370 1910 9410 1950
rect 9480 1910 9520 1950
rect 9700 1910 9740 1950
rect 8920 1740 8960 1780
rect 9150 1570 9190 1610
rect 9370 1570 9410 1610
rect 9590 1570 9630 1610
rect 9810 1570 9850 1610
rect 36620 1840 36660 1860
rect 10040 1740 10080 1780
rect 36620 1820 36660 1840
rect 35540 1700 35580 1740
rect 35660 1700 35700 1740
rect 35900 1700 35940 1740
rect 36140 1700 36180 1740
rect 36260 1700 36300 1740
rect 36380 1700 36420 1740
rect 36620 1700 36660 1740
rect 36860 1700 36900 1740
rect 36980 1700 37020 1740
rect 37100 1700 37140 1740
rect 37340 1700 37380 1740
rect 37580 1700 37620 1740
rect 37700 1700 37740 1740
rect 35600 1360 35640 1400
rect 35780 1360 35820 1400
rect 36020 1360 36060 1400
rect 36260 1360 36300 1400
rect 36500 1360 36540 1400
rect 36740 1360 36780 1400
rect 36980 1360 37020 1400
rect 37220 1360 37260 1400
rect 37460 1360 37500 1400
rect 37640 1360 37680 1400
rect 38700 1820 38740 1860
rect 38940 1820 38980 1860
rect 39180 1820 39220 1860
rect 39420 1820 39460 1860
rect 39660 1840 39700 1860
rect 39660 1820 39700 1840
rect 39900 1820 39940 1860
rect 40140 1820 40180 1860
rect 40380 1820 40420 1860
rect 40620 1820 40660 1860
rect 38580 1700 38620 1740
rect 38700 1700 38740 1740
rect 38940 1700 38980 1740
rect 39180 1700 39220 1740
rect 39300 1700 39340 1740
rect 39420 1700 39460 1740
rect 39660 1700 39700 1740
rect 39900 1700 39940 1740
rect 40020 1700 40060 1740
rect 40140 1700 40180 1740
rect 40380 1700 40420 1740
rect 40620 1700 40660 1740
rect 40740 1700 40780 1740
rect 38640 1360 38680 1400
rect 38820 1360 38860 1400
rect 39060 1360 39100 1400
rect 39300 1360 39340 1400
rect 39540 1360 39580 1400
rect 39780 1360 39820 1400
rect 40020 1360 40060 1400
rect 40260 1360 40300 1400
rect 40500 1360 40540 1400
rect 40680 1360 40720 1400
rect 36400 1040 36440 1080
rect 36280 950 36320 990
rect 36520 950 36560 990
rect 36760 950 36800 990
rect 37000 950 37040 990
rect 37240 950 37280 990
rect 37480 950 37520 990
rect 39880 1040 39920 1080
rect 38800 950 38840 990
rect 39040 950 39080 990
rect 39280 950 39320 990
rect 39520 950 39560 990
rect 39760 950 39800 990
rect 40000 950 40040 990
rect 37600 830 37640 870
rect 38680 830 38720 870
rect 36280 710 36320 750
rect 36400 710 36440 750
rect 36640 710 36680 750
rect 36880 710 36920 750
rect 37120 710 37160 750
rect 37360 710 37400 750
rect 38920 710 38960 750
rect 39160 710 39200 750
rect 39400 710 39440 750
rect 39640 710 39680 750
rect 39880 710 39920 750
rect 40000 710 40040 750
rect 35800 360 35840 400
rect 35980 390 36020 430
rect 36220 390 36260 430
rect 36460 390 36500 430
rect 36700 390 36740 430
rect 37180 390 37220 430
rect 37420 390 37460 430
rect 37660 390 37700 430
rect 37960 360 38000 400
rect 36880 -240 36920 -200
rect 38320 360 38360 400
rect 38620 390 38660 430
rect 38860 390 38900 430
rect 39100 390 39140 430
rect 39580 390 39620 430
rect 39820 390 39860 430
rect 40060 390 40100 430
rect 40300 390 40340 430
rect 40480 360 40520 400
rect 39400 -240 39440 -200
rect 38140 -440 38180 -400
rect 36060 -540 36100 -500
rect 36220 -540 36260 -500
rect 36380 -540 36420 -500
rect 36540 -540 36580 -500
rect 36700 -540 36740 -500
rect 36860 -540 36900 -500
rect 37020 -540 37060 -500
rect 37180 -540 37220 -500
rect 37340 -540 37380 -500
rect 37500 -540 37540 -500
rect 37660 -540 37700 -500
rect 37820 -540 37860 -500
rect 37980 -540 38020 -500
rect 38140 -540 38180 -500
rect 38300 -540 38340 -500
rect 38460 -540 38500 -500
rect 38620 -540 38660 -500
rect 38780 -540 38820 -500
rect 38940 -540 38980 -500
rect 39100 -540 39140 -500
rect 39260 -540 39300 -500
rect 39420 -540 39460 -500
rect 39580 -540 39620 -500
rect 39740 -540 39780 -500
rect 39900 -540 39940 -500
rect 40060 -540 40100 -500
rect 35980 -710 36020 -670
rect 40290 -710 40330 -670
rect 36580 -1090 36620 -1050
rect 36800 -1090 36840 -1050
rect 36910 -1090 36950 -1050
rect 37020 -1090 37060 -1050
rect 36470 -1430 36510 -1390
rect 36690 -1430 36730 -1390
rect 36910 -1430 36950 -1390
rect 37130 -1430 37170 -1390
rect 37360 -1260 37400 -1220
rect 37810 -1090 37850 -1050
rect 38030 -1090 38070 -1050
rect 38140 -1090 38180 -1050
rect 38250 -1090 38290 -1050
rect 38470 -1090 38510 -1050
rect 37470 -1260 37510 -1220
rect 37750 -1430 37790 -1390
rect 37920 -1430 37960 -1390
rect 38140 -1430 38180 -1390
rect 38360 -1430 38400 -1390
rect 38580 -1430 38620 -1390
rect 38810 -1260 38850 -1220
rect 39260 -1090 39300 -1050
rect 39370 -1090 39410 -1050
rect 39480 -1090 39520 -1050
rect 39700 -1090 39740 -1050
rect 38920 -1260 38960 -1220
rect 39150 -1430 39190 -1390
rect 39370 -1430 39410 -1390
rect 39590 -1430 39630 -1390
rect 39810 -1430 39850 -1390
rect 40040 -1260 40080 -1220
rect 44152 -2880 44202 -2830
rect 44152 -3000 44202 -2950
rect 44152 -3410 44202 -3360
rect 44152 -3530 44202 -3480
rect 46722 -3150 46772 -3100
rect 46722 -3270 46772 -3220
rect 46390 -3470 46410 -3430
rect 46410 -3470 46430 -3430
rect 46600 -3470 46620 -3430
rect 46620 -3470 46640 -3430
rect 45210 -3640 45250 -3620
rect 45210 -3660 45250 -3640
rect 44542 -3940 44592 -3890
rect 45888 -3940 45938 -3890
rect 48860 -3630 48910 -3580
rect 48860 -3750 48910 -3700
rect 34000 -4636 34006 -4630
rect 34006 -4636 34034 -4630
rect 34000 -4664 34034 -4636
rect 34100 -4664 34134 -4630
rect 34200 -4664 34234 -4630
rect 34300 -4636 34332 -4630
rect 34332 -4636 34334 -4630
rect 34400 -4636 34422 -4630
rect 34422 -4636 34434 -4630
rect 34500 -4636 34512 -4630
rect 34512 -4636 34534 -4630
rect 34300 -4664 34334 -4636
rect 34400 -4664 34434 -4636
rect 34500 -4664 34534 -4636
rect 34000 -4764 34034 -4730
rect 34100 -4764 34134 -4730
rect 34200 -4764 34234 -4730
rect 34300 -4764 34334 -4730
rect 34400 -4764 34434 -4730
rect 34500 -4764 34534 -4730
rect 34000 -4864 34034 -4830
rect 34100 -4864 34134 -4830
rect 34200 -4864 34234 -4830
rect 34300 -4864 34334 -4830
rect 34400 -4864 34434 -4830
rect 34500 -4864 34534 -4830
rect 34000 -4962 34034 -4930
rect 34000 -4964 34006 -4962
rect 34006 -4964 34034 -4962
rect 34100 -4964 34134 -4930
rect 34200 -4964 34234 -4930
rect 34300 -4962 34334 -4930
rect 34400 -4962 34434 -4930
rect 34500 -4962 34534 -4930
rect 34300 -4964 34332 -4962
rect 34332 -4964 34334 -4962
rect 34400 -4964 34422 -4962
rect 34422 -4964 34434 -4962
rect 34500 -4964 34512 -4962
rect 34512 -4964 34534 -4962
rect 34000 -5052 34034 -5030
rect 34000 -5064 34006 -5052
rect 34006 -5064 34034 -5052
rect 34100 -5064 34134 -5030
rect 34200 -5064 34234 -5030
rect 34300 -5052 34334 -5030
rect 34400 -5052 34434 -5030
rect 34500 -5052 34534 -5030
rect 34300 -5064 34332 -5052
rect 34332 -5064 34334 -5052
rect 34400 -5064 34422 -5052
rect 34422 -5064 34434 -5052
rect 34500 -5064 34512 -5052
rect 34512 -5064 34534 -5052
rect 34000 -5142 34034 -5130
rect 34000 -5164 34006 -5142
rect 34006 -5164 34034 -5142
rect 34100 -5164 34134 -5130
rect 34200 -5164 34234 -5130
rect 34300 -5142 34334 -5130
rect 34400 -5142 34434 -5130
rect 34500 -5142 34534 -5130
rect 34300 -5164 34332 -5142
rect 34332 -5164 34334 -5142
rect 34400 -5164 34422 -5142
rect 34422 -5164 34434 -5142
rect 34500 -5164 34512 -5142
rect 34512 -5164 34534 -5142
rect 35360 -4636 35366 -4630
rect 35366 -4636 35394 -4630
rect 35360 -4664 35394 -4636
rect 35460 -4664 35494 -4630
rect 35560 -4664 35594 -4630
rect 35660 -4636 35692 -4630
rect 35692 -4636 35694 -4630
rect 35760 -4636 35782 -4630
rect 35782 -4636 35794 -4630
rect 35860 -4636 35872 -4630
rect 35872 -4636 35894 -4630
rect 35660 -4664 35694 -4636
rect 35760 -4664 35794 -4636
rect 35860 -4664 35894 -4636
rect 35360 -4764 35394 -4730
rect 35460 -4764 35494 -4730
rect 35560 -4764 35594 -4730
rect 35660 -4764 35694 -4730
rect 35760 -4764 35794 -4730
rect 35860 -4764 35894 -4730
rect 35360 -4864 35394 -4830
rect 35460 -4864 35494 -4830
rect 35560 -4864 35594 -4830
rect 35660 -4864 35694 -4830
rect 35760 -4864 35794 -4830
rect 35860 -4864 35894 -4830
rect 35360 -4962 35394 -4930
rect 35360 -4964 35366 -4962
rect 35366 -4964 35394 -4962
rect 35460 -4964 35494 -4930
rect 35560 -4964 35594 -4930
rect 35660 -4962 35694 -4930
rect 35760 -4962 35794 -4930
rect 35860 -4962 35894 -4930
rect 35660 -4964 35692 -4962
rect 35692 -4964 35694 -4962
rect 35760 -4964 35782 -4962
rect 35782 -4964 35794 -4962
rect 35860 -4964 35872 -4962
rect 35872 -4964 35894 -4962
rect 35360 -5052 35394 -5030
rect 35360 -5064 35366 -5052
rect 35366 -5064 35394 -5052
rect 35460 -5064 35494 -5030
rect 35560 -5064 35594 -5030
rect 35660 -5052 35694 -5030
rect 35760 -5052 35794 -5030
rect 35860 -5052 35894 -5030
rect 35660 -5064 35692 -5052
rect 35692 -5064 35694 -5052
rect 35760 -5064 35782 -5052
rect 35782 -5064 35794 -5052
rect 35860 -5064 35872 -5052
rect 35872 -5064 35894 -5052
rect 35360 -5142 35394 -5130
rect 35360 -5164 35366 -5142
rect 35366 -5164 35394 -5142
rect 35460 -5164 35494 -5130
rect 35560 -5164 35594 -5130
rect 35660 -5142 35694 -5130
rect 35760 -5142 35794 -5130
rect 35860 -5142 35894 -5130
rect 35660 -5164 35692 -5142
rect 35692 -5164 35694 -5142
rect 35760 -5164 35782 -5142
rect 35782 -5164 35794 -5142
rect 35860 -5164 35872 -5142
rect 35872 -5164 35894 -5142
rect 36720 -4636 36726 -4630
rect 36726 -4636 36754 -4630
rect 36720 -4664 36754 -4636
rect 36820 -4664 36854 -4630
rect 36920 -4664 36954 -4630
rect 37020 -4636 37052 -4630
rect 37052 -4636 37054 -4630
rect 37120 -4636 37142 -4630
rect 37142 -4636 37154 -4630
rect 37220 -4636 37232 -4630
rect 37232 -4636 37254 -4630
rect 37020 -4664 37054 -4636
rect 37120 -4664 37154 -4636
rect 37220 -4664 37254 -4636
rect 36720 -4764 36754 -4730
rect 36820 -4764 36854 -4730
rect 36920 -4764 36954 -4730
rect 37020 -4764 37054 -4730
rect 37120 -4764 37154 -4730
rect 37220 -4764 37254 -4730
rect 36720 -4864 36754 -4830
rect 36820 -4864 36854 -4830
rect 36920 -4864 36954 -4830
rect 37020 -4864 37054 -4830
rect 37120 -4864 37154 -4830
rect 37220 -4864 37254 -4830
rect 36720 -4962 36754 -4930
rect 36720 -4964 36726 -4962
rect 36726 -4964 36754 -4962
rect 36820 -4964 36854 -4930
rect 36920 -4964 36954 -4930
rect 37020 -4962 37054 -4930
rect 37120 -4962 37154 -4930
rect 37220 -4962 37254 -4930
rect 37020 -4964 37052 -4962
rect 37052 -4964 37054 -4962
rect 37120 -4964 37142 -4962
rect 37142 -4964 37154 -4962
rect 37220 -4964 37232 -4962
rect 37232 -4964 37254 -4962
rect 36720 -5052 36754 -5030
rect 36720 -5064 36726 -5052
rect 36726 -5064 36754 -5052
rect 36820 -5064 36854 -5030
rect 36920 -5064 36954 -5030
rect 37020 -5052 37054 -5030
rect 37120 -5052 37154 -5030
rect 37220 -5052 37254 -5030
rect 37020 -5064 37052 -5052
rect 37052 -5064 37054 -5052
rect 37120 -5064 37142 -5052
rect 37142 -5064 37154 -5052
rect 37220 -5064 37232 -5052
rect 37232 -5064 37254 -5052
rect 36720 -5142 36754 -5130
rect 36720 -5164 36726 -5142
rect 36726 -5164 36754 -5142
rect 36820 -5164 36854 -5130
rect 36920 -5164 36954 -5130
rect 37020 -5142 37054 -5130
rect 37120 -5142 37154 -5130
rect 37220 -5142 37254 -5130
rect 37020 -5164 37052 -5142
rect 37052 -5164 37054 -5142
rect 37120 -5164 37142 -5142
rect 37142 -5164 37154 -5142
rect 37220 -5164 37232 -5142
rect 37232 -5164 37254 -5142
rect 44542 -4360 44592 -4310
rect 45888 -4360 45938 -4310
rect 47052 -4160 47102 -4110
rect 48450 -4160 48500 -4110
rect 34000 -5996 34006 -5990
rect 34006 -5996 34034 -5990
rect 34000 -6024 34034 -5996
rect 34100 -6024 34134 -5990
rect 34200 -6024 34234 -5990
rect 34300 -5996 34332 -5990
rect 34332 -5996 34334 -5990
rect 34400 -5996 34422 -5990
rect 34422 -5996 34434 -5990
rect 34500 -5996 34512 -5990
rect 34512 -5996 34534 -5990
rect 34300 -6024 34334 -5996
rect 34400 -6024 34434 -5996
rect 34500 -6024 34534 -5996
rect 34000 -6124 34034 -6090
rect 34100 -6124 34134 -6090
rect 34200 -6124 34234 -6090
rect 34300 -6124 34334 -6090
rect 34400 -6124 34434 -6090
rect 34500 -6124 34534 -6090
rect 34000 -6224 34034 -6190
rect 34100 -6224 34134 -6190
rect 34200 -6224 34234 -6190
rect 34300 -6224 34334 -6190
rect 34400 -6224 34434 -6190
rect 34500 -6224 34534 -6190
rect 34000 -6322 34034 -6290
rect 34000 -6324 34006 -6322
rect 34006 -6324 34034 -6322
rect 34100 -6324 34134 -6290
rect 34200 -6324 34234 -6290
rect 34300 -6322 34334 -6290
rect 34400 -6322 34434 -6290
rect 34500 -6322 34534 -6290
rect 34300 -6324 34332 -6322
rect 34332 -6324 34334 -6322
rect 34400 -6324 34422 -6322
rect 34422 -6324 34434 -6322
rect 34500 -6324 34512 -6322
rect 34512 -6324 34534 -6322
rect 34000 -6412 34034 -6390
rect 34000 -6424 34006 -6412
rect 34006 -6424 34034 -6412
rect 34100 -6424 34134 -6390
rect 34200 -6424 34234 -6390
rect 34300 -6412 34334 -6390
rect 34400 -6412 34434 -6390
rect 34500 -6412 34534 -6390
rect 34300 -6424 34332 -6412
rect 34332 -6424 34334 -6412
rect 34400 -6424 34422 -6412
rect 34422 -6424 34434 -6412
rect 34500 -6424 34512 -6412
rect 34512 -6424 34534 -6412
rect 34000 -6502 34034 -6490
rect 34000 -6524 34006 -6502
rect 34006 -6524 34034 -6502
rect 34100 -6524 34134 -6490
rect 34200 -6524 34234 -6490
rect 34300 -6502 34334 -6490
rect 34400 -6502 34434 -6490
rect 34500 -6502 34534 -6490
rect 34300 -6524 34332 -6502
rect 34332 -6524 34334 -6502
rect 34400 -6524 34422 -6502
rect 34422 -6524 34434 -6502
rect 34500 -6524 34512 -6502
rect 34512 -6524 34534 -6502
rect 35360 -5996 35366 -5990
rect 35366 -5996 35394 -5990
rect 35360 -6024 35394 -5996
rect 35460 -6024 35494 -5990
rect 35560 -6024 35594 -5990
rect 35660 -5996 35692 -5990
rect 35692 -5996 35694 -5990
rect 35760 -5996 35782 -5990
rect 35782 -5996 35794 -5990
rect 35860 -5996 35872 -5990
rect 35872 -5996 35894 -5990
rect 35660 -6024 35694 -5996
rect 35760 -6024 35794 -5996
rect 35860 -6024 35894 -5996
rect 35360 -6124 35394 -6090
rect 35460 -6124 35494 -6090
rect 35560 -6124 35594 -6090
rect 35660 -6124 35694 -6090
rect 35760 -6124 35794 -6090
rect 35860 -6124 35894 -6090
rect 35360 -6224 35394 -6190
rect 35460 -6224 35494 -6190
rect 35560 -6224 35594 -6190
rect 35660 -6224 35694 -6190
rect 35760 -6224 35794 -6190
rect 35860 -6224 35894 -6190
rect 35360 -6322 35394 -6290
rect 35360 -6324 35366 -6322
rect 35366 -6324 35394 -6322
rect 35460 -6324 35494 -6290
rect 35560 -6324 35594 -6290
rect 35660 -6322 35694 -6290
rect 35760 -6322 35794 -6290
rect 35860 -6322 35894 -6290
rect 35660 -6324 35692 -6322
rect 35692 -6324 35694 -6322
rect 35760 -6324 35782 -6322
rect 35782 -6324 35794 -6322
rect 35860 -6324 35872 -6322
rect 35872 -6324 35894 -6322
rect 35360 -6412 35394 -6390
rect 35360 -6424 35366 -6412
rect 35366 -6424 35394 -6412
rect 35460 -6424 35494 -6390
rect 35560 -6424 35594 -6390
rect 35660 -6412 35694 -6390
rect 35760 -6412 35794 -6390
rect 35860 -6412 35894 -6390
rect 35660 -6424 35692 -6412
rect 35692 -6424 35694 -6412
rect 35760 -6424 35782 -6412
rect 35782 -6424 35794 -6412
rect 35860 -6424 35872 -6412
rect 35872 -6424 35894 -6412
rect 35360 -6502 35394 -6490
rect 35360 -6524 35366 -6502
rect 35366 -6524 35394 -6502
rect 35460 -6524 35494 -6490
rect 35560 -6524 35594 -6490
rect 35660 -6502 35694 -6490
rect 35760 -6502 35794 -6490
rect 35860 -6502 35894 -6490
rect 35660 -6524 35692 -6502
rect 35692 -6524 35694 -6502
rect 35760 -6524 35782 -6502
rect 35782 -6524 35794 -6502
rect 35860 -6524 35872 -6502
rect 35872 -6524 35894 -6502
rect 36720 -5996 36726 -5990
rect 36726 -5996 36754 -5990
rect 36720 -6024 36754 -5996
rect 36820 -6024 36854 -5990
rect 36920 -6024 36954 -5990
rect 37020 -5996 37052 -5990
rect 37052 -5996 37054 -5990
rect 37120 -5996 37142 -5990
rect 37142 -5996 37154 -5990
rect 37220 -5996 37232 -5990
rect 37232 -5996 37254 -5990
rect 37020 -6024 37054 -5996
rect 37120 -6024 37154 -5996
rect 37220 -6024 37254 -5996
rect 36720 -6124 36754 -6090
rect 36820 -6124 36854 -6090
rect 36920 -6124 36954 -6090
rect 37020 -6124 37054 -6090
rect 37120 -6124 37154 -6090
rect 37220 -6124 37254 -6090
rect 36720 -6224 36754 -6190
rect 36820 -6224 36854 -6190
rect 36920 -6224 36954 -6190
rect 37020 -6224 37054 -6190
rect 37120 -6224 37154 -6190
rect 37220 -6224 37254 -6190
rect 36720 -6322 36754 -6290
rect 36720 -6324 36726 -6322
rect 36726 -6324 36754 -6322
rect 36820 -6324 36854 -6290
rect 36920 -6324 36954 -6290
rect 37020 -6322 37054 -6290
rect 37120 -6322 37154 -6290
rect 37220 -6322 37254 -6290
rect 37020 -6324 37052 -6322
rect 37052 -6324 37054 -6322
rect 37120 -6324 37142 -6322
rect 37142 -6324 37154 -6322
rect 37220 -6324 37232 -6322
rect 37232 -6324 37254 -6322
rect 36720 -6412 36754 -6390
rect 36720 -6424 36726 -6412
rect 36726 -6424 36754 -6412
rect 36820 -6424 36854 -6390
rect 36920 -6424 36954 -6390
rect 37020 -6412 37054 -6390
rect 37120 -6412 37154 -6390
rect 37220 -6412 37254 -6390
rect 37020 -6424 37052 -6412
rect 37052 -6424 37054 -6412
rect 37120 -6424 37142 -6412
rect 37142 -6424 37154 -6412
rect 37220 -6424 37232 -6412
rect 37232 -6424 37254 -6412
rect 36720 -6502 36754 -6490
rect 36720 -6524 36726 -6502
rect 36726 -6524 36754 -6502
rect 36820 -6524 36854 -6490
rect 36920 -6524 36954 -6490
rect 37020 -6502 37054 -6490
rect 37120 -6502 37154 -6490
rect 37220 -6502 37254 -6490
rect 37020 -6524 37052 -6502
rect 37052 -6524 37054 -6502
rect 37120 -6524 37142 -6502
rect 37142 -6524 37154 -6502
rect 37220 -6524 37232 -6502
rect 37232 -6524 37254 -6502
rect 34000 -7356 34006 -7350
rect 34006 -7356 34034 -7350
rect 34000 -7384 34034 -7356
rect 34100 -7384 34134 -7350
rect 34200 -7384 34234 -7350
rect 34300 -7356 34332 -7350
rect 34332 -7356 34334 -7350
rect 34400 -7356 34422 -7350
rect 34422 -7356 34434 -7350
rect 34500 -7356 34512 -7350
rect 34512 -7356 34534 -7350
rect 34300 -7384 34334 -7356
rect 34400 -7384 34434 -7356
rect 34500 -7384 34534 -7356
rect 34000 -7484 34034 -7450
rect 34100 -7484 34134 -7450
rect 34200 -7484 34234 -7450
rect 34300 -7484 34334 -7450
rect 34400 -7484 34434 -7450
rect 34500 -7484 34534 -7450
rect 34000 -7584 34034 -7550
rect 34100 -7584 34134 -7550
rect 34200 -7584 34234 -7550
rect 34300 -7584 34334 -7550
rect 34400 -7584 34434 -7550
rect 34500 -7584 34534 -7550
rect 34000 -7682 34034 -7650
rect 34000 -7684 34006 -7682
rect 34006 -7684 34034 -7682
rect 34100 -7684 34134 -7650
rect 34200 -7684 34234 -7650
rect 34300 -7682 34334 -7650
rect 34400 -7682 34434 -7650
rect 34500 -7682 34534 -7650
rect 34300 -7684 34332 -7682
rect 34332 -7684 34334 -7682
rect 34400 -7684 34422 -7682
rect 34422 -7684 34434 -7682
rect 34500 -7684 34512 -7682
rect 34512 -7684 34534 -7682
rect 34000 -7772 34034 -7750
rect 34000 -7784 34006 -7772
rect 34006 -7784 34034 -7772
rect 34100 -7784 34134 -7750
rect 34200 -7784 34234 -7750
rect 34300 -7772 34334 -7750
rect 34400 -7772 34434 -7750
rect 34500 -7772 34534 -7750
rect 34300 -7784 34332 -7772
rect 34332 -7784 34334 -7772
rect 34400 -7784 34422 -7772
rect 34422 -7784 34434 -7772
rect 34500 -7784 34512 -7772
rect 34512 -7784 34534 -7772
rect 34000 -7862 34034 -7850
rect 34000 -7884 34006 -7862
rect 34006 -7884 34034 -7862
rect 34100 -7884 34134 -7850
rect 34200 -7884 34234 -7850
rect 34300 -7862 34334 -7850
rect 34400 -7862 34434 -7850
rect 34500 -7862 34534 -7850
rect 34300 -7884 34332 -7862
rect 34332 -7884 34334 -7862
rect 34400 -7884 34422 -7862
rect 34422 -7884 34434 -7862
rect 34500 -7884 34512 -7862
rect 34512 -7884 34534 -7862
rect 35360 -7356 35366 -7350
rect 35366 -7356 35394 -7350
rect 35360 -7384 35394 -7356
rect 35460 -7384 35494 -7350
rect 35560 -7384 35594 -7350
rect 35660 -7356 35692 -7350
rect 35692 -7356 35694 -7350
rect 35760 -7356 35782 -7350
rect 35782 -7356 35794 -7350
rect 35860 -7356 35872 -7350
rect 35872 -7356 35894 -7350
rect 35660 -7384 35694 -7356
rect 35760 -7384 35794 -7356
rect 35860 -7384 35894 -7356
rect 35360 -7484 35394 -7450
rect 35460 -7484 35494 -7450
rect 35560 -7484 35594 -7450
rect 35660 -7484 35694 -7450
rect 35760 -7484 35794 -7450
rect 35860 -7484 35894 -7450
rect 35360 -7584 35394 -7550
rect 35460 -7584 35494 -7550
rect 35560 -7584 35594 -7550
rect 35660 -7584 35694 -7550
rect 35760 -7584 35794 -7550
rect 35860 -7584 35894 -7550
rect 35360 -7682 35394 -7650
rect 35360 -7684 35366 -7682
rect 35366 -7684 35394 -7682
rect 35460 -7684 35494 -7650
rect 35560 -7684 35594 -7650
rect 35660 -7682 35694 -7650
rect 35760 -7682 35794 -7650
rect 35860 -7682 35894 -7650
rect 35660 -7684 35692 -7682
rect 35692 -7684 35694 -7682
rect 35760 -7684 35782 -7682
rect 35782 -7684 35794 -7682
rect 35860 -7684 35872 -7682
rect 35872 -7684 35894 -7682
rect 35360 -7772 35394 -7750
rect 35360 -7784 35366 -7772
rect 35366 -7784 35394 -7772
rect 35460 -7784 35494 -7750
rect 35560 -7784 35594 -7750
rect 35660 -7772 35694 -7750
rect 35760 -7772 35794 -7750
rect 35860 -7772 35894 -7750
rect 35660 -7784 35692 -7772
rect 35692 -7784 35694 -7772
rect 35760 -7784 35782 -7772
rect 35782 -7784 35794 -7772
rect 35860 -7784 35872 -7772
rect 35872 -7784 35894 -7772
rect 35360 -7862 35394 -7850
rect 35360 -7884 35366 -7862
rect 35366 -7884 35394 -7862
rect 35460 -7884 35494 -7850
rect 35560 -7884 35594 -7850
rect 35660 -7862 35694 -7850
rect 35760 -7862 35794 -7850
rect 35860 -7862 35894 -7850
rect 35660 -7884 35692 -7862
rect 35692 -7884 35694 -7862
rect 35760 -7884 35782 -7862
rect 35782 -7884 35794 -7862
rect 35860 -7884 35872 -7862
rect 35872 -7884 35894 -7862
rect 36720 -7356 36726 -7350
rect 36726 -7356 36754 -7350
rect 36720 -7384 36754 -7356
rect 36820 -7384 36854 -7350
rect 36920 -7384 36954 -7350
rect 37020 -7356 37052 -7350
rect 37052 -7356 37054 -7350
rect 37120 -7356 37142 -7350
rect 37142 -7356 37154 -7350
rect 37220 -7356 37232 -7350
rect 37232 -7356 37254 -7350
rect 37020 -7384 37054 -7356
rect 37120 -7384 37154 -7356
rect 37220 -7384 37254 -7356
rect 36720 -7484 36754 -7450
rect 36820 -7484 36854 -7450
rect 36920 -7484 36954 -7450
rect 37020 -7484 37054 -7450
rect 37120 -7484 37154 -7450
rect 37220 -7484 37254 -7450
rect 36720 -7584 36754 -7550
rect 36820 -7584 36854 -7550
rect 36920 -7584 36954 -7550
rect 37020 -7584 37054 -7550
rect 37120 -7584 37154 -7550
rect 37220 -7584 37254 -7550
rect 36720 -7682 36754 -7650
rect 36720 -7684 36726 -7682
rect 36726 -7684 36754 -7682
rect 36820 -7684 36854 -7650
rect 36920 -7684 36954 -7650
rect 37020 -7682 37054 -7650
rect 37120 -7682 37154 -7650
rect 37220 -7682 37254 -7650
rect 37020 -7684 37052 -7682
rect 37052 -7684 37054 -7682
rect 37120 -7684 37142 -7682
rect 37142 -7684 37154 -7682
rect 37220 -7684 37232 -7682
rect 37232 -7684 37254 -7682
rect 36720 -7772 36754 -7750
rect 36720 -7784 36726 -7772
rect 36726 -7784 36754 -7772
rect 36820 -7784 36854 -7750
rect 36920 -7784 36954 -7750
rect 37020 -7772 37054 -7750
rect 37120 -7772 37154 -7750
rect 37220 -7772 37254 -7750
rect 37020 -7784 37052 -7772
rect 37052 -7784 37054 -7772
rect 37120 -7784 37142 -7772
rect 37142 -7784 37154 -7772
rect 37220 -7784 37232 -7772
rect 37232 -7784 37254 -7772
rect 36720 -7862 36754 -7850
rect 36720 -7884 36726 -7862
rect 36726 -7884 36754 -7862
rect 36820 -7884 36854 -7850
rect 36920 -7884 36954 -7850
rect 37020 -7862 37054 -7850
rect 37120 -7862 37154 -7850
rect 37220 -7862 37254 -7850
rect 37020 -7884 37052 -7862
rect 37052 -7884 37054 -7862
rect 37120 -7884 37142 -7862
rect 37142 -7884 37154 -7862
rect 37220 -7884 37232 -7862
rect 37232 -7884 37254 -7862
rect 35580 -8580 35620 -8540
<< metal1 >>
rect 2700 7750 2780 7760
rect 2700 7690 2710 7750
rect 2770 7690 2780 7750
rect 32700 7750 32780 7760
rect 2700 7680 2780 7690
rect 8880 7690 8960 7700
rect -30 7590 50 7600
rect -30 7530 -20 7590
rect 40 7530 50 7590
rect -30 7520 50 7530
rect 1880 7590 1960 7600
rect 1880 7530 1890 7590
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect -120 7480 -40 7490
rect -120 7420 -110 7480
rect -50 7420 -40 7480
rect -120 7410 -40 7420
rect -100 6120 -60 7410
rect -120 6110 -40 6120
rect -120 6050 -110 6110
rect -50 6050 -40 6110
rect -120 6040 -40 6050
rect -10 5710 30 7520
rect 2510 7380 2590 7390
rect 2510 7320 2520 7380
rect 2580 7320 2590 7380
rect 2510 7310 2590 7320
rect 140 7280 220 7290
rect 140 7220 150 7280
rect 210 7220 220 7280
rect 140 7210 220 7220
rect 150 7180 200 7210
rect 132 7110 142 7180
rect 212 7110 222 7180
rect 132 6990 142 7060
rect 212 6990 222 7060
rect 2530 6760 2570 7310
rect 2720 6910 2760 7680
rect 8880 7630 8890 7690
rect 8950 7630 8960 7690
rect 32700 7690 32710 7750
rect 32770 7690 32780 7750
rect 32700 7680 32780 7690
rect 38880 7690 38960 7700
rect 8880 7620 8960 7630
rect 3270 7590 3370 7610
rect 3270 7530 3290 7590
rect 3350 7530 3370 7590
rect 5020 7600 5100 7610
rect 5020 7540 5030 7600
rect 5090 7540 5100 7600
rect 5020 7530 5100 7540
rect 9310 7590 9390 7600
rect 9310 7530 9320 7590
rect 9380 7530 9390 7590
rect 3270 7510 3370 7530
rect 2702 6840 2712 6910
rect 2782 6840 2792 6910
rect 2722 6790 2762 6840
rect 140 6750 220 6760
rect 140 6690 150 6750
rect 210 6690 220 6750
rect 140 6680 220 6690
rect 2510 6750 2590 6760
rect 2510 6690 2520 6750
rect 2580 6690 2590 6750
rect 2702 6720 2712 6790
rect 2782 6720 2792 6790
rect 2510 6680 2590 6690
rect 150 6650 200 6680
rect 132 6580 142 6650
rect 212 6580 222 6650
rect 2370 6580 2450 6590
rect 132 6460 142 6530
rect 212 6460 222 6530
rect 2370 6520 2380 6580
rect 2440 6520 2450 6580
rect 2370 6510 2450 6520
rect 2580 6580 2660 6590
rect 2580 6520 2590 6580
rect 2650 6520 2660 6580
rect 2580 6510 2660 6520
rect 1190 6390 1270 6400
rect 1190 6330 1200 6390
rect 1260 6330 1270 6390
rect 4840 6360 4850 6430
rect 4920 6360 4930 6430
rect 1190 6320 1270 6330
rect 4840 6310 4930 6320
rect 4840 6240 4850 6310
rect 4920 6240 4930 6310
rect 4840 6230 4930 6240
rect 522 6050 532 6120
rect 602 6050 612 6120
rect 1868 6050 1878 6120
rect 1948 6050 1958 6120
rect 2420 6110 2500 6120
rect 2420 6050 2430 6110
rect 2490 6050 2500 6110
rect 2420 6040 2500 6050
rect 2210 5900 2290 5910
rect 2210 5840 2220 5900
rect 2280 5840 2290 5900
rect 2210 5830 2290 5840
rect -30 5700 50 5710
rect -30 5640 -20 5700
rect 40 5640 50 5700
rect -30 5630 50 5640
rect 522 5630 532 5700
rect 602 5630 612 5700
rect 1868 5630 1878 5700
rect 1948 5630 1958 5700
rect 2230 5100 2270 5830
rect 2440 5610 2480 6040
rect 4860 5900 4900 6230
rect 3032 5830 3042 5900
rect 3112 5830 3122 5900
rect 4430 5830 4440 5900
rect 4510 5830 4520 5900
rect 4840 5890 4920 5900
rect 4840 5830 4850 5890
rect 4910 5830 4920 5890
rect 4840 5820 4920 5830
rect 2420 5600 2500 5610
rect 2420 5540 2430 5600
rect 2490 5540 2500 5600
rect 2420 5530 2500 5540
rect 4750 5600 4830 5610
rect 4750 5540 4760 5600
rect 4820 5540 4830 5600
rect 4750 5530 4830 5540
rect 4660 5280 4740 5290
rect 4660 5220 4670 5280
rect 4730 5220 4740 5280
rect 4660 5210 4740 5220
rect 4550 5190 4630 5200
rect 4550 5130 4560 5190
rect 4620 5130 4630 5190
rect 4550 5120 4630 5130
rect 550 4400 3970 5100
rect -220 3440 -140 3450
rect -220 3380 -210 3440
rect -150 3430 -140 3440
rect -90 3440 -10 3450
rect -90 3430 -80 3440
rect -150 3390 -80 3430
rect -150 3380 -140 3390
rect -220 3370 -140 3380
rect -90 3380 -80 3390
rect -20 3380 -10 3440
rect -90 3370 -10 3380
rect 550 2380 1250 4400
rect 1904 3420 2604 3740
rect 1904 3360 2540 3420
rect 2594 3360 2604 3420
rect 1904 3040 2604 3360
rect 3270 2380 3970 4400
rect 550 1680 3970 2380
rect 4570 2350 4610 5120
rect 4680 4100 4720 5210
rect 4770 5010 4810 5530
rect 4860 5400 4900 5820
rect 4930 5690 5010 5700
rect 4930 5630 4940 5690
rect 5000 5630 5010 5690
rect 4930 5620 5010 5630
rect 4840 5390 4920 5400
rect 4840 5330 4850 5390
rect 4910 5330 4920 5390
rect 4840 5320 4920 5330
rect 4750 5000 4830 5010
rect 4750 4940 4760 5000
rect 4820 4940 4830 5000
rect 4750 4930 4830 4940
rect 4660 4090 4740 4100
rect 4660 4030 4670 4090
rect 4730 4030 4740 4090
rect 4660 4020 4740 4030
rect 4680 3430 4720 4020
rect 4860 3770 4900 5320
rect 4950 4760 4990 5620
rect 4930 4750 5010 4760
rect 4930 4690 4940 4750
rect 5000 4690 5010 4750
rect 4930 4680 5010 4690
rect 5040 4300 5080 7530
rect 9310 7520 9390 7530
rect 10270 7590 10370 7610
rect 10270 7530 10290 7590
rect 10350 7530 10370 7590
rect 5380 7480 5460 7490
rect 5380 7420 5390 7480
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7480 6870 7500
rect 6770 7420 6790 7480
rect 6850 7420 6870 7480
rect 6770 7400 6870 7420
rect 9220 7480 9300 7490
rect 9220 7420 9230 7480
rect 9290 7420 9300 7480
rect 9220 7410 9300 7420
rect 8560 7380 8640 7390
rect 8560 7320 8570 7380
rect 8630 7320 8640 7380
rect 8560 7310 8640 7320
rect 5110 7280 5190 7290
rect 5110 7220 5120 7280
rect 5180 7220 5190 7280
rect 5110 7210 5190 7220
rect 6620 7270 6700 7280
rect 6620 7210 6630 7270
rect 6690 7210 6700 7270
rect 5130 6520 5170 7210
rect 6620 7200 6700 7210
rect 6400 7180 6480 7190
rect 6400 7120 6410 7180
rect 6470 7120 6480 7180
rect 6400 7110 6480 7120
rect 6420 7070 6460 7110
rect 6640 7070 6680 7200
rect 8120 7180 8200 7190
rect 8120 7120 8130 7180
rect 8190 7120 8200 7180
rect 8120 7110 8200 7120
rect 8140 7070 8180 7110
rect 8580 7070 8620 7310
rect 9130 7180 9210 7190
rect 9130 7120 9140 7180
rect 9200 7120 9210 7180
rect 9130 7110 9210 7120
rect 6070 7060 6150 7070
rect 6070 7000 6080 7060
rect 6140 7000 6150 7060
rect 6070 6990 6150 7000
rect 6290 7060 6370 7070
rect 6290 7000 6300 7060
rect 6360 7000 6370 7060
rect 6290 6990 6370 7000
rect 6410 7050 6470 7070
rect 6410 7010 6420 7050
rect 6460 7010 6470 7050
rect 6410 6990 6470 7010
rect 6510 7060 6590 7070
rect 6510 7000 6520 7060
rect 6580 7000 6590 7060
rect 6510 6990 6590 7000
rect 6630 7050 6690 7070
rect 6630 7010 6640 7050
rect 6680 7010 6690 7050
rect 6630 6990 6690 7010
rect 6730 7060 6810 7070
rect 6730 7000 6740 7060
rect 6800 7000 6810 7060
rect 6730 6990 6810 7000
rect 7350 7060 7430 7070
rect 7350 7000 7360 7060
rect 7420 7000 7430 7060
rect 7350 6990 7430 7000
rect 7570 7060 7650 7070
rect 7570 7000 7580 7060
rect 7640 7000 7650 7060
rect 7570 6990 7650 7000
rect 7790 7060 7870 7070
rect 7790 7000 7800 7060
rect 7860 7000 7870 7060
rect 7790 6990 7870 7000
rect 8010 7060 8090 7070
rect 8010 7000 8020 7060
rect 8080 7000 8090 7060
rect 8010 6990 8090 7000
rect 8130 7050 8190 7070
rect 8130 7010 8140 7050
rect 8180 7010 8190 7050
rect 8130 6990 8190 7010
rect 8230 7060 8310 7070
rect 8230 7000 8240 7060
rect 8300 7000 8310 7060
rect 8230 6990 8310 7000
rect 8450 7060 8530 7070
rect 8450 7000 8460 7060
rect 8520 7000 8530 7060
rect 8450 6990 8530 7000
rect 8570 7050 8630 7070
rect 8570 7010 8580 7050
rect 8620 7010 8630 7050
rect 8570 6990 8630 7010
rect 8670 7060 8750 7070
rect 8670 7000 8680 7060
rect 8740 7000 8750 7060
rect 8670 6990 8750 7000
rect 6180 6720 6260 6730
rect 6180 6660 6190 6720
rect 6250 6660 6260 6720
rect 6180 6650 6260 6660
rect 6400 6720 6480 6730
rect 6400 6660 6410 6720
rect 6470 6660 6480 6720
rect 6400 6650 6480 6660
rect 6620 6720 6700 6730
rect 6620 6660 6630 6720
rect 6690 6660 6700 6720
rect 6620 6650 6700 6660
rect 7460 6710 7540 6730
rect 7460 6670 7480 6710
rect 7520 6670 7540 6710
rect 7460 6650 7540 6670
rect 7680 6720 7760 6730
rect 7680 6660 7690 6720
rect 7750 6660 7760 6720
rect 7680 6650 7760 6660
rect 7900 6720 7980 6730
rect 7900 6660 7910 6720
rect 7970 6660 7980 6720
rect 7900 6650 7980 6660
rect 8120 6720 8200 6730
rect 8120 6660 8130 6720
rect 8190 6660 8200 6720
rect 8120 6650 8200 6660
rect 8340 6720 8420 6730
rect 8340 6660 8350 6720
rect 8410 6660 8420 6720
rect 8340 6650 8420 6660
rect 8560 6710 8640 6730
rect 8560 6670 8580 6710
rect 8620 6670 8640 6710
rect 8560 6650 8640 6670
rect 5110 6510 5190 6520
rect 5110 6450 5120 6510
rect 5180 6450 5190 6510
rect 5110 6440 5190 6450
rect 5220 6510 5300 6520
rect 5220 6450 5230 6510
rect 5290 6450 5300 6510
rect 5220 6440 5300 6450
rect 5110 6330 5190 6340
rect 5110 6270 5120 6330
rect 5180 6270 5190 6330
rect 5110 6260 5190 6270
rect 5020 4290 5100 4300
rect 5020 4230 5030 4290
rect 5090 4230 5100 4290
rect 5020 4220 5100 4230
rect 4840 3760 4920 3770
rect 4840 3700 4850 3760
rect 4910 3700 4920 3760
rect 4840 3690 4920 3700
rect 4660 3420 4740 3430
rect 4660 3360 4670 3420
rect 4730 3360 4740 3420
rect 4660 3350 4740 3360
rect 4550 2340 4630 2350
rect 4550 2280 4560 2340
rect 4620 2280 4630 2340
rect 4550 2270 4630 2280
rect 5130 1430 5170 6260
rect 5240 5110 5280 6440
rect 6120 6420 6200 6430
rect 6120 6360 6130 6420
rect 6190 6360 6200 6420
rect 6120 6350 6200 6360
rect 5650 6050 5730 6060
rect 5650 5990 5660 6050
rect 5720 5990 5730 6050
rect 5650 5980 5730 5990
rect 6140 5940 6180 6350
rect 7480 6340 7520 6650
rect 7460 6330 7540 6340
rect 7460 6270 7470 6330
rect 7530 6270 7540 6330
rect 7460 6260 7540 6270
rect 8140 6260 8180 6650
rect 8580 6330 8620 6650
rect 9150 6640 9190 7110
rect 9130 6630 9210 6640
rect 9130 6570 9140 6630
rect 9200 6570 9210 6630
rect 9130 6560 9210 6570
rect 9240 6530 9280 7410
rect 9220 6520 9300 6530
rect 9220 6460 9230 6520
rect 9290 6460 9300 6520
rect 9220 6450 9300 6460
rect 9330 6420 9370 7520
rect 10270 7510 10370 7530
rect 29970 7590 30050 7600
rect 29970 7530 29980 7590
rect 30040 7530 30050 7590
rect 29970 7520 30050 7530
rect 31880 7590 31960 7600
rect 31880 7530 31890 7590
rect 31950 7530 31960 7590
rect 31880 7520 31960 7530
rect 29880 7480 29960 7490
rect 29880 7420 29890 7480
rect 29950 7420 29960 7480
rect 29880 7410 29960 7420
rect 29900 7380 29940 7410
rect 29990 7380 30030 7520
rect 32720 7380 32760 7680
rect 38880 7630 38890 7690
rect 38950 7630 38960 7690
rect 38880 7620 38960 7630
rect 33270 7590 33370 7610
rect 33270 7530 33290 7590
rect 33350 7530 33370 7590
rect 35020 7600 35100 7610
rect 35020 7540 35030 7600
rect 35090 7540 35100 7600
rect 35020 7530 35100 7540
rect 39310 7590 39390 7600
rect 39310 7530 39320 7590
rect 39380 7530 39390 7590
rect 33270 7510 33370 7530
rect 35040 7380 35080 7530
rect 39310 7520 39390 7530
rect 40270 7590 40370 7610
rect 40270 7530 40290 7590
rect 40350 7530 40370 7590
rect 35380 7480 35460 7490
rect 35380 7420 35390 7480
rect 35450 7420 35460 7480
rect 35380 7410 35460 7420
rect 36770 7480 36870 7500
rect 36770 7420 36790 7480
rect 36850 7420 36870 7480
rect 36770 7400 36870 7420
rect 39220 7480 39300 7490
rect 39220 7420 39230 7480
rect 39290 7420 39300 7480
rect 39220 7410 39300 7420
rect 38560 7380 38640 7390
rect 38560 7320 38570 7380
rect 38630 7320 38640 7380
rect 38560 7310 38640 7320
rect 9840 7180 9920 7190
rect 9840 7120 9850 7180
rect 9910 7120 9920 7180
rect 9840 7110 9920 7120
rect 9860 7070 9900 7110
rect 9510 7060 9590 7070
rect 9510 7000 9520 7060
rect 9580 7000 9590 7060
rect 9510 6990 9590 7000
rect 9730 7060 9810 7070
rect 9730 7000 9740 7060
rect 9800 7000 9810 7060
rect 9730 6990 9810 7000
rect 9850 7050 9910 7070
rect 9850 7010 9860 7050
rect 9900 7010 9910 7050
rect 9850 6990 9910 7010
rect 9950 7060 10030 7070
rect 9950 7000 9960 7060
rect 10020 7000 10030 7060
rect 9950 6990 10030 7000
rect 10170 7060 10250 7070
rect 10170 7000 10180 7060
rect 10240 7000 10250 7060
rect 10170 6990 10250 7000
rect 9620 6720 9700 6730
rect 9620 6660 9630 6720
rect 9690 6660 9700 6720
rect 9620 6650 9700 6660
rect 9840 6720 9920 6730
rect 9840 6660 9850 6720
rect 9910 6660 9920 6720
rect 9840 6650 9920 6660
rect 10060 6720 10140 6730
rect 10060 6660 10070 6720
rect 10130 6660 10140 6720
rect 10060 6650 10140 6660
rect 9940 6610 10020 6620
rect 9940 6550 9950 6610
rect 10010 6550 10020 6610
rect 9940 6540 10020 6550
rect 9310 6410 9390 6420
rect 9310 6350 9320 6410
rect 9380 6350 9390 6410
rect 9310 6340 9390 6350
rect 8560 6320 8640 6330
rect 8560 6260 8570 6320
rect 8630 6260 8640 6320
rect 8120 6250 8200 6260
rect 8560 6250 8640 6260
rect 8120 6190 8130 6250
rect 8190 6190 8200 6250
rect 8120 6180 8200 6190
rect 6500 6130 6580 6140
rect 6500 6070 6510 6130
rect 6570 6070 6580 6130
rect 6500 6060 6580 6070
rect 6860 6130 6940 6140
rect 6860 6070 6870 6130
rect 6930 6070 6940 6130
rect 6860 6060 6940 6070
rect 7220 6130 7300 6140
rect 7220 6070 7230 6130
rect 7290 6070 7300 6130
rect 7220 6060 7300 6070
rect 7580 6130 7660 6140
rect 7580 6070 7590 6130
rect 7650 6070 7660 6130
rect 7580 6060 7660 6070
rect 7940 6130 8020 6140
rect 7940 6070 7950 6130
rect 8010 6070 8020 6130
rect 7940 6060 8020 6070
rect 8300 6130 8380 6140
rect 8300 6070 8310 6130
rect 8370 6070 8380 6130
rect 8300 6060 8380 6070
rect 8660 6130 8740 6140
rect 8660 6070 8670 6130
rect 8730 6070 8740 6130
rect 8660 6060 8740 6070
rect 9020 6130 9100 6140
rect 9020 6070 9030 6130
rect 9090 6070 9100 6130
rect 9020 6060 9100 6070
rect 9380 6130 9460 6140
rect 9380 6070 9390 6130
rect 9450 6070 9460 6130
rect 9380 6060 9460 6070
rect 9740 6130 9820 6140
rect 9740 6070 9750 6130
rect 9810 6070 9820 6130
rect 9740 6060 9820 6070
rect 5650 5930 5730 5940
rect 5650 5870 5660 5930
rect 5720 5870 5730 5930
rect 5650 5860 5730 5870
rect 6120 5930 6200 5940
rect 6120 5870 6130 5930
rect 6190 5870 6200 5930
rect 6120 5860 6200 5870
rect 5520 5590 5600 5600
rect 5520 5530 5530 5590
rect 5590 5530 5600 5590
rect 5520 5520 5600 5530
rect 5650 5580 5730 5600
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 5780 5590 5860 5600
rect 5780 5530 5790 5590
rect 5850 5530 5860 5590
rect 5780 5520 5860 5530
rect 5670 5200 5710 5520
rect 6140 5290 6180 5860
rect 6240 5590 6320 5600
rect 6240 5530 6250 5590
rect 6310 5530 6320 5590
rect 6240 5520 6320 5530
rect 6120 5280 6200 5290
rect 6120 5220 6130 5280
rect 6190 5220 6200 5280
rect 6120 5210 6200 5220
rect 5650 5190 5730 5200
rect 5650 5130 5660 5190
rect 5720 5130 5730 5190
rect 5650 5120 5730 5130
rect 5220 5100 5300 5110
rect 5220 5040 5230 5100
rect 5290 5040 5300 5100
rect 5220 5030 5300 5040
rect 5640 4870 5720 4880
rect 5640 4810 5650 4870
rect 5710 4810 5720 4870
rect 5640 4800 5720 4810
rect 5880 4870 5960 4880
rect 5880 4810 5890 4870
rect 5950 4810 5960 4870
rect 5880 4800 5960 4810
rect 6120 4870 6200 4880
rect 6120 4810 6130 4870
rect 6190 4810 6200 4870
rect 6120 4800 6200 4810
rect 5660 4760 5700 4800
rect 5900 4760 5940 4800
rect 6140 4760 6180 4800
rect 6260 4760 6300 5520
rect 6680 5380 6760 5400
rect 6680 5340 6700 5380
rect 6740 5340 6760 5380
rect 6680 5320 6760 5340
rect 7040 5380 7120 5400
rect 7040 5340 7060 5380
rect 7100 5340 7120 5380
rect 7040 5320 7120 5340
rect 7400 5380 7480 5400
rect 7400 5340 7420 5380
rect 7460 5340 7480 5380
rect 7400 5320 7480 5340
rect 7760 5390 7840 5400
rect 7760 5330 7770 5390
rect 7830 5330 7840 5390
rect 7760 5320 7840 5330
rect 7940 5380 8020 5400
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 8120 5380 8200 5400
rect 8120 5340 8140 5380
rect 8180 5340 8200 5380
rect 8120 5320 8200 5340
rect 8480 5390 8560 5400
rect 8480 5330 8490 5390
rect 8550 5330 8560 5390
rect 8480 5320 8560 5330
rect 8840 5380 8920 5400
rect 8840 5340 8860 5380
rect 8900 5340 8920 5380
rect 8840 5320 8920 5340
rect 9200 5380 9280 5400
rect 9200 5340 9220 5380
rect 9260 5340 9280 5380
rect 9200 5320 9280 5340
rect 9380 5380 9460 5400
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 9560 5380 9640 5400
rect 9560 5340 9580 5380
rect 9620 5340 9640 5380
rect 9560 5320 9640 5340
rect 6700 5110 6740 5320
rect 7060 5200 7100 5320
rect 7420 5290 7460 5320
rect 7400 5280 7480 5290
rect 7400 5220 7410 5280
rect 7470 5220 7480 5280
rect 7400 5210 7480 5220
rect 7040 5190 7120 5200
rect 7040 5130 7050 5190
rect 7110 5130 7120 5190
rect 7040 5120 7120 5130
rect 6680 5100 6760 5110
rect 6680 5040 6690 5100
rect 6750 5040 6760 5100
rect 6680 5030 6760 5040
rect 6360 4870 6440 4880
rect 6360 4810 6370 4870
rect 6430 4810 6440 4870
rect 6360 4800 6440 4810
rect 6600 4870 6680 4880
rect 6600 4810 6610 4870
rect 6670 4810 6680 4870
rect 6600 4800 6680 4810
rect 6840 4870 6920 4880
rect 6840 4810 6850 4870
rect 6910 4810 6920 4870
rect 6840 4800 6920 4810
rect 7080 4870 7160 4880
rect 7080 4810 7090 4870
rect 7150 4810 7160 4870
rect 7080 4800 7160 4810
rect 7320 4870 7400 4880
rect 7320 4810 7330 4870
rect 7390 4810 7400 4870
rect 7320 4800 7400 4810
rect 7560 4870 7640 4880
rect 7560 4810 7570 4870
rect 7630 4810 7640 4870
rect 7560 4800 7640 4810
rect 6380 4760 6420 4800
rect 6620 4760 6660 4800
rect 6860 4760 6900 4800
rect 7100 4760 7140 4800
rect 7340 4760 7380 4800
rect 7580 4760 7620 4800
rect 7960 4760 8000 5320
rect 8140 5110 8180 5320
rect 8860 5290 8900 5320
rect 8840 5280 8920 5290
rect 8840 5220 8850 5280
rect 8910 5220 8920 5280
rect 8840 5210 8920 5220
rect 9220 5200 9260 5320
rect 9400 5200 9440 5320
rect 9200 5190 9280 5200
rect 9200 5130 9210 5190
rect 9270 5130 9280 5190
rect 9200 5120 9280 5130
rect 9380 5190 9460 5200
rect 9380 5130 9390 5190
rect 9450 5130 9460 5190
rect 9380 5120 9460 5130
rect 9580 5110 9620 5320
rect 8120 5100 8200 5110
rect 8120 5040 8130 5100
rect 8190 5040 8200 5100
rect 8120 5030 8200 5040
rect 9560 5100 9640 5110
rect 9560 5040 9570 5100
rect 9630 5040 9640 5100
rect 9560 5030 9640 5040
rect 9960 5010 10000 6540
rect 10120 6520 10200 6530
rect 10120 6460 10130 6520
rect 10190 6460 10200 6520
rect 10120 6450 10200 6460
rect 10030 6410 10110 6420
rect 10030 6350 10040 6410
rect 10100 6350 10110 6410
rect 10030 6340 10110 6350
rect 10050 5200 10090 6340
rect 10140 5310 10180 6450
rect 11230 6320 11310 6330
rect 11230 6260 11240 6320
rect 11300 6260 11310 6320
rect 11230 6250 11310 6260
rect 10580 6050 10660 6080
rect 10580 5990 10590 6050
rect 10650 5990 10660 6050
rect 10580 5980 10660 5990
rect 10600 5940 10640 5980
rect 10580 5930 10660 5940
rect 10580 5870 10590 5930
rect 10650 5870 10660 5930
rect 10580 5860 10660 5870
rect 10450 5590 10530 5600
rect 10450 5530 10460 5590
rect 10520 5530 10530 5590
rect 10450 5520 10530 5530
rect 10580 5580 10660 5600
rect 10580 5540 10600 5580
rect 10640 5540 10660 5580
rect 10580 5520 10660 5540
rect 10710 5590 10790 5600
rect 10710 5530 10720 5590
rect 10780 5530 10790 5590
rect 10710 5520 10790 5530
rect 10120 5300 10200 5310
rect 10120 5240 10130 5300
rect 10190 5240 10200 5300
rect 10120 5230 10200 5240
rect 10030 5190 10110 5200
rect 10030 5130 10040 5190
rect 10100 5130 10110 5190
rect 10030 5120 10110 5130
rect 10600 5010 10640 5520
rect 11050 5300 11130 5310
rect 11050 5240 11060 5300
rect 11120 5240 11130 5300
rect 11050 5230 11130 5240
rect 8560 5000 8640 5010
rect 8560 4940 8570 5000
rect 8630 4940 8640 5000
rect 8560 4930 8640 4940
rect 9940 5000 10020 5010
rect 9940 4940 9950 5000
rect 10010 4940 10020 5000
rect 9940 4930 10020 4940
rect 10580 5000 10660 5010
rect 10580 4940 10590 5000
rect 10650 4940 10660 5000
rect 10580 4930 10660 4940
rect 8580 4760 8620 4930
rect 8680 4870 8760 4880
rect 8680 4810 8690 4870
rect 8750 4810 8760 4870
rect 8680 4800 8760 4810
rect 8920 4870 9000 4880
rect 8920 4810 8930 4870
rect 8990 4810 9000 4870
rect 8920 4800 9000 4810
rect 9160 4870 9240 4880
rect 9160 4810 9170 4870
rect 9230 4810 9240 4870
rect 9160 4800 9240 4810
rect 9400 4870 9480 4880
rect 9400 4810 9410 4870
rect 9470 4810 9480 4870
rect 9400 4800 9480 4810
rect 9640 4870 9720 4880
rect 9640 4810 9650 4870
rect 9710 4810 9720 4870
rect 9640 4800 9720 4810
rect 9880 4870 9960 4880
rect 9880 4810 9890 4870
rect 9950 4810 9960 4870
rect 9880 4800 9960 4810
rect 10120 4870 10200 4880
rect 10120 4810 10130 4870
rect 10190 4810 10200 4870
rect 10120 4800 10200 4810
rect 10360 4870 10440 4880
rect 10360 4810 10370 4870
rect 10430 4810 10440 4870
rect 10360 4800 10440 4810
rect 10600 4870 10680 4880
rect 10600 4810 10610 4870
rect 10670 4810 10680 4870
rect 10600 4800 10680 4810
rect 8700 4760 8740 4800
rect 8940 4760 8980 4800
rect 9180 4760 9220 4800
rect 9420 4760 9460 4800
rect 9660 4760 9700 4800
rect 9900 4760 9940 4800
rect 10140 4760 10180 4800
rect 10380 4760 10420 4800
rect 10620 4760 10660 4800
rect 5520 4750 5600 4760
rect 5520 4690 5530 4750
rect 5590 4690 5600 4750
rect 5520 4680 5600 4690
rect 5650 4740 5710 4760
rect 5650 4700 5660 4740
rect 5700 4700 5710 4740
rect 5650 4680 5710 4700
rect 5890 4740 5950 4760
rect 5890 4700 5900 4740
rect 5940 4700 5950 4740
rect 5890 4680 5950 4700
rect 6130 4740 6190 4760
rect 6130 4700 6140 4740
rect 6180 4700 6190 4740
rect 6130 4680 6190 4700
rect 6240 4750 6320 4760
rect 6240 4690 6250 4750
rect 6310 4690 6320 4750
rect 6240 4680 6320 4690
rect 6370 4740 6430 4760
rect 6370 4700 6380 4740
rect 6420 4700 6430 4740
rect 6370 4680 6430 4700
rect 6610 4740 6670 4760
rect 6610 4700 6620 4740
rect 6660 4700 6670 4740
rect 6610 4680 6670 4700
rect 6850 4740 6910 4760
rect 6850 4700 6860 4740
rect 6900 4700 6910 4740
rect 6850 4680 6910 4700
rect 6960 4750 7040 4760
rect 6960 4690 6970 4750
rect 7030 4690 7040 4750
rect 6960 4680 7040 4690
rect 7090 4740 7150 4760
rect 7090 4700 7100 4740
rect 7140 4700 7150 4740
rect 7090 4680 7150 4700
rect 7330 4740 7390 4760
rect 7330 4700 7340 4740
rect 7380 4700 7390 4740
rect 7330 4680 7390 4700
rect 7570 4740 7630 4760
rect 7570 4700 7580 4740
rect 7620 4700 7630 4740
rect 7570 4680 7630 4700
rect 7680 4750 7760 4760
rect 7680 4690 7690 4750
rect 7750 4690 7760 4750
rect 7680 4680 7760 4690
rect 7940 4750 8020 4760
rect 7940 4690 7950 4750
rect 8010 4690 8020 4750
rect 7940 4680 8020 4690
rect 8300 4750 8380 4760
rect 8300 4690 8310 4750
rect 8370 4690 8380 4750
rect 8300 4680 8380 4690
rect 8560 4750 8640 4760
rect 8560 4690 8570 4750
rect 8630 4690 8640 4750
rect 8560 4680 8640 4690
rect 8690 4740 8750 4760
rect 8690 4700 8700 4740
rect 8740 4700 8750 4740
rect 8690 4680 8750 4700
rect 8930 4740 8990 4760
rect 8930 4700 8940 4740
rect 8980 4700 8990 4740
rect 8930 4680 8990 4700
rect 9170 4740 9230 4760
rect 9170 4700 9180 4740
rect 9220 4700 9230 4740
rect 9170 4680 9230 4700
rect 9280 4750 9360 4760
rect 9280 4690 9290 4750
rect 9350 4690 9360 4750
rect 9280 4680 9360 4690
rect 9410 4740 9470 4760
rect 9410 4700 9420 4740
rect 9460 4700 9470 4740
rect 9410 4680 9470 4700
rect 9650 4740 9710 4760
rect 9650 4700 9660 4740
rect 9700 4700 9710 4740
rect 9650 4680 9710 4700
rect 9890 4740 9950 4760
rect 9890 4700 9900 4740
rect 9940 4700 9950 4740
rect 9890 4680 9950 4700
rect 10000 4750 10080 4760
rect 10000 4690 10010 4750
rect 10070 4690 10080 4750
rect 10000 4680 10080 4690
rect 10130 4740 10190 4760
rect 10130 4700 10140 4740
rect 10180 4700 10190 4740
rect 10130 4680 10190 4700
rect 10370 4740 10430 4760
rect 10370 4700 10380 4740
rect 10420 4700 10430 4740
rect 10370 4680 10430 4700
rect 10610 4740 10670 4760
rect 10610 4700 10620 4740
rect 10660 4700 10670 4740
rect 10610 4680 10670 4700
rect 10720 4750 10800 4760
rect 10720 4690 10730 4750
rect 10790 4690 10800 4750
rect 10720 4680 10800 4690
rect 5580 4400 5660 4420
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4410 5840 4420
rect 5760 4350 5770 4410
rect 5830 4350 5840 4410
rect 5760 4340 5840 4350
rect 6000 4400 6080 4420
rect 6000 4360 6020 4400
rect 6060 4360 6080 4400
rect 6000 4340 6080 4360
rect 6240 4400 6320 4420
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4410 6560 4420
rect 6480 4350 6490 4410
rect 6550 4350 6560 4410
rect 6480 4340 6560 4350
rect 6720 4400 6800 4420
rect 6720 4360 6740 4400
rect 6780 4360 6800 4400
rect 6720 4340 6800 4360
rect 6960 4400 7040 4420
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4410 7280 4420
rect 7200 4350 7210 4410
rect 7270 4350 7280 4410
rect 7200 4340 7280 4350
rect 7440 4400 7520 4420
rect 7440 4360 7460 4400
rect 7500 4360 7520 4400
rect 7440 4340 7520 4360
rect 7630 4400 7690 4420
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 5600 4300 5640 4340
rect 6020 4300 6060 4340
rect 6260 4300 6300 4340
rect 5580 4290 5660 4300
rect 5580 4230 5590 4290
rect 5650 4230 5660 4290
rect 5580 4220 5660 4230
rect 6000 4290 6080 4300
rect 6000 4230 6010 4290
rect 6070 4230 6080 4290
rect 6000 4220 6080 4230
rect 6240 4290 6320 4300
rect 6240 4230 6250 4290
rect 6310 4230 6320 4290
rect 6240 4220 6320 4230
rect 6520 4130 6560 4340
rect 6740 4300 6780 4340
rect 6980 4300 7020 4340
rect 7460 4300 7500 4340
rect 7640 4300 7680 4340
rect 6720 4290 6800 4300
rect 6720 4230 6730 4290
rect 6790 4230 6800 4290
rect 6720 4220 6800 4230
rect 6960 4290 7040 4300
rect 6960 4230 6970 4290
rect 7030 4230 7040 4290
rect 6960 4220 7040 4230
rect 7440 4290 7520 4300
rect 7440 4230 7450 4290
rect 7510 4230 7520 4290
rect 7440 4220 7520 4230
rect 7620 4290 7700 4300
rect 7620 4230 7630 4290
rect 7690 4230 7700 4290
rect 7620 4220 7700 4230
rect 6500 4120 6580 4130
rect 6380 4090 6460 4100
rect 6380 4030 6390 4090
rect 6450 4030 6460 4090
rect 6500 4060 6510 4120
rect 6570 4060 6580 4120
rect 6500 4050 6580 4060
rect 6380 4020 6460 4030
rect 6520 4010 6560 4050
rect 6740 4010 6780 4220
rect 6980 4120 7060 4130
rect 6980 4060 6990 4120
rect 7050 4060 7060 4120
rect 6980 4050 7060 4060
rect 7460 4120 7540 4130
rect 7460 4060 7470 4120
rect 7530 4060 7540 4120
rect 7460 4050 7540 4060
rect 7000 4010 7040 4050
rect 7480 4010 7520 4050
rect 6260 4000 6340 4010
rect 6260 3940 6270 4000
rect 6330 3940 6340 4000
rect 6260 3930 6340 3940
rect 6510 3990 6570 4010
rect 6510 3950 6520 3990
rect 6560 3950 6570 3990
rect 6510 3930 6570 3950
rect 6740 4000 6820 4010
rect 6740 3940 6750 4000
rect 6810 3940 6820 4000
rect 6740 3930 6820 3940
rect 6990 3990 7050 4010
rect 6990 3950 7000 3990
rect 7040 3950 7050 3990
rect 6990 3930 7050 3950
rect 7220 4000 7300 4010
rect 7220 3940 7230 4000
rect 7290 3940 7300 4000
rect 7220 3930 7300 3940
rect 7470 3990 7530 4010
rect 7470 3950 7480 3990
rect 7520 3950 7530 3990
rect 7470 3930 7530 3950
rect 7580 3880 7660 3890
rect 7580 3820 7590 3880
rect 7650 3820 7660 3880
rect 7580 3810 7660 3820
rect 6260 3760 6340 3770
rect 6260 3700 6270 3760
rect 6330 3700 6340 3760
rect 6260 3690 6340 3700
rect 6390 3750 6450 3770
rect 6390 3710 6400 3750
rect 6440 3710 6450 3750
rect 6390 3690 6450 3710
rect 6630 3750 6690 3770
rect 6630 3710 6640 3750
rect 6680 3710 6690 3750
rect 6630 3690 6690 3710
rect 6870 3750 6930 3770
rect 6870 3710 6880 3750
rect 6920 3710 6930 3750
rect 6870 3690 6930 3710
rect 7110 3750 7170 3770
rect 7110 3710 7120 3750
rect 7160 3710 7170 3750
rect 7110 3690 7170 3710
rect 7350 3750 7410 3770
rect 7350 3710 7360 3750
rect 7400 3710 7410 3750
rect 7350 3690 7410 3710
rect 6400 3650 6440 3690
rect 6640 3650 6680 3690
rect 6880 3650 6920 3690
rect 7120 3650 7160 3690
rect 7360 3650 7400 3690
rect 5780 3640 5860 3650
rect 5780 3580 5790 3640
rect 5850 3580 5860 3640
rect 5780 3570 5860 3580
rect 6380 3640 6460 3650
rect 6380 3580 6390 3640
rect 6450 3580 6460 3640
rect 6380 3570 6460 3580
rect 6620 3640 6700 3650
rect 6620 3580 6630 3640
rect 6690 3580 6700 3640
rect 6620 3570 6700 3580
rect 6860 3640 6940 3650
rect 6860 3580 6870 3640
rect 6930 3580 6940 3640
rect 6860 3570 6940 3580
rect 7100 3640 7180 3650
rect 7100 3580 7110 3640
rect 7170 3580 7180 3640
rect 7100 3570 7180 3580
rect 7340 3640 7420 3650
rect 7340 3580 7350 3640
rect 7410 3580 7420 3640
rect 7340 3570 7420 3580
rect 5800 3420 5840 3570
rect 5960 3440 6040 3450
rect 5780 3400 5860 3420
rect 5780 3360 5800 3400
rect 5840 3360 5860 3400
rect 5960 3380 5970 3440
rect 6030 3380 6040 3440
rect 5960 3370 6040 3380
rect 6200 3440 6280 3450
rect 6200 3380 6210 3440
rect 6270 3380 6280 3440
rect 6200 3370 6280 3380
rect 6440 3440 6520 3450
rect 6440 3380 6450 3440
rect 6510 3380 6520 3440
rect 6440 3370 6520 3380
rect 6680 3440 6760 3450
rect 6680 3380 6690 3440
rect 6750 3380 6760 3440
rect 6680 3370 6760 3380
rect 7160 3440 7240 3450
rect 7160 3380 7170 3440
rect 7230 3380 7240 3440
rect 7160 3370 7240 3380
rect 7400 3440 7480 3450
rect 7400 3380 7410 3440
rect 7470 3380 7480 3440
rect 7400 3370 7480 3380
rect 7640 3440 7720 3450
rect 7640 3380 7650 3440
rect 7710 3380 7720 3440
rect 7960 3420 8000 4680
rect 8120 3880 8200 3890
rect 8120 3820 8130 3880
rect 8190 3820 8200 3880
rect 8120 3810 8200 3820
rect 7640 3370 7720 3380
rect 7940 3400 8020 3420
rect 5780 3340 5860 3360
rect 7940 3360 7960 3400
rect 8000 3360 8020 3400
rect 7940 3340 8020 3360
rect 8140 2820 8180 3810
rect 8320 3420 8360 4680
rect 8630 4400 8690 4420
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 8800 4400 8880 4420
rect 8800 4360 8820 4400
rect 8860 4360 8880 4400
rect 8800 4340 8880 4360
rect 9040 4410 9120 4420
rect 9040 4350 9050 4410
rect 9110 4350 9120 4410
rect 9040 4340 9120 4350
rect 9280 4400 9360 4420
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9520 4400 9600 4420
rect 9520 4360 9540 4400
rect 9580 4360 9600 4400
rect 9520 4340 9600 4360
rect 9760 4410 9840 4420
rect 9760 4350 9770 4410
rect 9830 4350 9840 4410
rect 9760 4340 9840 4350
rect 10000 4400 10080 4420
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10240 4400 10320 4420
rect 10240 4360 10260 4400
rect 10300 4360 10320 4400
rect 10240 4340 10320 4360
rect 10480 4410 10560 4420
rect 10480 4350 10490 4410
rect 10550 4350 10560 4410
rect 10480 4340 10560 4350
rect 10660 4400 10740 4420
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 8640 4300 8680 4340
rect 8820 4300 8860 4340
rect 9300 4300 9340 4340
rect 9540 4300 9580 4340
rect 8620 4290 8700 4300
rect 8620 4230 8630 4290
rect 8690 4230 8700 4290
rect 8620 4220 8700 4230
rect 8800 4290 8880 4300
rect 8800 4230 8810 4290
rect 8870 4230 8880 4290
rect 8800 4220 8880 4230
rect 9280 4290 9360 4300
rect 9280 4230 9290 4290
rect 9350 4230 9360 4290
rect 9280 4220 9360 4230
rect 9520 4290 9600 4300
rect 9520 4230 9530 4290
rect 9590 4230 9600 4290
rect 9520 4220 9600 4230
rect 8780 4120 8860 4130
rect 8780 4060 8790 4120
rect 8850 4060 8860 4120
rect 8780 4050 8860 4060
rect 9260 4120 9340 4130
rect 9260 4060 9270 4120
rect 9330 4060 9340 4120
rect 9260 4050 9340 4060
rect 8800 4010 8840 4050
rect 9280 4010 9320 4050
rect 9520 4010 9560 4220
rect 9760 4130 9800 4340
rect 10020 4300 10060 4340
rect 10260 4300 10300 4340
rect 10680 4300 10720 4340
rect 11070 4300 11110 5230
rect 11140 5100 11220 5110
rect 11140 5040 11150 5100
rect 11210 5040 11220 5100
rect 11140 5030 11220 5040
rect 10000 4290 10080 4300
rect 10000 4230 10010 4290
rect 10070 4230 10080 4290
rect 10000 4220 10080 4230
rect 10240 4290 10320 4300
rect 10240 4230 10250 4290
rect 10310 4230 10320 4290
rect 10240 4220 10320 4230
rect 10660 4290 10740 4300
rect 10660 4230 10670 4290
rect 10730 4230 10740 4290
rect 10660 4220 10740 4230
rect 11050 4290 11130 4300
rect 11050 4230 11060 4290
rect 11120 4230 11130 4290
rect 11050 4220 11130 4230
rect 9740 4120 9820 4130
rect 9740 4060 9750 4120
rect 9810 4060 9820 4120
rect 11160 4100 11200 5030
rect 9740 4050 9820 4060
rect 9860 4090 9940 4100
rect 9760 4010 9800 4050
rect 9860 4030 9870 4090
rect 9930 4030 9940 4090
rect 9860 4020 9940 4030
rect 11140 4090 11220 4100
rect 11140 4030 11150 4090
rect 11210 4030 11220 4090
rect 11140 4020 11220 4030
rect 8790 3990 8850 4010
rect 8790 3950 8800 3990
rect 8840 3950 8850 3990
rect 8790 3930 8850 3950
rect 9020 4000 9100 4010
rect 9020 3940 9030 4000
rect 9090 3940 9100 4000
rect 9020 3930 9100 3940
rect 9270 3990 9330 4010
rect 9270 3950 9280 3990
rect 9320 3950 9330 3990
rect 9270 3930 9330 3950
rect 9500 4000 9580 4010
rect 9500 3940 9510 4000
rect 9570 3940 9580 4000
rect 9500 3930 9580 3940
rect 9750 3990 9810 4010
rect 9750 3950 9760 3990
rect 9800 3950 9810 3990
rect 9750 3930 9810 3950
rect 9980 4000 10060 4010
rect 9980 3940 9990 4000
rect 10050 3940 10060 4000
rect 9980 3930 10060 3940
rect 8660 3880 8740 3890
rect 8660 3820 8670 3880
rect 8730 3820 8740 3880
rect 8660 3810 8740 3820
rect 11250 3770 11290 6250
rect 38580 6200 38620 7310
rect 39240 6200 39280 7410
rect 39330 6200 39370 7520
rect 40270 7510 40370 7530
rect 36620 4270 36700 4280
rect 36620 4210 36630 4270
rect 36690 4210 36700 4270
rect 36620 4200 36700 4210
rect 36400 4180 36480 4190
rect 36400 4120 36410 4180
rect 36470 4120 36480 4180
rect 36400 4110 36480 4120
rect 36420 4070 36460 4110
rect 36640 4070 36680 4200
rect 38120 4180 38200 4190
rect 38120 4120 38130 4180
rect 38190 4120 38200 4180
rect 38120 4110 38200 4120
rect 38140 4070 38180 4110
rect 38580 4070 38620 4370
rect 39130 4180 39210 4190
rect 39130 4120 39140 4180
rect 39200 4120 39210 4180
rect 39130 4110 39210 4120
rect 36070 4060 36150 4070
rect 36070 4000 36080 4060
rect 36140 4000 36150 4060
rect 36070 3990 36150 4000
rect 36290 4060 36370 4070
rect 36290 4000 36300 4060
rect 36360 4000 36370 4060
rect 36290 3990 36370 4000
rect 36410 4050 36470 4070
rect 36410 4010 36420 4050
rect 36460 4010 36470 4050
rect 36410 3990 36470 4010
rect 36510 4060 36590 4070
rect 36510 4000 36520 4060
rect 36580 4000 36590 4060
rect 36510 3990 36590 4000
rect 36630 4050 36690 4070
rect 36630 4010 36640 4050
rect 36680 4010 36690 4050
rect 36630 3990 36690 4010
rect 36730 4060 36810 4070
rect 36730 4000 36740 4060
rect 36800 4000 36810 4060
rect 36730 3990 36810 4000
rect 37350 4060 37430 4070
rect 37350 4000 37360 4060
rect 37420 4000 37430 4060
rect 37350 3990 37430 4000
rect 37570 4060 37650 4070
rect 37570 4000 37580 4060
rect 37640 4000 37650 4060
rect 37570 3990 37650 4000
rect 37790 4060 37870 4070
rect 37790 4000 37800 4060
rect 37860 4000 37870 4060
rect 37790 3990 37870 4000
rect 38010 4060 38090 4070
rect 38010 4000 38020 4060
rect 38080 4000 38090 4060
rect 38010 3990 38090 4000
rect 38130 4050 38190 4070
rect 38130 4010 38140 4050
rect 38180 4010 38190 4050
rect 38130 3990 38190 4010
rect 38230 4060 38310 4070
rect 38230 4000 38240 4060
rect 38300 4000 38310 4060
rect 38230 3990 38310 4000
rect 38450 4060 38530 4070
rect 38450 4000 38460 4060
rect 38520 4000 38530 4060
rect 38450 3990 38530 4000
rect 38570 4050 38630 4070
rect 38570 4010 38580 4050
rect 38620 4010 38630 4050
rect 38570 3990 38630 4010
rect 38670 4060 38750 4070
rect 38670 4000 38680 4060
rect 38740 4000 38750 4060
rect 38670 3990 38750 4000
rect 8910 3750 8970 3770
rect 8910 3710 8920 3750
rect 8960 3710 8970 3750
rect 8910 3690 8970 3710
rect 9150 3750 9210 3770
rect 9150 3710 9160 3750
rect 9200 3710 9210 3750
rect 9150 3690 9210 3710
rect 9390 3750 9450 3770
rect 9390 3710 9400 3750
rect 9440 3710 9450 3750
rect 9390 3690 9450 3710
rect 9630 3750 9690 3770
rect 9630 3710 9640 3750
rect 9680 3710 9690 3750
rect 9630 3690 9690 3710
rect 9870 3750 9930 3770
rect 9870 3710 9880 3750
rect 9920 3710 9930 3750
rect 9870 3690 9930 3710
rect 9980 3760 10060 3770
rect 9980 3700 9990 3760
rect 10050 3700 10060 3760
rect 9980 3690 10060 3700
rect 11230 3760 11310 3770
rect 11230 3700 11240 3760
rect 11300 3700 11310 3760
rect 11230 3690 11310 3700
rect 36180 3720 36260 3730
rect 8920 3650 8960 3690
rect 9160 3650 9200 3690
rect 9400 3650 9440 3690
rect 9640 3650 9680 3690
rect 9880 3650 9920 3690
rect 36180 3660 36190 3720
rect 36250 3660 36260 3720
rect 36180 3650 36260 3660
rect 36400 3720 36480 3730
rect 36400 3660 36410 3720
rect 36470 3660 36480 3720
rect 36400 3650 36480 3660
rect 36620 3720 36700 3730
rect 36620 3660 36630 3720
rect 36690 3660 36700 3720
rect 36620 3650 36700 3660
rect 37460 3710 37540 3730
rect 37460 3670 37480 3710
rect 37520 3670 37540 3710
rect 37460 3650 37540 3670
rect 37680 3720 37760 3730
rect 37680 3660 37690 3720
rect 37750 3660 37760 3720
rect 37680 3650 37760 3660
rect 37900 3720 37980 3730
rect 37900 3660 37910 3720
rect 37970 3660 37980 3720
rect 37900 3650 37980 3660
rect 38120 3720 38200 3730
rect 38120 3660 38130 3720
rect 38190 3660 38200 3720
rect 38120 3650 38200 3660
rect 38340 3720 38420 3730
rect 38340 3660 38350 3720
rect 38410 3660 38420 3720
rect 38340 3650 38420 3660
rect 38560 3710 38640 3730
rect 38560 3670 38580 3710
rect 38620 3670 38640 3710
rect 38560 3650 38640 3670
rect 8900 3640 8980 3650
rect 8900 3580 8910 3640
rect 8970 3580 8980 3640
rect 8900 3570 8980 3580
rect 9140 3640 9220 3650
rect 9140 3580 9150 3640
rect 9210 3580 9220 3640
rect 9140 3570 9220 3580
rect 9380 3640 9460 3650
rect 9380 3580 9390 3640
rect 9450 3580 9460 3640
rect 9380 3570 9460 3580
rect 9620 3640 9700 3650
rect 9620 3580 9630 3640
rect 9690 3580 9700 3640
rect 9620 3570 9700 3580
rect 9860 3640 9940 3650
rect 9860 3580 9870 3640
rect 9930 3580 9940 3640
rect 9860 3570 9940 3580
rect 10460 3640 10540 3650
rect 10460 3580 10470 3640
rect 10530 3580 10540 3640
rect 10460 3570 10540 3580
rect 8600 3440 8680 3450
rect 8300 3400 8380 3420
rect 8300 3360 8320 3400
rect 8360 3360 8380 3400
rect 8600 3380 8610 3440
rect 8670 3380 8680 3440
rect 8600 3370 8680 3380
rect 8840 3440 8920 3450
rect 8840 3380 8850 3440
rect 8910 3380 8920 3440
rect 8840 3370 8920 3380
rect 9080 3440 9160 3450
rect 9080 3380 9090 3440
rect 9150 3380 9160 3440
rect 9080 3370 9160 3380
rect 9560 3440 9640 3450
rect 9560 3380 9570 3440
rect 9630 3380 9640 3440
rect 9560 3370 9640 3380
rect 9800 3440 9880 3450
rect 9800 3380 9810 3440
rect 9870 3380 9880 3440
rect 9800 3370 9880 3380
rect 10040 3440 10120 3450
rect 10040 3380 10050 3440
rect 10110 3380 10120 3440
rect 10040 3370 10120 3380
rect 10280 3440 10360 3450
rect 10280 3380 10290 3440
rect 10350 3380 10360 3440
rect 10480 3420 10520 3570
rect 10280 3370 10360 3380
rect 10460 3400 10540 3420
rect 8300 3340 8380 3360
rect 10460 3360 10480 3400
rect 10520 3360 10540 3400
rect 10460 3340 10540 3360
rect 6860 2810 6940 2820
rect 6860 2750 6870 2810
rect 6930 2750 6940 2810
rect 6860 2740 6940 2750
rect 8120 2810 8200 2820
rect 8120 2750 8130 2810
rect 8190 2750 8200 2810
rect 8120 2740 8200 2750
rect 9380 2810 9460 2820
rect 9380 2750 9390 2810
rect 9450 2750 9460 2810
rect 9380 2740 9460 2750
rect 8140 2630 8180 2740
rect 8120 2620 8200 2630
rect 8120 2560 8130 2620
rect 8190 2560 8200 2620
rect 8120 2550 8200 2560
rect 6040 2510 6120 2520
rect 6040 2450 6050 2510
rect 6110 2450 6120 2510
rect 6040 2440 6120 2450
rect 6200 2510 6280 2520
rect 6200 2450 6210 2510
rect 6270 2450 6280 2510
rect 6200 2440 6280 2450
rect 6360 2510 6440 2520
rect 6360 2450 6370 2510
rect 6430 2450 6440 2510
rect 6360 2440 6440 2450
rect 6520 2510 6600 2520
rect 6520 2450 6530 2510
rect 6590 2450 6600 2510
rect 6520 2440 6600 2450
rect 6680 2510 6760 2520
rect 6680 2450 6690 2510
rect 6750 2450 6760 2510
rect 6680 2440 6760 2450
rect 6840 2510 6920 2520
rect 6840 2450 6850 2510
rect 6910 2450 6920 2510
rect 6840 2440 6920 2450
rect 7000 2510 7080 2520
rect 7000 2450 7010 2510
rect 7070 2450 7080 2510
rect 7000 2440 7080 2450
rect 7160 2510 7240 2520
rect 7160 2450 7170 2510
rect 7230 2450 7240 2510
rect 7160 2440 7240 2450
rect 7320 2510 7400 2520
rect 7320 2450 7330 2510
rect 7390 2450 7400 2510
rect 7320 2440 7400 2450
rect 7480 2510 7560 2520
rect 7480 2450 7490 2510
rect 7550 2450 7560 2510
rect 7480 2440 7560 2450
rect 7640 2510 7720 2520
rect 7640 2450 7650 2510
rect 7710 2450 7720 2510
rect 7640 2440 7720 2450
rect 7800 2510 7880 2520
rect 7800 2450 7810 2510
rect 7870 2450 7880 2510
rect 7800 2440 7880 2450
rect 7960 2510 8040 2520
rect 7960 2450 7970 2510
rect 8030 2450 8040 2510
rect 7960 2440 8040 2450
rect 8120 2510 8200 2520
rect 8120 2450 8130 2510
rect 8190 2450 8200 2510
rect 8120 2440 8200 2450
rect 8280 2510 8360 2520
rect 8280 2450 8290 2510
rect 8350 2450 8360 2510
rect 8280 2440 8360 2450
rect 8440 2510 8520 2520
rect 8440 2450 8450 2510
rect 8510 2450 8520 2510
rect 8440 2440 8520 2450
rect 8600 2510 8680 2520
rect 8600 2450 8610 2510
rect 8670 2450 8680 2510
rect 8600 2440 8680 2450
rect 8760 2510 8840 2520
rect 8760 2450 8770 2510
rect 8830 2450 8840 2510
rect 8760 2440 8840 2450
rect 8920 2510 9000 2520
rect 8920 2450 8930 2510
rect 8990 2450 9000 2510
rect 8920 2440 9000 2450
rect 9080 2510 9160 2520
rect 9080 2450 9090 2510
rect 9150 2450 9160 2510
rect 9080 2440 9160 2450
rect 9240 2510 9320 2520
rect 9240 2450 9250 2510
rect 9310 2450 9320 2510
rect 9240 2440 9320 2450
rect 9400 2510 9480 2520
rect 9400 2450 9410 2510
rect 9470 2450 9480 2510
rect 9400 2440 9480 2450
rect 9560 2510 9640 2520
rect 9560 2450 9570 2510
rect 9630 2450 9640 2510
rect 9560 2440 9640 2450
rect 9720 2510 9800 2520
rect 9720 2450 9730 2510
rect 9790 2450 9800 2510
rect 9720 2440 9800 2450
rect 9880 2510 9960 2520
rect 9880 2450 9890 2510
rect 9950 2450 9960 2510
rect 9880 2440 9960 2450
rect 10040 2510 10120 2520
rect 10040 2450 10050 2510
rect 10110 2450 10120 2510
rect 35250 2460 35280 3430
rect 36120 3420 36200 3430
rect 36120 3360 36130 3420
rect 36190 3360 36200 3420
rect 36120 3350 36200 3360
rect 35650 3050 35730 3060
rect 35650 2990 35660 3050
rect 35720 2990 35730 3050
rect 35650 2980 35730 2990
rect 36140 2940 36180 3350
rect 37480 3340 37520 3650
rect 37460 3330 37540 3340
rect 37460 3270 37470 3330
rect 37530 3270 37540 3330
rect 37460 3260 37540 3270
rect 38140 3260 38180 3650
rect 38580 3330 38620 3650
rect 39150 3640 39190 4110
rect 39130 3630 39210 3640
rect 39130 3570 39140 3630
rect 39200 3570 39210 3630
rect 39130 3560 39210 3570
rect 39240 3530 39280 4370
rect 39220 3520 39300 3530
rect 39220 3460 39230 3520
rect 39290 3460 39300 3520
rect 39220 3450 39300 3460
rect 39330 3420 39370 4370
rect 39840 4180 39920 4190
rect 39840 4120 39850 4180
rect 39910 4120 39920 4180
rect 39840 4110 39920 4120
rect 39860 4070 39900 4110
rect 39510 4060 39590 4070
rect 39510 4000 39520 4060
rect 39580 4000 39590 4060
rect 39510 3990 39590 4000
rect 39730 4060 39810 4070
rect 39730 4000 39740 4060
rect 39800 4000 39810 4060
rect 39730 3990 39810 4000
rect 39850 4050 39910 4070
rect 39850 4010 39860 4050
rect 39900 4010 39910 4050
rect 39850 3990 39910 4010
rect 39950 4060 40030 4070
rect 39950 4000 39960 4060
rect 40020 4000 40030 4060
rect 39950 3990 40030 4000
rect 40170 4060 40250 4070
rect 40170 4000 40180 4060
rect 40240 4000 40250 4060
rect 40170 3990 40250 4000
rect 39620 3720 39700 3730
rect 39620 3660 39630 3720
rect 39690 3660 39700 3720
rect 39620 3650 39700 3660
rect 39840 3720 39920 3730
rect 39840 3660 39850 3720
rect 39910 3660 39920 3720
rect 39840 3650 39920 3660
rect 40060 3720 40140 3730
rect 40060 3660 40070 3720
rect 40130 3660 40140 3720
rect 40060 3650 40140 3660
rect 39940 3610 40020 3620
rect 39940 3550 39950 3610
rect 40010 3550 40020 3610
rect 39940 3540 40020 3550
rect 39310 3410 39390 3420
rect 39310 3350 39320 3410
rect 39380 3350 39390 3410
rect 39310 3340 39390 3350
rect 38560 3320 38640 3330
rect 38560 3260 38570 3320
rect 38630 3260 38640 3320
rect 38120 3250 38200 3260
rect 38560 3250 38640 3260
rect 38120 3190 38130 3250
rect 38190 3190 38200 3250
rect 38120 3180 38200 3190
rect 36500 3130 36580 3140
rect 36500 3070 36510 3130
rect 36570 3070 36580 3130
rect 36500 3060 36580 3070
rect 36860 3130 36940 3140
rect 36860 3070 36870 3130
rect 36930 3070 36940 3130
rect 36860 3060 36940 3070
rect 37220 3130 37300 3140
rect 37220 3070 37230 3130
rect 37290 3070 37300 3130
rect 37220 3060 37300 3070
rect 37580 3130 37660 3140
rect 37580 3070 37590 3130
rect 37650 3070 37660 3130
rect 37580 3060 37660 3070
rect 37940 3130 38020 3140
rect 37940 3070 37950 3130
rect 38010 3070 38020 3130
rect 37940 3060 38020 3070
rect 38300 3130 38380 3140
rect 38300 3070 38310 3130
rect 38370 3070 38380 3130
rect 38300 3060 38380 3070
rect 38660 3130 38740 3140
rect 38660 3070 38670 3130
rect 38730 3070 38740 3130
rect 38660 3060 38740 3070
rect 39020 3130 39100 3140
rect 39020 3070 39030 3130
rect 39090 3070 39100 3130
rect 39020 3060 39100 3070
rect 39380 3130 39460 3140
rect 39380 3070 39390 3130
rect 39450 3070 39460 3130
rect 39380 3060 39460 3070
rect 39740 3130 39820 3140
rect 39740 3070 39750 3130
rect 39810 3070 39820 3130
rect 39740 3060 39820 3070
rect 35650 2930 35730 2940
rect 35650 2870 35660 2930
rect 35720 2870 35730 2930
rect 35650 2860 35730 2870
rect 36120 2930 36200 2940
rect 36120 2870 36130 2930
rect 36190 2870 36200 2930
rect 36120 2860 36200 2870
rect 35520 2590 35600 2600
rect 35520 2530 35530 2590
rect 35590 2530 35600 2590
rect 35520 2520 35600 2530
rect 35650 2580 35730 2600
rect 35650 2540 35670 2580
rect 35710 2540 35730 2580
rect 35650 2520 35730 2540
rect 35780 2590 35860 2600
rect 35780 2530 35790 2590
rect 35850 2530 35860 2590
rect 35780 2520 35860 2530
rect 10040 2440 10120 2450
rect 5960 2340 6040 2350
rect 5960 2280 5970 2340
rect 6030 2280 6040 2340
rect 5960 2270 6040 2280
rect 10270 2340 10350 2350
rect 10270 2280 10280 2340
rect 10340 2280 10350 2340
rect 10270 2270 10350 2280
rect 34660 2280 34740 2290
rect 34660 2220 34670 2280
rect 34730 2220 34740 2280
rect 34660 2210 34740 2220
rect 34550 2190 34630 2200
rect 34550 2130 34560 2190
rect 34620 2130 34630 2190
rect 34550 2120 34630 2130
rect 6890 2100 6970 2110
rect 6890 2040 6900 2100
rect 6960 2040 6970 2100
rect 6890 2030 6970 2040
rect 8120 2100 8200 2110
rect 8120 2040 8130 2100
rect 8190 2040 8200 2100
rect 8120 2030 8200 2040
rect 9350 2100 9430 2110
rect 9350 2040 9360 2100
rect 9420 2040 9430 2100
rect 9350 2030 9430 2040
rect 6910 1970 6950 2030
rect 8140 1970 8180 2030
rect 9370 1970 9410 2030
rect 6560 1960 6640 1970
rect 6560 1900 6570 1960
rect 6630 1900 6640 1960
rect 6560 1890 6640 1900
rect 6780 1960 6860 1970
rect 6780 1900 6790 1960
rect 6850 1900 6860 1960
rect 6780 1890 6860 1900
rect 6900 1950 6960 1970
rect 6900 1910 6910 1950
rect 6950 1910 6960 1950
rect 6900 1890 6960 1910
rect 7000 1960 7080 1970
rect 7000 1900 7010 1960
rect 7070 1900 7080 1960
rect 7000 1890 7080 1900
rect 7790 1960 7870 1970
rect 7790 1900 7800 1960
rect 7860 1900 7870 1960
rect 7790 1890 7870 1900
rect 8010 1960 8090 1970
rect 8010 1900 8020 1960
rect 8080 1900 8090 1960
rect 8010 1890 8090 1900
rect 8130 1950 8190 1970
rect 8130 1910 8140 1950
rect 8180 1910 8190 1950
rect 8130 1890 8190 1910
rect 8230 1960 8310 1970
rect 8230 1900 8240 1960
rect 8300 1900 8310 1960
rect 8230 1890 8310 1900
rect 8450 1960 8530 1970
rect 8450 1900 8460 1960
rect 8520 1900 8530 1960
rect 8450 1890 8530 1900
rect 9240 1960 9320 1970
rect 9240 1900 9250 1960
rect 9310 1900 9320 1960
rect 9240 1890 9320 1900
rect 9360 1950 9420 1970
rect 9360 1910 9370 1950
rect 9410 1910 9420 1950
rect 9360 1890 9420 1910
rect 9460 1960 9540 1970
rect 9460 1900 9470 1960
rect 9530 1900 9540 1960
rect 9460 1890 9540 1900
rect 9680 1960 9760 1970
rect 9680 1900 9690 1960
rect 9750 1900 9760 1960
rect 9680 1890 9760 1900
rect 7340 1790 7420 1800
rect 7340 1730 7350 1790
rect 7410 1730 7420 1790
rect 7340 1720 7420 1730
rect 7450 1790 7530 1800
rect 7450 1730 7460 1790
rect 7520 1730 7530 1790
rect 7450 1720 7530 1730
rect 8790 1790 8870 1800
rect 8790 1730 8800 1790
rect 8860 1730 8870 1790
rect 8790 1720 8870 1730
rect 8900 1790 8980 1800
rect 8900 1730 8910 1790
rect 8970 1730 8980 1790
rect 8900 1720 8980 1730
rect 10020 1790 10100 1800
rect 10020 1730 10030 1790
rect 10090 1730 10100 1790
rect 10020 1720 10100 1730
rect 6450 1620 6530 1630
rect 6450 1560 6460 1620
rect 6520 1560 6530 1620
rect 6450 1550 6530 1560
rect 6670 1620 6750 1630
rect 6670 1560 6680 1620
rect 6740 1560 6750 1620
rect 6670 1550 6750 1560
rect 6890 1620 6970 1630
rect 6890 1560 6900 1620
rect 6960 1560 6970 1620
rect 6890 1550 6970 1560
rect 7110 1620 7190 1630
rect 7110 1560 7120 1620
rect 7180 1560 7190 1620
rect 7110 1550 7190 1560
rect 7730 1610 7810 1630
rect 7730 1570 7750 1610
rect 7790 1570 7810 1610
rect 7730 1550 7810 1570
rect 7900 1610 7980 1630
rect 7900 1570 7920 1610
rect 7960 1570 7980 1610
rect 7900 1550 7980 1570
rect 8120 1620 8200 1630
rect 8120 1560 8130 1620
rect 8190 1560 8200 1620
rect 8120 1550 8200 1560
rect 8340 1620 8420 1630
rect 8340 1560 8350 1620
rect 8410 1560 8420 1620
rect 8340 1550 8420 1560
rect 8560 1620 8640 1630
rect 8560 1560 8570 1620
rect 8630 1560 8640 1620
rect 8560 1550 8640 1560
rect 9130 1620 9210 1630
rect 9130 1560 9140 1620
rect 9200 1560 9210 1620
rect 9130 1550 9210 1560
rect 9350 1610 9430 1630
rect 9350 1570 9370 1610
rect 9410 1570 9430 1610
rect 9350 1550 9430 1570
rect 9570 1620 9650 1630
rect 9570 1560 9580 1620
rect 9640 1560 9650 1620
rect 9570 1550 9650 1560
rect 9790 1610 9870 1630
rect 9790 1570 9810 1610
rect 9850 1570 9870 1610
rect 9790 1550 9870 1570
rect 5110 1420 5190 1430
rect 5110 1360 5120 1420
rect 5180 1360 5190 1420
rect 5110 1350 5190 1360
rect 6690 1100 6730 1550
rect 7750 1430 7790 1550
rect 7730 1420 7810 1430
rect 7730 1360 7740 1420
rect 7800 1360 7810 1420
rect 7730 1350 7810 1360
rect 7920 1100 7960 1550
rect 8360 1100 8400 1550
rect 9370 1520 9410 1550
rect 9350 1510 9430 1520
rect 9350 1450 9360 1510
rect 9420 1450 9430 1510
rect 9350 1440 9430 1450
rect 9370 1100 9410 1440
rect 9590 1100 9630 1550
rect 9810 1520 9850 1550
rect 9790 1510 9870 1520
rect 9790 1450 9800 1510
rect 9860 1450 9870 1510
rect 9790 1440 9870 1450
rect 34570 -650 34610 2120
rect 34680 1100 34720 2210
rect 34770 2010 34810 2460
rect 34860 2400 34900 2460
rect 34840 2390 34920 2400
rect 34840 2330 34850 2390
rect 34910 2330 34920 2390
rect 34840 2320 34920 2330
rect 34750 2000 34830 2010
rect 34750 1940 34760 2000
rect 34820 1940 34830 2000
rect 34750 1930 34830 1940
rect 34660 1090 34740 1100
rect 34660 1030 34670 1090
rect 34730 1030 34740 1090
rect 34660 1020 34740 1030
rect 34680 430 34720 1020
rect 34860 770 34900 2320
rect 34950 1760 34990 2460
rect 34930 1750 35010 1760
rect 34930 1690 34940 1750
rect 35000 1690 35010 1750
rect 34930 1680 35010 1690
rect 35040 1300 35080 2460
rect 35020 1290 35100 1300
rect 35020 1230 35030 1290
rect 35090 1230 35100 1290
rect 35020 1220 35100 1230
rect 34840 760 34920 770
rect 34840 700 34850 760
rect 34910 700 34920 760
rect 34840 690 34920 700
rect 34660 420 34740 430
rect 34660 360 34670 420
rect 34730 360 34740 420
rect 34660 350 34740 360
rect 34550 -660 34630 -650
rect 34550 -720 34560 -660
rect 34620 -720 34630 -660
rect 34550 -730 34630 -720
rect 35130 -1570 35170 2460
rect 35240 2110 35280 2460
rect 35670 2200 35710 2520
rect 36140 2290 36180 2860
rect 36240 2590 36320 2600
rect 36240 2530 36250 2590
rect 36310 2530 36320 2590
rect 36240 2520 36320 2530
rect 36120 2280 36200 2290
rect 36120 2220 36130 2280
rect 36190 2220 36200 2280
rect 36120 2210 36200 2220
rect 35650 2190 35730 2200
rect 35650 2130 35660 2190
rect 35720 2130 35730 2190
rect 35650 2120 35730 2130
rect 35220 2100 35300 2110
rect 35220 2040 35230 2100
rect 35290 2040 35300 2100
rect 35220 2030 35300 2040
rect 35640 1870 35720 1880
rect 35640 1810 35650 1870
rect 35710 1810 35720 1870
rect 35640 1800 35720 1810
rect 35880 1870 35960 1880
rect 35880 1810 35890 1870
rect 35950 1810 35960 1870
rect 35880 1800 35960 1810
rect 36120 1870 36200 1880
rect 36120 1810 36130 1870
rect 36190 1810 36200 1870
rect 36120 1800 36200 1810
rect 35660 1760 35700 1800
rect 35900 1760 35940 1800
rect 36140 1760 36180 1800
rect 36260 1760 36300 2520
rect 36680 2380 36760 2400
rect 36680 2340 36700 2380
rect 36740 2340 36760 2380
rect 36680 2320 36760 2340
rect 37040 2380 37120 2400
rect 37040 2340 37060 2380
rect 37100 2340 37120 2380
rect 37040 2320 37120 2340
rect 37400 2380 37480 2400
rect 37400 2340 37420 2380
rect 37460 2340 37480 2380
rect 37400 2320 37480 2340
rect 37760 2390 37840 2400
rect 37760 2330 37770 2390
rect 37830 2330 37840 2390
rect 37760 2320 37840 2330
rect 37940 2380 38020 2400
rect 37940 2340 37960 2380
rect 38000 2340 38020 2380
rect 37940 2320 38020 2340
rect 38120 2380 38200 2400
rect 38120 2340 38140 2380
rect 38180 2340 38200 2380
rect 38120 2320 38200 2340
rect 38480 2390 38560 2400
rect 38480 2330 38490 2390
rect 38550 2330 38560 2390
rect 38480 2320 38560 2330
rect 38840 2380 38920 2400
rect 38840 2340 38860 2380
rect 38900 2340 38920 2380
rect 38840 2320 38920 2340
rect 39200 2380 39280 2400
rect 39200 2340 39220 2380
rect 39260 2340 39280 2380
rect 39200 2320 39280 2340
rect 39380 2380 39460 2400
rect 39380 2340 39400 2380
rect 39440 2340 39460 2380
rect 39380 2320 39460 2340
rect 39560 2380 39640 2400
rect 39560 2340 39580 2380
rect 39620 2340 39640 2380
rect 39560 2320 39640 2340
rect 36700 2110 36740 2320
rect 37060 2200 37100 2320
rect 37420 2290 37460 2320
rect 37400 2280 37480 2290
rect 37400 2220 37410 2280
rect 37470 2220 37480 2280
rect 37400 2210 37480 2220
rect 37040 2190 37120 2200
rect 37040 2130 37050 2190
rect 37110 2130 37120 2190
rect 37040 2120 37120 2130
rect 36680 2100 36760 2110
rect 36680 2040 36690 2100
rect 36750 2040 36760 2100
rect 36680 2030 36760 2040
rect 36360 1870 36440 1880
rect 36360 1810 36370 1870
rect 36430 1810 36440 1870
rect 36360 1800 36440 1810
rect 36600 1870 36680 1880
rect 36600 1810 36610 1870
rect 36670 1810 36680 1870
rect 36600 1800 36680 1810
rect 36840 1870 36920 1880
rect 36840 1810 36850 1870
rect 36910 1810 36920 1870
rect 36840 1800 36920 1810
rect 37080 1870 37160 1880
rect 37080 1810 37090 1870
rect 37150 1810 37160 1870
rect 37080 1800 37160 1810
rect 37320 1870 37400 1880
rect 37320 1810 37330 1870
rect 37390 1810 37400 1870
rect 37320 1800 37400 1810
rect 37560 1870 37640 1880
rect 37560 1810 37570 1870
rect 37630 1810 37640 1870
rect 37560 1800 37640 1810
rect 36380 1760 36420 1800
rect 36620 1760 36660 1800
rect 36860 1760 36900 1800
rect 37100 1760 37140 1800
rect 37340 1760 37380 1800
rect 37580 1760 37620 1800
rect 37960 1760 38000 2320
rect 38140 2110 38180 2320
rect 38860 2290 38900 2320
rect 38840 2280 38920 2290
rect 38840 2220 38850 2280
rect 38910 2220 38920 2280
rect 38840 2210 38920 2220
rect 39220 2200 39260 2320
rect 39400 2200 39440 2320
rect 39200 2190 39280 2200
rect 39200 2130 39210 2190
rect 39270 2130 39280 2190
rect 39200 2120 39280 2130
rect 39380 2190 39460 2200
rect 39380 2130 39390 2190
rect 39450 2130 39460 2190
rect 39380 2120 39460 2130
rect 39580 2110 39620 2320
rect 38120 2100 38200 2110
rect 38120 2040 38130 2100
rect 38190 2040 38200 2100
rect 38120 2030 38200 2040
rect 39560 2100 39640 2110
rect 39560 2040 39570 2100
rect 39630 2040 39640 2100
rect 39560 2030 39640 2040
rect 39960 2010 40000 3540
rect 40120 3520 40200 3530
rect 40120 3460 40130 3520
rect 40190 3460 40200 3520
rect 40120 3450 40200 3460
rect 40030 3410 40110 3420
rect 40030 3350 40040 3410
rect 40100 3350 40110 3410
rect 40030 3340 40110 3350
rect 40050 2200 40090 3340
rect 40140 2310 40180 3450
rect 41230 3320 41310 3330
rect 41230 3260 41240 3320
rect 41300 3260 41310 3320
rect 41230 3250 41310 3260
rect 40580 3050 40660 3080
rect 40580 2990 40590 3050
rect 40650 2990 40660 3050
rect 40580 2980 40660 2990
rect 40600 2940 40640 2980
rect 40580 2930 40660 2940
rect 40580 2870 40590 2930
rect 40650 2870 40660 2930
rect 40580 2860 40660 2870
rect 40450 2590 40530 2600
rect 40450 2530 40460 2590
rect 40520 2530 40530 2590
rect 40450 2520 40530 2530
rect 40580 2580 40660 2600
rect 40580 2540 40600 2580
rect 40640 2540 40660 2580
rect 40580 2520 40660 2540
rect 40710 2590 40790 2600
rect 40710 2530 40720 2590
rect 40780 2530 40790 2590
rect 40710 2520 40790 2530
rect 40120 2300 40200 2310
rect 40120 2240 40130 2300
rect 40190 2240 40200 2300
rect 40120 2230 40200 2240
rect 40030 2190 40110 2200
rect 40030 2130 40040 2190
rect 40100 2130 40110 2190
rect 40030 2120 40110 2130
rect 40600 2010 40640 2520
rect 41050 2300 41130 2310
rect 41050 2240 41060 2300
rect 41120 2240 41130 2300
rect 41050 2230 41130 2240
rect 38560 2000 38640 2010
rect 38560 1940 38570 2000
rect 38630 1940 38640 2000
rect 38560 1930 38640 1940
rect 39940 2000 40020 2010
rect 39940 1940 39950 2000
rect 40010 1940 40020 2000
rect 39940 1930 40020 1940
rect 40580 2000 40660 2010
rect 40580 1940 40590 2000
rect 40650 1940 40660 2000
rect 40580 1930 40660 1940
rect 38580 1760 38620 1930
rect 38680 1870 38760 1880
rect 38680 1810 38690 1870
rect 38750 1810 38760 1870
rect 38680 1800 38760 1810
rect 38920 1870 39000 1880
rect 38920 1810 38930 1870
rect 38990 1810 39000 1870
rect 38920 1800 39000 1810
rect 39160 1870 39240 1880
rect 39160 1810 39170 1870
rect 39230 1810 39240 1870
rect 39160 1800 39240 1810
rect 39400 1870 39480 1880
rect 39400 1810 39410 1870
rect 39470 1810 39480 1870
rect 39400 1800 39480 1810
rect 39640 1870 39720 1880
rect 39640 1810 39650 1870
rect 39710 1810 39720 1870
rect 39640 1800 39720 1810
rect 39880 1870 39960 1880
rect 39880 1810 39890 1870
rect 39950 1810 39960 1870
rect 39880 1800 39960 1810
rect 40120 1870 40200 1880
rect 40120 1810 40130 1870
rect 40190 1810 40200 1870
rect 40120 1800 40200 1810
rect 40360 1870 40440 1880
rect 40360 1810 40370 1870
rect 40430 1810 40440 1870
rect 40360 1800 40440 1810
rect 40600 1870 40680 1880
rect 40600 1810 40610 1870
rect 40670 1810 40680 1870
rect 40600 1800 40680 1810
rect 38700 1760 38740 1800
rect 38940 1760 38980 1800
rect 39180 1760 39220 1800
rect 39420 1760 39460 1800
rect 39660 1760 39700 1800
rect 39900 1760 39940 1800
rect 40140 1760 40180 1800
rect 40380 1760 40420 1800
rect 40620 1760 40660 1800
rect 35520 1750 35600 1760
rect 35520 1690 35530 1750
rect 35590 1690 35600 1750
rect 35520 1680 35600 1690
rect 35650 1740 35710 1760
rect 35650 1700 35660 1740
rect 35700 1700 35710 1740
rect 35650 1680 35710 1700
rect 35890 1740 35950 1760
rect 35890 1700 35900 1740
rect 35940 1700 35950 1740
rect 35890 1680 35950 1700
rect 36130 1740 36190 1760
rect 36130 1700 36140 1740
rect 36180 1700 36190 1740
rect 36130 1680 36190 1700
rect 36240 1750 36320 1760
rect 36240 1690 36250 1750
rect 36310 1690 36320 1750
rect 36240 1680 36320 1690
rect 36370 1740 36430 1760
rect 36370 1700 36380 1740
rect 36420 1700 36430 1740
rect 36370 1680 36430 1700
rect 36610 1740 36670 1760
rect 36610 1700 36620 1740
rect 36660 1700 36670 1740
rect 36610 1680 36670 1700
rect 36850 1740 36910 1760
rect 36850 1700 36860 1740
rect 36900 1700 36910 1740
rect 36850 1680 36910 1700
rect 36960 1750 37040 1760
rect 36960 1690 36970 1750
rect 37030 1690 37040 1750
rect 36960 1680 37040 1690
rect 37090 1740 37150 1760
rect 37090 1700 37100 1740
rect 37140 1700 37150 1740
rect 37090 1680 37150 1700
rect 37330 1740 37390 1760
rect 37330 1700 37340 1740
rect 37380 1700 37390 1740
rect 37330 1680 37390 1700
rect 37570 1740 37630 1760
rect 37570 1700 37580 1740
rect 37620 1700 37630 1740
rect 37570 1680 37630 1700
rect 37680 1750 37760 1760
rect 37680 1690 37690 1750
rect 37750 1690 37760 1750
rect 37680 1680 37760 1690
rect 37940 1750 38020 1760
rect 37940 1690 37950 1750
rect 38010 1690 38020 1750
rect 37940 1680 38020 1690
rect 38300 1750 38380 1760
rect 38300 1690 38310 1750
rect 38370 1690 38380 1750
rect 38300 1680 38380 1690
rect 38560 1750 38640 1760
rect 38560 1690 38570 1750
rect 38630 1690 38640 1750
rect 38560 1680 38640 1690
rect 38690 1740 38750 1760
rect 38690 1700 38700 1740
rect 38740 1700 38750 1740
rect 38690 1680 38750 1700
rect 38930 1740 38990 1760
rect 38930 1700 38940 1740
rect 38980 1700 38990 1740
rect 38930 1680 38990 1700
rect 39170 1740 39230 1760
rect 39170 1700 39180 1740
rect 39220 1700 39230 1740
rect 39170 1680 39230 1700
rect 39280 1750 39360 1760
rect 39280 1690 39290 1750
rect 39350 1690 39360 1750
rect 39280 1680 39360 1690
rect 39410 1740 39470 1760
rect 39410 1700 39420 1740
rect 39460 1700 39470 1740
rect 39410 1680 39470 1700
rect 39650 1740 39710 1760
rect 39650 1700 39660 1740
rect 39700 1700 39710 1740
rect 39650 1680 39710 1700
rect 39890 1740 39950 1760
rect 39890 1700 39900 1740
rect 39940 1700 39950 1740
rect 39890 1680 39950 1700
rect 40000 1750 40080 1760
rect 40000 1690 40010 1750
rect 40070 1690 40080 1750
rect 40000 1680 40080 1690
rect 40130 1740 40190 1760
rect 40130 1700 40140 1740
rect 40180 1700 40190 1740
rect 40130 1680 40190 1700
rect 40370 1740 40430 1760
rect 40370 1700 40380 1740
rect 40420 1700 40430 1740
rect 40370 1680 40430 1700
rect 40610 1740 40670 1760
rect 40610 1700 40620 1740
rect 40660 1700 40670 1740
rect 40610 1680 40670 1700
rect 40720 1750 40800 1760
rect 40720 1690 40730 1750
rect 40790 1690 40800 1750
rect 40720 1680 40800 1690
rect 35580 1400 35660 1420
rect 35580 1360 35600 1400
rect 35640 1360 35660 1400
rect 35580 1340 35660 1360
rect 35760 1410 35840 1420
rect 35760 1350 35770 1410
rect 35830 1350 35840 1410
rect 35760 1340 35840 1350
rect 36000 1400 36080 1420
rect 36000 1360 36020 1400
rect 36060 1360 36080 1400
rect 36000 1340 36080 1360
rect 36240 1400 36320 1420
rect 36240 1360 36260 1400
rect 36300 1360 36320 1400
rect 36240 1340 36320 1360
rect 36480 1410 36560 1420
rect 36480 1350 36490 1410
rect 36550 1350 36560 1410
rect 36480 1340 36560 1350
rect 36720 1400 36800 1420
rect 36720 1360 36740 1400
rect 36780 1360 36800 1400
rect 36720 1340 36800 1360
rect 36960 1400 37040 1420
rect 36960 1360 36980 1400
rect 37020 1360 37040 1400
rect 36960 1340 37040 1360
rect 37200 1410 37280 1420
rect 37200 1350 37210 1410
rect 37270 1350 37280 1410
rect 37200 1340 37280 1350
rect 37440 1400 37520 1420
rect 37440 1360 37460 1400
rect 37500 1360 37520 1400
rect 37440 1340 37520 1360
rect 37630 1400 37690 1420
rect 37630 1360 37640 1400
rect 37680 1360 37690 1400
rect 37630 1340 37690 1360
rect 35600 1300 35640 1340
rect 36020 1300 36060 1340
rect 36260 1300 36300 1340
rect 35580 1290 35660 1300
rect 35580 1230 35590 1290
rect 35650 1230 35660 1290
rect 35580 1220 35660 1230
rect 36000 1290 36080 1300
rect 36000 1230 36010 1290
rect 36070 1230 36080 1290
rect 36000 1220 36080 1230
rect 36240 1290 36320 1300
rect 36240 1230 36250 1290
rect 36310 1230 36320 1290
rect 36240 1220 36320 1230
rect 36520 1130 36560 1340
rect 36740 1300 36780 1340
rect 36980 1300 37020 1340
rect 37460 1300 37500 1340
rect 37640 1300 37680 1340
rect 36720 1290 36800 1300
rect 36720 1230 36730 1290
rect 36790 1230 36800 1290
rect 36720 1220 36800 1230
rect 36960 1290 37040 1300
rect 36960 1230 36970 1290
rect 37030 1230 37040 1290
rect 36960 1220 37040 1230
rect 37440 1290 37520 1300
rect 37440 1230 37450 1290
rect 37510 1230 37520 1290
rect 37440 1220 37520 1230
rect 37620 1290 37700 1300
rect 37620 1230 37630 1290
rect 37690 1230 37700 1290
rect 37620 1220 37700 1230
rect 36500 1120 36580 1130
rect 36380 1090 36460 1100
rect 36380 1030 36390 1090
rect 36450 1030 36460 1090
rect 36500 1060 36510 1120
rect 36570 1060 36580 1120
rect 36500 1050 36580 1060
rect 36380 1020 36460 1030
rect 36520 1010 36560 1050
rect 36740 1010 36780 1220
rect 36980 1120 37060 1130
rect 36980 1060 36990 1120
rect 37050 1060 37060 1120
rect 36980 1050 37060 1060
rect 37460 1120 37540 1130
rect 37460 1060 37470 1120
rect 37530 1060 37540 1120
rect 37460 1050 37540 1060
rect 37000 1010 37040 1050
rect 37480 1010 37520 1050
rect 36260 1000 36340 1010
rect 36260 940 36270 1000
rect 36330 940 36340 1000
rect 36260 930 36340 940
rect 36510 990 36570 1010
rect 36510 950 36520 990
rect 36560 950 36570 990
rect 36510 930 36570 950
rect 36740 1000 36820 1010
rect 36740 940 36750 1000
rect 36810 940 36820 1000
rect 36740 930 36820 940
rect 36990 990 37050 1010
rect 36990 950 37000 990
rect 37040 950 37050 990
rect 36990 930 37050 950
rect 37220 1000 37300 1010
rect 37220 940 37230 1000
rect 37290 940 37300 1000
rect 37220 930 37300 940
rect 37470 990 37530 1010
rect 37470 950 37480 990
rect 37520 950 37530 990
rect 37470 930 37530 950
rect 37580 880 37660 890
rect 37580 820 37590 880
rect 37650 820 37660 880
rect 37580 810 37660 820
rect 36260 760 36340 770
rect 36260 700 36270 760
rect 36330 700 36340 760
rect 36260 690 36340 700
rect 36390 750 36450 770
rect 36390 710 36400 750
rect 36440 710 36450 750
rect 36390 690 36450 710
rect 36630 750 36690 770
rect 36630 710 36640 750
rect 36680 710 36690 750
rect 36630 690 36690 710
rect 36870 750 36930 770
rect 36870 710 36880 750
rect 36920 710 36930 750
rect 36870 690 36930 710
rect 37110 750 37170 770
rect 37110 710 37120 750
rect 37160 710 37170 750
rect 37110 690 37170 710
rect 37350 750 37410 770
rect 37350 710 37360 750
rect 37400 710 37410 750
rect 37350 690 37410 710
rect 36400 650 36440 690
rect 36640 650 36680 690
rect 36880 650 36920 690
rect 37120 650 37160 690
rect 37360 650 37400 690
rect 35780 640 35860 650
rect 35780 580 35790 640
rect 35850 580 35860 640
rect 35780 570 35860 580
rect 36380 640 36460 650
rect 36380 580 36390 640
rect 36450 580 36460 640
rect 36380 570 36460 580
rect 36620 640 36700 650
rect 36620 580 36630 640
rect 36690 580 36700 640
rect 36620 570 36700 580
rect 36860 640 36940 650
rect 36860 580 36870 640
rect 36930 580 36940 640
rect 36860 570 36940 580
rect 37100 640 37180 650
rect 37100 580 37110 640
rect 37170 580 37180 640
rect 37100 570 37180 580
rect 37340 640 37420 650
rect 37340 580 37350 640
rect 37410 580 37420 640
rect 37340 570 37420 580
rect 35800 420 35840 570
rect 35960 440 36040 450
rect 35780 400 35860 420
rect 35780 360 35800 400
rect 35840 360 35860 400
rect 35960 380 35970 440
rect 36030 380 36040 440
rect 35960 370 36040 380
rect 36200 440 36280 450
rect 36200 380 36210 440
rect 36270 380 36280 440
rect 36200 370 36280 380
rect 36440 440 36520 450
rect 36440 380 36450 440
rect 36510 380 36520 440
rect 36440 370 36520 380
rect 36680 440 36760 450
rect 36680 380 36690 440
rect 36750 380 36760 440
rect 36680 370 36760 380
rect 37160 440 37240 450
rect 37160 380 37170 440
rect 37230 380 37240 440
rect 37160 370 37240 380
rect 37400 440 37480 450
rect 37400 380 37410 440
rect 37470 380 37480 440
rect 37400 370 37480 380
rect 37640 440 37720 450
rect 37640 380 37650 440
rect 37710 380 37720 440
rect 37960 420 38000 1680
rect 38120 880 38200 890
rect 38120 820 38130 880
rect 38190 820 38200 880
rect 38120 810 38200 820
rect 37640 370 37720 380
rect 37940 400 38020 420
rect 35780 340 35860 360
rect 37940 360 37960 400
rect 38000 360 38020 400
rect 37940 340 38020 360
rect 38140 -180 38180 810
rect 38320 420 38360 1680
rect 38630 1400 38690 1420
rect 38630 1360 38640 1400
rect 38680 1360 38690 1400
rect 38630 1340 38690 1360
rect 38800 1400 38880 1420
rect 38800 1360 38820 1400
rect 38860 1360 38880 1400
rect 38800 1340 38880 1360
rect 39040 1410 39120 1420
rect 39040 1350 39050 1410
rect 39110 1350 39120 1410
rect 39040 1340 39120 1350
rect 39280 1400 39360 1420
rect 39280 1360 39300 1400
rect 39340 1360 39360 1400
rect 39280 1340 39360 1360
rect 39520 1400 39600 1420
rect 39520 1360 39540 1400
rect 39580 1360 39600 1400
rect 39520 1340 39600 1360
rect 39760 1410 39840 1420
rect 39760 1350 39770 1410
rect 39830 1350 39840 1410
rect 39760 1340 39840 1350
rect 40000 1400 40080 1420
rect 40000 1360 40020 1400
rect 40060 1360 40080 1400
rect 40000 1340 40080 1360
rect 40240 1400 40320 1420
rect 40240 1360 40260 1400
rect 40300 1360 40320 1400
rect 40240 1340 40320 1360
rect 40480 1410 40560 1420
rect 40480 1350 40490 1410
rect 40550 1350 40560 1410
rect 40480 1340 40560 1350
rect 40660 1400 40740 1420
rect 40660 1360 40680 1400
rect 40720 1360 40740 1400
rect 40660 1340 40740 1360
rect 38640 1300 38680 1340
rect 38820 1300 38860 1340
rect 39300 1300 39340 1340
rect 39540 1300 39580 1340
rect 38620 1290 38700 1300
rect 38620 1230 38630 1290
rect 38690 1230 38700 1290
rect 38620 1220 38700 1230
rect 38800 1290 38880 1300
rect 38800 1230 38810 1290
rect 38870 1230 38880 1290
rect 38800 1220 38880 1230
rect 39280 1290 39360 1300
rect 39280 1230 39290 1290
rect 39350 1230 39360 1290
rect 39280 1220 39360 1230
rect 39520 1290 39600 1300
rect 39520 1230 39530 1290
rect 39590 1230 39600 1290
rect 39520 1220 39600 1230
rect 38780 1120 38860 1130
rect 38780 1060 38790 1120
rect 38850 1060 38860 1120
rect 38780 1050 38860 1060
rect 39260 1120 39340 1130
rect 39260 1060 39270 1120
rect 39330 1060 39340 1120
rect 39260 1050 39340 1060
rect 38800 1010 38840 1050
rect 39280 1010 39320 1050
rect 39520 1010 39560 1220
rect 39760 1130 39800 1340
rect 40020 1300 40060 1340
rect 40260 1300 40300 1340
rect 40680 1300 40720 1340
rect 41070 1300 41110 2230
rect 41140 2100 41220 2110
rect 41140 2040 41150 2100
rect 41210 2040 41220 2100
rect 41140 2030 41220 2040
rect 40000 1290 40080 1300
rect 40000 1230 40010 1290
rect 40070 1230 40080 1290
rect 40000 1220 40080 1230
rect 40240 1290 40320 1300
rect 40240 1230 40250 1290
rect 40310 1230 40320 1290
rect 40240 1220 40320 1230
rect 40660 1290 40740 1300
rect 40660 1230 40670 1290
rect 40730 1230 40740 1290
rect 40660 1220 40740 1230
rect 41050 1290 41130 1300
rect 41050 1230 41060 1290
rect 41120 1230 41130 1290
rect 41050 1220 41130 1230
rect 39740 1120 39820 1130
rect 39740 1060 39750 1120
rect 39810 1060 39820 1120
rect 41160 1100 41200 2030
rect 39740 1050 39820 1060
rect 39860 1090 39940 1100
rect 39760 1010 39800 1050
rect 39860 1030 39870 1090
rect 39930 1030 39940 1090
rect 39860 1020 39940 1030
rect 41140 1090 41220 1100
rect 41140 1030 41150 1090
rect 41210 1030 41220 1090
rect 41140 1020 41220 1030
rect 38790 990 38850 1010
rect 38790 950 38800 990
rect 38840 950 38850 990
rect 38790 930 38850 950
rect 39020 1000 39100 1010
rect 39020 940 39030 1000
rect 39090 940 39100 1000
rect 39020 930 39100 940
rect 39270 990 39330 1010
rect 39270 950 39280 990
rect 39320 950 39330 990
rect 39270 930 39330 950
rect 39500 1000 39580 1010
rect 39500 940 39510 1000
rect 39570 940 39580 1000
rect 39500 930 39580 940
rect 39750 990 39810 1010
rect 39750 950 39760 990
rect 39800 950 39810 990
rect 39750 930 39810 950
rect 39980 1000 40060 1010
rect 39980 940 39990 1000
rect 40050 940 40060 1000
rect 39980 930 40060 940
rect 38660 880 38740 890
rect 38660 820 38670 880
rect 38730 820 38740 880
rect 38660 810 38740 820
rect 41250 770 41290 3250
rect 38910 750 38970 770
rect 38910 710 38920 750
rect 38960 710 38970 750
rect 38910 690 38970 710
rect 39150 750 39210 770
rect 39150 710 39160 750
rect 39200 710 39210 750
rect 39150 690 39210 710
rect 39390 750 39450 770
rect 39390 710 39400 750
rect 39440 710 39450 750
rect 39390 690 39450 710
rect 39630 750 39690 770
rect 39630 710 39640 750
rect 39680 710 39690 750
rect 39630 690 39690 710
rect 39870 750 39930 770
rect 39870 710 39880 750
rect 39920 710 39930 750
rect 39870 690 39930 710
rect 39980 760 40060 770
rect 39980 700 39990 760
rect 40050 700 40060 760
rect 39980 690 40060 700
rect 41230 760 41310 770
rect 41230 700 41240 760
rect 41300 700 41310 760
rect 41230 690 41310 700
rect 38920 650 38960 690
rect 39160 650 39200 690
rect 39400 650 39440 690
rect 39640 650 39680 690
rect 39880 650 39920 690
rect 38900 640 38980 650
rect 38900 580 38910 640
rect 38970 580 38980 640
rect 38900 570 38980 580
rect 39140 640 39220 650
rect 39140 580 39150 640
rect 39210 580 39220 640
rect 39140 570 39220 580
rect 39380 640 39460 650
rect 39380 580 39390 640
rect 39450 580 39460 640
rect 39380 570 39460 580
rect 39620 640 39700 650
rect 39620 580 39630 640
rect 39690 580 39700 640
rect 39620 570 39700 580
rect 39860 640 39940 650
rect 39860 580 39870 640
rect 39930 580 39940 640
rect 39860 570 39940 580
rect 40460 640 40540 650
rect 40460 580 40470 640
rect 40530 580 40540 640
rect 40460 570 40540 580
rect 38600 440 38680 450
rect 38300 400 38380 420
rect 38300 360 38320 400
rect 38360 360 38380 400
rect 38600 380 38610 440
rect 38670 380 38680 440
rect 38600 370 38680 380
rect 38840 440 38920 450
rect 38840 380 38850 440
rect 38910 380 38920 440
rect 38840 370 38920 380
rect 39080 440 39160 450
rect 39080 380 39090 440
rect 39150 380 39160 440
rect 39080 370 39160 380
rect 39560 440 39640 450
rect 39560 380 39570 440
rect 39630 380 39640 440
rect 39560 370 39640 380
rect 39800 440 39880 450
rect 39800 380 39810 440
rect 39870 380 39880 440
rect 39800 370 39880 380
rect 40040 440 40120 450
rect 40040 380 40050 440
rect 40110 380 40120 440
rect 40040 370 40120 380
rect 40280 440 40360 450
rect 40280 380 40290 440
rect 40350 380 40360 440
rect 40480 420 40520 570
rect 40280 370 40360 380
rect 40460 400 40540 420
rect 38300 340 38380 360
rect 40460 360 40480 400
rect 40520 360 40540 400
rect 40460 340 40540 360
rect 36860 -190 36940 -180
rect 36860 -250 36870 -190
rect 36930 -250 36940 -190
rect 36860 -260 36940 -250
rect 38120 -190 38200 -180
rect 38120 -250 38130 -190
rect 38190 -250 38200 -190
rect 38120 -260 38200 -250
rect 39380 -190 39460 -180
rect 39380 -250 39390 -190
rect 39450 -250 39460 -190
rect 39380 -260 39460 -250
rect 38140 -370 38180 -260
rect 38120 -380 38200 -370
rect 38120 -440 38130 -380
rect 38190 -440 38200 -380
rect 38120 -450 38200 -440
rect 36040 -490 36120 -480
rect 36040 -550 36050 -490
rect 36110 -550 36120 -490
rect 36040 -560 36120 -550
rect 36200 -490 36280 -480
rect 36200 -550 36210 -490
rect 36270 -550 36280 -490
rect 36200 -560 36280 -550
rect 36360 -490 36440 -480
rect 36360 -550 36370 -490
rect 36430 -550 36440 -490
rect 36360 -560 36440 -550
rect 36520 -490 36600 -480
rect 36520 -550 36530 -490
rect 36590 -550 36600 -490
rect 36520 -560 36600 -550
rect 36680 -490 36760 -480
rect 36680 -550 36690 -490
rect 36750 -550 36760 -490
rect 36680 -560 36760 -550
rect 36840 -490 36920 -480
rect 36840 -550 36850 -490
rect 36910 -550 36920 -490
rect 36840 -560 36920 -550
rect 37000 -490 37080 -480
rect 37000 -550 37010 -490
rect 37070 -550 37080 -490
rect 37000 -560 37080 -550
rect 37160 -490 37240 -480
rect 37160 -550 37170 -490
rect 37230 -550 37240 -490
rect 37160 -560 37240 -550
rect 37320 -490 37400 -480
rect 37320 -550 37330 -490
rect 37390 -550 37400 -490
rect 37320 -560 37400 -550
rect 37480 -490 37560 -480
rect 37480 -550 37490 -490
rect 37550 -550 37560 -490
rect 37480 -560 37560 -550
rect 37640 -490 37720 -480
rect 37640 -550 37650 -490
rect 37710 -550 37720 -490
rect 37640 -560 37720 -550
rect 37800 -490 37880 -480
rect 37800 -550 37810 -490
rect 37870 -550 37880 -490
rect 37800 -560 37880 -550
rect 37960 -490 38040 -480
rect 37960 -550 37970 -490
rect 38030 -550 38040 -490
rect 37960 -560 38040 -550
rect 38120 -490 38200 -480
rect 38120 -550 38130 -490
rect 38190 -550 38200 -490
rect 38120 -560 38200 -550
rect 38280 -490 38360 -480
rect 38280 -550 38290 -490
rect 38350 -550 38360 -490
rect 38280 -560 38360 -550
rect 38440 -490 38520 -480
rect 38440 -550 38450 -490
rect 38510 -550 38520 -490
rect 38440 -560 38520 -550
rect 38600 -490 38680 -480
rect 38600 -550 38610 -490
rect 38670 -550 38680 -490
rect 38600 -560 38680 -550
rect 38760 -490 38840 -480
rect 38760 -550 38770 -490
rect 38830 -550 38840 -490
rect 38760 -560 38840 -550
rect 38920 -490 39000 -480
rect 38920 -550 38930 -490
rect 38990 -550 39000 -490
rect 38920 -560 39000 -550
rect 39080 -490 39160 -480
rect 39080 -550 39090 -490
rect 39150 -550 39160 -490
rect 39080 -560 39160 -550
rect 39240 -490 39320 -480
rect 39240 -550 39250 -490
rect 39310 -550 39320 -490
rect 39240 -560 39320 -550
rect 39400 -490 39480 -480
rect 39400 -550 39410 -490
rect 39470 -550 39480 -490
rect 39400 -560 39480 -550
rect 39560 -490 39640 -480
rect 39560 -550 39570 -490
rect 39630 -550 39640 -490
rect 39560 -560 39640 -550
rect 39720 -490 39800 -480
rect 39720 -550 39730 -490
rect 39790 -550 39800 -490
rect 39720 -560 39800 -550
rect 39880 -490 39960 -480
rect 39880 -550 39890 -490
rect 39950 -550 39960 -490
rect 39880 -560 39960 -550
rect 40040 -490 40120 -480
rect 40040 -550 40050 -490
rect 40110 -550 40120 -490
rect 40040 -560 40120 -550
rect 35960 -660 36040 -650
rect 35960 -720 35970 -660
rect 36030 -720 36040 -660
rect 35960 -730 36040 -720
rect 40270 -660 40350 -650
rect 40270 -720 40280 -660
rect 40340 -720 40350 -660
rect 40270 -730 40350 -720
rect 36890 -900 36970 -890
rect 36890 -960 36900 -900
rect 36960 -960 36970 -900
rect 36890 -970 36970 -960
rect 38120 -900 38200 -890
rect 38120 -960 38130 -900
rect 38190 -960 38200 -900
rect 38120 -970 38200 -960
rect 39350 -900 39430 -890
rect 39350 -960 39360 -900
rect 39420 -960 39430 -900
rect 39350 -970 39430 -960
rect 36910 -1030 36950 -970
rect 38140 -1030 38180 -970
rect 39370 -1030 39410 -970
rect 36560 -1040 36640 -1030
rect 36560 -1100 36570 -1040
rect 36630 -1100 36640 -1040
rect 36560 -1110 36640 -1100
rect 36780 -1040 36860 -1030
rect 36780 -1100 36790 -1040
rect 36850 -1100 36860 -1040
rect 36780 -1110 36860 -1100
rect 36900 -1050 36960 -1030
rect 36900 -1090 36910 -1050
rect 36950 -1090 36960 -1050
rect 36900 -1110 36960 -1090
rect 37000 -1040 37080 -1030
rect 37000 -1100 37010 -1040
rect 37070 -1100 37080 -1040
rect 37000 -1110 37080 -1100
rect 37790 -1040 37870 -1030
rect 37790 -1100 37800 -1040
rect 37860 -1100 37870 -1040
rect 37790 -1110 37870 -1100
rect 38010 -1040 38090 -1030
rect 38010 -1100 38020 -1040
rect 38080 -1100 38090 -1040
rect 38010 -1110 38090 -1100
rect 38130 -1050 38190 -1030
rect 38130 -1090 38140 -1050
rect 38180 -1090 38190 -1050
rect 38130 -1110 38190 -1090
rect 38230 -1040 38310 -1030
rect 38230 -1100 38240 -1040
rect 38300 -1100 38310 -1040
rect 38230 -1110 38310 -1100
rect 38450 -1040 38530 -1030
rect 38450 -1100 38460 -1040
rect 38520 -1100 38530 -1040
rect 38450 -1110 38530 -1100
rect 39240 -1040 39320 -1030
rect 39240 -1100 39250 -1040
rect 39310 -1100 39320 -1040
rect 39240 -1110 39320 -1100
rect 39360 -1050 39420 -1030
rect 39360 -1090 39370 -1050
rect 39410 -1090 39420 -1050
rect 39360 -1110 39420 -1090
rect 39460 -1040 39540 -1030
rect 39460 -1100 39470 -1040
rect 39530 -1100 39540 -1040
rect 39460 -1110 39540 -1100
rect 39680 -1040 39760 -1030
rect 39680 -1100 39690 -1040
rect 39750 -1100 39760 -1040
rect 39680 -1110 39760 -1100
rect 37340 -1210 37420 -1200
rect 37340 -1270 37350 -1210
rect 37410 -1270 37420 -1210
rect 37340 -1280 37420 -1270
rect 37450 -1210 37530 -1200
rect 37450 -1270 37460 -1210
rect 37520 -1270 37530 -1210
rect 37450 -1280 37530 -1270
rect 38790 -1210 38870 -1200
rect 38790 -1270 38800 -1210
rect 38860 -1270 38870 -1210
rect 38790 -1280 38870 -1270
rect 38900 -1210 38980 -1200
rect 38900 -1270 38910 -1210
rect 38970 -1270 38980 -1210
rect 38900 -1280 38980 -1270
rect 40020 -1210 40100 -1200
rect 40020 -1270 40030 -1210
rect 40090 -1270 40100 -1210
rect 40020 -1280 40100 -1270
rect 36450 -1380 36530 -1370
rect 36450 -1440 36460 -1380
rect 36520 -1440 36530 -1380
rect 36450 -1450 36530 -1440
rect 36670 -1380 36750 -1370
rect 36670 -1440 36680 -1380
rect 36740 -1440 36750 -1380
rect 36670 -1450 36750 -1440
rect 36890 -1380 36970 -1370
rect 36890 -1440 36900 -1380
rect 36960 -1440 36970 -1380
rect 36890 -1450 36970 -1440
rect 37110 -1380 37190 -1370
rect 37110 -1440 37120 -1380
rect 37180 -1440 37190 -1380
rect 37110 -1450 37190 -1440
rect 37730 -1390 37810 -1370
rect 37730 -1430 37750 -1390
rect 37790 -1430 37810 -1390
rect 37730 -1450 37810 -1430
rect 37900 -1390 37980 -1370
rect 37900 -1430 37920 -1390
rect 37960 -1430 37980 -1390
rect 37900 -1450 37980 -1430
rect 38120 -1380 38200 -1370
rect 38120 -1440 38130 -1380
rect 38190 -1440 38200 -1380
rect 38120 -1450 38200 -1440
rect 38340 -1380 38420 -1370
rect 38340 -1440 38350 -1380
rect 38410 -1440 38420 -1380
rect 38340 -1450 38420 -1440
rect 38560 -1380 38640 -1370
rect 38560 -1440 38570 -1380
rect 38630 -1440 38640 -1380
rect 38560 -1450 38640 -1440
rect 39130 -1380 39210 -1370
rect 39130 -1440 39140 -1380
rect 39200 -1440 39210 -1380
rect 39130 -1450 39210 -1440
rect 39350 -1390 39430 -1370
rect 39350 -1430 39370 -1390
rect 39410 -1430 39430 -1390
rect 39350 -1450 39430 -1430
rect 39570 -1380 39650 -1370
rect 39570 -1440 39580 -1380
rect 39640 -1440 39650 -1380
rect 39570 -1450 39650 -1440
rect 39790 -1390 39870 -1370
rect 39790 -1430 39810 -1390
rect 39850 -1430 39870 -1390
rect 39790 -1450 39870 -1430
rect 35110 -1580 35190 -1570
rect 35110 -1640 35120 -1580
rect 35180 -1640 35190 -1580
rect 35110 -1650 35190 -1640
rect 36690 -1900 36730 -1450
rect 37750 -1570 37790 -1450
rect 37730 -1580 37810 -1570
rect 37730 -1640 37740 -1580
rect 37800 -1640 37810 -1580
rect 37730 -1650 37810 -1640
rect 37920 -1900 37960 -1450
rect 38360 -1900 38400 -1450
rect 39370 -1480 39410 -1450
rect 39350 -1490 39430 -1480
rect 39350 -1550 39360 -1490
rect 39420 -1550 39430 -1490
rect 39350 -1560 39430 -1550
rect 39370 -1900 39410 -1560
rect 39590 -1900 39630 -1450
rect 39810 -1480 39850 -1450
rect 39790 -1490 39870 -1480
rect 39790 -1550 39800 -1490
rect 39860 -1550 39870 -1490
rect 39790 -1560 39870 -1550
rect 46510 -2620 46590 -2610
rect 43900 -3880 43940 -2620
rect 43880 -3890 43960 -3880
rect 43880 -3950 43890 -3890
rect 43950 -3950 43960 -3890
rect 43880 -3960 43960 -3950
rect 43990 -4290 44030 -2620
rect 46510 -2680 46520 -2620
rect 46580 -2680 46590 -2620
rect 46510 -2690 46590 -2680
rect 44140 -2720 44220 -2710
rect 44140 -2780 44150 -2720
rect 44210 -2780 44220 -2720
rect 44140 -2790 44220 -2780
rect 44150 -2820 44200 -2790
rect 44132 -2890 44142 -2820
rect 44212 -2890 44222 -2820
rect 44132 -3010 44142 -2940
rect 44212 -3010 44222 -2940
rect 46530 -3240 46570 -2690
rect 46720 -3090 46760 -2620
rect 46702 -3160 46712 -3090
rect 46782 -3160 46792 -3090
rect 46722 -3210 46762 -3160
rect 44140 -3250 44220 -3240
rect 44140 -3310 44150 -3250
rect 44210 -3310 44220 -3250
rect 44140 -3320 44220 -3310
rect 46510 -3250 46590 -3240
rect 46510 -3310 46520 -3250
rect 46580 -3310 46590 -3250
rect 46702 -3280 46712 -3210
rect 46782 -3280 46792 -3210
rect 46510 -3320 46590 -3310
rect 44150 -3350 44200 -3320
rect 44132 -3420 44142 -3350
rect 44212 -3420 44222 -3350
rect 46370 -3420 46450 -3410
rect 44132 -3540 44142 -3470
rect 44212 -3540 44222 -3470
rect 46370 -3480 46380 -3420
rect 46440 -3480 46450 -3420
rect 46370 -3490 46450 -3480
rect 46580 -3420 46660 -3410
rect 46580 -3480 46590 -3420
rect 46650 -3480 46660 -3420
rect 46580 -3490 46660 -3480
rect 45190 -3610 45270 -3600
rect 45190 -3670 45200 -3610
rect 45260 -3670 45270 -3610
rect 48840 -3640 48850 -3570
rect 48920 -3640 48930 -3570
rect 45190 -3680 45270 -3670
rect 48840 -3690 48930 -3680
rect 48840 -3760 48850 -3690
rect 48920 -3760 48930 -3690
rect 48840 -3770 48930 -3760
rect 44522 -3950 44532 -3880
rect 44602 -3950 44612 -3880
rect 45868 -3950 45878 -3880
rect 45948 -3950 45958 -3880
rect 46420 -3890 46500 -3880
rect 46420 -3950 46430 -3890
rect 46490 -3950 46500 -3890
rect 46420 -3960 46500 -3950
rect 46210 -4100 46290 -4090
rect 46210 -4160 46220 -4100
rect 46280 -4160 46290 -4100
rect 46210 -4170 46290 -4160
rect 43970 -4300 44050 -4290
rect 43970 -4360 43980 -4300
rect 44040 -4360 44050 -4300
rect 43970 -4370 44050 -4360
rect 44522 -4370 44532 -4300
rect 44602 -4370 44612 -4300
rect 45868 -4370 45878 -4300
rect 45948 -4370 45958 -4300
rect 46230 -4530 46270 -4170
rect 46440 -4390 46480 -3960
rect 48860 -4100 48900 -3770
rect 47032 -4170 47042 -4100
rect 47112 -4170 47122 -4100
rect 48430 -4170 48440 -4100
rect 48510 -4170 48520 -4100
rect 48840 -4110 48920 -4100
rect 48840 -4170 48850 -4110
rect 48910 -4170 48920 -4110
rect 48840 -4180 48920 -4170
rect 46420 -4400 46500 -4390
rect 46420 -4460 46430 -4400
rect 46490 -4460 46500 -4400
rect 46420 -4470 46500 -4460
rect 48750 -4400 48830 -4390
rect 48750 -4460 48760 -4400
rect 48820 -4460 48830 -4400
rect 48750 -4470 48830 -4460
rect 48770 -4540 48810 -4470
rect 48860 -4540 48900 -4180
rect 48930 -4310 49010 -4300
rect 48930 -4370 48940 -4310
rect 49000 -4370 49010 -4310
rect 48930 -4380 49010 -4370
rect 48950 -4540 48990 -4380
rect 49040 -4540 49080 -2620
rect 49110 -2720 49190 -2710
rect 49110 -2780 49120 -2720
rect 49180 -2780 49190 -2720
rect 49110 -2790 49190 -2780
rect 49130 -3480 49170 -2790
rect 49110 -3490 49190 -3480
rect 49110 -3550 49120 -3490
rect 49180 -3550 49190 -3490
rect 49110 -3560 49190 -3550
rect 49220 -3490 49250 -3480
rect 49220 -3550 49230 -3490
rect 49220 -3560 49250 -3550
rect 49110 -3670 49190 -3660
rect 49110 -3730 49120 -3670
rect 49180 -3730 49190 -3670
rect 49110 -3740 49190 -3730
rect 49130 -4540 49170 -3740
rect 49240 -4540 49250 -3560
rect 33910 -4630 37330 -4540
rect 33910 -4664 34000 -4630
rect 34034 -4664 34100 -4630
rect 34134 -4664 34200 -4630
rect 34234 -4664 34300 -4630
rect 34334 -4664 34400 -4630
rect 34434 -4664 34500 -4630
rect 34534 -4664 35360 -4630
rect 35394 -4664 35460 -4630
rect 35494 -4664 35560 -4630
rect 35594 -4664 35660 -4630
rect 35694 -4664 35760 -4630
rect 35794 -4664 35860 -4630
rect 35894 -4664 36720 -4630
rect 36754 -4664 36820 -4630
rect 36854 -4664 36920 -4630
rect 36954 -4664 37020 -4630
rect 37054 -4664 37120 -4630
rect 37154 -4664 37220 -4630
rect 37254 -4664 37330 -4630
rect 33910 -4730 37330 -4664
rect 33910 -4764 34000 -4730
rect 34034 -4764 34100 -4730
rect 34134 -4764 34200 -4730
rect 34234 -4764 34300 -4730
rect 34334 -4764 34400 -4730
rect 34434 -4764 34500 -4730
rect 34534 -4764 35360 -4730
rect 35394 -4764 35460 -4730
rect 35494 -4764 35560 -4730
rect 35594 -4764 35660 -4730
rect 35694 -4764 35760 -4730
rect 35794 -4764 35860 -4730
rect 35894 -4764 36720 -4730
rect 36754 -4764 36820 -4730
rect 36854 -4764 36920 -4730
rect 36954 -4764 37020 -4730
rect 37054 -4764 37120 -4730
rect 37154 -4764 37220 -4730
rect 37254 -4764 37330 -4730
rect 33910 -4830 37330 -4764
rect 33910 -4864 34000 -4830
rect 34034 -4864 34100 -4830
rect 34134 -4864 34200 -4830
rect 34234 -4864 34300 -4830
rect 34334 -4864 34400 -4830
rect 34434 -4864 34500 -4830
rect 34534 -4864 35360 -4830
rect 35394 -4864 35460 -4830
rect 35494 -4864 35560 -4830
rect 35594 -4864 35660 -4830
rect 35694 -4864 35760 -4830
rect 35794 -4864 35860 -4830
rect 35894 -4864 36720 -4830
rect 36754 -4864 36820 -4830
rect 36854 -4864 36920 -4830
rect 36954 -4864 37020 -4830
rect 37054 -4864 37120 -4830
rect 37154 -4864 37220 -4830
rect 37254 -4864 37330 -4830
rect 33910 -4930 37330 -4864
rect 33910 -4964 34000 -4930
rect 34034 -4964 34100 -4930
rect 34134 -4964 34200 -4930
rect 34234 -4964 34300 -4930
rect 34334 -4964 34400 -4930
rect 34434 -4964 34500 -4930
rect 34534 -4964 35360 -4930
rect 35394 -4964 35460 -4930
rect 35494 -4964 35560 -4930
rect 35594 -4964 35660 -4930
rect 35694 -4964 35760 -4930
rect 35794 -4964 35860 -4930
rect 35894 -4964 36720 -4930
rect 36754 -4964 36820 -4930
rect 36854 -4964 36920 -4930
rect 36954 -4964 37020 -4930
rect 37054 -4964 37120 -4930
rect 37154 -4964 37220 -4930
rect 37254 -4964 37330 -4930
rect 33910 -5030 37330 -4964
rect 33910 -5064 34000 -5030
rect 34034 -5064 34100 -5030
rect 34134 -5064 34200 -5030
rect 34234 -5064 34300 -5030
rect 34334 -5064 34400 -5030
rect 34434 -5064 34500 -5030
rect 34534 -5064 35360 -5030
rect 35394 -5064 35460 -5030
rect 35494 -5064 35560 -5030
rect 35594 -5064 35660 -5030
rect 35694 -5064 35760 -5030
rect 35794 -5064 35860 -5030
rect 35894 -5064 36720 -5030
rect 36754 -5064 36820 -5030
rect 36854 -5064 36920 -5030
rect 36954 -5064 37020 -5030
rect 37054 -5064 37120 -5030
rect 37154 -5064 37220 -5030
rect 37254 -5064 37330 -5030
rect 33910 -5130 37330 -5064
rect 33910 -5164 34000 -5130
rect 34034 -5164 34100 -5130
rect 34134 -5164 34200 -5130
rect 34234 -5164 34300 -5130
rect 34334 -5164 34400 -5130
rect 34434 -5164 34500 -5130
rect 34534 -5164 35360 -5130
rect 35394 -5164 35460 -5130
rect 35494 -5164 35560 -5130
rect 35594 -5164 35660 -5130
rect 35694 -5164 35760 -5130
rect 35794 -5164 35860 -5130
rect 35894 -5164 36720 -5130
rect 36754 -5164 36820 -5130
rect 36854 -5164 36920 -5130
rect 36954 -5164 37020 -5130
rect 37054 -5164 37120 -5130
rect 37154 -5164 37220 -5130
rect 37254 -5164 37330 -5130
rect 33910 -5240 37330 -5164
rect 33910 -5990 34610 -5240
rect 33910 -6024 34000 -5990
rect 34034 -6024 34100 -5990
rect 34134 -6024 34200 -5990
rect 34234 -6024 34300 -5990
rect 34334 -6024 34400 -5990
rect 34434 -6024 34500 -5990
rect 34534 -6024 34610 -5990
rect 33910 -6090 34610 -6024
rect 33910 -6124 34000 -6090
rect 34034 -6124 34100 -6090
rect 34134 -6124 34200 -6090
rect 34234 -6124 34300 -6090
rect 34334 -6124 34400 -6090
rect 34434 -6124 34500 -6090
rect 34534 -6124 34610 -6090
rect 33910 -6190 34610 -6124
rect 33910 -6224 34000 -6190
rect 34034 -6224 34100 -6190
rect 34134 -6224 34200 -6190
rect 34234 -6224 34300 -6190
rect 34334 -6224 34400 -6190
rect 34434 -6224 34500 -6190
rect 34534 -6224 34610 -6190
rect 33910 -6240 34610 -6224
rect 33580 -6280 34610 -6240
rect 33910 -6290 34610 -6280
rect 33910 -6324 34000 -6290
rect 34034 -6324 34100 -6290
rect 34134 -6324 34200 -6290
rect 34234 -6324 34300 -6290
rect 34334 -6324 34400 -6290
rect 34434 -6324 34500 -6290
rect 34534 -6324 34610 -6290
rect 33910 -6390 34610 -6324
rect 33910 -6424 34000 -6390
rect 34034 -6424 34100 -6390
rect 34134 -6424 34200 -6390
rect 34234 -6424 34300 -6390
rect 34334 -6424 34400 -6390
rect 34434 -6424 34500 -6390
rect 34534 -6424 34610 -6390
rect 33910 -6490 34610 -6424
rect 33910 -6524 34000 -6490
rect 34034 -6524 34100 -6490
rect 34134 -6524 34200 -6490
rect 34234 -6524 34300 -6490
rect 34334 -6524 34400 -6490
rect 34434 -6524 34500 -6490
rect 34534 -6524 34610 -6490
rect 29780 -6560 29860 -6550
rect 29780 -6620 29790 -6560
rect 29850 -6570 29860 -6560
rect 29850 -6610 29880 -6570
rect 29850 -6620 29860 -6610
rect 29780 -6630 29860 -6620
rect 33910 -7260 34610 -6524
rect 35270 -5916 35970 -5906
rect 35270 -5970 35590 -5916
rect 35650 -5970 35970 -5916
rect 35270 -5990 35970 -5970
rect 35270 -6024 35360 -5990
rect 35394 -6024 35460 -5990
rect 35494 -6024 35560 -5990
rect 35594 -6024 35660 -5990
rect 35694 -6024 35760 -5990
rect 35794 -6024 35860 -5990
rect 35894 -6024 35970 -5990
rect 35270 -6090 35970 -6024
rect 35270 -6124 35360 -6090
rect 35394 -6124 35460 -6090
rect 35494 -6124 35560 -6090
rect 35594 -6124 35660 -6090
rect 35694 -6124 35760 -6090
rect 35794 -6124 35860 -6090
rect 35894 -6124 35970 -6090
rect 35270 -6190 35970 -6124
rect 35270 -6224 35360 -6190
rect 35394 -6224 35460 -6190
rect 35494 -6224 35560 -6190
rect 35594 -6224 35660 -6190
rect 35694 -6224 35760 -6190
rect 35794 -6224 35860 -6190
rect 35894 -6224 35970 -6190
rect 35270 -6290 35970 -6224
rect 35270 -6324 35360 -6290
rect 35394 -6324 35460 -6290
rect 35494 -6324 35560 -6290
rect 35594 -6324 35660 -6290
rect 35694 -6324 35760 -6290
rect 35794 -6324 35860 -6290
rect 35894 -6324 35970 -6290
rect 35270 -6390 35970 -6324
rect 35270 -6424 35360 -6390
rect 35394 -6424 35460 -6390
rect 35494 -6424 35560 -6390
rect 35594 -6424 35660 -6390
rect 35694 -6424 35760 -6390
rect 35794 -6424 35860 -6390
rect 35894 -6424 35970 -6390
rect 35270 -6490 35970 -6424
rect 35270 -6524 35360 -6490
rect 35394 -6524 35460 -6490
rect 35494 -6524 35560 -6490
rect 35594 -6524 35660 -6490
rect 35694 -6524 35760 -6490
rect 35794 -6524 35860 -6490
rect 35894 -6524 35970 -6490
rect 35270 -6606 35970 -6524
rect 36630 -5990 37330 -5240
rect 36630 -6024 36720 -5990
rect 36754 -6024 36820 -5990
rect 36854 -6024 36920 -5990
rect 36954 -6024 37020 -5990
rect 37054 -6024 37120 -5990
rect 37154 -6024 37220 -5990
rect 37254 -6024 37330 -5990
rect 36630 -6090 37330 -6024
rect 36630 -6124 36720 -6090
rect 36754 -6124 36820 -6090
rect 36854 -6124 36920 -6090
rect 36954 -6124 37020 -6090
rect 37054 -6124 37120 -6090
rect 37154 -6124 37220 -6090
rect 37254 -6124 37330 -6090
rect 36630 -6190 37330 -6124
rect 36630 -6224 36720 -6190
rect 36754 -6224 36820 -6190
rect 36854 -6224 36920 -6190
rect 36954 -6224 37020 -6190
rect 37054 -6224 37120 -6190
rect 37154 -6224 37220 -6190
rect 37254 -6224 37330 -6190
rect 36630 -6290 37330 -6224
rect 36630 -6324 36720 -6290
rect 36754 -6324 36820 -6290
rect 36854 -6324 36920 -6290
rect 36954 -6324 37020 -6290
rect 37054 -6324 37120 -6290
rect 37154 -6324 37220 -6290
rect 37254 -6324 37330 -6290
rect 36630 -6390 37330 -6324
rect 36630 -6424 36720 -6390
rect 36754 -6424 36820 -6390
rect 36854 -6424 36920 -6390
rect 36954 -6424 37020 -6390
rect 37054 -6424 37120 -6390
rect 37154 -6424 37220 -6390
rect 37254 -6424 37330 -6390
rect 36630 -6490 37330 -6424
rect 36630 -6524 36720 -6490
rect 36754 -6524 36820 -6490
rect 36854 -6524 36920 -6490
rect 36954 -6524 37020 -6490
rect 37054 -6524 37120 -6490
rect 37154 -6524 37220 -6490
rect 37254 -6524 37330 -6490
rect 36630 -7260 37330 -6524
rect 33910 -7350 37330 -7260
rect 33910 -7384 34000 -7350
rect 34034 -7384 34100 -7350
rect 34134 -7384 34200 -7350
rect 34234 -7384 34300 -7350
rect 34334 -7384 34400 -7350
rect 34434 -7384 34500 -7350
rect 34534 -7384 35360 -7350
rect 35394 -7384 35460 -7350
rect 35494 -7384 35560 -7350
rect 35594 -7384 35660 -7350
rect 35694 -7384 35760 -7350
rect 35794 -7384 35860 -7350
rect 35894 -7384 36720 -7350
rect 36754 -7384 36820 -7350
rect 36854 -7384 36920 -7350
rect 36954 -7384 37020 -7350
rect 37054 -7384 37120 -7350
rect 37154 -7384 37220 -7350
rect 37254 -7384 37330 -7350
rect 33910 -7450 37330 -7384
rect 33910 -7484 34000 -7450
rect 34034 -7484 34100 -7450
rect 34134 -7484 34200 -7450
rect 34234 -7484 34300 -7450
rect 34334 -7484 34400 -7450
rect 34434 -7484 34500 -7450
rect 34534 -7484 35360 -7450
rect 35394 -7484 35460 -7450
rect 35494 -7484 35560 -7450
rect 35594 -7484 35660 -7450
rect 35694 -7484 35760 -7450
rect 35794 -7484 35860 -7450
rect 35894 -7484 36720 -7450
rect 36754 -7484 36820 -7450
rect 36854 -7484 36920 -7450
rect 36954 -7484 37020 -7450
rect 37054 -7484 37120 -7450
rect 37154 -7484 37220 -7450
rect 37254 -7484 37330 -7450
rect 33910 -7550 37330 -7484
rect 33910 -7584 34000 -7550
rect 34034 -7584 34100 -7550
rect 34134 -7584 34200 -7550
rect 34234 -7584 34300 -7550
rect 34334 -7584 34400 -7550
rect 34434 -7584 34500 -7550
rect 34534 -7584 35360 -7550
rect 35394 -7584 35460 -7550
rect 35494 -7584 35560 -7550
rect 35594 -7584 35660 -7550
rect 35694 -7584 35760 -7550
rect 35794 -7584 35860 -7550
rect 35894 -7584 36720 -7550
rect 36754 -7584 36820 -7550
rect 36854 -7584 36920 -7550
rect 36954 -7584 37020 -7550
rect 37054 -7584 37120 -7550
rect 37154 -7584 37220 -7550
rect 37254 -7584 37330 -7550
rect 33910 -7650 37330 -7584
rect 33910 -7684 34000 -7650
rect 34034 -7684 34100 -7650
rect 34134 -7684 34200 -7650
rect 34234 -7684 34300 -7650
rect 34334 -7684 34400 -7650
rect 34434 -7684 34500 -7650
rect 34534 -7684 35360 -7650
rect 35394 -7684 35460 -7650
rect 35494 -7684 35560 -7650
rect 35594 -7684 35660 -7650
rect 35694 -7684 35760 -7650
rect 35794 -7684 35860 -7650
rect 35894 -7684 36720 -7650
rect 36754 -7684 36820 -7650
rect 36854 -7684 36920 -7650
rect 36954 -7684 37020 -7650
rect 37054 -7684 37120 -7650
rect 37154 -7684 37220 -7650
rect 37254 -7684 37330 -7650
rect 33910 -7750 37330 -7684
rect 33910 -7784 34000 -7750
rect 34034 -7784 34100 -7750
rect 34134 -7784 34200 -7750
rect 34234 -7784 34300 -7750
rect 34334 -7784 34400 -7750
rect 34434 -7784 34500 -7750
rect 34534 -7784 35360 -7750
rect 35394 -7784 35460 -7750
rect 35494 -7784 35560 -7750
rect 35594 -7784 35660 -7750
rect 35694 -7784 35760 -7750
rect 35794 -7784 35860 -7750
rect 35894 -7784 36720 -7750
rect 36754 -7784 36820 -7750
rect 36854 -7784 36920 -7750
rect 36954 -7784 37020 -7750
rect 37054 -7784 37120 -7750
rect 37154 -7784 37220 -7750
rect 37254 -7784 37330 -7750
rect 33910 -7850 37330 -7784
rect 33910 -7884 34000 -7850
rect 34034 -7884 34100 -7850
rect 34134 -7884 34200 -7850
rect 34234 -7884 34300 -7850
rect 34334 -7884 34400 -7850
rect 34434 -7884 34500 -7850
rect 34534 -7884 35360 -7850
rect 35394 -7884 35460 -7850
rect 35494 -7884 35560 -7850
rect 35594 -7884 35660 -7850
rect 35694 -7884 35760 -7850
rect 35794 -7884 35860 -7850
rect 35894 -7884 36720 -7850
rect 36754 -7884 36820 -7850
rect 36854 -7884 36920 -7850
rect 36954 -7884 37020 -7850
rect 37054 -7884 37120 -7850
rect 37154 -7884 37220 -7850
rect 37254 -7884 37330 -7850
rect 33910 -7960 37330 -7884
rect 35560 -8530 35640 -8520
rect 35560 -8590 35570 -8530
rect 35630 -8590 35640 -8530
rect 35560 -8600 35640 -8590
rect 35580 -8630 35620 -8600
<< via1 >>
rect 2710 7690 2770 7750
rect -20 7530 40 7590
rect 1890 7530 1950 7590
rect -110 7420 -50 7480
rect -110 6050 -50 6110
rect 2520 7320 2580 7380
rect 150 7220 210 7280
rect 142 7170 212 7180
rect 142 7120 152 7170
rect 152 7120 202 7170
rect 202 7120 212 7170
rect 142 7110 212 7120
rect 142 7050 212 7060
rect 142 7000 152 7050
rect 152 7000 202 7050
rect 202 7000 212 7050
rect 142 6990 212 7000
rect 8890 7630 8950 7690
rect 32710 7690 32770 7750
rect 3290 7530 3350 7590
rect 5030 7540 5090 7600
rect 9320 7530 9380 7590
rect 2712 6900 2782 6910
rect 2712 6850 2722 6900
rect 2722 6850 2772 6900
rect 2772 6850 2782 6900
rect 2712 6840 2782 6850
rect 150 6690 210 6750
rect 2520 6690 2580 6750
rect 2712 6780 2782 6790
rect 2712 6730 2722 6780
rect 2722 6730 2772 6780
rect 2772 6730 2782 6780
rect 2712 6720 2782 6730
rect 142 6640 212 6650
rect 142 6590 152 6640
rect 152 6590 202 6640
rect 202 6590 212 6640
rect 142 6580 212 6590
rect 142 6520 212 6530
rect 142 6470 152 6520
rect 152 6470 202 6520
rect 202 6470 212 6520
rect 142 6460 212 6470
rect 2380 6570 2440 6580
rect 2380 6530 2390 6570
rect 2390 6530 2430 6570
rect 2430 6530 2440 6570
rect 2380 6520 2440 6530
rect 2590 6570 2650 6580
rect 2590 6530 2600 6570
rect 2600 6530 2640 6570
rect 2640 6530 2650 6570
rect 2590 6520 2650 6530
rect 1200 6380 1260 6390
rect 1200 6340 1210 6380
rect 1210 6340 1250 6380
rect 1250 6340 1260 6380
rect 1200 6330 1260 6340
rect 4850 6420 4920 6430
rect 4850 6370 4860 6420
rect 4860 6370 4910 6420
rect 4910 6370 4920 6420
rect 4850 6360 4920 6370
rect 4850 6300 4920 6310
rect 4850 6250 4860 6300
rect 4860 6250 4910 6300
rect 4910 6250 4920 6300
rect 4850 6240 4920 6250
rect 532 6110 602 6120
rect 532 6060 542 6110
rect 542 6060 592 6110
rect 592 6060 602 6110
rect 532 6050 602 6060
rect 1878 6110 1948 6120
rect 1878 6060 1888 6110
rect 1888 6060 1938 6110
rect 1938 6060 1948 6110
rect 1878 6050 1948 6060
rect 2430 6050 2490 6110
rect 2220 5840 2280 5900
rect -20 5640 40 5700
rect 532 5690 602 5700
rect 532 5640 542 5690
rect 542 5640 592 5690
rect 592 5640 602 5690
rect 532 5630 602 5640
rect 1878 5690 1948 5700
rect 1878 5640 1888 5690
rect 1888 5640 1938 5690
rect 1938 5640 1948 5690
rect 1878 5630 1948 5640
rect 3042 5890 3112 5900
rect 3042 5840 3052 5890
rect 3052 5840 3102 5890
rect 3102 5840 3112 5890
rect 3042 5830 3112 5840
rect 4440 5890 4510 5900
rect 4440 5840 4450 5890
rect 4450 5840 4500 5890
rect 4500 5840 4510 5890
rect 4440 5830 4510 5840
rect 4850 5830 4910 5890
rect 2430 5540 2490 5600
rect 4760 5540 4820 5600
rect 4670 5220 4730 5280
rect 4560 5130 4620 5190
rect -210 3380 -150 3440
rect -80 3430 -20 3440
rect -80 3390 -70 3430
rect -70 3390 -30 3430
rect -30 3390 -20 3430
rect -80 3380 -20 3390
rect 2540 3360 2594 3420
rect 4940 5630 5000 5690
rect 4850 5330 4910 5390
rect 4760 4940 4820 5000
rect 4670 4030 4730 4090
rect 4940 4690 5000 4750
rect 10290 7530 10350 7590
rect 5390 7420 5450 7480
rect 6790 7420 6850 7480
rect 9230 7420 9290 7480
rect 8570 7320 8630 7380
rect 5120 7220 5180 7280
rect 6630 7210 6690 7270
rect 6410 7120 6470 7180
rect 8130 7120 8190 7180
rect 9140 7120 9200 7180
rect 6080 7050 6140 7060
rect 6080 7010 6090 7050
rect 6090 7010 6130 7050
rect 6130 7010 6140 7050
rect 6080 7000 6140 7010
rect 6300 7050 6360 7060
rect 6300 7010 6310 7050
rect 6310 7010 6350 7050
rect 6350 7010 6360 7050
rect 6300 7000 6360 7010
rect 6520 7050 6580 7060
rect 6520 7010 6530 7050
rect 6530 7010 6570 7050
rect 6570 7010 6580 7050
rect 6520 7000 6580 7010
rect 6740 7050 6800 7060
rect 6740 7010 6750 7050
rect 6750 7010 6790 7050
rect 6790 7010 6800 7050
rect 6740 7000 6800 7010
rect 7360 7050 7420 7060
rect 7360 7010 7370 7050
rect 7370 7010 7410 7050
rect 7410 7010 7420 7050
rect 7360 7000 7420 7010
rect 7580 7050 7640 7060
rect 7580 7010 7590 7050
rect 7590 7010 7630 7050
rect 7630 7010 7640 7050
rect 7580 7000 7640 7010
rect 7800 7050 7860 7060
rect 7800 7010 7810 7050
rect 7810 7010 7850 7050
rect 7850 7010 7860 7050
rect 7800 7000 7860 7010
rect 8020 7050 8080 7060
rect 8020 7010 8030 7050
rect 8030 7010 8070 7050
rect 8070 7010 8080 7050
rect 8020 7000 8080 7010
rect 8240 7050 8300 7060
rect 8240 7010 8250 7050
rect 8250 7010 8290 7050
rect 8290 7010 8300 7050
rect 8240 7000 8300 7010
rect 8460 7050 8520 7060
rect 8460 7010 8470 7050
rect 8470 7010 8510 7050
rect 8510 7010 8520 7050
rect 8460 7000 8520 7010
rect 8680 7050 8740 7060
rect 8680 7010 8690 7050
rect 8690 7010 8730 7050
rect 8730 7010 8740 7050
rect 8680 7000 8740 7010
rect 6190 6710 6250 6720
rect 6190 6670 6200 6710
rect 6200 6670 6240 6710
rect 6240 6670 6250 6710
rect 6190 6660 6250 6670
rect 6410 6710 6470 6720
rect 6410 6670 6420 6710
rect 6420 6670 6460 6710
rect 6460 6670 6470 6710
rect 6410 6660 6470 6670
rect 6630 6710 6690 6720
rect 6630 6670 6640 6710
rect 6640 6670 6680 6710
rect 6680 6670 6690 6710
rect 6630 6660 6690 6670
rect 7690 6710 7750 6720
rect 7690 6670 7700 6710
rect 7700 6670 7740 6710
rect 7740 6670 7750 6710
rect 7690 6660 7750 6670
rect 7910 6710 7970 6720
rect 7910 6670 7920 6710
rect 7920 6670 7960 6710
rect 7960 6670 7970 6710
rect 7910 6660 7970 6670
rect 8130 6710 8190 6720
rect 8130 6670 8140 6710
rect 8140 6670 8180 6710
rect 8180 6670 8190 6710
rect 8130 6660 8190 6670
rect 8350 6710 8410 6720
rect 8350 6670 8360 6710
rect 8360 6670 8400 6710
rect 8400 6670 8410 6710
rect 8350 6660 8410 6670
rect 5120 6450 5180 6510
rect 5230 6450 5290 6510
rect 5120 6270 5180 6330
rect 5030 4230 5090 4290
rect 4850 3700 4910 3760
rect 4670 3360 4730 3420
rect 4560 2280 4620 2340
rect 6130 6360 6190 6420
rect 5660 6040 5720 6050
rect 5660 6000 5670 6040
rect 5670 6000 5710 6040
rect 5710 6000 5720 6040
rect 5660 5990 5720 6000
rect 7470 6270 7530 6330
rect 9140 6570 9200 6630
rect 9230 6460 9290 6520
rect 29980 7530 30040 7590
rect 31890 7530 31950 7590
rect 29890 7420 29950 7480
rect 38890 7630 38950 7690
rect 33290 7530 33350 7590
rect 35030 7540 35090 7600
rect 39320 7530 39380 7590
rect 40290 7530 40350 7590
rect 35390 7420 35450 7480
rect 36790 7420 36850 7480
rect 39230 7420 39290 7480
rect 38570 7320 38630 7380
rect 9850 7120 9910 7180
rect 9520 7050 9580 7060
rect 9520 7010 9530 7050
rect 9530 7010 9570 7050
rect 9570 7010 9580 7050
rect 9520 7000 9580 7010
rect 9740 7050 9800 7060
rect 9740 7010 9750 7050
rect 9750 7010 9790 7050
rect 9790 7010 9800 7050
rect 9740 7000 9800 7010
rect 9960 7050 10020 7060
rect 9960 7010 9970 7050
rect 9970 7010 10010 7050
rect 10010 7010 10020 7050
rect 9960 7000 10020 7010
rect 10180 7050 10240 7060
rect 10180 7010 10190 7050
rect 10190 7010 10230 7050
rect 10230 7010 10240 7050
rect 10180 7000 10240 7010
rect 9630 6710 9690 6720
rect 9630 6670 9640 6710
rect 9640 6670 9680 6710
rect 9680 6670 9690 6710
rect 9630 6660 9690 6670
rect 9850 6710 9910 6720
rect 9850 6670 9860 6710
rect 9860 6670 9900 6710
rect 9900 6670 9910 6710
rect 9850 6660 9910 6670
rect 10070 6710 10130 6720
rect 10070 6670 10080 6710
rect 10080 6670 10120 6710
rect 10120 6670 10130 6710
rect 10070 6660 10130 6670
rect 9950 6550 10010 6610
rect 9320 6350 9380 6410
rect 8570 6260 8630 6320
rect 8130 6190 8190 6250
rect 6510 6120 6570 6130
rect 6510 6080 6520 6120
rect 6520 6080 6560 6120
rect 6560 6080 6570 6120
rect 6510 6070 6570 6080
rect 6870 6120 6930 6130
rect 6870 6080 6880 6120
rect 6880 6080 6920 6120
rect 6920 6080 6930 6120
rect 6870 6070 6930 6080
rect 7230 6120 7290 6130
rect 7230 6080 7240 6120
rect 7240 6080 7280 6120
rect 7280 6080 7290 6120
rect 7230 6070 7290 6080
rect 7590 6120 7650 6130
rect 7590 6080 7600 6120
rect 7600 6080 7640 6120
rect 7640 6080 7650 6120
rect 7590 6070 7650 6080
rect 7950 6120 8010 6130
rect 7950 6080 7960 6120
rect 7960 6080 8000 6120
rect 8000 6080 8010 6120
rect 7950 6070 8010 6080
rect 8310 6120 8370 6130
rect 8310 6080 8320 6120
rect 8320 6080 8360 6120
rect 8360 6080 8370 6120
rect 8310 6070 8370 6080
rect 8670 6120 8730 6130
rect 8670 6080 8680 6120
rect 8680 6080 8720 6120
rect 8720 6080 8730 6120
rect 8670 6070 8730 6080
rect 9030 6120 9090 6130
rect 9030 6080 9040 6120
rect 9040 6080 9080 6120
rect 9080 6080 9090 6120
rect 9030 6070 9090 6080
rect 9390 6120 9450 6130
rect 9390 6080 9400 6120
rect 9400 6080 9440 6120
rect 9440 6080 9450 6120
rect 9390 6070 9450 6080
rect 9750 6120 9810 6130
rect 9750 6080 9760 6120
rect 9760 6080 9800 6120
rect 9800 6080 9810 6120
rect 9750 6070 9810 6080
rect 5660 5920 5720 5930
rect 5660 5880 5670 5920
rect 5670 5880 5710 5920
rect 5710 5880 5720 5920
rect 5660 5870 5720 5880
rect 6130 5870 6190 5930
rect 5530 5580 5590 5590
rect 5530 5540 5540 5580
rect 5540 5540 5580 5580
rect 5580 5540 5590 5580
rect 5530 5530 5590 5540
rect 5790 5580 5850 5590
rect 5790 5540 5800 5580
rect 5800 5540 5840 5580
rect 5840 5540 5850 5580
rect 5790 5530 5850 5540
rect 6250 5530 6310 5590
rect 6130 5220 6190 5280
rect 5660 5130 5720 5190
rect 5230 5040 5290 5100
rect 5650 4810 5710 4870
rect 5890 4810 5950 4870
rect 6130 4810 6190 4870
rect 7770 5380 7830 5390
rect 7770 5340 7780 5380
rect 7780 5340 7820 5380
rect 7820 5340 7830 5380
rect 7770 5330 7830 5340
rect 8490 5380 8550 5390
rect 8490 5340 8500 5380
rect 8500 5340 8540 5380
rect 8540 5340 8550 5380
rect 8490 5330 8550 5340
rect 7410 5220 7470 5280
rect 7050 5130 7110 5190
rect 6690 5040 6750 5100
rect 6370 4810 6430 4870
rect 6610 4860 6670 4870
rect 6610 4820 6620 4860
rect 6620 4820 6660 4860
rect 6660 4820 6670 4860
rect 6610 4810 6670 4820
rect 6850 4810 6910 4870
rect 7090 4810 7150 4870
rect 7330 4810 7390 4870
rect 7570 4810 7630 4870
rect 8850 5220 8910 5280
rect 9210 5130 9270 5190
rect 9390 5130 9450 5190
rect 8130 5040 8190 5100
rect 9570 5040 9630 5100
rect 10130 6460 10190 6520
rect 10040 6350 10100 6410
rect 11240 6260 11300 6320
rect 10590 6040 10650 6050
rect 10590 6000 10600 6040
rect 10600 6000 10640 6040
rect 10640 6000 10650 6040
rect 10590 5990 10650 6000
rect 10590 5920 10650 5930
rect 10590 5880 10600 5920
rect 10600 5880 10640 5920
rect 10640 5880 10650 5920
rect 10590 5870 10650 5880
rect 10460 5580 10520 5590
rect 10460 5540 10470 5580
rect 10470 5540 10510 5580
rect 10510 5540 10520 5580
rect 10460 5530 10520 5540
rect 10720 5580 10780 5590
rect 10720 5540 10730 5580
rect 10730 5540 10770 5580
rect 10770 5540 10780 5580
rect 10720 5530 10780 5540
rect 10130 5240 10190 5300
rect 10040 5130 10100 5190
rect 11060 5240 11120 5300
rect 8570 4940 8630 5000
rect 9950 4940 10010 5000
rect 10590 4940 10650 5000
rect 8690 4860 8750 4870
rect 8690 4820 8700 4860
rect 8700 4820 8740 4860
rect 8740 4820 8750 4860
rect 8690 4810 8750 4820
rect 8930 4860 8990 4870
rect 8930 4820 8940 4860
rect 8940 4820 8980 4860
rect 8980 4820 8990 4860
rect 8930 4810 8990 4820
rect 9170 4860 9230 4870
rect 9170 4820 9180 4860
rect 9180 4820 9220 4860
rect 9220 4820 9230 4860
rect 9170 4810 9230 4820
rect 9410 4860 9470 4870
rect 9410 4820 9420 4860
rect 9420 4820 9460 4860
rect 9460 4820 9470 4860
rect 9410 4810 9470 4820
rect 9650 4860 9710 4870
rect 9650 4820 9660 4860
rect 9660 4820 9700 4860
rect 9700 4820 9710 4860
rect 9650 4810 9710 4820
rect 9890 4860 9950 4870
rect 9890 4820 9900 4860
rect 9900 4820 9940 4860
rect 9940 4820 9950 4860
rect 9890 4810 9950 4820
rect 10130 4860 10190 4870
rect 10130 4820 10140 4860
rect 10140 4820 10180 4860
rect 10180 4820 10190 4860
rect 10130 4810 10190 4820
rect 10370 4860 10430 4870
rect 10370 4820 10380 4860
rect 10380 4820 10420 4860
rect 10420 4820 10430 4860
rect 10370 4810 10430 4820
rect 10610 4860 10670 4870
rect 10610 4820 10620 4860
rect 10620 4820 10660 4860
rect 10660 4820 10670 4860
rect 10610 4810 10670 4820
rect 5530 4740 5590 4750
rect 5530 4700 5540 4740
rect 5540 4700 5580 4740
rect 5580 4700 5590 4740
rect 5530 4690 5590 4700
rect 6250 4740 6310 4750
rect 6250 4700 6260 4740
rect 6260 4700 6300 4740
rect 6300 4700 6310 4740
rect 6250 4690 6310 4700
rect 6970 4740 7030 4750
rect 6970 4700 6980 4740
rect 6980 4700 7020 4740
rect 7020 4700 7030 4740
rect 6970 4690 7030 4700
rect 7690 4740 7750 4750
rect 7690 4700 7700 4740
rect 7700 4700 7740 4740
rect 7740 4700 7750 4740
rect 7690 4690 7750 4700
rect 7950 4690 8010 4750
rect 8310 4690 8370 4750
rect 8570 4740 8630 4750
rect 8570 4700 8580 4740
rect 8580 4700 8620 4740
rect 8620 4700 8630 4740
rect 8570 4690 8630 4700
rect 9290 4740 9350 4750
rect 9290 4700 9300 4740
rect 9300 4700 9340 4740
rect 9340 4700 9350 4740
rect 9290 4690 9350 4700
rect 10010 4740 10070 4750
rect 10010 4700 10020 4740
rect 10020 4700 10060 4740
rect 10060 4700 10070 4740
rect 10010 4690 10070 4700
rect 10730 4740 10790 4750
rect 10730 4700 10740 4740
rect 10740 4700 10780 4740
rect 10780 4700 10790 4740
rect 10730 4690 10790 4700
rect 5770 4400 5830 4410
rect 5770 4360 5780 4400
rect 5780 4360 5820 4400
rect 5820 4360 5830 4400
rect 5770 4350 5830 4360
rect 6490 4400 6550 4410
rect 6490 4360 6500 4400
rect 6500 4360 6540 4400
rect 6540 4360 6550 4400
rect 6490 4350 6550 4360
rect 7210 4400 7270 4410
rect 7210 4360 7220 4400
rect 7220 4360 7260 4400
rect 7260 4360 7270 4400
rect 7210 4350 7270 4360
rect 5590 4230 5650 4290
rect 6010 4230 6070 4290
rect 6250 4230 6310 4290
rect 6730 4230 6790 4290
rect 6970 4230 7030 4290
rect 7450 4230 7510 4290
rect 7630 4230 7690 4290
rect 6390 4080 6450 4090
rect 6390 4040 6400 4080
rect 6400 4040 6440 4080
rect 6440 4040 6450 4080
rect 6390 4030 6450 4040
rect 6510 4060 6570 4120
rect 6990 4060 7050 4120
rect 7470 4060 7530 4120
rect 6270 3990 6330 4000
rect 6270 3950 6280 3990
rect 6280 3950 6320 3990
rect 6320 3950 6330 3990
rect 6270 3940 6330 3950
rect 6750 3990 6810 4000
rect 6750 3950 6760 3990
rect 6760 3950 6800 3990
rect 6800 3950 6810 3990
rect 6750 3940 6810 3950
rect 7230 3990 7290 4000
rect 7230 3950 7240 3990
rect 7240 3950 7280 3990
rect 7280 3950 7290 3990
rect 7230 3940 7290 3950
rect 7590 3870 7650 3880
rect 7590 3830 7600 3870
rect 7600 3830 7640 3870
rect 7640 3830 7650 3870
rect 7590 3820 7650 3830
rect 6270 3750 6330 3760
rect 6270 3710 6280 3750
rect 6280 3710 6320 3750
rect 6320 3710 6330 3750
rect 6270 3700 6330 3710
rect 5790 3580 5850 3640
rect 6390 3580 6450 3640
rect 6630 3580 6690 3640
rect 6870 3580 6930 3640
rect 7110 3580 7170 3640
rect 7350 3580 7410 3640
rect 5970 3430 6030 3440
rect 5970 3390 5980 3430
rect 5980 3390 6020 3430
rect 6020 3390 6030 3430
rect 5970 3380 6030 3390
rect 6210 3430 6270 3440
rect 6210 3390 6220 3430
rect 6220 3390 6260 3430
rect 6260 3390 6270 3430
rect 6210 3380 6270 3390
rect 6450 3430 6510 3440
rect 6450 3390 6460 3430
rect 6460 3390 6500 3430
rect 6500 3390 6510 3430
rect 6450 3380 6510 3390
rect 6690 3430 6750 3440
rect 6690 3390 6700 3430
rect 6700 3390 6740 3430
rect 6740 3390 6750 3430
rect 6690 3380 6750 3390
rect 7170 3430 7230 3440
rect 7170 3390 7180 3430
rect 7180 3390 7220 3430
rect 7220 3390 7230 3430
rect 7170 3380 7230 3390
rect 7410 3430 7470 3440
rect 7410 3390 7420 3430
rect 7420 3390 7460 3430
rect 7460 3390 7470 3430
rect 7410 3380 7470 3390
rect 7650 3430 7710 3440
rect 7650 3390 7660 3430
rect 7660 3390 7700 3430
rect 7700 3390 7710 3430
rect 7650 3380 7710 3390
rect 8130 3820 8190 3880
rect 9050 4400 9110 4410
rect 9050 4360 9060 4400
rect 9060 4360 9100 4400
rect 9100 4360 9110 4400
rect 9050 4350 9110 4360
rect 9770 4400 9830 4410
rect 9770 4360 9780 4400
rect 9780 4360 9820 4400
rect 9820 4360 9830 4400
rect 9770 4350 9830 4360
rect 10490 4400 10550 4410
rect 10490 4360 10500 4400
rect 10500 4360 10540 4400
rect 10540 4360 10550 4400
rect 10490 4350 10550 4360
rect 8630 4230 8690 4290
rect 8810 4230 8870 4290
rect 9290 4230 9350 4290
rect 9530 4230 9590 4290
rect 8790 4060 8850 4120
rect 9270 4060 9330 4120
rect 11150 5040 11210 5100
rect 10010 4230 10070 4290
rect 10250 4230 10310 4290
rect 10670 4230 10730 4290
rect 11060 4230 11120 4290
rect 9750 4060 9810 4120
rect 9870 4080 9930 4090
rect 9870 4040 9880 4080
rect 9880 4040 9920 4080
rect 9920 4040 9930 4080
rect 9870 4030 9930 4040
rect 11150 4030 11210 4090
rect 9030 3990 9090 4000
rect 9030 3950 9040 3990
rect 9040 3950 9080 3990
rect 9080 3950 9090 3990
rect 9030 3940 9090 3950
rect 9510 3990 9570 4000
rect 9510 3950 9520 3990
rect 9520 3950 9560 3990
rect 9560 3950 9570 3990
rect 9510 3940 9570 3950
rect 9990 3990 10050 4000
rect 9990 3950 10000 3990
rect 10000 3950 10040 3990
rect 10040 3950 10050 3990
rect 9990 3940 10050 3950
rect 8670 3870 8730 3880
rect 8670 3830 8680 3870
rect 8680 3830 8720 3870
rect 8720 3830 8730 3870
rect 8670 3820 8730 3830
rect 36630 4210 36690 4270
rect 36410 4120 36470 4180
rect 38130 4120 38190 4180
rect 39140 4120 39200 4180
rect 36080 4050 36140 4060
rect 36080 4010 36090 4050
rect 36090 4010 36130 4050
rect 36130 4010 36140 4050
rect 36080 4000 36140 4010
rect 36300 4050 36360 4060
rect 36300 4010 36310 4050
rect 36310 4010 36350 4050
rect 36350 4010 36360 4050
rect 36300 4000 36360 4010
rect 36520 4050 36580 4060
rect 36520 4010 36530 4050
rect 36530 4010 36570 4050
rect 36570 4010 36580 4050
rect 36520 4000 36580 4010
rect 36740 4050 36800 4060
rect 36740 4010 36750 4050
rect 36750 4010 36790 4050
rect 36790 4010 36800 4050
rect 36740 4000 36800 4010
rect 37360 4050 37420 4060
rect 37360 4010 37370 4050
rect 37370 4010 37410 4050
rect 37410 4010 37420 4050
rect 37360 4000 37420 4010
rect 37580 4050 37640 4060
rect 37580 4010 37590 4050
rect 37590 4010 37630 4050
rect 37630 4010 37640 4050
rect 37580 4000 37640 4010
rect 37800 4050 37860 4060
rect 37800 4010 37810 4050
rect 37810 4010 37850 4050
rect 37850 4010 37860 4050
rect 37800 4000 37860 4010
rect 38020 4050 38080 4060
rect 38020 4010 38030 4050
rect 38030 4010 38070 4050
rect 38070 4010 38080 4050
rect 38020 4000 38080 4010
rect 38240 4050 38300 4060
rect 38240 4010 38250 4050
rect 38250 4010 38290 4050
rect 38290 4010 38300 4050
rect 38240 4000 38300 4010
rect 38460 4050 38520 4060
rect 38460 4010 38470 4050
rect 38470 4010 38510 4050
rect 38510 4010 38520 4050
rect 38460 4000 38520 4010
rect 38680 4050 38740 4060
rect 38680 4010 38690 4050
rect 38690 4010 38730 4050
rect 38730 4010 38740 4050
rect 38680 4000 38740 4010
rect 9990 3750 10050 3760
rect 9990 3710 10000 3750
rect 10000 3710 10040 3750
rect 10040 3710 10050 3750
rect 9990 3700 10050 3710
rect 11240 3700 11300 3760
rect 36190 3710 36250 3720
rect 36190 3670 36200 3710
rect 36200 3670 36240 3710
rect 36240 3670 36250 3710
rect 36190 3660 36250 3670
rect 36410 3710 36470 3720
rect 36410 3670 36420 3710
rect 36420 3670 36460 3710
rect 36460 3670 36470 3710
rect 36410 3660 36470 3670
rect 36630 3710 36690 3720
rect 36630 3670 36640 3710
rect 36640 3670 36680 3710
rect 36680 3670 36690 3710
rect 36630 3660 36690 3670
rect 37690 3710 37750 3720
rect 37690 3670 37700 3710
rect 37700 3670 37740 3710
rect 37740 3670 37750 3710
rect 37690 3660 37750 3670
rect 37910 3710 37970 3720
rect 37910 3670 37920 3710
rect 37920 3670 37960 3710
rect 37960 3670 37970 3710
rect 37910 3660 37970 3670
rect 38130 3710 38190 3720
rect 38130 3670 38140 3710
rect 38140 3670 38180 3710
rect 38180 3670 38190 3710
rect 38130 3660 38190 3670
rect 38350 3710 38410 3720
rect 38350 3670 38360 3710
rect 38360 3670 38400 3710
rect 38400 3670 38410 3710
rect 38350 3660 38410 3670
rect 8910 3580 8970 3640
rect 9150 3580 9210 3640
rect 9390 3580 9450 3640
rect 9630 3580 9690 3640
rect 9870 3580 9930 3640
rect 10470 3580 10530 3640
rect 8610 3430 8670 3440
rect 8610 3390 8620 3430
rect 8620 3390 8660 3430
rect 8660 3390 8670 3430
rect 8610 3380 8670 3390
rect 8850 3430 8910 3440
rect 8850 3390 8860 3430
rect 8860 3390 8900 3430
rect 8900 3390 8910 3430
rect 8850 3380 8910 3390
rect 9090 3430 9150 3440
rect 9090 3390 9100 3430
rect 9100 3390 9140 3430
rect 9140 3390 9150 3430
rect 9090 3380 9150 3390
rect 9570 3430 9630 3440
rect 9570 3390 9580 3430
rect 9580 3390 9620 3430
rect 9620 3390 9630 3430
rect 9570 3380 9630 3390
rect 9810 3430 9870 3440
rect 9810 3390 9820 3430
rect 9820 3390 9860 3430
rect 9860 3390 9870 3430
rect 9810 3380 9870 3390
rect 10050 3430 10110 3440
rect 10050 3390 10060 3430
rect 10060 3390 10100 3430
rect 10100 3390 10110 3430
rect 10050 3380 10110 3390
rect 10290 3430 10350 3440
rect 10290 3390 10300 3430
rect 10300 3390 10340 3430
rect 10340 3390 10350 3430
rect 10290 3380 10350 3390
rect 6870 2800 6930 2810
rect 6870 2760 6880 2800
rect 6880 2760 6920 2800
rect 6920 2760 6930 2800
rect 6870 2750 6930 2760
rect 8130 2750 8190 2810
rect 9390 2800 9450 2810
rect 9390 2760 9400 2800
rect 9400 2760 9440 2800
rect 9440 2760 9450 2800
rect 9390 2750 9450 2760
rect 8130 2600 8190 2620
rect 8130 2560 8140 2600
rect 8140 2560 8180 2600
rect 8180 2560 8190 2600
rect 6050 2500 6110 2510
rect 6050 2460 6060 2500
rect 6060 2460 6100 2500
rect 6100 2460 6110 2500
rect 6050 2450 6110 2460
rect 6210 2500 6270 2510
rect 6210 2460 6220 2500
rect 6220 2460 6260 2500
rect 6260 2460 6270 2500
rect 6210 2450 6270 2460
rect 6370 2500 6430 2510
rect 6370 2460 6380 2500
rect 6380 2460 6420 2500
rect 6420 2460 6430 2500
rect 6370 2450 6430 2460
rect 6530 2500 6590 2510
rect 6530 2460 6540 2500
rect 6540 2460 6580 2500
rect 6580 2460 6590 2500
rect 6530 2450 6590 2460
rect 6690 2500 6750 2510
rect 6690 2460 6700 2500
rect 6700 2460 6740 2500
rect 6740 2460 6750 2500
rect 6690 2450 6750 2460
rect 6850 2500 6910 2510
rect 6850 2460 6860 2500
rect 6860 2460 6900 2500
rect 6900 2460 6910 2500
rect 6850 2450 6910 2460
rect 7010 2500 7070 2510
rect 7010 2460 7020 2500
rect 7020 2460 7060 2500
rect 7060 2460 7070 2500
rect 7010 2450 7070 2460
rect 7170 2500 7230 2510
rect 7170 2460 7180 2500
rect 7180 2460 7220 2500
rect 7220 2460 7230 2500
rect 7170 2450 7230 2460
rect 7330 2500 7390 2510
rect 7330 2460 7340 2500
rect 7340 2460 7380 2500
rect 7380 2460 7390 2500
rect 7330 2450 7390 2460
rect 7490 2500 7550 2510
rect 7490 2460 7500 2500
rect 7500 2460 7540 2500
rect 7540 2460 7550 2500
rect 7490 2450 7550 2460
rect 7650 2500 7710 2510
rect 7650 2460 7660 2500
rect 7660 2460 7700 2500
rect 7700 2460 7710 2500
rect 7650 2450 7710 2460
rect 7810 2500 7870 2510
rect 7810 2460 7820 2500
rect 7820 2460 7860 2500
rect 7860 2460 7870 2500
rect 7810 2450 7870 2460
rect 7970 2500 8030 2510
rect 7970 2460 7980 2500
rect 7980 2460 8020 2500
rect 8020 2460 8030 2500
rect 7970 2450 8030 2460
rect 8130 2500 8190 2510
rect 8130 2460 8140 2500
rect 8140 2460 8180 2500
rect 8180 2460 8190 2500
rect 8130 2450 8190 2460
rect 8290 2500 8350 2510
rect 8290 2460 8300 2500
rect 8300 2460 8340 2500
rect 8340 2460 8350 2500
rect 8290 2450 8350 2460
rect 8450 2500 8510 2510
rect 8450 2460 8460 2500
rect 8460 2460 8500 2500
rect 8500 2460 8510 2500
rect 8450 2450 8510 2460
rect 8610 2500 8670 2510
rect 8610 2460 8620 2500
rect 8620 2460 8660 2500
rect 8660 2460 8670 2500
rect 8610 2450 8670 2460
rect 8770 2500 8830 2510
rect 8770 2460 8780 2500
rect 8780 2460 8820 2500
rect 8820 2460 8830 2500
rect 8770 2450 8830 2460
rect 8930 2500 8990 2510
rect 8930 2460 8940 2500
rect 8940 2460 8980 2500
rect 8980 2460 8990 2500
rect 8930 2450 8990 2460
rect 9090 2500 9150 2510
rect 9090 2460 9100 2500
rect 9100 2460 9140 2500
rect 9140 2460 9150 2500
rect 9090 2450 9150 2460
rect 9250 2500 9310 2510
rect 9250 2460 9260 2500
rect 9260 2460 9300 2500
rect 9300 2460 9310 2500
rect 9250 2450 9310 2460
rect 9410 2500 9470 2510
rect 9410 2460 9420 2500
rect 9420 2460 9460 2500
rect 9460 2460 9470 2500
rect 9410 2450 9470 2460
rect 9570 2500 9630 2510
rect 9570 2460 9580 2500
rect 9580 2460 9620 2500
rect 9620 2460 9630 2500
rect 9570 2450 9630 2460
rect 9730 2500 9790 2510
rect 9730 2460 9740 2500
rect 9740 2460 9780 2500
rect 9780 2460 9790 2500
rect 9730 2450 9790 2460
rect 9890 2500 9950 2510
rect 9890 2460 9900 2500
rect 9900 2460 9940 2500
rect 9940 2460 9950 2500
rect 9890 2450 9950 2460
rect 10050 2500 10110 2510
rect 10050 2460 10060 2500
rect 10060 2460 10100 2500
rect 10100 2460 10110 2500
rect 10050 2450 10110 2460
rect 36130 3360 36190 3420
rect 35660 3040 35720 3050
rect 35660 3000 35670 3040
rect 35670 3000 35710 3040
rect 35710 3000 35720 3040
rect 35660 2990 35720 3000
rect 37470 3270 37530 3330
rect 39140 3570 39200 3630
rect 39230 3460 39290 3520
rect 39850 4120 39910 4180
rect 39520 4050 39580 4060
rect 39520 4010 39530 4050
rect 39530 4010 39570 4050
rect 39570 4010 39580 4050
rect 39520 4000 39580 4010
rect 39740 4050 39800 4060
rect 39740 4010 39750 4050
rect 39750 4010 39790 4050
rect 39790 4010 39800 4050
rect 39740 4000 39800 4010
rect 39960 4050 40020 4060
rect 39960 4010 39970 4050
rect 39970 4010 40010 4050
rect 40010 4010 40020 4050
rect 39960 4000 40020 4010
rect 40180 4050 40240 4060
rect 40180 4010 40190 4050
rect 40190 4010 40230 4050
rect 40230 4010 40240 4050
rect 40180 4000 40240 4010
rect 39630 3710 39690 3720
rect 39630 3670 39640 3710
rect 39640 3670 39680 3710
rect 39680 3670 39690 3710
rect 39630 3660 39690 3670
rect 39850 3710 39910 3720
rect 39850 3670 39860 3710
rect 39860 3670 39900 3710
rect 39900 3670 39910 3710
rect 39850 3660 39910 3670
rect 40070 3710 40130 3720
rect 40070 3670 40080 3710
rect 40080 3670 40120 3710
rect 40120 3670 40130 3710
rect 40070 3660 40130 3670
rect 39950 3550 40010 3610
rect 39320 3350 39380 3410
rect 38570 3260 38630 3320
rect 38130 3190 38190 3250
rect 36510 3120 36570 3130
rect 36510 3080 36520 3120
rect 36520 3080 36560 3120
rect 36560 3080 36570 3120
rect 36510 3070 36570 3080
rect 36870 3120 36930 3130
rect 36870 3080 36880 3120
rect 36880 3080 36920 3120
rect 36920 3080 36930 3120
rect 36870 3070 36930 3080
rect 37230 3120 37290 3130
rect 37230 3080 37240 3120
rect 37240 3080 37280 3120
rect 37280 3080 37290 3120
rect 37230 3070 37290 3080
rect 37590 3120 37650 3130
rect 37590 3080 37600 3120
rect 37600 3080 37640 3120
rect 37640 3080 37650 3120
rect 37590 3070 37650 3080
rect 37950 3120 38010 3130
rect 37950 3080 37960 3120
rect 37960 3080 38000 3120
rect 38000 3080 38010 3120
rect 37950 3070 38010 3080
rect 38310 3120 38370 3130
rect 38310 3080 38320 3120
rect 38320 3080 38360 3120
rect 38360 3080 38370 3120
rect 38310 3070 38370 3080
rect 38670 3120 38730 3130
rect 38670 3080 38680 3120
rect 38680 3080 38720 3120
rect 38720 3080 38730 3120
rect 38670 3070 38730 3080
rect 39030 3120 39090 3130
rect 39030 3080 39040 3120
rect 39040 3080 39080 3120
rect 39080 3080 39090 3120
rect 39030 3070 39090 3080
rect 39390 3120 39450 3130
rect 39390 3080 39400 3120
rect 39400 3080 39440 3120
rect 39440 3080 39450 3120
rect 39390 3070 39450 3080
rect 39750 3120 39810 3130
rect 39750 3080 39760 3120
rect 39760 3080 39800 3120
rect 39800 3080 39810 3120
rect 39750 3070 39810 3080
rect 35660 2920 35720 2930
rect 35660 2880 35670 2920
rect 35670 2880 35710 2920
rect 35710 2880 35720 2920
rect 35660 2870 35720 2880
rect 36130 2870 36190 2930
rect 35530 2580 35590 2590
rect 35530 2540 35540 2580
rect 35540 2540 35580 2580
rect 35580 2540 35590 2580
rect 35530 2530 35590 2540
rect 35790 2580 35850 2590
rect 35790 2540 35800 2580
rect 35800 2540 35840 2580
rect 35840 2540 35850 2580
rect 35790 2530 35850 2540
rect 5970 2330 6030 2340
rect 5970 2290 5980 2330
rect 5980 2290 6020 2330
rect 6020 2290 6030 2330
rect 5970 2280 6030 2290
rect 10280 2330 10340 2340
rect 10280 2290 10290 2330
rect 10290 2290 10330 2330
rect 10330 2290 10340 2330
rect 10280 2280 10340 2290
rect 34670 2220 34730 2280
rect 34560 2130 34620 2190
rect 6900 2040 6960 2100
rect 8130 2040 8190 2100
rect 9360 2040 9420 2100
rect 6570 1950 6630 1960
rect 6570 1910 6580 1950
rect 6580 1910 6620 1950
rect 6620 1910 6630 1950
rect 6570 1900 6630 1910
rect 6790 1950 6850 1960
rect 6790 1910 6800 1950
rect 6800 1910 6840 1950
rect 6840 1910 6850 1950
rect 6790 1900 6850 1910
rect 7010 1950 7070 1960
rect 7010 1910 7020 1950
rect 7020 1910 7060 1950
rect 7060 1910 7070 1950
rect 7010 1900 7070 1910
rect 7800 1950 7860 1960
rect 7800 1910 7810 1950
rect 7810 1910 7850 1950
rect 7850 1910 7860 1950
rect 7800 1900 7860 1910
rect 8020 1950 8080 1960
rect 8020 1910 8030 1950
rect 8030 1910 8070 1950
rect 8070 1910 8080 1950
rect 8020 1900 8080 1910
rect 8240 1950 8300 1960
rect 8240 1910 8250 1950
rect 8250 1910 8290 1950
rect 8290 1910 8300 1950
rect 8240 1900 8300 1910
rect 8460 1950 8520 1960
rect 8460 1910 8470 1950
rect 8470 1910 8510 1950
rect 8510 1910 8520 1950
rect 8460 1900 8520 1910
rect 9250 1950 9310 1960
rect 9250 1910 9260 1950
rect 9260 1910 9300 1950
rect 9300 1910 9310 1950
rect 9250 1900 9310 1910
rect 9470 1950 9530 1960
rect 9470 1910 9480 1950
rect 9480 1910 9520 1950
rect 9520 1910 9530 1950
rect 9470 1900 9530 1910
rect 9690 1950 9750 1960
rect 9690 1910 9700 1950
rect 9700 1910 9740 1950
rect 9740 1910 9750 1950
rect 9690 1900 9750 1910
rect 7350 1780 7410 1790
rect 7350 1740 7360 1780
rect 7360 1740 7400 1780
rect 7400 1740 7410 1780
rect 7350 1730 7410 1740
rect 7460 1780 7520 1790
rect 7460 1740 7470 1780
rect 7470 1740 7510 1780
rect 7510 1740 7520 1780
rect 7460 1730 7520 1740
rect 8800 1780 8860 1790
rect 8800 1740 8810 1780
rect 8810 1740 8850 1780
rect 8850 1740 8860 1780
rect 8800 1730 8860 1740
rect 8910 1780 8970 1790
rect 8910 1740 8920 1780
rect 8920 1740 8960 1780
rect 8960 1740 8970 1780
rect 8910 1730 8970 1740
rect 10030 1780 10090 1790
rect 10030 1740 10040 1780
rect 10040 1740 10080 1780
rect 10080 1740 10090 1780
rect 10030 1730 10090 1740
rect 6460 1610 6520 1620
rect 6460 1570 6470 1610
rect 6470 1570 6510 1610
rect 6510 1570 6520 1610
rect 6460 1560 6520 1570
rect 6680 1610 6740 1620
rect 6680 1570 6690 1610
rect 6690 1570 6730 1610
rect 6730 1570 6740 1610
rect 6680 1560 6740 1570
rect 6900 1610 6960 1620
rect 6900 1570 6910 1610
rect 6910 1570 6950 1610
rect 6950 1570 6960 1610
rect 6900 1560 6960 1570
rect 7120 1610 7180 1620
rect 7120 1570 7130 1610
rect 7130 1570 7170 1610
rect 7170 1570 7180 1610
rect 7120 1560 7180 1570
rect 8130 1610 8190 1620
rect 8130 1570 8140 1610
rect 8140 1570 8180 1610
rect 8180 1570 8190 1610
rect 8130 1560 8190 1570
rect 8350 1610 8410 1620
rect 8350 1570 8360 1610
rect 8360 1570 8400 1610
rect 8400 1570 8410 1610
rect 8350 1560 8410 1570
rect 8570 1610 8630 1620
rect 8570 1570 8580 1610
rect 8580 1570 8620 1610
rect 8620 1570 8630 1610
rect 8570 1560 8630 1570
rect 9140 1610 9200 1620
rect 9140 1570 9150 1610
rect 9150 1570 9190 1610
rect 9190 1570 9200 1610
rect 9140 1560 9200 1570
rect 9580 1610 9640 1620
rect 9580 1570 9590 1610
rect 9590 1570 9630 1610
rect 9630 1570 9640 1610
rect 9580 1560 9640 1570
rect 5120 1360 5180 1420
rect 7740 1360 7800 1420
rect 9360 1450 9420 1510
rect 9800 1450 9860 1510
rect 34850 2330 34910 2390
rect 34760 1940 34820 2000
rect 34670 1030 34730 1090
rect 34940 1690 35000 1750
rect 35030 1230 35090 1290
rect 34850 700 34910 760
rect 34670 360 34730 420
rect 34560 -720 34620 -660
rect 36250 2530 36310 2590
rect 36130 2220 36190 2280
rect 35660 2130 35720 2190
rect 35230 2040 35290 2100
rect 35650 1810 35710 1870
rect 35890 1810 35950 1870
rect 36130 1810 36190 1870
rect 37770 2380 37830 2390
rect 37770 2340 37780 2380
rect 37780 2340 37820 2380
rect 37820 2340 37830 2380
rect 37770 2330 37830 2340
rect 38490 2380 38550 2390
rect 38490 2340 38500 2380
rect 38500 2340 38540 2380
rect 38540 2340 38550 2380
rect 38490 2330 38550 2340
rect 37410 2220 37470 2280
rect 37050 2130 37110 2190
rect 36690 2040 36750 2100
rect 36370 1810 36430 1870
rect 36610 1860 36670 1870
rect 36610 1820 36620 1860
rect 36620 1820 36660 1860
rect 36660 1820 36670 1860
rect 36610 1810 36670 1820
rect 36850 1810 36910 1870
rect 37090 1810 37150 1870
rect 37330 1810 37390 1870
rect 37570 1810 37630 1870
rect 38850 2220 38910 2280
rect 39210 2130 39270 2190
rect 39390 2130 39450 2190
rect 38130 2040 38190 2100
rect 39570 2040 39630 2100
rect 40130 3460 40190 3520
rect 40040 3350 40100 3410
rect 41240 3260 41300 3320
rect 40590 3040 40650 3050
rect 40590 3000 40600 3040
rect 40600 3000 40640 3040
rect 40640 3000 40650 3040
rect 40590 2990 40650 3000
rect 40590 2920 40650 2930
rect 40590 2880 40600 2920
rect 40600 2880 40640 2920
rect 40640 2880 40650 2920
rect 40590 2870 40650 2880
rect 40460 2580 40520 2590
rect 40460 2540 40470 2580
rect 40470 2540 40510 2580
rect 40510 2540 40520 2580
rect 40460 2530 40520 2540
rect 40720 2580 40780 2590
rect 40720 2540 40730 2580
rect 40730 2540 40770 2580
rect 40770 2540 40780 2580
rect 40720 2530 40780 2540
rect 40130 2240 40190 2300
rect 40040 2130 40100 2190
rect 41060 2240 41120 2300
rect 38570 1940 38630 2000
rect 39950 1940 40010 2000
rect 40590 1940 40650 2000
rect 38690 1860 38750 1870
rect 38690 1820 38700 1860
rect 38700 1820 38740 1860
rect 38740 1820 38750 1860
rect 38690 1810 38750 1820
rect 38930 1860 38990 1870
rect 38930 1820 38940 1860
rect 38940 1820 38980 1860
rect 38980 1820 38990 1860
rect 38930 1810 38990 1820
rect 39170 1860 39230 1870
rect 39170 1820 39180 1860
rect 39180 1820 39220 1860
rect 39220 1820 39230 1860
rect 39170 1810 39230 1820
rect 39410 1860 39470 1870
rect 39410 1820 39420 1860
rect 39420 1820 39460 1860
rect 39460 1820 39470 1860
rect 39410 1810 39470 1820
rect 39650 1860 39710 1870
rect 39650 1820 39660 1860
rect 39660 1820 39700 1860
rect 39700 1820 39710 1860
rect 39650 1810 39710 1820
rect 39890 1860 39950 1870
rect 39890 1820 39900 1860
rect 39900 1820 39940 1860
rect 39940 1820 39950 1860
rect 39890 1810 39950 1820
rect 40130 1860 40190 1870
rect 40130 1820 40140 1860
rect 40140 1820 40180 1860
rect 40180 1820 40190 1860
rect 40130 1810 40190 1820
rect 40370 1860 40430 1870
rect 40370 1820 40380 1860
rect 40380 1820 40420 1860
rect 40420 1820 40430 1860
rect 40370 1810 40430 1820
rect 40610 1860 40670 1870
rect 40610 1820 40620 1860
rect 40620 1820 40660 1860
rect 40660 1820 40670 1860
rect 40610 1810 40670 1820
rect 35530 1740 35590 1750
rect 35530 1700 35540 1740
rect 35540 1700 35580 1740
rect 35580 1700 35590 1740
rect 35530 1690 35590 1700
rect 36250 1740 36310 1750
rect 36250 1700 36260 1740
rect 36260 1700 36300 1740
rect 36300 1700 36310 1740
rect 36250 1690 36310 1700
rect 36970 1740 37030 1750
rect 36970 1700 36980 1740
rect 36980 1700 37020 1740
rect 37020 1700 37030 1740
rect 36970 1690 37030 1700
rect 37690 1740 37750 1750
rect 37690 1700 37700 1740
rect 37700 1700 37740 1740
rect 37740 1700 37750 1740
rect 37690 1690 37750 1700
rect 37950 1690 38010 1750
rect 38310 1690 38370 1750
rect 38570 1740 38630 1750
rect 38570 1700 38580 1740
rect 38580 1700 38620 1740
rect 38620 1700 38630 1740
rect 38570 1690 38630 1700
rect 39290 1740 39350 1750
rect 39290 1700 39300 1740
rect 39300 1700 39340 1740
rect 39340 1700 39350 1740
rect 39290 1690 39350 1700
rect 40010 1740 40070 1750
rect 40010 1700 40020 1740
rect 40020 1700 40060 1740
rect 40060 1700 40070 1740
rect 40010 1690 40070 1700
rect 40730 1740 40790 1750
rect 40730 1700 40740 1740
rect 40740 1700 40780 1740
rect 40780 1700 40790 1740
rect 40730 1690 40790 1700
rect 35770 1400 35830 1410
rect 35770 1360 35780 1400
rect 35780 1360 35820 1400
rect 35820 1360 35830 1400
rect 35770 1350 35830 1360
rect 36490 1400 36550 1410
rect 36490 1360 36500 1400
rect 36500 1360 36540 1400
rect 36540 1360 36550 1400
rect 36490 1350 36550 1360
rect 37210 1400 37270 1410
rect 37210 1360 37220 1400
rect 37220 1360 37260 1400
rect 37260 1360 37270 1400
rect 37210 1350 37270 1360
rect 35590 1230 35650 1290
rect 36010 1230 36070 1290
rect 36250 1230 36310 1290
rect 36730 1230 36790 1290
rect 36970 1230 37030 1290
rect 37450 1230 37510 1290
rect 37630 1230 37690 1290
rect 36390 1080 36450 1090
rect 36390 1040 36400 1080
rect 36400 1040 36440 1080
rect 36440 1040 36450 1080
rect 36390 1030 36450 1040
rect 36510 1060 36570 1120
rect 36990 1060 37050 1120
rect 37470 1060 37530 1120
rect 36270 990 36330 1000
rect 36270 950 36280 990
rect 36280 950 36320 990
rect 36320 950 36330 990
rect 36270 940 36330 950
rect 36750 990 36810 1000
rect 36750 950 36760 990
rect 36760 950 36800 990
rect 36800 950 36810 990
rect 36750 940 36810 950
rect 37230 990 37290 1000
rect 37230 950 37240 990
rect 37240 950 37280 990
rect 37280 950 37290 990
rect 37230 940 37290 950
rect 37590 870 37650 880
rect 37590 830 37600 870
rect 37600 830 37640 870
rect 37640 830 37650 870
rect 37590 820 37650 830
rect 36270 750 36330 760
rect 36270 710 36280 750
rect 36280 710 36320 750
rect 36320 710 36330 750
rect 36270 700 36330 710
rect 35790 580 35850 640
rect 36390 580 36450 640
rect 36630 580 36690 640
rect 36870 580 36930 640
rect 37110 580 37170 640
rect 37350 580 37410 640
rect 35970 430 36030 440
rect 35970 390 35980 430
rect 35980 390 36020 430
rect 36020 390 36030 430
rect 35970 380 36030 390
rect 36210 430 36270 440
rect 36210 390 36220 430
rect 36220 390 36260 430
rect 36260 390 36270 430
rect 36210 380 36270 390
rect 36450 430 36510 440
rect 36450 390 36460 430
rect 36460 390 36500 430
rect 36500 390 36510 430
rect 36450 380 36510 390
rect 36690 430 36750 440
rect 36690 390 36700 430
rect 36700 390 36740 430
rect 36740 390 36750 430
rect 36690 380 36750 390
rect 37170 430 37230 440
rect 37170 390 37180 430
rect 37180 390 37220 430
rect 37220 390 37230 430
rect 37170 380 37230 390
rect 37410 430 37470 440
rect 37410 390 37420 430
rect 37420 390 37460 430
rect 37460 390 37470 430
rect 37410 380 37470 390
rect 37650 430 37710 440
rect 37650 390 37660 430
rect 37660 390 37700 430
rect 37700 390 37710 430
rect 37650 380 37710 390
rect 38130 820 38190 880
rect 39050 1400 39110 1410
rect 39050 1360 39060 1400
rect 39060 1360 39100 1400
rect 39100 1360 39110 1400
rect 39050 1350 39110 1360
rect 39770 1400 39830 1410
rect 39770 1360 39780 1400
rect 39780 1360 39820 1400
rect 39820 1360 39830 1400
rect 39770 1350 39830 1360
rect 40490 1400 40550 1410
rect 40490 1360 40500 1400
rect 40500 1360 40540 1400
rect 40540 1360 40550 1400
rect 40490 1350 40550 1360
rect 38630 1230 38690 1290
rect 38810 1230 38870 1290
rect 39290 1230 39350 1290
rect 39530 1230 39590 1290
rect 38790 1060 38850 1120
rect 39270 1060 39330 1120
rect 41150 2040 41210 2100
rect 40010 1230 40070 1290
rect 40250 1230 40310 1290
rect 40670 1230 40730 1290
rect 41060 1230 41120 1290
rect 39750 1060 39810 1120
rect 39870 1080 39930 1090
rect 39870 1040 39880 1080
rect 39880 1040 39920 1080
rect 39920 1040 39930 1080
rect 39870 1030 39930 1040
rect 41150 1030 41210 1090
rect 39030 990 39090 1000
rect 39030 950 39040 990
rect 39040 950 39080 990
rect 39080 950 39090 990
rect 39030 940 39090 950
rect 39510 990 39570 1000
rect 39510 950 39520 990
rect 39520 950 39560 990
rect 39560 950 39570 990
rect 39510 940 39570 950
rect 39990 990 40050 1000
rect 39990 950 40000 990
rect 40000 950 40040 990
rect 40040 950 40050 990
rect 39990 940 40050 950
rect 38670 870 38730 880
rect 38670 830 38680 870
rect 38680 830 38720 870
rect 38720 830 38730 870
rect 38670 820 38730 830
rect 39990 750 40050 760
rect 39990 710 40000 750
rect 40000 710 40040 750
rect 40040 710 40050 750
rect 39990 700 40050 710
rect 41240 700 41300 760
rect 38910 580 38970 640
rect 39150 580 39210 640
rect 39390 580 39450 640
rect 39630 580 39690 640
rect 39870 580 39930 640
rect 40470 580 40530 640
rect 38610 430 38670 440
rect 38610 390 38620 430
rect 38620 390 38660 430
rect 38660 390 38670 430
rect 38610 380 38670 390
rect 38850 430 38910 440
rect 38850 390 38860 430
rect 38860 390 38900 430
rect 38900 390 38910 430
rect 38850 380 38910 390
rect 39090 430 39150 440
rect 39090 390 39100 430
rect 39100 390 39140 430
rect 39140 390 39150 430
rect 39090 380 39150 390
rect 39570 430 39630 440
rect 39570 390 39580 430
rect 39580 390 39620 430
rect 39620 390 39630 430
rect 39570 380 39630 390
rect 39810 430 39870 440
rect 39810 390 39820 430
rect 39820 390 39860 430
rect 39860 390 39870 430
rect 39810 380 39870 390
rect 40050 430 40110 440
rect 40050 390 40060 430
rect 40060 390 40100 430
rect 40100 390 40110 430
rect 40050 380 40110 390
rect 40290 430 40350 440
rect 40290 390 40300 430
rect 40300 390 40340 430
rect 40340 390 40350 430
rect 40290 380 40350 390
rect 36870 -200 36930 -190
rect 36870 -240 36880 -200
rect 36880 -240 36920 -200
rect 36920 -240 36930 -200
rect 36870 -250 36930 -240
rect 38130 -250 38190 -190
rect 39390 -200 39450 -190
rect 39390 -240 39400 -200
rect 39400 -240 39440 -200
rect 39440 -240 39450 -200
rect 39390 -250 39450 -240
rect 38130 -400 38190 -380
rect 38130 -440 38140 -400
rect 38140 -440 38180 -400
rect 38180 -440 38190 -400
rect 36050 -500 36110 -490
rect 36050 -540 36060 -500
rect 36060 -540 36100 -500
rect 36100 -540 36110 -500
rect 36050 -550 36110 -540
rect 36210 -500 36270 -490
rect 36210 -540 36220 -500
rect 36220 -540 36260 -500
rect 36260 -540 36270 -500
rect 36210 -550 36270 -540
rect 36370 -500 36430 -490
rect 36370 -540 36380 -500
rect 36380 -540 36420 -500
rect 36420 -540 36430 -500
rect 36370 -550 36430 -540
rect 36530 -500 36590 -490
rect 36530 -540 36540 -500
rect 36540 -540 36580 -500
rect 36580 -540 36590 -500
rect 36530 -550 36590 -540
rect 36690 -500 36750 -490
rect 36690 -540 36700 -500
rect 36700 -540 36740 -500
rect 36740 -540 36750 -500
rect 36690 -550 36750 -540
rect 36850 -500 36910 -490
rect 36850 -540 36860 -500
rect 36860 -540 36900 -500
rect 36900 -540 36910 -500
rect 36850 -550 36910 -540
rect 37010 -500 37070 -490
rect 37010 -540 37020 -500
rect 37020 -540 37060 -500
rect 37060 -540 37070 -500
rect 37010 -550 37070 -540
rect 37170 -500 37230 -490
rect 37170 -540 37180 -500
rect 37180 -540 37220 -500
rect 37220 -540 37230 -500
rect 37170 -550 37230 -540
rect 37330 -500 37390 -490
rect 37330 -540 37340 -500
rect 37340 -540 37380 -500
rect 37380 -540 37390 -500
rect 37330 -550 37390 -540
rect 37490 -500 37550 -490
rect 37490 -540 37500 -500
rect 37500 -540 37540 -500
rect 37540 -540 37550 -500
rect 37490 -550 37550 -540
rect 37650 -500 37710 -490
rect 37650 -540 37660 -500
rect 37660 -540 37700 -500
rect 37700 -540 37710 -500
rect 37650 -550 37710 -540
rect 37810 -500 37870 -490
rect 37810 -540 37820 -500
rect 37820 -540 37860 -500
rect 37860 -540 37870 -500
rect 37810 -550 37870 -540
rect 37970 -500 38030 -490
rect 37970 -540 37980 -500
rect 37980 -540 38020 -500
rect 38020 -540 38030 -500
rect 37970 -550 38030 -540
rect 38130 -500 38190 -490
rect 38130 -540 38140 -500
rect 38140 -540 38180 -500
rect 38180 -540 38190 -500
rect 38130 -550 38190 -540
rect 38290 -500 38350 -490
rect 38290 -540 38300 -500
rect 38300 -540 38340 -500
rect 38340 -540 38350 -500
rect 38290 -550 38350 -540
rect 38450 -500 38510 -490
rect 38450 -540 38460 -500
rect 38460 -540 38500 -500
rect 38500 -540 38510 -500
rect 38450 -550 38510 -540
rect 38610 -500 38670 -490
rect 38610 -540 38620 -500
rect 38620 -540 38660 -500
rect 38660 -540 38670 -500
rect 38610 -550 38670 -540
rect 38770 -500 38830 -490
rect 38770 -540 38780 -500
rect 38780 -540 38820 -500
rect 38820 -540 38830 -500
rect 38770 -550 38830 -540
rect 38930 -500 38990 -490
rect 38930 -540 38940 -500
rect 38940 -540 38980 -500
rect 38980 -540 38990 -500
rect 38930 -550 38990 -540
rect 39090 -500 39150 -490
rect 39090 -540 39100 -500
rect 39100 -540 39140 -500
rect 39140 -540 39150 -500
rect 39090 -550 39150 -540
rect 39250 -500 39310 -490
rect 39250 -540 39260 -500
rect 39260 -540 39300 -500
rect 39300 -540 39310 -500
rect 39250 -550 39310 -540
rect 39410 -500 39470 -490
rect 39410 -540 39420 -500
rect 39420 -540 39460 -500
rect 39460 -540 39470 -500
rect 39410 -550 39470 -540
rect 39570 -500 39630 -490
rect 39570 -540 39580 -500
rect 39580 -540 39620 -500
rect 39620 -540 39630 -500
rect 39570 -550 39630 -540
rect 39730 -500 39790 -490
rect 39730 -540 39740 -500
rect 39740 -540 39780 -500
rect 39780 -540 39790 -500
rect 39730 -550 39790 -540
rect 39890 -500 39950 -490
rect 39890 -540 39900 -500
rect 39900 -540 39940 -500
rect 39940 -540 39950 -500
rect 39890 -550 39950 -540
rect 40050 -500 40110 -490
rect 40050 -540 40060 -500
rect 40060 -540 40100 -500
rect 40100 -540 40110 -500
rect 40050 -550 40110 -540
rect 35970 -670 36030 -660
rect 35970 -710 35980 -670
rect 35980 -710 36020 -670
rect 36020 -710 36030 -670
rect 35970 -720 36030 -710
rect 40280 -670 40340 -660
rect 40280 -710 40290 -670
rect 40290 -710 40330 -670
rect 40330 -710 40340 -670
rect 40280 -720 40340 -710
rect 36900 -960 36960 -900
rect 38130 -960 38190 -900
rect 39360 -960 39420 -900
rect 36570 -1050 36630 -1040
rect 36570 -1090 36580 -1050
rect 36580 -1090 36620 -1050
rect 36620 -1090 36630 -1050
rect 36570 -1100 36630 -1090
rect 36790 -1050 36850 -1040
rect 36790 -1090 36800 -1050
rect 36800 -1090 36840 -1050
rect 36840 -1090 36850 -1050
rect 36790 -1100 36850 -1090
rect 37010 -1050 37070 -1040
rect 37010 -1090 37020 -1050
rect 37020 -1090 37060 -1050
rect 37060 -1090 37070 -1050
rect 37010 -1100 37070 -1090
rect 37800 -1050 37860 -1040
rect 37800 -1090 37810 -1050
rect 37810 -1090 37850 -1050
rect 37850 -1090 37860 -1050
rect 37800 -1100 37860 -1090
rect 38020 -1050 38080 -1040
rect 38020 -1090 38030 -1050
rect 38030 -1090 38070 -1050
rect 38070 -1090 38080 -1050
rect 38020 -1100 38080 -1090
rect 38240 -1050 38300 -1040
rect 38240 -1090 38250 -1050
rect 38250 -1090 38290 -1050
rect 38290 -1090 38300 -1050
rect 38240 -1100 38300 -1090
rect 38460 -1050 38520 -1040
rect 38460 -1090 38470 -1050
rect 38470 -1090 38510 -1050
rect 38510 -1090 38520 -1050
rect 38460 -1100 38520 -1090
rect 39250 -1050 39310 -1040
rect 39250 -1090 39260 -1050
rect 39260 -1090 39300 -1050
rect 39300 -1090 39310 -1050
rect 39250 -1100 39310 -1090
rect 39470 -1050 39530 -1040
rect 39470 -1090 39480 -1050
rect 39480 -1090 39520 -1050
rect 39520 -1090 39530 -1050
rect 39470 -1100 39530 -1090
rect 39690 -1050 39750 -1040
rect 39690 -1090 39700 -1050
rect 39700 -1090 39740 -1050
rect 39740 -1090 39750 -1050
rect 39690 -1100 39750 -1090
rect 37350 -1220 37410 -1210
rect 37350 -1260 37360 -1220
rect 37360 -1260 37400 -1220
rect 37400 -1260 37410 -1220
rect 37350 -1270 37410 -1260
rect 37460 -1220 37520 -1210
rect 37460 -1260 37470 -1220
rect 37470 -1260 37510 -1220
rect 37510 -1260 37520 -1220
rect 37460 -1270 37520 -1260
rect 38800 -1220 38860 -1210
rect 38800 -1260 38810 -1220
rect 38810 -1260 38850 -1220
rect 38850 -1260 38860 -1220
rect 38800 -1270 38860 -1260
rect 38910 -1220 38970 -1210
rect 38910 -1260 38920 -1220
rect 38920 -1260 38960 -1220
rect 38960 -1260 38970 -1220
rect 38910 -1270 38970 -1260
rect 40030 -1220 40090 -1210
rect 40030 -1260 40040 -1220
rect 40040 -1260 40080 -1220
rect 40080 -1260 40090 -1220
rect 40030 -1270 40090 -1260
rect 36460 -1390 36520 -1380
rect 36460 -1430 36470 -1390
rect 36470 -1430 36510 -1390
rect 36510 -1430 36520 -1390
rect 36460 -1440 36520 -1430
rect 36680 -1390 36740 -1380
rect 36680 -1430 36690 -1390
rect 36690 -1430 36730 -1390
rect 36730 -1430 36740 -1390
rect 36680 -1440 36740 -1430
rect 36900 -1390 36960 -1380
rect 36900 -1430 36910 -1390
rect 36910 -1430 36950 -1390
rect 36950 -1430 36960 -1390
rect 36900 -1440 36960 -1430
rect 37120 -1390 37180 -1380
rect 37120 -1430 37130 -1390
rect 37130 -1430 37170 -1390
rect 37170 -1430 37180 -1390
rect 37120 -1440 37180 -1430
rect 38130 -1390 38190 -1380
rect 38130 -1430 38140 -1390
rect 38140 -1430 38180 -1390
rect 38180 -1430 38190 -1390
rect 38130 -1440 38190 -1430
rect 38350 -1390 38410 -1380
rect 38350 -1430 38360 -1390
rect 38360 -1430 38400 -1390
rect 38400 -1430 38410 -1390
rect 38350 -1440 38410 -1430
rect 38570 -1390 38630 -1380
rect 38570 -1430 38580 -1390
rect 38580 -1430 38620 -1390
rect 38620 -1430 38630 -1390
rect 38570 -1440 38630 -1430
rect 39140 -1390 39200 -1380
rect 39140 -1430 39150 -1390
rect 39150 -1430 39190 -1390
rect 39190 -1430 39200 -1390
rect 39140 -1440 39200 -1430
rect 39580 -1390 39640 -1380
rect 39580 -1430 39590 -1390
rect 39590 -1430 39630 -1390
rect 39630 -1430 39640 -1390
rect 39580 -1440 39640 -1430
rect 35120 -1640 35180 -1580
rect 37740 -1640 37800 -1580
rect 39360 -1550 39420 -1490
rect 39800 -1550 39860 -1490
rect 43890 -3950 43950 -3890
rect 46520 -2680 46580 -2620
rect 44150 -2780 44210 -2720
rect 44142 -2830 44212 -2820
rect 44142 -2880 44152 -2830
rect 44152 -2880 44202 -2830
rect 44202 -2880 44212 -2830
rect 44142 -2890 44212 -2880
rect 44142 -2950 44212 -2940
rect 44142 -3000 44152 -2950
rect 44152 -3000 44202 -2950
rect 44202 -3000 44212 -2950
rect 44142 -3010 44212 -3000
rect 46712 -3100 46782 -3090
rect 46712 -3150 46722 -3100
rect 46722 -3150 46772 -3100
rect 46772 -3150 46782 -3100
rect 46712 -3160 46782 -3150
rect 44150 -3310 44210 -3250
rect 46520 -3310 46580 -3250
rect 46712 -3220 46782 -3210
rect 46712 -3270 46722 -3220
rect 46722 -3270 46772 -3220
rect 46772 -3270 46782 -3220
rect 46712 -3280 46782 -3270
rect 44142 -3360 44212 -3350
rect 44142 -3410 44152 -3360
rect 44152 -3410 44202 -3360
rect 44202 -3410 44212 -3360
rect 44142 -3420 44212 -3410
rect 44142 -3480 44212 -3470
rect 44142 -3530 44152 -3480
rect 44152 -3530 44202 -3480
rect 44202 -3530 44212 -3480
rect 44142 -3540 44212 -3530
rect 46380 -3430 46440 -3420
rect 46380 -3470 46390 -3430
rect 46390 -3470 46430 -3430
rect 46430 -3470 46440 -3430
rect 46380 -3480 46440 -3470
rect 46590 -3430 46650 -3420
rect 46590 -3470 46600 -3430
rect 46600 -3470 46640 -3430
rect 46640 -3470 46650 -3430
rect 46590 -3480 46650 -3470
rect 45200 -3620 45260 -3610
rect 45200 -3660 45210 -3620
rect 45210 -3660 45250 -3620
rect 45250 -3660 45260 -3620
rect 45200 -3670 45260 -3660
rect 48850 -3580 48920 -3570
rect 48850 -3630 48860 -3580
rect 48860 -3630 48910 -3580
rect 48910 -3630 48920 -3580
rect 48850 -3640 48920 -3630
rect 48850 -3700 48920 -3690
rect 48850 -3750 48860 -3700
rect 48860 -3750 48910 -3700
rect 48910 -3750 48920 -3700
rect 48850 -3760 48920 -3750
rect 44532 -3890 44602 -3880
rect 44532 -3940 44542 -3890
rect 44542 -3940 44592 -3890
rect 44592 -3940 44602 -3890
rect 44532 -3950 44602 -3940
rect 45878 -3890 45948 -3880
rect 45878 -3940 45888 -3890
rect 45888 -3940 45938 -3890
rect 45938 -3940 45948 -3890
rect 45878 -3950 45948 -3940
rect 46430 -3950 46490 -3890
rect 46220 -4160 46280 -4100
rect 43980 -4360 44040 -4300
rect 44532 -4310 44602 -4300
rect 44532 -4360 44542 -4310
rect 44542 -4360 44592 -4310
rect 44592 -4360 44602 -4310
rect 44532 -4370 44602 -4360
rect 45878 -4310 45948 -4300
rect 45878 -4360 45888 -4310
rect 45888 -4360 45938 -4310
rect 45938 -4360 45948 -4310
rect 45878 -4370 45948 -4360
rect 47042 -4110 47112 -4100
rect 47042 -4160 47052 -4110
rect 47052 -4160 47102 -4110
rect 47102 -4160 47112 -4110
rect 47042 -4170 47112 -4160
rect 48440 -4110 48510 -4100
rect 48440 -4160 48450 -4110
rect 48450 -4160 48500 -4110
rect 48500 -4160 48510 -4110
rect 48440 -4170 48510 -4160
rect 48850 -4170 48910 -4110
rect 46430 -4460 46490 -4400
rect 48760 -4460 48820 -4400
rect 48940 -4370 49000 -4310
rect 49120 -2780 49180 -2720
rect 49120 -3550 49180 -3490
rect 49230 -3550 49250 -3490
rect 49120 -3730 49180 -3670
rect 29790 -6620 29850 -6560
rect 35590 -5970 35650 -5916
rect 35570 -8540 35630 -8530
rect 35570 -8580 35580 -8540
rect 35580 -8580 35620 -8540
rect 35620 -8580 35630 -8540
rect 35570 -8590 35630 -8580
<< metal2 >>
rect -220 7750 -140 7760
rect -220 7690 -210 7750
rect -150 7740 -140 7750
rect 2700 7750 2780 7760
rect 2700 7740 2710 7750
rect -150 7700 2710 7740
rect -150 7690 -140 7700
rect -220 7680 -140 7690
rect 2700 7690 2710 7700
rect 2770 7690 2780 7750
rect 29780 7750 29860 7760
rect 2700 7680 2780 7690
rect 8880 7690 8960 7700
rect 8880 7630 8890 7690
rect 8950 7680 8960 7690
rect 11500 7690 11580 7700
rect 11500 7680 11510 7690
rect 8950 7640 11510 7680
rect 8950 7630 8960 7640
rect 8880 7620 8960 7630
rect 11500 7630 11510 7640
rect 11570 7630 11580 7690
rect 29780 7690 29790 7750
rect 29850 7740 29860 7750
rect 32700 7750 32780 7760
rect 32700 7740 32710 7750
rect 29850 7700 32710 7740
rect 29850 7690 29860 7700
rect 29780 7680 29860 7690
rect 32700 7690 32710 7700
rect 32770 7690 32780 7750
rect 32700 7680 32780 7690
rect 38880 7690 38960 7700
rect 11500 7620 11580 7630
rect 38880 7630 38890 7690
rect 38950 7680 38960 7690
rect 41500 7690 41580 7700
rect 41500 7680 41510 7690
rect 38950 7640 41510 7680
rect 38950 7630 38960 7640
rect 38880 7620 38960 7630
rect 41500 7630 41510 7640
rect 41570 7630 41580 7690
rect 41500 7620 41580 7630
rect -30 7590 50 7600
rect -30 7530 -20 7590
rect 40 7580 50 7590
rect 1880 7590 1960 7600
rect 1880 7580 1890 7590
rect 40 7540 1890 7580
rect 40 7530 50 7540
rect -30 7520 50 7530
rect 1880 7530 1890 7540
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect 3270 7590 3370 7610
rect 5020 7600 5100 7610
rect 5020 7590 5030 7600
rect 3270 7530 3290 7590
rect 3350 7550 5030 7590
rect 3350 7530 3370 7550
rect 5020 7540 5030 7550
rect 5090 7540 5100 7600
rect 5020 7530 5100 7540
rect 9310 7590 9390 7600
rect 9310 7530 9320 7590
rect 9380 7580 9390 7590
rect 10270 7590 10370 7610
rect 10270 7580 10290 7590
rect 9380 7540 10290 7580
rect 9380 7530 9390 7540
rect 3270 7510 3370 7530
rect 9310 7520 9390 7530
rect 10270 7530 10290 7540
rect 10350 7530 10370 7590
rect 10270 7510 10370 7530
rect 29970 7590 30050 7600
rect 29970 7530 29980 7590
rect 30040 7580 30050 7590
rect 31880 7590 31960 7600
rect 31880 7580 31890 7590
rect 30040 7540 31890 7580
rect 30040 7530 30050 7540
rect 29970 7520 30050 7530
rect 31880 7530 31890 7540
rect 31950 7530 31960 7590
rect 31880 7520 31960 7530
rect 33270 7590 33370 7610
rect 35020 7600 35100 7610
rect 35020 7590 35030 7600
rect 33270 7530 33290 7590
rect 33350 7550 35030 7590
rect 33350 7530 33370 7550
rect 35020 7540 35030 7550
rect 35090 7540 35100 7600
rect 35020 7530 35100 7540
rect 39310 7590 39390 7600
rect 39310 7530 39320 7590
rect 39380 7580 39390 7590
rect 40270 7590 40370 7610
rect 40270 7580 40290 7590
rect 39380 7540 40290 7580
rect 39380 7530 39390 7540
rect 33270 7510 33370 7530
rect 39310 7520 39390 7530
rect 40270 7530 40290 7540
rect 40350 7530 40370 7590
rect 40270 7510 40370 7530
rect -120 7480 -40 7490
rect -120 7420 -110 7480
rect -50 7470 -40 7480
rect 5380 7480 5460 7490
rect 5380 7470 5390 7480
rect -50 7430 5390 7470
rect -50 7420 -40 7430
rect -120 7410 -40 7420
rect 5380 7420 5390 7430
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7480 6870 7500
rect 6770 7420 6790 7480
rect 6850 7470 6870 7480
rect 9220 7480 9300 7490
rect 9220 7470 9230 7480
rect 6850 7430 9230 7470
rect 6850 7420 6870 7430
rect 6770 7400 6870 7420
rect 9220 7420 9230 7430
rect 9290 7420 9300 7480
rect 9220 7410 9300 7420
rect 29880 7480 29960 7490
rect 29880 7420 29890 7480
rect 29950 7470 29960 7480
rect 35380 7480 35460 7490
rect 35380 7470 35390 7480
rect 29950 7430 35390 7470
rect 29950 7420 29960 7430
rect 29880 7410 29960 7420
rect 35380 7420 35390 7430
rect 35450 7420 35460 7480
rect 35380 7410 35460 7420
rect 36770 7480 36870 7500
rect 36770 7420 36790 7480
rect 36850 7470 36870 7480
rect 39220 7480 39300 7490
rect 39220 7470 39230 7480
rect 36850 7430 39230 7470
rect 36850 7420 36870 7430
rect 36770 7400 36870 7420
rect 39220 7420 39230 7430
rect 39290 7420 39300 7480
rect 39220 7410 39300 7420
rect 2510 7380 2590 7390
rect 2510 7320 2520 7380
rect 2580 7370 2590 7380
rect 8560 7380 8640 7390
rect 8560 7370 8570 7380
rect 2580 7330 8570 7370
rect 2580 7320 2590 7330
rect 2510 7310 2590 7320
rect 8560 7320 8570 7330
rect 8630 7320 8640 7380
rect 38560 7380 38640 7390
rect 38560 7370 38570 7380
rect 35250 7330 38570 7370
rect 8560 7310 8640 7320
rect 38560 7320 38570 7330
rect 38630 7320 38640 7380
rect 38560 7310 38640 7320
rect 140 7280 220 7290
rect 140 7220 150 7280
rect 210 7270 220 7280
rect 5110 7280 5190 7290
rect 5110 7270 5120 7280
rect 210 7230 5120 7270
rect 210 7220 220 7230
rect 140 7210 220 7220
rect 5110 7220 5120 7230
rect 5180 7220 5190 7280
rect 5110 7210 5190 7220
rect 6620 7270 6700 7280
rect 6620 7210 6630 7270
rect 6690 7260 6700 7270
rect 6690 7220 12200 7260
rect 6690 7210 6700 7220
rect 6620 7200 6700 7210
rect 6400 7180 6480 7190
rect 132 7110 142 7180
rect 212 7110 222 7180
rect 6400 7120 6410 7180
rect 6470 7170 6480 7180
rect 8120 7180 8200 7190
rect 8120 7170 8130 7180
rect 6470 7130 8130 7170
rect 6470 7120 6480 7130
rect 6400 7110 6480 7120
rect 8120 7120 8130 7130
rect 8190 7170 8200 7180
rect 9130 7180 9210 7190
rect 9130 7170 9140 7180
rect 8190 7130 9140 7170
rect 8190 7120 8200 7130
rect 8120 7110 8200 7120
rect 9130 7120 9140 7130
rect 9200 7170 9210 7180
rect 9840 7180 9920 7190
rect 9840 7170 9850 7180
rect 9200 7130 9850 7170
rect 9200 7120 9210 7130
rect 9130 7110 9210 7120
rect 9840 7120 9850 7130
rect 9910 7120 9920 7180
rect 9840 7110 9920 7120
rect 6070 7060 6150 7070
rect -220 7050 -140 7060
rect -220 6990 -210 7050
rect -150 7040 -140 7050
rect 132 7040 142 7060
rect -150 7000 142 7040
rect -150 6990 -140 7000
rect 132 6990 142 7000
rect 212 6990 222 7060
rect 6070 7000 6080 7060
rect 6140 7050 6150 7060
rect 6290 7060 6370 7070
rect 6290 7050 6300 7060
rect 6140 7010 6300 7050
rect 6140 7000 6150 7010
rect 6070 6990 6150 7000
rect 6290 7000 6300 7010
rect 6360 7050 6370 7060
rect 6510 7060 6590 7070
rect 6510 7050 6520 7060
rect 6360 7010 6520 7050
rect 6360 7000 6370 7010
rect 6290 6990 6370 7000
rect 6510 7000 6520 7010
rect 6580 7050 6590 7060
rect 6730 7060 6810 7070
rect 6730 7050 6740 7060
rect 6580 7010 6740 7050
rect 6580 7000 6590 7010
rect 6510 6990 6590 7000
rect 6730 7000 6740 7010
rect 6800 7050 6810 7060
rect 7350 7060 7430 7070
rect 7350 7050 7360 7060
rect 6800 7010 7360 7050
rect 6800 7000 6810 7010
rect 6730 6990 6810 7000
rect 7350 7000 7360 7010
rect 7420 7050 7430 7060
rect 7570 7060 7650 7070
rect 7570 7050 7580 7060
rect 7420 7010 7580 7050
rect 7420 7000 7430 7010
rect 7350 6990 7430 7000
rect 7570 7000 7580 7010
rect 7640 7050 7650 7060
rect 7790 7060 7870 7070
rect 7790 7050 7800 7060
rect 7640 7010 7800 7050
rect 7640 7000 7650 7010
rect 7570 6990 7650 7000
rect 7790 7000 7800 7010
rect 7860 7050 7870 7060
rect 8010 7060 8090 7070
rect 8010 7050 8020 7060
rect 7860 7010 8020 7050
rect 7860 7000 7870 7010
rect 7790 6990 7870 7000
rect 8010 7000 8020 7010
rect 8080 7050 8090 7060
rect 8230 7060 8310 7070
rect 8230 7050 8240 7060
rect 8080 7010 8240 7050
rect 8080 7000 8090 7010
rect 8010 6990 8090 7000
rect 8230 7000 8240 7010
rect 8300 7050 8310 7060
rect 8450 7060 8530 7070
rect 8450 7050 8460 7060
rect 8300 7010 8460 7050
rect 8300 7000 8310 7010
rect 8230 6990 8310 7000
rect 8450 7000 8460 7010
rect 8520 7050 8530 7060
rect 8670 7060 8750 7070
rect 8670 7050 8680 7060
rect 8520 7010 8680 7050
rect 8520 7000 8530 7010
rect 8450 6990 8530 7000
rect 8670 7000 8680 7010
rect 8740 7050 8750 7060
rect 9510 7060 9590 7070
rect 9510 7050 9520 7060
rect 8740 7010 9520 7050
rect 8740 7000 8750 7010
rect 8670 6990 8750 7000
rect 9510 7000 9520 7010
rect 9580 7050 9590 7060
rect 9730 7060 9810 7070
rect 9730 7050 9740 7060
rect 9580 7010 9740 7050
rect 9580 7000 9590 7010
rect 9510 6990 9590 7000
rect 9730 7000 9740 7010
rect 9800 7050 9810 7060
rect 9950 7060 10030 7070
rect 9950 7050 9960 7060
rect 9800 7010 9960 7050
rect 9800 7000 9810 7010
rect 9730 6990 9810 7000
rect 9950 7000 9960 7010
rect 10020 7050 10030 7060
rect 10170 7060 10250 7070
rect 10170 7050 10180 7060
rect 10020 7010 10180 7050
rect 10020 7000 10030 7010
rect 9950 6990 10030 7000
rect 10170 7000 10180 7010
rect 10240 7050 10250 7060
rect 11500 7060 11580 7070
rect 11500 7050 11510 7060
rect 10240 7010 11510 7050
rect 10240 7000 10250 7010
rect 10170 6990 10250 7000
rect 11500 7000 11510 7010
rect 11570 7000 11580 7060
rect 11500 6990 11580 7000
rect -220 6980 -140 6990
rect 2702 6840 2712 6910
rect 2782 6840 2792 6910
rect 140 6750 220 6760
rect 140 6690 150 6750
rect 210 6740 220 6750
rect 2510 6750 2590 6760
rect 2510 6740 2520 6750
rect 210 6700 2520 6740
rect 210 6690 220 6700
rect 140 6680 220 6690
rect 2510 6690 2520 6700
rect 2580 6690 2590 6750
rect 2702 6720 2712 6790
rect 2782 6720 2792 6790
rect 6180 6720 6260 6730
rect 2510 6680 2590 6690
rect 6180 6660 6190 6720
rect 6250 6710 6260 6720
rect 6400 6720 6480 6730
rect 6400 6710 6410 6720
rect 6250 6670 6410 6710
rect 6250 6660 6260 6670
rect 6180 6650 6260 6660
rect 6400 6660 6410 6670
rect 6470 6710 6480 6720
rect 6620 6720 6700 6730
rect 6620 6710 6630 6720
rect 6470 6670 6630 6710
rect 6470 6660 6480 6670
rect 6400 6650 6480 6660
rect 6620 6660 6630 6670
rect 6690 6660 6700 6720
rect 6620 6650 6700 6660
rect 7680 6720 7760 6730
rect 7680 6660 7690 6720
rect 7750 6710 7760 6720
rect 7900 6720 7980 6730
rect 7900 6710 7910 6720
rect 7750 6670 7910 6710
rect 7750 6660 7760 6670
rect 7680 6650 7760 6660
rect 7900 6660 7910 6670
rect 7970 6710 7980 6720
rect 8120 6720 8200 6730
rect 8120 6710 8130 6720
rect 7970 6670 8130 6710
rect 7970 6660 7980 6670
rect 7900 6650 7980 6660
rect 8120 6660 8130 6670
rect 8190 6710 8200 6720
rect 8340 6720 8420 6730
rect 8340 6710 8350 6720
rect 8190 6670 8350 6710
rect 8190 6660 8200 6670
rect 8120 6650 8200 6660
rect 8340 6660 8350 6670
rect 8410 6660 8420 6720
rect 8340 6650 8420 6660
rect 9620 6720 9700 6730
rect 9620 6660 9630 6720
rect 9690 6710 9700 6720
rect 9840 6720 9920 6730
rect 9840 6710 9850 6720
rect 9690 6670 9850 6710
rect 9690 6660 9700 6670
rect 9620 6650 9700 6660
rect 9840 6660 9850 6670
rect 9910 6710 9920 6720
rect 10060 6720 10140 6730
rect 10060 6710 10070 6720
rect 9910 6670 10070 6710
rect 9910 6660 9920 6670
rect 9840 6650 9920 6660
rect 10060 6660 10070 6670
rect 10130 6710 10140 6720
rect 10130 6670 12200 6710
rect 10130 6660 10140 6670
rect 10060 6650 10140 6660
rect 132 6580 142 6650
rect 212 6580 222 6650
rect 9130 6630 9210 6640
rect 2370 6580 2450 6590
rect -220 6520 -140 6530
rect -220 6460 -210 6520
rect -150 6510 -140 6520
rect 132 6510 142 6530
rect -150 6470 142 6510
rect -150 6460 -140 6470
rect 132 6460 142 6470
rect 212 6460 222 6530
rect 2370 6520 2380 6580
rect 2440 6570 2450 6580
rect 2580 6580 2660 6590
rect 2580 6570 2590 6580
rect 2440 6530 2590 6570
rect 2440 6520 2450 6530
rect 2370 6510 2450 6520
rect 2580 6520 2590 6530
rect 2650 6520 2660 6580
rect 9130 6570 9140 6630
rect 9200 6620 9210 6630
rect 9200 6610 10020 6620
rect 9200 6580 9950 6610
rect 9200 6570 9210 6580
rect 9130 6560 9210 6570
rect 9940 6550 9950 6580
rect 10010 6550 10020 6610
rect 9940 6540 10020 6550
rect 9220 6520 9300 6530
rect 2580 6510 2660 6520
rect 5110 6510 5190 6520
rect -220 6450 -140 6460
rect 5110 6450 5120 6510
rect 5180 6500 5190 6510
rect 5220 6510 5300 6520
rect 5220 6500 5230 6510
rect 5180 6460 5230 6500
rect 5180 6450 5190 6460
rect 5110 6440 5190 6450
rect 5220 6450 5230 6460
rect 5290 6450 5300 6510
rect 9220 6460 9230 6520
rect 9290 6510 9300 6520
rect 10120 6520 10200 6530
rect 10120 6510 10130 6520
rect 9290 6470 10130 6510
rect 9290 6460 9300 6470
rect 9220 6450 9300 6460
rect 10120 6460 10130 6470
rect 10190 6460 10200 6520
rect 10120 6450 10200 6460
rect 5220 6440 5300 6450
rect -220 6390 -140 6400
rect -220 6330 -210 6390
rect -150 6380 -140 6390
rect 1190 6390 1270 6400
rect 1190 6380 1200 6390
rect -150 6340 1200 6380
rect -150 6330 -140 6340
rect -220 6320 -140 6330
rect 1190 6330 1200 6340
rect 1260 6330 1270 6390
rect 4840 6360 4850 6430
rect 4920 6410 4930 6430
rect 6120 6420 6200 6430
rect 6120 6410 6130 6420
rect 4920 6370 6130 6410
rect 4920 6360 4930 6370
rect 6120 6360 6130 6370
rect 6190 6360 6200 6420
rect 6120 6350 6200 6360
rect 9310 6410 9390 6420
rect 9310 6350 9320 6410
rect 9380 6400 9390 6410
rect 10030 6410 10110 6420
rect 10030 6400 10040 6410
rect 9380 6360 10040 6400
rect 9380 6350 9390 6360
rect 9310 6340 9390 6350
rect 10030 6350 10040 6360
rect 10100 6350 10110 6410
rect 10030 6340 10110 6350
rect 1190 6320 1270 6330
rect 5110 6330 5190 6340
rect 4840 6310 4930 6320
rect 4840 6240 4850 6310
rect 4920 6240 4930 6310
rect 5110 6270 5120 6330
rect 5180 6320 5190 6330
rect 7460 6330 7540 6340
rect 7460 6320 7470 6330
rect 5180 6280 7470 6320
rect 5180 6270 5190 6280
rect 5110 6260 5190 6270
rect 7460 6270 7470 6280
rect 7530 6270 7540 6330
rect 7460 6260 7540 6270
rect 8560 6320 8640 6330
rect 8560 6260 8570 6320
rect 8630 6310 8640 6320
rect 11230 6320 11310 6330
rect 11230 6310 11240 6320
rect 8630 6270 11240 6310
rect 8630 6260 8640 6270
rect 4840 6230 4930 6240
rect 8120 6250 8200 6260
rect 8560 6250 8640 6260
rect 11230 6260 11240 6270
rect 11300 6260 11310 6320
rect 11230 6250 11310 6260
rect 8120 6190 8130 6250
rect 8190 6220 8200 6250
rect 8190 6190 12200 6220
rect 8120 6180 12200 6190
rect 6500 6130 6580 6140
rect -120 6110 -40 6120
rect -120 6050 -110 6110
rect -50 6100 -40 6110
rect 522 6100 532 6120
rect -50 6060 532 6100
rect -50 6050 -40 6060
rect 522 6050 532 6060
rect 602 6050 612 6120
rect 1868 6050 1878 6120
rect 1948 6100 1958 6120
rect 2420 6110 2500 6120
rect 2420 6100 2430 6110
rect 1948 6060 2430 6100
rect 1948 6050 1958 6060
rect 2420 6050 2430 6060
rect 2490 6050 2500 6110
rect 6500 6100 6510 6130
rect -120 6040 -40 6050
rect 2420 6040 2500 6050
rect 5650 6070 6510 6100
rect 6570 6120 6580 6130
rect 6860 6130 6940 6140
rect 6860 6120 6870 6130
rect 6570 6080 6870 6120
rect 6570 6070 6580 6080
rect 5650 6060 6580 6070
rect 6860 6070 6870 6080
rect 6930 6120 6940 6130
rect 7220 6130 7300 6140
rect 7220 6120 7230 6130
rect 6930 6080 7230 6120
rect 6930 6070 6940 6080
rect 6860 6060 6940 6070
rect 7220 6070 7230 6080
rect 7290 6120 7300 6130
rect 7580 6130 7660 6140
rect 7580 6120 7590 6130
rect 7290 6080 7590 6120
rect 7290 6070 7300 6080
rect 7220 6060 7300 6070
rect 7580 6070 7590 6080
rect 7650 6120 7660 6130
rect 7940 6130 8020 6140
rect 7940 6120 7950 6130
rect 7650 6080 7950 6120
rect 7650 6070 7660 6080
rect 7580 6060 7660 6070
rect 7940 6070 7950 6080
rect 8010 6120 8020 6130
rect 8300 6130 8380 6140
rect 8300 6120 8310 6130
rect 8010 6080 8310 6120
rect 8010 6070 8020 6080
rect 7940 6060 8020 6070
rect 8300 6070 8310 6080
rect 8370 6120 8380 6130
rect 8660 6130 8740 6140
rect 8660 6120 8670 6130
rect 8370 6080 8670 6120
rect 8370 6070 8380 6080
rect 8300 6060 8380 6070
rect 8660 6070 8670 6080
rect 8730 6120 8740 6130
rect 9020 6130 9100 6140
rect 9020 6120 9030 6130
rect 8730 6080 9030 6120
rect 8730 6070 8740 6080
rect 8660 6060 8740 6070
rect 9020 6070 9030 6080
rect 9090 6120 9100 6130
rect 9380 6130 9460 6140
rect 9380 6120 9390 6130
rect 9090 6080 9390 6120
rect 9090 6070 9100 6080
rect 9020 6060 9100 6070
rect 9380 6070 9390 6080
rect 9450 6120 9460 6130
rect 9740 6130 9820 6140
rect 9740 6120 9750 6130
rect 9450 6080 9750 6120
rect 9450 6070 9460 6080
rect 9380 6060 9460 6070
rect 9740 6070 9750 6080
rect 9810 6120 9820 6130
rect 11500 6130 11580 6140
rect 11500 6120 11510 6130
rect 9810 6080 11510 6120
rect 9810 6070 9820 6080
rect 9740 6060 9820 6070
rect 5650 6050 5730 6060
rect 5650 5990 5660 6050
rect 5720 5990 5730 6050
rect 5650 5980 5730 5990
rect 10580 6050 10660 6080
rect 11500 6070 11510 6080
rect 11570 6070 11580 6130
rect 11500 6060 11580 6070
rect 10580 5990 10590 6050
rect 10650 5990 10660 6050
rect 10580 5980 10660 5990
rect 5650 5930 5730 5940
rect 2210 5900 2290 5910
rect 2210 5840 2220 5900
rect 2280 5890 2290 5900
rect 3032 5890 3042 5900
rect 2280 5850 3042 5890
rect 2280 5840 2290 5850
rect 2210 5830 2290 5840
rect 3032 5830 3042 5850
rect 3112 5830 3122 5900
rect 4430 5830 4440 5900
rect 4510 5880 4520 5900
rect 4840 5890 4920 5900
rect 4840 5880 4850 5890
rect 4510 5840 4850 5880
rect 4510 5830 4520 5840
rect 4840 5830 4850 5840
rect 4910 5830 4920 5890
rect 5650 5870 5660 5930
rect 5720 5920 5730 5930
rect 6120 5930 6200 5940
rect 6120 5920 6130 5930
rect 5720 5880 6130 5920
rect 5720 5870 5730 5880
rect 5650 5860 5730 5870
rect 6120 5870 6130 5880
rect 6190 5870 6200 5930
rect 6120 5860 6200 5870
rect 10580 5930 10660 5940
rect 10580 5870 10590 5930
rect 10650 5870 10660 5930
rect 10580 5860 10660 5870
rect 4840 5820 4920 5830
rect -30 5700 50 5710
rect -30 5640 -20 5700
rect 40 5680 50 5700
rect 522 5680 532 5700
rect 40 5640 532 5680
rect -30 5630 50 5640
rect 522 5630 532 5640
rect 602 5630 612 5700
rect 1868 5630 1878 5700
rect 1948 5680 1958 5700
rect 4930 5690 5010 5700
rect 4930 5680 4940 5690
rect 1948 5640 4940 5680
rect 1948 5630 1958 5640
rect 4930 5630 4940 5640
rect 5000 5630 5010 5690
rect 4930 5620 5010 5630
rect 2420 5600 2500 5610
rect 2420 5540 2430 5600
rect 2490 5590 2500 5600
rect 4750 5600 4830 5610
rect 4750 5590 4760 5600
rect 2490 5550 4760 5590
rect 2490 5540 2500 5550
rect 2420 5530 2500 5540
rect 4750 5540 4760 5550
rect 4820 5540 4830 5600
rect 4750 5530 4830 5540
rect 5520 5590 5600 5600
rect 5520 5530 5530 5590
rect 5590 5580 5600 5590
rect 5780 5590 5860 5600
rect 5780 5580 5790 5590
rect 5590 5540 5790 5580
rect 5590 5530 5600 5540
rect 5520 5520 5600 5530
rect 5780 5530 5790 5540
rect 5850 5580 5860 5590
rect 6240 5590 6320 5600
rect 6240 5580 6250 5590
rect 5850 5540 6250 5580
rect 5850 5530 5860 5540
rect 5780 5520 5860 5530
rect 6240 5530 6250 5540
rect 6310 5530 6320 5590
rect 6240 5520 6320 5530
rect 10450 5590 10530 5600
rect 10450 5530 10460 5590
rect 10520 5580 10530 5590
rect 10710 5590 10790 5600
rect 10710 5580 10720 5590
rect 10520 5540 10720 5580
rect 10520 5530 10530 5540
rect 10450 5520 10530 5530
rect 10710 5530 10720 5540
rect 10780 5580 10790 5590
rect 10780 5540 12200 5580
rect 10780 5530 10790 5540
rect 10710 5520 10790 5530
rect 4840 5390 4920 5400
rect 4840 5330 4850 5390
rect 4910 5380 4920 5390
rect 7760 5390 7840 5400
rect 7760 5380 7770 5390
rect 4910 5340 7770 5380
rect 4910 5330 4920 5340
rect 4840 5320 4920 5330
rect 7760 5330 7770 5340
rect 7830 5380 7840 5390
rect 8480 5390 8560 5400
rect 8480 5380 8490 5390
rect 7830 5340 8490 5380
rect 7830 5330 7840 5340
rect 7760 5320 7840 5330
rect 8480 5330 8490 5340
rect 8550 5330 8560 5390
rect 8480 5320 8560 5330
rect 10120 5300 10200 5310
rect 4660 5280 4740 5290
rect 4660 5220 4670 5280
rect 4730 5270 4740 5280
rect 6120 5280 6200 5290
rect 6120 5270 6130 5280
rect 4730 5230 6130 5270
rect 4730 5220 4740 5230
rect 4660 5210 4740 5220
rect 6120 5220 6130 5230
rect 6190 5270 6200 5280
rect 7400 5280 7480 5290
rect 7400 5270 7410 5280
rect 6190 5230 7410 5270
rect 6190 5220 6200 5230
rect 6120 5210 6200 5220
rect 7400 5220 7410 5230
rect 7470 5270 7480 5280
rect 8840 5280 8920 5290
rect 8840 5270 8850 5280
rect 7470 5230 8850 5270
rect 7470 5220 7480 5230
rect 7400 5210 7480 5220
rect 8840 5220 8850 5230
rect 8910 5220 8920 5280
rect 10120 5240 10130 5300
rect 10190 5290 10200 5300
rect 11050 5300 11130 5310
rect 11050 5290 11060 5300
rect 10190 5250 11060 5290
rect 10190 5240 10200 5250
rect 10120 5230 10200 5240
rect 11050 5240 11060 5250
rect 11120 5240 11130 5300
rect 11050 5230 11130 5240
rect 8840 5210 8920 5220
rect 4550 5190 4630 5200
rect 4550 5130 4560 5190
rect 4620 5180 4630 5190
rect 5650 5190 5730 5200
rect 5650 5180 5660 5190
rect 4620 5140 5660 5180
rect 4620 5130 4630 5140
rect 4550 5120 4630 5130
rect 5650 5130 5660 5140
rect 5720 5180 5730 5190
rect 7040 5190 7120 5200
rect 7040 5180 7050 5190
rect 5720 5140 7050 5180
rect 5720 5130 5730 5140
rect 5650 5120 5730 5130
rect 7040 5130 7050 5140
rect 7110 5180 7120 5190
rect 9200 5190 9280 5200
rect 9200 5180 9210 5190
rect 7110 5140 9210 5180
rect 7110 5130 7120 5140
rect 7040 5120 7120 5130
rect 9200 5130 9210 5140
rect 9270 5130 9280 5190
rect 9200 5120 9280 5130
rect 9380 5190 9460 5200
rect 9380 5130 9390 5190
rect 9450 5180 9460 5190
rect 10030 5190 10110 5200
rect 10030 5180 10040 5190
rect 9450 5140 10040 5180
rect 9450 5130 9460 5140
rect 9380 5120 9460 5130
rect 10030 5130 10040 5140
rect 10100 5130 10110 5190
rect 10030 5120 10110 5130
rect 5220 5100 5300 5110
rect 5220 5040 5230 5100
rect 5290 5090 5300 5100
rect 6680 5100 6760 5110
rect 6680 5090 6690 5100
rect 5290 5050 6690 5090
rect 5290 5040 5300 5050
rect 5220 5030 5300 5040
rect 6680 5040 6690 5050
rect 6750 5090 6760 5100
rect 8120 5100 8200 5110
rect 8120 5090 8130 5100
rect 6750 5050 8130 5090
rect 6750 5040 6760 5050
rect 6680 5030 6760 5040
rect 8120 5040 8130 5050
rect 8190 5090 8200 5100
rect 9560 5100 9640 5110
rect 9560 5090 9570 5100
rect 8190 5050 9570 5090
rect 8190 5040 8200 5050
rect 8120 5030 8200 5040
rect 9560 5040 9570 5050
rect 9630 5090 9640 5100
rect 11140 5100 11220 5110
rect 11140 5090 11150 5100
rect 9630 5050 11150 5090
rect 9630 5040 9640 5050
rect 9560 5030 9640 5040
rect 11140 5040 11150 5050
rect 11210 5040 11220 5100
rect 11140 5030 11220 5040
rect 4750 5000 4830 5010
rect 4750 4940 4760 5000
rect 4820 4990 4830 5000
rect 8560 5000 8640 5010
rect 8560 4990 8570 5000
rect 4820 4950 8570 4990
rect 4820 4940 4830 4950
rect 4750 4930 4830 4940
rect 8560 4940 8570 4950
rect 8630 4990 8640 5000
rect 9940 5000 10020 5010
rect 9940 4990 9950 5000
rect 8630 4950 9950 4990
rect 8630 4940 8640 4950
rect 8560 4930 8640 4940
rect 9940 4940 9950 4950
rect 10010 4990 10020 5000
rect 10580 5000 10660 5010
rect 10580 4990 10590 5000
rect 10010 4950 10590 4990
rect 10010 4940 10020 4950
rect 9940 4930 10020 4940
rect 10580 4940 10590 4950
rect 10650 4940 10660 5000
rect 10580 4930 10660 4940
rect 5640 4870 5720 4880
rect 5640 4810 5650 4870
rect 5710 4860 5720 4870
rect 5880 4870 5960 4880
rect 5880 4860 5890 4870
rect 5710 4820 5890 4860
rect 5710 4810 5720 4820
rect 5640 4800 5720 4810
rect 5880 4810 5890 4820
rect 5950 4860 5960 4870
rect 6120 4870 6200 4880
rect 6120 4860 6130 4870
rect 5950 4820 6130 4860
rect 5950 4810 5960 4820
rect 5880 4800 5960 4810
rect 6120 4810 6130 4820
rect 6190 4860 6200 4870
rect 6360 4870 6440 4880
rect 6360 4860 6370 4870
rect 6190 4820 6370 4860
rect 6190 4810 6200 4820
rect 6120 4800 6200 4810
rect 6360 4810 6370 4820
rect 6430 4860 6440 4870
rect 6600 4870 6680 4880
rect 6600 4860 6610 4870
rect 6430 4820 6610 4860
rect 6430 4810 6440 4820
rect 6360 4800 6440 4810
rect 6600 4810 6610 4820
rect 6670 4860 6680 4870
rect 6840 4870 6920 4880
rect 6840 4860 6850 4870
rect 6670 4820 6850 4860
rect 6670 4810 6680 4820
rect 6600 4800 6680 4810
rect 6840 4810 6850 4820
rect 6910 4860 6920 4870
rect 7080 4870 7160 4880
rect 7080 4860 7090 4870
rect 6910 4820 7090 4860
rect 6910 4810 6920 4820
rect 6840 4800 6920 4810
rect 7080 4810 7090 4820
rect 7150 4860 7160 4870
rect 7320 4870 7400 4880
rect 7320 4860 7330 4870
rect 7150 4820 7330 4860
rect 7150 4810 7160 4820
rect 7080 4800 7160 4810
rect 7320 4810 7330 4820
rect 7390 4860 7400 4870
rect 7560 4870 7640 4880
rect 7560 4860 7570 4870
rect 7390 4820 7570 4860
rect 7390 4810 7400 4820
rect 7320 4800 7400 4810
rect 7560 4810 7570 4820
rect 7630 4860 7640 4870
rect 8680 4870 8760 4880
rect 8680 4860 8690 4870
rect 7630 4820 8690 4860
rect 7630 4810 7640 4820
rect 7560 4800 7640 4810
rect 8680 4810 8690 4820
rect 8750 4860 8760 4870
rect 8920 4870 9000 4880
rect 8920 4860 8930 4870
rect 8750 4820 8930 4860
rect 8750 4810 8760 4820
rect 8680 4800 8760 4810
rect 8920 4810 8930 4820
rect 8990 4860 9000 4870
rect 9160 4870 9240 4880
rect 9160 4860 9170 4870
rect 8990 4820 9170 4860
rect 8990 4810 9000 4820
rect 8920 4800 9000 4810
rect 9160 4810 9170 4820
rect 9230 4860 9240 4870
rect 9400 4870 9480 4880
rect 9400 4860 9410 4870
rect 9230 4820 9410 4860
rect 9230 4810 9240 4820
rect 9160 4800 9240 4810
rect 9400 4810 9410 4820
rect 9470 4860 9480 4870
rect 9640 4870 9720 4880
rect 9640 4860 9650 4870
rect 9470 4820 9650 4860
rect 9470 4810 9480 4820
rect 9400 4800 9480 4810
rect 9640 4810 9650 4820
rect 9710 4860 9720 4870
rect 9880 4870 9960 4880
rect 9880 4860 9890 4870
rect 9710 4820 9890 4860
rect 9710 4810 9720 4820
rect 9640 4800 9720 4810
rect 9880 4810 9890 4820
rect 9950 4860 9960 4870
rect 10120 4870 10200 4880
rect 10120 4860 10130 4870
rect 9950 4820 10130 4860
rect 9950 4810 9960 4820
rect 9880 4800 9960 4810
rect 10120 4810 10130 4820
rect 10190 4860 10200 4870
rect 10360 4870 10440 4880
rect 10360 4860 10370 4870
rect 10190 4820 10370 4860
rect 10190 4810 10200 4820
rect 10120 4800 10200 4810
rect 10360 4810 10370 4820
rect 10430 4860 10440 4870
rect 10600 4870 10680 4880
rect 10600 4860 10610 4870
rect 10430 4820 10610 4860
rect 10430 4810 10440 4820
rect 10360 4800 10440 4810
rect 10600 4810 10610 4820
rect 10670 4860 10680 4870
rect 11500 4870 11580 4880
rect 11500 4860 11510 4870
rect 10670 4820 11510 4860
rect 10670 4810 10680 4820
rect 10600 4800 10680 4810
rect 11500 4810 11510 4820
rect 11570 4810 11580 4870
rect 11500 4800 11580 4810
rect 4930 4750 5010 4760
rect 4930 4690 4940 4750
rect 5000 4740 5010 4750
rect 5520 4750 5600 4760
rect 5520 4740 5530 4750
rect 5000 4700 5530 4740
rect 5000 4690 5010 4700
rect 4930 4680 5010 4690
rect 5520 4690 5530 4700
rect 5590 4740 5600 4750
rect 6240 4750 6320 4760
rect 6240 4740 6250 4750
rect 5590 4700 6250 4740
rect 5590 4690 5600 4700
rect 5520 4680 5600 4690
rect 6240 4690 6250 4700
rect 6310 4740 6320 4750
rect 6960 4750 7040 4760
rect 6960 4740 6970 4750
rect 6310 4700 6970 4740
rect 6310 4690 6320 4700
rect 6240 4680 6320 4690
rect 6960 4690 6970 4700
rect 7030 4740 7040 4750
rect 7680 4750 7760 4760
rect 7680 4740 7690 4750
rect 7030 4700 7690 4740
rect 7030 4690 7040 4700
rect 6960 4680 7040 4690
rect 7680 4690 7690 4700
rect 7750 4740 7760 4750
rect 7940 4750 8020 4760
rect 7940 4740 7950 4750
rect 7750 4700 7950 4740
rect 7750 4690 7760 4700
rect 7680 4680 7760 4690
rect 7940 4690 7950 4700
rect 8010 4690 8020 4750
rect 7940 4680 8020 4690
rect 8300 4750 8380 4760
rect 8300 4690 8310 4750
rect 8370 4740 8380 4750
rect 8560 4750 8640 4760
rect 8560 4740 8570 4750
rect 8370 4700 8570 4740
rect 8370 4690 8380 4700
rect 8300 4680 8380 4690
rect 8560 4690 8570 4700
rect 8630 4740 8640 4750
rect 9280 4750 9360 4760
rect 9280 4740 9290 4750
rect 8630 4700 9290 4740
rect 8630 4690 8640 4700
rect 8560 4680 8640 4690
rect 9280 4690 9290 4700
rect 9350 4740 9360 4750
rect 10000 4750 10080 4760
rect 10000 4740 10010 4750
rect 9350 4700 10010 4740
rect 9350 4690 9360 4700
rect 9280 4680 9360 4690
rect 10000 4690 10010 4700
rect 10070 4740 10080 4750
rect 10720 4750 10800 4760
rect 10720 4740 10730 4750
rect 10070 4700 10730 4740
rect 10070 4690 10080 4700
rect 10000 4680 10080 4690
rect 10720 4690 10730 4700
rect 10790 4690 10800 4750
rect 10720 4680 10800 4690
rect 5760 4410 5840 4420
rect 5760 4350 5770 4410
rect 5830 4400 5840 4410
rect 6000 4400 6080 4420
rect 6480 4410 6560 4420
rect 6480 4400 6490 4410
rect 5830 4360 6490 4400
rect 5830 4350 5840 4360
rect 5760 4340 5840 4350
rect 6000 4340 6080 4360
rect 6480 4350 6490 4360
rect 6550 4400 6560 4410
rect 6720 4400 6800 4420
rect 7200 4410 7280 4420
rect 7200 4400 7210 4410
rect 6550 4360 7210 4400
rect 6550 4350 6560 4360
rect 6480 4340 6560 4350
rect 6720 4340 6800 4360
rect 7200 4350 7210 4360
rect 7270 4350 7280 4410
rect 7200 4340 7280 4350
rect 7440 4340 7520 4420
rect 8800 4340 8880 4420
rect 9040 4410 9120 4420
rect 9040 4350 9050 4410
rect 9110 4400 9120 4410
rect 9520 4400 9600 4420
rect 9760 4410 9840 4420
rect 9760 4400 9770 4410
rect 9110 4360 9770 4400
rect 9110 4350 9120 4360
rect 9040 4340 9120 4350
rect 9520 4340 9600 4360
rect 9760 4350 9770 4360
rect 9830 4400 9840 4410
rect 10240 4400 10320 4420
rect 10480 4410 10560 4420
rect 10480 4400 10490 4410
rect 9830 4360 10490 4400
rect 9830 4350 9840 4360
rect 9760 4340 9840 4350
rect 10240 4340 10320 4360
rect 10480 4350 10490 4360
rect 10550 4350 10560 4410
rect 10480 4340 10560 4350
rect 5020 4290 5100 4300
rect 5020 4230 5030 4290
rect 5090 4280 5100 4290
rect 5580 4290 5660 4300
rect 5580 4280 5590 4290
rect 5090 4240 5590 4280
rect 5090 4230 5100 4240
rect 5020 4220 5100 4230
rect 5580 4230 5590 4240
rect 5650 4280 5660 4290
rect 6000 4290 6080 4300
rect 6000 4280 6010 4290
rect 5650 4240 6010 4280
rect 5650 4230 5660 4240
rect 5580 4220 5660 4230
rect 6000 4230 6010 4240
rect 6070 4280 6080 4290
rect 6240 4290 6320 4300
rect 6240 4280 6250 4290
rect 6070 4240 6250 4280
rect 6070 4230 6080 4240
rect 6000 4220 6080 4230
rect 6240 4230 6250 4240
rect 6310 4280 6320 4290
rect 6720 4290 6800 4300
rect 6720 4280 6730 4290
rect 6310 4240 6730 4280
rect 6310 4230 6320 4240
rect 6240 4220 6320 4230
rect 6720 4230 6730 4240
rect 6790 4280 6800 4290
rect 6960 4290 7040 4300
rect 6960 4280 6970 4290
rect 6790 4240 6970 4280
rect 6790 4230 6800 4240
rect 6720 4220 6800 4230
rect 6960 4230 6970 4240
rect 7030 4280 7040 4290
rect 7440 4290 7520 4300
rect 7440 4280 7450 4290
rect 7030 4240 7450 4280
rect 7030 4230 7040 4240
rect 6960 4220 7040 4230
rect 7440 4230 7450 4240
rect 7510 4280 7520 4290
rect 7620 4290 7700 4300
rect 7620 4280 7630 4290
rect 7510 4240 7630 4280
rect 7510 4230 7520 4240
rect 7440 4220 7520 4230
rect 7620 4230 7630 4240
rect 7690 4230 7700 4290
rect 7620 4220 7700 4230
rect 8620 4290 8700 4300
rect 8620 4230 8630 4290
rect 8690 4280 8700 4290
rect 8800 4290 8880 4300
rect 8800 4280 8810 4290
rect 8690 4240 8810 4280
rect 8690 4230 8700 4240
rect 8620 4220 8700 4230
rect 8800 4230 8810 4240
rect 8870 4280 8880 4290
rect 9280 4290 9360 4300
rect 9280 4280 9290 4290
rect 8870 4240 9290 4280
rect 8870 4230 8880 4240
rect 8800 4220 8880 4230
rect 9280 4230 9290 4240
rect 9350 4280 9360 4290
rect 9520 4290 9600 4300
rect 9520 4280 9530 4290
rect 9350 4240 9530 4280
rect 9350 4230 9360 4240
rect 9280 4220 9360 4230
rect 9520 4230 9530 4240
rect 9590 4280 9600 4290
rect 10000 4290 10080 4300
rect 10000 4280 10010 4290
rect 9590 4240 10010 4280
rect 9590 4230 9600 4240
rect 9520 4220 9600 4230
rect 10000 4230 10010 4240
rect 10070 4280 10080 4290
rect 10240 4290 10320 4300
rect 10240 4280 10250 4290
rect 10070 4240 10250 4280
rect 10070 4230 10080 4240
rect 10000 4220 10080 4230
rect 10240 4230 10250 4240
rect 10310 4280 10320 4290
rect 10660 4290 10740 4300
rect 10660 4280 10670 4290
rect 10310 4240 10670 4280
rect 10310 4230 10320 4240
rect 10240 4220 10320 4230
rect 10660 4230 10670 4240
rect 10730 4280 10740 4290
rect 11050 4290 11130 4300
rect 11050 4280 11060 4290
rect 10730 4240 11060 4280
rect 10730 4230 10740 4240
rect 10660 4220 10740 4230
rect 11050 4230 11060 4240
rect 11120 4230 11130 4290
rect 11050 4220 11130 4230
rect 36620 4270 36700 4280
rect 36620 4210 36630 4270
rect 36690 4260 36700 4270
rect 36690 4220 42200 4260
rect 36690 4210 36700 4220
rect 36620 4200 36700 4210
rect 36400 4180 36480 4190
rect 6500 4120 6580 4130
rect 4660 4090 4740 4100
rect 4660 4030 4670 4090
rect 4730 4080 4740 4090
rect 6380 4090 6460 4100
rect 6380 4080 6390 4090
rect 4730 4040 6390 4080
rect 4730 4030 4740 4040
rect 4660 4020 4740 4030
rect 6380 4030 6390 4040
rect 6450 4030 6460 4090
rect 6500 4060 6510 4120
rect 6570 4110 6580 4120
rect 6980 4120 7060 4130
rect 6980 4110 6990 4120
rect 6570 4070 6990 4110
rect 6570 4060 6580 4070
rect 6500 4050 6580 4060
rect 6980 4060 6990 4070
rect 7050 4110 7060 4120
rect 7460 4120 7540 4130
rect 7460 4110 7470 4120
rect 7050 4070 7470 4110
rect 7050 4060 7060 4070
rect 6980 4050 7060 4060
rect 7460 4060 7470 4070
rect 7530 4060 7540 4120
rect 7460 4050 7540 4060
rect 8780 4120 8860 4130
rect 8780 4060 8790 4120
rect 8850 4110 8860 4120
rect 9260 4120 9340 4130
rect 9260 4110 9270 4120
rect 8850 4070 9270 4110
rect 8850 4060 8860 4070
rect 8780 4050 8860 4060
rect 9260 4060 9270 4070
rect 9330 4110 9340 4120
rect 9740 4120 9820 4130
rect 9740 4110 9750 4120
rect 9330 4070 9750 4110
rect 9330 4060 9340 4070
rect 9260 4050 9340 4060
rect 9740 4060 9750 4070
rect 9810 4060 9820 4120
rect 36400 4120 36410 4180
rect 36470 4170 36480 4180
rect 38120 4180 38200 4190
rect 38120 4170 38130 4180
rect 36470 4130 38130 4170
rect 36470 4120 36480 4130
rect 36400 4110 36480 4120
rect 38120 4120 38130 4130
rect 38190 4170 38200 4180
rect 39130 4180 39210 4190
rect 39130 4170 39140 4180
rect 38190 4130 39140 4170
rect 38190 4120 38200 4130
rect 38120 4110 38200 4120
rect 39130 4120 39140 4130
rect 39200 4170 39210 4180
rect 39840 4180 39920 4190
rect 39840 4170 39850 4180
rect 39200 4130 39850 4170
rect 39200 4120 39210 4130
rect 39130 4110 39210 4120
rect 39840 4120 39850 4130
rect 39910 4120 39920 4180
rect 39840 4110 39920 4120
rect 9740 4050 9820 4060
rect 9860 4090 9940 4100
rect 6380 4020 6460 4030
rect 9860 4030 9870 4090
rect 9930 4080 9940 4090
rect 11140 4090 11220 4100
rect 11140 4080 11150 4090
rect 9930 4040 11150 4080
rect 9930 4030 9940 4040
rect 9860 4020 9940 4030
rect 11140 4030 11150 4040
rect 11210 4080 11220 4090
rect 11210 4040 12200 4080
rect 36070 4060 36150 4070
rect 11210 4030 11220 4040
rect 11140 4020 11220 4030
rect 6260 4000 6340 4010
rect 6260 3940 6270 4000
rect 6330 3990 6340 4000
rect 6740 4000 6820 4010
rect 6740 3990 6750 4000
rect 6330 3950 6750 3990
rect 6330 3940 6340 3950
rect 6260 3930 6340 3940
rect 6740 3940 6750 3950
rect 6810 3990 6820 4000
rect 7220 4000 7300 4010
rect 7220 3990 7230 4000
rect 6810 3950 7230 3990
rect 6810 3940 6820 3950
rect 6740 3930 6820 3940
rect 7220 3940 7230 3950
rect 7290 3940 7300 4000
rect 7220 3930 7300 3940
rect 9020 4000 9100 4010
rect 9020 3940 9030 4000
rect 9090 3990 9100 4000
rect 9500 4000 9580 4010
rect 9500 3990 9510 4000
rect 9090 3950 9510 3990
rect 9090 3940 9100 3950
rect 9020 3930 9100 3940
rect 9500 3940 9510 3950
rect 9570 3990 9580 4000
rect 9980 4000 10060 4010
rect 9980 3990 9990 4000
rect 9570 3950 9990 3990
rect 9570 3940 9580 3950
rect 9500 3930 9580 3940
rect 9980 3940 9990 3950
rect 10050 3940 10060 4000
rect 36070 4000 36080 4060
rect 36140 4050 36150 4060
rect 36290 4060 36370 4070
rect 36290 4050 36300 4060
rect 36140 4010 36300 4050
rect 36140 4000 36150 4010
rect 36070 3990 36150 4000
rect 36290 4000 36300 4010
rect 36360 4050 36370 4060
rect 36510 4060 36590 4070
rect 36510 4050 36520 4060
rect 36360 4010 36520 4050
rect 36360 4000 36370 4010
rect 36290 3990 36370 4000
rect 36510 4000 36520 4010
rect 36580 4050 36590 4060
rect 36730 4060 36810 4070
rect 36730 4050 36740 4060
rect 36580 4010 36740 4050
rect 36580 4000 36590 4010
rect 36510 3990 36590 4000
rect 36730 4000 36740 4010
rect 36800 4050 36810 4060
rect 37350 4060 37430 4070
rect 37350 4050 37360 4060
rect 36800 4010 37360 4050
rect 36800 4000 36810 4010
rect 36730 3990 36810 4000
rect 37350 4000 37360 4010
rect 37420 4050 37430 4060
rect 37570 4060 37650 4070
rect 37570 4050 37580 4060
rect 37420 4010 37580 4050
rect 37420 4000 37430 4010
rect 37350 3990 37430 4000
rect 37570 4000 37580 4010
rect 37640 4050 37650 4060
rect 37790 4060 37870 4070
rect 37790 4050 37800 4060
rect 37640 4010 37800 4050
rect 37640 4000 37650 4010
rect 37570 3990 37650 4000
rect 37790 4000 37800 4010
rect 37860 4050 37870 4060
rect 38010 4060 38090 4070
rect 38010 4050 38020 4060
rect 37860 4010 38020 4050
rect 37860 4000 37870 4010
rect 37790 3990 37870 4000
rect 38010 4000 38020 4010
rect 38080 4050 38090 4060
rect 38230 4060 38310 4070
rect 38230 4050 38240 4060
rect 38080 4010 38240 4050
rect 38080 4000 38090 4010
rect 38010 3990 38090 4000
rect 38230 4000 38240 4010
rect 38300 4050 38310 4060
rect 38450 4060 38530 4070
rect 38450 4050 38460 4060
rect 38300 4010 38460 4050
rect 38300 4000 38310 4010
rect 38230 3990 38310 4000
rect 38450 4000 38460 4010
rect 38520 4050 38530 4060
rect 38670 4060 38750 4070
rect 38670 4050 38680 4060
rect 38520 4010 38680 4050
rect 38520 4000 38530 4010
rect 38450 3990 38530 4000
rect 38670 4000 38680 4010
rect 38740 4050 38750 4060
rect 39510 4060 39590 4070
rect 39510 4050 39520 4060
rect 38740 4010 39520 4050
rect 38740 4000 38750 4010
rect 38670 3990 38750 4000
rect 39510 4000 39520 4010
rect 39580 4050 39590 4060
rect 39730 4060 39810 4070
rect 39730 4050 39740 4060
rect 39580 4010 39740 4050
rect 39580 4000 39590 4010
rect 39510 3990 39590 4000
rect 39730 4000 39740 4010
rect 39800 4050 39810 4060
rect 39950 4060 40030 4070
rect 39950 4050 39960 4060
rect 39800 4010 39960 4050
rect 39800 4000 39810 4010
rect 39730 3990 39810 4000
rect 39950 4000 39960 4010
rect 40020 4050 40030 4060
rect 40170 4060 40250 4070
rect 40170 4050 40180 4060
rect 40020 4010 40180 4050
rect 40020 4000 40030 4010
rect 39950 3990 40030 4000
rect 40170 4000 40180 4010
rect 40240 4050 40250 4060
rect 41500 4060 41580 4070
rect 41500 4050 41510 4060
rect 40240 4010 41510 4050
rect 40240 4000 40250 4010
rect 40170 3990 40250 4000
rect 41500 4000 41510 4010
rect 41570 4000 41580 4060
rect 41500 3990 41580 4000
rect 9980 3930 10060 3940
rect 7580 3880 7660 3890
rect 7580 3820 7590 3880
rect 7650 3870 7660 3880
rect 8120 3880 8200 3890
rect 8120 3870 8130 3880
rect 7650 3830 8130 3870
rect 7650 3820 7660 3830
rect 7580 3810 7660 3820
rect 8120 3820 8130 3830
rect 8190 3870 8200 3880
rect 8660 3880 8740 3890
rect 8660 3870 8670 3880
rect 8190 3830 8670 3870
rect 8190 3820 8200 3830
rect 8120 3810 8200 3820
rect 8660 3820 8670 3830
rect 8730 3820 8740 3880
rect 8660 3810 8740 3820
rect 4840 3760 4920 3770
rect 4840 3700 4850 3760
rect 4910 3750 4920 3760
rect 6260 3760 6340 3770
rect 6260 3750 6270 3760
rect 4910 3710 6270 3750
rect 4910 3700 4920 3710
rect 4840 3690 4920 3700
rect 6260 3700 6270 3710
rect 6330 3700 6340 3760
rect 6260 3690 6340 3700
rect 9980 3760 10060 3770
rect 9980 3700 9990 3760
rect 10050 3750 10060 3760
rect 11230 3760 11310 3770
rect 11230 3750 11240 3760
rect 10050 3710 11240 3750
rect 10050 3700 10060 3710
rect 9980 3690 10060 3700
rect 11230 3700 11240 3710
rect 11300 3700 11310 3760
rect 11230 3690 11310 3700
rect 36180 3720 36260 3730
rect 36180 3660 36190 3720
rect 36250 3710 36260 3720
rect 36400 3720 36480 3730
rect 36400 3710 36410 3720
rect 36250 3670 36410 3710
rect 36250 3660 36260 3670
rect 36180 3650 36260 3660
rect 36400 3660 36410 3670
rect 36470 3710 36480 3720
rect 36620 3720 36700 3730
rect 36620 3710 36630 3720
rect 36470 3670 36630 3710
rect 36470 3660 36480 3670
rect 36400 3650 36480 3660
rect 36620 3660 36630 3670
rect 36690 3660 36700 3720
rect 36620 3650 36700 3660
rect 37680 3720 37760 3730
rect 37680 3660 37690 3720
rect 37750 3710 37760 3720
rect 37900 3720 37980 3730
rect 37900 3710 37910 3720
rect 37750 3670 37910 3710
rect 37750 3660 37760 3670
rect 37680 3650 37760 3660
rect 37900 3660 37910 3670
rect 37970 3710 37980 3720
rect 38120 3720 38200 3730
rect 38120 3710 38130 3720
rect 37970 3670 38130 3710
rect 37970 3660 37980 3670
rect 37900 3650 37980 3660
rect 38120 3660 38130 3670
rect 38190 3710 38200 3720
rect 38340 3720 38420 3730
rect 38340 3710 38350 3720
rect 38190 3670 38350 3710
rect 38190 3660 38200 3670
rect 38120 3650 38200 3660
rect 38340 3660 38350 3670
rect 38410 3660 38420 3720
rect 38340 3650 38420 3660
rect 39620 3720 39700 3730
rect 39620 3660 39630 3720
rect 39690 3710 39700 3720
rect 39840 3720 39920 3730
rect 39840 3710 39850 3720
rect 39690 3670 39850 3710
rect 39690 3660 39700 3670
rect 39620 3650 39700 3660
rect 39840 3660 39850 3670
rect 39910 3710 39920 3720
rect 40060 3720 40140 3730
rect 40060 3710 40070 3720
rect 39910 3670 40070 3710
rect 39910 3660 39920 3670
rect 39840 3650 39920 3660
rect 40060 3660 40070 3670
rect 40130 3710 40140 3720
rect 40130 3670 42200 3710
rect 40130 3660 40140 3670
rect 40060 3650 40140 3660
rect 5780 3640 5860 3650
rect 5780 3580 5790 3640
rect 5850 3630 5860 3640
rect 6380 3640 6460 3650
rect 6380 3630 6390 3640
rect 5850 3590 6390 3630
rect 5850 3580 5860 3590
rect 5780 3570 5860 3580
rect 6380 3580 6390 3590
rect 6450 3630 6460 3640
rect 6620 3640 6700 3650
rect 6620 3630 6630 3640
rect 6450 3590 6630 3630
rect 6450 3580 6460 3590
rect 6380 3570 6460 3580
rect 6620 3580 6630 3590
rect 6690 3630 6700 3640
rect 6860 3640 6940 3650
rect 6860 3630 6870 3640
rect 6690 3590 6870 3630
rect 6690 3580 6700 3590
rect 6620 3570 6700 3580
rect 6860 3580 6870 3590
rect 6930 3630 6940 3640
rect 7100 3640 7180 3650
rect 7100 3630 7110 3640
rect 6930 3590 7110 3630
rect 6930 3580 6940 3590
rect 6860 3570 6940 3580
rect 7100 3580 7110 3590
rect 7170 3630 7180 3640
rect 7340 3640 7420 3650
rect 7340 3630 7350 3640
rect 7170 3590 7350 3630
rect 7170 3580 7180 3590
rect 7100 3570 7180 3580
rect 7340 3580 7350 3590
rect 7410 3580 7420 3640
rect 7340 3570 7420 3580
rect 8900 3640 8980 3650
rect 8900 3580 8910 3640
rect 8970 3630 8980 3640
rect 9140 3640 9220 3650
rect 9140 3630 9150 3640
rect 8970 3590 9150 3630
rect 8970 3580 8980 3590
rect 8900 3570 8980 3580
rect 9140 3580 9150 3590
rect 9210 3630 9220 3640
rect 9380 3640 9460 3650
rect 9380 3630 9390 3640
rect 9210 3590 9390 3630
rect 9210 3580 9220 3590
rect 9140 3570 9220 3580
rect 9380 3580 9390 3590
rect 9450 3630 9460 3640
rect 9620 3640 9700 3650
rect 9620 3630 9630 3640
rect 9450 3590 9630 3630
rect 9450 3580 9460 3590
rect 9380 3570 9460 3580
rect 9620 3580 9630 3590
rect 9690 3630 9700 3640
rect 9860 3640 9940 3650
rect 9860 3630 9870 3640
rect 9690 3590 9870 3630
rect 9690 3580 9700 3590
rect 9620 3570 9700 3580
rect 9860 3580 9870 3590
rect 9930 3630 9940 3640
rect 10460 3640 10540 3650
rect 10460 3630 10470 3640
rect 9930 3590 10470 3630
rect 9930 3580 9940 3590
rect 9860 3570 9940 3580
rect 10460 3580 10470 3590
rect 10530 3580 10540 3640
rect 10460 3570 10540 3580
rect 39130 3630 39210 3640
rect 39130 3570 39140 3630
rect 39200 3620 39210 3630
rect 39200 3610 40020 3620
rect 39200 3580 39950 3610
rect 39200 3570 39210 3580
rect 39130 3560 39210 3570
rect 39940 3550 39950 3580
rect 40010 3550 40020 3610
rect 39940 3540 40020 3550
rect 39220 3520 39300 3530
rect 39220 3460 39230 3520
rect 39290 3510 39300 3520
rect 40120 3520 40200 3530
rect 40120 3510 40130 3520
rect 39290 3470 40130 3510
rect 39290 3460 39300 3470
rect 39220 3450 39300 3460
rect 40120 3460 40130 3470
rect 40190 3460 40200 3520
rect 40120 3450 40200 3460
rect -220 3440 -140 3450
rect -220 3380 -210 3440
rect -150 3380 -140 3440
rect -220 3370 -140 3380
rect -90 3440 -10 3450
rect -90 3380 -80 3440
rect -20 3380 -10 3440
rect 5960 3440 6040 3450
rect -90 3370 -10 3380
rect 2524 3420 2604 3430
rect 2524 3360 2540 3420
rect 2594 3410 2604 3420
rect 4660 3420 4740 3430
rect 4660 3410 4670 3420
rect 2594 3370 4670 3410
rect 2594 3360 2604 3370
rect 2524 3350 2604 3360
rect 4660 3360 4670 3370
rect 4730 3360 4740 3420
rect 5960 3380 5970 3440
rect 6030 3430 6040 3440
rect 6200 3440 6280 3450
rect 6200 3430 6210 3440
rect 6030 3390 6210 3430
rect 6030 3380 6040 3390
rect 5960 3370 6040 3380
rect 6200 3380 6210 3390
rect 6270 3430 6280 3440
rect 6440 3440 6520 3450
rect 6440 3430 6450 3440
rect 6270 3390 6450 3430
rect 6270 3380 6280 3390
rect 6200 3370 6280 3380
rect 6440 3380 6450 3390
rect 6510 3430 6520 3440
rect 6680 3440 6760 3450
rect 6680 3430 6690 3440
rect 6510 3390 6690 3430
rect 6510 3380 6520 3390
rect 6440 3370 6520 3380
rect 6680 3380 6690 3390
rect 6750 3430 6760 3440
rect 7160 3440 7240 3450
rect 7160 3430 7170 3440
rect 6750 3390 7170 3430
rect 6750 3380 6760 3390
rect 6680 3370 6760 3380
rect 7160 3380 7170 3390
rect 7230 3430 7240 3440
rect 7400 3440 7480 3450
rect 7400 3430 7410 3440
rect 7230 3390 7410 3430
rect 7230 3380 7240 3390
rect 7160 3370 7240 3380
rect 7400 3380 7410 3390
rect 7470 3430 7480 3440
rect 7640 3440 7720 3450
rect 7640 3430 7650 3440
rect 7470 3390 7650 3430
rect 7470 3380 7480 3390
rect 7400 3370 7480 3380
rect 7640 3380 7650 3390
rect 7710 3430 7720 3440
rect 8600 3440 8680 3450
rect 8600 3430 8610 3440
rect 7710 3390 8610 3430
rect 7710 3380 7720 3390
rect 7640 3370 7720 3380
rect 8600 3380 8610 3390
rect 8670 3430 8680 3440
rect 8840 3440 8920 3450
rect 8840 3430 8850 3440
rect 8670 3390 8850 3430
rect 8670 3380 8680 3390
rect 8600 3370 8680 3380
rect 8840 3380 8850 3390
rect 8910 3430 8920 3440
rect 9080 3440 9160 3450
rect 9080 3430 9090 3440
rect 8910 3390 9090 3430
rect 8910 3380 8920 3390
rect 8840 3370 8920 3380
rect 9080 3380 9090 3390
rect 9150 3430 9160 3440
rect 9560 3440 9640 3450
rect 9560 3430 9570 3440
rect 9150 3390 9570 3430
rect 9150 3380 9160 3390
rect 9080 3370 9160 3380
rect 9560 3380 9570 3390
rect 9630 3430 9640 3440
rect 9800 3440 9880 3450
rect 9800 3430 9810 3440
rect 9630 3390 9810 3430
rect 9630 3380 9640 3390
rect 9560 3370 9640 3380
rect 9800 3380 9810 3390
rect 9870 3430 9880 3440
rect 10040 3440 10120 3450
rect 10040 3430 10050 3440
rect 9870 3390 10050 3430
rect 9870 3380 9880 3390
rect 9800 3370 9880 3380
rect 10040 3380 10050 3390
rect 10110 3430 10120 3440
rect 10280 3440 10360 3450
rect 10280 3430 10290 3440
rect 10110 3390 10290 3430
rect 10110 3380 10120 3390
rect 10040 3370 10120 3380
rect 10280 3380 10290 3390
rect 10350 3430 10360 3440
rect 11500 3440 11580 3450
rect 11500 3430 11510 3440
rect 10350 3390 11510 3430
rect 10350 3380 10360 3390
rect 10280 3370 10360 3380
rect 11500 3380 11510 3390
rect 11570 3380 11580 3440
rect 36120 3420 36200 3430
rect 36120 3410 36130 3420
rect 11500 3370 11580 3380
rect 35250 3370 36130 3410
rect 4660 3350 4740 3360
rect 36120 3360 36130 3370
rect 36190 3360 36200 3420
rect 36120 3350 36200 3360
rect 39310 3410 39390 3420
rect 39310 3350 39320 3410
rect 39380 3400 39390 3410
rect 40030 3410 40110 3420
rect 40030 3400 40040 3410
rect 39380 3360 40040 3400
rect 39380 3350 39390 3360
rect 39310 3340 39390 3350
rect 40030 3350 40040 3360
rect 40100 3350 40110 3410
rect 40030 3340 40110 3350
rect 37460 3330 37540 3340
rect 37460 3320 37470 3330
rect 35250 3280 37470 3320
rect 37460 3270 37470 3280
rect 37530 3270 37540 3330
rect 37460 3260 37540 3270
rect 38560 3320 38640 3330
rect 38560 3260 38570 3320
rect 38630 3310 38640 3320
rect 41230 3320 41310 3330
rect 41230 3310 41240 3320
rect 38630 3270 41240 3310
rect 38630 3260 38640 3270
rect 38120 3250 38200 3260
rect 38560 3250 38640 3260
rect 41230 3260 41240 3270
rect 41300 3260 41310 3320
rect 41230 3250 41310 3260
rect 38120 3190 38130 3250
rect 38190 3220 38200 3250
rect 38190 3190 42200 3220
rect 38120 3180 42200 3190
rect 36500 3130 36580 3140
rect 36500 3100 36510 3130
rect 35650 3070 36510 3100
rect 36570 3120 36580 3130
rect 36860 3130 36940 3140
rect 36860 3120 36870 3130
rect 36570 3080 36870 3120
rect 36570 3070 36580 3080
rect 35650 3060 36580 3070
rect 36860 3070 36870 3080
rect 36930 3120 36940 3130
rect 37220 3130 37300 3140
rect 37220 3120 37230 3130
rect 36930 3080 37230 3120
rect 36930 3070 36940 3080
rect 36860 3060 36940 3070
rect 37220 3070 37230 3080
rect 37290 3120 37300 3130
rect 37580 3130 37660 3140
rect 37580 3120 37590 3130
rect 37290 3080 37590 3120
rect 37290 3070 37300 3080
rect 37220 3060 37300 3070
rect 37580 3070 37590 3080
rect 37650 3120 37660 3130
rect 37940 3130 38020 3140
rect 37940 3120 37950 3130
rect 37650 3080 37950 3120
rect 37650 3070 37660 3080
rect 37580 3060 37660 3070
rect 37940 3070 37950 3080
rect 38010 3120 38020 3130
rect 38300 3130 38380 3140
rect 38300 3120 38310 3130
rect 38010 3080 38310 3120
rect 38010 3070 38020 3080
rect 37940 3060 38020 3070
rect 38300 3070 38310 3080
rect 38370 3120 38380 3130
rect 38660 3130 38740 3140
rect 38660 3120 38670 3130
rect 38370 3080 38670 3120
rect 38370 3070 38380 3080
rect 38300 3060 38380 3070
rect 38660 3070 38670 3080
rect 38730 3120 38740 3130
rect 39020 3130 39100 3140
rect 39020 3120 39030 3130
rect 38730 3080 39030 3120
rect 38730 3070 38740 3080
rect 38660 3060 38740 3070
rect 39020 3070 39030 3080
rect 39090 3120 39100 3130
rect 39380 3130 39460 3140
rect 39380 3120 39390 3130
rect 39090 3080 39390 3120
rect 39090 3070 39100 3080
rect 39020 3060 39100 3070
rect 39380 3070 39390 3080
rect 39450 3120 39460 3130
rect 39740 3130 39820 3140
rect 39740 3120 39750 3130
rect 39450 3080 39750 3120
rect 39450 3070 39460 3080
rect 39380 3060 39460 3070
rect 39740 3070 39750 3080
rect 39810 3120 39820 3130
rect 41500 3130 41580 3140
rect 41500 3120 41510 3130
rect 39810 3080 41510 3120
rect 39810 3070 39820 3080
rect 39740 3060 39820 3070
rect 35650 3050 35730 3060
rect 35650 2990 35660 3050
rect 35720 2990 35730 3050
rect 35650 2980 35730 2990
rect 40580 3050 40660 3080
rect 41500 3070 41510 3080
rect 41570 3070 41580 3130
rect 41500 3060 41580 3070
rect 40580 2990 40590 3050
rect 40650 2990 40660 3050
rect 40580 2980 40660 2990
rect 35650 2930 35730 2940
rect 35650 2870 35660 2930
rect 35720 2920 35730 2930
rect 36120 2930 36200 2940
rect 36120 2920 36130 2930
rect 35720 2880 36130 2920
rect 35720 2870 35730 2880
rect 35650 2860 35730 2870
rect 36120 2870 36130 2880
rect 36190 2870 36200 2930
rect 36120 2860 36200 2870
rect 40580 2930 40660 2940
rect 40580 2870 40590 2930
rect 40650 2870 40660 2930
rect 40580 2860 40660 2870
rect 6860 2810 6940 2820
rect 6860 2750 6870 2810
rect 6930 2800 6940 2810
rect 8120 2810 8200 2820
rect 8120 2800 8130 2810
rect 6930 2760 8130 2800
rect 6930 2750 6940 2760
rect 6860 2740 6940 2750
rect 8120 2750 8130 2760
rect 8190 2800 8200 2810
rect 9380 2810 9460 2820
rect 9380 2800 9390 2810
rect 8190 2760 9390 2800
rect 8190 2750 8200 2760
rect 8120 2740 8200 2750
rect 9380 2750 9390 2760
rect 9450 2800 9460 2810
rect 11330 2810 11410 2820
rect 11330 2800 11340 2810
rect 9450 2760 11340 2800
rect 9450 2750 9460 2760
rect 9380 2740 9460 2750
rect 11330 2750 11340 2760
rect 11400 2750 11410 2810
rect 11330 2740 11410 2750
rect 8120 2620 8200 2630
rect 8120 2560 8130 2620
rect 8190 2560 8200 2620
rect 8120 2550 8200 2560
rect 35520 2590 35600 2600
rect 35520 2530 35530 2590
rect 35590 2580 35600 2590
rect 35780 2590 35860 2600
rect 35780 2580 35790 2590
rect 35590 2540 35790 2580
rect 35590 2530 35600 2540
rect 35520 2520 35600 2530
rect 35780 2530 35790 2540
rect 35850 2580 35860 2590
rect 36240 2590 36320 2600
rect 36240 2580 36250 2590
rect 35850 2540 36250 2580
rect 35850 2530 35860 2540
rect 35780 2520 35860 2530
rect 36240 2530 36250 2540
rect 36310 2530 36320 2590
rect 36240 2520 36320 2530
rect 40450 2590 40530 2600
rect 40450 2530 40460 2590
rect 40520 2580 40530 2590
rect 40710 2590 40790 2600
rect 40710 2580 40720 2590
rect 40520 2540 40720 2580
rect 40520 2530 40530 2540
rect 40450 2520 40530 2530
rect 40710 2530 40720 2540
rect 40780 2580 40790 2590
rect 40780 2540 42200 2580
rect 40780 2530 40790 2540
rect 40710 2520 40790 2530
rect 6040 2510 6120 2520
rect 6040 2450 6050 2510
rect 6110 2500 6120 2510
rect 6200 2510 6280 2520
rect 6200 2500 6210 2510
rect 6110 2460 6210 2500
rect 6110 2450 6120 2460
rect 6040 2440 6120 2450
rect 6200 2450 6210 2460
rect 6270 2500 6280 2510
rect 6360 2510 6440 2520
rect 6360 2500 6370 2510
rect 6270 2460 6370 2500
rect 6270 2450 6280 2460
rect 6200 2440 6280 2450
rect 6360 2450 6370 2460
rect 6430 2500 6440 2510
rect 6520 2510 6600 2520
rect 6520 2500 6530 2510
rect 6430 2460 6530 2500
rect 6430 2450 6440 2460
rect 6360 2440 6440 2450
rect 6520 2450 6530 2460
rect 6590 2500 6600 2510
rect 6680 2510 6760 2520
rect 6680 2500 6690 2510
rect 6590 2460 6690 2500
rect 6590 2450 6600 2460
rect 6520 2440 6600 2450
rect 6680 2450 6690 2460
rect 6750 2500 6760 2510
rect 6840 2510 6920 2520
rect 6840 2500 6850 2510
rect 6750 2460 6850 2500
rect 6750 2450 6760 2460
rect 6680 2440 6760 2450
rect 6840 2450 6850 2460
rect 6910 2500 6920 2510
rect 7000 2510 7080 2520
rect 7000 2500 7010 2510
rect 6910 2460 7010 2500
rect 6910 2450 6920 2460
rect 6840 2440 6920 2450
rect 7000 2450 7010 2460
rect 7070 2500 7080 2510
rect 7160 2510 7240 2520
rect 7160 2500 7170 2510
rect 7070 2460 7170 2500
rect 7070 2450 7080 2460
rect 7000 2440 7080 2450
rect 7160 2450 7170 2460
rect 7230 2500 7240 2510
rect 7320 2510 7400 2520
rect 7320 2500 7330 2510
rect 7230 2460 7330 2500
rect 7230 2450 7240 2460
rect 7160 2440 7240 2450
rect 7320 2450 7330 2460
rect 7390 2500 7400 2510
rect 7480 2510 7560 2520
rect 7480 2500 7490 2510
rect 7390 2460 7490 2500
rect 7390 2450 7400 2460
rect 7320 2440 7400 2450
rect 7480 2450 7490 2460
rect 7550 2500 7560 2510
rect 7640 2510 7720 2520
rect 7640 2500 7650 2510
rect 7550 2460 7650 2500
rect 7550 2450 7560 2460
rect 7480 2440 7560 2450
rect 7640 2450 7650 2460
rect 7710 2500 7720 2510
rect 7800 2510 7880 2520
rect 7800 2500 7810 2510
rect 7710 2460 7810 2500
rect 7710 2450 7720 2460
rect 7640 2440 7720 2450
rect 7800 2450 7810 2460
rect 7870 2500 7880 2510
rect 7960 2510 8040 2520
rect 7960 2500 7970 2510
rect 7870 2460 7970 2500
rect 7870 2450 7880 2460
rect 7800 2440 7880 2450
rect 7960 2450 7970 2460
rect 8030 2450 8040 2510
rect 7960 2440 8040 2450
rect 8120 2510 8200 2520
rect 8120 2450 8130 2510
rect 8190 2500 8200 2510
rect 8280 2510 8360 2520
rect 8280 2500 8290 2510
rect 8190 2460 8290 2500
rect 8190 2450 8200 2460
rect 8120 2440 8200 2450
rect 8280 2450 8290 2460
rect 8350 2500 8360 2510
rect 8440 2510 8520 2520
rect 8440 2500 8450 2510
rect 8350 2460 8450 2500
rect 8350 2450 8360 2460
rect 8280 2440 8360 2450
rect 8440 2450 8450 2460
rect 8510 2500 8520 2510
rect 8600 2510 8680 2520
rect 8600 2500 8610 2510
rect 8510 2460 8610 2500
rect 8510 2450 8520 2460
rect 8440 2440 8520 2450
rect 8600 2450 8610 2460
rect 8670 2500 8680 2510
rect 8760 2510 8840 2520
rect 8760 2500 8770 2510
rect 8670 2460 8770 2500
rect 8670 2450 8680 2460
rect 8600 2440 8680 2450
rect 8760 2450 8770 2460
rect 8830 2500 8840 2510
rect 8920 2510 9000 2520
rect 8920 2500 8930 2510
rect 8830 2460 8930 2500
rect 8830 2450 8840 2460
rect 8760 2440 8840 2450
rect 8920 2450 8930 2460
rect 8990 2500 9000 2510
rect 9080 2510 9160 2520
rect 9080 2500 9090 2510
rect 8990 2460 9090 2500
rect 8990 2450 9000 2460
rect 8920 2440 9000 2450
rect 9080 2450 9090 2460
rect 9150 2500 9160 2510
rect 9240 2510 9320 2520
rect 9240 2500 9250 2510
rect 9150 2460 9250 2500
rect 9150 2450 9160 2460
rect 9080 2440 9160 2450
rect 9240 2450 9250 2460
rect 9310 2500 9320 2510
rect 9400 2510 9480 2520
rect 9400 2500 9410 2510
rect 9310 2460 9410 2500
rect 9310 2450 9320 2460
rect 9240 2440 9320 2450
rect 9400 2450 9410 2460
rect 9470 2500 9480 2510
rect 9560 2510 9640 2520
rect 9560 2500 9570 2510
rect 9470 2460 9570 2500
rect 9470 2450 9480 2460
rect 9400 2440 9480 2450
rect 9560 2450 9570 2460
rect 9630 2500 9640 2510
rect 9720 2510 9800 2520
rect 9720 2500 9730 2510
rect 9630 2460 9730 2500
rect 9630 2450 9640 2460
rect 9560 2440 9640 2450
rect 9720 2450 9730 2460
rect 9790 2500 9800 2510
rect 9880 2510 9960 2520
rect 9880 2500 9890 2510
rect 9790 2460 9890 2500
rect 9790 2450 9800 2460
rect 9720 2440 9800 2450
rect 9880 2450 9890 2460
rect 9950 2500 9960 2510
rect 10040 2510 10120 2520
rect 10040 2500 10050 2510
rect 9950 2460 10050 2500
rect 9950 2450 9960 2460
rect 9880 2440 9960 2450
rect 10040 2450 10050 2460
rect 10110 2450 10120 2510
rect 10040 2440 10120 2450
rect 34840 2390 34920 2400
rect 4550 2340 4630 2350
rect 4550 2280 4560 2340
rect 4620 2330 4630 2340
rect 5960 2340 6040 2350
rect 5960 2330 5970 2340
rect 4620 2290 5970 2330
rect 4620 2280 4630 2290
rect 4550 2270 4630 2280
rect 5960 2280 5970 2290
rect 6030 2280 6040 2340
rect 5960 2270 6040 2280
rect 10270 2340 10350 2350
rect 10270 2280 10280 2340
rect 10340 2330 10350 2340
rect 11330 2340 11410 2350
rect 11330 2330 11340 2340
rect 10340 2290 11340 2330
rect 10340 2280 10350 2290
rect 10270 2270 10350 2280
rect 11330 2280 11340 2290
rect 11400 2280 11410 2340
rect 34840 2330 34850 2390
rect 34910 2380 34920 2390
rect 37760 2390 37840 2400
rect 37760 2380 37770 2390
rect 34910 2340 37770 2380
rect 34910 2330 34920 2340
rect 34840 2320 34920 2330
rect 37760 2330 37770 2340
rect 37830 2380 37840 2390
rect 38480 2390 38560 2400
rect 38480 2380 38490 2390
rect 37830 2340 38490 2380
rect 37830 2330 37840 2340
rect 37760 2320 37840 2330
rect 38480 2330 38490 2340
rect 38550 2330 38560 2390
rect 38480 2320 38560 2330
rect 40120 2300 40200 2310
rect 11330 2270 11410 2280
rect 34660 2280 34740 2290
rect 34660 2220 34670 2280
rect 34730 2270 34740 2280
rect 36120 2280 36200 2290
rect 36120 2270 36130 2280
rect 34730 2230 36130 2270
rect 34730 2220 34740 2230
rect 34660 2210 34740 2220
rect 36120 2220 36130 2230
rect 36190 2270 36200 2280
rect 37400 2280 37480 2290
rect 37400 2270 37410 2280
rect 36190 2230 37410 2270
rect 36190 2220 36200 2230
rect 36120 2210 36200 2220
rect 37400 2220 37410 2230
rect 37470 2270 37480 2280
rect 38840 2280 38920 2290
rect 38840 2270 38850 2280
rect 37470 2230 38850 2270
rect 37470 2220 37480 2230
rect 37400 2210 37480 2220
rect 38840 2220 38850 2230
rect 38910 2220 38920 2280
rect 40120 2240 40130 2300
rect 40190 2290 40200 2300
rect 41050 2300 41130 2310
rect 41050 2290 41060 2300
rect 40190 2250 41060 2290
rect 40190 2240 40200 2250
rect 40120 2230 40200 2240
rect 41050 2240 41060 2250
rect 41120 2240 41130 2300
rect 41050 2230 41130 2240
rect 38840 2210 38920 2220
rect 34550 2190 34630 2200
rect 34550 2130 34560 2190
rect 34620 2180 34630 2190
rect 35650 2190 35730 2200
rect 35650 2180 35660 2190
rect 34620 2140 35660 2180
rect 34620 2130 34630 2140
rect 34550 2120 34630 2130
rect 35650 2130 35660 2140
rect 35720 2180 35730 2190
rect 37040 2190 37120 2200
rect 37040 2180 37050 2190
rect 35720 2140 37050 2180
rect 35720 2130 35730 2140
rect 35650 2120 35730 2130
rect 37040 2130 37050 2140
rect 37110 2180 37120 2190
rect 39200 2190 39280 2200
rect 39200 2180 39210 2190
rect 37110 2140 39210 2180
rect 37110 2130 37120 2140
rect 37040 2120 37120 2130
rect 39200 2130 39210 2140
rect 39270 2130 39280 2190
rect 39200 2120 39280 2130
rect 39380 2190 39460 2200
rect 39380 2130 39390 2190
rect 39450 2180 39460 2190
rect 40030 2190 40110 2200
rect 40030 2180 40040 2190
rect 39450 2140 40040 2180
rect 39450 2130 39460 2140
rect 39380 2120 39460 2130
rect 40030 2130 40040 2140
rect 40100 2130 40110 2190
rect 40030 2120 40110 2130
rect 6890 2100 6970 2110
rect 6890 2040 6900 2100
rect 6960 2090 6970 2100
rect 8120 2100 8200 2110
rect 8120 2090 8130 2100
rect 6960 2050 8130 2090
rect 6960 2040 6970 2050
rect 6890 2030 6970 2040
rect 8120 2040 8130 2050
rect 8190 2090 8200 2100
rect 9350 2100 9430 2110
rect 9350 2090 9360 2100
rect 8190 2050 9360 2090
rect 8190 2040 8200 2050
rect 8120 2030 8200 2040
rect 9350 2040 9360 2050
rect 9420 2040 9430 2100
rect 9350 2030 9430 2040
rect 35220 2100 35300 2110
rect 35220 2040 35230 2100
rect 35290 2090 35300 2100
rect 36680 2100 36760 2110
rect 36680 2090 36690 2100
rect 35290 2050 36690 2090
rect 35290 2040 35300 2050
rect 35220 2030 35300 2040
rect 36680 2040 36690 2050
rect 36750 2090 36760 2100
rect 38120 2100 38200 2110
rect 38120 2090 38130 2100
rect 36750 2050 38130 2090
rect 36750 2040 36760 2050
rect 36680 2030 36760 2040
rect 38120 2040 38130 2050
rect 38190 2090 38200 2100
rect 39560 2100 39640 2110
rect 39560 2090 39570 2100
rect 38190 2050 39570 2090
rect 38190 2040 38200 2050
rect 38120 2030 38200 2040
rect 39560 2040 39570 2050
rect 39630 2090 39640 2100
rect 41140 2100 41220 2110
rect 41140 2090 41150 2100
rect 39630 2050 41150 2090
rect 39630 2040 39640 2050
rect 39560 2030 39640 2040
rect 41140 2040 41150 2050
rect 41210 2040 41220 2100
rect 41140 2030 41220 2040
rect 34750 2000 34830 2010
rect 6560 1960 6640 1970
rect 6560 1900 6570 1960
rect 6630 1950 6640 1960
rect 6780 1960 6860 1970
rect 6780 1950 6790 1960
rect 6630 1910 6790 1950
rect 6630 1900 6640 1910
rect 6560 1890 6640 1900
rect 6780 1900 6790 1910
rect 6850 1950 6860 1960
rect 7000 1960 7080 1970
rect 7000 1950 7010 1960
rect 6850 1910 7010 1950
rect 6850 1900 6860 1910
rect 6780 1890 6860 1900
rect 7000 1900 7010 1910
rect 7070 1950 7080 1960
rect 7790 1960 7870 1970
rect 7790 1950 7800 1960
rect 7070 1910 7800 1950
rect 7070 1900 7080 1910
rect 7000 1890 7080 1900
rect 7790 1900 7800 1910
rect 7860 1950 7870 1960
rect 8010 1960 8090 1970
rect 8010 1950 8020 1960
rect 7860 1910 8020 1950
rect 7860 1900 7870 1910
rect 7790 1890 7870 1900
rect 8010 1900 8020 1910
rect 8080 1950 8090 1960
rect 8230 1960 8310 1970
rect 8230 1950 8240 1960
rect 8080 1910 8240 1950
rect 8080 1900 8090 1910
rect 8010 1890 8090 1900
rect 8230 1900 8240 1910
rect 8300 1950 8310 1960
rect 8450 1960 8530 1970
rect 8450 1950 8460 1960
rect 8300 1910 8460 1950
rect 8300 1900 8310 1910
rect 8230 1890 8310 1900
rect 8450 1900 8460 1910
rect 8520 1950 8530 1960
rect 9240 1960 9320 1970
rect 9240 1950 9250 1960
rect 8520 1910 9250 1950
rect 8520 1900 8530 1910
rect 8450 1890 8530 1900
rect 9240 1900 9250 1910
rect 9310 1950 9320 1960
rect 9460 1960 9540 1970
rect 9460 1950 9470 1960
rect 9310 1910 9470 1950
rect 9310 1900 9320 1910
rect 9240 1890 9320 1900
rect 9460 1900 9470 1910
rect 9530 1950 9540 1960
rect 9680 1960 9760 1970
rect 9680 1950 9690 1960
rect 9530 1910 9690 1950
rect 9530 1900 9540 1910
rect 9460 1890 9540 1900
rect 9680 1900 9690 1910
rect 9750 1950 9760 1960
rect 11330 1960 11410 1970
rect 11330 1950 11340 1960
rect 9750 1910 11340 1950
rect 9750 1900 9760 1910
rect 9680 1890 9760 1900
rect 11330 1900 11340 1910
rect 11400 1900 11410 1960
rect 34750 1940 34760 2000
rect 34820 1990 34830 2000
rect 38560 2000 38640 2010
rect 38560 1990 38570 2000
rect 34820 1950 38570 1990
rect 34820 1940 34830 1950
rect 34750 1930 34830 1940
rect 38560 1940 38570 1950
rect 38630 1990 38640 2000
rect 39940 2000 40020 2010
rect 39940 1990 39950 2000
rect 38630 1950 39950 1990
rect 38630 1940 38640 1950
rect 38560 1930 38640 1940
rect 39940 1940 39950 1950
rect 40010 1990 40020 2000
rect 40580 2000 40660 2010
rect 40580 1990 40590 2000
rect 40010 1950 40590 1990
rect 40010 1940 40020 1950
rect 39940 1930 40020 1940
rect 40580 1940 40590 1950
rect 40650 1940 40660 2000
rect 40580 1930 40660 1940
rect 11330 1890 11410 1900
rect 35640 1870 35720 1880
rect 35640 1810 35650 1870
rect 35710 1860 35720 1870
rect 35880 1870 35960 1880
rect 35880 1860 35890 1870
rect 35710 1820 35890 1860
rect 35710 1810 35720 1820
rect 35640 1800 35720 1810
rect 35880 1810 35890 1820
rect 35950 1860 35960 1870
rect 36120 1870 36200 1880
rect 36120 1860 36130 1870
rect 35950 1820 36130 1860
rect 35950 1810 35960 1820
rect 35880 1800 35960 1810
rect 36120 1810 36130 1820
rect 36190 1860 36200 1870
rect 36360 1870 36440 1880
rect 36360 1860 36370 1870
rect 36190 1820 36370 1860
rect 36190 1810 36200 1820
rect 36120 1800 36200 1810
rect 36360 1810 36370 1820
rect 36430 1860 36440 1870
rect 36600 1870 36680 1880
rect 36600 1860 36610 1870
rect 36430 1820 36610 1860
rect 36430 1810 36440 1820
rect 36360 1800 36440 1810
rect 36600 1810 36610 1820
rect 36670 1860 36680 1870
rect 36840 1870 36920 1880
rect 36840 1860 36850 1870
rect 36670 1820 36850 1860
rect 36670 1810 36680 1820
rect 36600 1800 36680 1810
rect 36840 1810 36850 1820
rect 36910 1860 36920 1870
rect 37080 1870 37160 1880
rect 37080 1860 37090 1870
rect 36910 1820 37090 1860
rect 36910 1810 36920 1820
rect 36840 1800 36920 1810
rect 37080 1810 37090 1820
rect 37150 1860 37160 1870
rect 37320 1870 37400 1880
rect 37320 1860 37330 1870
rect 37150 1820 37330 1860
rect 37150 1810 37160 1820
rect 37080 1800 37160 1810
rect 37320 1810 37330 1820
rect 37390 1860 37400 1870
rect 37560 1870 37640 1880
rect 37560 1860 37570 1870
rect 37390 1820 37570 1860
rect 37390 1810 37400 1820
rect 37320 1800 37400 1810
rect 37560 1810 37570 1820
rect 37630 1860 37640 1870
rect 38680 1870 38760 1880
rect 38680 1860 38690 1870
rect 37630 1820 38690 1860
rect 37630 1810 37640 1820
rect 37560 1800 37640 1810
rect 38680 1810 38690 1820
rect 38750 1860 38760 1870
rect 38920 1870 39000 1880
rect 38920 1860 38930 1870
rect 38750 1820 38930 1860
rect 38750 1810 38760 1820
rect 38680 1800 38760 1810
rect 38920 1810 38930 1820
rect 38990 1860 39000 1870
rect 39160 1870 39240 1880
rect 39160 1860 39170 1870
rect 38990 1820 39170 1860
rect 38990 1810 39000 1820
rect 38920 1800 39000 1810
rect 39160 1810 39170 1820
rect 39230 1860 39240 1870
rect 39400 1870 39480 1880
rect 39400 1860 39410 1870
rect 39230 1820 39410 1860
rect 39230 1810 39240 1820
rect 39160 1800 39240 1810
rect 39400 1810 39410 1820
rect 39470 1860 39480 1870
rect 39640 1870 39720 1880
rect 39640 1860 39650 1870
rect 39470 1820 39650 1860
rect 39470 1810 39480 1820
rect 39400 1800 39480 1810
rect 39640 1810 39650 1820
rect 39710 1860 39720 1870
rect 39880 1870 39960 1880
rect 39880 1860 39890 1870
rect 39710 1820 39890 1860
rect 39710 1810 39720 1820
rect 39640 1800 39720 1810
rect 39880 1810 39890 1820
rect 39950 1860 39960 1870
rect 40120 1870 40200 1880
rect 40120 1860 40130 1870
rect 39950 1820 40130 1860
rect 39950 1810 39960 1820
rect 39880 1800 39960 1810
rect 40120 1810 40130 1820
rect 40190 1860 40200 1870
rect 40360 1870 40440 1880
rect 40360 1860 40370 1870
rect 40190 1820 40370 1860
rect 40190 1810 40200 1820
rect 40120 1800 40200 1810
rect 40360 1810 40370 1820
rect 40430 1860 40440 1870
rect 40600 1870 40680 1880
rect 40600 1860 40610 1870
rect 40430 1820 40610 1860
rect 40430 1810 40440 1820
rect 40360 1800 40440 1810
rect 40600 1810 40610 1820
rect 40670 1860 40680 1870
rect 41500 1870 41580 1880
rect 41500 1860 41510 1870
rect 40670 1820 41510 1860
rect 40670 1810 40680 1820
rect 40600 1800 40680 1810
rect 41500 1810 41510 1820
rect 41570 1810 41580 1870
rect 41500 1800 41580 1810
rect 7340 1790 7420 1800
rect 7340 1730 7350 1790
rect 7410 1780 7420 1790
rect 7450 1790 7530 1800
rect 7450 1780 7460 1790
rect 7410 1740 7460 1780
rect 7410 1730 7420 1740
rect 7340 1720 7420 1730
rect 7450 1730 7460 1740
rect 7520 1730 7530 1790
rect 7450 1720 7530 1730
rect 8790 1790 8870 1800
rect 8790 1730 8800 1790
rect 8860 1780 8870 1790
rect 8900 1790 8980 1800
rect 8900 1780 8910 1790
rect 8860 1740 8910 1780
rect 8860 1730 8870 1740
rect 8790 1720 8870 1730
rect 8900 1730 8910 1740
rect 8970 1730 8980 1790
rect 8900 1720 8980 1730
rect 10020 1790 10100 1800
rect 10020 1730 10030 1790
rect 10090 1780 10100 1790
rect 11330 1790 11410 1800
rect 11330 1780 11340 1790
rect 10090 1740 11340 1780
rect 10090 1730 10100 1740
rect 10020 1720 10100 1730
rect 11330 1730 11340 1740
rect 11400 1730 11410 1790
rect 11330 1720 11410 1730
rect 34930 1750 35010 1760
rect 34930 1690 34940 1750
rect 35000 1740 35010 1750
rect 35520 1750 35600 1760
rect 35520 1740 35530 1750
rect 35000 1700 35530 1740
rect 35000 1690 35010 1700
rect 34930 1680 35010 1690
rect 35520 1690 35530 1700
rect 35590 1740 35600 1750
rect 36240 1750 36320 1760
rect 36240 1740 36250 1750
rect 35590 1700 36250 1740
rect 35590 1690 35600 1700
rect 35520 1680 35600 1690
rect 36240 1690 36250 1700
rect 36310 1740 36320 1750
rect 36960 1750 37040 1760
rect 36960 1740 36970 1750
rect 36310 1700 36970 1740
rect 36310 1690 36320 1700
rect 36240 1680 36320 1690
rect 36960 1690 36970 1700
rect 37030 1740 37040 1750
rect 37680 1750 37760 1760
rect 37680 1740 37690 1750
rect 37030 1700 37690 1740
rect 37030 1690 37040 1700
rect 36960 1680 37040 1690
rect 37680 1690 37690 1700
rect 37750 1740 37760 1750
rect 37940 1750 38020 1760
rect 37940 1740 37950 1750
rect 37750 1700 37950 1740
rect 37750 1690 37760 1700
rect 37680 1680 37760 1690
rect 37940 1690 37950 1700
rect 38010 1690 38020 1750
rect 37940 1680 38020 1690
rect 38300 1750 38380 1760
rect 38300 1690 38310 1750
rect 38370 1740 38380 1750
rect 38560 1750 38640 1760
rect 38560 1740 38570 1750
rect 38370 1700 38570 1740
rect 38370 1690 38380 1700
rect 38300 1680 38380 1690
rect 38560 1690 38570 1700
rect 38630 1740 38640 1750
rect 39280 1750 39360 1760
rect 39280 1740 39290 1750
rect 38630 1700 39290 1740
rect 38630 1690 38640 1700
rect 38560 1680 38640 1690
rect 39280 1690 39290 1700
rect 39350 1740 39360 1750
rect 40000 1750 40080 1760
rect 40000 1740 40010 1750
rect 39350 1700 40010 1740
rect 39350 1690 39360 1700
rect 39280 1680 39360 1690
rect 40000 1690 40010 1700
rect 40070 1740 40080 1750
rect 40720 1750 40800 1760
rect 40720 1740 40730 1750
rect 40070 1700 40730 1740
rect 40070 1690 40080 1700
rect 40000 1680 40080 1690
rect 40720 1690 40730 1700
rect 40790 1690 40800 1750
rect 40720 1680 40800 1690
rect 6450 1620 6530 1630
rect 6450 1560 6460 1620
rect 6520 1610 6530 1620
rect 6670 1620 6750 1630
rect 6670 1610 6680 1620
rect 6520 1570 6680 1610
rect 6520 1560 6530 1570
rect 6450 1550 6530 1560
rect 6670 1560 6680 1570
rect 6740 1610 6750 1620
rect 6890 1620 6970 1630
rect 6890 1610 6900 1620
rect 6740 1570 6900 1610
rect 6740 1560 6750 1570
rect 6670 1550 6750 1560
rect 6890 1560 6900 1570
rect 6960 1610 6970 1620
rect 7110 1620 7190 1630
rect 7110 1610 7120 1620
rect 6960 1570 7120 1610
rect 6960 1560 6970 1570
rect 6890 1550 6970 1560
rect 7110 1560 7120 1570
rect 7180 1560 7190 1620
rect 7110 1550 7190 1560
rect 8120 1620 8200 1630
rect 8120 1560 8130 1620
rect 8190 1610 8200 1620
rect 8340 1620 8420 1630
rect 8340 1610 8350 1620
rect 8190 1570 8350 1610
rect 8190 1560 8200 1570
rect 8120 1550 8200 1560
rect 8340 1560 8350 1570
rect 8410 1610 8420 1620
rect 8560 1620 8640 1630
rect 8560 1610 8570 1620
rect 8410 1570 8570 1610
rect 8410 1560 8420 1570
rect 8340 1550 8420 1560
rect 8560 1560 8570 1570
rect 8630 1560 8640 1620
rect 8560 1550 8640 1560
rect 9130 1620 9210 1630
rect 9130 1560 9140 1620
rect 9200 1610 9210 1620
rect 9570 1620 9650 1630
rect 9570 1610 9580 1620
rect 9200 1570 9580 1610
rect 9200 1560 9210 1570
rect 9130 1550 9210 1560
rect 9570 1560 9580 1570
rect 9640 1560 9650 1620
rect 9570 1550 9650 1560
rect 9350 1510 9430 1520
rect 9350 1450 9360 1510
rect 9420 1500 9430 1510
rect 9790 1510 9870 1520
rect 9790 1500 9800 1510
rect 9420 1460 9800 1500
rect 9420 1450 9430 1460
rect 9350 1440 9430 1450
rect 9790 1450 9800 1460
rect 9860 1450 9870 1510
rect 9790 1440 9870 1450
rect 5110 1420 5190 1430
rect 5110 1360 5120 1420
rect 5180 1410 5190 1420
rect 7730 1420 7810 1430
rect 7730 1410 7740 1420
rect 5180 1370 7740 1410
rect 5180 1360 5190 1370
rect 5110 1350 5190 1360
rect 7730 1360 7740 1370
rect 7800 1360 7810 1420
rect 7730 1350 7810 1360
rect 35760 1410 35840 1420
rect 35760 1350 35770 1410
rect 35830 1400 35840 1410
rect 36000 1400 36080 1420
rect 36480 1410 36560 1420
rect 36480 1400 36490 1410
rect 35830 1360 36490 1400
rect 35830 1350 35840 1360
rect 35760 1340 35840 1350
rect 36000 1340 36080 1360
rect 36480 1350 36490 1360
rect 36550 1400 36560 1410
rect 36720 1400 36800 1420
rect 37200 1410 37280 1420
rect 37200 1400 37210 1410
rect 36550 1360 37210 1400
rect 36550 1350 36560 1360
rect 36480 1340 36560 1350
rect 36720 1340 36800 1360
rect 37200 1350 37210 1360
rect 37270 1350 37280 1410
rect 37200 1340 37280 1350
rect 37440 1340 37520 1420
rect 38800 1340 38880 1420
rect 39040 1410 39120 1420
rect 39040 1350 39050 1410
rect 39110 1400 39120 1410
rect 39520 1400 39600 1420
rect 39760 1410 39840 1420
rect 39760 1400 39770 1410
rect 39110 1360 39770 1400
rect 39110 1350 39120 1360
rect 39040 1340 39120 1350
rect 39520 1340 39600 1360
rect 39760 1350 39770 1360
rect 39830 1400 39840 1410
rect 40240 1400 40320 1420
rect 40480 1410 40560 1420
rect 40480 1400 40490 1410
rect 39830 1360 40490 1400
rect 39830 1350 39840 1360
rect 39760 1340 39840 1350
rect 40240 1340 40320 1360
rect 40480 1350 40490 1360
rect 40550 1350 40560 1410
rect 40480 1340 40560 1350
rect 35020 1290 35100 1300
rect 35020 1230 35030 1290
rect 35090 1280 35100 1290
rect 35580 1290 35660 1300
rect 35580 1280 35590 1290
rect 35090 1240 35590 1280
rect 35090 1230 35100 1240
rect 35020 1220 35100 1230
rect 35580 1230 35590 1240
rect 35650 1280 35660 1290
rect 36000 1290 36080 1300
rect 36000 1280 36010 1290
rect 35650 1240 36010 1280
rect 35650 1230 35660 1240
rect 35580 1220 35660 1230
rect 36000 1230 36010 1240
rect 36070 1280 36080 1290
rect 36240 1290 36320 1300
rect 36240 1280 36250 1290
rect 36070 1240 36250 1280
rect 36070 1230 36080 1240
rect 36000 1220 36080 1230
rect 36240 1230 36250 1240
rect 36310 1280 36320 1290
rect 36720 1290 36800 1300
rect 36720 1280 36730 1290
rect 36310 1240 36730 1280
rect 36310 1230 36320 1240
rect 36240 1220 36320 1230
rect 36720 1230 36730 1240
rect 36790 1280 36800 1290
rect 36960 1290 37040 1300
rect 36960 1280 36970 1290
rect 36790 1240 36970 1280
rect 36790 1230 36800 1240
rect 36720 1220 36800 1230
rect 36960 1230 36970 1240
rect 37030 1280 37040 1290
rect 37440 1290 37520 1300
rect 37440 1280 37450 1290
rect 37030 1240 37450 1280
rect 37030 1230 37040 1240
rect 36960 1220 37040 1230
rect 37440 1230 37450 1240
rect 37510 1280 37520 1290
rect 37620 1290 37700 1300
rect 37620 1280 37630 1290
rect 37510 1240 37630 1280
rect 37510 1230 37520 1240
rect 37440 1220 37520 1230
rect 37620 1230 37630 1240
rect 37690 1230 37700 1290
rect 37620 1220 37700 1230
rect 38620 1290 38700 1300
rect 38620 1230 38630 1290
rect 38690 1280 38700 1290
rect 38800 1290 38880 1300
rect 38800 1280 38810 1290
rect 38690 1240 38810 1280
rect 38690 1230 38700 1240
rect 38620 1220 38700 1230
rect 38800 1230 38810 1240
rect 38870 1280 38880 1290
rect 39280 1290 39360 1300
rect 39280 1280 39290 1290
rect 38870 1240 39290 1280
rect 38870 1230 38880 1240
rect 38800 1220 38880 1230
rect 39280 1230 39290 1240
rect 39350 1280 39360 1290
rect 39520 1290 39600 1300
rect 39520 1280 39530 1290
rect 39350 1240 39530 1280
rect 39350 1230 39360 1240
rect 39280 1220 39360 1230
rect 39520 1230 39530 1240
rect 39590 1280 39600 1290
rect 40000 1290 40080 1300
rect 40000 1280 40010 1290
rect 39590 1240 40010 1280
rect 39590 1230 39600 1240
rect 39520 1220 39600 1230
rect 40000 1230 40010 1240
rect 40070 1280 40080 1290
rect 40240 1290 40320 1300
rect 40240 1280 40250 1290
rect 40070 1240 40250 1280
rect 40070 1230 40080 1240
rect 40000 1220 40080 1230
rect 40240 1230 40250 1240
rect 40310 1280 40320 1290
rect 40660 1290 40740 1300
rect 40660 1280 40670 1290
rect 40310 1240 40670 1280
rect 40310 1230 40320 1240
rect 40240 1220 40320 1230
rect 40660 1230 40670 1240
rect 40730 1280 40740 1290
rect 41050 1290 41130 1300
rect 41050 1280 41060 1290
rect 40730 1240 41060 1280
rect 40730 1230 40740 1240
rect 40660 1220 40740 1230
rect 41050 1230 41060 1240
rect 41120 1230 41130 1290
rect 41050 1220 41130 1230
rect 36500 1120 36580 1130
rect 34660 1090 34740 1100
rect 34660 1030 34670 1090
rect 34730 1080 34740 1090
rect 36380 1090 36460 1100
rect 36380 1080 36390 1090
rect 34730 1040 36390 1080
rect 34730 1030 34740 1040
rect 34660 1020 34740 1030
rect 36380 1030 36390 1040
rect 36450 1030 36460 1090
rect 36500 1060 36510 1120
rect 36570 1110 36580 1120
rect 36980 1120 37060 1130
rect 36980 1110 36990 1120
rect 36570 1070 36990 1110
rect 36570 1060 36580 1070
rect 36500 1050 36580 1060
rect 36980 1060 36990 1070
rect 37050 1110 37060 1120
rect 37460 1120 37540 1130
rect 37460 1110 37470 1120
rect 37050 1070 37470 1110
rect 37050 1060 37060 1070
rect 36980 1050 37060 1060
rect 37460 1060 37470 1070
rect 37530 1060 37540 1120
rect 37460 1050 37540 1060
rect 38780 1120 38860 1130
rect 38780 1060 38790 1120
rect 38850 1110 38860 1120
rect 39260 1120 39340 1130
rect 39260 1110 39270 1120
rect 38850 1070 39270 1110
rect 38850 1060 38860 1070
rect 38780 1050 38860 1060
rect 39260 1060 39270 1070
rect 39330 1110 39340 1120
rect 39740 1120 39820 1130
rect 39740 1110 39750 1120
rect 39330 1070 39750 1110
rect 39330 1060 39340 1070
rect 39260 1050 39340 1060
rect 39740 1060 39750 1070
rect 39810 1060 39820 1120
rect 39740 1050 39820 1060
rect 39860 1090 39940 1100
rect 36380 1020 36460 1030
rect 39860 1030 39870 1090
rect 39930 1080 39940 1090
rect 41140 1090 41220 1100
rect 41140 1080 41150 1090
rect 39930 1040 41150 1080
rect 39930 1030 39940 1040
rect 39860 1020 39940 1030
rect 41140 1030 41150 1040
rect 41210 1080 41220 1090
rect 41210 1040 42200 1080
rect 41210 1030 41220 1040
rect 41140 1020 41220 1030
rect 36260 1000 36340 1010
rect 36260 940 36270 1000
rect 36330 990 36340 1000
rect 36740 1000 36820 1010
rect 36740 990 36750 1000
rect 36330 950 36750 990
rect 36330 940 36340 950
rect 36260 930 36340 940
rect 36740 940 36750 950
rect 36810 990 36820 1000
rect 37220 1000 37300 1010
rect 37220 990 37230 1000
rect 36810 950 37230 990
rect 36810 940 36820 950
rect 36740 930 36820 940
rect 37220 940 37230 950
rect 37290 940 37300 1000
rect 37220 930 37300 940
rect 39020 1000 39100 1010
rect 39020 940 39030 1000
rect 39090 990 39100 1000
rect 39500 1000 39580 1010
rect 39500 990 39510 1000
rect 39090 950 39510 990
rect 39090 940 39100 950
rect 39020 930 39100 940
rect 39500 940 39510 950
rect 39570 990 39580 1000
rect 39980 1000 40060 1010
rect 39980 990 39990 1000
rect 39570 950 39990 990
rect 39570 940 39580 950
rect 39500 930 39580 940
rect 39980 940 39990 950
rect 40050 940 40060 1000
rect 39980 930 40060 940
rect 37580 880 37660 890
rect 37580 820 37590 880
rect 37650 870 37660 880
rect 38120 880 38200 890
rect 38120 870 38130 880
rect 37650 830 38130 870
rect 37650 820 37660 830
rect 37580 810 37660 820
rect 38120 820 38130 830
rect 38190 870 38200 880
rect 38660 880 38740 890
rect 38660 870 38670 880
rect 38190 830 38670 870
rect 38190 820 38200 830
rect 38120 810 38200 820
rect 38660 820 38670 830
rect 38730 820 38740 880
rect 38660 810 38740 820
rect 34840 760 34920 770
rect 34840 700 34850 760
rect 34910 750 34920 760
rect 36260 760 36340 770
rect 36260 750 36270 760
rect 34910 710 36270 750
rect 34910 700 34920 710
rect 34840 690 34920 700
rect 36260 700 36270 710
rect 36330 700 36340 760
rect 36260 690 36340 700
rect 39980 760 40060 770
rect 39980 700 39990 760
rect 40050 750 40060 760
rect 41230 760 41310 770
rect 41230 750 41240 760
rect 40050 710 41240 750
rect 40050 700 40060 710
rect 39980 690 40060 700
rect 41230 700 41240 710
rect 41300 700 41310 760
rect 41230 690 41310 700
rect 35780 640 35860 650
rect 35780 580 35790 640
rect 35850 630 35860 640
rect 36380 640 36460 650
rect 36380 630 36390 640
rect 35850 590 36390 630
rect 35850 580 35860 590
rect 35780 570 35860 580
rect 36380 580 36390 590
rect 36450 630 36460 640
rect 36620 640 36700 650
rect 36620 630 36630 640
rect 36450 590 36630 630
rect 36450 580 36460 590
rect 36380 570 36460 580
rect 36620 580 36630 590
rect 36690 630 36700 640
rect 36860 640 36940 650
rect 36860 630 36870 640
rect 36690 590 36870 630
rect 36690 580 36700 590
rect 36620 570 36700 580
rect 36860 580 36870 590
rect 36930 630 36940 640
rect 37100 640 37180 650
rect 37100 630 37110 640
rect 36930 590 37110 630
rect 36930 580 36940 590
rect 36860 570 36940 580
rect 37100 580 37110 590
rect 37170 630 37180 640
rect 37340 640 37420 650
rect 37340 630 37350 640
rect 37170 590 37350 630
rect 37170 580 37180 590
rect 37100 570 37180 580
rect 37340 580 37350 590
rect 37410 580 37420 640
rect 37340 570 37420 580
rect 38900 640 38980 650
rect 38900 580 38910 640
rect 38970 630 38980 640
rect 39140 640 39220 650
rect 39140 630 39150 640
rect 38970 590 39150 630
rect 38970 580 38980 590
rect 38900 570 38980 580
rect 39140 580 39150 590
rect 39210 630 39220 640
rect 39380 640 39460 650
rect 39380 630 39390 640
rect 39210 590 39390 630
rect 39210 580 39220 590
rect 39140 570 39220 580
rect 39380 580 39390 590
rect 39450 630 39460 640
rect 39620 640 39700 650
rect 39620 630 39630 640
rect 39450 590 39630 630
rect 39450 580 39460 590
rect 39380 570 39460 580
rect 39620 580 39630 590
rect 39690 630 39700 640
rect 39860 640 39940 650
rect 39860 630 39870 640
rect 39690 590 39870 630
rect 39690 580 39700 590
rect 39620 570 39700 580
rect 39860 580 39870 590
rect 39930 630 39940 640
rect 40460 640 40540 650
rect 40460 630 40470 640
rect 39930 590 40470 630
rect 39930 580 39940 590
rect 39860 570 39940 580
rect 40460 580 40470 590
rect 40530 580 40540 640
rect 40460 570 40540 580
rect 35960 440 36040 450
rect 34660 420 34740 430
rect 34660 410 34670 420
rect 34500 370 34670 410
rect 34660 360 34670 370
rect 34730 360 34740 420
rect 35960 380 35970 440
rect 36030 430 36040 440
rect 36200 440 36280 450
rect 36200 430 36210 440
rect 36030 390 36210 430
rect 36030 380 36040 390
rect 35960 370 36040 380
rect 36200 380 36210 390
rect 36270 430 36280 440
rect 36440 440 36520 450
rect 36440 430 36450 440
rect 36270 390 36450 430
rect 36270 380 36280 390
rect 36200 370 36280 380
rect 36440 380 36450 390
rect 36510 430 36520 440
rect 36680 440 36760 450
rect 36680 430 36690 440
rect 36510 390 36690 430
rect 36510 380 36520 390
rect 36440 370 36520 380
rect 36680 380 36690 390
rect 36750 430 36760 440
rect 37160 440 37240 450
rect 37160 430 37170 440
rect 36750 390 37170 430
rect 36750 380 36760 390
rect 36680 370 36760 380
rect 37160 380 37170 390
rect 37230 430 37240 440
rect 37400 440 37480 450
rect 37400 430 37410 440
rect 37230 390 37410 430
rect 37230 380 37240 390
rect 37160 370 37240 380
rect 37400 380 37410 390
rect 37470 430 37480 440
rect 37640 440 37720 450
rect 37640 430 37650 440
rect 37470 390 37650 430
rect 37470 380 37480 390
rect 37400 370 37480 380
rect 37640 380 37650 390
rect 37710 430 37720 440
rect 38600 440 38680 450
rect 38600 430 38610 440
rect 37710 390 38610 430
rect 37710 380 37720 390
rect 37640 370 37720 380
rect 38600 380 38610 390
rect 38670 430 38680 440
rect 38840 440 38920 450
rect 38840 430 38850 440
rect 38670 390 38850 430
rect 38670 380 38680 390
rect 38600 370 38680 380
rect 38840 380 38850 390
rect 38910 430 38920 440
rect 39080 440 39160 450
rect 39080 430 39090 440
rect 38910 390 39090 430
rect 38910 380 38920 390
rect 38840 370 38920 380
rect 39080 380 39090 390
rect 39150 430 39160 440
rect 39560 440 39640 450
rect 39560 430 39570 440
rect 39150 390 39570 430
rect 39150 380 39160 390
rect 39080 370 39160 380
rect 39560 380 39570 390
rect 39630 430 39640 440
rect 39800 440 39880 450
rect 39800 430 39810 440
rect 39630 390 39810 430
rect 39630 380 39640 390
rect 39560 370 39640 380
rect 39800 380 39810 390
rect 39870 430 39880 440
rect 40040 440 40120 450
rect 40040 430 40050 440
rect 39870 390 40050 430
rect 39870 380 39880 390
rect 39800 370 39880 380
rect 40040 380 40050 390
rect 40110 430 40120 440
rect 40280 440 40360 450
rect 40280 430 40290 440
rect 40110 390 40290 430
rect 40110 380 40120 390
rect 40040 370 40120 380
rect 40280 380 40290 390
rect 40350 430 40360 440
rect 41500 440 41580 450
rect 41500 430 41510 440
rect 40350 390 41510 430
rect 40350 380 40360 390
rect 40280 370 40360 380
rect 41500 380 41510 390
rect 41570 380 41580 440
rect 41500 370 41580 380
rect 34660 350 34740 360
rect 36860 -190 36940 -180
rect 36860 -250 36870 -190
rect 36930 -200 36940 -190
rect 38120 -190 38200 -180
rect 38120 -200 38130 -190
rect 36930 -240 38130 -200
rect 36930 -250 36940 -240
rect 36860 -260 36940 -250
rect 38120 -250 38130 -240
rect 38190 -200 38200 -190
rect 39380 -190 39460 -180
rect 39380 -200 39390 -190
rect 38190 -240 39390 -200
rect 38190 -250 38200 -240
rect 38120 -260 38200 -250
rect 39380 -250 39390 -240
rect 39450 -200 39460 -190
rect 41330 -190 41410 -180
rect 41330 -200 41340 -190
rect 39450 -240 41340 -200
rect 39450 -250 39460 -240
rect 39380 -260 39460 -250
rect 41330 -250 41340 -240
rect 41400 -250 41410 -190
rect 41330 -260 41410 -250
rect 38120 -380 38200 -370
rect 38120 -440 38130 -380
rect 38190 -440 38200 -380
rect 38120 -450 38200 -440
rect 36040 -490 36120 -480
rect 36040 -550 36050 -490
rect 36110 -500 36120 -490
rect 36200 -490 36280 -480
rect 36200 -500 36210 -490
rect 36110 -540 36210 -500
rect 36110 -550 36120 -540
rect 36040 -560 36120 -550
rect 36200 -550 36210 -540
rect 36270 -500 36280 -490
rect 36360 -490 36440 -480
rect 36360 -500 36370 -490
rect 36270 -540 36370 -500
rect 36270 -550 36280 -540
rect 36200 -560 36280 -550
rect 36360 -550 36370 -540
rect 36430 -500 36440 -490
rect 36520 -490 36600 -480
rect 36520 -500 36530 -490
rect 36430 -540 36530 -500
rect 36430 -550 36440 -540
rect 36360 -560 36440 -550
rect 36520 -550 36530 -540
rect 36590 -500 36600 -490
rect 36680 -490 36760 -480
rect 36680 -500 36690 -490
rect 36590 -540 36690 -500
rect 36590 -550 36600 -540
rect 36520 -560 36600 -550
rect 36680 -550 36690 -540
rect 36750 -500 36760 -490
rect 36840 -490 36920 -480
rect 36840 -500 36850 -490
rect 36750 -540 36850 -500
rect 36750 -550 36760 -540
rect 36680 -560 36760 -550
rect 36840 -550 36850 -540
rect 36910 -500 36920 -490
rect 37000 -490 37080 -480
rect 37000 -500 37010 -490
rect 36910 -540 37010 -500
rect 36910 -550 36920 -540
rect 36840 -560 36920 -550
rect 37000 -550 37010 -540
rect 37070 -500 37080 -490
rect 37160 -490 37240 -480
rect 37160 -500 37170 -490
rect 37070 -540 37170 -500
rect 37070 -550 37080 -540
rect 37000 -560 37080 -550
rect 37160 -550 37170 -540
rect 37230 -500 37240 -490
rect 37320 -490 37400 -480
rect 37320 -500 37330 -490
rect 37230 -540 37330 -500
rect 37230 -550 37240 -540
rect 37160 -560 37240 -550
rect 37320 -550 37330 -540
rect 37390 -500 37400 -490
rect 37480 -490 37560 -480
rect 37480 -500 37490 -490
rect 37390 -540 37490 -500
rect 37390 -550 37400 -540
rect 37320 -560 37400 -550
rect 37480 -550 37490 -540
rect 37550 -500 37560 -490
rect 37640 -490 37720 -480
rect 37640 -500 37650 -490
rect 37550 -540 37650 -500
rect 37550 -550 37560 -540
rect 37480 -560 37560 -550
rect 37640 -550 37650 -540
rect 37710 -500 37720 -490
rect 37800 -490 37880 -480
rect 37800 -500 37810 -490
rect 37710 -540 37810 -500
rect 37710 -550 37720 -540
rect 37640 -560 37720 -550
rect 37800 -550 37810 -540
rect 37870 -500 37880 -490
rect 37960 -490 38040 -480
rect 37960 -500 37970 -490
rect 37870 -540 37970 -500
rect 37870 -550 37880 -540
rect 37800 -560 37880 -550
rect 37960 -550 37970 -540
rect 38030 -550 38040 -490
rect 37960 -560 38040 -550
rect 38120 -490 38200 -480
rect 38120 -550 38130 -490
rect 38190 -500 38200 -490
rect 38280 -490 38360 -480
rect 38280 -500 38290 -490
rect 38190 -540 38290 -500
rect 38190 -550 38200 -540
rect 38120 -560 38200 -550
rect 38280 -550 38290 -540
rect 38350 -500 38360 -490
rect 38440 -490 38520 -480
rect 38440 -500 38450 -490
rect 38350 -540 38450 -500
rect 38350 -550 38360 -540
rect 38280 -560 38360 -550
rect 38440 -550 38450 -540
rect 38510 -500 38520 -490
rect 38600 -490 38680 -480
rect 38600 -500 38610 -490
rect 38510 -540 38610 -500
rect 38510 -550 38520 -540
rect 38440 -560 38520 -550
rect 38600 -550 38610 -540
rect 38670 -500 38680 -490
rect 38760 -490 38840 -480
rect 38760 -500 38770 -490
rect 38670 -540 38770 -500
rect 38670 -550 38680 -540
rect 38600 -560 38680 -550
rect 38760 -550 38770 -540
rect 38830 -500 38840 -490
rect 38920 -490 39000 -480
rect 38920 -500 38930 -490
rect 38830 -540 38930 -500
rect 38830 -550 38840 -540
rect 38760 -560 38840 -550
rect 38920 -550 38930 -540
rect 38990 -500 39000 -490
rect 39080 -490 39160 -480
rect 39080 -500 39090 -490
rect 38990 -540 39090 -500
rect 38990 -550 39000 -540
rect 38920 -560 39000 -550
rect 39080 -550 39090 -540
rect 39150 -500 39160 -490
rect 39240 -490 39320 -480
rect 39240 -500 39250 -490
rect 39150 -540 39250 -500
rect 39150 -550 39160 -540
rect 39080 -560 39160 -550
rect 39240 -550 39250 -540
rect 39310 -500 39320 -490
rect 39400 -490 39480 -480
rect 39400 -500 39410 -490
rect 39310 -540 39410 -500
rect 39310 -550 39320 -540
rect 39240 -560 39320 -550
rect 39400 -550 39410 -540
rect 39470 -500 39480 -490
rect 39560 -490 39640 -480
rect 39560 -500 39570 -490
rect 39470 -540 39570 -500
rect 39470 -550 39480 -540
rect 39400 -560 39480 -550
rect 39560 -550 39570 -540
rect 39630 -500 39640 -490
rect 39720 -490 39800 -480
rect 39720 -500 39730 -490
rect 39630 -540 39730 -500
rect 39630 -550 39640 -540
rect 39560 -560 39640 -550
rect 39720 -550 39730 -540
rect 39790 -500 39800 -490
rect 39880 -490 39960 -480
rect 39880 -500 39890 -490
rect 39790 -540 39890 -500
rect 39790 -550 39800 -540
rect 39720 -560 39800 -550
rect 39880 -550 39890 -540
rect 39950 -500 39960 -490
rect 40040 -490 40120 -480
rect 40040 -500 40050 -490
rect 39950 -540 40050 -500
rect 39950 -550 39960 -540
rect 39880 -560 39960 -550
rect 40040 -550 40050 -540
rect 40110 -550 40120 -490
rect 40040 -560 40120 -550
rect 34550 -660 34630 -650
rect 34550 -720 34560 -660
rect 34620 -670 34630 -660
rect 35960 -660 36040 -650
rect 35960 -670 35970 -660
rect 34620 -710 35970 -670
rect 34620 -720 34630 -710
rect 34550 -730 34630 -720
rect 35960 -720 35970 -710
rect 36030 -720 36040 -660
rect 35960 -730 36040 -720
rect 40270 -660 40350 -650
rect 40270 -720 40280 -660
rect 40340 -670 40350 -660
rect 41330 -660 41410 -650
rect 41330 -670 41340 -660
rect 40340 -710 41340 -670
rect 40340 -720 40350 -710
rect 40270 -730 40350 -720
rect 41330 -720 41340 -710
rect 41400 -720 41410 -660
rect 41330 -730 41410 -720
rect 36890 -900 36970 -890
rect 36890 -960 36900 -900
rect 36960 -910 36970 -900
rect 38120 -900 38200 -890
rect 38120 -910 38130 -900
rect 36960 -950 38130 -910
rect 36960 -960 36970 -950
rect 36890 -970 36970 -960
rect 38120 -960 38130 -950
rect 38190 -910 38200 -900
rect 39350 -900 39430 -890
rect 39350 -910 39360 -900
rect 38190 -950 39360 -910
rect 38190 -960 38200 -950
rect 38120 -970 38200 -960
rect 39350 -960 39360 -950
rect 39420 -960 39430 -900
rect 39350 -970 39430 -960
rect 36560 -1040 36640 -1030
rect 36560 -1100 36570 -1040
rect 36630 -1050 36640 -1040
rect 36780 -1040 36860 -1030
rect 36780 -1050 36790 -1040
rect 36630 -1090 36790 -1050
rect 36630 -1100 36640 -1090
rect 36560 -1110 36640 -1100
rect 36780 -1100 36790 -1090
rect 36850 -1050 36860 -1040
rect 37000 -1040 37080 -1030
rect 37000 -1050 37010 -1040
rect 36850 -1090 37010 -1050
rect 36850 -1100 36860 -1090
rect 36780 -1110 36860 -1100
rect 37000 -1100 37010 -1090
rect 37070 -1050 37080 -1040
rect 37790 -1040 37870 -1030
rect 37790 -1050 37800 -1040
rect 37070 -1090 37800 -1050
rect 37070 -1100 37080 -1090
rect 37000 -1110 37080 -1100
rect 37790 -1100 37800 -1090
rect 37860 -1050 37870 -1040
rect 38010 -1040 38090 -1030
rect 38010 -1050 38020 -1040
rect 37860 -1090 38020 -1050
rect 37860 -1100 37870 -1090
rect 37790 -1110 37870 -1100
rect 38010 -1100 38020 -1090
rect 38080 -1050 38090 -1040
rect 38230 -1040 38310 -1030
rect 38230 -1050 38240 -1040
rect 38080 -1090 38240 -1050
rect 38080 -1100 38090 -1090
rect 38010 -1110 38090 -1100
rect 38230 -1100 38240 -1090
rect 38300 -1050 38310 -1040
rect 38450 -1040 38530 -1030
rect 38450 -1050 38460 -1040
rect 38300 -1090 38460 -1050
rect 38300 -1100 38310 -1090
rect 38230 -1110 38310 -1100
rect 38450 -1100 38460 -1090
rect 38520 -1050 38530 -1040
rect 39240 -1040 39320 -1030
rect 39240 -1050 39250 -1040
rect 38520 -1090 39250 -1050
rect 38520 -1100 38530 -1090
rect 38450 -1110 38530 -1100
rect 39240 -1100 39250 -1090
rect 39310 -1050 39320 -1040
rect 39460 -1040 39540 -1030
rect 39460 -1050 39470 -1040
rect 39310 -1090 39470 -1050
rect 39310 -1100 39320 -1090
rect 39240 -1110 39320 -1100
rect 39460 -1100 39470 -1090
rect 39530 -1050 39540 -1040
rect 39680 -1040 39760 -1030
rect 39680 -1050 39690 -1040
rect 39530 -1090 39690 -1050
rect 39530 -1100 39540 -1090
rect 39460 -1110 39540 -1100
rect 39680 -1100 39690 -1090
rect 39750 -1050 39760 -1040
rect 41330 -1040 41410 -1030
rect 41330 -1050 41340 -1040
rect 39750 -1090 41340 -1050
rect 39750 -1100 39760 -1090
rect 39680 -1110 39760 -1100
rect 41330 -1100 41340 -1090
rect 41400 -1100 41410 -1040
rect 41330 -1110 41410 -1100
rect 37340 -1210 37420 -1200
rect 37340 -1270 37350 -1210
rect 37410 -1220 37420 -1210
rect 37450 -1210 37530 -1200
rect 37450 -1220 37460 -1210
rect 37410 -1260 37460 -1220
rect 37410 -1270 37420 -1260
rect 37340 -1280 37420 -1270
rect 37450 -1270 37460 -1260
rect 37520 -1270 37530 -1210
rect 37450 -1280 37530 -1270
rect 38790 -1210 38870 -1200
rect 38790 -1270 38800 -1210
rect 38860 -1220 38870 -1210
rect 38900 -1210 38980 -1200
rect 38900 -1220 38910 -1210
rect 38860 -1260 38910 -1220
rect 38860 -1270 38870 -1260
rect 38790 -1280 38870 -1270
rect 38900 -1270 38910 -1260
rect 38970 -1270 38980 -1210
rect 38900 -1280 38980 -1270
rect 40020 -1210 40100 -1200
rect 40020 -1270 40030 -1210
rect 40090 -1220 40100 -1210
rect 41330 -1210 41410 -1200
rect 41330 -1220 41340 -1210
rect 40090 -1260 41340 -1220
rect 40090 -1270 40100 -1260
rect 40020 -1280 40100 -1270
rect 41330 -1270 41340 -1260
rect 41400 -1270 41410 -1210
rect 41330 -1280 41410 -1270
rect 36450 -1380 36530 -1370
rect 36450 -1440 36460 -1380
rect 36520 -1390 36530 -1380
rect 36670 -1380 36750 -1370
rect 36670 -1390 36680 -1380
rect 36520 -1430 36680 -1390
rect 36520 -1440 36530 -1430
rect 36450 -1450 36530 -1440
rect 36670 -1440 36680 -1430
rect 36740 -1390 36750 -1380
rect 36890 -1380 36970 -1370
rect 36890 -1390 36900 -1380
rect 36740 -1430 36900 -1390
rect 36740 -1440 36750 -1430
rect 36670 -1450 36750 -1440
rect 36890 -1440 36900 -1430
rect 36960 -1390 36970 -1380
rect 37110 -1380 37190 -1370
rect 37110 -1390 37120 -1380
rect 36960 -1430 37120 -1390
rect 36960 -1440 36970 -1430
rect 36890 -1450 36970 -1440
rect 37110 -1440 37120 -1430
rect 37180 -1440 37190 -1380
rect 37110 -1450 37190 -1440
rect 38120 -1380 38200 -1370
rect 38120 -1440 38130 -1380
rect 38190 -1390 38200 -1380
rect 38340 -1380 38420 -1370
rect 38340 -1390 38350 -1380
rect 38190 -1430 38350 -1390
rect 38190 -1440 38200 -1430
rect 38120 -1450 38200 -1440
rect 38340 -1440 38350 -1430
rect 38410 -1390 38420 -1380
rect 38560 -1380 38640 -1370
rect 38560 -1390 38570 -1380
rect 38410 -1430 38570 -1390
rect 38410 -1440 38420 -1430
rect 38340 -1450 38420 -1440
rect 38560 -1440 38570 -1430
rect 38630 -1440 38640 -1380
rect 38560 -1450 38640 -1440
rect 39130 -1380 39210 -1370
rect 39130 -1440 39140 -1380
rect 39200 -1390 39210 -1380
rect 39570 -1380 39650 -1370
rect 39570 -1390 39580 -1380
rect 39200 -1430 39580 -1390
rect 39200 -1440 39210 -1430
rect 39130 -1450 39210 -1440
rect 39570 -1440 39580 -1430
rect 39640 -1440 39650 -1380
rect 39570 -1450 39650 -1440
rect 39350 -1490 39430 -1480
rect 39350 -1550 39360 -1490
rect 39420 -1500 39430 -1490
rect 39790 -1490 39870 -1480
rect 39790 -1500 39800 -1490
rect 39420 -1540 39800 -1500
rect 39420 -1550 39430 -1540
rect 39350 -1560 39430 -1550
rect 39790 -1550 39800 -1540
rect 39860 -1550 39870 -1490
rect 39790 -1560 39870 -1550
rect 35110 -1580 35190 -1570
rect 35110 -1640 35120 -1580
rect 35180 -1590 35190 -1580
rect 37730 -1580 37810 -1570
rect 37730 -1590 37740 -1580
rect 35180 -1630 37740 -1590
rect 35180 -1640 35190 -1630
rect 35110 -1650 35190 -1640
rect 37730 -1640 37740 -1630
rect 37800 -1640 37810 -1580
rect 37730 -1650 37810 -1640
rect 46510 -2620 46590 -2610
rect 46510 -2680 46520 -2620
rect 46580 -2630 46590 -2620
rect 46580 -2670 49250 -2630
rect 46580 -2680 46590 -2670
rect 46510 -2690 46590 -2680
rect 44140 -2720 44220 -2710
rect 44140 -2780 44150 -2720
rect 44210 -2730 44220 -2720
rect 49110 -2720 49190 -2710
rect 49110 -2730 49120 -2720
rect 44210 -2770 49120 -2730
rect 44210 -2780 44220 -2770
rect 44140 -2790 44220 -2780
rect 49110 -2780 49120 -2770
rect 49180 -2780 49190 -2720
rect 49110 -2790 49190 -2780
rect 44132 -2890 44142 -2820
rect 44212 -2890 44222 -2820
rect 43780 -2950 43860 -2940
rect 43780 -3010 43790 -2950
rect 43850 -2960 43860 -2950
rect 44132 -2960 44142 -2940
rect 43850 -3000 44142 -2960
rect 43850 -3010 43860 -3000
rect 44132 -3010 44142 -3000
rect 44212 -3010 44222 -2940
rect 43780 -3020 43860 -3010
rect 46702 -3160 46712 -3090
rect 46782 -3160 46792 -3090
rect 44140 -3250 44220 -3240
rect 44140 -3310 44150 -3250
rect 44210 -3260 44220 -3250
rect 46510 -3250 46590 -3240
rect 46510 -3260 46520 -3250
rect 44210 -3300 46520 -3260
rect 44210 -3310 44220 -3300
rect 44140 -3320 44220 -3310
rect 46510 -3310 46520 -3300
rect 46580 -3310 46590 -3250
rect 46702 -3280 46712 -3210
rect 46782 -3280 46792 -3210
rect 46510 -3320 46590 -3310
rect 44132 -3420 44142 -3350
rect 44212 -3420 44222 -3350
rect 46370 -3420 46450 -3410
rect 43780 -3480 43860 -3470
rect 43780 -3540 43790 -3480
rect 43850 -3490 43860 -3480
rect 44132 -3490 44142 -3470
rect 43850 -3530 44142 -3490
rect 43850 -3540 43860 -3530
rect 44132 -3540 44142 -3530
rect 44212 -3540 44222 -3470
rect 46370 -3480 46380 -3420
rect 46440 -3430 46450 -3420
rect 46580 -3420 46660 -3410
rect 46580 -3430 46590 -3420
rect 46440 -3470 46590 -3430
rect 46440 -3480 46450 -3470
rect 46370 -3490 46450 -3480
rect 46580 -3480 46590 -3470
rect 46650 -3480 46660 -3420
rect 46580 -3490 46660 -3480
rect 49110 -3490 49190 -3480
rect 43780 -3550 43860 -3540
rect 49110 -3550 49120 -3490
rect 49180 -3500 49190 -3490
rect 49220 -3490 49250 -3480
rect 49220 -3500 49230 -3490
rect 49180 -3540 49230 -3500
rect 49180 -3550 49190 -3540
rect 49110 -3560 49190 -3550
rect 49220 -3550 49230 -3540
rect 49220 -3560 49250 -3550
rect 43780 -3610 43860 -3600
rect 43780 -3670 43790 -3610
rect 43850 -3620 43860 -3610
rect 45190 -3610 45270 -3600
rect 45190 -3620 45200 -3610
rect 43850 -3660 45200 -3620
rect 43850 -3670 43860 -3660
rect 43780 -3680 43860 -3670
rect 45190 -3670 45200 -3660
rect 45260 -3670 45270 -3610
rect 48840 -3640 48850 -3570
rect 48920 -3590 48930 -3570
rect 48920 -3630 49250 -3590
rect 48920 -3640 48930 -3630
rect 45190 -3680 45270 -3670
rect 49110 -3670 49190 -3660
rect 48840 -3690 48930 -3680
rect 48840 -3760 48850 -3690
rect 48920 -3760 48930 -3690
rect 49110 -3730 49120 -3670
rect 49180 -3680 49190 -3670
rect 49180 -3720 49250 -3680
rect 49180 -3730 49190 -3720
rect 49110 -3740 49190 -3730
rect 48840 -3770 48930 -3760
rect 43880 -3890 43960 -3880
rect 43880 -3950 43890 -3890
rect 43950 -3900 43960 -3890
rect 44522 -3900 44532 -3880
rect 43950 -3940 44532 -3900
rect 43950 -3950 43960 -3940
rect 44522 -3950 44532 -3940
rect 44602 -3950 44612 -3880
rect 45868 -3950 45878 -3880
rect 45948 -3900 45958 -3880
rect 46420 -3890 46500 -3880
rect 46420 -3900 46430 -3890
rect 45948 -3940 46430 -3900
rect 45948 -3950 45958 -3940
rect 46420 -3950 46430 -3940
rect 46490 -3950 46500 -3890
rect 43880 -3960 43960 -3950
rect 46420 -3960 46500 -3950
rect 46210 -4100 46290 -4090
rect 35600 -5906 35640 -4140
rect 46210 -4160 46220 -4100
rect 46280 -4110 46290 -4100
rect 47032 -4110 47042 -4100
rect 46280 -4150 47042 -4110
rect 46280 -4160 46290 -4150
rect 46210 -4170 46290 -4160
rect 47032 -4170 47042 -4150
rect 47112 -4170 47122 -4100
rect 48430 -4170 48440 -4100
rect 48510 -4120 48520 -4100
rect 48840 -4110 48920 -4100
rect 48840 -4120 48850 -4110
rect 48510 -4160 48850 -4120
rect 48510 -4170 48520 -4160
rect 48840 -4170 48850 -4160
rect 48910 -4170 48920 -4110
rect 48840 -4180 48920 -4170
rect 43970 -4300 44050 -4290
rect 43970 -4360 43980 -4300
rect 44040 -4320 44050 -4300
rect 44522 -4320 44532 -4300
rect 44040 -4360 44532 -4320
rect 43970 -4370 44050 -4360
rect 44522 -4370 44532 -4360
rect 44602 -4370 44612 -4300
rect 45868 -4370 45878 -4300
rect 45948 -4320 45958 -4300
rect 48930 -4310 49010 -4300
rect 48930 -4320 48940 -4310
rect 45948 -4360 48940 -4320
rect 45948 -4370 45958 -4360
rect 48930 -4370 48940 -4360
rect 49000 -4370 49010 -4310
rect 48930 -4380 49010 -4370
rect 46420 -4400 46500 -4390
rect 46420 -4460 46430 -4400
rect 46490 -4410 46500 -4400
rect 48750 -4400 48830 -4390
rect 48750 -4410 48760 -4400
rect 46490 -4450 48760 -4410
rect 46490 -4460 46500 -4450
rect 46420 -4470 46500 -4460
rect 48750 -4460 48760 -4450
rect 48820 -4460 48830 -4400
rect 48750 -4470 48830 -4460
rect 35580 -5916 35660 -5906
rect 35580 -5970 35590 -5916
rect 35650 -5970 35660 -5916
rect 35580 -5986 35660 -5970
rect 29780 -6560 29860 -6550
rect 29780 -6620 29790 -6560
rect 29850 -6620 29860 -6560
rect 29780 -6630 29860 -6620
rect 35560 -8530 35640 -8520
rect 35560 -8590 35570 -8530
rect 35630 -8590 35640 -8530
rect 35560 -8600 35640 -8590
<< via2 >>
rect -210 7690 -150 7750
rect 8890 7630 8950 7690
rect 11510 7630 11570 7690
rect 29790 7690 29850 7750
rect 38890 7630 38950 7690
rect 41510 7630 41570 7690
rect 1890 7530 1950 7590
rect 3290 7530 3350 7590
rect 10290 7530 10350 7590
rect 31890 7530 31950 7590
rect 33290 7530 33350 7590
rect 40290 7530 40350 7590
rect 5390 7420 5450 7480
rect 6790 7420 6850 7480
rect 35390 7420 35450 7480
rect 36790 7420 36850 7480
rect -210 6990 -150 7050
rect 11510 7000 11570 7060
rect -210 6460 -150 6520
rect -210 6330 -150 6390
rect 11510 6070 11570 6130
rect 11510 4810 11570 4870
rect 41510 4000 41570 4060
rect -210 3380 -150 3440
rect 11510 3380 11570 3440
rect 41510 3070 41570 3130
rect 11340 2750 11400 2810
rect 11340 2280 11400 2340
rect 11340 1900 11400 1960
rect 41510 1810 41570 1870
rect 11340 1730 11400 1790
rect 41510 380 41570 440
rect 41340 -250 41400 -190
rect 41340 -720 41400 -660
rect 41340 -1100 41400 -1040
rect 41340 -1270 41400 -1210
rect 43790 -3010 43850 -2950
rect 43790 -3540 43850 -3480
rect 43790 -3670 43850 -3610
rect 29790 -6620 29850 -6560
<< metal3 >>
rect -400 10690 -300 10700
rect -400 10610 -390 10690
rect -310 10610 -300 10690
rect -400 10600 -300 10610
rect 11490 10690 11590 10700
rect 11490 10610 11500 10690
rect 11580 10610 11590 10690
rect 11490 10600 11590 10610
rect 29600 10690 29700 10700
rect 29600 10610 29610 10690
rect 29690 10610 29700 10690
rect 29600 10600 29700 10610
rect 41490 10690 41590 10700
rect 41490 10610 41500 10690
rect 41580 10610 41590 10690
rect 41490 10600 41590 10610
rect -390 1170 -310 10600
rect -230 10520 -130 10530
rect -230 10440 -220 10520
rect -140 10440 -130 10520
rect -230 10430 -130 10440
rect 11320 10520 11420 10530
rect 11320 10440 11330 10520
rect 11410 10440 11420 10520
rect 11320 10430 11420 10440
rect -220 7750 -140 10430
rect 290 10240 750 10410
rect 990 10240 1450 10410
rect 1690 10240 2150 10410
rect 2390 10240 2850 10410
rect 3090 10240 3550 10410
rect 290 10140 3550 10240
rect 290 9950 750 10140
rect 990 9950 1450 10140
rect 1690 9950 2150 10140
rect 2390 9950 2850 10140
rect 3090 9950 3550 10140
rect 3790 10240 4250 10410
rect 4490 10240 4950 10410
rect 5190 10240 5650 10410
rect 5890 10240 6350 10410
rect 6590 10240 7050 10410
rect 3790 10140 7050 10240
rect 3790 9950 4250 10140
rect 4490 9950 4950 10140
rect 5190 9950 5650 10140
rect 5890 9950 6350 10140
rect 6590 9950 7050 10140
rect 7290 10240 7750 10410
rect 7990 10240 8450 10410
rect 8690 10240 9150 10410
rect 9390 10240 9850 10410
rect 10090 10240 10550 10410
rect 7290 10140 10550 10240
rect 7290 9950 7750 10140
rect 7990 9950 8450 10140
rect 8690 9950 9150 10140
rect 9390 9950 9850 10140
rect 10090 9950 10550 10140
rect 1870 9710 1970 9950
rect 5370 9710 5470 9950
rect 8870 9710 8970 9950
rect 290 9540 750 9710
rect 990 9540 1450 9710
rect 1690 9540 2150 9710
rect 2390 9540 2850 9710
rect 3090 9540 3550 9710
rect 290 9440 3550 9540
rect 290 9250 750 9440
rect 990 9250 1450 9440
rect 1690 9250 2150 9440
rect 2390 9250 2850 9440
rect 3090 9250 3550 9440
rect 3790 9540 4250 9710
rect 4490 9540 4950 9710
rect 5190 9540 5650 9710
rect 5890 9540 6350 9710
rect 6590 9540 7050 9710
rect 3790 9440 7050 9540
rect 3790 9250 4250 9440
rect 4490 9250 4950 9440
rect 5190 9250 5650 9440
rect 5890 9250 6350 9440
rect 6590 9250 7050 9440
rect 7290 9540 7750 9710
rect 7990 9540 8450 9710
rect 8690 9540 9150 9710
rect 9390 9540 9850 9710
rect 10090 9540 10550 9710
rect 7290 9440 10550 9540
rect 7290 9250 7750 9440
rect 7990 9250 8450 9440
rect 8690 9250 9150 9440
rect 9390 9250 9850 9440
rect 10090 9250 10550 9440
rect 1870 9010 1970 9250
rect 5370 9010 5470 9250
rect 8870 9010 8970 9250
rect 290 8840 750 9010
rect 990 8840 1450 9010
rect 1690 8840 2150 9010
rect 2390 8840 2850 9010
rect 3090 8840 3550 9010
rect 290 8740 3550 8840
rect 290 8550 750 8740
rect 990 8550 1450 8740
rect 1690 8550 2150 8740
rect 2390 8550 2850 8740
rect 3090 8550 3550 8740
rect 3790 8840 4250 9010
rect 4490 8840 4950 9010
rect 5190 8840 5650 9010
rect 5890 8840 6350 9010
rect 6590 8840 7050 9010
rect 3790 8740 7050 8840
rect 3790 8550 4250 8740
rect 4490 8550 4950 8740
rect 5190 8550 5650 8740
rect 5890 8550 6350 8740
rect 6590 8550 7050 8740
rect 7290 8840 7750 9010
rect 7990 8840 8450 9010
rect 8690 8840 9150 9010
rect 9390 8840 9850 9010
rect 10090 8840 10550 9010
rect 7290 8740 10550 8840
rect 7290 8550 7750 8740
rect 7990 8550 8450 8740
rect 8690 8550 9150 8740
rect 9390 8550 9850 8740
rect 10090 8550 10550 8740
rect 1870 8310 1970 8550
rect 5370 8310 5470 8550
rect 8870 8310 8970 8550
rect 290 8140 750 8310
rect 990 8140 1450 8310
rect 1690 8140 2150 8310
rect 2390 8140 2850 8310
rect 3090 8140 3550 8310
rect 290 8040 3550 8140
rect 290 7850 750 8040
rect 990 7850 1450 8040
rect 1690 7850 2150 8040
rect 2390 7850 2850 8040
rect 3090 7850 3550 8040
rect 3790 8140 4250 8310
rect 4490 8140 4950 8310
rect 5190 8140 5650 8310
rect 5890 8140 6350 8310
rect 6590 8140 7050 8310
rect 3790 8040 7050 8140
rect 3790 7850 4250 8040
rect 4490 7850 4950 8040
rect 5190 7850 5650 8040
rect 5890 7850 6350 8040
rect 6590 7850 7050 8040
rect 7290 8140 7750 8310
rect 7990 8140 8450 8310
rect 8690 8140 9150 8310
rect 9390 8140 9850 8310
rect 10090 8140 10550 8310
rect 7290 8040 10550 8140
rect 7290 7850 7750 8040
rect 7990 7850 8450 8040
rect 8690 7850 9150 8040
rect 9390 7850 9850 8040
rect 10090 7850 10550 8040
rect -220 7690 -210 7750
rect -150 7690 -140 7750
rect -220 7050 -140 7690
rect 1880 7590 1960 7850
rect 1880 7530 1890 7590
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect 3270 7600 3370 7610
rect 3270 7520 3280 7600
rect 3360 7520 3370 7600
rect 3270 7510 3370 7520
rect 5380 7480 5460 7850
rect 8880 7690 8960 7850
rect 8880 7630 8890 7690
rect 8950 7630 8960 7690
rect 8880 7620 8960 7630
rect 10270 7600 10370 7610
rect 10270 7520 10280 7600
rect 10360 7520 10370 7600
rect 10270 7510 10370 7520
rect 5380 7420 5390 7480
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7490 6870 7500
rect 6770 7410 6780 7490
rect 6860 7410 6870 7490
rect 6770 7400 6870 7410
rect -220 6990 -210 7050
rect -150 6990 -140 7050
rect -220 6520 -140 6990
rect -220 6460 -210 6520
rect -150 6460 -140 6520
rect -220 6390 -140 6460
rect -220 6330 -210 6390
rect -150 6330 -140 6390
rect -220 3440 -140 6330
rect -220 3380 -210 3440
rect -150 3380 -140 3440
rect -220 1330 -140 3380
rect 11330 2810 11410 10430
rect 11330 2750 11340 2810
rect 11400 2750 11410 2810
rect 11330 2340 11410 2750
rect 11330 2280 11340 2340
rect 11400 2280 11410 2340
rect 11330 1960 11410 2280
rect 11330 1900 11340 1960
rect 11400 1900 11410 1960
rect 11330 1790 11410 1900
rect 11330 1730 11340 1790
rect 11400 1730 11410 1790
rect 11330 1330 11410 1730
rect 11500 7690 11580 10600
rect 11500 7630 11510 7690
rect 11570 7630 11580 7690
rect 11500 7060 11580 7630
rect 11500 7000 11510 7060
rect 11570 7000 11580 7060
rect 11500 6130 11580 7000
rect 11500 6070 11510 6130
rect 11570 6070 11580 6130
rect 11500 4870 11580 6070
rect 11500 4810 11510 4870
rect 11570 4810 11580 4870
rect 11500 3440 11580 4810
rect 11500 3380 11510 3440
rect 11570 3380 11580 3440
rect -230 1320 -130 1330
rect -230 1240 -220 1320
rect -140 1240 -130 1320
rect -230 1230 -130 1240
rect 11320 1320 11420 1330
rect 11320 1240 11330 1320
rect 11410 1240 11420 1320
rect 11320 1230 11420 1240
rect 11500 1170 11580 3380
rect -400 1160 -300 1170
rect -400 1080 -390 1160
rect -310 1080 -300 1160
rect -400 1070 -300 1080
rect 11490 1160 11590 1170
rect 11490 1080 11500 1160
rect 11580 1080 11590 1160
rect 11490 1070 11590 1080
rect 29610 -8830 29690 10600
rect 29770 10520 29870 10530
rect 29770 10440 29780 10520
rect 29860 10440 29870 10520
rect 29770 10430 29870 10440
rect 41320 10520 41420 10530
rect 41320 10440 41330 10520
rect 41410 10440 41420 10520
rect 41320 10430 41420 10440
rect 29780 7750 29860 10430
rect 30290 10240 30750 10410
rect 30990 10240 31450 10410
rect 31690 10240 32150 10410
rect 32390 10240 32850 10410
rect 33090 10240 33550 10410
rect 30290 10140 33550 10240
rect 30290 9950 30750 10140
rect 30990 9950 31450 10140
rect 31690 9950 32150 10140
rect 32390 9950 32850 10140
rect 33090 9950 33550 10140
rect 33790 10240 34250 10410
rect 34490 10240 34950 10410
rect 35190 10240 35650 10410
rect 35890 10240 36350 10410
rect 36590 10240 37050 10410
rect 33790 10140 37050 10240
rect 33790 9950 34250 10140
rect 34490 9950 34950 10140
rect 35190 9950 35650 10140
rect 35890 9950 36350 10140
rect 36590 9950 37050 10140
rect 37290 10240 37750 10410
rect 37990 10240 38450 10410
rect 38690 10240 39150 10410
rect 39390 10240 39850 10410
rect 40090 10240 40550 10410
rect 37290 10140 40550 10240
rect 37290 9950 37750 10140
rect 37990 9950 38450 10140
rect 38690 9950 39150 10140
rect 39390 9950 39850 10140
rect 40090 9950 40550 10140
rect 31870 9710 31970 9950
rect 35370 9710 35470 9950
rect 38870 9710 38970 9950
rect 30290 9540 30750 9710
rect 30990 9540 31450 9710
rect 31690 9540 32150 9710
rect 32390 9540 32850 9710
rect 33090 9540 33550 9710
rect 30290 9440 33550 9540
rect 30290 9250 30750 9440
rect 30990 9250 31450 9440
rect 31690 9250 32150 9440
rect 32390 9250 32850 9440
rect 33090 9250 33550 9440
rect 33790 9540 34250 9710
rect 34490 9540 34950 9710
rect 35190 9540 35650 9710
rect 35890 9540 36350 9710
rect 36590 9540 37050 9710
rect 33790 9440 37050 9540
rect 33790 9250 34250 9440
rect 34490 9250 34950 9440
rect 35190 9250 35650 9440
rect 35890 9250 36350 9440
rect 36590 9250 37050 9440
rect 37290 9540 37750 9710
rect 37990 9540 38450 9710
rect 38690 9540 39150 9710
rect 39390 9540 39850 9710
rect 40090 9540 40550 9710
rect 37290 9440 40550 9540
rect 37290 9250 37750 9440
rect 37990 9250 38450 9440
rect 38690 9250 39150 9440
rect 39390 9250 39850 9440
rect 40090 9250 40550 9440
rect 31870 9010 31970 9250
rect 35370 9010 35470 9250
rect 38870 9010 38970 9250
rect 30290 8840 30750 9010
rect 30990 8840 31450 9010
rect 31690 8840 32150 9010
rect 32390 8840 32850 9010
rect 33090 8840 33550 9010
rect 30290 8740 33550 8840
rect 30290 8550 30750 8740
rect 30990 8550 31450 8740
rect 31690 8550 32150 8740
rect 32390 8550 32850 8740
rect 33090 8550 33550 8740
rect 33790 8840 34250 9010
rect 34490 8840 34950 9010
rect 35190 8840 35650 9010
rect 35890 8840 36350 9010
rect 36590 8840 37050 9010
rect 33790 8740 37050 8840
rect 33790 8550 34250 8740
rect 34490 8550 34950 8740
rect 35190 8550 35650 8740
rect 35890 8550 36350 8740
rect 36590 8550 37050 8740
rect 37290 8840 37750 9010
rect 37990 8840 38450 9010
rect 38690 8840 39150 9010
rect 39390 8840 39850 9010
rect 40090 8840 40550 9010
rect 37290 8740 40550 8840
rect 37290 8550 37750 8740
rect 37990 8550 38450 8740
rect 38690 8550 39150 8740
rect 39390 8550 39850 8740
rect 40090 8550 40550 8740
rect 31870 8310 31970 8550
rect 35370 8310 35470 8550
rect 38870 8310 38970 8550
rect 30290 8140 30750 8310
rect 30990 8140 31450 8310
rect 31690 8140 32150 8310
rect 32390 8140 32850 8310
rect 33090 8140 33550 8310
rect 30290 8040 33550 8140
rect 30290 7850 30750 8040
rect 30990 7850 31450 8040
rect 31690 7850 32150 8040
rect 32390 7850 32850 8040
rect 33090 7850 33550 8040
rect 33790 8140 34250 8310
rect 34490 8140 34950 8310
rect 35190 8140 35650 8310
rect 35890 8140 36350 8310
rect 36590 8140 37050 8310
rect 33790 8040 37050 8140
rect 33790 7850 34250 8040
rect 34490 7850 34950 8040
rect 35190 7850 35650 8040
rect 35890 7850 36350 8040
rect 36590 7850 37050 8040
rect 37290 8140 37750 8310
rect 37990 8140 38450 8310
rect 38690 8140 39150 8310
rect 39390 8140 39850 8310
rect 40090 8140 40550 8310
rect 37290 8040 40550 8140
rect 37290 7850 37750 8040
rect 37990 7850 38450 8040
rect 38690 7850 39150 8040
rect 39390 7850 39850 8040
rect 40090 7850 40550 8040
rect 29780 7690 29790 7750
rect 29850 7690 29860 7750
rect 29780 -6560 29860 7690
rect 31880 7590 31960 7850
rect 31880 7530 31890 7590
rect 31950 7530 31960 7590
rect 31880 7520 31960 7530
rect 33270 7600 33370 7610
rect 33270 7520 33280 7600
rect 33360 7520 33370 7600
rect 33270 7510 33370 7520
rect 35380 7480 35460 7850
rect 38880 7690 38960 7850
rect 38880 7630 38890 7690
rect 38950 7630 38960 7690
rect 38880 7620 38960 7630
rect 40270 7600 40370 7610
rect 40270 7520 40280 7600
rect 40360 7520 40370 7600
rect 40270 7510 40370 7520
rect 35380 7420 35390 7480
rect 35450 7420 35460 7480
rect 35380 7410 35460 7420
rect 36770 7490 36870 7500
rect 36770 7410 36780 7490
rect 36860 7410 36870 7490
rect 36770 7400 36870 7410
rect 29780 -6620 29790 -6560
rect 29850 -6620 29860 -6560
rect 29780 -8670 29860 -6620
rect 41330 -190 41410 10430
rect 41330 -250 41340 -190
rect 41400 -250 41410 -190
rect 41330 -660 41410 -250
rect 41330 -720 41340 -660
rect 41400 -720 41410 -660
rect 41330 -1040 41410 -720
rect 41330 -1100 41340 -1040
rect 41400 -1100 41410 -1040
rect 41330 -1210 41410 -1100
rect 41330 -1270 41340 -1210
rect 41400 -1270 41410 -1210
rect 41330 -8670 41410 -1270
rect 41500 7690 41580 10600
rect 41500 7630 41510 7690
rect 41570 7630 41580 7690
rect 41500 4060 41580 7630
rect 41500 4000 41510 4060
rect 41570 4000 41580 4060
rect 41500 3130 41580 4000
rect 41500 3070 41510 3130
rect 41570 3070 41580 3130
rect 41500 1870 41580 3070
rect 41500 1810 41510 1870
rect 41570 1810 41580 1870
rect 41500 440 41580 1810
rect 41500 380 41510 440
rect 41570 380 41580 440
rect 29770 -8680 29870 -8670
rect 29770 -8760 29780 -8680
rect 29860 -8760 29870 -8680
rect 29770 -8770 29870 -8760
rect 41320 -8680 41420 -8670
rect 41320 -8760 41330 -8680
rect 41410 -8760 41420 -8680
rect 41320 -8770 41420 -8760
rect 41500 -8830 41580 380
rect 43780 -2950 43860 -2550
rect 43780 -3010 43790 -2950
rect 43850 -3010 43860 -2950
rect 43780 -3480 43860 -3010
rect 43780 -3540 43790 -3480
rect 43850 -3540 43860 -3480
rect 43780 -3610 43860 -3540
rect 43780 -3670 43790 -3610
rect 43850 -3670 43860 -3610
rect 43780 -4550 43860 -3670
rect 29600 -8840 29700 -8830
rect 29600 -8920 29610 -8840
rect 29690 -8920 29700 -8840
rect 29600 -8930 29700 -8920
rect 41490 -8840 41590 -8830
rect 41490 -8920 41500 -8840
rect 41580 -8920 41590 -8840
rect 41490 -8930 41590 -8920
<< via3 >>
rect -390 10610 -310 10690
rect 11500 10610 11580 10690
rect 29610 10610 29690 10690
rect 41500 10610 41580 10690
rect -220 10440 -140 10520
rect 11330 10440 11410 10520
rect 3280 7590 3360 7600
rect 3280 7530 3290 7590
rect 3290 7530 3350 7590
rect 3350 7530 3360 7590
rect 3280 7520 3360 7530
rect 10280 7590 10360 7600
rect 10280 7530 10290 7590
rect 10290 7530 10350 7590
rect 10350 7530 10360 7590
rect 10280 7520 10360 7530
rect 6780 7480 6860 7490
rect 6780 7420 6790 7480
rect 6790 7420 6850 7480
rect 6850 7420 6860 7480
rect 6780 7410 6860 7420
rect -220 1240 -140 1320
rect 11330 1240 11410 1320
rect -390 1080 -310 1160
rect 11500 1080 11580 1160
rect 29780 10440 29860 10520
rect 41330 10440 41410 10520
rect 33280 7590 33360 7600
rect 33280 7530 33290 7590
rect 33290 7530 33350 7590
rect 33350 7530 33360 7590
rect 33280 7520 33360 7530
rect 40280 7590 40360 7600
rect 40280 7530 40290 7590
rect 40290 7530 40350 7590
rect 40350 7530 40360 7590
rect 40280 7520 40360 7530
rect 36780 7480 36860 7490
rect 36780 7420 36790 7480
rect 36790 7420 36850 7480
rect 36850 7420 36860 7480
rect 36780 7410 36860 7420
rect 29780 -8760 29860 -8680
rect 41330 -8760 41410 -8680
rect 29610 -8920 29690 -8840
rect 41500 -8920 41580 -8840
<< mimcap >>
rect 320 10230 720 10380
rect 320 10150 480 10230
rect 560 10150 720 10230
rect 320 9980 720 10150
rect 1020 10230 1420 10380
rect 1020 10150 1180 10230
rect 1260 10150 1420 10230
rect 1020 9980 1420 10150
rect 1720 10230 2120 10380
rect 1720 10150 1880 10230
rect 1960 10150 2120 10230
rect 1720 9980 2120 10150
rect 2420 10230 2820 10380
rect 2420 10150 2580 10230
rect 2660 10150 2820 10230
rect 2420 9980 2820 10150
rect 3120 10230 3520 10380
rect 3120 10150 3280 10230
rect 3360 10150 3520 10230
rect 3120 9980 3520 10150
rect 3820 10230 4220 10380
rect 3820 10150 3980 10230
rect 4060 10150 4220 10230
rect 3820 9980 4220 10150
rect 4520 10230 4920 10380
rect 4520 10150 4680 10230
rect 4760 10150 4920 10230
rect 4520 9980 4920 10150
rect 5220 10230 5620 10380
rect 5220 10150 5380 10230
rect 5460 10150 5620 10230
rect 5220 9980 5620 10150
rect 5920 10230 6320 10380
rect 5920 10150 6080 10230
rect 6160 10150 6320 10230
rect 5920 9980 6320 10150
rect 6620 10230 7020 10380
rect 6620 10150 6780 10230
rect 6860 10150 7020 10230
rect 6620 9980 7020 10150
rect 7320 10230 7720 10380
rect 7320 10150 7480 10230
rect 7560 10150 7720 10230
rect 7320 9980 7720 10150
rect 8020 10230 8420 10380
rect 8020 10150 8180 10230
rect 8260 10150 8420 10230
rect 8020 9980 8420 10150
rect 8720 10230 9120 10380
rect 8720 10150 8880 10230
rect 8960 10150 9120 10230
rect 8720 9980 9120 10150
rect 9420 10230 9820 10380
rect 9420 10150 9580 10230
rect 9660 10150 9820 10230
rect 9420 9980 9820 10150
rect 10120 10230 10520 10380
rect 10120 10150 10280 10230
rect 10360 10150 10520 10230
rect 10120 9980 10520 10150
rect 30320 10230 30720 10380
rect 30320 10150 30480 10230
rect 30560 10150 30720 10230
rect 30320 9980 30720 10150
rect 31020 10230 31420 10380
rect 31020 10150 31180 10230
rect 31260 10150 31420 10230
rect 31020 9980 31420 10150
rect 31720 10230 32120 10380
rect 31720 10150 31880 10230
rect 31960 10150 32120 10230
rect 31720 9980 32120 10150
rect 32420 10230 32820 10380
rect 32420 10150 32580 10230
rect 32660 10150 32820 10230
rect 32420 9980 32820 10150
rect 33120 10230 33520 10380
rect 33120 10150 33280 10230
rect 33360 10150 33520 10230
rect 33120 9980 33520 10150
rect 33820 10230 34220 10380
rect 33820 10150 33980 10230
rect 34060 10150 34220 10230
rect 33820 9980 34220 10150
rect 34520 10230 34920 10380
rect 34520 10150 34680 10230
rect 34760 10150 34920 10230
rect 34520 9980 34920 10150
rect 35220 10230 35620 10380
rect 35220 10150 35380 10230
rect 35460 10150 35620 10230
rect 35220 9980 35620 10150
rect 35920 10230 36320 10380
rect 35920 10150 36080 10230
rect 36160 10150 36320 10230
rect 35920 9980 36320 10150
rect 36620 10230 37020 10380
rect 36620 10150 36780 10230
rect 36860 10150 37020 10230
rect 36620 9980 37020 10150
rect 37320 10230 37720 10380
rect 37320 10150 37480 10230
rect 37560 10150 37720 10230
rect 37320 9980 37720 10150
rect 38020 10230 38420 10380
rect 38020 10150 38180 10230
rect 38260 10150 38420 10230
rect 38020 9980 38420 10150
rect 38720 10230 39120 10380
rect 38720 10150 38880 10230
rect 38960 10150 39120 10230
rect 38720 9980 39120 10150
rect 39420 10230 39820 10380
rect 39420 10150 39580 10230
rect 39660 10150 39820 10230
rect 39420 9980 39820 10150
rect 40120 10230 40520 10380
rect 40120 10150 40280 10230
rect 40360 10150 40520 10230
rect 40120 9980 40520 10150
rect 320 9530 720 9680
rect 320 9450 480 9530
rect 560 9450 720 9530
rect 320 9280 720 9450
rect 1020 9530 1420 9680
rect 1020 9450 1180 9530
rect 1260 9450 1420 9530
rect 1020 9280 1420 9450
rect 1720 9530 2120 9680
rect 1720 9450 1880 9530
rect 1960 9450 2120 9530
rect 1720 9280 2120 9450
rect 2420 9530 2820 9680
rect 2420 9450 2580 9530
rect 2660 9450 2820 9530
rect 2420 9280 2820 9450
rect 3120 9530 3520 9680
rect 3120 9450 3280 9530
rect 3360 9450 3520 9530
rect 3120 9280 3520 9450
rect 3820 9530 4220 9680
rect 3820 9450 3980 9530
rect 4060 9450 4220 9530
rect 3820 9280 4220 9450
rect 4520 9530 4920 9680
rect 4520 9450 4680 9530
rect 4760 9450 4920 9530
rect 4520 9280 4920 9450
rect 5220 9530 5620 9680
rect 5220 9450 5380 9530
rect 5460 9450 5620 9530
rect 5220 9280 5620 9450
rect 5920 9530 6320 9680
rect 5920 9450 6080 9530
rect 6160 9450 6320 9530
rect 5920 9280 6320 9450
rect 6620 9530 7020 9680
rect 6620 9450 6780 9530
rect 6860 9450 7020 9530
rect 6620 9280 7020 9450
rect 7320 9530 7720 9680
rect 7320 9450 7480 9530
rect 7560 9450 7720 9530
rect 7320 9280 7720 9450
rect 8020 9530 8420 9680
rect 8020 9450 8180 9530
rect 8260 9450 8420 9530
rect 8020 9280 8420 9450
rect 8720 9530 9120 9680
rect 8720 9450 8880 9530
rect 8960 9450 9120 9530
rect 8720 9280 9120 9450
rect 9420 9530 9820 9680
rect 9420 9450 9580 9530
rect 9660 9450 9820 9530
rect 9420 9280 9820 9450
rect 10120 9530 10520 9680
rect 10120 9450 10280 9530
rect 10360 9450 10520 9530
rect 10120 9280 10520 9450
rect 30320 9530 30720 9680
rect 30320 9450 30480 9530
rect 30560 9450 30720 9530
rect 30320 9280 30720 9450
rect 31020 9530 31420 9680
rect 31020 9450 31180 9530
rect 31260 9450 31420 9530
rect 31020 9280 31420 9450
rect 31720 9530 32120 9680
rect 31720 9450 31880 9530
rect 31960 9450 32120 9530
rect 31720 9280 32120 9450
rect 32420 9530 32820 9680
rect 32420 9450 32580 9530
rect 32660 9450 32820 9530
rect 32420 9280 32820 9450
rect 33120 9530 33520 9680
rect 33120 9450 33280 9530
rect 33360 9450 33520 9530
rect 33120 9280 33520 9450
rect 33820 9530 34220 9680
rect 33820 9450 33980 9530
rect 34060 9450 34220 9530
rect 33820 9280 34220 9450
rect 34520 9530 34920 9680
rect 34520 9450 34680 9530
rect 34760 9450 34920 9530
rect 34520 9280 34920 9450
rect 35220 9530 35620 9680
rect 35220 9450 35380 9530
rect 35460 9450 35620 9530
rect 35220 9280 35620 9450
rect 35920 9530 36320 9680
rect 35920 9450 36080 9530
rect 36160 9450 36320 9530
rect 35920 9280 36320 9450
rect 36620 9530 37020 9680
rect 36620 9450 36780 9530
rect 36860 9450 37020 9530
rect 36620 9280 37020 9450
rect 37320 9530 37720 9680
rect 37320 9450 37480 9530
rect 37560 9450 37720 9530
rect 37320 9280 37720 9450
rect 38020 9530 38420 9680
rect 38020 9450 38180 9530
rect 38260 9450 38420 9530
rect 38020 9280 38420 9450
rect 38720 9530 39120 9680
rect 38720 9450 38880 9530
rect 38960 9450 39120 9530
rect 38720 9280 39120 9450
rect 39420 9530 39820 9680
rect 39420 9450 39580 9530
rect 39660 9450 39820 9530
rect 39420 9280 39820 9450
rect 40120 9530 40520 9680
rect 40120 9450 40280 9530
rect 40360 9450 40520 9530
rect 40120 9280 40520 9450
rect 320 8830 720 8980
rect 320 8750 480 8830
rect 560 8750 720 8830
rect 320 8580 720 8750
rect 1020 8830 1420 8980
rect 1020 8750 1180 8830
rect 1260 8750 1420 8830
rect 1020 8580 1420 8750
rect 1720 8830 2120 8980
rect 1720 8750 1880 8830
rect 1960 8750 2120 8830
rect 1720 8580 2120 8750
rect 2420 8830 2820 8980
rect 2420 8750 2580 8830
rect 2660 8750 2820 8830
rect 2420 8580 2820 8750
rect 3120 8830 3520 8980
rect 3120 8750 3280 8830
rect 3360 8750 3520 8830
rect 3120 8580 3520 8750
rect 3820 8830 4220 8980
rect 3820 8750 3980 8830
rect 4060 8750 4220 8830
rect 3820 8580 4220 8750
rect 4520 8830 4920 8980
rect 4520 8750 4680 8830
rect 4760 8750 4920 8830
rect 4520 8580 4920 8750
rect 5220 8830 5620 8980
rect 5220 8750 5380 8830
rect 5460 8750 5620 8830
rect 5220 8580 5620 8750
rect 5920 8830 6320 8980
rect 5920 8750 6080 8830
rect 6160 8750 6320 8830
rect 5920 8580 6320 8750
rect 6620 8830 7020 8980
rect 6620 8750 6780 8830
rect 6860 8750 7020 8830
rect 6620 8580 7020 8750
rect 7320 8830 7720 8980
rect 7320 8750 7480 8830
rect 7560 8750 7720 8830
rect 7320 8580 7720 8750
rect 8020 8830 8420 8980
rect 8020 8750 8180 8830
rect 8260 8750 8420 8830
rect 8020 8580 8420 8750
rect 8720 8830 9120 8980
rect 8720 8750 8880 8830
rect 8960 8750 9120 8830
rect 8720 8580 9120 8750
rect 9420 8830 9820 8980
rect 9420 8750 9580 8830
rect 9660 8750 9820 8830
rect 9420 8580 9820 8750
rect 10120 8830 10520 8980
rect 10120 8750 10280 8830
rect 10360 8750 10520 8830
rect 10120 8580 10520 8750
rect 30320 8830 30720 8980
rect 30320 8750 30480 8830
rect 30560 8750 30720 8830
rect 30320 8580 30720 8750
rect 31020 8830 31420 8980
rect 31020 8750 31180 8830
rect 31260 8750 31420 8830
rect 31020 8580 31420 8750
rect 31720 8830 32120 8980
rect 31720 8750 31880 8830
rect 31960 8750 32120 8830
rect 31720 8580 32120 8750
rect 32420 8830 32820 8980
rect 32420 8750 32580 8830
rect 32660 8750 32820 8830
rect 32420 8580 32820 8750
rect 33120 8830 33520 8980
rect 33120 8750 33280 8830
rect 33360 8750 33520 8830
rect 33120 8580 33520 8750
rect 33820 8830 34220 8980
rect 33820 8750 33980 8830
rect 34060 8750 34220 8830
rect 33820 8580 34220 8750
rect 34520 8830 34920 8980
rect 34520 8750 34680 8830
rect 34760 8750 34920 8830
rect 34520 8580 34920 8750
rect 35220 8830 35620 8980
rect 35220 8750 35380 8830
rect 35460 8750 35620 8830
rect 35220 8580 35620 8750
rect 35920 8830 36320 8980
rect 35920 8750 36080 8830
rect 36160 8750 36320 8830
rect 35920 8580 36320 8750
rect 36620 8830 37020 8980
rect 36620 8750 36780 8830
rect 36860 8750 37020 8830
rect 36620 8580 37020 8750
rect 37320 8830 37720 8980
rect 37320 8750 37480 8830
rect 37560 8750 37720 8830
rect 37320 8580 37720 8750
rect 38020 8830 38420 8980
rect 38020 8750 38180 8830
rect 38260 8750 38420 8830
rect 38020 8580 38420 8750
rect 38720 8830 39120 8980
rect 38720 8750 38880 8830
rect 38960 8750 39120 8830
rect 38720 8580 39120 8750
rect 39420 8830 39820 8980
rect 39420 8750 39580 8830
rect 39660 8750 39820 8830
rect 39420 8580 39820 8750
rect 40120 8830 40520 8980
rect 40120 8750 40280 8830
rect 40360 8750 40520 8830
rect 40120 8580 40520 8750
rect 320 8130 720 8280
rect 320 8050 480 8130
rect 560 8050 720 8130
rect 320 7880 720 8050
rect 1020 8130 1420 8280
rect 1020 8050 1180 8130
rect 1260 8050 1420 8130
rect 1020 7880 1420 8050
rect 1720 8130 2120 8280
rect 1720 8050 1880 8130
rect 1960 8050 2120 8130
rect 1720 7880 2120 8050
rect 2420 8130 2820 8280
rect 2420 8050 2580 8130
rect 2660 8050 2820 8130
rect 2420 7880 2820 8050
rect 3120 8130 3520 8280
rect 3120 8050 3280 8130
rect 3360 8050 3520 8130
rect 3120 7880 3520 8050
rect 3820 8130 4220 8280
rect 3820 8050 3980 8130
rect 4060 8050 4220 8130
rect 3820 7880 4220 8050
rect 4520 8130 4920 8280
rect 4520 8050 4680 8130
rect 4760 8050 4920 8130
rect 4520 7880 4920 8050
rect 5220 8130 5620 8280
rect 5220 8050 5380 8130
rect 5460 8050 5620 8130
rect 5220 7880 5620 8050
rect 5920 8130 6320 8280
rect 5920 8050 6080 8130
rect 6160 8050 6320 8130
rect 5920 7880 6320 8050
rect 6620 8130 7020 8280
rect 6620 8050 6780 8130
rect 6860 8050 7020 8130
rect 6620 7880 7020 8050
rect 7320 8130 7720 8280
rect 7320 8050 7480 8130
rect 7560 8050 7720 8130
rect 7320 7880 7720 8050
rect 8020 8130 8420 8280
rect 8020 8050 8180 8130
rect 8260 8050 8420 8130
rect 8020 7880 8420 8050
rect 8720 8130 9120 8280
rect 8720 8050 8880 8130
rect 8960 8050 9120 8130
rect 8720 7880 9120 8050
rect 9420 8130 9820 8280
rect 9420 8050 9580 8130
rect 9660 8050 9820 8130
rect 9420 7880 9820 8050
rect 10120 8130 10520 8280
rect 10120 8050 10280 8130
rect 10360 8050 10520 8130
rect 10120 7880 10520 8050
rect 30320 8130 30720 8280
rect 30320 8050 30480 8130
rect 30560 8050 30720 8130
rect 30320 7880 30720 8050
rect 31020 8130 31420 8280
rect 31020 8050 31180 8130
rect 31260 8050 31420 8130
rect 31020 7880 31420 8050
rect 31720 8130 32120 8280
rect 31720 8050 31880 8130
rect 31960 8050 32120 8130
rect 31720 7880 32120 8050
rect 32420 8130 32820 8280
rect 32420 8050 32580 8130
rect 32660 8050 32820 8130
rect 32420 7880 32820 8050
rect 33120 8130 33520 8280
rect 33120 8050 33280 8130
rect 33360 8050 33520 8130
rect 33120 7880 33520 8050
rect 33820 8130 34220 8280
rect 33820 8050 33980 8130
rect 34060 8050 34220 8130
rect 33820 7880 34220 8050
rect 34520 8130 34920 8280
rect 34520 8050 34680 8130
rect 34760 8050 34920 8130
rect 34520 7880 34920 8050
rect 35220 8130 35620 8280
rect 35220 8050 35380 8130
rect 35460 8050 35620 8130
rect 35220 7880 35620 8050
rect 35920 8130 36320 8280
rect 35920 8050 36080 8130
rect 36160 8050 36320 8130
rect 35920 7880 36320 8050
rect 36620 8130 37020 8280
rect 36620 8050 36780 8130
rect 36860 8050 37020 8130
rect 36620 7880 37020 8050
rect 37320 8130 37720 8280
rect 37320 8050 37480 8130
rect 37560 8050 37720 8130
rect 37320 7880 37720 8050
rect 38020 8130 38420 8280
rect 38020 8050 38180 8130
rect 38260 8050 38420 8130
rect 38020 7880 38420 8050
rect 38720 8130 39120 8280
rect 38720 8050 38880 8130
rect 38960 8050 39120 8130
rect 38720 7880 39120 8050
rect 39420 8130 39820 8280
rect 39420 8050 39580 8130
rect 39660 8050 39820 8130
rect 39420 7880 39820 8050
rect 40120 8130 40520 8280
rect 40120 8050 40280 8130
rect 40360 8050 40520 8130
rect 40120 7880 40520 8050
<< mimcapcontact >>
rect 480 10150 560 10230
rect 1180 10150 1260 10230
rect 1880 10150 1960 10230
rect 2580 10150 2660 10230
rect 3280 10150 3360 10230
rect 3980 10150 4060 10230
rect 4680 10150 4760 10230
rect 5380 10150 5460 10230
rect 6080 10150 6160 10230
rect 6780 10150 6860 10230
rect 7480 10150 7560 10230
rect 8180 10150 8260 10230
rect 8880 10150 8960 10230
rect 9580 10150 9660 10230
rect 10280 10150 10360 10230
rect 30480 10150 30560 10230
rect 31180 10150 31260 10230
rect 31880 10150 31960 10230
rect 32580 10150 32660 10230
rect 33280 10150 33360 10230
rect 33980 10150 34060 10230
rect 34680 10150 34760 10230
rect 35380 10150 35460 10230
rect 36080 10150 36160 10230
rect 36780 10150 36860 10230
rect 37480 10150 37560 10230
rect 38180 10150 38260 10230
rect 38880 10150 38960 10230
rect 39580 10150 39660 10230
rect 40280 10150 40360 10230
rect 480 9450 560 9530
rect 1180 9450 1260 9530
rect 1880 9450 1960 9530
rect 2580 9450 2660 9530
rect 3280 9450 3360 9530
rect 3980 9450 4060 9530
rect 4680 9450 4760 9530
rect 5380 9450 5460 9530
rect 6080 9450 6160 9530
rect 6780 9450 6860 9530
rect 7480 9450 7560 9530
rect 8180 9450 8260 9530
rect 8880 9450 8960 9530
rect 9580 9450 9660 9530
rect 10280 9450 10360 9530
rect 30480 9450 30560 9530
rect 31180 9450 31260 9530
rect 31880 9450 31960 9530
rect 32580 9450 32660 9530
rect 33280 9450 33360 9530
rect 33980 9450 34060 9530
rect 34680 9450 34760 9530
rect 35380 9450 35460 9530
rect 36080 9450 36160 9530
rect 36780 9450 36860 9530
rect 37480 9450 37560 9530
rect 38180 9450 38260 9530
rect 38880 9450 38960 9530
rect 39580 9450 39660 9530
rect 40280 9450 40360 9530
rect 480 8750 560 8830
rect 1180 8750 1260 8830
rect 1880 8750 1960 8830
rect 2580 8750 2660 8830
rect 3280 8750 3360 8830
rect 3980 8750 4060 8830
rect 4680 8750 4760 8830
rect 5380 8750 5460 8830
rect 6080 8750 6160 8830
rect 6780 8750 6860 8830
rect 7480 8750 7560 8830
rect 8180 8750 8260 8830
rect 8880 8750 8960 8830
rect 9580 8750 9660 8830
rect 10280 8750 10360 8830
rect 30480 8750 30560 8830
rect 31180 8750 31260 8830
rect 31880 8750 31960 8830
rect 32580 8750 32660 8830
rect 33280 8750 33360 8830
rect 33980 8750 34060 8830
rect 34680 8750 34760 8830
rect 35380 8750 35460 8830
rect 36080 8750 36160 8830
rect 36780 8750 36860 8830
rect 37480 8750 37560 8830
rect 38180 8750 38260 8830
rect 38880 8750 38960 8830
rect 39580 8750 39660 8830
rect 40280 8750 40360 8830
rect 480 8050 560 8130
rect 1180 8050 1260 8130
rect 1880 8050 1960 8130
rect 2580 8050 2660 8130
rect 3280 8050 3360 8130
rect 3980 8050 4060 8130
rect 4680 8050 4760 8130
rect 5380 8050 5460 8130
rect 6080 8050 6160 8130
rect 6780 8050 6860 8130
rect 7480 8050 7560 8130
rect 8180 8050 8260 8130
rect 8880 8050 8960 8130
rect 9580 8050 9660 8130
rect 10280 8050 10360 8130
rect 30480 8050 30560 8130
rect 31180 8050 31260 8130
rect 31880 8050 31960 8130
rect 32580 8050 32660 8130
rect 33280 8050 33360 8130
rect 33980 8050 34060 8130
rect 34680 8050 34760 8130
rect 35380 8050 35460 8130
rect 36080 8050 36160 8130
rect 36780 8050 36860 8130
rect 37480 8050 37560 8130
rect 38180 8050 38260 8130
rect 38880 8050 38960 8130
rect 39580 8050 39660 8130
rect 40280 8050 40360 8130
<< metal4 >>
rect -400 10690 11590 10700
rect -400 10610 -390 10690
rect -310 10610 11500 10690
rect 11580 10610 11590 10690
rect -400 10600 11590 10610
rect 29600 10690 41590 10700
rect 29600 10610 29610 10690
rect 29690 10610 41500 10690
rect 41580 10610 41590 10690
rect 29600 10600 41590 10610
rect -230 10520 11420 10530
rect -230 10440 -220 10520
rect -140 10440 11330 10520
rect 11410 10440 11420 10520
rect -230 10430 11420 10440
rect 29770 10520 41420 10530
rect 29770 10440 29780 10520
rect 29860 10440 41330 10520
rect 41410 10440 41420 10520
rect 29770 10430 41420 10440
rect 470 10230 3370 10240
rect 470 10150 480 10230
rect 560 10150 1180 10230
rect 1260 10150 1880 10230
rect 1960 10150 2580 10230
rect 2660 10150 3280 10230
rect 3360 10150 3370 10230
rect 470 10140 3370 10150
rect 3970 10230 6870 10240
rect 3970 10150 3980 10230
rect 4060 10150 4680 10230
rect 4760 10150 5380 10230
rect 5460 10150 6080 10230
rect 6160 10150 6780 10230
rect 6860 10150 6870 10230
rect 3970 10140 6870 10150
rect 7470 10230 10370 10240
rect 7470 10150 7480 10230
rect 7560 10150 8180 10230
rect 8260 10150 8880 10230
rect 8960 10150 9580 10230
rect 9660 10150 10280 10230
rect 10360 10150 10370 10230
rect 7470 10140 10370 10150
rect 30470 10230 33370 10240
rect 30470 10150 30480 10230
rect 30560 10150 31180 10230
rect 31260 10150 31880 10230
rect 31960 10150 32580 10230
rect 32660 10150 33280 10230
rect 33360 10150 33370 10230
rect 30470 10140 33370 10150
rect 33970 10230 36870 10240
rect 33970 10150 33980 10230
rect 34060 10150 34680 10230
rect 34760 10150 35380 10230
rect 35460 10150 36080 10230
rect 36160 10150 36780 10230
rect 36860 10150 36870 10230
rect 33970 10140 36870 10150
rect 37470 10230 40370 10240
rect 37470 10150 37480 10230
rect 37560 10150 38180 10230
rect 38260 10150 38880 10230
rect 38960 10150 39580 10230
rect 39660 10150 40280 10230
rect 40360 10150 40370 10230
rect 37470 10140 40370 10150
rect 1870 9540 1970 10140
rect 5370 9540 5470 10140
rect 8870 9540 8970 10140
rect 31870 9540 31970 10140
rect 35370 9540 35470 10140
rect 38870 9540 38970 10140
rect 470 9530 3370 9540
rect 470 9450 480 9530
rect 560 9450 1180 9530
rect 1260 9450 1880 9530
rect 1960 9450 2580 9530
rect 2660 9450 3280 9530
rect 3360 9450 3370 9530
rect 470 9440 3370 9450
rect 3970 9530 6870 9540
rect 3970 9450 3980 9530
rect 4060 9450 4680 9530
rect 4760 9450 5380 9530
rect 5460 9450 6080 9530
rect 6160 9450 6780 9530
rect 6860 9450 6870 9530
rect 3970 9440 6870 9450
rect 7470 9530 10370 9540
rect 7470 9450 7480 9530
rect 7560 9450 8180 9530
rect 8260 9450 8880 9530
rect 8960 9450 9580 9530
rect 9660 9450 10280 9530
rect 10360 9450 10370 9530
rect 7470 9440 10370 9450
rect 30470 9530 33370 9540
rect 30470 9450 30480 9530
rect 30560 9450 31180 9530
rect 31260 9450 31880 9530
rect 31960 9450 32580 9530
rect 32660 9450 33280 9530
rect 33360 9450 33370 9530
rect 30470 9440 33370 9450
rect 33970 9530 36870 9540
rect 33970 9450 33980 9530
rect 34060 9450 34680 9530
rect 34760 9450 35380 9530
rect 35460 9450 36080 9530
rect 36160 9450 36780 9530
rect 36860 9450 36870 9530
rect 33970 9440 36870 9450
rect 37470 9530 40370 9540
rect 37470 9450 37480 9530
rect 37560 9450 38180 9530
rect 38260 9450 38880 9530
rect 38960 9450 39580 9530
rect 39660 9450 40280 9530
rect 40360 9450 40370 9530
rect 37470 9440 40370 9450
rect 1870 8840 1970 9440
rect 5370 8840 5470 9440
rect 8870 8840 8970 9440
rect 31870 8840 31970 9440
rect 35370 8840 35470 9440
rect 38870 8840 38970 9440
rect 470 8830 3370 8840
rect 470 8750 480 8830
rect 560 8750 1180 8830
rect 1260 8750 1880 8830
rect 1960 8750 2580 8830
rect 2660 8750 3280 8830
rect 3360 8750 3370 8830
rect 470 8740 3370 8750
rect 3970 8830 6870 8840
rect 3970 8750 3980 8830
rect 4060 8750 4680 8830
rect 4760 8750 5380 8830
rect 5460 8750 6080 8830
rect 6160 8750 6780 8830
rect 6860 8750 6870 8830
rect 3970 8740 6870 8750
rect 7470 8830 10370 8840
rect 7470 8750 7480 8830
rect 7560 8750 8180 8830
rect 8260 8750 8880 8830
rect 8960 8750 9580 8830
rect 9660 8750 10280 8830
rect 10360 8750 10370 8830
rect 7470 8740 10370 8750
rect 30470 8830 33370 8840
rect 30470 8750 30480 8830
rect 30560 8750 31180 8830
rect 31260 8750 31880 8830
rect 31960 8750 32580 8830
rect 32660 8750 33280 8830
rect 33360 8750 33370 8830
rect 30470 8740 33370 8750
rect 33970 8830 36870 8840
rect 33970 8750 33980 8830
rect 34060 8750 34680 8830
rect 34760 8750 35380 8830
rect 35460 8750 36080 8830
rect 36160 8750 36780 8830
rect 36860 8750 36870 8830
rect 33970 8740 36870 8750
rect 37470 8830 40370 8840
rect 37470 8750 37480 8830
rect 37560 8750 38180 8830
rect 38260 8750 38880 8830
rect 38960 8750 39580 8830
rect 39660 8750 40280 8830
rect 40360 8750 40370 8830
rect 37470 8740 40370 8750
rect 1870 8140 1970 8740
rect 5370 8140 5470 8740
rect 8870 8140 8970 8740
rect 31870 8140 31970 8740
rect 35370 8140 35470 8740
rect 38870 8140 38970 8740
rect 470 8130 3370 8140
rect 470 8050 480 8130
rect 560 8050 1180 8130
rect 1260 8050 1880 8130
rect 1960 8050 2580 8130
rect 2660 8050 3280 8130
rect 3360 8050 3370 8130
rect 470 8040 3370 8050
rect 3970 8130 6870 8140
rect 3970 8050 3980 8130
rect 4060 8050 4680 8130
rect 4760 8050 5380 8130
rect 5460 8050 6080 8130
rect 6160 8050 6780 8130
rect 6860 8050 6870 8130
rect 3970 8040 6870 8050
rect 7470 8130 10370 8140
rect 7470 8050 7480 8130
rect 7560 8050 8180 8130
rect 8260 8050 8880 8130
rect 8960 8050 9580 8130
rect 9660 8050 10280 8130
rect 10360 8050 10370 8130
rect 7470 8040 10370 8050
rect 30470 8130 33370 8140
rect 30470 8050 30480 8130
rect 30560 8050 31180 8130
rect 31260 8050 31880 8130
rect 31960 8050 32580 8130
rect 32660 8050 33280 8130
rect 33360 8050 33370 8130
rect 30470 8040 33370 8050
rect 33970 8130 36870 8140
rect 33970 8050 33980 8130
rect 34060 8050 34680 8130
rect 34760 8050 35380 8130
rect 35460 8050 36080 8130
rect 36160 8050 36780 8130
rect 36860 8050 36870 8130
rect 33970 8040 36870 8050
rect 37470 8130 40370 8140
rect 37470 8050 37480 8130
rect 37560 8050 38180 8130
rect 38260 8050 38880 8130
rect 38960 8050 39580 8130
rect 39660 8050 40280 8130
rect 40360 8050 40370 8130
rect 37470 8040 40370 8050
rect 3270 7600 3370 8040
rect 3270 7520 3280 7600
rect 3360 7520 3370 7600
rect 3270 7510 3370 7520
rect 6770 7490 6870 8040
rect 10270 7600 10370 8040
rect 10270 7520 10280 7600
rect 10360 7520 10370 7600
rect 10270 7510 10370 7520
rect 33270 7600 33370 8040
rect 33270 7520 33280 7600
rect 33360 7520 33370 7600
rect 33270 7510 33370 7520
rect 6770 7410 6780 7490
rect 6860 7410 6870 7490
rect 6770 7400 6870 7410
rect 36770 7490 36870 8040
rect 40270 7600 40370 8040
rect 40270 7520 40280 7600
rect 40360 7520 40370 7600
rect 40270 7510 40370 7520
rect 36770 7410 36780 7490
rect 36860 7410 36870 7490
rect 36770 7400 36870 7410
rect -230 1320 11420 1330
rect -230 1240 -220 1320
rect -140 1240 11330 1320
rect 11410 1240 11420 1320
rect -230 1230 11420 1240
rect -400 1160 11590 1170
rect -400 1080 -390 1160
rect -310 1080 11500 1160
rect 11580 1080 11590 1160
rect -400 1070 11590 1080
rect 29770 -8680 41420 -8670
rect 29770 -8760 29780 -8680
rect 29860 -8760 41330 -8680
rect 41410 -8760 41420 -8680
rect 29770 -8770 41420 -8760
rect 29600 -8840 41590 -8830
rect 29600 -8920 29610 -8840
rect 29690 -8920 41500 -8840
rect 41580 -8920 41590 -8840
rect 29600 -8930 41590 -8920
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 2950 0 1 2720
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1723858470
transform 1 0 2950 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11
timestamp 1723858470
transform 1 0 2950 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12
timestamp 1723858470
transform 1 0 230 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13
timestamp 1723858470
transform 1 0 230 0 1 2720
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14
timestamp 1723858470
transform 1 0 230 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15
timestamp 1723858470
transform 1 0 1590 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16
timestamp 1723858470
transform 1 0 1590 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17
timestamp 1723858470
transform 1 0 1590 0 1 2720
box 0 0 1340 1340
<< labels >>
flabel metal2 910 7580 910 7580 1 FreeSans 800 0 0 80 cap_res1
flabel metal3 5460 7450 5460 7450 3 FreeSans 800 0 80 0 cap_res2
flabel metal1 3970 4740 3970 4740 3 FreeSans 800 0 80 0 Vbe2
flabel poly 9420 5380 9420 5380 5 FreeSans 800 0 0 -80 V_TOP
flabel metal1 10120 2480 10120 2480 3 FreeSans 800 0 400 0 START_UP_NFET1
flabel metal2 10420 3750 10420 3750 1 FreeSans 800 0 0 160 V_CUR_REF_REG
flabel metal2 10520 4340 10520 4340 5 FreeSans 800 0 0 -80 V_mir2
flabel metal1 5170 1990 5170 1990 3 FreeSans 800 0 80 0 NFET_GATE_10uA
flabel metal2 12200 6200 12200 6200 3 FreeSans 800 0 400 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 12200 7240 12200 7240 3 FreeSans 800 0 400 0 V_CMFB_S1
port 10 e
flabel metal2 12200 4060 12200 4060 3 FreeSans 800 0 400 0 ERR_AMP_REF
port 3 e
flabel metal3 11580 9500 11580 9500 3 FreeSans 800 0 400 0 VDDA
port 4 e
flabel metal3 11410 9050 11410 9050 3 FreeSans 800 0 400 0 GNDA
port 2 e
flabel metal2 5900 3750 5900 3750 1 FreeSans 800 0 0 160 Vin+
flabel metal2 5890 4040 5890 4040 5 FreeSans 800 0 0 -160 Vin-
flabel metal1 4610 2910 4610 2910 3 FreeSans 800 0 400 0 START_UP
flabel metal2 8620 4260 8620 4260 7 FreeSans 480 0 -240 0 1st_Vout_2
flabel metal2 8900 3570 8900 3570 7 FreeSans 800 0 -400 0 V_p_2
flabel metal2 7420 3570 7420 3570 3 FreeSans 800 0 400 0 V_p_1
flabel metal2 5800 4340 5800 4340 5 FreeSans 800 0 0 -80 V_mir1
flabel metal2 7700 4260 7700 4260 3 FreeSans 480 0 240 0 1st_Vout_1
flabel metal2 12200 5560 12200 5560 3 FreeSans 800 0 400 0 VB1_CUR_BIAS
port 1 e
flabel metal2 12200 6690 12200 6690 3 FreeSans 800 0 400 0 V_CMFB_S3
port 12 e
flabel via1 8160 7170 8160 7170 1 FreeSans 800 0 0 400 PFET_GATE_10uA
flabel metal1 9610 1100 9610 1100 5 FreeSans 800 0 0 -400 V_CMFB_S4
port 11 s
flabel metal1 8400 1170 8400 1170 3 FreeSans 800 0 400 0 VB3_CUR_BIAS
port 6 e
flabel metal1 7920 1170 7920 1170 7 FreeSans 800 0 -400 0 ERR_AMP_CUR_BIAS
port 7 w
flabel metal1 6710 1100 6710 1100 5 FreeSans 800 0 0 -400 VB2_CUR_BIAS
port 5 s
flabel metal1 9390 1100 9390 1100 5 FreeSans 800 0 0 -400 V_CMFB_S2
port 8 s
flabel metal2 30910 7580 30910 7580 1 FreeSans 800 0 0 80 cap_res1
flabel metal3 35460 7450 35460 7450 3 FreeSans 800 0 80 0 cap_res2
flabel metal3 41580 9500 41580 9500 3 FreeSans 800 0 400 0 VDDA
port 4 e
flabel metal3 41410 9050 41410 9050 3 FreeSans 800 0 400 0 GNDA
port 2 e
flabel space 39610 -8900 39610 -8900 5 FreeSans 800 0 0 -400 V_CMFB_S4
port 11 s
flabel space 38400 -8830 38400 -8830 3 FreeSans 800 0 400 0 VB3_CUR_BIAS
port 6 e
flabel space 37920 -8830 37920 -8830 7 FreeSans 800 0 -400 0 ERR_AMP_CUR_BIAS
port 7 w
flabel space 36710 -8900 36710 -8900 5 FreeSans 800 0 0 -400 VB2_CUR_BIAS
port 5 s
flabel space 39390 -8900 39390 -8900 5 FreeSans 800 0 0 -400 V_CMFB_S2
port 8 s
flabel via1 38160 4170 38160 4170 1 FreeSans 800 0 0 400 PFET_GATE_10uA
flabel metal2 42200 3690 42200 3690 3 FreeSans 800 0 400 0 V_CMFB_S3
port 12 e
flabel metal2 42200 2560 42200 2560 3 FreeSans 800 0 400 0 VB1_CUR_BIAS
port 1 e
flabel metal2 37700 1260 37700 1260 3 FreeSans 480 0 240 0 1st_Vout_1
flabel metal2 35800 1340 35800 1340 5 FreeSans 800 0 0 -80 V_mir1
flabel metal2 37420 570 37420 570 3 FreeSans 800 0 400 0 V_p_1
flabel metal2 38900 570 38900 570 7 FreeSans 800 0 -400 0 V_p_2
flabel metal2 38620 1260 38620 1260 7 FreeSans 480 0 -240 0 1st_Vout_2
flabel metal2 35890 1040 35890 1040 5 FreeSans 800 0 0 -160 Vin-
flabel metal2 35900 750 35900 750 1 FreeSans 800 0 0 160 Vin+
flabel metal2 42200 1060 42200 1060 3 FreeSans 800 0 400 0 ERR_AMP_REF
port 3 e
flabel metal2 42200 4240 42200 4240 3 FreeSans 800 0 400 0 V_CMFB_S1
port 10 e
flabel metal2 42200 3200 42200 3200 3 FreeSans 800 0 400 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 40520 1340 40520 1340 5 FreeSans 800 0 0 -80 V_mir2
flabel metal2 40420 750 40420 750 1 FreeSans 800 0 0 160 V_CUR_REF_REG
flabel metal1 40120 -520 40120 -520 3 FreeSans 800 0 400 0 START_UP_NFET1
flabel poly 39420 2380 39420 2380 5 FreeSans 800 0 0 -80 V_TOP
flabel locali s 35148 -4970 35188 -4852 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 34989 -4947 35038 -4846 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 35560 -5006 35664 -4758 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 36508 -4970 36548 -4852 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 36349 -4947 36398 -4846 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 36920 -5006 37024 -4758 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 33788 -4970 33828 -4852 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 33629 -4947 33678 -4846 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 34200 -5006 34304 -4758 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 36508 -7690 36548 -7572 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 36349 -7667 36398 -7566 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 36920 -7726 37024 -7478 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 35148 -7690 35188 -7572 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 34989 -7667 35038 -7566 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 35560 -7726 35664 -7478 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 33788 -7690 33828 -7572 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 33629 -7667 33678 -7566 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 34200 -7726 34304 -7478 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 36508 -6330 36548 -6212 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 36349 -6307 36398 -6206 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 36920 -6366 37024 -6118 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 33788 -6330 33828 -6212 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 33629 -6307 33678 -6206 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 34200 -6366 34304 -6118 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel locali s 35148 -6330 35188 -6212 0 FreeSans 400 270 0 0 Base
port 4 nsew
flabel locali s 34989 -6307 35038 -6206 0 FreeSans 400 270 0 0 Collector
port 3 nsew
flabel locali s 35560 -6366 35664 -6118 0 FreeSans 400 270 0 0 Emitter
port 2 nsew
flabel metal1 34270 -4540 34270 -4540 1 FreeSans 800 270 0 80 Vbe2
flabel metal1 35170 -1010 35170 -1010 3 FreeSans 800 0 80 0 NFET_GATE_10uA
flabel metal1 34610 -90 34610 -90 3 FreeSans 800 0 400 0 START_UP
<< end >>
