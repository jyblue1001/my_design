magic
tech sky130A
timestamp 1738185398
<< nwell >>
rect -2400 460 -2160 545
rect -3070 220 -1755 460
rect -1625 230 385 370
<< pwell >>
rect -2565 120 -2550 125
rect -3070 -90 -1755 115
rect -2100 -165 -2080 -90
<< nmos >>
rect -3000 10 -2985 110
rect -2855 10 -2840 110
rect -2710 10 -2695 110
rect -2565 10 -2550 110
rect -2420 10 -2405 110
rect -2275 10 -2260 110
rect -2130 10 -2115 110
rect -1985 10 -1970 110
rect -1840 10 -1825 110
rect -1505 0 -1445 100
rect -1395 0 -1335 100
rect -1285 0 -1225 100
rect -1175 0 -1115 100
rect -845 0 -785 100
rect -735 0 -675 100
rect -625 0 -565 100
rect -515 0 -455 100
rect -75 0 -15 100
rect 35 0 95 100
rect 145 0 205 100
rect 255 0 315 100
<< pmos >>
rect -3000 240 -2985 440
rect -2855 240 -2840 440
rect -2710 240 -2695 440
rect -2565 240 -2550 440
rect -2420 240 -2405 440
rect -2275 240 -2260 440
rect -2130 240 -2115 440
rect -1985 240 -1970 440
rect -1840 240 -1825 440
rect -1555 250 -1495 350
rect -1445 250 -1385 350
rect -1335 250 -1275 350
rect -1225 250 -1165 350
rect -1115 250 -1055 350
rect -1005 250 -945 350
rect -895 250 -835 350
rect -785 250 -725 350
rect -515 250 -455 350
rect -405 250 -345 350
rect -295 250 -235 350
rect -185 250 -125 350
rect -75 250 -15 350
rect 35 250 95 350
rect 145 250 205 350
rect 255 250 315 350
<< ndiff >>
rect -3050 95 -3000 110
rect -3050 25 -3035 95
rect -3015 25 -3000 95
rect -3050 10 -3000 25
rect -2985 95 -2935 110
rect -2985 25 -2970 95
rect -2950 25 -2935 95
rect -2985 10 -2935 25
rect -2905 95 -2855 110
rect -2905 25 -2890 95
rect -2870 25 -2855 95
rect -2905 10 -2855 25
rect -2840 95 -2790 110
rect -2840 25 -2825 95
rect -2805 25 -2790 95
rect -2840 10 -2790 25
rect -2760 95 -2710 110
rect -2760 25 -2745 95
rect -2725 25 -2710 95
rect -2760 10 -2710 25
rect -2695 95 -2645 110
rect -2695 25 -2680 95
rect -2660 25 -2645 95
rect -2695 10 -2645 25
rect -2615 95 -2565 110
rect -2615 25 -2600 95
rect -2580 25 -2565 95
rect -2615 10 -2565 25
rect -2550 95 -2500 110
rect -2550 25 -2535 95
rect -2515 25 -2500 95
rect -2550 10 -2500 25
rect -2470 95 -2420 110
rect -2470 25 -2455 95
rect -2435 25 -2420 95
rect -2470 10 -2420 25
rect -2405 95 -2355 110
rect -2405 25 -2390 95
rect -2370 25 -2355 95
rect -2405 10 -2355 25
rect -2325 95 -2275 110
rect -2325 25 -2310 95
rect -2290 25 -2275 95
rect -2325 10 -2275 25
rect -2260 95 -2210 110
rect -2260 25 -2245 95
rect -2225 25 -2210 95
rect -2260 10 -2210 25
rect -2180 95 -2130 110
rect -2180 25 -2165 95
rect -2145 25 -2130 95
rect -2180 10 -2130 25
rect -2115 95 -2065 110
rect -2115 25 -2100 95
rect -2080 25 -2065 95
rect -2115 10 -2065 25
rect -2035 95 -1985 110
rect -2035 25 -2020 95
rect -2000 25 -1985 95
rect -2035 10 -1985 25
rect -1970 95 -1920 110
rect -1970 25 -1955 95
rect -1935 25 -1920 95
rect -1970 10 -1920 25
rect -1890 95 -1840 110
rect -1890 25 -1875 95
rect -1855 25 -1840 95
rect -1890 10 -1840 25
rect -1825 95 -1775 110
rect -1825 25 -1810 95
rect -1790 25 -1775 95
rect -1825 10 -1775 25
rect -1555 85 -1505 100
rect -1555 15 -1540 85
rect -1520 15 -1505 85
rect -1555 0 -1505 15
rect -1445 85 -1395 100
rect -1445 15 -1430 85
rect -1410 15 -1395 85
rect -1445 0 -1395 15
rect -1335 85 -1285 100
rect -1335 15 -1320 85
rect -1300 15 -1285 85
rect -1335 0 -1285 15
rect -1225 85 -1175 100
rect -1225 15 -1210 85
rect -1190 15 -1175 85
rect -1225 0 -1175 15
rect -1115 85 -1065 100
rect -1115 15 -1100 85
rect -1080 15 -1065 85
rect -1115 0 -1065 15
rect -895 85 -845 100
rect -895 15 -880 85
rect -860 15 -845 85
rect -895 0 -845 15
rect -785 85 -735 100
rect -785 15 -770 85
rect -750 15 -735 85
rect -785 0 -735 15
rect -675 85 -625 100
rect -675 15 -660 85
rect -640 15 -625 85
rect -675 0 -625 15
rect -565 85 -515 100
rect -565 15 -550 85
rect -530 15 -515 85
rect -565 0 -515 15
rect -455 85 -405 100
rect -455 15 -440 85
rect -420 15 -405 85
rect -455 0 -405 15
rect -125 85 -75 100
rect -125 15 -110 85
rect -90 15 -75 85
rect -125 0 -75 15
rect -15 85 35 100
rect -15 15 0 85
rect 20 15 35 85
rect -15 0 35 15
rect 95 85 145 100
rect 95 15 110 85
rect 130 15 145 85
rect 95 0 145 15
rect 205 85 255 100
rect 205 15 220 85
rect 240 15 255 85
rect 205 0 255 15
rect 315 85 365 100
rect 315 15 330 85
rect 350 15 365 85
rect 315 0 365 15
<< pdiff >>
rect -3050 425 -3000 440
rect -3050 255 -3035 425
rect -3015 255 -3000 425
rect -3050 240 -3000 255
rect -2985 425 -2935 440
rect -2985 255 -2970 425
rect -2950 255 -2935 425
rect -2985 240 -2935 255
rect -2905 425 -2855 440
rect -2905 255 -2890 425
rect -2870 255 -2855 425
rect -2905 240 -2855 255
rect -2840 425 -2790 440
rect -2840 255 -2825 425
rect -2805 255 -2790 425
rect -2840 240 -2790 255
rect -2760 425 -2710 440
rect -2760 255 -2745 425
rect -2725 255 -2710 425
rect -2760 240 -2710 255
rect -2695 425 -2645 440
rect -2695 255 -2680 425
rect -2660 255 -2645 425
rect -2695 240 -2645 255
rect -2615 425 -2565 440
rect -2615 255 -2600 425
rect -2580 255 -2565 425
rect -2615 240 -2565 255
rect -2550 425 -2500 440
rect -2550 255 -2535 425
rect -2515 255 -2500 425
rect -2550 240 -2500 255
rect -2470 425 -2420 440
rect -2470 255 -2455 425
rect -2435 255 -2420 425
rect -2470 240 -2420 255
rect -2405 425 -2355 440
rect -2405 255 -2390 425
rect -2370 255 -2355 425
rect -2405 240 -2355 255
rect -2325 425 -2275 440
rect -2325 255 -2310 425
rect -2290 255 -2275 425
rect -2325 240 -2275 255
rect -2260 425 -2210 440
rect -2260 255 -2245 425
rect -2225 255 -2210 425
rect -2260 240 -2210 255
rect -2180 425 -2130 440
rect -2180 255 -2165 425
rect -2145 255 -2130 425
rect -2180 240 -2130 255
rect -2115 425 -2065 440
rect -2115 255 -2100 425
rect -2080 255 -2065 425
rect -2115 240 -2065 255
rect -2035 425 -1985 440
rect -2035 255 -2020 425
rect -2000 255 -1985 425
rect -2035 240 -1985 255
rect -1970 425 -1920 440
rect -1970 255 -1955 425
rect -1935 255 -1920 425
rect -1970 240 -1920 255
rect -1890 425 -1840 440
rect -1890 255 -1875 425
rect -1855 255 -1840 425
rect -1890 240 -1840 255
rect -1825 425 -1775 440
rect -1825 255 -1810 425
rect -1790 255 -1775 425
rect -1825 240 -1775 255
rect -1605 335 -1555 350
rect -1605 265 -1590 335
rect -1570 265 -1555 335
rect -1605 250 -1555 265
rect -1495 335 -1445 350
rect -1495 265 -1480 335
rect -1460 265 -1445 335
rect -1495 250 -1445 265
rect -1385 335 -1335 350
rect -1385 265 -1370 335
rect -1350 265 -1335 335
rect -1385 250 -1335 265
rect -1275 335 -1225 350
rect -1275 265 -1260 335
rect -1240 265 -1225 335
rect -1275 250 -1225 265
rect -1165 335 -1115 350
rect -1165 265 -1150 335
rect -1130 265 -1115 335
rect -1165 250 -1115 265
rect -1055 335 -1005 350
rect -1055 265 -1040 335
rect -1020 265 -1005 335
rect -1055 250 -1005 265
rect -945 335 -895 350
rect -945 265 -930 335
rect -910 265 -895 335
rect -945 250 -895 265
rect -835 335 -785 350
rect -835 265 -820 335
rect -800 265 -785 335
rect -835 250 -785 265
rect -725 335 -675 350
rect -725 265 -710 335
rect -690 265 -675 335
rect -725 250 -675 265
rect -565 335 -515 350
rect -565 265 -550 335
rect -530 265 -515 335
rect -565 250 -515 265
rect -455 335 -405 350
rect -455 265 -440 335
rect -420 265 -405 335
rect -455 250 -405 265
rect -345 335 -295 350
rect -345 265 -330 335
rect -310 265 -295 335
rect -345 250 -295 265
rect -235 335 -185 350
rect -235 265 -220 335
rect -200 265 -185 335
rect -235 250 -185 265
rect -125 335 -75 350
rect -125 265 -110 335
rect -90 265 -75 335
rect -125 250 -75 265
rect -15 335 35 350
rect -15 265 0 335
rect 20 265 35 335
rect -15 250 35 265
rect 95 335 145 350
rect 95 265 110 335
rect 130 265 145 335
rect 95 250 145 265
rect 205 335 255 350
rect 205 265 220 335
rect 240 265 255 335
rect 205 250 255 265
rect 315 335 365 350
rect 315 265 330 335
rect 350 265 365 335
rect 315 250 365 265
<< ndiffc >>
rect -3035 25 -3015 95
rect -2970 25 -2950 95
rect -2890 25 -2870 95
rect -2825 25 -2805 95
rect -2745 25 -2725 95
rect -2680 25 -2660 95
rect -2600 25 -2580 95
rect -2535 25 -2515 95
rect -2455 25 -2435 95
rect -2390 25 -2370 95
rect -2310 25 -2290 95
rect -2245 25 -2225 95
rect -2165 25 -2145 95
rect -2100 25 -2080 95
rect -2020 25 -2000 95
rect -1955 25 -1935 95
rect -1875 25 -1855 95
rect -1810 25 -1790 95
rect -1540 15 -1520 85
rect -1430 15 -1410 85
rect -1320 15 -1300 85
rect -1210 15 -1190 85
rect -1100 15 -1080 85
rect -880 15 -860 85
rect -770 15 -750 85
rect -660 15 -640 85
rect -550 15 -530 85
rect -440 15 -420 85
rect -110 15 -90 85
rect 0 15 20 85
rect 110 15 130 85
rect 220 15 240 85
rect 330 15 350 85
<< pdiffc >>
rect -3035 255 -3015 425
rect -2970 255 -2950 425
rect -2890 255 -2870 425
rect -2825 255 -2805 425
rect -2745 255 -2725 425
rect -2680 255 -2660 425
rect -2600 255 -2580 425
rect -2535 255 -2515 425
rect -2455 255 -2435 425
rect -2390 255 -2370 425
rect -2310 255 -2290 425
rect -2245 255 -2225 425
rect -2165 255 -2145 425
rect -2100 255 -2080 425
rect -2020 255 -2000 425
rect -1955 255 -1935 425
rect -1875 255 -1855 425
rect -1810 255 -1790 425
rect -1590 265 -1570 335
rect -1480 265 -1460 335
rect -1370 265 -1350 335
rect -1260 265 -1240 335
rect -1150 265 -1130 335
rect -1040 265 -1020 335
rect -930 265 -910 335
rect -820 265 -800 335
rect -710 265 -690 335
rect -550 265 -530 335
rect -440 265 -420 335
rect -330 265 -310 335
rect -220 265 -200 335
rect -110 265 -90 335
rect 0 265 20 335
rect 110 265 130 335
rect 220 265 240 335
rect 330 265 350 335
<< psubdiff >>
rect -2590 -40 -2490 -25
rect -2590 -60 -2575 -40
rect -2505 -60 -2490 -40
rect -2590 -75 -2490 -60
rect -1030 85 -980 100
rect -1030 15 -1015 85
rect -995 15 -980 85
rect -1030 0 -980 15
rect -375 85 -325 100
rect -375 15 -360 85
rect -340 15 -325 85
rect -375 0 -325 15
<< nsubdiff >>
rect -2380 510 -2180 525
rect -2380 490 -2365 510
rect -2195 490 -2180 510
rect -2380 475 -2180 490
rect -645 335 -595 350
rect -645 265 -630 335
rect -610 265 -595 335
rect -645 250 -595 265
<< psubdiffcont >>
rect -2575 -60 -2505 -40
rect -1015 15 -995 85
rect -360 15 -340 85
<< nsubdiffcont >>
rect -2365 490 -2195 510
rect -630 265 -610 335
<< poly >>
rect 435 875 475 885
rect -2670 860 445 875
rect -2670 700 -2655 860
rect 435 855 445 860
rect 465 855 475 875
rect 435 845 475 855
rect -2690 690 -2650 700
rect -2690 670 -2680 690
rect -2660 670 -2650 690
rect -2690 660 -2650 670
rect -2610 690 -1615 700
rect -2610 670 -2600 690
rect -2580 685 -1615 690
rect -2580 670 -2570 685
rect -2610 660 -2570 670
rect -2530 650 -1655 660
rect -2530 630 -2520 650
rect -2500 645 -1655 650
rect -2500 630 -2490 645
rect -2530 620 -2490 630
rect -2710 580 -1825 595
rect -3000 440 -2985 455
rect -2855 440 -2840 455
rect -2710 440 -2695 580
rect -2565 440 -2550 455
rect -2420 440 -2405 455
rect -2275 440 -2260 455
rect -2130 440 -2115 455
rect -1985 440 -1970 455
rect -1840 440 -1825 580
rect -3000 185 -2985 240
rect -2855 200 -2840 240
rect -2710 200 -2695 240
rect -2565 225 -2550 240
rect -3065 170 -2985 185
rect -3000 110 -2985 170
rect -2880 190 -2840 200
rect -2880 170 -2870 190
rect -2850 170 -2840 190
rect -2880 160 -2840 170
rect -2735 190 -2695 200
rect -2735 170 -2725 190
rect -2705 170 -2695 190
rect -2670 215 -2550 225
rect -2670 195 -2660 215
rect -2640 210 -2550 215
rect -2640 195 -2630 210
rect -2670 185 -2630 195
rect -2735 160 -2695 170
rect -2855 110 -2840 160
rect -2710 135 -2695 160
rect -2710 120 -2550 135
rect -2710 110 -2695 120
rect -2565 110 -2550 120
rect -2420 110 -2405 240
rect -2275 230 -2260 240
rect -2355 215 -2260 230
rect -2235 215 -2195 225
rect -2130 215 -2115 240
rect -1985 215 -1970 240
rect -1840 225 -1825 240
rect -2355 165 -2340 215
rect -2235 195 -2225 215
rect -2205 200 -1860 215
rect -2205 195 -2195 200
rect -2235 190 -2195 195
rect -2380 155 -2340 165
rect -2195 160 -2155 165
rect -2380 135 -2370 155
rect -2350 135 -2340 155
rect -2380 125 -2340 135
rect -2275 155 -2155 160
rect -2275 145 -2185 155
rect -2275 110 -2260 145
rect -2195 135 -2185 145
rect -2165 135 -2155 155
rect -2195 125 -2155 135
rect -2130 110 -2115 200
rect -1875 165 -1860 200
rect -1670 195 -1655 645
rect -1630 235 -1615 685
rect -1555 350 -1495 365
rect -1445 350 -1385 365
rect -1335 350 -1275 365
rect -1225 350 -1165 365
rect -1115 350 -1055 365
rect -1005 350 -945 365
rect -895 350 -835 365
rect -785 350 -725 365
rect -515 350 -455 365
rect -405 350 -345 365
rect -295 350 -235 365
rect -185 350 -125 365
rect -75 350 -15 365
rect 35 350 95 365
rect 145 350 205 365
rect 255 350 315 365
rect -1555 240 -1495 250
rect -1445 240 -1385 250
rect -1335 240 -1275 250
rect -1225 240 -1165 250
rect -1115 240 -1055 250
rect -1005 240 -945 250
rect -895 240 -835 250
rect -785 240 -725 250
rect -1555 235 -725 240
rect -1630 220 -725 235
rect -515 240 -455 250
rect -405 240 -345 250
rect -295 240 -235 250
rect -185 240 -125 250
rect -75 240 -15 250
rect 35 240 95 250
rect 145 240 205 250
rect 255 240 315 250
rect 435 245 475 255
rect 435 240 445 245
rect -515 225 445 240
rect 465 225 475 245
rect -515 195 -500 225
rect 435 215 475 225
rect -1670 180 -500 195
rect -2090 150 -2050 160
rect -1875 150 -1825 165
rect -2090 130 -2080 150
rect -2060 135 -2050 150
rect -2060 130 -1970 135
rect -2090 120 -1970 130
rect -1985 110 -1970 120
rect -1840 110 -1825 150
rect -1550 145 -1510 155
rect -1550 135 -1540 145
rect -1755 125 -1540 135
rect -1520 135 -1510 145
rect -1330 145 -1290 155
rect -1330 135 -1320 145
rect -1520 125 -1320 135
rect -1300 135 -1290 145
rect -1110 145 -1070 155
rect -1110 135 -1100 145
rect -1300 125 -1100 135
rect -1080 135 -1070 145
rect -1080 125 -455 135
rect 435 125 475 135
rect -1755 110 -455 125
rect -3000 -5 -2985 10
rect -2855 -5 -2840 10
rect -2710 -5 -2695 10
rect -2565 -5 -2550 10
rect -2420 -120 -2405 10
rect -2275 -5 -2260 10
rect -2130 -5 -2115 10
rect -1985 -5 -1970 10
rect -1840 -5 -1825 10
rect -1945 -15 -1905 -5
rect -1945 -35 -1935 -15
rect -1915 -30 -1905 -15
rect -1755 -30 -1740 110
rect -1505 100 -1445 110
rect -1395 100 -1335 110
rect -1285 100 -1225 110
rect -1175 100 -1115 110
rect -845 100 -785 110
rect -735 100 -675 110
rect -625 100 -565 110
rect -515 100 -455 110
rect -170 110 445 125
rect -1505 -15 -1445 0
rect -1395 -15 -1335 0
rect -1285 -15 -1225 0
rect -1175 -15 -1115 0
rect -845 -15 -785 0
rect -735 -15 -675 0
rect -625 -15 -565 0
rect -515 -15 -455 0
rect -1915 -35 -1740 -30
rect -1945 -45 -1740 -35
rect -2040 -80 -1725 -70
rect -2040 -100 -2030 -80
rect -2010 -85 -1810 -80
rect -2010 -100 -2000 -85
rect -2040 -110 -2000 -100
rect -1820 -100 -1810 -85
rect -1790 -85 -1725 -80
rect -1790 -100 -1780 -85
rect -1820 -110 -1780 -100
rect -3065 -135 -2405 -120
rect -1740 -120 -1725 -85
rect -170 -120 -155 110
rect -75 100 -15 110
rect 35 100 95 110
rect 145 100 205 110
rect 255 100 315 110
rect 435 105 445 110
rect 465 105 475 125
rect 435 95 475 105
rect -75 -15 -15 0
rect 35 -15 95 0
rect 145 -15 205 0
rect 255 -15 315 0
rect -2120 -135 -2080 -125
rect -1740 -135 -155 -120
rect -2120 -155 -2110 -135
rect -2090 -150 -2080 -135
rect -2090 -155 -1805 -150
rect -2120 -160 -1805 -155
rect 435 -155 475 -145
rect 435 -160 445 -155
rect -2120 -165 445 -160
rect -1820 -175 445 -165
rect 465 -175 475 -155
rect 435 -185 475 -175
<< polycont >>
rect 445 855 465 875
rect -2680 670 -2660 690
rect -2600 670 -2580 690
rect -2520 630 -2500 650
rect -2870 170 -2850 190
rect -2725 170 -2705 190
rect -2660 195 -2640 215
rect -2225 195 -2205 215
rect -2370 135 -2350 155
rect -2185 135 -2165 155
rect 445 225 465 245
rect -2080 130 -2060 150
rect -1540 125 -1520 145
rect -1320 125 -1300 145
rect -1100 125 -1080 145
rect -1935 -35 -1915 -15
rect -2030 -100 -2010 -80
rect -1810 -100 -1790 -80
rect 445 105 465 125
rect -2110 -155 -2090 -135
rect 445 -175 465 -155
<< locali >>
rect 515 890 570 900
rect 435 875 475 885
rect 515 875 525 890
rect 435 855 445 875
rect 465 855 525 875
rect 560 855 570 890
rect 435 845 475 855
rect 515 845 570 855
rect -2690 690 -2650 700
rect -2690 670 -2680 690
rect -2660 670 -2650 690
rect -2690 660 -2650 670
rect -2670 435 -2650 660
rect -3045 425 -3005 435
rect -3045 255 -3035 425
rect -3015 255 -3005 425
rect -3045 245 -3005 255
rect -2980 425 -2940 435
rect -2980 255 -2970 425
rect -2950 255 -2940 425
rect -2980 245 -2940 255
rect -2900 425 -2860 435
rect -2900 255 -2890 425
rect -2870 255 -2860 425
rect -2900 245 -2860 255
rect -2835 425 -2795 435
rect -2835 255 -2825 425
rect -2805 255 -2795 425
rect -2835 245 -2795 255
rect -2755 425 -2715 435
rect -2755 255 -2745 425
rect -2725 255 -2715 425
rect -2755 245 -2715 255
rect -2690 425 -2650 435
rect -2690 255 -2680 425
rect -2660 255 -2650 425
rect -2690 245 -2650 255
rect -2610 690 -2570 700
rect -2610 670 -2600 690
rect -2580 670 -2570 690
rect -2610 660 -2570 670
rect -2610 435 -2590 660
rect -2530 650 -2490 660
rect -2530 630 -2520 650
rect -2500 630 -2490 650
rect -2530 620 -2490 630
rect -2530 435 -2510 620
rect -2375 510 -2185 520
rect -2375 490 -2365 510
rect -2195 490 -2185 510
rect -2375 480 -2185 490
rect -2610 425 -2570 435
rect -2610 255 -2600 425
rect -2580 255 -2570 425
rect -2610 245 -2570 255
rect -2545 425 -2505 435
rect -2545 255 -2535 425
rect -2515 255 -2505 425
rect -2545 245 -2505 255
rect -2465 425 -2425 435
rect -2465 255 -2455 425
rect -2435 255 -2425 425
rect -2465 245 -2425 255
rect -2400 425 -2360 435
rect -2400 255 -2390 425
rect -2370 275 -2360 425
rect -2320 425 -2280 435
rect -2370 255 -2355 275
rect -2400 245 -2355 255
rect -2320 255 -2310 425
rect -2290 255 -2280 425
rect -2320 245 -2280 255
rect -2255 425 -2215 435
rect -2255 255 -2245 425
rect -2225 255 -2215 425
rect -2255 245 -2215 255
rect -2175 425 -2135 435
rect -2175 255 -2165 425
rect -2145 255 -2135 425
rect -2175 245 -2135 255
rect -2110 425 -2070 435
rect -2110 255 -2100 425
rect -2080 255 -2070 425
rect -2110 245 -2070 255
rect -2030 425 -1990 435
rect -2030 255 -2020 425
rect -2000 255 -1990 425
rect -2030 245 -1990 255
rect -1965 425 -1925 435
rect -1965 255 -1955 425
rect -1935 255 -1925 425
rect -1965 245 -1925 255
rect -1885 425 -1845 435
rect -1885 255 -1875 425
rect -1855 255 -1845 425
rect -1885 245 -1845 255
rect -1820 425 -1780 435
rect -1820 255 -1810 425
rect -1790 255 -1780 425
rect -1590 365 -690 385
rect -1590 345 -1570 365
rect -1370 345 -1350 365
rect -1150 345 -1130 365
rect -930 345 -910 365
rect -710 345 -690 365
rect -550 365 350 385
rect -550 345 -530 365
rect -330 345 -310 365
rect -110 345 -90 365
rect 110 345 130 365
rect 330 345 350 365
rect -1600 335 -1560 345
rect -1600 265 -1590 335
rect -1570 265 -1560 335
rect -1600 255 -1560 265
rect -1490 335 -1450 345
rect -1490 265 -1480 335
rect -1460 265 -1450 335
rect -1490 255 -1450 265
rect -1380 335 -1340 345
rect -1380 265 -1370 335
rect -1350 265 -1340 335
rect -1380 255 -1340 265
rect -1270 335 -1230 345
rect -1270 265 -1260 335
rect -1240 265 -1230 335
rect -1270 255 -1230 265
rect -1160 335 -1120 345
rect -1160 265 -1150 335
rect -1130 265 -1120 335
rect -1160 255 -1120 265
rect -1050 335 -1010 345
rect -1050 265 -1040 335
rect -1020 265 -1010 335
rect -1050 255 -1010 265
rect -940 335 -900 345
rect -940 265 -930 335
rect -910 265 -900 335
rect -940 255 -900 265
rect -830 335 -790 345
rect -830 265 -820 335
rect -800 265 -790 335
rect -830 255 -790 265
rect -720 335 -680 345
rect -720 265 -710 335
rect -690 265 -680 335
rect -720 255 -680 265
rect -640 335 -600 345
rect -640 265 -630 335
rect -610 265 -600 335
rect -640 255 -600 265
rect -560 335 -520 345
rect -560 265 -550 335
rect -530 265 -520 335
rect -560 255 -520 265
rect -450 335 -410 345
rect -450 265 -440 335
rect -420 265 -410 335
rect -450 255 -410 265
rect -340 335 -300 345
rect -340 265 -330 335
rect -310 265 -300 335
rect -340 255 -300 265
rect -230 335 -190 345
rect -230 265 -220 335
rect -200 265 -190 335
rect -230 255 -190 265
rect -120 335 -80 345
rect -120 265 -110 335
rect -90 265 -80 335
rect -120 255 -80 265
rect -10 335 30 345
rect -10 265 0 335
rect 20 265 30 335
rect -10 255 30 265
rect 100 335 140 345
rect 100 265 110 335
rect 130 265 140 335
rect 100 255 140 265
rect 210 335 250 345
rect 210 265 220 335
rect 240 265 250 335
rect 210 255 250 265
rect 320 335 360 345
rect 320 265 330 335
rect 350 265 360 335
rect 320 255 360 265
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect -1820 245 -1780 255
rect -2960 190 -2940 245
rect -2880 190 -2840 200
rect -2960 170 -2870 190
rect -2850 170 -2840 190
rect -2960 105 -2940 170
rect -2880 160 -2840 170
rect -2815 190 -2795 245
rect -2670 225 -2650 245
rect -2670 215 -2630 225
rect -2735 190 -2695 200
rect -2815 170 -2725 190
rect -2705 170 -2695 190
rect -2815 105 -2795 170
rect -2735 160 -2695 170
rect -2670 195 -2660 215
rect -2640 195 -2630 215
rect -2670 185 -2630 195
rect -2670 105 -2650 185
rect -2600 105 -2580 245
rect -2545 105 -2525 245
rect -2445 225 -2425 245
rect -2310 225 -2290 245
rect -2445 205 -2290 225
rect -2445 105 -2425 205
rect -2380 155 -2340 165
rect -2380 135 -2370 155
rect -2350 135 -2340 155
rect -2380 125 -2340 135
rect -2380 105 -2360 125
rect -2310 105 -2290 205
rect -2245 225 -2225 245
rect -2245 215 -2195 225
rect -2245 195 -2225 215
rect -2205 195 -2195 215
rect -2245 190 -2195 195
rect -2245 105 -2225 190
rect -2170 165 -2150 245
rect -2195 155 -2150 165
rect -2195 135 -2185 155
rect -2165 135 -2150 155
rect -2195 125 -2150 135
rect -2090 160 -2070 245
rect -2090 150 -2050 160
rect -2090 130 -2080 150
rect -2060 130 -2050 150
rect -2090 120 -2050 130
rect -2090 105 -2070 120
rect -2020 105 -2000 245
rect -1955 105 -1935 245
rect -710 225 -690 255
rect -710 205 -640 225
rect -1550 145 -1510 155
rect -1550 125 -1540 145
rect -1520 125 -1510 145
rect -1550 115 -1510 125
rect -1330 145 -1290 155
rect -1330 125 -1320 145
rect -1300 125 -1290 145
rect -1330 115 -1290 125
rect -1110 145 -1070 155
rect -1110 125 -1100 145
rect -1080 125 -1070 145
rect -1110 115 -1070 125
rect -3045 95 -3005 105
rect -3045 25 -3035 95
rect -3015 25 -3005 95
rect -3045 15 -3005 25
rect -2980 95 -2940 105
rect -2980 25 -2970 95
rect -2950 25 -2940 95
rect -2980 15 -2940 25
rect -2900 95 -2860 105
rect -2900 25 -2890 95
rect -2870 25 -2860 95
rect -2900 15 -2860 25
rect -2835 95 -2795 105
rect -2835 25 -2825 95
rect -2805 25 -2795 95
rect -2835 15 -2795 25
rect -2755 95 -2715 105
rect -2755 25 -2745 95
rect -2725 25 -2715 95
rect -2755 15 -2715 25
rect -2690 95 -2650 105
rect -2690 25 -2680 95
rect -2660 25 -2650 95
rect -2690 15 -2650 25
rect -2610 95 -2570 105
rect -2610 25 -2600 95
rect -2580 25 -2570 95
rect -2610 15 -2570 25
rect -2545 95 -2505 105
rect -2545 25 -2535 95
rect -2515 25 -2505 95
rect -2545 15 -2505 25
rect -2465 95 -2425 105
rect -2465 25 -2455 95
rect -2435 25 -2425 95
rect -2465 15 -2425 25
rect -2400 95 -2360 105
rect -2400 25 -2390 95
rect -2370 25 -2360 95
rect -2400 15 -2360 25
rect -2320 95 -2280 105
rect -2320 25 -2310 95
rect -2290 25 -2280 95
rect -2320 15 -2280 25
rect -2255 95 -2215 105
rect -2255 25 -2245 95
rect -2225 25 -2215 95
rect -2255 15 -2215 25
rect -2175 95 -2135 105
rect -2175 25 -2165 95
rect -2145 25 -2135 95
rect -2175 15 -2135 25
rect -2110 95 -2070 105
rect -2110 25 -2100 95
rect -2080 25 -2070 95
rect -2110 15 -2070 25
rect -2030 95 -1990 105
rect -2030 25 -2020 95
rect -2000 25 -1990 95
rect -2030 15 -1990 25
rect -1965 95 -1920 105
rect -1965 25 -1955 95
rect -1935 25 -1920 95
rect -1965 15 -1920 25
rect -1885 95 -1845 105
rect -1885 25 -1875 95
rect -1855 25 -1845 95
rect -1885 15 -1845 25
rect -1820 95 -1780 105
rect -1540 95 -1520 115
rect -1320 95 -1300 115
rect -1100 95 -1080 115
rect -660 95 -640 205
rect 330 185 350 255
rect 435 250 475 255
rect 515 250 570 260
rect 435 245 540 250
rect 435 225 445 245
rect 465 230 540 245
rect 465 225 475 230
rect 435 215 475 225
rect 330 165 1250 185
rect 330 95 350 165
rect 435 125 475 135
rect 435 105 445 125
rect 465 120 475 125
rect 465 105 550 120
rect 435 100 550 105
rect 435 95 475 100
rect -1820 25 -1810 95
rect -1790 25 -1780 95
rect -1820 15 -1780 25
rect -1550 85 -1510 95
rect -1550 15 -1540 85
rect -1520 15 -1510 85
rect -2585 -40 -2495 -30
rect -2585 -60 -2575 -40
rect -2505 -60 -2495 -40
rect -2585 -70 -2495 -60
rect -2100 -125 -2080 15
rect -2020 -70 -2000 15
rect -1945 -5 -1925 15
rect -1945 -15 -1905 -5
rect -1945 -35 -1935 -15
rect -1915 -35 -1905 -15
rect -1945 -45 -1905 -35
rect -1810 -70 -1790 15
rect -1550 5 -1510 15
rect -1440 85 -1400 95
rect -1440 15 -1430 85
rect -1410 15 -1400 85
rect -1440 5 -1400 15
rect -1330 85 -1290 95
rect -1330 15 -1320 85
rect -1300 15 -1290 85
rect -1330 5 -1290 15
rect -1220 85 -1180 95
rect -1220 15 -1210 85
rect -1190 15 -1180 85
rect -1220 5 -1180 15
rect -1110 85 -1070 95
rect -1110 15 -1100 85
rect -1080 15 -1070 85
rect -1110 5 -1070 15
rect -1025 85 -985 95
rect -1025 15 -1015 85
rect -995 15 -985 85
rect -1025 5 -985 15
rect -890 85 -850 95
rect -890 15 -880 85
rect -860 15 -850 85
rect -890 5 -850 15
rect -780 85 -740 95
rect -780 15 -770 85
rect -750 15 -740 85
rect -780 5 -740 15
rect -670 85 -630 95
rect -670 15 -660 85
rect -640 15 -630 85
rect -670 5 -630 15
rect -560 85 -520 95
rect -560 15 -550 85
rect -530 15 -520 85
rect -560 5 -520 15
rect -450 85 -410 95
rect -450 15 -440 85
rect -420 15 -410 85
rect -450 5 -410 15
rect -370 85 -330 95
rect -370 15 -360 85
rect -340 15 -330 85
rect -370 5 -330 15
rect -120 85 -80 95
rect -120 15 -110 85
rect -90 15 -80 85
rect -120 5 -80 15
rect -10 85 30 95
rect -10 15 0 85
rect 20 15 30 85
rect -10 5 30 15
rect 100 85 140 95
rect 100 15 110 85
rect 130 15 140 85
rect 100 5 140 15
rect 210 85 250 95
rect 210 15 220 85
rect 240 15 250 85
rect 210 5 250 15
rect 320 85 360 95
rect 320 15 330 85
rect 350 15 360 85
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect 320 5 360 15
rect -1540 -15 -1520 5
rect -1320 -15 -1300 5
rect -1100 -15 -1080 5
rect -1710 -35 -1080 -15
rect -880 -15 -860 5
rect -660 -15 -640 5
rect -440 -15 -420 5
rect -880 -35 -420 -15
rect -110 -15 -90 5
rect 110 -15 130 5
rect 330 -15 350 5
rect -110 -35 350 -15
rect -2040 -80 -2000 -70
rect -2040 -100 -2030 -80
rect -2010 -100 -2000 -80
rect -2040 -110 -2000 -100
rect -1820 -80 -1780 -70
rect -1820 -100 -1810 -80
rect -1790 -100 -1780 -80
rect -1820 -110 -1780 -100
rect -2120 -135 -2080 -125
rect -2120 -155 -2110 -135
rect -2090 -155 -2080 -135
rect -2120 -165 -2080 -155
rect -1710 -210 -1690 -35
rect 515 -130 570 -120
rect 435 -155 475 -145
rect 515 -155 525 -130
rect 435 -175 445 -155
rect 465 -165 525 -155
rect 560 -165 570 -130
rect 465 -175 570 -165
rect 435 -185 475 -175
rect -3065 -230 -1690 -210
<< viali >>
rect 525 855 560 890
rect -3035 255 -3015 425
rect -2890 255 -2870 425
rect -2745 255 -2725 425
rect -2365 490 -2195 510
rect -2390 255 -2370 425
rect -2165 255 -2145 425
rect -1875 255 -1855 425
rect -1480 265 -1460 335
rect -1260 265 -1240 335
rect -1040 265 -1020 335
rect -820 265 -800 335
rect -630 265 -610 335
rect -440 265 -420 335
rect -220 265 -200 335
rect 0 265 20 335
rect 220 265 240 335
rect 525 260 560 295
rect -3035 25 -3015 95
rect -2890 25 -2870 95
rect -2745 25 -2725 95
rect -2390 25 -2370 95
rect -2165 25 -2145 95
rect -1875 25 -1855 95
rect -2575 -60 -2505 -40
rect -1430 15 -1410 85
rect -1210 15 -1190 85
rect -1015 15 -995 85
rect -770 15 -750 85
rect -550 15 -530 85
rect -360 15 -340 85
rect 0 15 20 85
rect 220 15 240 85
rect 525 55 560 90
rect 525 -165 560 -130
<< metal1 >>
rect 515 890 570 900
rect 515 855 525 890
rect 560 855 570 890
rect 515 845 570 855
rect -2380 510 -2180 525
rect -2380 490 -2365 510
rect -2195 490 -2180 510
rect -2380 440 -2180 490
rect -3100 425 365 440
rect -3100 255 -3035 425
rect -3015 255 -2890 425
rect -2870 255 -2745 425
rect -2725 255 -2390 425
rect -2370 255 -2165 425
rect -2145 255 -1875 425
rect -1855 335 365 425
rect -1855 265 -1480 335
rect -1460 265 -1260 335
rect -1240 265 -1040 335
rect -1020 265 -820 335
rect -800 265 -630 335
rect -610 265 -440 335
rect -420 265 -220 335
rect -200 265 0 335
rect 20 265 220 335
rect 240 265 365 335
rect -1855 255 365 265
rect -3100 240 365 255
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect 515 250 570 260
rect -3100 95 365 110
rect -3100 25 -3035 95
rect -3015 25 -2890 95
rect -2870 25 -2745 95
rect -2725 25 -2390 95
rect -2370 25 -2165 95
rect -2145 25 -1875 95
rect -1855 85 365 95
rect -1855 25 -1430 85
rect -3100 15 -1430 25
rect -1410 15 -1210 85
rect -1190 15 -1015 85
rect -995 15 -770 85
rect -750 15 -550 85
rect -530 15 -360 85
rect -340 15 0 85
rect 20 15 220 85
rect 240 15 365 85
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect -3100 0 365 15
rect -2590 -40 -2485 0
rect -2590 -60 -2575 -40
rect -2505 -60 -2485 -40
rect -2590 -75 -2485 -60
rect 515 -130 570 -120
rect 515 -165 525 -130
rect 560 -165 570 -130
rect 515 -175 570 -165
<< via1 >>
rect 525 855 560 890
rect 525 260 560 295
rect 525 55 560 90
rect 525 -165 560 -130
<< metal2 >>
rect 515 890 570 900
rect 515 855 525 890
rect 560 855 570 890
rect 515 845 570 855
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect 515 250 570 260
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect 515 -130 570 -120
rect 515 -165 525 -130
rect 560 -165 570 -130
rect 515 -175 570 -165
<< via2 >>
rect 525 855 560 890
rect 525 260 560 295
rect 525 55 560 90
rect 525 -165 560 -130
<< metal3 >>
rect 690 900 1140 925
rect 515 890 1140 900
rect 515 855 525 890
rect 560 855 1140 890
rect 515 845 1140 855
rect 690 305 1140 845
rect 515 295 1140 305
rect 515 260 525 295
rect 560 260 1140 295
rect 515 250 1140 260
rect 690 235 1140 250
rect 690 100 980 115
rect 515 90 980 100
rect 515 55 525 90
rect 560 55 980 90
rect 515 45 980 55
rect 690 -120 980 45
rect 515 -130 980 -120
rect 515 -165 525 -130
rect 560 -165 980 -130
rect 515 -175 980 -165
<< via3 >>
rect 525 260 560 295
rect 525 55 560 90
<< mimcap >>
rect 705 295 1125 910
rect 705 260 715 295
rect 750 260 1125 295
rect 705 250 1125 260
rect 705 90 965 100
rect 705 55 715 90
rect 750 55 965 90
rect 705 -160 965 55
<< mimcapcontact >>
rect 715 260 750 295
rect 715 55 750 90
<< metal4 >>
rect 515 295 760 305
rect 515 260 525 295
rect 560 260 715 295
rect 750 260 760 295
rect 515 250 760 260
rect 515 90 760 100
rect 515 55 525 90
rect 560 55 715 90
rect 750 55 760 90
rect 515 45 760 55
<< labels >>
flabel locali -3065 -220 -3065 -220 7 FreeSans 400 0 -200 0 I_IN
flabel poly -3065 -125 -3065 -125 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel poly -3065 175 -3065 175 7 FreeSans 400 0 -200 0 UP_PFD
flabel metal1 -3100 340 -3100 340 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 -3100 60 -3100 60 7 FreeSans 400 0 -200 0 GNDA
flabel locali 1250 175 1250 175 3 FreeSans 400 0 80 0 VOUT
flabel poly -1620 590 -1615 590 3 FreeSans 400 0 200 0 OPAMP_OUT
flabel poly -2130 -5 -2130 -5 7 FreeSans 400 0 -200 -200 DOWN_b
flabel poly -500 190 -500 190 3 FreeSans 400 0 200 0 UP_input
flabel poly -2670 820 -2670 820 7 FreeSans 400 0 -200 0 UP_b
flabel poly -2120 -165 -2120 -165 7 FreeSans 400 0 -200 -200 DOWN
flabel poly -155 -135 -155 -135 3 FreeSans 400 0 200 0 DOWN_input
flabel poly -2710 595 -2710 595 7 FreeSans 400 0 -200 0 UP
<< end >>
