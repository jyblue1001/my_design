* PEX produced on Tue Feb 18 05:55:46 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from div120_2.ext - technology: sky130A

.subckt div120_2 VOUT VIN VDDA GNDA
X0 div2_4_1.C.t3 div2_4_1.A.t2 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1 div5_2_0.D.t2 div5_2_0.B.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X2 GNDA.t43 div5_2_0.Q2_b.t2 div5_2_0.M.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 div3_3_0.CLK.t2 div8.t2 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 VDDA.t76 div24.t3 div3_3_0.A.t0 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X5 GNDA.t6 div2.t2 a_1320_n1010.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 GNDA.t4 div3_3_0.I.t2 div3_3_0.G.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X7 VDDA.t40 VIN.t0 a_20_n1010.t2 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X8 VDDA.t17 div4.t2 a_2620_n1010.t2 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X9 div2_4_1.B.t1 div2.t3 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X10 GNDA.t31 a_20_n1010.t3 div2_4_1.C.t2 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 div2_4_0.A.t0 a_2620_n1010.t3 div2_4_0.B.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X12 div3_3_0.F.t1 div3_3_0.CLK.t3 div3_3_0.E.t2 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X13 div3_3_0.I.t0 div3_3_0.H.t4 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 div5_2_0.A.t0 div5_2_0.Q2_b.t3 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X15 GNDA.t53 div24.t4 div5_2_0.D.t1 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X16 div8.t0 a_2620_n1010.t4 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X17 VDDA.t38 div3_3_0.D.t2 div3_3_0.E.t0 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 div5_2_0.A.t2 div5_2_0.Q2_b.t4 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X19 GNDA.t57 div3_3_0.CLK.t4 div3_3_0.C.t3 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X20 GNDA.t88 div24.t5 div5_2_0.D.t3 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X21 GNDA.t50 div24.t6 div5_2_0.J.t3 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 div5_2_0.K.t0 div5_2_0.Q2_b.t5 div5_2_0.L.t1 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 GNDA.t38 div5_2_0.Q2_b.t6 div5_2_0.M.t1 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X24 div5_2_0.Q2_b.t1 div24.t7 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X25 div4.t0 div2_4_2.C.t4 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X26 GNDA.t12 a_2620_n1010.t5 div2_4_0.C.t2 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X27 GNDA.t90 div3_3_0.CLK.t5 div3_3_0.C.t2 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X28 a_1320_n1010.t2 div2.t4 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X29 div2_4_0.C.t3 div2_4_0.A.t2 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X30 div3_3_0.D.t1 div3_3_0.CLK.t6 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X31 VDDA.t36 VOUT.t2 div5_2_0.K.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X32 GNDA.t63 div3_3_0.CLK.t7 div3_3_0.H.t3 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X33 VDDA.t32 div4.t3 div2_4_2.A.t0 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X34 VOUT.t0 div5_2_0.Q2_b.t7 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X35 div2_4_2.A.t1 a_1320_n1010.t3 div2_4_2.B.t1 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X36 GNDA.t92 a_1320_n1010.t4 div2_4_2.C.t3 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X37 GNDA.t27 div5_2_0.E.t2 div5_2_0.I.t2 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X38 div5_2_0.G.t0 VOUT.t3 div5_2_0.F.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X39 GNDA.t8 VIN.t1 a_20_n1010.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X40 div2_4_1.C.t0 a_20_n1010.t4 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X41 div2_4_0.B.t1 div8.t3 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X42 GNDA.t103 div3_3_0.CLK.t8 div3_3_0.H.t2 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X43 div3_3_0.I.t1 div3_3_0.CLK.t9 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X44 div5_2_0.E.t1 div24.t8 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X45 div3_3_0.B.t0 div24.t9 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X46 div5_2_0.B.t1 div24.t10 div5_2_0.C.t1 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 GNDA.t98 div24.t11 div5_2_0.J.t2 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X48 div24.t2 div3_3_0.I.t3 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X49 VDDA.t54 div5_2_0.Q2_b.t8 div5_2_0.G.t1 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X50 VOUT.t1 div5_2_0.M.t4 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X51 a_20_n1010.t1 VIN.t2 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X52 a_2620_n1010.t1 div4.t4 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X53 div3_3_0.C.t0 div3_3_0.A.t2 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X54 VDDA.t24 div2.t5 div2_4_1.A.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X55 VDDA.t46 div8.t4 div3_3_0.CLK.t1 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X56 VDDA.t56 div5_2_0.A.t3 div5_2_0.B.t0 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X57 GNDA.t19 a_1320_n1010.t5 div2_4_2.C.t2 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X58 div3_3_0.G.t0 div3_3_0.D.t3 div3_3_0.F.t0 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X59 div5_2_0.E.t0 div5_2_0.D.t4 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X60 div3_3_0.E.t1 div3_3_0.I.t4 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X61 div2_4_0.C.t1 a_2620_n1010.t6 GNDA.t73 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X62 div5_2_0.J.t1 div24.t12 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X63 div3_3_0.D.t0 div3_3_0.C.t4 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X64 div5_2_0.D.t0 div24.t13 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X65 div5_2_0.M.t2 div5_2_0.Q2_b.t9 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 VDDA.t52 div5_2_0.Q2_b.t10 div5_2_0.A.t1 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X67 div2_4_2.B.t0 div4.t5 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X68 div5_2_0.H.t1 div24.t14 div5_2_0.G.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X69 div2_4_1.A.t1 a_20_n1010.t5 div2_4_1.B.t0 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X70 GNDA.t23 a_20_n1010.t6 div2_4_1.C.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X71 div2.t1 div2_4_1.C.t4 GNDA.t82 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X72 GNDA.t46 div4.t6 a_2620_n1010.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X73 div3_3_0.C.t1 div3_3_0.CLK.t10 GNDA.t94 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X74 div5_2_0.L.t0 VOUT.t4 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X75 VDDA.t1 div5_2_0.G.t3 div5_2_0.J.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X76 div5_2_0.M.t3 div5_2_0.K.t2 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X77 div2.t0 a_20_n1010.t7 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X78 div2_4_2.C.t0 div2_4_2.A.t2 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X79 div5_2_0.I.t0 VOUT.t5 GNDA.t76 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X80 div3_3_0.H.t1 div3_3_0.CLK.t11 GNDA.t96 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X81 VDDA.t11 div2.t6 a_1320_n1010.t1 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X82 VDDA.t42 div8.t5 div2_4_0.A.t1 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X83 div24.t0 div3_3_0.I.t5 GNDA.t21 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X84 div5_2_0.I.t1 div5_2_0.Q2_b.t11 div5_2_0.H.t0 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X85 VDDA.t22 div3_3_0.I.t6 div24.t1 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X86 div2_4_2.C.t1 a_1320_n1010.t6 GNDA.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X87 div3_3_0.A.t1 div3_3_0.CLK.t12 div3_3_0.B.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X88 div5_2_0.Q2_b.t0 div5_2_0.J.t4 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X89 div5_2_0.F.t1 div5_2_0.E.t3 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X90 GNDA.t10 a_2620_n1010.t7 div2_4_0.C.t0 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X91 div8.t1 div2_4_0.C.t4 GNDA.t67 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X92 div4.t1 a_1320_n1010.t7 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X93 VDDA.t66 div3_3_0.E.t3 div3_3_0.H.t0 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X94 GNDA.t71 div8.t6 div3_3_0.CLK.t0 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X95 div5_2_0.C.t0 div5_2_0.A.t4 GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 div2_4_1.A.n0 div2_4_1.A.t0 713.933
R1 div2_4_1.A.t1 div2_4_1.A.n0 337
R2 div2_4_1.A.n0 div2_4_1.A.t2 314.233
R3 VDDA.t53 VDDA.t29 2804.76
R4 VDDA.t35 VDDA.t67 2533.33
R5 VDDA.t71 VDDA.t37 2307.14
R6 VDDA.t33 VDDA.t45 2216.67
R7 VDDA.t14 VDDA.t16 2216.67
R8 VDDA.t8 VDDA.t10 2216.67
R9 VDDA.t69 VDDA.t57 2126.19
R10 VDDA.t49 VDDA.t55 1538.1
R11 VDDA.t0 VDDA.t18 1492.86
R12 VDDA.t47 VDDA.t65 1492.86
R13 VDDA.n58 VDDA.t61 1289.29
R14 VDDA.t2 VDDA.n117 1289.29
R15 VDDA.t21 VDDA.t51 1130.95
R16 VDDA.t73 VDDA.t75 1130.95
R17 VDDA.t4 VDDA.t41 1130.95
R18 VDDA.t12 VDDA.t31 1130.95
R19 VDDA.t23 VDDA.t59 1130.95
R20 VDDA.t6 VDDA.n119 927.381
R21 VDDA.t19 VDDA.n120 927.381
R22 VDDA.t27 VDDA.n122 927.381
R23 VDDA.n123 VDDA.t63 927.381
R24 VDDA.n3 VDDA.t58 726.734
R25 VDDA.n236 VDDA.t22 726.734
R26 VDDA.n124 VDDA.t9 663.801
R27 VDDA.n121 VDDA.t15 663.801
R28 VDDA.n24 VDDA.t34 663.801
R29 VDDA.n118 VDDA.t72 663.801
R30 VDDA.n116 VDDA.t30 663.801
R31 VDDA.n59 VDDA.t44 663.801
R32 VDDA.n131 VDDA.n130 647.933
R33 VDDA.n137 VDDA.n127 647.933
R34 VDDA.n40 VDDA.n39 647.933
R35 VDDA.n38 VDDA.n37 647.933
R36 VDDA.n174 VDDA.n30 647.933
R37 VDDA.n180 VDDA.n27 647.933
R38 VDDA.n20 VDDA.n19 647.933
R39 VDDA.n18 VDDA.n17 647.933
R40 VDDA.n217 VDDA.n10 647.933
R41 VDDA.n224 VDDA.n7 647.933
R42 VDDA.n101 VDDA.n98 647.933
R43 VDDA.n108 VDDA.n95 647.933
R44 VDDA.n71 VDDA.n70 647.933
R45 VDDA.n57 VDDA.n56 647.933
R46 VDDA.n83 VDDA.n49 646.715
R47 VDDA.n58 VDDA.t43 610.715
R48 VDDA.n117 VDDA.t29 610.715
R49 VDDA.n119 VDDA.t71 610.715
R50 VDDA.n120 VDDA.t33 610.715
R51 VDDA.n122 VDDA.t14 610.715
R52 VDDA.n123 VDDA.t8 610.715
R53 VDDA.t61 VDDA.t35 497.62
R54 VDDA.t67 VDDA.t0 497.62
R55 VDDA.t18 VDDA.t25 497.62
R56 VDDA.t25 VDDA.t53 497.62
R57 VDDA.t55 VDDA.t2 497.62
R58 VDDA.t51 VDDA.t49 497.62
R59 VDDA.t57 VDDA.t21 497.62
R60 VDDA.t65 VDDA.t69 497.62
R61 VDDA.t37 VDDA.t47 497.62
R62 VDDA.t75 VDDA.t6 497.62
R63 VDDA.t45 VDDA.t73 497.62
R64 VDDA.t41 VDDA.t19 497.62
R65 VDDA.t16 VDDA.t4 497.62
R66 VDDA.t31 VDDA.t27 497.62
R67 VDDA.t10 VDDA.t12 497.62
R68 VDDA.t63 VDDA.t23 497.62
R69 VDDA.t59 VDDA.t39 497.62
R70 VDDA.n124 VDDA.n123 382.8
R71 VDDA.n122 VDDA.n121 382.8
R72 VDDA.n120 VDDA.n24 382.8
R73 VDDA.n119 VDDA.n118 382.8
R74 VDDA.n117 VDDA.n116 382.8
R75 VDDA.n59 VDDA.n58 382.8
R76 VDDA.n130 VDDA.t60 78.8005
R77 VDDA.n130 VDDA.t40 78.8005
R78 VDDA.n127 VDDA.t64 78.8005
R79 VDDA.n127 VDDA.t24 78.8005
R80 VDDA.n39 VDDA.t13 78.8005
R81 VDDA.n39 VDDA.t11 78.8005
R82 VDDA.n37 VDDA.t28 78.8005
R83 VDDA.n37 VDDA.t32 78.8005
R84 VDDA.n30 VDDA.t5 78.8005
R85 VDDA.n30 VDDA.t17 78.8005
R86 VDDA.n27 VDDA.t20 78.8005
R87 VDDA.n27 VDDA.t42 78.8005
R88 VDDA.n19 VDDA.t74 78.8005
R89 VDDA.n19 VDDA.t46 78.8005
R90 VDDA.n17 VDDA.t7 78.8005
R91 VDDA.n17 VDDA.t76 78.8005
R92 VDDA.n10 VDDA.t48 78.8005
R93 VDDA.n10 VDDA.t38 78.8005
R94 VDDA.n7 VDDA.t70 78.8005
R95 VDDA.n7 VDDA.t66 78.8005
R96 VDDA.n98 VDDA.t50 78.8005
R97 VDDA.n98 VDDA.t52 78.8005
R98 VDDA.n95 VDDA.t3 78.8005
R99 VDDA.n95 VDDA.t56 78.8005
R100 VDDA.n49 VDDA.t26 78.8005
R101 VDDA.n49 VDDA.t54 78.8005
R102 VDDA.n70 VDDA.t68 78.8005
R103 VDDA.n70 VDDA.t1 78.8005
R104 VDDA.n56 VDDA.t62 78.8005
R105 VDDA.n56 VDDA.t36 78.8005
R106 VDDA.n60 VDDA.n59 66.5733
R107 VDDA.n144 VDDA.n124 54.4005
R108 VDDA.n121 VDDA.n33 54.4005
R109 VDDA.n187 VDDA.n24 54.4005
R110 VDDA.n118 VDDA.n13 54.4005
R111 VDDA.n116 VDDA.n115 54.4005
R112 VDDA.n63 VDDA.n62 32.0005
R113 VDDA.n64 VDDA.n63 32.0005
R114 VDDA.n64 VDDA.n54 32.0005
R115 VDDA.n68 VDDA.n54 32.0005
R116 VDDA.n69 VDDA.n68 32.0005
R117 VDDA.n72 VDDA.n69 32.0005
R118 VDDA.n76 VDDA.n52 32.0005
R119 VDDA.n77 VDDA.n76 32.0005
R120 VDDA.n78 VDDA.n77 32.0005
R121 VDDA.n78 VDDA.n50 32.0005
R122 VDDA.n82 VDDA.n50 32.0005
R123 VDDA.n85 VDDA.n84 32.0005
R124 VDDA.n85 VDDA.n47 32.0005
R125 VDDA.n89 VDDA.n47 32.0005
R126 VDDA.n90 VDDA.n89 32.0005
R127 VDDA.n91 VDDA.n90 32.0005
R128 VDDA.n91 VDDA.n44 32.0005
R129 VDDA.n114 VDDA.n45 32.0005
R130 VDDA.n110 VDDA.n45 32.0005
R131 VDDA.n110 VDDA.n109 32.0005
R132 VDDA.n107 VDDA.n96 32.0005
R133 VDDA.n103 VDDA.n96 32.0005
R134 VDDA.n103 VDDA.n102 32.0005
R135 VDDA.n100 VDDA.n2 32.0005
R136 VDDA.n237 VDDA.n2 32.0005
R137 VDDA.n235 VDDA.n234 32.0005
R138 VDDA.n231 VDDA.n230 32.0005
R139 VDDA.n230 VDDA.n229 32.0005
R140 VDDA.n229 VDDA.n5 32.0005
R141 VDDA.n225 VDDA.n5 32.0005
R142 VDDA.n223 VDDA.n222 32.0005
R143 VDDA.n222 VDDA.n8 32.0005
R144 VDDA.n218 VDDA.n8 32.0005
R145 VDDA.n216 VDDA.n215 32.0005
R146 VDDA.n215 VDDA.n11 32.0005
R147 VDDA.n211 VDDA.n11 32.0005
R148 VDDA.n211 VDDA.n210 32.0005
R149 VDDA.n210 VDDA.n209 32.0005
R150 VDDA.n206 VDDA.n205 32.0005
R151 VDDA.n205 VDDA.n204 32.0005
R152 VDDA.n204 VDDA.n15 32.0005
R153 VDDA.n200 VDDA.n199 32.0005
R154 VDDA.n199 VDDA.n198 32.0005
R155 VDDA.n195 VDDA.n194 32.0005
R156 VDDA.n194 VDDA.n193 32.0005
R157 VDDA.n193 VDDA.n22 32.0005
R158 VDDA.n189 VDDA.n22 32.0005
R159 VDDA.n189 VDDA.n188 32.0005
R160 VDDA.n186 VDDA.n25 32.0005
R161 VDDA.n182 VDDA.n25 32.0005
R162 VDDA.n182 VDDA.n181 32.0005
R163 VDDA.n179 VDDA.n28 32.0005
R164 VDDA.n175 VDDA.n28 32.0005
R165 VDDA.n173 VDDA.n172 32.0005
R166 VDDA.n172 VDDA.n31 32.0005
R167 VDDA.n168 VDDA.n31 32.0005
R168 VDDA.n168 VDDA.n167 32.0005
R169 VDDA.n167 VDDA.n166 32.0005
R170 VDDA.n163 VDDA.n162 32.0005
R171 VDDA.n162 VDDA.n161 32.0005
R172 VDDA.n161 VDDA.n35 32.0005
R173 VDDA.n157 VDDA.n156 32.0005
R174 VDDA.n156 VDDA.n155 32.0005
R175 VDDA.n152 VDDA.n151 32.0005
R176 VDDA.n151 VDDA.n150 32.0005
R177 VDDA.n150 VDDA.n42 32.0005
R178 VDDA.n146 VDDA.n42 32.0005
R179 VDDA.n146 VDDA.n145 32.0005
R180 VDDA.n143 VDDA.n125 32.0005
R181 VDDA.n139 VDDA.n125 32.0005
R182 VDDA.n139 VDDA.n138 32.0005
R183 VDDA.n136 VDDA.n128 32.0005
R184 VDDA.n132 VDDA.n128 32.0005
R185 VDDA.n60 VDDA.n57 29.8684
R186 VDDA.n84 VDDA.n83 28.8005
R187 VDDA.n102 VDDA.n101 28.8005
R188 VDDA.n209 VDDA.n13 28.8005
R189 VDDA.n198 VDDA.n20 28.8005
R190 VDDA.n188 VDDA.n187 28.8005
R191 VDDA.n175 VDDA.n174 28.8005
R192 VDDA.n166 VDDA.n33 28.8005
R193 VDDA.n155 VDDA.n40 28.8005
R194 VDDA.n145 VDDA.n144 28.8005
R195 VDDA.n132 VDDA.n131 28.8005
R196 VDDA.n115 VDDA.n114 25.6005
R197 VDDA.n224 VDDA.n223 22.4005
R198 VDDA.n218 VDDA.n217 22.4005
R199 VDDA.n200 VDDA.n18 22.4005
R200 VDDA.n180 VDDA.n179 22.4005
R201 VDDA.n157 VDDA.n38 22.4005
R202 VDDA.n137 VDDA.n136 22.4005
R203 VDDA.n71 VDDA.n52 19.2005
R204 VDDA.n236 VDDA.n235 19.2005
R205 VDDA.n234 VDDA.n3 19.2005
R206 VDDA.n109 VDDA.n108 16.0005
R207 VDDA.n108 VDDA.n107 16.0005
R208 VDDA.n72 VDDA.n71 12.8005
R209 VDDA.n237 VDDA.n236 12.8005
R210 VDDA.n231 VDDA.n3 12.8005
R211 VDDA.n131 VDDA.n129 10.7683
R212 VDDA.n62 VDDA.n57 9.6005
R213 VDDA.n225 VDDA.n224 9.6005
R214 VDDA.n217 VDDA.n216 9.6005
R215 VDDA.n18 VDDA.n15 9.6005
R216 VDDA.n181 VDDA.n180 9.6005
R217 VDDA.n38 VDDA.n35 9.6005
R218 VDDA.n138 VDDA.n137 9.6005
R219 VDDA.n62 VDDA.n61 9.3005
R220 VDDA.n63 VDDA.n55 9.3005
R221 VDDA.n65 VDDA.n64 9.3005
R222 VDDA.n66 VDDA.n54 9.3005
R223 VDDA.n68 VDDA.n67 9.3005
R224 VDDA.n69 VDDA.n53 9.3005
R225 VDDA.n73 VDDA.n72 9.3005
R226 VDDA.n74 VDDA.n52 9.3005
R227 VDDA.n76 VDDA.n75 9.3005
R228 VDDA.n77 VDDA.n51 9.3005
R229 VDDA.n79 VDDA.n78 9.3005
R230 VDDA.n80 VDDA.n50 9.3005
R231 VDDA.n82 VDDA.n81 9.3005
R232 VDDA.n84 VDDA.n48 9.3005
R233 VDDA.n86 VDDA.n85 9.3005
R234 VDDA.n87 VDDA.n47 9.3005
R235 VDDA.n89 VDDA.n88 9.3005
R236 VDDA.n90 VDDA.n46 9.3005
R237 VDDA.n92 VDDA.n91 9.3005
R238 VDDA.n93 VDDA.n44 9.3005
R239 VDDA.n114 VDDA.n113 9.3005
R240 VDDA.n112 VDDA.n45 9.3005
R241 VDDA.n111 VDDA.n110 9.3005
R242 VDDA.n109 VDDA.n94 9.3005
R243 VDDA.n107 VDDA.n106 9.3005
R244 VDDA.n105 VDDA.n96 9.3005
R245 VDDA.n104 VDDA.n103 9.3005
R246 VDDA.n102 VDDA.n97 9.3005
R247 VDDA.n100 VDDA.n99 9.3005
R248 VDDA.n2 VDDA.n0 9.3005
R249 VDDA.n238 VDDA.n237 9.3005
R250 VDDA.n235 VDDA.n1 9.3005
R251 VDDA.n234 VDDA.n233 9.3005
R252 VDDA.n232 VDDA.n231 9.3005
R253 VDDA.n230 VDDA.n4 9.3005
R254 VDDA.n229 VDDA.n228 9.3005
R255 VDDA.n227 VDDA.n5 9.3005
R256 VDDA.n226 VDDA.n225 9.3005
R257 VDDA.n223 VDDA.n6 9.3005
R258 VDDA.n222 VDDA.n221 9.3005
R259 VDDA.n220 VDDA.n8 9.3005
R260 VDDA.n219 VDDA.n218 9.3005
R261 VDDA.n216 VDDA.n9 9.3005
R262 VDDA.n215 VDDA.n214 9.3005
R263 VDDA.n213 VDDA.n11 9.3005
R264 VDDA.n212 VDDA.n211 9.3005
R265 VDDA.n210 VDDA.n12 9.3005
R266 VDDA.n209 VDDA.n208 9.3005
R267 VDDA.n207 VDDA.n206 9.3005
R268 VDDA.n205 VDDA.n14 9.3005
R269 VDDA.n204 VDDA.n203 9.3005
R270 VDDA.n202 VDDA.n15 9.3005
R271 VDDA.n201 VDDA.n200 9.3005
R272 VDDA.n199 VDDA.n16 9.3005
R273 VDDA.n198 VDDA.n197 9.3005
R274 VDDA.n196 VDDA.n195 9.3005
R275 VDDA.n194 VDDA.n21 9.3005
R276 VDDA.n193 VDDA.n192 9.3005
R277 VDDA.n191 VDDA.n22 9.3005
R278 VDDA.n190 VDDA.n189 9.3005
R279 VDDA.n188 VDDA.n23 9.3005
R280 VDDA.n186 VDDA.n185 9.3005
R281 VDDA.n184 VDDA.n25 9.3005
R282 VDDA.n183 VDDA.n182 9.3005
R283 VDDA.n181 VDDA.n26 9.3005
R284 VDDA.n179 VDDA.n178 9.3005
R285 VDDA.n177 VDDA.n28 9.3005
R286 VDDA.n176 VDDA.n175 9.3005
R287 VDDA.n173 VDDA.n29 9.3005
R288 VDDA.n172 VDDA.n171 9.3005
R289 VDDA.n170 VDDA.n31 9.3005
R290 VDDA.n169 VDDA.n168 9.3005
R291 VDDA.n167 VDDA.n32 9.3005
R292 VDDA.n166 VDDA.n165 9.3005
R293 VDDA.n164 VDDA.n163 9.3005
R294 VDDA.n162 VDDA.n34 9.3005
R295 VDDA.n161 VDDA.n160 9.3005
R296 VDDA.n159 VDDA.n35 9.3005
R297 VDDA.n158 VDDA.n157 9.3005
R298 VDDA.n156 VDDA.n36 9.3005
R299 VDDA.n155 VDDA.n154 9.3005
R300 VDDA.n153 VDDA.n152 9.3005
R301 VDDA.n151 VDDA.n41 9.3005
R302 VDDA.n150 VDDA.n149 9.3005
R303 VDDA.n148 VDDA.n42 9.3005
R304 VDDA.n147 VDDA.n146 9.3005
R305 VDDA.n145 VDDA.n43 9.3005
R306 VDDA.n143 VDDA.n142 9.3005
R307 VDDA.n141 VDDA.n125 9.3005
R308 VDDA.n140 VDDA.n139 9.3005
R309 VDDA.n138 VDDA.n126 9.3005
R310 VDDA.n136 VDDA.n135 9.3005
R311 VDDA.n134 VDDA.n128 9.3005
R312 VDDA.n133 VDDA.n132 9.3005
R313 VDDA.n115 VDDA.n44 6.4005
R314 VDDA.n83 VDDA.n82 3.2005
R315 VDDA.n101 VDDA.n100 3.2005
R316 VDDA.n206 VDDA.n13 3.2005
R317 VDDA.n195 VDDA.n20 3.2005
R318 VDDA.n187 VDDA.n186 3.2005
R319 VDDA.n174 VDDA.n173 3.2005
R320 VDDA.n163 VDDA.n33 3.2005
R321 VDDA.n152 VDDA.n40 3.2005
R322 VDDA.n144 VDDA.n143 3.2005
R323 VDDA.n129 VDDA 0.25314
R324 VDDA.n61 VDDA.n60 0.224489
R325 VDDA.n133 VDDA.n129 0.185879
R326 VDDA.n61 VDDA.n55 0.15675
R327 VDDA.n65 VDDA.n55 0.15675
R328 VDDA.n66 VDDA.n65 0.15675
R329 VDDA.n67 VDDA.n66 0.15675
R330 VDDA.n67 VDDA.n53 0.15675
R331 VDDA.n73 VDDA.n53 0.15675
R332 VDDA.n74 VDDA.n73 0.15675
R333 VDDA.n75 VDDA.n74 0.15675
R334 VDDA.n75 VDDA.n51 0.15675
R335 VDDA.n79 VDDA.n51 0.15675
R336 VDDA.n80 VDDA.n79 0.15675
R337 VDDA.n81 VDDA.n80 0.15675
R338 VDDA.n81 VDDA.n48 0.15675
R339 VDDA.n86 VDDA.n48 0.15675
R340 VDDA.n87 VDDA.n86 0.15675
R341 VDDA.n88 VDDA.n87 0.15675
R342 VDDA.n88 VDDA.n46 0.15675
R343 VDDA.n92 VDDA.n46 0.15675
R344 VDDA.n93 VDDA.n92 0.15675
R345 VDDA.n113 VDDA.n93 0.15675
R346 VDDA.n113 VDDA.n112 0.15675
R347 VDDA.n112 VDDA.n111 0.15675
R348 VDDA.n111 VDDA.n94 0.15675
R349 VDDA.n106 VDDA.n94 0.15675
R350 VDDA.n106 VDDA.n105 0.15675
R351 VDDA.n105 VDDA.n104 0.15675
R352 VDDA.n104 VDDA.n97 0.15675
R353 VDDA.n99 VDDA.n97 0.15675
R354 VDDA.n99 VDDA.n0 0.15675
R355 VDDA.n238 VDDA.n1 0.15675
R356 VDDA.n233 VDDA.n1 0.15675
R357 VDDA.n233 VDDA.n232 0.15675
R358 VDDA.n232 VDDA.n4 0.15675
R359 VDDA.n228 VDDA.n4 0.15675
R360 VDDA.n228 VDDA.n227 0.15675
R361 VDDA.n227 VDDA.n226 0.15675
R362 VDDA.n226 VDDA.n6 0.15675
R363 VDDA.n221 VDDA.n6 0.15675
R364 VDDA.n221 VDDA.n220 0.15675
R365 VDDA.n220 VDDA.n219 0.15675
R366 VDDA.n219 VDDA.n9 0.15675
R367 VDDA.n214 VDDA.n9 0.15675
R368 VDDA.n214 VDDA.n213 0.15675
R369 VDDA.n213 VDDA.n212 0.15675
R370 VDDA.n212 VDDA.n12 0.15675
R371 VDDA.n208 VDDA.n12 0.15675
R372 VDDA.n208 VDDA.n207 0.15675
R373 VDDA.n207 VDDA.n14 0.15675
R374 VDDA.n203 VDDA.n14 0.15675
R375 VDDA.n203 VDDA.n202 0.15675
R376 VDDA.n202 VDDA.n201 0.15675
R377 VDDA.n201 VDDA.n16 0.15675
R378 VDDA.n197 VDDA.n16 0.15675
R379 VDDA.n197 VDDA.n196 0.15675
R380 VDDA.n196 VDDA.n21 0.15675
R381 VDDA.n192 VDDA.n191 0.15675
R382 VDDA.n191 VDDA.n190 0.15675
R383 VDDA.n190 VDDA.n23 0.15675
R384 VDDA.n185 VDDA.n23 0.15675
R385 VDDA.n185 VDDA.n184 0.15675
R386 VDDA.n184 VDDA.n183 0.15675
R387 VDDA.n183 VDDA.n26 0.15675
R388 VDDA.n178 VDDA.n26 0.15675
R389 VDDA.n178 VDDA.n177 0.15675
R390 VDDA.n177 VDDA.n176 0.15675
R391 VDDA.n176 VDDA.n29 0.15675
R392 VDDA.n171 VDDA.n29 0.15675
R393 VDDA.n170 VDDA.n169 0.15675
R394 VDDA.n169 VDDA.n32 0.15675
R395 VDDA.n165 VDDA.n32 0.15675
R396 VDDA.n165 VDDA.n164 0.15675
R397 VDDA.n164 VDDA.n34 0.15675
R398 VDDA.n160 VDDA.n34 0.15675
R399 VDDA.n160 VDDA.n159 0.15675
R400 VDDA.n159 VDDA.n158 0.15675
R401 VDDA.n158 VDDA.n36 0.15675
R402 VDDA.n154 VDDA.n36 0.15675
R403 VDDA.n154 VDDA.n153 0.15675
R404 VDDA.n153 VDDA.n41 0.15675
R405 VDDA.n149 VDDA.n148 0.15675
R406 VDDA.n148 VDDA.n147 0.15675
R407 VDDA.n147 VDDA.n43 0.15675
R408 VDDA.n142 VDDA.n43 0.15675
R409 VDDA.n142 VDDA.n141 0.15675
R410 VDDA.n141 VDDA.n140 0.15675
R411 VDDA.n140 VDDA.n126 0.15675
R412 VDDA.n135 VDDA.n126 0.15675
R413 VDDA.n135 VDDA.n134 0.15675
R414 VDDA.n134 VDDA.n133 0.15675
R415 VDDA VDDA.n0 0.1255
R416 VDDA VDDA.n21 0.1255
R417 VDDA.n171 VDDA 0.1255
R418 VDDA VDDA.n41 0.1255
R419 VDDA VDDA.n238 0.03175
R420 VDDA.n192 VDDA 0.03175
R421 VDDA VDDA.n170 0.03175
R422 VDDA.n149 VDDA 0.03175
R423 div2_4_1.C.n0 div2_4_1.C.t3 750.201
R424 div2_4_1.C.n1 div2_4_1.C.t4 349.433
R425 div2_4_1.C.n0 div2_4_1.C.t1 276.733
R426 div2_4_1.C.n2 div2_4_1.C.n1 206.333
R427 div2_4_1.C.n1 div2_4_1.C.n0 48.0005
R428 div2_4_1.C.n2 div2_4_1.C.t2 48.0005
R429 div2_4_1.C.t0 div2_4_1.C.n2 48.0005
R430 div5_2_0.B.n0 div5_2_0.B.t0 663.801
R431 div5_2_0.B.n0 div5_2_0.B.t2 348.851
R432 div5_2_0.B div5_2_0.B.t1 282.921
R433 div5_2_0.B div5_2_0.B.n0 114.133
R434 div5_2_0.D.n0 div5_2_0.D.t2 761.4
R435 div5_2_0.D.n1 div5_2_0.D.t4 350.349
R436 div5_2_0.D.n0 div5_2_0.D.t3 254.333
R437 div5_2_0.D.n2 div5_2_0.D.n1 206.333
R438 div5_2_0.D.n1 div5_2_0.D.n0 70.4005
R439 div5_2_0.D.n2 div5_2_0.D.t1 48.0005
R440 div5_2_0.D.t0 div5_2_0.D.n2 48.0005
R441 div5_2_0.Q2_b.n4 div5_2_0.Q2_b.t1 777.4
R442 div5_2_0.Q2_b.t11 div5_2_0.Q2_b.t8 514.134
R443 div5_2_0.Q2_b.n3 div5_2_0.Q2_b.n2 364.178
R444 div5_2_0.Q2_b.n0 div5_2_0.Q2_b.t7 353.467
R445 div5_2_0.Q2_b.t3 div5_2_0.Q2_b.n5 353.467
R446 div5_2_0.Q2_b.n6 div5_2_0.Q2_b.t3 318.702
R447 div5_2_0.Q2_b.n6 div5_2_0.Q2_b.t11 307.909
R448 div5_2_0.Q2_b.n5 div5_2_0.Q2_b.t4 289.2
R449 div5_2_0.Q2_b.n4 div5_2_0.Q2_b.n3 257.079
R450 div5_2_0.Q2_b.t0 div5_2_0.Q2_b.n7 233
R451 div5_2_0.Q2_b.n0 div5_2_0.Q2_b.t2 192.8
R452 div5_2_0.Q2_b.n2 div5_2_0.Q2_b.n1 176.733
R453 div5_2_0.Q2_b.n2 div5_2_0.Q2_b.t6 112.468
R454 div5_2_0.Q2_b.n1 div5_2_0.Q2_b.t9 112.468
R455 div5_2_0.Q2_b.n3 div5_2_0.Q2_b.t5 112.468
R456 div5_2_0.Q2_b.n5 div5_2_0.Q2_b.t10 112.468
R457 div5_2_0.Q2_b.n1 div5_2_0.Q2_b.n0 96.4005
R458 div5_2_0.Q2_b.n7 div5_2_0.Q2_b.n6 38.2642
R459 div5_2_0.Q2_b.n7 div5_2_0.Q2_b.n4 21.3338
R460 div5_2_0.M.n0 div5_2_0.M.t3 761.4
R461 div5_2_0.M.n1 div5_2_0.M.t4 349.433
R462 div5_2_0.M.n0 div5_2_0.M.t1 254.333
R463 div5_2_0.M.n2 div5_2_0.M.n1 206.333
R464 div5_2_0.M.n1 div5_2_0.M.n0 70.4005
R465 div5_2_0.M.t0 div5_2_0.M.n2 48.0005
R466 div5_2_0.M.n2 div5_2_0.M.t2 48.0005
R467 GNDA.t20 GNDA.t40 3168
R468 GNDA.t83 GNDA.t0 3080
R469 GNDA.t68 GNDA.t32 2992
R470 GNDA.t75 GNDA.t49 2904
R471 GNDA.t16 GNDA.t44 2904
R472 GNDA.t51 GNDA.t89 2904
R473 GNDA.t13 GNDA.t9 2904
R474 GNDA.t60 GNDA.t91 2904
R475 GNDA.t22 GNDA.t74 2904
R476 GNDA.t40 GNDA.n128 2772
R477 GNDA.t39 GNDA.t37 2200
R478 GNDA.t99 GNDA.t87 2200
R479 GNDA.t64 GNDA.t20 2200
R480 GNDA.n130 GNDA.t70 1980
R481 GNDA.n131 GNDA.t45 1980
R482 GNDA.n132 GNDA.t5 1980
R483 GNDA.n129 GNDA.t102 1716
R484 GNDA.t66 GNDA.n130 1716
R485 GNDA.t77 GNDA.n131 1716
R486 GNDA.n132 GNDA.t81 1716
R487 GNDA.n131 GNDA.n35 1204.13
R488 GNDA.n130 GNDA.n24 1204.13
R489 GNDA.n133 GNDA.n132 1204.13
R490 GNDA.n128 GNDA.t24 1188
R491 GNDA.t3 GNDA.n129 1188
R492 GNDA.n129 GNDA.n11 1182.8
R493 GNDA.n128 GNDA.n127 1182.8
R494 GNDA.t42 GNDA.t79 968
R495 GNDA.t35 GNDA.t42 968
R496 GNDA.t37 GNDA.t35 968
R497 GNDA.t32 GNDA.t39 968
R498 GNDA.t97 GNDA.t68 968
R499 GNDA.t85 GNDA.t97 968
R500 GNDA.t49 GNDA.t85 968
R501 GNDA.t26 GNDA.t75 968
R502 GNDA.t34 GNDA.t26 968
R503 GNDA.t0 GNDA.t34 968
R504 GNDA.t52 GNDA.t83 968
R505 GNDA.t47 GNDA.t52 968
R506 GNDA.t87 GNDA.t47 968
R507 GNDA.t24 GNDA.t99 968
R508 GNDA.t62 GNDA.t64 968
R509 GNDA.t95 GNDA.t62 968
R510 GNDA.t102 GNDA.t95 968
R511 GNDA.t61 GNDA.t3 968
R512 GNDA.t44 GNDA.t61 968
R513 GNDA.t56 GNDA.t16 968
R514 GNDA.t93 GNDA.t56 968
R515 GNDA.t89 GNDA.t93 968
R516 GNDA.t100 GNDA.t51 968
R517 GNDA.t70 GNDA.t100 968
R518 GNDA.t11 GNDA.t66 968
R519 GNDA.t72 GNDA.t11 968
R520 GNDA.t9 GNDA.t72 968
R521 GNDA.t28 GNDA.t13 968
R522 GNDA.t45 GNDA.t28 968
R523 GNDA.t18 GNDA.t77 968
R524 GNDA.t1 GNDA.t18 968
R525 GNDA.t91 GNDA.t1 968
R526 GNDA.t54 GNDA.t60 968
R527 GNDA.t5 GNDA.t54 968
R528 GNDA.t81 GNDA.t30 968
R529 GNDA.t30 GNDA.t14 968
R530 GNDA.t14 GNDA.t22 968
R531 GNDA.t74 GNDA.t58 968
R532 GNDA.t58 GNDA.t7 968
R533 GNDA.n74 GNDA.t33 295.933
R534 GNDA.n2 GNDA.t41 295.933
R535 GNDA.n3 GNDA.t21 295.933
R536 GNDA.n69 GNDA.n68 256.207
R537 GNDA.n67 GNDA.n66 247.934
R538 GNDA.n61 GNDA.n60 247.934
R539 GNDA.n86 GNDA.n59 247.934
R540 GNDA.n93 GNDA.n56 247.934
R541 GNDA.n105 GNDA.n51 247.934
R542 GNDA.n108 GNDA.n107 247.934
R543 GNDA.n6 GNDA.n5 247.934
R544 GNDA.n238 GNDA.n8 247.934
R545 GNDA.n17 GNDA.n16 247.934
R546 GNDA.n218 GNDA.n18 247.934
R547 GNDA.n23 GNDA.n22 246.714
R548 GNDA.n11 GNDA.t4 233
R549 GNDA.n127 GNDA.t25 233
R550 GNDA.n27 GNDA.n26 219.133
R551 GNDA.n196 GNDA.n29 219.133
R552 GNDA.n33 GNDA.n32 219.133
R553 GNDA.n38 GNDA.n37 219.133
R554 GNDA.n174 GNDA.n40 219.133
R555 GNDA.n44 GNDA.n43 219.133
R556 GNDA.n136 GNDA.n135 219.133
R557 GNDA.n152 GNDA.n138 219.133
R558 GNDA.n142 GNDA.n141 219.133
R559 GNDA.n232 GNDA.n11 54.4005
R560 GNDA.n127 GNDA.n126 54.4005
R561 GNDA.n68 GNDA.t80 48.0005
R562 GNDA.n68 GNDA.t43 48.0005
R563 GNDA.n66 GNDA.t36 48.0005
R564 GNDA.n66 GNDA.t38 48.0005
R565 GNDA.n60 GNDA.t69 48.0005
R566 GNDA.n60 GNDA.t98 48.0005
R567 GNDA.n59 GNDA.t86 48.0005
R568 GNDA.n59 GNDA.t50 48.0005
R569 GNDA.n56 GNDA.t76 48.0005
R570 GNDA.n56 GNDA.t27 48.0005
R571 GNDA.n51 GNDA.t84 48.0005
R572 GNDA.n51 GNDA.t53 48.0005
R573 GNDA.n107 GNDA.t48 48.0005
R574 GNDA.n107 GNDA.t88 48.0005
R575 GNDA.n5 GNDA.t65 48.0005
R576 GNDA.n5 GNDA.t63 48.0005
R577 GNDA.n8 GNDA.t96 48.0005
R578 GNDA.n8 GNDA.t103 48.0005
R579 GNDA.n16 GNDA.t17 48.0005
R580 GNDA.n16 GNDA.t57 48.0005
R581 GNDA.n18 GNDA.t94 48.0005
R582 GNDA.n18 GNDA.t90 48.0005
R583 GNDA.n22 GNDA.t101 48.0005
R584 GNDA.n22 GNDA.t71 48.0005
R585 GNDA.n26 GNDA.t67 48.0005
R586 GNDA.n26 GNDA.t12 48.0005
R587 GNDA.n29 GNDA.t73 48.0005
R588 GNDA.n29 GNDA.t10 48.0005
R589 GNDA.n32 GNDA.t29 48.0005
R590 GNDA.n32 GNDA.t46 48.0005
R591 GNDA.n37 GNDA.t78 48.0005
R592 GNDA.n37 GNDA.t19 48.0005
R593 GNDA.n40 GNDA.t2 48.0005
R594 GNDA.n40 GNDA.t92 48.0005
R595 GNDA.n43 GNDA.t55 48.0005
R596 GNDA.n43 GNDA.t6 48.0005
R597 GNDA.n135 GNDA.t82 48.0005
R598 GNDA.n135 GNDA.t31 48.0005
R599 GNDA.n138 GNDA.t15 48.0005
R600 GNDA.n138 GNDA.t23 48.0005
R601 GNDA.n141 GNDA.t59 48.0005
R602 GNDA.n141 GNDA.t8 48.0005
R603 GNDA.n72 GNDA.n65 32.0005
R604 GNDA.n73 GNDA.n72 32.0005
R605 GNDA.n75 GNDA.n73 32.0005
R606 GNDA.n79 GNDA.n63 32.0005
R607 GNDA.n80 GNDA.n79 32.0005
R608 GNDA.n81 GNDA.n80 32.0005
R609 GNDA.n85 GNDA.n84 32.0005
R610 GNDA.n87 GNDA.n57 32.0005
R611 GNDA.n91 GNDA.n57 32.0005
R612 GNDA.n92 GNDA.n91 32.0005
R613 GNDA.n94 GNDA.n54 32.0005
R614 GNDA.n98 GNDA.n54 32.0005
R615 GNDA.n99 GNDA.n98 32.0005
R616 GNDA.n100 GNDA.n99 32.0005
R617 GNDA.n100 GNDA.n52 32.0005
R618 GNDA.n104 GNDA.n52 32.0005
R619 GNDA.n109 GNDA.n106 32.0005
R620 GNDA.n113 GNDA.n49 32.0005
R621 GNDA.n114 GNDA.n113 32.0005
R622 GNDA.n115 GNDA.n114 32.0005
R623 GNDA.n115 GNDA.n46 32.0005
R624 GNDA.n125 GNDA.n47 32.0005
R625 GNDA.n121 GNDA.n47 32.0005
R626 GNDA.n121 GNDA.n120 32.0005
R627 GNDA.n120 GNDA.n119 32.0005
R628 GNDA.n250 GNDA.n249 32.0005
R629 GNDA.n249 GNDA.n248 32.0005
R630 GNDA.n245 GNDA.n244 32.0005
R631 GNDA.n244 GNDA.n243 32.0005
R632 GNDA.n240 GNDA.n239 32.0005
R633 GNDA.n237 GNDA.n9 32.0005
R634 GNDA.n233 GNDA.n9 32.0005
R635 GNDA.n231 GNDA.n230 32.0005
R636 GNDA.n230 GNDA.n12 32.0005
R637 GNDA.n226 GNDA.n12 32.0005
R638 GNDA.n226 GNDA.n225 32.0005
R639 GNDA.n225 GNDA.n224 32.0005
R640 GNDA.n224 GNDA.n14 32.0005
R641 GNDA.n220 GNDA.n219 32.0005
R642 GNDA.n217 GNDA.n19 32.0005
R643 GNDA.n213 GNDA.n19 32.0005
R644 GNDA.n213 GNDA.n212 32.0005
R645 GNDA.n212 GNDA.n211 32.0005
R646 GNDA.n211 GNDA.n21 32.0005
R647 GNDA.n207 GNDA.n206 32.0005
R648 GNDA.n203 GNDA.n202 32.0005
R649 GNDA.n202 GNDA.n201 32.0005
R650 GNDA.n198 GNDA.n197 32.0005
R651 GNDA.n195 GNDA.n30 32.0005
R652 GNDA.n191 GNDA.n30 32.0005
R653 GNDA.n191 GNDA.n190 32.0005
R654 GNDA.n190 GNDA.n189 32.0005
R655 GNDA.n186 GNDA.n185 32.0005
R656 GNDA.n185 GNDA.n184 32.0005
R657 GNDA.n181 GNDA.n180 32.0005
R658 GNDA.n180 GNDA.n179 32.0005
R659 GNDA.n176 GNDA.n175 32.0005
R660 GNDA.n173 GNDA.n41 32.0005
R661 GNDA.n169 GNDA.n41 32.0005
R662 GNDA.n169 GNDA.n168 32.0005
R663 GNDA.n168 GNDA.n167 32.0005
R664 GNDA.n164 GNDA.n163 32.0005
R665 GNDA.n163 GNDA.n162 32.0005
R666 GNDA.n159 GNDA.n158 32.0005
R667 GNDA.n158 GNDA.n157 32.0005
R668 GNDA.n154 GNDA.n153 32.0005
R669 GNDA.n151 GNDA.n139 32.0005
R670 GNDA.n147 GNDA.n139 32.0005
R671 GNDA.n147 GNDA.n146 32.0005
R672 GNDA.n146 GNDA.n145 32.0005
R673 GNDA.n67 GNDA.n65 28.8005
R674 GNDA.n250 GNDA.n2 28.8005
R675 GNDA.n240 GNDA.n6 28.8005
R676 GNDA.n207 GNDA.n23 28.8005
R677 GNDA.n189 GNDA.n33 28.8005
R678 GNDA.n167 GNDA.n44 28.8005
R679 GNDA.n145 GNDA.n142 28.8005
R680 GNDA.n75 GNDA.n74 25.6005
R681 GNDA.n84 GNDA.n61 25.6005
R682 GNDA.n93 GNDA.n92 25.6005
R683 GNDA.n109 GNDA.n108 25.6005
R684 GNDA.n220 GNDA.n17 25.6005
R685 GNDA.n198 GNDA.n27 25.6005
R686 GNDA.n176 GNDA.n38 25.6005
R687 GNDA.n154 GNDA.n136 25.6005
R688 GNDA.n238 GNDA.n237 22.4005
R689 GNDA.n206 GNDA.n24 22.4005
R690 GNDA.n184 GNDA.n35 22.4005
R691 GNDA.n162 GNDA.n133 22.4005
R692 GNDA.n87 GNDA.n86 19.2005
R693 GNDA.n105 GNDA.n104 19.2005
R694 GNDA.n248 GNDA.n3 19.2005
R695 GNDA.n233 GNDA.n232 19.2005
R696 GNDA.n218 GNDA.n217 19.2005
R697 GNDA.n196 GNDA.n195 19.2005
R698 GNDA.n174 GNDA.n173 19.2005
R699 GNDA.n152 GNDA.n151 19.2005
R700 GNDA.n126 GNDA.n46 16.0005
R701 GNDA.n126 GNDA.n125 16.0005
R702 GNDA.n86 GNDA.n85 12.8005
R703 GNDA.n106 GNDA.n105 12.8005
R704 GNDA.n245 GNDA.n3 12.8005
R705 GNDA.n232 GNDA.n231 12.8005
R706 GNDA.n219 GNDA.n218 12.8005
R707 GNDA.n197 GNDA.n196 12.8005
R708 GNDA.n175 GNDA.n174 12.8005
R709 GNDA.n153 GNDA.n152 12.8005
R710 GNDA.n143 GNDA.n142 10.7683
R711 GNDA.n69 GNDA.n67 10.4505
R712 GNDA.n239 GNDA.n238 9.6005
R713 GNDA.n203 GNDA.n24 9.6005
R714 GNDA.n181 GNDA.n35 9.6005
R715 GNDA.n159 GNDA.n133 9.6005
R716 GNDA.n145 GNDA.n144 9.3005
R717 GNDA.n146 GNDA.n140 9.3005
R718 GNDA.n148 GNDA.n147 9.3005
R719 GNDA.n149 GNDA.n139 9.3005
R720 GNDA.n151 GNDA.n150 9.3005
R721 GNDA.n153 GNDA.n137 9.3005
R722 GNDA.n155 GNDA.n154 9.3005
R723 GNDA.n157 GNDA.n156 9.3005
R724 GNDA.n158 GNDA.n134 9.3005
R725 GNDA.n160 GNDA.n159 9.3005
R726 GNDA.n162 GNDA.n161 9.3005
R727 GNDA.n163 GNDA.n45 9.3005
R728 GNDA.n165 GNDA.n164 9.3005
R729 GNDA.n167 GNDA.n166 9.3005
R730 GNDA.n168 GNDA.n42 9.3005
R731 GNDA.n170 GNDA.n169 9.3005
R732 GNDA.n171 GNDA.n41 9.3005
R733 GNDA.n173 GNDA.n172 9.3005
R734 GNDA.n175 GNDA.n39 9.3005
R735 GNDA.n177 GNDA.n176 9.3005
R736 GNDA.n179 GNDA.n178 9.3005
R737 GNDA.n180 GNDA.n36 9.3005
R738 GNDA.n182 GNDA.n181 9.3005
R739 GNDA.n184 GNDA.n183 9.3005
R740 GNDA.n185 GNDA.n34 9.3005
R741 GNDA.n187 GNDA.n186 9.3005
R742 GNDA.n189 GNDA.n188 9.3005
R743 GNDA.n190 GNDA.n31 9.3005
R744 GNDA.n192 GNDA.n191 9.3005
R745 GNDA.n193 GNDA.n30 9.3005
R746 GNDA.n195 GNDA.n194 9.3005
R747 GNDA.n197 GNDA.n28 9.3005
R748 GNDA.n199 GNDA.n198 9.3005
R749 GNDA.n201 GNDA.n200 9.3005
R750 GNDA.n202 GNDA.n25 9.3005
R751 GNDA.n204 GNDA.n203 9.3005
R752 GNDA.n206 GNDA.n205 9.3005
R753 GNDA.n208 GNDA.n207 9.3005
R754 GNDA.n70 GNDA.n65 9.3005
R755 GNDA.n72 GNDA.n71 9.3005
R756 GNDA.n73 GNDA.n64 9.3005
R757 GNDA.n76 GNDA.n75 9.3005
R758 GNDA.n77 GNDA.n63 9.3005
R759 GNDA.n79 GNDA.n78 9.3005
R760 GNDA.n80 GNDA.n62 9.3005
R761 GNDA.n82 GNDA.n81 9.3005
R762 GNDA.n84 GNDA.n83 9.3005
R763 GNDA.n85 GNDA.n58 9.3005
R764 GNDA.n88 GNDA.n87 9.3005
R765 GNDA.n89 GNDA.n57 9.3005
R766 GNDA.n91 GNDA.n90 9.3005
R767 GNDA.n92 GNDA.n55 9.3005
R768 GNDA.n95 GNDA.n94 9.3005
R769 GNDA.n96 GNDA.n54 9.3005
R770 GNDA.n98 GNDA.n97 9.3005
R771 GNDA.n99 GNDA.n53 9.3005
R772 GNDA.n101 GNDA.n100 9.3005
R773 GNDA.n102 GNDA.n52 9.3005
R774 GNDA.n104 GNDA.n103 9.3005
R775 GNDA.n106 GNDA.n50 9.3005
R776 GNDA.n110 GNDA.n109 9.3005
R777 GNDA.n111 GNDA.n49 9.3005
R778 GNDA.n113 GNDA.n112 9.3005
R779 GNDA.n114 GNDA.n48 9.3005
R780 GNDA.n116 GNDA.n115 9.3005
R781 GNDA.n117 GNDA.n46 9.3005
R782 GNDA.n125 GNDA.n124 9.3005
R783 GNDA.n123 GNDA.n47 9.3005
R784 GNDA.n122 GNDA.n121 9.3005
R785 GNDA.n120 GNDA.n118 9.3005
R786 GNDA.n119 GNDA.n0 9.3005
R787 GNDA.n251 GNDA.n250 9.3005
R788 GNDA.n249 GNDA.n1 9.3005
R789 GNDA.n248 GNDA.n247 9.3005
R790 GNDA.n246 GNDA.n245 9.3005
R791 GNDA.n244 GNDA.n4 9.3005
R792 GNDA.n243 GNDA.n242 9.3005
R793 GNDA.n241 GNDA.n240 9.3005
R794 GNDA.n239 GNDA.n7 9.3005
R795 GNDA.n237 GNDA.n236 9.3005
R796 GNDA.n235 GNDA.n9 9.3005
R797 GNDA.n234 GNDA.n233 9.3005
R798 GNDA.n231 GNDA.n10 9.3005
R799 GNDA.n230 GNDA.n229 9.3005
R800 GNDA.n228 GNDA.n12 9.3005
R801 GNDA.n227 GNDA.n226 9.3005
R802 GNDA.n225 GNDA.n13 9.3005
R803 GNDA.n224 GNDA.n223 9.3005
R804 GNDA.n222 GNDA.n14 9.3005
R805 GNDA.n221 GNDA.n220 9.3005
R806 GNDA.n219 GNDA.n15 9.3005
R807 GNDA.n217 GNDA.n216 9.3005
R808 GNDA.n215 GNDA.n19 9.3005
R809 GNDA.n214 GNDA.n213 9.3005
R810 GNDA.n212 GNDA.n20 9.3005
R811 GNDA.n211 GNDA.n210 9.3005
R812 GNDA.n209 GNDA.n21 9.3005
R813 GNDA.n74 GNDA.n63 6.4005
R814 GNDA.n81 GNDA.n61 6.4005
R815 GNDA.n94 GNDA.n93 6.4005
R816 GNDA.n108 GNDA.n49 6.4005
R817 GNDA.n17 GNDA.n14 6.4005
R818 GNDA.n201 GNDA.n27 6.4005
R819 GNDA.n179 GNDA.n38 6.4005
R820 GNDA.n157 GNDA.n136 6.4005
R821 GNDA.n119 GNDA.n2 3.2005
R822 GNDA.n243 GNDA.n6 3.2005
R823 GNDA.n23 GNDA.n21 3.2005
R824 GNDA.n186 GNDA.n33 3.2005
R825 GNDA.n164 GNDA.n44 3.2005
R826 GNDA.n70 GNDA.n69 0.442364
R827 GNDA.n143 GNDA 0.25314
R828 GNDA.n144 GNDA.n143 0.185879
R829 GNDA.n71 GNDA.n70 0.15675
R830 GNDA.n71 GNDA.n64 0.15675
R831 GNDA.n76 GNDA.n64 0.15675
R832 GNDA.n77 GNDA.n76 0.15675
R833 GNDA.n78 GNDA.n77 0.15675
R834 GNDA.n78 GNDA.n62 0.15675
R835 GNDA.n82 GNDA.n62 0.15675
R836 GNDA.n83 GNDA.n82 0.15675
R837 GNDA.n83 GNDA.n58 0.15675
R838 GNDA.n88 GNDA.n58 0.15675
R839 GNDA.n89 GNDA.n88 0.15675
R840 GNDA.n90 GNDA.n89 0.15675
R841 GNDA.n90 GNDA.n55 0.15675
R842 GNDA.n95 GNDA.n55 0.15675
R843 GNDA.n96 GNDA.n95 0.15675
R844 GNDA.n97 GNDA.n96 0.15675
R845 GNDA.n97 GNDA.n53 0.15675
R846 GNDA.n101 GNDA.n53 0.15675
R847 GNDA.n102 GNDA.n101 0.15675
R848 GNDA.n103 GNDA.n102 0.15675
R849 GNDA.n103 GNDA.n50 0.15675
R850 GNDA.n110 GNDA.n50 0.15675
R851 GNDA.n111 GNDA.n110 0.15675
R852 GNDA.n112 GNDA.n111 0.15675
R853 GNDA.n112 GNDA.n48 0.15675
R854 GNDA.n116 GNDA.n48 0.15675
R855 GNDA.n117 GNDA.n116 0.15675
R856 GNDA.n124 GNDA.n117 0.15675
R857 GNDA.n124 GNDA.n123 0.15675
R858 GNDA.n123 GNDA.n122 0.15675
R859 GNDA.n122 GNDA.n118 0.15675
R860 GNDA.n118 GNDA.n0 0.15675
R861 GNDA.n251 GNDA.n1 0.15675
R862 GNDA.n247 GNDA.n1 0.15675
R863 GNDA.n247 GNDA.n246 0.15675
R864 GNDA.n246 GNDA.n4 0.15675
R865 GNDA.n242 GNDA.n4 0.15675
R866 GNDA.n242 GNDA.n241 0.15675
R867 GNDA.n241 GNDA.n7 0.15675
R868 GNDA.n236 GNDA.n7 0.15675
R869 GNDA.n236 GNDA.n235 0.15675
R870 GNDA.n235 GNDA.n234 0.15675
R871 GNDA.n234 GNDA.n10 0.15675
R872 GNDA.n229 GNDA.n10 0.15675
R873 GNDA.n229 GNDA.n228 0.15675
R874 GNDA.n228 GNDA.n227 0.15675
R875 GNDA.n227 GNDA.n13 0.15675
R876 GNDA.n223 GNDA.n13 0.15675
R877 GNDA.n223 GNDA.n222 0.15675
R878 GNDA.n222 GNDA.n221 0.15675
R879 GNDA.n221 GNDA.n15 0.15675
R880 GNDA.n216 GNDA.n15 0.15675
R881 GNDA.n216 GNDA.n215 0.15675
R882 GNDA.n215 GNDA.n214 0.15675
R883 GNDA.n214 GNDA.n20 0.15675
R884 GNDA.n210 GNDA.n20 0.15675
R885 GNDA.n210 GNDA.n209 0.15675
R886 GNDA.n209 GNDA.n208 0.15675
R887 GNDA.n205 GNDA.n204 0.15675
R888 GNDA.n204 GNDA.n25 0.15675
R889 GNDA.n200 GNDA.n25 0.15675
R890 GNDA.n200 GNDA.n199 0.15675
R891 GNDA.n199 GNDA.n28 0.15675
R892 GNDA.n194 GNDA.n28 0.15675
R893 GNDA.n194 GNDA.n193 0.15675
R894 GNDA.n193 GNDA.n192 0.15675
R895 GNDA.n192 GNDA.n31 0.15675
R896 GNDA.n188 GNDA.n31 0.15675
R897 GNDA.n188 GNDA.n187 0.15675
R898 GNDA.n187 GNDA.n34 0.15675
R899 GNDA.n183 GNDA.n182 0.15675
R900 GNDA.n182 GNDA.n36 0.15675
R901 GNDA.n178 GNDA.n36 0.15675
R902 GNDA.n178 GNDA.n177 0.15675
R903 GNDA.n177 GNDA.n39 0.15675
R904 GNDA.n172 GNDA.n39 0.15675
R905 GNDA.n172 GNDA.n171 0.15675
R906 GNDA.n171 GNDA.n170 0.15675
R907 GNDA.n170 GNDA.n42 0.15675
R908 GNDA.n166 GNDA.n42 0.15675
R909 GNDA.n166 GNDA.n165 0.15675
R910 GNDA.n165 GNDA.n45 0.15675
R911 GNDA.n161 GNDA.n160 0.15675
R912 GNDA.n160 GNDA.n134 0.15675
R913 GNDA.n156 GNDA.n134 0.15675
R914 GNDA.n156 GNDA.n155 0.15675
R915 GNDA.n155 GNDA.n137 0.15675
R916 GNDA.n150 GNDA.n137 0.15675
R917 GNDA.n150 GNDA.n149 0.15675
R918 GNDA.n149 GNDA.n148 0.15675
R919 GNDA.n148 GNDA.n140 0.15675
R920 GNDA.n144 GNDA.n140 0.15675
R921 GNDA GNDA.n0 0.1255
R922 GNDA.n208 GNDA 0.1255
R923 GNDA GNDA.n34 0.1255
R924 GNDA GNDA.n45 0.1255
R925 GNDA GNDA.n251 0.03175
R926 GNDA.n205 GNDA 0.03175
R927 GNDA.n183 GNDA 0.03175
R928 GNDA.n161 GNDA 0.03175
R929 div8.t5 div8.t3 1012.2
R930 div8.n1 div8.t0 663.801
R931 div8.t4 div8.t2 401.668
R932 div8.n1 div8.t5 361.692
R933 div8.n2 div8.t1 298.921
R934 div8.n0 div8.t4 257.067
R935 div3_3_0.VIN div8.n0 216.9
R936 div8.n0 div8.t6 208.868
R937 div2_4_0.VOUT div3_3_0.VIN 177.701
R938 div8.n2 div8.n1 67.2005
R939 div2_4_0.VOUT div8.n2 36.8005
R940 div3_3_0.CLK.n3 div3_3_0.CLK.n2 742.51
R941 div3_3_0.CLK.n8 div3_3_0.CLK.t1 723.534
R942 div3_3_0.CLK.t2 div3_3_0.CLK.n9 723.534
R943 div3_3_0.CLK.n2 div3_3_0.CLK.n1 684.806
R944 div3_3_0.CLK.n7 div3_3_0.CLK.n6 366.856
R945 div3_3_0.CLK.n0 div3_3_0.CLK.t9 337.401
R946 div3_3_0.CLK.n0 div3_3_0.CLK.t7 305.267
R947 div3_3_0.CLK.n8 div3_3_0.CLK.t0 254.333
R948 div3_3_0.CLK.n4 div3_3_0.CLK.n3 224.934
R949 div3_3_0.CLK.n7 div3_3_0.CLK.t12 190.123
R950 div3_3_0.CLK.n9 div3_3_0.CLK.n7 187.201
R951 div3_3_0.CLK.n1 div3_3_0.CLK.n0 176.733
R952 div3_3_0.CLK.n5 div3_3_0.CLK.n4 176.733
R953 div3_3_0.CLK.n6 div3_3_0.CLK.n5 176.733
R954 div3_3_0.CLK.n3 div3_3_0.CLK.t6 144.601
R955 div3_3_0.CLK.n2 div3_3_0.CLK.t3 131.976
R956 div3_3_0.CLK.n0 div3_3_0.CLK.t11 128.534
R957 div3_3_0.CLK.n1 div3_3_0.CLK.t8 128.534
R958 div3_3_0.CLK.n4 div3_3_0.CLK.t4 112.468
R959 div3_3_0.CLK.n6 div3_3_0.CLK.t5 112.468
R960 div3_3_0.CLK.n5 div3_3_0.CLK.t10 112.468
R961 div3_3_0.CLK.n9 div3_3_0.CLK.n8 70.4005
R962 div24.n3 div24.n2 919.244
R963 div3_3_0.VOUT div24.n7 886.702
R964 div24.t9 div24.t3 819.4
R965 div24.n9 div24.n8 628.734
R966 div24.n2 div24.n1 520.361
R967 div24.n7 div24.n6 364.178
R968 div24.n0 div24.t7 337.401
R969 div24.n10 div24.t9 336.25
R970 div24.n0 div24.t11 305.267
R971 div24.n9 div24.t0 257.534
R972 div24.n4 div24.t4 192.8
R973 div24.n1 div24.n0 176.733
R974 div24.n6 div24.n5 176.733
R975 div24.n4 div24.n3 160.667
R976 div24.n3 div24.t8 144.601
R977 div24.n2 div24.t14 131.976
R978 div24.n0 div24.t12 128.534
R979 div24.n1 div24.t6 128.534
R980 div24.n6 div24.t5 112.468
R981 div24.n5 div24.t13 112.468
R982 div24.n7 div24.t10 112.468
R983 div24.n5 div24.n4 96.4005
R984 div24.n8 div24.t1 78.8005
R985 div24.n8 div24.t2 78.8005
R986 div5_2_0.VIN div24.n10 25.6005
R987 div24.n10 div24.n9 11.2005
R988 div5_2_0.VIN div3_3_0.VOUT 6.4005
R989 div3_3_0.A.n0 div3_3_0.A.t0 713.933
R990 div3_3_0.A.n0 div3_3_0.A.t2 314.233
R991 div3_3_0.A.t1 div3_3_0.A.n0 308.2
R992 div2.t5 div2.t3 1012.2
R993 div2.n1 div2.t0 663.801
R994 div2.t6 div2.t4 401.668
R995 div2.n1 div2.t5 361.692
R996 div2.n0 div2.t2 353.467
R997 div2.n2 div2.t1 298.921
R998 div2.n0 div2.t6 257.067
R999 div2_4_2.VIN div2.n0 216.9
R1000 div2_4_1.VOUT div2_4_2.VIN 177.701
R1001 div2.n2 div2.n1 67.2005
R1002 div2_4_1.VOUT div2.n2 36.8005
R1003 a_1320_n1010.n4 a_1320_n1010.t1 752.333
R1004 a_1320_n1010.t2 a_1320_n1010.n5 752.333
R1005 a_1320_n1010.n0 a_1320_n1010.t7 514.134
R1006 a_1320_n1010.n3 a_1320_n1010.n2 366.856
R1007 a_1320_n1010.n4 a_1320_n1010.t0 254.333
R1008 a_1320_n1010.n3 a_1320_n1010.t3 190.123
R1009 a_1320_n1010.n5 a_1320_n1010.n3 187.201
R1010 a_1320_n1010.n1 a_1320_n1010.n0 176.733
R1011 a_1320_n1010.n2 a_1320_n1010.n1 176.733
R1012 a_1320_n1010.n0 a_1320_n1010.t5 112.468
R1013 a_1320_n1010.n2 a_1320_n1010.t4 112.468
R1014 a_1320_n1010.n1 a_1320_n1010.t6 112.468
R1015 a_1320_n1010.n5 a_1320_n1010.n4 70.4005
R1016 div3_3_0.I.n0 div3_3_0.I.t1 663.801
R1017 div3_3_0.I.t4 div3_3_0.I.t2 514.134
R1018 div3_3_0.I.n0 div3_3_0.I.t4 479.284
R1019 div3_3_0.I.n3 div3_3_0.I.n2 344.8
R1020 div3_3_0.I.n1 div3_3_0.I.t6 289.2
R1021 div3_3_0.I.t0 div3_3_0.I.n3 275.454
R1022 div3_3_0.I.n2 div3_3_0.I.t5 241
R1023 div3_3_0.I.n1 div3_3_0.I.t3 112.468
R1024 div3_3_0.I.n3 div3_3_0.I.n0 97.9205
R1025 div3_3_0.I.n2 div3_3_0.I.n1 64.2672
R1026 div3_3_0.G.t0 div3_3_0.G.t1 96.0005
R1027 VIN.t0 VIN.t2 401.668
R1028 VIN.n0 VIN.t1 353.467
R1029 VIN.n0 VIN.t0 257.067
R1030 VIN VIN.n0 216.9
R1031 a_20_n1010.n4 a_20_n1010.t1 752.333
R1032 a_20_n1010.t2 a_20_n1010.n5 752.333
R1033 a_20_n1010.n0 a_20_n1010.t7 514.134
R1034 a_20_n1010.n3 a_20_n1010.n2 366.856
R1035 a_20_n1010.n5 a_20_n1010.t0 254.333
R1036 a_20_n1010.n3 a_20_n1010.t5 190.123
R1037 a_20_n1010.n4 a_20_n1010.n3 187.201
R1038 a_20_n1010.n1 a_20_n1010.n0 176.733
R1039 a_20_n1010.n2 a_20_n1010.n1 176.733
R1040 a_20_n1010.n0 a_20_n1010.t3 112.468
R1041 a_20_n1010.n2 a_20_n1010.t6 112.468
R1042 a_20_n1010.n1 a_20_n1010.t4 112.468
R1043 a_20_n1010.n5 a_20_n1010.n4 70.4005
R1044 div4.t3 div4.t5 1012.2
R1045 div4.n1 div4.t1 663.801
R1046 div4.t2 div4.t4 401.668
R1047 div4.n1 div4.t3 361.692
R1048 div4.n0 div4.t6 353.467
R1049 div4.n2 div4.t0 298.921
R1050 div4.n0 div4.t2 257.067
R1051 div2_4_0.VIN div4.n0 216.9
R1052 div2_4_2.VOUT div2_4_0.VIN 177.701
R1053 div4.n2 div4.n1 67.2005
R1054 div2_4_2.VOUT div4.n2 36.8005
R1055 a_2620_n1010.n4 a_2620_n1010.t1 752.333
R1056 a_2620_n1010.t2 a_2620_n1010.n5 752.333
R1057 a_2620_n1010.n0 a_2620_n1010.t4 514.134
R1058 a_2620_n1010.n3 a_2620_n1010.n2 366.856
R1059 a_2620_n1010.n5 a_2620_n1010.t0 254.333
R1060 a_2620_n1010.n3 a_2620_n1010.t3 190.123
R1061 a_2620_n1010.n4 a_2620_n1010.n3 187.201
R1062 a_2620_n1010.n1 a_2620_n1010.n0 176.733
R1063 a_2620_n1010.n2 a_2620_n1010.n1 176.733
R1064 a_2620_n1010.n0 a_2620_n1010.t5 112.468
R1065 a_2620_n1010.n2 a_2620_n1010.t7 112.468
R1066 a_2620_n1010.n1 a_2620_n1010.t6 112.468
R1067 a_2620_n1010.n5 a_2620_n1010.n4 70.4005
R1068 div2_4_1.B.t0 div2_4_1.B.t1 96.0005
R1069 div2_4_0.B.t0 div2_4_0.B.t1 96.0005
R1070 div2_4_0.A.n0 div2_4_0.A.t1 713.933
R1071 div2_4_0.A.t0 div2_4_0.A.n0 337
R1072 div2_4_0.A.n0 div2_4_0.A.t2 314.233
R1073 div3_3_0.E.n0 div3_3_0.E.t1 685.134
R1074 div3_3_0.E.n1 div3_3_0.E.t0 663.801
R1075 div3_3_0.E.n0 div3_3_0.E.t3 534.268
R1076 div3_3_0.E.t2 div3_3_0.E.n1 362.921
R1077 div3_3_0.E.n1 div3_3_0.E.n0 91.7338
R1078 div3_3_0.F.t0 div3_3_0.F.t1 96.0005
R1079 div3_3_0.H.n0 div3_3_0.H.t0 723.534
R1080 div3_3_0.H.n1 div3_3_0.H.t4 553.534
R1081 div3_3_0.H.n0 div3_3_0.H.t2 254.333
R1082 div3_3_0.H.n2 div3_3_0.H.n1 206.333
R1083 div3_3_0.H.n1 div3_3_0.H.n0 70.4005
R1084 div3_3_0.H.t3 div3_3_0.H.n2 48.0005
R1085 div3_3_0.H.n2 div3_3_0.H.t1 48.0005
R1086 div5_2_0.A.n2 div5_2_0.A.t1 755.534
R1087 div5_2_0.A.t2 div5_2_0.A.n2 685.134
R1088 div5_2_0.A.n1 div5_2_0.A.n0 389.733
R1089 div5_2_0.A.n1 div5_2_0.A.t0 340.2
R1090 div5_2_0.A.n0 div5_2_0.A.t4 321.334
R1091 div5_2_0.A.n0 div5_2_0.A.t3 144.601
R1092 div5_2_0.A.n2 div5_2_0.A.n1 19.2005
R1093 div3_3_0.D.n1 div3_3_0.D.n0 701.467
R1094 div3_3_0.D.n1 div3_3_0.D.t1 694.201
R1095 div3_3_0.D.n0 div3_3_0.D.t3 321.334
R1096 div3_3_0.D.t0 div3_3_0.D.n1 314.921
R1097 div3_3_0.D.n0 div3_3_0.D.t2 144.601
R1098 div3_3_0.C.n0 div3_3_0.C.t0 721.4
R1099 div3_3_0.C.n1 div3_3_0.C.t4 350.349
R1100 div3_3_0.C.n0 div3_3_0.C.t2 276.733
R1101 div3_3_0.C.n2 div3_3_0.C.n1 206.333
R1102 div3_3_0.C.n1 div3_3_0.C.n0 48.0005
R1103 div3_3_0.C.t3 div3_3_0.C.n2 48.0005
R1104 div3_3_0.C.n2 div3_3_0.C.t1 48.0005
R1105 div5_2_0.J.n2 div5_2_0.J.t0 723.534
R1106 div5_2_0.J.n1 div5_2_0.J.t4 553.534
R1107 div5_2_0.J.t3 div5_2_0.J.n2 254.333
R1108 div5_2_0.J.n1 div5_2_0.J.n0 206.333
R1109 div5_2_0.J.n2 div5_2_0.J.n1 70.4005
R1110 div5_2_0.J.n0 div5_2_0.J.t2 48.0005
R1111 div5_2_0.J.n0 div5_2_0.J.t1 48.0005
R1112 div5_2_0.L.t0 div5_2_0.L.t1 96.0005
R1113 div5_2_0.K.n0 div5_2_0.K.t1 663.801
R1114 div5_2_0.K.t0 div5_2_0.K.n0 397.053
R1115 div5_2_0.K.n0 div5_2_0.K.t2 355.378
R1116 div2_4_2.C.n2 div2_4_2.C.t0 750.201
R1117 div2_4_2.C.n1 div2_4_2.C.t4 349.433
R1118 div2_4_2.C.t3 div2_4_2.C.n2 276.733
R1119 div2_4_2.C.n1 div2_4_2.C.n0 206.333
R1120 div2_4_2.C.n0 div2_4_2.C.t2 48.0005
R1121 div2_4_2.C.n0 div2_4_2.C.t1 48.0005
R1122 div2_4_2.C.n2 div2_4_2.C.n1 48.0005
R1123 div2_4_0.C.n0 div2_4_0.C.t3 750.201
R1124 div2_4_0.C.n1 div2_4_0.C.t4 349.433
R1125 div2_4_0.C.n0 div2_4_0.C.t0 276.733
R1126 div2_4_0.C.n2 div2_4_0.C.n1 206.333
R1127 div2_4_0.C.n1 div2_4_0.C.n0 48.0005
R1128 div2_4_0.C.t2 div2_4_0.C.n2 48.0005
R1129 div2_4_0.C.n2 div2_4_0.C.t1 48.0005
R1130 VOUT.n1 VOUT.t3 772.196
R1131 VOUT.n3 VOUT.t0 751.801
R1132 VOUT.n2 VOUT.n1 607.465
R1133 VOUT.t3 VOUT.t5 514.134
R1134 VOUT.n0 VOUT.t4 289.2
R1135 VOUT.n2 VOUT.t1 233
R1136 VOUT.n1 VOUT.n0 208.868
R1137 VOUT.n0 VOUT.t2 176.733
R1138 VOUT.n3 VOUT.n2 40.3205
R1139 VOUT VOUT.n3 32.0005
R1140 div2_4_2.A.n0 div2_4_2.A.t0 713.933
R1141 div2_4_2.A.t1 div2_4_2.A.n0 337
R1142 div2_4_2.A.n0 div2_4_2.A.t2 314.233
R1143 div2_4_2.B.t0 div2_4_2.B.t1 96.0005
R1144 div5_2_0.E.n0 div5_2_0.E.t1 723
R1145 div5_2_0.E.t3 div5_2_0.E.t2 514.134
R1146 div5_2_0.E.n0 div5_2_0.E.t3 335.983
R1147 div5_2_0.E.t0 div5_2_0.E.n0 314.921
R1148 div5_2_0.I.t0 div5_2_0.I.n0 531.067
R1149 div5_2_0.I.n0 div5_2_0.I.t2 48.0005
R1150 div5_2_0.I.n0 div5_2_0.I.t1 48.0005
R1151 div5_2_0.F.t0 div5_2_0.F.t1 157.601
R1152 div5_2_0.G.n0 div5_2_0.G.t0 685.134
R1153 div5_2_0.G.n1 div5_2_0.G.t1 685.134
R1154 div5_2_0.G.n0 div5_2_0.G.t3 534.268
R1155 div5_2_0.G.t2 div5_2_0.G.n1 340.521
R1156 div5_2_0.G.n1 div5_2_0.G.n0 105.6
R1157 div3_3_0.B.t0 div3_3_0.B.t1 96.0005
R1158 div5_2_0.C.t0 div5_2_0.C.t1 96.0005
R1159 div5_2_0.H.t0 div5_2_0.H.t1 96.0005
C0 VDDA VOUT 1.02478f
C1 VDDA VIN 0.138342f
C2 div5_2_0.B VDDA 0.506749f
C3 VOUT GNDA 1.84912f
C4 VIN GNDA 0.344458f
C5 VDDA GNDA 12.908f
C6 div5_2_0.B GNDA 0.178977f
.ends

