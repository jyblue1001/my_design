magic
tech sky130A
timestamp 1752572815
<< metal1 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6655 2990 6685
rect 2950 6650 2990 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6040 6685 6080 6690
rect 6040 6655 6045 6685
rect 6075 6655 6080 6685
rect 3030 6650 3070 6655
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6550 2945 6580
rect 2905 6545 2945 6550
rect 2915 3090 2935 6545
rect 2960 3140 2980 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 3955 6645 3995 6650
rect 3955 6615 3960 6645
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3965 5280 3985 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 4000 6475 4040 6480
rect 4000 6445 4005 6475
rect 4035 6445 4040 6475
rect 4000 6440 4040 6445
rect 4010 5405 4030 6440
rect 4000 5400 4040 5405
rect 4000 5370 4005 5400
rect 4035 5370 4040 5400
rect 4000 5365 4040 5370
rect 4075 5400 4115 5405
rect 4075 5370 4080 5400
rect 4110 5370 4115 5400
rect 4075 5365 4115 5370
rect 3965 5275 4040 5280
rect 3965 5245 3985 5275
rect 4015 5245 4040 5275
rect 3965 5240 4040 5245
rect 4020 3635 4040 5240
rect 4010 3630 4050 3635
rect 4010 3600 4015 3630
rect 4045 3600 4050 3630
rect 4010 3595 4050 3600
rect 4085 3375 4105 5365
rect 5085 5340 5105 6655
rect 5730 6585 5750 6655
rect 6040 6650 6080 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5385 5420 5405 6485
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5385 5415 5415
rect 5375 5380 5415 5385
rect 5495 5415 5535 5420
rect 5495 5385 5500 5415
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 5075 5335 5115 5340
rect 5075 5305 5080 5335
rect 5110 5305 5115 5335
rect 5075 5300 5115 5305
rect 5505 4720 5525 5380
rect 5995 5335 6035 5340
rect 5995 5305 6000 5335
rect 6030 5305 6035 5335
rect 5995 5300 6035 5305
rect 5495 4715 5535 4720
rect 5495 4685 5500 4715
rect 5530 4685 5535 4715
rect 5495 4680 5535 4685
rect 6005 3530 6025 5300
rect 6050 3685 6070 6650
rect 6785 5090 6805 6660
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 7020 6650 7060 6655
rect 7100 6685 7140 6690
rect 7100 6655 7105 6685
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5055 6450 5085
rect 6410 5050 6450 5055
rect 6775 5085 6815 5090
rect 6775 5055 6780 5085
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 6420 4775 6440 5050
rect 6410 4770 6450 4775
rect 6410 4740 6415 4770
rect 6445 4740 6450 4770
rect 6410 4735 6450 4740
rect 6040 3680 6080 3685
rect 6040 3650 6045 3680
rect 6075 3650 6080 3680
rect 6040 3645 6080 3650
rect 5215 3525 5255 3530
rect 5215 3495 5220 3525
rect 5250 3495 5255 3525
rect 5215 3490 5255 3495
rect 5995 3525 6035 3530
rect 5995 3495 6000 3525
rect 6030 3495 6035 3525
rect 5995 3490 6035 3495
rect 4075 3370 4115 3375
rect 4075 3340 4080 3370
rect 4110 3340 4115 3370
rect 4075 3335 4115 3340
rect 2950 3135 3005 3140
rect 2950 3105 2955 3135
rect 2905 3085 2960 3090
rect 2905 3055 2910 3085
rect 2940 3055 2960 3085
rect 2905 3050 2960 3055
rect 2940 2865 2960 3050
rect 2985 2755 3005 3135
rect 5225 2590 5245 3490
rect 7110 3140 7130 6650
rect 7145 6580 7185 6585
rect 7145 6550 7150 6580
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 7085 3135 7140 3140
rect 7085 2755 7105 3135
rect 7135 3105 7140 3135
rect 7155 3090 7175 6545
rect 7130 3085 7185 3090
rect 7130 3055 7150 3085
rect 7180 3055 7185 3085
rect 7130 3050 7185 3055
rect 7130 2865 7150 3050
rect 5205 2585 5245 2590
rect 5205 2555 5210 2585
rect 5240 2555 5245 2585
rect 5205 2550 5245 2555
rect 2440 1800 2480 1830
<< via1 >>
rect 2955 6655 2985 6685
rect 3035 6655 3065 6685
rect 6045 6655 6075 6685
rect 2910 6550 2940 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 3960 6615 3990 6645
rect 3550 6445 3580 6475
rect 4335 6550 4365 6580
rect 4005 6445 4035 6475
rect 4005 5370 4035 5400
rect 4080 5370 4110 5400
rect 3985 5245 4015 5275
rect 4015 3600 4045 3630
rect 6705 6655 6735 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 5380 5385 5410 5415
rect 5500 5385 5530 5415
rect 5080 5305 5110 5335
rect 6000 5305 6030 5335
rect 5500 4685 5530 4715
rect 7025 6655 7055 6685
rect 7105 6655 7135 6685
rect 6415 5055 6445 5085
rect 6780 5055 6810 5085
rect 6415 4740 6445 4770
rect 6045 3650 6075 3680
rect 5220 3495 5250 3525
rect 6000 3495 6030 3525
rect 4080 3340 4110 3370
rect 2955 3105 2985 3135
rect 2910 3055 2940 3085
rect 7150 6550 7180 6580
rect 7105 3105 7135 3135
rect 7150 3055 7180 3085
rect 5210 2555 5240 2585
<< metal2 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6680 2990 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2985 6660 3035 6680
rect 2985 6655 2990 6660
rect 2950 6650 2990 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6040 6685 6080 6690
rect 6040 6655 6045 6685
rect 6075 6680 6080 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6075 6660 6705 6680
rect 6075 6655 6080 6660
rect 6040 6650 6080 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 6700 6650 6740 6655
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6680 7060 6685
rect 7100 6685 7140 6690
rect 7100 6680 7105 6685
rect 7055 6660 7105 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7100 6655 7105 6660
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 3955 6645 3995 6650
rect 3955 6640 3960 6645
rect 3435 6620 3960 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 3955 6615 3960 6620
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6575 2945 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2940 6555 4335 6575
rect 2940 6550 2945 6555
rect 2905 6545 2945 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7145 6580 7185 6585
rect 7145 6575 7150 6580
rect 5755 6555 7150 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7145 6550 7150 6555
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 4000 6475 4040 6480
rect 4000 6470 4005 6475
rect 3580 6450 4005 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 4000 6445 4005 6450
rect 4035 6445 4040 6475
rect 4000 6440 4040 6445
rect 5375 5415 5415 5420
rect 4000 5400 4040 5405
rect 4000 5370 4005 5400
rect 4035 5395 4040 5400
rect 4075 5400 4115 5405
rect 4075 5395 4080 5400
rect 4035 5375 4080 5395
rect 4035 5370 4040 5375
rect 4000 5365 4040 5370
rect 4075 5370 4080 5375
rect 4110 5370 4115 5400
rect 5375 5385 5380 5415
rect 5410 5410 5415 5415
rect 5495 5415 5535 5420
rect 5495 5410 5500 5415
rect 5410 5390 5500 5410
rect 5410 5385 5415 5390
rect 5375 5380 5415 5385
rect 5495 5385 5500 5390
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 4075 5365 4115 5370
rect 5075 5335 5115 5340
rect 5075 5305 5080 5335
rect 5110 5330 5115 5335
rect 5995 5335 6035 5340
rect 5995 5330 6000 5335
rect 5110 5310 6000 5330
rect 5110 5305 5115 5310
rect 5075 5300 5115 5305
rect 5995 5305 6000 5310
rect 6030 5305 6035 5335
rect 5995 5300 6035 5305
rect 3980 5275 4020 5280
rect 3980 5245 3985 5275
rect 4015 5245 4020 5275
rect 3980 5240 4020 5245
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5080 6450 5085
rect 6775 5085 6815 5090
rect 6775 5080 6780 5085
rect 6445 5060 6780 5080
rect 6445 5055 6450 5060
rect 6410 5050 6450 5055
rect 6775 5055 6780 5060
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 6410 4770 6450 4775
rect 6410 4765 6415 4770
rect 5745 4745 6415 4765
rect 6410 4740 6415 4745
rect 6445 4740 6450 4770
rect 6410 4735 6450 4740
rect 5495 4715 5535 4720
rect 5495 4685 5500 4715
rect 5530 4685 5535 4715
rect 5495 4680 5535 4685
rect 6040 3680 6080 3685
rect 6040 3675 6045 3680
rect 5270 3655 6045 3675
rect 6040 3650 6045 3655
rect 6075 3650 6080 3680
rect 6040 3645 6080 3650
rect 4010 3630 4050 3635
rect 4010 3600 4015 3630
rect 4045 3615 4050 3630
rect 4045 3600 4510 3615
rect 4010 3595 4510 3600
rect 5215 3525 5255 3530
rect 5215 3495 5220 3525
rect 5250 3520 5255 3525
rect 5995 3525 6035 3530
rect 5995 3520 6000 3525
rect 5250 3500 6000 3520
rect 5250 3495 5255 3500
rect 5215 3490 5255 3495
rect 5995 3495 6000 3500
rect 6030 3495 6035 3525
rect 5995 3490 6035 3495
rect 4075 3370 4115 3375
rect 4075 3340 4080 3370
rect 4110 3340 4115 3370
rect 4075 3335 4115 3340
rect 2950 3135 2990 3140
rect 2950 3105 2955 3135
rect 2985 3105 2990 3135
rect 7100 3135 7140 3140
rect 7100 3105 7105 3135
rect 7135 3105 7140 3135
rect 2905 3085 2945 3090
rect 2905 3055 2910 3085
rect 2940 3055 2945 3085
rect 2905 3050 2945 3055
rect 7145 3085 7185 3090
rect 7145 3055 7150 3085
rect 7180 3055 7185 3085
rect 7145 3050 7185 3055
rect 4080 2945 4100 2965
rect 5990 2945 6010 2965
rect 5205 2585 5245 2590
rect 5205 2580 5210 2585
rect 5035 2560 5210 2580
rect 5205 2555 5210 2560
rect 5240 2555 5245 2585
rect 5205 2550 5245 2555
rect 5035 2455 5055 2475
rect 2815 2140 2835 2160
rect 7220 2140 7240 2160
rect 2440 1800 2480 1830
<< metal3 >>
rect 9335 14460 9385 14465
rect 9335 14420 9340 14460
rect 9380 14420 9385 14460
rect 9335 14415 9385 14420
rect 9340 50 9380 14415
rect 9335 45 9385 50
rect 9335 5 9340 45
rect 9380 5 9385 45
rect 9335 0 9385 5
<< via3 >>
rect 9340 14420 9380 14460
rect 9340 5 9380 45
<< metal4 >>
rect 7255 14460 9385 14465
rect 7255 14420 9340 14460
rect 9380 14420 9385 14460
rect 7255 14415 9385 14420
rect 540 6700 590 6750
rect 540 0 590 50
rect 9325 45 9385 50
rect 9325 5 9340 45
rect 9380 5 9385 45
rect 9325 0 9385 5
use bgr_7  bgr_7_0
timestamp 1752484787
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic_14  two_stage_opamp_dummy_magic_14_0
timestamp 1752571794
transform 1 0 4200 0 1 2465
box -3850 -2465 5140 4285
<< labels >>
flabel metal4 565 0 565 0 5 FreeSans 800 0 0 -320 GNDA
port 2 s
flabel metal2 2825 2140 2825 2140 5 FreeSans 800 0 0 -320 VOUT+
port 3 s
flabel metal2 7230 2140 7230 2140 5 FreeSans 800 0 0 -320 VOUT-
port 4 s
flabel metal4 565 6750 565 6750 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 4080 2955 4080 2955 7 FreeSans 800 0 -320 0 VIN+
port 5 w
flabel metal2 6010 2955 6010 2955 3 FreeSans 800 0 320 0 VIN-
port 6 e
<< end >>
