magic
tech sky130A
timestamp 1737957840
<< nwell >>
rect 970 225 2110 730
<< nmos >>
rect 1040 20 1055 70
rect 1105 20 1120 70
rect 1170 20 1185 70
rect 1235 20 1250 70
rect 1400 20 1415 70
rect 1465 20 1480 70
rect 1530 20 1545 70
rect 1595 20 1610 70
rect 1780 20 1795 70
rect 1845 20 1860 70
rect 1910 20 1925 70
rect 1975 20 1990 70
rect 1605 -380 1655 -130
rect 1705 -380 1755 -130
rect 1805 -380 1855 -130
rect 1905 -380 1955 -130
<< pmos >>
rect 1060 460 1110 710
rect 1160 460 1210 710
rect 1260 460 1310 710
rect 1360 460 1410 710
rect 1460 460 1510 710
rect 1560 460 1610 710
rect 1660 460 1710 710
rect 1760 460 1810 710
rect 1040 245 1055 345
rect 1105 245 1120 345
rect 1170 245 1185 345
rect 1235 245 1250 345
rect 1400 245 1415 345
rect 1465 245 1480 345
rect 1530 245 1545 345
rect 1595 245 1610 345
rect 1780 245 1795 345
rect 1845 245 1860 345
rect 1910 245 1925 345
rect 1975 245 1990 345
<< ndiff >>
rect 990 55 1040 70
rect 990 35 1005 55
rect 1025 35 1040 55
rect 990 20 1040 35
rect 1055 55 1105 70
rect 1055 35 1070 55
rect 1090 35 1105 55
rect 1055 20 1105 35
rect 1120 55 1170 70
rect 1120 35 1135 55
rect 1155 35 1170 55
rect 1120 20 1170 35
rect 1185 55 1235 70
rect 1185 35 1200 55
rect 1220 35 1235 55
rect 1185 20 1235 35
rect 1250 55 1300 70
rect 1350 55 1400 70
rect 1250 35 1265 55
rect 1285 35 1300 55
rect 1350 35 1365 55
rect 1385 35 1400 55
rect 1250 20 1300 35
rect 1350 20 1400 35
rect 1415 55 1465 70
rect 1415 35 1430 55
rect 1450 35 1465 55
rect 1415 20 1465 35
rect 1480 55 1530 70
rect 1480 35 1495 55
rect 1515 35 1530 55
rect 1480 20 1530 35
rect 1545 55 1595 70
rect 1545 35 1560 55
rect 1580 35 1595 55
rect 1545 20 1595 35
rect 1610 55 1660 70
rect 1610 35 1625 55
rect 1645 35 1660 55
rect 1610 20 1660 35
rect 1730 55 1780 70
rect 1730 35 1745 55
rect 1765 35 1780 55
rect 1730 20 1780 35
rect 1795 55 1845 70
rect 1795 35 1810 55
rect 1830 35 1845 55
rect 1795 20 1845 35
rect 1860 55 1910 70
rect 1860 35 1875 55
rect 1895 35 1910 55
rect 1860 20 1910 35
rect 1925 55 1975 70
rect 1925 35 1940 55
rect 1960 35 1975 55
rect 1925 20 1975 35
rect 1990 55 2040 70
rect 1990 35 2005 55
rect 2025 35 2040 55
rect 1990 20 2040 35
rect 1555 -145 1605 -130
rect 1555 -365 1570 -145
rect 1590 -365 1605 -145
rect 1555 -380 1605 -365
rect 1655 -145 1705 -130
rect 1655 -365 1670 -145
rect 1690 -365 1705 -145
rect 1655 -380 1705 -365
rect 1755 -145 1805 -130
rect 1755 -365 1770 -145
rect 1790 -365 1805 -145
rect 1755 -380 1805 -365
rect 1855 -145 1905 -130
rect 1855 -365 1870 -145
rect 1890 -365 1905 -145
rect 1855 -380 1905 -365
rect 1955 -145 2005 -130
rect 1955 -365 1970 -145
rect 1990 -365 2005 -145
rect 1955 -380 2005 -365
<< pdiff >>
rect 1010 695 1060 710
rect 1010 475 1025 695
rect 1045 475 1060 695
rect 1010 460 1060 475
rect 1110 695 1160 710
rect 1110 475 1125 695
rect 1145 475 1160 695
rect 1110 460 1160 475
rect 1210 695 1260 710
rect 1210 475 1225 695
rect 1245 475 1260 695
rect 1210 460 1260 475
rect 1310 695 1360 710
rect 1310 475 1325 695
rect 1345 475 1360 695
rect 1310 460 1360 475
rect 1410 695 1460 710
rect 1410 475 1425 695
rect 1445 475 1460 695
rect 1410 460 1460 475
rect 1510 695 1560 710
rect 1510 475 1525 695
rect 1545 475 1560 695
rect 1510 460 1560 475
rect 1610 695 1660 710
rect 1610 475 1625 695
rect 1645 475 1660 695
rect 1610 460 1660 475
rect 1710 695 1760 710
rect 1710 475 1725 695
rect 1745 475 1760 695
rect 1710 460 1760 475
rect 1810 695 1860 710
rect 1810 475 1825 695
rect 1845 475 1860 695
rect 1810 460 1860 475
rect 990 330 1040 345
rect 990 260 1005 330
rect 1025 260 1040 330
rect 990 245 1040 260
rect 1055 330 1105 345
rect 1055 260 1070 330
rect 1090 260 1105 330
rect 1055 245 1105 260
rect 1120 330 1170 345
rect 1120 260 1135 330
rect 1155 260 1170 330
rect 1120 245 1170 260
rect 1185 330 1235 345
rect 1185 260 1200 330
rect 1220 260 1235 330
rect 1185 245 1235 260
rect 1250 330 1300 345
rect 1350 330 1400 345
rect 1250 260 1265 330
rect 1285 260 1300 330
rect 1350 260 1365 330
rect 1385 260 1400 330
rect 1250 245 1300 260
rect 1350 245 1400 260
rect 1415 330 1465 345
rect 1415 260 1430 330
rect 1450 260 1465 330
rect 1415 245 1465 260
rect 1480 330 1530 345
rect 1480 260 1495 330
rect 1515 260 1530 330
rect 1480 245 1530 260
rect 1545 330 1595 345
rect 1545 260 1560 330
rect 1580 260 1595 330
rect 1545 245 1595 260
rect 1610 330 1660 345
rect 1610 260 1625 330
rect 1645 260 1660 330
rect 1610 245 1660 260
rect 1730 330 1780 345
rect 1730 260 1745 330
rect 1765 260 1780 330
rect 1730 245 1780 260
rect 1795 330 1845 345
rect 1795 260 1810 330
rect 1830 260 1845 330
rect 1795 245 1845 260
rect 1860 330 1910 345
rect 1860 260 1875 330
rect 1895 260 1910 330
rect 1860 245 1910 260
rect 1925 330 1975 345
rect 1925 260 1940 330
rect 1960 260 1975 330
rect 1925 245 1975 260
rect 1990 330 2040 345
rect 1990 260 2005 330
rect 2025 260 2040 330
rect 1990 245 2040 260
<< ndiffc >>
rect 1005 35 1025 55
rect 1070 35 1090 55
rect 1135 35 1155 55
rect 1200 35 1220 55
rect 1265 35 1285 55
rect 1365 35 1385 55
rect 1430 35 1450 55
rect 1495 35 1515 55
rect 1560 35 1580 55
rect 1625 35 1645 55
rect 1745 35 1765 55
rect 1810 35 1830 55
rect 1875 35 1895 55
rect 1940 35 1960 55
rect 2005 35 2025 55
rect 1570 -365 1590 -145
rect 1670 -365 1690 -145
rect 1770 -365 1790 -145
rect 1870 -365 1890 -145
rect 1970 -365 1990 -145
<< pdiffc >>
rect 1025 475 1045 695
rect 1125 475 1145 695
rect 1225 475 1245 695
rect 1325 475 1345 695
rect 1425 475 1445 695
rect 1525 475 1545 695
rect 1625 475 1645 695
rect 1725 475 1745 695
rect 1825 475 1845 695
rect 1005 260 1025 330
rect 1070 260 1090 330
rect 1135 260 1155 330
rect 1200 260 1220 330
rect 1265 260 1285 330
rect 1365 260 1385 330
rect 1430 260 1450 330
rect 1495 260 1515 330
rect 1560 260 1580 330
rect 1625 260 1645 330
rect 1745 260 1765 330
rect 1810 260 1830 330
rect 1875 260 1895 330
rect 1940 260 1960 330
rect 2005 260 2025 330
<< psubdiff >>
rect 1300 55 1350 70
rect 1300 35 1315 55
rect 1335 35 1350 55
rect 1300 20 1350 35
<< nsubdiff >>
rect 1300 330 1350 345
rect 1300 260 1315 330
rect 1335 260 1350 330
rect 1300 245 1350 260
<< psubdiffcont >>
rect 1315 35 1335 55
<< nsubdiffcont >>
rect 1315 260 1335 330
<< poly >>
rect 1215 755 1255 765
rect 1215 735 1225 755
rect 1245 735 1255 755
rect 1615 755 1655 765
rect 1615 735 1625 755
rect 1645 735 1655 755
rect 1060 720 1810 735
rect 1060 710 1110 720
rect 1160 710 1210 720
rect 1260 710 1310 720
rect 1360 710 1410 720
rect 1460 710 1510 720
rect 1560 710 1610 720
rect 1660 710 1710 720
rect 1760 710 1810 720
rect 1060 445 1110 460
rect 1160 445 1210 460
rect 1260 445 1310 460
rect 1360 445 1410 460
rect 1460 445 1510 460
rect 1560 445 1610 460
rect 1660 445 1710 460
rect 1760 445 1810 460
rect 845 385 1250 400
rect 1040 345 1055 385
rect 1105 345 1120 360
rect 1170 345 1185 360
rect 1235 345 1250 385
rect 1400 345 1415 360
rect 1465 345 1480 360
rect 1530 345 1545 360
rect 1595 345 1610 360
rect 1780 345 1795 360
rect 1845 345 1860 360
rect 1910 345 1925 360
rect 1975 345 1990 360
rect 2105 250 2145 260
rect 1040 225 1055 245
rect 1105 235 1120 245
rect 1170 235 1185 245
rect 1105 220 1185 235
rect 1235 220 1250 245
rect 1400 235 1415 245
rect 1465 235 1480 245
rect 1530 235 1545 245
rect 1595 235 1610 245
rect 1780 235 1795 245
rect 1845 235 1860 245
rect 1910 235 1925 245
rect 1975 235 1990 245
rect 2105 235 2115 250
rect 1400 220 1610 235
rect 1685 230 2115 235
rect 2135 230 2145 250
rect 1685 225 2145 230
rect 1105 200 1120 220
rect 1235 205 1320 220
rect 965 185 1120 200
rect 965 -65 980 185
rect 1125 145 1165 155
rect 1125 95 1135 145
rect 1155 95 1165 145
rect 1305 125 1320 205
rect 1485 200 1495 220
rect 1515 200 1525 220
rect 1485 190 1525 200
rect 1685 205 1695 225
rect 1715 220 2145 225
rect 1715 205 1725 220
rect 1685 195 1725 205
rect 1355 180 1395 190
rect 1355 160 1365 180
rect 1385 165 1395 180
rect 1385 160 1650 165
rect 1355 150 1650 160
rect 1715 150 1755 155
rect 1635 145 1755 150
rect 1635 135 1725 145
rect 1305 110 1480 125
rect 1465 95 1480 110
rect 1715 95 1725 135
rect 1745 95 1755 145
rect 1040 80 1250 95
rect 1040 70 1055 80
rect 1105 70 1120 80
rect 1170 70 1185 80
rect 1235 70 1250 80
rect 1400 70 1415 85
rect 1465 80 1545 95
rect 1715 85 2145 95
rect 1465 70 1480 80
rect 1530 70 1545 80
rect 1595 70 1610 85
rect 1715 80 2115 85
rect 1780 70 1795 80
rect 1845 70 1860 80
rect 1910 70 1925 80
rect 1975 70 1990 80
rect 2105 65 2115 80
rect 2135 65 2145 85
rect 2105 55 2145 65
rect 1040 5 1055 20
rect 1105 5 1120 20
rect 1170 5 1185 20
rect 1235 5 1250 20
rect 1400 -20 1415 20
rect 1465 5 1480 20
rect 1530 5 1545 20
rect 1595 -20 1610 20
rect 1780 5 1795 20
rect 1845 5 1860 20
rect 1910 5 1925 20
rect 1975 5 1990 20
rect 1400 -35 1610 -20
rect 1495 -65 1510 -35
rect 850 -80 1510 -65
rect 1605 -130 1655 -115
rect 1705 -130 1755 -115
rect 1805 -130 1855 -115
rect 1905 -130 1955 -115
rect 1605 -390 1655 -380
rect 1705 -390 1755 -380
rect 1805 -390 1855 -380
rect 1905 -390 1955 -380
rect 1605 -405 1955 -390
rect 1760 -425 1770 -405
rect 1790 -425 1800 -405
rect 1760 -435 1800 -425
<< polycont >>
rect 1225 735 1245 755
rect 1625 735 1645 755
rect 2115 230 2135 250
rect 1135 95 1155 145
rect 1495 200 1515 220
rect 1695 205 1715 225
rect 1365 160 1385 180
rect 1725 95 1745 145
rect 2115 65 2135 85
rect 1770 -425 1790 -405
<< xpolycontact >>
rect 2110 745 2145 965
rect 2110 410 2145 630
rect 1010 -415 1230 -130
rect 1280 -415 1500 -130
rect 2110 -260 2145 -40
rect 2110 -565 2145 -345
<< xpolyres >>
rect 2110 630 2145 745
rect 1230 -415 1280 -130
rect 2110 -345 2145 -260
<< locali >>
rect 2165 1070 2205 1080
rect 2125 1050 2175 1070
rect 2195 1050 2205 1070
rect 2125 965 2145 1050
rect 2165 1040 2205 1050
rect 1215 755 1255 765
rect 1215 745 1225 755
rect 955 735 1225 745
rect 1245 745 1255 755
rect 1615 755 1655 765
rect 1615 745 1625 755
rect 1245 735 1625 745
rect 1645 745 1655 755
rect 1645 735 1845 745
rect 955 725 1845 735
rect 955 -130 975 725
rect 1015 695 1055 705
rect 1015 475 1025 695
rect 1045 475 1055 695
rect 1015 465 1055 475
rect 1115 695 1155 705
rect 1115 475 1125 695
rect 1145 475 1155 695
rect 1115 465 1155 475
rect 1215 695 1255 725
rect 1215 475 1225 695
rect 1245 475 1255 695
rect 1215 465 1255 475
rect 1315 695 1355 705
rect 1315 475 1325 695
rect 1345 475 1355 695
rect 1315 465 1355 475
rect 1415 695 1455 705
rect 1415 475 1425 695
rect 1445 475 1455 695
rect 1415 465 1455 475
rect 1515 695 1555 705
rect 1515 475 1525 695
rect 1545 475 1555 695
rect 1515 465 1555 475
rect 1615 695 1655 725
rect 1825 705 1845 725
rect 1615 475 1625 695
rect 1645 475 1655 695
rect 1615 465 1655 475
rect 1715 695 1755 705
rect 1715 475 1725 695
rect 1745 475 1755 695
rect 1715 465 1755 475
rect 1815 695 1855 705
rect 1815 475 1825 695
rect 1845 475 1855 695
rect 1815 465 1855 475
rect 1025 440 1045 465
rect 1425 440 1445 465
rect 1825 440 1845 465
rect 1025 420 1845 440
rect 1225 380 1245 420
rect 2125 380 2145 410
rect 1005 360 1285 380
rect 1005 340 1025 360
rect 1265 340 1285 360
rect 1365 360 1645 380
rect 1365 340 1385 360
rect 1625 340 1645 360
rect 1810 360 2145 380
rect 1810 340 1830 360
rect 1940 340 1960 360
rect 995 330 1035 340
rect 995 260 1005 330
rect 1025 260 1035 330
rect 995 250 1035 260
rect 1060 330 1100 340
rect 1060 260 1070 330
rect 1090 260 1100 330
rect 1060 250 1100 260
rect 1125 330 1165 340
rect 1125 260 1135 330
rect 1155 260 1165 330
rect 1125 250 1165 260
rect 1190 330 1230 340
rect 1190 260 1200 330
rect 1220 260 1230 330
rect 1190 250 1230 260
rect 1255 330 1395 340
rect 1255 260 1265 330
rect 1285 260 1315 330
rect 1335 260 1365 330
rect 1385 260 1395 330
rect 1255 250 1395 260
rect 1420 330 1460 340
rect 1420 260 1430 330
rect 1450 260 1460 330
rect 1420 250 1460 260
rect 1485 330 1525 340
rect 1485 260 1495 330
rect 1515 260 1525 330
rect 1135 155 1155 250
rect 1265 180 1285 250
rect 1485 220 1525 260
rect 1550 330 1590 340
rect 1550 260 1560 330
rect 1580 260 1590 330
rect 1550 250 1590 260
rect 1615 330 1655 340
rect 1615 260 1625 330
rect 1645 260 1655 330
rect 1615 250 1655 260
rect 1735 330 1775 340
rect 1735 260 1745 330
rect 1765 260 1775 330
rect 1735 250 1775 260
rect 1800 330 1840 340
rect 1800 260 1810 330
rect 1830 260 1840 330
rect 1800 250 1840 260
rect 1865 330 1905 340
rect 1865 260 1875 330
rect 1895 260 1905 330
rect 1865 250 1905 260
rect 1930 330 1970 340
rect 1930 260 1940 330
rect 1960 260 1970 330
rect 1930 250 1970 260
rect 1995 330 2035 340
rect 1995 260 2005 330
rect 2025 260 2035 330
rect 2165 305 2205 315
rect 2165 285 2175 305
rect 2195 285 2205 305
rect 2165 275 2205 285
rect 2165 260 2185 275
rect 1995 250 2035 260
rect 2105 250 2185 260
rect 1485 200 1495 220
rect 1515 200 1525 220
rect 1485 190 1525 200
rect 1625 230 1645 250
rect 1685 230 1725 235
rect 1625 225 1725 230
rect 1625 210 1695 225
rect 1355 180 1395 190
rect 1265 160 1365 180
rect 1385 160 1395 180
rect 1125 145 1165 155
rect 1125 95 1135 145
rect 1155 95 1165 145
rect 1125 85 1165 95
rect 1135 65 1155 85
rect 1265 65 1285 160
rect 1355 150 1395 160
rect 1495 65 1515 190
rect 1625 65 1645 210
rect 1685 205 1695 210
rect 1715 205 1725 225
rect 2105 230 2115 250
rect 2135 240 2185 250
rect 2135 230 2145 240
rect 2105 220 2145 230
rect 1685 195 1725 205
rect 2165 185 2185 240
rect 2165 165 3095 185
rect 1715 145 1755 155
rect 1715 95 1725 145
rect 1745 95 1755 145
rect 2165 95 2185 165
rect 1715 85 1755 95
rect 2105 85 2185 95
rect 2105 65 2115 85
rect 2135 75 2185 85
rect 2135 65 2145 75
rect 995 55 1035 65
rect 995 35 1005 55
rect 1025 35 1035 55
rect 995 25 1035 35
rect 1060 55 1100 65
rect 1060 35 1070 55
rect 1090 35 1100 55
rect 1060 25 1100 35
rect 1125 55 1165 65
rect 1125 35 1135 55
rect 1155 35 1165 55
rect 1125 25 1165 35
rect 1190 55 1230 65
rect 1190 35 1200 55
rect 1220 35 1230 55
rect 1190 25 1230 35
rect 1255 55 1395 65
rect 1255 35 1265 55
rect 1285 35 1315 55
rect 1335 35 1365 55
rect 1385 35 1395 55
rect 1255 25 1395 35
rect 1420 55 1460 65
rect 1420 35 1430 55
rect 1450 35 1460 55
rect 1420 25 1460 35
rect 1485 55 1525 65
rect 1485 35 1495 55
rect 1515 35 1525 55
rect 1485 25 1525 35
rect 1550 55 1590 65
rect 1550 35 1560 55
rect 1580 35 1590 55
rect 1550 25 1590 35
rect 1615 55 1655 65
rect 1615 35 1625 55
rect 1645 35 1655 55
rect 1615 25 1655 35
rect 1735 55 1775 65
rect 1735 35 1745 55
rect 1765 35 1775 55
rect 1735 25 1775 35
rect 1800 55 1840 65
rect 1800 35 1810 55
rect 1830 35 1840 55
rect 1800 25 1840 35
rect 1865 55 1905 65
rect 1865 35 1875 55
rect 1895 35 1905 55
rect 1865 25 1905 35
rect 1930 55 1970 65
rect 1930 35 1940 55
rect 1960 35 1970 55
rect 1930 25 1970 35
rect 1995 55 2035 65
rect 2105 55 2145 65
rect 1995 35 2005 55
rect 2025 35 2035 55
rect 1995 25 2035 35
rect 2165 40 2185 75
rect 2165 30 2205 40
rect 1005 5 1025 25
rect 1265 5 1285 25
rect 1005 -15 1285 5
rect 1365 5 1385 25
rect 1495 5 1515 25
rect 1625 5 1645 25
rect 1365 -15 1645 5
rect 1810 5 1830 25
rect 1940 5 1960 25
rect 2165 10 2175 30
rect 2195 10 2205 30
rect 1810 -15 2145 5
rect 2165 0 2205 10
rect 1625 -35 1645 -15
rect 1625 -55 1790 -35
rect 2125 -40 2145 -15
rect 1770 -90 1790 -55
rect 1570 -110 1990 -90
rect 955 -150 1010 -130
rect 1570 -135 1590 -110
rect 1970 -135 1990 -110
rect 1560 -145 1600 -135
rect 1560 -365 1570 -145
rect 1590 -365 1600 -145
rect 1560 -375 1600 -365
rect 1660 -145 1700 -135
rect 1660 -365 1670 -145
rect 1690 -365 1700 -145
rect 1660 -375 1700 -365
rect 1760 -145 1800 -135
rect 1760 -365 1770 -145
rect 1790 -365 1800 -145
rect 1760 -375 1800 -365
rect 1860 -145 1900 -135
rect 1860 -365 1870 -145
rect 1890 -365 1900 -145
rect 1860 -375 1900 -365
rect 1960 -145 2000 -135
rect 1960 -365 1970 -145
rect 1990 -365 2000 -145
rect 1960 -375 2000 -365
rect 1770 -395 1790 -375
rect 1500 -405 1955 -395
rect 1500 -415 1770 -405
rect 1760 -425 1770 -415
rect 1790 -415 1955 -405
rect 1790 -425 1800 -415
rect 1760 -435 1800 -425
rect 2125 -735 2145 -565
rect 2165 -735 2205 -725
rect 2125 -755 2175 -735
rect 2195 -755 2205 -735
rect 2165 -765 2205 -755
<< viali >>
rect 2175 1050 2195 1070
rect 1125 475 1145 695
rect 1325 475 1345 695
rect 1525 475 1545 695
rect 1725 475 1745 695
rect 1315 260 1335 330
rect 1430 260 1450 330
rect 1560 260 1580 330
rect 1745 260 1765 330
rect 1875 260 1895 330
rect 2005 260 2025 330
rect 2175 285 2195 305
rect 1070 35 1090 55
rect 1200 35 1220 55
rect 1315 35 1335 55
rect 1745 35 1765 55
rect 1875 35 1895 55
rect 2005 35 2025 55
rect 2175 10 2195 30
rect 1670 -365 1690 -145
rect 1870 -365 1890 -145
rect 2175 -755 2195 -735
<< metal1 >>
rect 2165 1070 2205 1080
rect 2165 1050 2175 1070
rect 2195 1050 2205 1070
rect 2165 1040 2205 1050
rect 990 695 2040 710
rect 990 475 1125 695
rect 1145 475 1325 695
rect 1345 475 1525 695
rect 1545 475 1725 695
rect 1745 475 2040 695
rect 990 330 2040 475
rect 990 260 1315 330
rect 1335 260 1430 330
rect 1450 260 1560 330
rect 1580 260 1745 330
rect 1765 260 1875 330
rect 1895 260 2005 330
rect 2025 260 2040 330
rect 2165 305 2205 315
rect 2165 285 2175 305
rect 2195 285 2205 305
rect 2165 275 2205 285
rect 990 245 2040 260
rect 990 55 2040 70
rect 990 35 1070 55
rect 1090 35 1200 55
rect 1220 35 1315 55
rect 1335 35 1745 55
rect 1765 35 1875 55
rect 1895 35 2005 55
rect 2025 35 2040 55
rect 990 -145 2040 35
rect 2165 30 2205 40
rect 2165 10 2175 30
rect 2195 10 2205 30
rect 2165 0 2205 10
rect 990 -365 1670 -145
rect 1690 -365 1870 -145
rect 1890 -365 2040 -145
rect 990 -380 2040 -365
rect 2165 -735 2205 -725
rect 2165 -755 2175 -735
rect 2195 -755 2205 -735
rect 2165 -765 2205 -755
<< metal3 >>
rect 2165 1040 3050 1085
rect 2220 255 3050 1040
rect 2220 -725 3050 60
rect 2165 -770 3050 -725
<< mimcap >>
rect 2235 315 3035 1070
rect 2235 280 2245 315
rect 2280 280 3035 315
rect 2235 270 3035 280
rect 2235 35 3035 45
rect 2235 0 2245 35
rect 2280 0 3035 35
rect 2235 -755 3035 0
<< mimcapcontact >>
rect 2245 280 2280 315
rect 2245 0 2280 35
<< metal4 >>
rect 2165 315 2285 320
rect 2165 280 2245 315
rect 2280 280 2285 315
rect 2165 275 2285 280
rect 2165 35 2285 40
rect 2165 0 2245 35
rect 2280 0 2285 35
rect 2165 -5 2285 0
<< labels >>
flabel metal1 990 580 990 580 7 FreeSans 400 0 0 0 VDDA
flabel poly 845 390 845 390 7 FreeSans 400 0 0 0 VIN+
flabel locali 3095 170 3095 170 3 FreeSans 400 0 0 0 VOUT
flabel poly 850 -70 850 -70 7 FreeSans 400 0 0 0 VIN-
flabel metal1 990 -270 990 -270 7 FreeSans 400 0 0 0 GNDA
<< end >>
