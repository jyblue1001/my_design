* PEX produced on Wed Jul  2 09:21:48 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA
X0 a_14640_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA.t323 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X1 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA.t217 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X2 two_stage_opamp_dummy_magic_0.VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 bgr_0.PFET_GATE_10uA.t10 VDDA.t417 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X4 bgr_0.V_mir2.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 bgr_0.V_p_2.t4 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X5 two_stage_opamp_dummy_magic_0.VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 two_stage_opamp_dummy_magic_0.VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 two_stage_opamp_dummy_magic_0.Vb1.t5 bgr_0.PFET_GATE_10uA.t11 VDDA.t415 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X8 two_stage_opamp_dummy_magic_0.VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_0.V_err_gate.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 two_stage_opamp_dummy_magic_0.VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDDA.t117 VDDA.t115 bgr_0.PFET_GATE_10uA.t6 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X13 GNDA.t48 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X14 two_stage_opamp_dummy_magic_0.X.t6 GNDA.t214 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X15 VDDA.t273 bgr_0.1st_Vout_1.t11 bgr_0.V_TOP.t10 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X16 two_stage_opamp_dummy_magic_0.VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 two_stage_opamp_dummy_magic_0.VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 two_stage_opamp_dummy_magic_0.VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VDDA.t127 two_stage_opamp_dummy_magic_0.X.t26 two_stage_opamp_dummy_magic_0.VOUT-.t2 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X20 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 two_stage_opamp_dummy_magic_0.Y.t25 VDDA.t278 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X21 bgr_0.PFET_GATE_10uA.t7 bgr_0.1st_Vout_2.t12 VDDA.t438 VDDA.t437 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X22 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 bgr_0.PFET_GATE_10uA.t12 VDDA.t413 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 two_stage_opamp_dummy_magic_0.VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_5750_2946.t0 GNDA.t258 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X25 two_stage_opamp_dummy_magic_0.VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 bgr_0.V_TOP.t14 VDDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 two_stage_opamp_dummy_magic_0.VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 two_stage_opamp_dummy_magic_0.VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDDA.t319 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X30 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t7 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X31 two_stage_opamp_dummy_magic_0.VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 two_stage_opamp_dummy_magic_0.VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_0.VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 GNDA.t295 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X35 two_stage_opamp_dummy_magic_0.VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 bgr_0.START_UP.t3 bgr_0.V_TOP.t15 VDDA.t300 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X37 VDDA.t172 two_stage_opamp_dummy_magic_0.Vb3.t8 two_stage_opamp_dummy_magic_0.VD3.t15 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X38 bgr_0.V_TOP.t16 VDDA.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VDDA.t114 VDDA.t112 two_stage_opamp_dummy_magic_0.V_err_gate.t1 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X40 two_stage_opamp_dummy_magic_0.VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 two_stage_opamp_dummy_magic_0.VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 two_stage_opamp_dummy_magic_0.Y.t5 GNDA.t211 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X44 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X45 two_stage_opamp_dummy_magic_0.VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 two_stage_opamp_dummy_magic_0.VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 two_stage_opamp_dummy_magic_0.V_err_p.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t277 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X48 two_stage_opamp_dummy_magic_0.VOUT-.t3 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X49 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 two_stage_opamp_dummy_magic_0.VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 bgr_0.1st_Vout_2.t10 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t10 GNDA.t354 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X52 bgr_0.PFET_GATE_10uA.t8 bgr_0.1st_Vout_2.t13 VDDA.t440 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t37 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X54 two_stage_opamp_dummy_magic_0.VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 two_stage_opamp_dummy_magic_0.VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 two_stage_opamp_dummy_magic_0.VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 two_stage_opamp_dummy_magic_0.V_err_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X59 two_stage_opamp_dummy_magic_0.VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 two_stage_opamp_dummy_magic_0.VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 GNDA.t33 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X62 two_stage_opamp_dummy_magic_0.VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 VDDA.t280 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t1 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X64 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t36 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X65 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 bgr_0.PFET_GATE_10uA.t13 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X66 bgr_0.V_TOP.t17 VDDA.t257 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 GNDA.t339 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 VDDA.t419 two_stage_opamp_dummy_magic_0.Vb3.t9 two_stage_opamp_dummy_magic_0.VD3.t29 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X69 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 two_stage_opamp_dummy_magic_0.VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_0.Vb1.t1 VDDA.t109 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X72 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X73 bgr_0.1st_Vout_1.t8 bgr_0.Vin+.t6 bgr_0.V_p_1.t9 GNDA.t327 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X74 two_stage_opamp_dummy_magic_0.VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 GNDA.t53 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 two_stage_opamp_dummy_magic_0.VOUT+.t3 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X76 GNDA.t284 two_stage_opamp_dummy_magic_0.X.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X77 GNDA.t237 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X78 VDDA.t108 VDDA.t106 bgr_0.V_TOP.t3 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X79 GNDA.t210 GNDA.t208 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X80 two_stage_opamp_dummy_magic_0.VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t15 VDDA.t442 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 two_stage_opamp_dummy_magic_0.VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 two_stage_opamp_dummy_magic_0.VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 two_stage_opamp_dummy_magic_0.VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t103 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X86 two_stage_opamp_dummy_magic_0.VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 GNDA.t73 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X88 two_stage_opamp_dummy_magic_0.VOUT+.t17 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X89 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t9 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X90 GNDA.t207 GNDA.t205 GNDA.t207 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X91 GNDA.t204 GNDA.t202 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X92 VDDA.t362 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X93 VDDA.t291 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t2 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X94 two_stage_opamp_dummy_magic_0.VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 GNDA.t201 GNDA.t199 two_stage_opamp_dummy_magic_0.VOUT+.t7 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X97 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t29 VDDA.t317 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X98 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X99 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t423 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X100 GNDA.t178 GNDA.t176 two_stage_opamp_dummy_magic_0.X.t5 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X101 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 bgr_0.V_TOP.t18 VDDA.t196 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X102 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t356 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X103 two_stage_opamp_dummy_magic_0.VOUT-.t4 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X104 two_stage_opamp_dummy_magic_0.VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 two_stage_opamp_dummy_magic_0.VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 two_stage_opamp_dummy_magic_0.VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 two_stage_opamp_dummy_magic_0.VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 two_stage_opamp_dummy_magic_0.VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 a_14640_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t244 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X111 two_stage_opamp_dummy_magic_0.VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 two_stage_opamp_dummy_magic_0.VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 two_stage_opamp_dummy_magic_0.VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 VDDA.t102 VDDA.t100 two_stage_opamp_dummy_magic_0.VD3.t1 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X115 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 bgr_0.NFET_GATE_10uA.t7 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_0.VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VDDA.t198 bgr_0.V_TOP.t19 bgr_0.START_UP.t2 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X118 GNDA.t286 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t324 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X119 two_stage_opamp_dummy_magic_0.VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VDDA.t138 two_stage_opamp_dummy_magic_0.X.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X121 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 bgr_0.PFET_GATE_10uA.t14 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X122 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X123 two_stage_opamp_dummy_magic_0.VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 GNDA.t198 GNDA.t196 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X125 GNDA.t46 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X126 GNDA.t239 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X127 two_stage_opamp_dummy_magic_0.VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 GNDA.t47 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X129 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X130 VDDA.t253 bgr_0.1st_Vout_2.t18 bgr_0.PFET_GATE_10uA.t3 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X131 two_stage_opamp_dummy_magic_0.VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 two_stage_opamp_dummy_magic_0.VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 bgr_0.Vin-.t7 bgr_0.START_UP.t6 bgr_0.V_TOP.t11 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X135 two_stage_opamp_dummy_magic_0.V_p.t9 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X136 two_stage_opamp_dummy_magic_0.VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 two_stage_opamp_dummy_magic_0.VOUT-.t16 a_5750_2946.t1 GNDA.t271 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X138 two_stage_opamp_dummy_magic_0.VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 two_stage_opamp_dummy_magic_0.VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 a_29640_9790.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X141 VDDA.t179 bgr_0.V_TOP.t20 bgr_0.Vin+.t5 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X142 two_stage_opamp_dummy_magic_0.VOUT+.t16 two_stage_opamp_dummy_magic_0.Y.t29 VDDA.t468 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X143 two_stage_opamp_dummy_magic_0.V_p.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X144 two_stage_opamp_dummy_magic_0.V_p.t8 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X145 two_stage_opamp_dummy_magic_0.VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 bgr_0.V_TOP.t21 VDDA.t180 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 two_stage_opamp_dummy_magic_0.VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X149 two_stage_opamp_dummy_magic_0.VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_0.V_p_1.t10 bgr_0.Vin-.t8 bgr_0.V_mir1.t16 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X151 two_stage_opamp_dummy_magic_0.VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 two_stage_opamp_dummy_magic_0.VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 two_stage_opamp_dummy_magic_0.Vb2.t6 bgr_0.NFET_GATE_10uA.t8 GNDA.t35 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X154 two_stage_opamp_dummy_magic_0.VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VDDA.t99 VDDA.t97 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X156 two_stage_opamp_dummy_magic_0.VOUT+.t6 GNDA.t193 GNDA.t195 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X157 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 VDDA.t94 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X158 two_stage_opamp_dummy_magic_0.VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 bgr_0.V_TOP.t22 VDDA.t274 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 two_stage_opamp_dummy_magic_0.VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 two_stage_opamp_dummy_magic_0.VD2.t18 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t20 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X162 GNDA.t346 bgr_0.NFET_GATE_10uA.t9 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X163 bgr_0.V_p_2.t1 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t6 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X164 two_stage_opamp_dummy_magic_0.VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 two_stage_opamp_dummy_magic_0.VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 two_stage_opamp_dummy_magic_0.VOUT-.t0 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X167 VDDA.t255 bgr_0.1st_Vout_2.t19 bgr_0.PFET_GATE_10uA.t4 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X168 two_stage_opamp_dummy_magic_0.VOUT-.t1 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t125 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X169 VDDA.t313 bgr_0.V_mir1.t14 bgr_0.V_mir1.t15 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 VDDA.t267 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X171 two_stage_opamp_dummy_magic_0.VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 two_stage_opamp_dummy_magic_0.VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 two_stage_opamp_dummy_magic_0.VOUT-.t9 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t100 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X174 two_stage_opamp_dummy_magic_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t10 GNDA.t294 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X175 bgr_0.V_mir1.t13 bgr_0.V_mir1.t12 VDDA.t430 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X176 bgr_0.V_TOP.t23 VDDA.t275 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t9 GNDA.t307 sky130_fd_pr__res_high_po_1p41 l=1.41
X178 two_stage_opamp_dummy_magic_0.VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 GNDA.t95 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X180 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 two_stage_opamp_dummy_magic_0.VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 GNDA.t137 GNDA.t181 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X183 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.Vb3.t11 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X184 two_stage_opamp_dummy_magic_0.VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X186 bgr_0.V_p_1.t8 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t7 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X187 two_stage_opamp_dummy_magic_0.err_amp_out.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t342 GNDA.t341 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X188 VDDA.t201 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X189 bgr_0.V_CUR_REF_REG.t0 VDDA.t63 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X190 two_stage_opamp_dummy_magic_0.VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 bgr_0.PFET_GATE_10uA.t15 VDDA.t407 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X192 two_stage_opamp_dummy_magic_0.VD1.t20 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t12 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X193 two_stage_opamp_dummy_magic_0.VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 two_stage_opamp_dummy_magic_0.VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VDDA.t93 VDDA.t91 two_stage_opamp_dummy_magic_0.V_err_p.t2 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X197 two_stage_opamp_dummy_magic_0.VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_0.VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 GNDA.t4 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X200 two_stage_opamp_dummy_magic_0.VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 GNDA.t137 GNDA.t192 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X202 two_stage_opamp_dummy_magic_0.err_amp_out.t11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X203 GNDA.t94 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X204 a_5230_5758.t1 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t254 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X205 bgr_0.Vin-.t5 bgr_0.V_TOP.t24 VDDA.t444 VDDA.t443 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X206 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 two_stage_opamp_dummy_magic_0.VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 two_stage_opamp_dummy_magic_0.VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 two_stage_opamp_dummy_magic_0.VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 two_stage_opamp_dummy_magic_0.VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 two_stage_opamp_dummy_magic_0.VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_0.V_p.t7 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X214 two_stage_opamp_dummy_magic_0.V_p.t23 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X215 two_stage_opamp_dummy_magic_0.VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VDDA.t185 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD4.t11 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X217 two_stage_opamp_dummy_magic_0.VOUT+.t15 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t302 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X218 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X219 two_stage_opamp_dummy_magic_0.V_p.t35 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X220 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA.t189 GNDA.t191 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X221 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t11 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X222 VDDA.t121 bgr_0.V_mir2.t8 bgr_0.V_mir2.t9 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X223 two_stage_opamp_dummy_magic_0.VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t9 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X225 two_stage_opamp_dummy_magic_0.VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 two_stage_opamp_dummy_magic_0.VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 two_stage_opamp_dummy_magic_0.VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 bgr_0.V_TOP.t25 VDDA.t445 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 two_stage_opamp_dummy_magic_0.VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 two_stage_opamp_dummy_magic_0.VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 GNDA.t314 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X233 a_14520_5738.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t270 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X234 two_stage_opamp_dummy_magic_0.VOUT-.t6 two_stage_opamp_dummy_magic_0.X.t38 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X235 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 bgr_0.V_TOP.t26 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X236 two_stage_opamp_dummy_magic_0.VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VDDA.t456 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA.t348 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X238 bgr_0.V_mir1.t9 bgr_0.V_mir1.t8 VDDA.t315 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X239 two_stage_opamp_dummy_magic_0.VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 bgr_0.V_TOP.t27 VDDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 two_stage_opamp_dummy_magic_0.VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 two_stage_opamp_dummy_magic_0.VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 two_stage_opamp_dummy_magic_0.VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 two_stage_opamp_dummy_magic_0.VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t88 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X246 GNDA.t288 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X247 two_stage_opamp_dummy_magic_0.VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 bgr_0.PFET_GATE_10uA.t5 VDDA.t85 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X250 GNDA.t224 VDDA.t469 bgr_0.V_TOP.t4 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X251 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 GNDA.t289 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t327 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X253 two_stage_opamp_dummy_magic_0.VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 two_stage_opamp_dummy_magic_0.VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X256 bgr_0.V_TOP.t28 VDDA.t207 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X258 VDDA.t161 two_stage_opamp_dummy_magic_0.X.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X259 two_stage_opamp_dummy_magic_0.VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X261 VDDA.t286 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X262 two_stage_opamp_dummy_magic_0.VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 two_stage_opamp_dummy_magic_0.VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 two_stage_opamp_dummy_magic_0.VD1.t19 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t16 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X266 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 two_stage_opamp_dummy_magic_0.VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VDDA.t358 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X269 bgr_0.V_TOP.t9 bgr_0.1st_Vout_1.t18 VDDA.t271 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X270 VDDA.t352 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X271 bgr_0.Vin-.t4 bgr_0.V_TOP.t29 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X272 GNDA.t231 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X273 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X274 GNDA.t246 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X275 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X276 two_stage_opamp_dummy_magic_0.V_p.t34 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X277 GNDA.t221 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X278 two_stage_opamp_dummy_magic_0.VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 bgr_0.V_TOP.t30 VDDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 a_29640_9790.t1 GNDA.t257 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X281 two_stage_opamp_dummy_magic_0.VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 two_stage_opamp_dummy_magic_0.VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 two_stage_opamp_dummy_magic_0.VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 bgr_0.V_mir2.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 bgr_0.V_p_2.t3 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X286 two_stage_opamp_dummy_magic_0.VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VDDA.t375 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD3.t26 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X288 two_stage_opamp_dummy_magic_0.VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 two_stage_opamp_dummy_magic_0.VOUT+.t14 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X290 bgr_0.1st_Vout_1.t6 bgr_0.Vin+.t8 bgr_0.V_p_1.t7 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X291 two_stage_opamp_dummy_magic_0.V_p.t33 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X292 two_stage_opamp_dummy_magic_0.V_p.t21 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA.t281 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X293 two_stage_opamp_dummy_magic_0.VOUT+.t13 two_stage_opamp_dummy_magic_0.Y.t37 VDDA.t321 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X294 two_stage_opamp_dummy_magic_0.VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 two_stage_opamp_dummy_magic_0.VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t186 GNDA.t188 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X299 VDDA.t84 VDDA.t82 bgr_0.NFET_GATE_10uA.t0 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X300 two_stage_opamp_dummy_magic_0.VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 two_stage_opamp_dummy_magic_0.VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t21 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X305 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X306 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 bgr_0.PFET_GATE_10uA.t16 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X307 GNDA.t15 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X308 GNDA.t185 GNDA.t183 bgr_0.NFET_GATE_10uA.t1 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X309 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X310 two_stage_opamp_dummy_magic_0.VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 two_stage_opamp_dummy_magic_0.VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VDDA.t311 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X314 two_stage_opamp_dummy_magic_0.VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 two_stage_opamp_dummy_magic_0.VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 two_stage_opamp_dummy_magic_0.VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VDDA.t462 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X318 two_stage_opamp_dummy_magic_0.VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_0.VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 two_stage_opamp_dummy_magic_0.VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VDDA.t81 VDDA.t79 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X322 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t76 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X323 bgr_0.V_mir1.t0 bgr_0.Vin-.t9 bgr_0.V_p_1.t1 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X324 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t354 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X325 GNDA.t267 VDDA.t73 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X326 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X327 two_stage_opamp_dummy_magic_0.VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 two_stage_opamp_dummy_magic_0.VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_0.VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VDDA.t287 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X332 two_stage_opamp_dummy_magic_0.VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VDDA.t308 bgr_0.V_TOP.t31 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X334 two_stage_opamp_dummy_magic_0.VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 two_stage_opamp_dummy_magic_0.VD1.t18 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.Y.t11 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X336 VDDA.t348 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X337 a_5350_5758.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t222 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X338 GNDA.t283 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_p_mir.t2 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X339 two_stage_opamp_dummy_magic_0.VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X342 two_stage_opamp_dummy_magic_0.VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 GNDA.t113 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X344 two_stage_opamp_dummy_magic_0.VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 two_stage_opamp_dummy_magic_0.VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_p.t18 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X347 VDDA.t200 bgr_0.V_mir1.t4 bgr_0.V_mir1.t5 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X348 two_stage_opamp_dummy_magic_0.V_p.t6 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X349 two_stage_opamp_dummy_magic_0.VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 two_stage_opamp_dummy_magic_0.VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GNDA.t137 GNDA.t179 bgr_0.Vin-.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X352 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.Vb3.t14 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X353 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X354 VDDA.t72 VDDA.t69 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X355 GNDA.t135 GNDA.t175 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X356 two_stage_opamp_dummy_magic_0.VOUT+.t2 VDDA.t66 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X357 two_stage_opamp_dummy_magic_0.V_p.t5 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X358 two_stage_opamp_dummy_magic_0.V_p.t19 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t115 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X359 two_stage_opamp_dummy_magic_0.VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 two_stage_opamp_dummy_magic_0.VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VDDA.t451 bgr_0.V_TOP.t32 bgr_0.Vin-.t3 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X362 GNDA.t137 GNDA.t182 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X363 two_stage_opamp_dummy_magic_0.VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 two_stage_opamp_dummy_magic_0.VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t8 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X367 two_stage_opamp_dummy_magic_0.VD2.t12 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t18 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X368 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 GNDA.t135 GNDA.t180 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X370 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 bgr_0.PFET_GATE_10uA.t17 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X371 two_stage_opamp_dummy_magic_0.VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 two_stage_opamp_dummy_magic_0.VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VDDA.t310 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X374 two_stage_opamp_dummy_magic_0.VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 GNDA.t39 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X376 VDDA.t325 two_stage_opamp_dummy_magic_0.Y.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X377 VDDA.t251 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t2 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X378 two_stage_opamp_dummy_magic_0.VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t22 GNDA.t350 sky130_fd_pr__res_high_po_1p41 l=1.41
X380 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X381 bgr_0.V_TOP.t33 VDDA.t452 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VDDA.t401 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X383 two_stage_opamp_dummy_magic_0.VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 two_stage_opamp_dummy_magic_0.V_err_p.t8 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t350 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X385 two_stage_opamp_dummy_magic_0.VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.VD3.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X387 two_stage_opamp_dummy_magic_0.VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 bgr_0.PFET_GATE_10uA.t1 VDDA.t470 GNDA.t225 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X389 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA.t269 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X390 two_stage_opamp_dummy_magic_0.VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VDDA.t62 VDDA.t60 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X392 VDDA.t206 bgr_0.1st_Vout_1.t24 bgr_0.V_TOP.t7 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X393 two_stage_opamp_dummy_magic_0.VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb3.t15 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X396 two_stage_opamp_dummy_magic_0.VD1.t17 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t18 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X397 VDDA.t364 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t7 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X398 a_27130_9400.t0 a_28738_9040.t0 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X399 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X400 two_stage_opamp_dummy_magic_0.VD1.t16 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X401 two_stage_opamp_dummy_magic_0.VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 two_stage_opamp_dummy_magic_0.VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 two_stage_opamp_dummy_magic_0.VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t174 GNDA.t171 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X405 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X406 GNDA.t17 VDDA.t57 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X407 bgr_0.Vin+.t1 a_28738_9040.t1 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X408 GNDA.t137 GNDA.t170 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X409 VDDA.t332 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X410 bgr_0.V_p_2.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 bgr_0.V_mir2.t14 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X411 two_stage_opamp_dummy_magic_0.VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 two_stage_opamp_dummy_magic_0.V_p.t32 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X413 bgr_0.V_p_1.t6 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t4 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X414 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 two_stage_opamp_dummy_magic_0.VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 two_stage_opamp_dummy_magic_0.VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 two_stage_opamp_dummy_magic_0.VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VDDA.t366 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VDDA.t56 VDDA.t54 GNDA.t75 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X420 two_stage_opamp_dummy_magic_0.VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 two_stage_opamp_dummy_magic_0.VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 GNDA.t265 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X423 two_stage_opamp_dummy_magic_0.VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 two_stage_opamp_dummy_magic_0.VOUT+.t0 a_14240_2946.t0 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X425 VDDA.t399 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X426 VDDA.t53 VDDA.t51 bgr_0.V_TOP.t2 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X427 two_stage_opamp_dummy_magic_0.VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 bgr_0.NFET_GATE_10uA.t15 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X429 VDDA.t397 bgr_0.PFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X430 two_stage_opamp_dummy_magic_0.VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 two_stage_opamp_dummy_magic_0.VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X433 two_stage_opamp_dummy_magic_0.VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 two_stage_opamp_dummy_magic_0.VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 two_stage_opamp_dummy_magic_0.VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t3 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X437 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X438 bgr_0.V_TOP.t6 bgr_0.1st_Vout_1.t26 VDDA.t204 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X439 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t42 GNDA.t42 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X440 two_stage_opamp_dummy_magic_0.VOUT-.t15 VDDA.t48 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X441 VDDA.t233 GNDA.t167 GNDA.t169 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X442 VDDA.t152 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.VD4.t8 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X443 bgr_0.V_p_1.t3 bgr_0.Vin-.t10 bgr_0.V_mir1.t2 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X444 two_stage_opamp_dummy_magic_0.VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 two_stage_opamp_dummy_magic_0.VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t45 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X447 VDDA.t395 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X448 bgr_0.START_UP.t1 bgr_0.V_TOP.t34 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X449 two_stage_opamp_dummy_magic_0.VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 bgr_0.NFET_GATE_10uA.t16 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X451 VDDA.t44 VDDA.t42 two_stage_opamp_dummy_magic_0.VOUT+.t1 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X452 two_stage_opamp_dummy_magic_0.VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X454 two_stage_opamp_dummy_magic_0.VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 two_stage_opamp_dummy_magic_0.VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA.t165 GNDA.t166 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X457 two_stage_opamp_dummy_magic_0.VOUT+.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t309 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X458 two_stage_opamp_dummy_magic_0.VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 two_stage_opamp_dummy_magic_0.VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 a_5350_5758.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA.t243 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X461 bgr_0.V_TOP.t35 VDDA.t246 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_0.VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 a_27130_9400.t1 GNDA.t251 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X464 VDDA.t119 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X465 two_stage_opamp_dummy_magic_0.V_err_gate.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X466 bgr_0.V_p_1.t0 VDDA.t471 GNDA.t227 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X467 two_stage_opamp_dummy_magic_0.VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VDDA.t218 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X469 VDDA.t158 two_stage_opamp_dummy_magic_0.X.t43 two_stage_opamp_dummy_magic_0.VOUT-.t5 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X470 bgr_0.Vin-.t0 a_28738_9160.t0 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X471 bgr_0.V_TOP.t13 bgr_0.cap_res1.t20 GNDA.t7 sky130_fd_pr__res_high_po_0p35 l=2.05
X472 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 VDDA.t39 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X473 VDDA.t465 two_stage_opamp_dummy_magic_0.Vb3.t18 two_stage_opamp_dummy_magic_0.VD4.t7 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X474 two_stage_opamp_dummy_magic_0.VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 two_stage_opamp_dummy_magic_0.VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 bgr_0.V_TOP.t36 VDDA.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 two_stage_opamp_dummy_magic_0.VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 two_stage_opamp_dummy_magic_0.Y.t0 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X479 two_stage_opamp_dummy_magic_0.V_p.t4 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X480 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X482 two_stage_opamp_dummy_magic_0.VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 GNDA.t164 GNDA.t162 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X484 two_stage_opamp_dummy_magic_0.VOUT+.t4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X485 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X486 two_stage_opamp_dummy_magic_0.VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 two_stage_opamp_dummy_magic_0.VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t353 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X489 two_stage_opamp_dummy_magic_0.VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 VDDA.t393 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X492 bgr_0.V_TOP.t37 VDDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 two_stage_opamp_dummy_magic_0.VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VDDA.t377 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.VD4.t6 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X496 VDDA.t38 VDDA.t36 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X497 two_stage_opamp_dummy_magic_0.VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 two_stage_opamp_dummy_magic_0.V_p.t18 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA.t88 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X499 two_stage_opamp_dummy_magic_0.V_p.t17 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X500 two_stage_opamp_dummy_magic_0.VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t44 GNDA.t261 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X502 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X503 bgr_0.V_mir2.t5 bgr_0.V_mir2.t4 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X504 VDDA.t35 VDDA.t33 GNDA.t266 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X505 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 two_stage_opamp_dummy_magic_0.VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 bgr_0.V_TOP.t12 bgr_0.START_UP.t7 bgr_0.Vin-.t6 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X508 two_stage_opamp_dummy_magic_0.VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 two_stage_opamp_dummy_magic_0.VD1.t7 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t31 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X511 two_stage_opamp_dummy_magic_0.VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 two_stage_opamp_dummy_magic_0.VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 bgr_0.V_TOP.t38 VDDA.t289 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 two_stage_opamp_dummy_magic_0.VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 two_stage_opamp_dummy_magic_0.VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 two_stage_opamp_dummy_magic_0.VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 two_stage_opamp_dummy_magic_0.VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X519 GNDA.t277 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA.t276 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X520 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA.t159 GNDA.t161 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X521 VDDA.t304 two_stage_opamp_dummy_magic_0.Y.t42 two_stage_opamp_dummy_magic_0.VOUT+.t12 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X522 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t297 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X523 two_stage_opamp_dummy_magic_0.VD1.t2 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t30 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X524 two_stage_opamp_dummy_magic_0.VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 two_stage_opamp_dummy_magic_0.VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 two_stage_opamp_dummy_magic_0.VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 two_stage_opamp_dummy_magic_0.VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 GNDA.t158 GNDA.t156 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X530 a_27130_9280.t1 GNDA.t242 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X531 two_stage_opamp_dummy_magic_0.VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 two_stage_opamp_dummy_magic_0.VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VDDA.t435 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t5 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X534 VDDA.t232 GNDA.t153 GNDA.t155 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X535 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X536 VDDA.t391 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X537 a_27130_9280.t0 a_28738_9160.t1 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X538 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X539 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t2 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X540 two_stage_opamp_dummy_magic_0.VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 two_stage_opamp_dummy_magic_0.V_err_gate.t13 bgr_0.NFET_GATE_10uA.t17 GNDA.t329 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X542 VDDA.t285 two_stage_opamp_dummy_magic_0.X.t45 two_stage_opamp_dummy_magic_0.VOUT-.t13 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X543 VDDA.t293 bgr_0.V_TOP.t39 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X544 two_stage_opamp_dummy_magic_0.VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VDDA.t32 VDDA.t30 two_stage_opamp_dummy_magic_0.VOUT-.t14 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X546 bgr_0.V_mir2.t3 bgr_0.V_mir2.t2 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X547 GNDA.t152 GNDA.t150 VDDA.t231 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X548 bgr_0.V_mir1.t3 bgr_0.Vin-.t11 bgr_0.V_p_1.t4 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X549 two_stage_opamp_dummy_magic_0.VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 two_stage_opamp_dummy_magic_0.VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VDDA.t295 bgr_0.V_TOP.t40 bgr_0.START_UP.t0 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X552 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_0.VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 two_stage_opamp_dummy_magic_0.VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 GNDA.t6 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X556 two_stage_opamp_dummy_magic_0.VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 two_stage_opamp_dummy_magic_0.VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_14240_2946.t1 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X559 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 two_stage_opamp_dummy_magic_0.Y.t43 GNDA.t305 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X560 two_stage_opamp_dummy_magic_0.VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 two_stage_opamp_dummy_magic_0.VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 two_stage_opamp_dummy_magic_0.VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 GNDA.t149 GNDA.t147 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X565 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X566 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t176 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X567 VDDA.t389 bgr_0.PFET_GATE_10uA.t24 bgr_0.V_CUR_REF_REG.t1 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X568 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t17 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X569 VDDA.t387 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X570 two_stage_opamp_dummy_magic_0.VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 two_stage_opamp_dummy_magic_0.VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X573 two_stage_opamp_dummy_magic_0.VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 GNDA.t344 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA.t343 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X576 two_stage_opamp_dummy_magic_0.VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 GNDA.t137 GNDA.t136 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X578 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X579 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t6 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X580 two_stage_opamp_dummy_magic_0.VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb3.t22 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X582 VDDA.t225 bgr_0.V_TOP.t41 bgr_0.Vin-.t2 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X583 two_stage_opamp_dummy_magic_0.VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 two_stage_opamp_dummy_magic_0.VD2.t15 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X585 bgr_0.1st_Vout_1.t9 bgr_0.Vin+.t10 bgr_0.V_p_1.t5 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X586 two_stage_opamp_dummy_magic_0.V_p.t15 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA.t279 GNDA.t278 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X587 GNDA.t135 GNDA.t134 bgr_0.Vbe2.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X588 VDDA.t29 VDDA.t27 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X589 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t47 GNDA.t67 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X590 VDDA.t447 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD3.t35 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X591 bgr_0.V_TOP.t1 VDDA.t24 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X592 GNDA.t98 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 two_stage_opamp_dummy_magic_0.VOUT+.t5 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X593 two_stage_opamp_dummy_magic_0.VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 bgr_0.Vin+.t0 bgr_0.Vbe2.t8 GNDA.t241 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X596 GNDA.t298 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X597 VDDA.t458 two_stage_opamp_dummy_magic_0.Y.t44 two_stage_opamp_dummy_magic_0.VOUT+.t11 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X598 a_5230_5758.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t250 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X599 GNDA.t146 GNDA.t144 two_stage_opamp_dummy_magic_0.VOUT-.t11 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X600 two_stage_opamp_dummy_magic_0.VD2.t5 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.V_p.t3 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X601 two_stage_opamp_dummy_magic_0.VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 bgr_0.1st_Vout_2.t4 bgr_0.V_mir2.t18 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X603 two_stage_opamp_dummy_magic_0.VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 GNDA.t77 bgr_0.NFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X605 bgr_0.PFET_GATE_10uA.t0 bgr_0.cap_res2.t0 GNDA.t7 sky130_fd_pr__res_high_po_0p35 l=2.05
X606 two_stage_opamp_dummy_magic_0.VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 two_stage_opamp_dummy_magic_0.V_err_gate.t5 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X609 two_stage_opamp_dummy_magic_0.VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 VDDA.t21 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X611 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X612 two_stage_opamp_dummy_magic_0.VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_0.VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 bgr_0.V_TOP.t42 VDDA.t226 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X616 two_stage_opamp_dummy_magic_0.Vb3.t2 bgr_0.NFET_GATE_10uA.t20 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X617 two_stage_opamp_dummy_magic_0.VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_0.VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 VDDA.t174 two_stage_opamp_dummy_magic_0.X.t48 two_stage_opamp_dummy_magic_0.VOUT-.t7 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X620 VDDA.t334 two_stage_opamp_dummy_magic_0.Vb3.t24 two_stage_opamp_dummy_magic_0.VD3.t23 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X621 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t309 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X622 a_29700_9260.t0 GNDA.t256 GNDA.t255 sky130_fd_pr__res_xhigh_po_0p35 l=6
X623 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.VD3.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X624 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X625 two_stage_opamp_dummy_magic_0.VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 GNDA.t11 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X627 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_0.Y.t46 GNDA.t29 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X628 two_stage_opamp_dummy_magic_0.VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_0.VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t306 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X631 two_stage_opamp_dummy_magic_0.VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X633 bgr_0.1st_Vout_2.t3 bgr_0.V_mir2.t19 VDDA.t344 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X634 two_stage_opamp_dummy_magic_0.VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 GNDA.t249 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X636 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t175 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X637 GNDA.t143 GNDA.t141 VDDA.t230 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X638 VDDA.t385 bgr_0.PFET_GATE_10uA.t26 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X639 two_stage_opamp_dummy_magic_0.VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 two_stage_opamp_dummy_magic_0.VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VDDA.t235 bgr_0.V_mir2.t0 bgr_0.V_mir2.t1 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X642 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X643 VDDA.t239 bgr_0.1st_Vout_1.t34 bgr_0.V_TOP.t5 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X644 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_0.VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 two_stage_opamp_dummy_magic_0.VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X648 two_stage_opamp_dummy_magic_0.V_p.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA.t300 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X649 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X650 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t315 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X651 two_stage_opamp_dummy_magic_0.VD2.t7 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.V_p.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X652 GNDA.t140 GNDA.t138 GNDA.t140 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X653 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X654 GNDA.t133 GNDA.t131 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X655 two_stage_opamp_dummy_magic_0.VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 two_stage_opamp_dummy_magic_0.VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VDDA.t449 bgr_0.V_mir1.t20 bgr_0.1st_Vout_1.t10 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X658 two_stage_opamp_dummy_magic_0.VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_0.VD3.t0 VDDA.t18 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X660 two_stage_opamp_dummy_magic_0.VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VDDA.t460 two_stage_opamp_dummy_magic_0.Y.t48 two_stage_opamp_dummy_magic_0.VOUT+.t10 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X662 two_stage_opamp_dummy_magic_0.VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 two_stage_opamp_dummy_magic_0.VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 two_stage_opamp_dummy_magic_0.VD2.t9 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.V_p.t1 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X665 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t370 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X666 VDDA.t455 two_stage_opamp_dummy_magic_0.Y.t49 two_stage_opamp_dummy_magic_0.VOUT+.t9 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X667 GNDA.t302 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X668 two_stage_opamp_dummy_magic_0.VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 a_14520_5738.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t96 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X670 GNDA.t292 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA.t291 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X671 bgr_0.Vin+.t4 bgr_0.V_TOP.t43 VDDA.t222 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X672 bgr_0.V_p_2.t8 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t8 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X673 two_stage_opamp_dummy_magic_0.VOUT-.t10 GNDA.t128 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X674 two_stage_opamp_dummy_magic_0.V_err_gate.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X675 bgr_0.V_p_1.t2 bgr_0.Vin-.t12 bgr_0.V_mir1.t1 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X676 VDDA.t17 VDDA.t15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X677 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X678 two_stage_opamp_dummy_magic_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t23 GNDA.t337 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X679 a_29700_9260.t1 bgr_0.V_CUR_REF_REG.t2 GNDA.t255 sky130_fd_pr__res_xhigh_po_0p35 l=6
X680 two_stage_opamp_dummy_magic_0.V_p.t40 two_stage_opamp_dummy_magic_0.Vb1.t2 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X681 VDDA.t426 two_stage_opamp_dummy_magic_0.X.t51 two_stage_opamp_dummy_magic_0.VOUT-.t17 VDDA.t425 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X682 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_0.Y.t50 VDDA.t328 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X683 two_stage_opamp_dummy_magic_0.VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 bgr_0.V_TOP.t0 VDDA.t12 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X685 two_stage_opamp_dummy_magic_0.VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 two_stage_opamp_dummy_magic_0.VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 two_stage_opamp_dummy_magic_0.VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 two_stage_opamp_dummy_magic_0.VOUT-.t8 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA.t79 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X689 two_stage_opamp_dummy_magic_0.VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VDDA.t263 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X691 VDDA.t346 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t2 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X692 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 two_stage_opamp_dummy_magic_0.Y.t51 GNDA.t30 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X693 two_stage_opamp_dummy_magic_0.VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X695 GNDA.t311 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X696 two_stage_opamp_dummy_magic_0.Vb2.t10 two_stage_opamp_dummy_magic_0.Vb2.t9 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X697 bgr_0.V_TOP.t44 VDDA.t223 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 bgr_0.Vin+.t3 bgr_0.V_TOP.t45 VDDA.t182 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X699 two_stage_opamp_dummy_magic_0.VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X700 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t427 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X701 two_stage_opamp_dummy_magic_0.VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X703 two_stage_opamp_dummy_magic_0.VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t265 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X705 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.Vb3.t27 VDDA.t188 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X706 two_stage_opamp_dummy_magic_0.VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X708 two_stage_opamp_dummy_magic_0.V_p.t11 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t304 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X709 two_stage_opamp_dummy_magic_0.V_err_p.t21 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t8 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X710 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA.t125 GNDA.t127 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X711 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 two_stage_opamp_dummy_magic_0.V_p_mir.t3 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X713 two_stage_opamp_dummy_magic_0.VD1.t1 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t29 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X714 two_stage_opamp_dummy_magic_0.VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 two_stage_opamp_dummy_magic_0.VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 two_stage_opamp_dummy_magic_0.VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 two_stage_opamp_dummy_magic_0.VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 bgr_0.V_p_2.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 bgr_0.V_mir2.t12 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X719 two_stage_opamp_dummy_magic_0.VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 two_stage_opamp_dummy_magic_0.VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VDDA.t133 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t1 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X722 VDDA.t212 two_stage_opamp_dummy_magic_0.Y.t52 two_stage_opamp_dummy_magic_0.VOUT+.t8 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X723 two_stage_opamp_dummy_magic_0.VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 two_stage_opamp_dummy_magic_0.VD1.t0 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.V_p.t28 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X725 GNDA.t69 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X726 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X727 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 bgr_0.NFET_GATE_10uA.t4 bgr_0.PFET_GATE_10uA.t27 VDDA.t383 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X729 two_stage_opamp_dummy_magic_0.VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 two_stage_opamp_dummy_magic_0.VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 bgr_0.V_TOP.t46 VDDA.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 bgr_0.1st_Vout_1.t0 bgr_0.V_mir1.t21 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X733 two_stage_opamp_dummy_magic_0.VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 two_stage_opamp_dummy_magic_0.VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 two_stage_opamp_dummy_magic_0.V_err_gate.t0 VDDA.t9 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X736 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X737 two_stage_opamp_dummy_magic_0.VD3.t30 two_stage_opamp_dummy_magic_0.Vb3.t28 VDDA.t421 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X738 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X739 VDDA.t381 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X740 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X741 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA.t122 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X742 bgr_0.V_TOP.t47 VDDA.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 two_stage_opamp_dummy_magic_0.VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.t2 GNDA.t352 GNDA.t351 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X745 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t453 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X746 two_stage_opamp_dummy_magic_0.VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 two_stage_opamp_dummy_magic_0.VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t463 GNDA.t349 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X749 two_stage_opamp_dummy_magic_0.VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_0.VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 two_stage_opamp_dummy_magic_0.VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VDDA.t8 VDDA.t6 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X753 two_stage_opamp_dummy_magic_0.VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 bgr_0.PFET_GATE_10uA.t29 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X755 VDDA.t135 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t0 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X756 two_stage_opamp_dummy_magic_0.VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 two_stage_opamp_dummy_magic_0.VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 two_stage_opamp_dummy_magic_0.VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VDDA.t165 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X760 two_stage_opamp_dummy_magic_0.VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X762 GNDA.t325 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X763 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 two_stage_opamp_dummy_magic_0.VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 two_stage_opamp_dummy_magic_0.VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 two_stage_opamp_dummy_magic_0.VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 bgr_0.1st_Vout_1.t5 bgr_0.V_mir1.t22 VDDA.t432 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X768 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t53 VDDA.t428 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X769 two_stage_opamp_dummy_magic_0.VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD1.t12 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X771 bgr_0.V_TOP.t48 VDDA.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t167 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X773 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.X.t22 two_stage_opamp_dummy_magic_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X774 two_stage_opamp_dummy_magic_0.VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t71 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X776 two_stage_opamp_dummy_magic_0.VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 two_stage_opamp_dummy_magic_0.VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 two_stage_opamp_dummy_magic_0.VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X780 two_stage_opamp_dummy_magic_0.V_err_p.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t7 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t252 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X782 two_stage_opamp_dummy_magic_0.VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t119 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X784 two_stage_opamp_dummy_magic_0.VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 GNDA.t340 VDDA.t472 bgr_0.V_p_2.t0 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X786 two_stage_opamp_dummy_magic_0.VD2.t6 two_stage_opamp_dummy_magic_0.VIN+ two_stage_opamp_dummy_magic_0.V_p.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X787 VDDA.t241 bgr_0.V_TOP.t49 bgr_0.Vin+.t2 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X788 VDDA.t5 VDDA.t3 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X789 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 two_stage_opamp_dummy_magic_0.VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 a_14640_5738.t0 a_14640_5738.t1 169.905
R1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 122.474
R10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 39.4005
R12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 39.4005
R13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 39.4005
R14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 39.4005
R16 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 32.2193
R17 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 19.7005
R18 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 19.7005
R19 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R20 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R22 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R24 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 19.7005
R25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R27 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 6.5005
R28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.1255
R29 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R30 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R32 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R33 GNDA.n1738 GNDA.n50 299369
R34 GNDA.n2487 GNDA.n41 68623.1
R35 GNDA.n1737 GNDA.n50 64900
R36 GNDA.n42 GNDA.n41 56607.7
R37 GNDA.n2452 GNDA.n2248 41223.8
R38 GNDA.n2488 GNDA.n40 35590.8
R39 GNDA.n2487 GNDA.n2486 33365.6
R40 GNDA.n2489 GNDA.n37 32661.5
R41 GNDA.n2489 GNDA.n38 32661.5
R42 GNDA.n1741 GNDA.n1740 30676.6
R43 GNDA.n1742 GNDA.n73 29091.6
R44 GNDA.n2465 GNDA.n2248 28430.8
R45 GNDA.n2319 GNDA.n2310 28430.8
R46 GNDA.n2488 GNDA.n39 28372.4
R47 GNDA.n1738 GNDA.n73 26648.4
R48 GNDA.n2490 GNDA.n2489 19630.8
R49 GNDA.n2489 GNDA.n2488 19630.8
R50 GNDA.n1742 GNDA.n1741 18723.2
R51 GNDA.n2483 GNDA.n41 18063.2
R52 GNDA.n1739 GNDA.n1737 17370.4
R53 GNDA.n2484 GNDA.n2483 15462.2
R54 GNDA.n39 GNDA.n37 14773.1
R55 GNDA.n2355 GNDA.n38 14314.3
R56 GNDA.n2486 GNDA.n42 13940.6
R57 GNDA.n2200 GNDA.n71 12361.8
R58 GNDA.n2200 GNDA.n72 12312.5
R59 GNDA.n2198 GNDA.n71 11918.5
R60 GNDA.n2198 GNDA.n72 11869.2
R61 GNDA.n1741 GNDA.n1735 11338.5
R62 GNDA.n1739 GNDA.n1738 11169.2
R63 GNDA.n2491 GNDA.n23 10835
R64 GNDA.n2491 GNDA.n24 10835
R65 GNDA.n36 GNDA.n23 10835
R66 GNDA.n36 GNDA.n24 10835
R67 GNDA.n1740 GNDA.n1739 10831.8
R68 GNDA.n2199 GNDA.n73 10371.4
R69 GNDA.n2431 GNDA.n2310 10371.4
R70 GNDA.n2488 GNDA.n2487 9476.92
R71 GNDA.n2281 GNDA.n7 9308.25
R72 GNDA.n2495 GNDA.n7 9308.25
R73 GNDA.n2281 GNDA.n8 9308.25
R74 GNDA.n2495 GNDA.n8 9308.25
R75 GNDA.n2434 GNDA.n2272 9259
R76 GNDA.n2434 GNDA.n2306 8914.25
R77 GNDA.n2484 GNDA.n42 8800
R78 GNDA.n2440 GNDA.n2272 8175.5
R79 GNDA.n1745 GNDA.n357 8175.5
R80 GNDA.n1745 GNDA.n358 8126.25
R81 GNDA.n2181 GNDA.n55 7880
R82 GNDA.n2238 GNDA.n55 7880
R83 GNDA.n2161 GNDA.n91 7880
R84 GNDA.n2163 GNDA.n91 7880
R85 GNDA.n2181 GNDA.n54 7830.75
R86 GNDA.n2238 GNDA.n54 7830.75
R87 GNDA.n2170 GNDA.n2161 7830.75
R88 GNDA.n2170 GNDA.n2163 7830.75
R89 GNDA.n2440 GNDA.n2306 7830.75
R90 GNDA.n2457 GNDA.n2264 7732.25
R91 GNDA.n2457 GNDA.n2265 7732.25
R92 GNDA.n2266 GNDA.n2264 7732.25
R93 GNDA.n2266 GNDA.n2265 7732.25
R94 GNDA.n2429 GNDA.n2312 7732.25
R95 GNDA.n2372 GNDA.n2312 7732.25
R96 GNDA.n2372 GNDA.n2313 7732.25
R97 GNDA.n2429 GNDA.n2313 7732.25
R98 GNDA.n1749 GNDA.n357 7732.25
R99 GNDA.n1749 GNDA.n358 7683
R100 GNDA.n2473 GNDA.n49 7338.25
R101 GNDA.n2363 GNDA.n2335 7338.25
R102 GNDA.n2363 GNDA.n2336 7289
R103 GNDA.n1740 GNDA.n1736 7287.5
R104 GNDA.n2473 GNDA.n48 7092
R105 GNDA.n2486 GNDA.n2485 6997.35
R106 GNDA.n1334 GNDA.n1327 6845.75
R107 GNDA.n1334 GNDA.n1328 6845.75
R108 GNDA.n1327 GNDA.n1141 6796.5
R109 GNDA.n1328 GNDA.n1141 6796.5
R110 GNDA.n1143 GNDA.n348 6698
R111 GNDA.n1759 GNDA.n348 6698
R112 GNDA.n1143 GNDA.n344 6648.75
R113 GNDA.n1759 GNDA.n344 6648.75
R114 GNDA.n2462 GNDA.n2250 6057.75
R115 GNDA.n2454 GNDA.n2250 6057.75
R116 GNDA.n2462 GNDA.n2251 6057.75
R117 GNDA.n2454 GNDA.n2251 6057.75
R118 GNDA.n2328 GNDA.n2320 6057.75
R119 GNDA.n2369 GNDA.n2320 6057.75
R120 GNDA.n2328 GNDA.n2322 6057.75
R121 GNDA.n2369 GNDA.n2322 6057.75
R122 GNDA.n2356 GNDA.n2355 5574.02
R123 GNDA.n1737 GNDA.n1736 5525.52
R124 GNDA.n1743 GNDA.n1735 5325.97
R125 GNDA.n2242 GNDA.n49 5319
R126 GNDA.n2365 GNDA.n2335 5319
R127 GNDA.n2242 GNDA.n48 5269.75
R128 GNDA.n2365 GNDA.n2336 5269.75
R129 GNDA.n2466 GNDA.n2244 5171.25
R130 GNDA.n2346 GNDA.n2341 5171.25
R131 GNDA.n2470 GNDA.n2244 5122
R132 GNDA.n2350 GNDA.n2341 5122
R133 GNDA.n85 GNDA.n84 4974.25
R134 GNDA.n2173 GNDA.n84 4974.25
R135 GNDA.n2466 GNDA.n2245 4944.7
R136 GNDA.n2346 GNDA.n2344 4944.7
R137 GNDA.n2285 GNDA.n2273 4925
R138 GNDA.n2299 GNDA.n2273 4925
R139 GNDA.n2470 GNDA.n2245 4895.45
R140 GNDA.n2350 GNDA.n2344 4895.45
R141 GNDA.n2285 GNDA.n2275 4728
R142 GNDA.n2299 GNDA.n2275 4728
R143 GNDA.n2482 GNDA.n39 4727.03
R144 GNDA.n764 GNDA.n560 4678.75
R145 GNDA.n760 GNDA.n560 4629.5
R146 GNDA.n764 GNDA.n561 4629.5
R147 GNDA.n1341 GNDA.n1132 4580.25
R148 GNDA.n1341 GNDA.n1133 4580.25
R149 GNDA.n760 GNDA.n561 4580.25
R150 GNDA.n1337 GNDA.n1131 4580.25
R151 GNDA.n1140 GNDA.n1131 4580.25
R152 GNDA.n2172 GNDA.n85 4531
R153 GNDA.n2173 GNDA.n2172 4531
R154 GNDA.n75 GNDA.n74 4531
R155 GNDA.n76 GNDA.n74 4531
R156 GNDA.n2196 GNDA.n75 4531
R157 GNDA.n2196 GNDA.n76 4531
R158 GNDA.n1162 GNDA.n1132 4481.75
R159 GNDA.n1162 GNDA.n1133 4481.75
R160 GNDA.n1337 GNDA.n1137 4481.75
R161 GNDA.n1140 GNDA.n1137 4481.75
R162 GNDA.n1743 GNDA.n1742 3770.78
R163 GNDA.n2449 GNDA.n2267 3595.25
R164 GNDA.n2443 GNDA.n2267 3595.25
R165 GNDA.n2498 GNDA.n5 3349
R166 GNDA.n2303 GNDA.n5 3299.75
R167 GNDA.n2449 GNDA.n2268 3250.5
R168 GNDA.n2443 GNDA.n2268 3250.5
R169 GNDA.n2498 GNDA.n6 3250.5
R170 GNDA.n2303 GNDA.n6 3201.25
R171 GNDA.n2485 GNDA.n2484 3174.4
R172 GNDA.n2310 GNDA.n38 2933.33
R173 GNDA.n2248 GNDA.n37 2933.33
R174 GNDA.n1736 GNDA.n1735 2569.8
R175 GNDA.n2240 GNDA.n2239 2403.7
R176 GNDA.n67 GNDA.n65 2371.15
R177 GNDA.n2206 GNDA.n65 2371.15
R178 GNDA.n51 GNDA.n44 2326.02
R179 GNDA.n2480 GNDA.n44 2326.02
R180 GNDA.n2354 GNDA.n2339 2326.02
R181 GNDA.n2358 GNDA.n2354 2326.02
R182 GNDA.n2240 GNDA.n50 2305.25
R183 GNDA.n2209 GNDA.n64 2142.38
R184 GNDA.n2156 GNDA.n83 2142.38
R185 GNDA.n2189 GNDA.n64 1846.88
R186 GNDA.n2177 GNDA.n83 1846.88
R187 GNDA.n2240 GNDA.n52 1775.62
R188 GNDA.n2241 GNDA.n2240 1532.48
R189 GNDA.n66 GNDA.n65 1301.55
R190 GNDA.n2477 GNDA.n44 1114.8
R191 GNDA.n2354 GNDA.n2353 1114.8
R192 GNDA.n2185 GNDA.n64 991.841
R193 GNDA.n89 GNDA.n83 991.841
R194 GNDA.n1695 GNDA.n384 949.682
R195 GNDA.n1782 GNDA.t137 949.682
R196 GNDA.n2201 GNDA.n69 803.201
R197 GNDA.n2201 GNDA.n70 800
R198 GNDA.n2197 GNDA.n69 774.4
R199 GNDA.n2197 GNDA.n70 771.201
R200 GNDA.n2323 GNDA.t153 734.418
R201 GNDA.n2325 GNDA.t141 734.418
R202 GNDA.n2256 GNDA.t167 734.418
R203 GNDA.n2252 GNDA.t150 734.418
R204 GNDA.n35 GNDA.n29 704
R205 GNDA.n35 GNDA.n34 697.601
R206 GNDA.n2309 GNDA.t171 682.201
R207 GNDA.n2271 GNDA.t125 682.201
R208 GNDA.n1765 GNDA.n336 669.307
R209 GNDA.n2308 GNDA.t205 666.134
R210 GNDA.n2270 GNDA.t138 666.134
R211 GNDA.n2160 GNDA.n2152 627.408
R212 GNDA.n2483 GNDA.n2482 624.324
R213 GNDA.n1707 GNDA.n1695 623.755
R214 GNDA.n1788 GNDA.t137 623.755
R215 GNDA.n2359 GNDA.n2338 617.601
R216 GNDA.n2479 GNDA.n45 617.601
R217 GNDA.n2493 GNDA.n18 604.801
R218 GNDA.n2494 GNDA.n2493 604.801
R219 GNDA.n2435 GNDA.n2307 601.601
R220 GNDA.n925 GNDA.n924 585
R221 GNDA.n922 GNDA.n897 585
R222 GNDA.n921 GNDA.n899 585
R223 GNDA.n919 GNDA.n918 585
R224 GNDA.n917 GNDA.n900 585
R225 GNDA.n916 GNDA.n915 585
R226 GNDA.n914 GNDA.n901 585
R227 GNDA.n912 GNDA.n911 585
R228 GNDA.n910 GNDA.n903 585
R229 GNDA.n909 GNDA.n908 585
R230 GNDA.n907 GNDA.n904 585
R231 GNDA.n210 GNDA.n208 585
R232 GNDA.n722 GNDA.n692 585
R233 GNDA.n721 GNDA.n720 585
R234 GNDA.n719 GNDA.n694 585
R235 GNDA.n717 GNDA.n716 585
R236 GNDA.n715 GNDA.n696 585
R237 GNDA.n714 GNDA.n713 585
R238 GNDA.n712 GNDA.n697 585
R239 GNDA.n710 GNDA.n709 585
R240 GNDA.n708 GNDA.n699 585
R241 GNDA.n707 GNDA.n706 585
R242 GNDA.n705 GNDA.n700 585
R243 GNDA.n703 GNDA.n702 585
R244 GNDA.n2150 GNDA.n2149 585
R245 GNDA.n2151 GNDA.n2150 585
R246 GNDA.n2115 GNDA.n2114 585
R247 GNDA.n2118 GNDA.n2117 585
R248 GNDA.n2120 GNDA.n2119 585
R249 GNDA.n2124 GNDA.n2123 585
R250 GNDA.n2122 GNDA.n115 585
R251 GNDA.n2131 GNDA.n2130 585
R252 GNDA.n2133 GNDA.n2132 585
R253 GNDA.n2137 GNDA.n2136 585
R254 GNDA.n2135 GNDA.n111 585
R255 GNDA.n2144 GNDA.n2143 585
R256 GNDA.n2146 GNDA.n2145 585
R257 GNDA.n2148 GNDA.n106 585
R258 GNDA.n1684 GNDA.n1683 585
R259 GNDA.n1588 GNDA.n99 585
R260 GNDA.n2151 GNDA.n99 585
R261 GNDA.n456 GNDA.n455 585
R262 GNDA.n1660 GNDA.n1659 585
R263 GNDA.n1662 GNDA.n1661 585
R264 GNDA.n453 GNDA.n452 585
R265 GNDA.n451 GNDA.n447 585
R266 GNDA.n1670 GNDA.n1669 585
R267 GNDA.n1672 GNDA.n1671 585
R268 GNDA.n445 GNDA.n444 585
R269 GNDA.n443 GNDA.n439 585
R270 GNDA.n1680 GNDA.n1679 585
R271 GNDA.n1682 GNDA.n1681 585
R272 GNDA.n834 GNDA.n833 585
R273 GNDA.n833 GNDA.n832 585
R274 GNDA.n524 GNDA.n520 585
R275 GNDA.n831 GNDA.n520 585
R276 GNDA.n829 GNDA.n828 585
R277 GNDA.n830 GNDA.n829 585
R278 GNDA.n537 GNDA.n522 585
R279 GNDA.n522 GNDA.n521 585
R280 GNDA.n536 GNDA.n535 585
R281 GNDA.n535 GNDA.n534 585
R282 GNDA.n533 GNDA.n532 585
R283 GNDA.n533 GNDA.n374 585
R284 GNDA.n527 GNDA.n370 585
R285 GNDA.n1723 GNDA.n370 585
R286 GNDA.n1726 GNDA.n1725 585
R287 GNDA.n1725 GNDA.n1724 585
R288 GNDA.n366 GNDA.n364 585
R289 GNDA.n364 GNDA.n362 585
R290 GNDA.n1733 GNDA.n1732 585
R291 GNDA.n1734 GNDA.n1733 585
R292 GNDA.n771 GNDA.n363 585
R293 GNDA.n363 GNDA.n361 585
R294 GNDA.n770 GNDA.n769 585
R295 GNDA.n769 GNDA.n768 585
R296 GNDA.n1948 GNDA.n1947 585
R297 GNDA.n1949 GNDA.n283 585
R298 GNDA.n1950 GNDA.n282 585
R299 GNDA.n279 GNDA.n278 585
R300 GNDA.n1955 GNDA.n277 585
R301 GNDA.n1956 GNDA.n276 585
R302 GNDA.n1957 GNDA.n275 585
R303 GNDA.n271 GNDA.n269 585
R304 GNDA.n1963 GNDA.n1962 585
R305 GNDA.n270 GNDA.n268 585
R306 GNDA.n1965 GNDA.n107 585
R307 GNDA.n1585 GNDA.n462 585
R308 GNDA.n461 GNDA.n460 585
R309 GNDA.n1579 GNDA.n1578 585
R310 GNDA.n1577 GNDA.n1576 585
R311 GNDA.n1575 GNDA.n466 585
R312 GNDA.n465 GNDA.n464 585
R313 GNDA.n1569 GNDA.n1568 585
R314 GNDA.n1567 GNDA.n1566 585
R315 GNDA.n1565 GNDA.n469 585
R316 GNDA.n468 GNDA.n257 585
R317 GNDA.n1965 GNDA.n257 585
R318 GNDA.n472 GNDA.n470 585
R319 GNDA.n472 GNDA.n204 585
R320 GNDA.n1948 GNDA.n285 585
R321 GNDA.n1949 GNDA.n281 585
R322 GNDA.n1951 GNDA.n1950 585
R323 GNDA.n1953 GNDA.n279 585
R324 GNDA.n1955 GNDA.n1954 585
R325 GNDA.n1956 GNDA.n274 585
R326 GNDA.n1958 GNDA.n1957 585
R327 GNDA.n1960 GNDA.n271 585
R328 GNDA.n1962 GNDA.n1961 585
R329 GNDA.n329 GNDA.n270 585
R330 GNDA.n458 GNDA.n273 585
R331 GNDA.n1585 GNDA.n1584 585
R332 GNDA.n1582 GNDA.n460 585
R333 GNDA.n1580 GNDA.n1579 585
R334 GNDA.n1576 GNDA.n463 585
R335 GNDA.n1575 GNDA.n1574 585
R336 GNDA.n1572 GNDA.n464 585
R337 GNDA.n1570 GNDA.n1569 585
R338 GNDA.n1566 GNDA.n467 585
R339 GNDA.n1565 GNDA.n1564 585
R340 GNDA.n1562 GNDA.n468 585
R341 GNDA.n1562 GNDA.n273 585
R342 GNDA.n1432 GNDA.n250 585
R343 GNDA.n1431 GNDA.n889 585
R344 GNDA.n888 GNDA.n887 585
R345 GNDA.n1426 GNDA.n1425 585
R346 GNDA.n1424 GNDA.n1423 585
R347 GNDA.n1422 GNDA.n893 585
R348 GNDA.n892 GNDA.n891 585
R349 GNDA.n1416 GNDA.n1415 585
R350 GNDA.n1414 GNDA.n1413 585
R351 GNDA.n1412 GNDA.n896 585
R352 GNDA.n898 GNDA.n895 585
R353 GNDA.n898 GNDA.n204 585
R354 GNDA.n1433 GNDA.n1432 585
R355 GNDA.n1431 GNDA.n1430 585
R356 GNDA.n1429 GNDA.n887 585
R357 GNDA.n1427 GNDA.n1426 585
R358 GNDA.n1423 GNDA.n890 585
R359 GNDA.n1422 GNDA.n1421 585
R360 GNDA.n1419 GNDA.n891 585
R361 GNDA.n1417 GNDA.n1416 585
R362 GNDA.n1413 GNDA.n894 585
R363 GNDA.n1412 GNDA.n1411 585
R364 GNDA.n1388 GNDA.n1387 585
R365 GNDA.n1389 GNDA.n933 585
R366 GNDA.n1391 GNDA.n1390 585
R367 GNDA.n1393 GNDA.n932 585
R368 GNDA.n1396 GNDA.n1395 585
R369 GNDA.n1397 GNDA.n931 585
R370 GNDA.n1399 GNDA.n1398 585
R371 GNDA.n1401 GNDA.n930 585
R372 GNDA.n1404 GNDA.n1403 585
R373 GNDA.n1405 GNDA.n929 585
R374 GNDA.n1407 GNDA.n1406 585
R375 GNDA.n1409 GNDA.n927 585
R376 GNDA.n1540 GNDA.n1539 585
R377 GNDA.n1541 GNDA.n509 585
R378 GNDA.n1543 GNDA.n1542 585
R379 GNDA.n1545 GNDA.n508 585
R380 GNDA.n1548 GNDA.n1547 585
R381 GNDA.n1549 GNDA.n507 585
R382 GNDA.n1551 GNDA.n1550 585
R383 GNDA.n1553 GNDA.n506 585
R384 GNDA.n1556 GNDA.n1555 585
R385 GNDA.n1557 GNDA.n505 585
R386 GNDA.n1559 GNDA.n1558 585
R387 GNDA.n1561 GNDA.n503 585
R388 GNDA.n1686 GNDA.n1685 585
R389 GNDA.n838 GNDA.n518 585
R390 GNDA.n841 GNDA.n517 585
R391 GNDA.n842 GNDA.n516 585
R392 GNDA.n845 GNDA.n515 585
R393 GNDA.n846 GNDA.n514 585
R394 GNDA.n849 GNDA.n513 585
R395 GNDA.n850 GNDA.n512 585
R396 GNDA.n853 GNDA.n511 585
R397 GNDA.n855 GNDA.n510 585
R398 GNDA.n856 GNDA.n430 585
R399 GNDA.n1686 GNDA.n430 585
R400 GNDA.n1537 GNDA.n857 585
R401 GNDA.n1537 GNDA.n1536 585
R402 GNDA.n1694 GNDA.n403 585
R403 GNDA.n839 GNDA.n838 585
R404 GNDA.n841 GNDA.n840 585
R405 GNDA.n843 GNDA.n842 585
R406 GNDA.n845 GNDA.n844 585
R407 GNDA.n847 GNDA.n846 585
R408 GNDA.n849 GNDA.n848 585
R409 GNDA.n851 GNDA.n850 585
R410 GNDA.n853 GNDA.n852 585
R411 GNDA.n855 GNDA.n854 585
R412 GNDA.n856 GNDA.n409 585
R413 GNDA.n1694 GNDA.n409 585
R414 GNDA.n1089 GNDA.n959 585
R415 GNDA.n957 GNDA.n954 585
R416 GNDA.n953 GNDA.n952 585
R417 GNDA.n951 GNDA.n948 585
R418 GNDA.n947 GNDA.n946 585
R419 GNDA.n945 GNDA.n942 585
R420 GNDA.n941 GNDA.n940 585
R421 GNDA.n939 GNDA.n936 585
R422 GNDA.n935 GNDA.n934 585
R423 GNDA.n389 GNDA.n387 585
R424 GNDA.n959 GNDA.n958 585
R425 GNDA.n957 GNDA.n956 585
R426 GNDA.n955 GNDA.n952 585
R427 GNDA.n951 GNDA.n950 585
R428 GNDA.n949 GNDA.n946 585
R429 GNDA.n945 GNDA.n944 585
R430 GNDA.n943 GNDA.n940 585
R431 GNDA.n939 GNDA.n938 585
R432 GNDA.n937 GNDA.n934 585
R433 GNDA.n397 GNDA.n387 585
R434 GNDA.n1945 GNDA.n287 585
R435 GNDA.n1946 GNDA.n1945 585
R436 GNDA.n1944 GNDA.n1943 585
R437 GNDA.n1943 GNDA.n204 585
R438 GNDA.n1846 GNDA.n1845 585
R439 GNDA.n309 GNDA.n308 585
R440 GNDA.n1918 GNDA.n1917 585
R441 GNDA.n1921 GNDA.n1920 585
R442 GNDA.n307 GNDA.n304 585
R443 GNDA.n300 GNDA.n299 585
R444 GNDA.n1929 GNDA.n1928 585
R445 GNDA.n1932 GNDA.n1931 585
R446 GNDA.n298 GNDA.n295 585
R447 GNDA.n291 GNDA.n289 585
R448 GNDA.n1940 GNDA.n1939 585
R449 GNDA.n1942 GNDA.n288 585
R450 GNDA.n1091 GNDA.n960 585
R451 GNDA.n1091 GNDA.n1090 585
R452 GNDA.n1088 GNDA.n859 585
R453 GNDA.n1536 GNDA.n859 585
R454 GNDA.n990 GNDA.n989 585
R455 GNDA.n982 GNDA.n981 585
R456 GNDA.n1062 GNDA.n1061 585
R457 GNDA.n1065 GNDA.n1064 585
R458 GNDA.n980 GNDA.n977 585
R459 GNDA.n973 GNDA.n972 585
R460 GNDA.n1073 GNDA.n1072 585
R461 GNDA.n1076 GNDA.n1075 585
R462 GNDA.n971 GNDA.n968 585
R463 GNDA.n964 GNDA.n963 585
R464 GNDA.n1084 GNDA.n1083 585
R465 GNDA.n1087 GNDA.n1086 585
R466 GNDA.n988 GNDA.n273 585
R467 GNDA.n986 GNDA.n273 585
R468 GNDA.n1200 GNDA.n1199 585
R469 GNDA.n1194 GNDA.n1193 585
R470 GNDA.n1272 GNDA.n1271 585
R471 GNDA.n1275 GNDA.n1274 585
R472 GNDA.n1192 GNDA.n1189 585
R473 GNDA.n1185 GNDA.n1184 585
R474 GNDA.n1283 GNDA.n1282 585
R475 GNDA.n1286 GNDA.n1285 585
R476 GNDA.n1183 GNDA.n1179 585
R477 GNDA.n1293 GNDA.n1292 585
R478 GNDA.n1295 GNDA.n1294 585
R479 GNDA.n1298 GNDA.n1297 585
R480 GNDA.n1694 GNDA.n396 585
R481 GNDA.n1694 GNDA.n410 585
R482 GNDA.n417 GNDA.n414 585
R483 GNDA.n1104 GNDA.n1103 585
R484 GNDA.n1107 GNDA.n1102 585
R485 GNDA.n1108 GNDA.n1101 585
R486 GNDA.n1111 GNDA.n1100 585
R487 GNDA.n1112 GNDA.n1099 585
R488 GNDA.n1115 GNDA.n1098 585
R489 GNDA.n1116 GNDA.n1097 585
R490 GNDA.n1119 GNDA.n1096 585
R491 GNDA.n1120 GNDA.n1095 585
R492 GNDA.n1093 GNDA.n858 585
R493 GNDA.n1536 GNDA.n858 585
R494 GNDA.n414 GNDA.n411 585
R495 GNDA.n1105 GNDA.n1104 585
R496 GNDA.n1107 GNDA.n1106 585
R497 GNDA.n1109 GNDA.n1108 585
R498 GNDA.n1111 GNDA.n1110 585
R499 GNDA.n1113 GNDA.n1112 585
R500 GNDA.n1115 GNDA.n1114 585
R501 GNDA.n1117 GNDA.n1116 585
R502 GNDA.n1119 GNDA.n1118 585
R503 GNDA.n1121 GNDA.n1120 585
R504 GNDA.n1362 GNDA.n1361 585
R505 GNDA.n1364 GNDA.n1126 585
R506 GNDA.n1367 GNDA.n1366 585
R507 GNDA.n1368 GNDA.n1125 585
R508 GNDA.n1370 GNDA.n1369 585
R509 GNDA.n1372 GNDA.n1124 585
R510 GNDA.n1375 GNDA.n1374 585
R511 GNDA.n1376 GNDA.n1123 585
R512 GNDA.n1378 GNDA.n1377 585
R513 GNDA.n1380 GNDA.n1122 585
R514 GNDA.n1381 GNDA.n1094 585
R515 GNDA.n1384 GNDA.n1383 585
R516 GNDA.n1968 GNDA.n249 585
R517 GNDA.n1968 GNDA.n1967 585
R518 GNDA.n1969 GNDA.n247 585
R519 GNDA.n247 GNDA.n204 585
R520 GNDA.n1689 GNDA.n415 585
R521 GNDA.n1689 GNDA.n1688 585
R522 GNDA.n1535 GNDA.n416 585
R523 GNDA.n1536 GNDA.n1535 585
R524 GNDA.n1438 GNDA.n1437 585
R525 GNDA.n882 GNDA.n881 585
R526 GNDA.n1510 GNDA.n1509 585
R527 GNDA.n1513 GNDA.n1512 585
R528 GNDA.n880 GNDA.n877 585
R529 GNDA.n873 GNDA.n872 585
R530 GNDA.n1521 GNDA.n1520 585
R531 GNDA.n1524 GNDA.n1523 585
R532 GNDA.n871 GNDA.n868 585
R533 GNDA.n864 GNDA.n862 585
R534 GNDA.n1532 GNDA.n1531 585
R535 GNDA.n1534 GNDA.n860 585
R536 GNDA.n1436 GNDA.n273 585
R537 GNDA.n1434 GNDA.n273 585
R538 GNDA.n587 GNDA.n412 585
R539 GNDA.n590 GNDA.n589 585
R540 GNDA.n663 GNDA.n662 585
R541 GNDA.n666 GNDA.n665 585
R542 GNDA.n586 GNDA.n583 585
R543 GNDA.n579 GNDA.n578 585
R544 GNDA.n674 GNDA.n673 585
R545 GNDA.n677 GNDA.n676 585
R546 GNDA.n577 GNDA.n574 585
R547 GNDA.n570 GNDA.n568 585
R548 GNDA.n685 GNDA.n684 585
R549 GNDA.n687 GNDA.n567 585
R550 GNDA.n1694 GNDA.n390 585
R551 GNDA.n1694 GNDA.n1693 585
R552 GNDA.n2065 GNDA.n219 585
R553 GNDA.n2063 GNDA.n2062 585
R554 GNDA.n2035 GNDA.n222 585
R555 GNDA.n2034 GNDA.n2030 585
R556 GNDA.n2041 GNDA.n2040 585
R557 GNDA.n2043 GNDA.n2028 585
R558 GNDA.n2045 GNDA.n2044 585
R559 GNDA.n2025 GNDA.n2024 585
R560 GNDA.n2051 GNDA.n2050 585
R561 GNDA.n2054 GNDA.n2053 585
R562 GNDA.n2023 GNDA.n245 585
R563 GNDA.n2021 GNDA.n2020 585
R564 GNDA.n501 GNDA.n500 585
R565 GNDA.n498 GNDA.n471 585
R566 GNDA.n497 GNDA.n496 585
R567 GNDA.n495 GNDA.n494 585
R568 GNDA.n493 GNDA.n474 585
R569 GNDA.n491 GNDA.n490 585
R570 GNDA.n489 GNDA.n475 585
R571 GNDA.n488 GNDA.n487 585
R572 GNDA.n485 GNDA.n476 585
R573 GNDA.n483 GNDA.n482 585
R574 GNDA.n481 GNDA.n477 585
R575 GNDA.n480 GNDA.n479 585
R576 GNDA.n1844 GNDA.n206 585
R577 GNDA.n1842 GNDA.n1841 585
R578 GNDA.n1836 GNDA.n313 585
R579 GNDA.n1840 GNDA.n313 585
R580 GNDA.n1838 GNDA.n1837 585
R581 GNDA.n1839 GNDA.n1838 585
R582 GNDA.n1835 GNDA.n315 585
R583 GNDA.n315 GNDA.n314 585
R584 GNDA.n1834 GNDA.n1833 585
R585 GNDA.n1833 GNDA.n1832 585
R586 GNDA.n317 GNDA.n316 585
R587 GNDA.n318 GNDA.n317 585
R588 GNDA.n1811 GNDA.n1810 585
R589 GNDA.n1810 GNDA.n1809 585
R590 GNDA.n1812 GNDA.n1808 585
R591 GNDA.n1808 GNDA.n1807 585
R592 GNDA.n1814 GNDA.n1813 585
R593 GNDA.n1815 GNDA.n1814 585
R594 GNDA.n1806 GNDA.n1805 585
R595 GNDA.n1816 GNDA.n1806 585
R596 GNDA.n1819 GNDA.n1818 585
R597 GNDA.n1818 GNDA.n1817 585
R598 GNDA.n2066 GNDA.n201 585
R599 GNDA.n221 GNDA.n220 585
R600 GNDA.n2069 GNDA.n218 585
R601 GNDA.n218 GNDA.n217 585
R602 GNDA.n2071 GNDA.n2070 585
R603 GNDA.n2072 GNDA.n2071 585
R604 GNDA.n216 GNDA.n215 585
R605 GNDA.n2073 GNDA.n216 585
R606 GNDA.n2076 GNDA.n2075 585
R607 GNDA.n2075 GNDA.n2074 585
R608 GNDA.n2077 GNDA.n214 585
R609 GNDA.n214 GNDA.n213 585
R610 GNDA.n2079 GNDA.n2078 585
R611 GNDA.n2080 GNDA.n2079 585
R612 GNDA.n212 GNDA.n211 585
R613 GNDA.n2081 GNDA.n212 585
R614 GNDA.n2084 GNDA.n2083 585
R615 GNDA.n2083 GNDA.n2082 585
R616 GNDA.n2085 GNDA.n209 585
R617 GNDA.n209 GNDA.n207 585
R618 GNDA.n2087 GNDA.n2086 585
R619 GNDA.n2088 GNDA.n2087 585
R620 GNDA.n2113 GNDA.n2112 585
R621 GNDA.n2111 GNDA.n2110 585
R622 GNDA.n2109 GNDA.n2108 585
R623 GNDA.n2109 GNDA.n191 585
R624 GNDA.n2107 GNDA.n192 585
R625 GNDA.n2103 GNDA.n192 585
R626 GNDA.n2106 GNDA.n2105 585
R627 GNDA.n2105 GNDA.n2104 585
R628 GNDA.n2101 GNDA.n193 585
R629 GNDA.n2102 GNDA.n2101 585
R630 GNDA.n2100 GNDA.n195 585
R631 GNDA.n2100 GNDA.n2099 585
R632 GNDA.n2094 GNDA.n194 585
R633 GNDA.n2098 GNDA.n194 585
R634 GNDA.n2096 GNDA.n2095 585
R635 GNDA.n2097 GNDA.n2096 585
R636 GNDA.n2093 GNDA.n197 585
R637 GNDA.n197 GNDA.n196 585
R638 GNDA.n2092 GNDA.n2091 585
R639 GNDA.n2091 GNDA.n2090 585
R640 GNDA.n199 GNDA.n198 585
R641 GNDA.n2089 GNDA.n199 585
R642 GNDA.n1787 GNDA.n1786 585
R643 GNDA.n1788 GNDA.n1787 585
R644 GNDA.n1791 GNDA.n1790 585
R645 GNDA.n1790 GNDA.n1789 585
R646 GNDA.n1792 GNDA.n326 585
R647 GNDA.n326 GNDA.n325 585
R648 GNDA.n1794 GNDA.n1793 585
R649 GNDA.n1795 GNDA.n1794 585
R650 GNDA.n324 GNDA.n323 585
R651 GNDA.n1796 GNDA.n324 585
R652 GNDA.n1799 GNDA.n1798 585
R653 GNDA.n1798 GNDA.n1797 585
R654 GNDA.n1800 GNDA.n321 585
R655 GNDA.n321 GNDA.n319 585
R656 GNDA.n1830 GNDA.n1829 585
R657 GNDA.n1831 GNDA.n1830 585
R658 GNDA.n1828 GNDA.n322 585
R659 GNDA.n322 GNDA.n320 585
R660 GNDA.n1827 GNDA.n1826 585
R661 GNDA.n1826 GNDA.n1825 585
R662 GNDA.n1802 GNDA.n1801 585
R663 GNDA.n1824 GNDA.n1802 585
R664 GNDA.n1822 GNDA.n1821 585
R665 GNDA.n1823 GNDA.n1822 585
R666 GNDA.n1820 GNDA.n1804 585
R667 GNDA.n1804 GNDA.n1803 585
R668 GNDA.n1766 GNDA.n337 585
R669 GNDA.n1768 GNDA.n1767 585
R670 GNDA.n1769 GNDA.n1768 585
R671 GNDA.n1709 GNDA.n1708 585
R672 GNDA.n1708 GNDA.n1707 585
R673 GNDA.n388 GNDA.n386 585
R674 GNDA.n1706 GNDA.n388 585
R675 GNDA.n1704 GNDA.n1703 585
R676 GNDA.n1705 GNDA.n1704 585
R677 GNDA.n1702 GNDA.n1697 585
R678 GNDA.n1697 GNDA.n1696 585
R679 GNDA.n1701 GNDA.n1700 585
R680 GNDA.n1700 GNDA.n1699 585
R681 GNDA.n1698 GNDA.n333 585
R682 GNDA.n335 GNDA.n333 585
R683 GNDA.n1771 GNDA.n334 585
R684 GNDA.n1771 GNDA.n1770 585
R685 GNDA.n1772 GNDA.n332 585
R686 GNDA.n1773 GNDA.n1772 585
R687 GNDA.n1776 GNDA.n1775 585
R688 GNDA.n1775 GNDA.n1774 585
R689 GNDA.n1777 GNDA.n331 585
R690 GNDA.n331 GNDA.n330 585
R691 GNDA.n1779 GNDA.n1778 585
R692 GNDA.n1780 GNDA.n1779 585
R693 GNDA.n328 GNDA.n327 585
R694 GNDA.n1781 GNDA.n328 585
R695 GNDA.n1784 GNDA.n1783 585
R696 GNDA.n1783 GNDA.n1782 585
R697 GNDA.n1159 GNDA.n1145 585
R698 GNDA.n1145 GNDA.n1142 585
R699 GNDA.n1158 GNDA.n1157 585
R700 GNDA.n1157 GNDA.n1156 585
R701 GNDA.n1148 GNDA.n1147 585
R702 GNDA.n1155 GNDA.n1148 585
R703 GNDA.n1153 GNDA.n1152 585
R704 GNDA.n1154 GNDA.n1153 585
R705 GNDA.n1151 GNDA.n1150 585
R706 GNDA.n1150 GNDA.n1149 585
R707 GNDA.n381 GNDA.n379 585
R708 GNDA.n379 GNDA.n377 585
R709 GNDA.n1721 GNDA.n1720 585
R710 GNDA.n1722 GNDA.n1721 585
R711 GNDA.n1719 GNDA.n380 585
R712 GNDA.n380 GNDA.n378 585
R713 GNDA.n1718 GNDA.n1717 585
R714 GNDA.n1717 GNDA.n1716 585
R715 GNDA.n383 GNDA.n382 585
R716 GNDA.n1715 GNDA.n383 585
R717 GNDA.n1713 GNDA.n1712 585
R718 GNDA.n1714 GNDA.n1713 585
R719 GNDA.n1711 GNDA.n385 585
R720 GNDA.n385 GNDA.n384 585
R721 GNDA.n1301 GNDA.n1300 585
R722 GNDA.n1303 GNDA.n1302 585
R723 GNDA.n1305 GNDA.n1304 585
R724 GNDA.n1304 GNDA.n1138 585
R725 GNDA.n1306 GNDA.n1169 585
R726 GNDA.n1169 GNDA.n1168 585
R727 GNDA.n1308 GNDA.n1307 585
R728 GNDA.n1309 GNDA.n1308 585
R729 GNDA.n1167 GNDA.n1166 585
R730 GNDA.n1310 GNDA.n1167 585
R731 GNDA.n1313 GNDA.n1312 585
R732 GNDA.n1312 GNDA.n1311 585
R733 GNDA.n1314 GNDA.n1165 585
R734 GNDA.n1165 GNDA.n1164 585
R735 GNDA.n1316 GNDA.n1315 585
R736 GNDA.n1317 GNDA.n1316 585
R737 GNDA.n1161 GNDA.n1160 585
R738 GNDA.n1318 GNDA.n1161 585
R739 GNDA.n1321 GNDA.n1320 585
R740 GNDA.n1320 GNDA.n1319 585
R741 GNDA.n1322 GNDA.n1146 585
R742 GNDA.n1146 GNDA.n1144 585
R743 GNDA.n1324 GNDA.n1323 585
R744 GNDA.n1325 GNDA.n1324 585
R745 GNDA.n1299 GNDA.n1174 585
R746 GNDA.n1299 GNDA.n1173 585
R747 GNDA.n565 GNDA.n563 585
R748 GNDA.n356 GNDA.n354 585
R749 GNDA.n1753 GNDA.n1752 585
R750 GNDA.n1752 GNDA.n1751 585
R751 GNDA.n1754 GNDA.n352 585
R752 GNDA.n355 GNDA.n352 585
R753 GNDA.n1756 GNDA.n1755 585
R754 GNDA.n1757 GNDA.n1756 585
R755 GNDA.n1344 GNDA.n351 585
R756 GNDA.n351 GNDA.n349 585
R757 GNDA.n1346 GNDA.n1345 585
R758 GNDA.n1348 GNDA.n1346 585
R759 GNDA.n1351 GNDA.n1350 585
R760 GNDA.n1350 GNDA.n1349 585
R761 GNDA.n1352 GNDA.n1343 585
R762 GNDA.n1347 GNDA.n1343 585
R763 GNDA.n1354 GNDA.n1353 585
R764 GNDA.n1355 GNDA.n1354 585
R765 GNDA.n1129 GNDA.n1128 585
R766 GNDA.n1356 GNDA.n1129 585
R767 GNDA.n1359 GNDA.n1358 585
R768 GNDA.n1358 GNDA.n1357 585
R769 GNDA.n1360 GNDA.n1127 585
R770 GNDA.n1130 GNDA.n1127 585
R771 GNDA.n688 GNDA.n566 585
R772 GNDA.n689 GNDA.n688 585
R773 GNDA.n559 GNDA.n558 585
R774 GNDA.n735 GNDA.n733 585
R775 GNDA.n738 GNDA.n737 585
R776 GNDA.n737 GNDA.n736 585
R777 GNDA.n739 GNDA.n730 585
R778 GNDA.n734 GNDA.n730 585
R779 GNDA.n741 GNDA.n740 585
R780 GNDA.n742 GNDA.n741 585
R781 GNDA.n728 GNDA.n727 585
R782 GNDA.n743 GNDA.n728 585
R783 GNDA.n746 GNDA.n745 585
R784 GNDA.n745 GNDA.n744 585
R785 GNDA.n747 GNDA.n726 585
R786 GNDA.n726 GNDA.n725 585
R787 GNDA.n749 GNDA.n748 585
R788 GNDA.n750 GNDA.n749 585
R789 GNDA.n724 GNDA.n723 585
R790 GNDA.n751 GNDA.n724 585
R791 GNDA.n754 GNDA.n753 585
R792 GNDA.n753 GNDA.n752 585
R793 GNDA.n755 GNDA.n693 585
R794 GNDA.n693 GNDA.n691 585
R795 GNDA.n757 GNDA.n756 585
R796 GNDA.n758 GNDA.n757 585
R797 GNDA.n767 GNDA.n557 585
R798 GNDA.n767 GNDA.n766 585
R799 GNDA.n2316 GNDA.t128 535.191
R800 GNDA.n2314 GNDA.t144 535.191
R801 GNDA.n2262 GNDA.t193 535.191
R802 GNDA.n2260 GNDA.t199 535.191
R803 GNDA.n2439 GNDA.n2307 531.201
R804 GNDA.n1747 GNDA.n1746 531.201
R805 GNDA.n1746 GNDA.n359 528
R806 GNDA.n2236 GNDA.n57 512
R807 GNDA.n2237 GNDA.n2236 512
R808 GNDA.n2167 GNDA.n2164 512
R809 GNDA.n2168 GNDA.n2167 512
R810 GNDA.n57 GNDA.n56 508.8
R811 GNDA.n2237 GNDA.n56 508.8
R812 GNDA.n2169 GNDA.n2164 508.8
R813 GNDA.n2169 GNDA.n2168 508.8
R814 GNDA.n1156 GNDA.n1142 505.748
R815 GNDA.n1156 GNDA.n1155 505.748
R816 GNDA.n1155 GNDA.n1154 505.748
R817 GNDA.n1154 GNDA.n1149 505.748
R818 GNDA.n1149 GNDA.n377 505.748
R819 GNDA.n1722 GNDA.n378 505.748
R820 GNDA.n1716 GNDA.n378 505.748
R821 GNDA.n1716 GNDA.n1715 505.748
R822 GNDA.n1715 GNDA.n1714 505.748
R823 GNDA.n1714 GNDA.n384 505.748
R824 GNDA.n1707 GNDA.n1706 505.748
R825 GNDA.n1706 GNDA.n1705 505.748
R826 GNDA.n1705 GNDA.n1696 505.748
R827 GNDA.n1699 GNDA.n1696 505.748
R828 GNDA.n1699 GNDA.n335 505.748
R829 GNDA.n1770 GNDA.n335 505.748
R830 GNDA.n1774 GNDA.n1773 505.748
R831 GNDA.n1774 GNDA.n330 505.748
R832 GNDA.n1780 GNDA.n330 505.748
R833 GNDA.n1781 GNDA.n1780 505.748
R834 GNDA.n1782 GNDA.n1781 505.748
R835 GNDA.n1789 GNDA.n1788 505.748
R836 GNDA.n1789 GNDA.n325 505.748
R837 GNDA.n1795 GNDA.n325 505.748
R838 GNDA.n1796 GNDA.n1795 505.748
R839 GNDA.n1797 GNDA.n1796 505.748
R840 GNDA.n1797 GNDA.n319 505.748
R841 GNDA.n1831 GNDA.n320 505.748
R842 GNDA.n1825 GNDA.n320 505.748
R843 GNDA.n1825 GNDA.n1824 505.748
R844 GNDA.n1824 GNDA.n1823 505.748
R845 GNDA.n1823 GNDA.n1803 505.748
R846 GNDA.n2428 GNDA.n2427 502.401
R847 GNDA.n1748 GNDA.n1747 499.2
R848 GNDA.t135 GNDA.n371 496.098
R849 GNDA.n2427 GNDA.n2373 496
R850 GNDA.n2377 GNDA.n2376 496
R851 GNDA.n9 GNDA.t214 493.418
R852 GNDA.n13 GNDA.t176 493.418
R853 GNDA.n12 GNDA.t211 493.418
R854 GNDA.n11 GNDA.t196 493.418
R855 GNDA.n30 GNDA.t217 493.418
R856 GNDA.n31 GNDA.t202 493.418
R857 GNDA.n21 GNDA.t189 493.418
R858 GNDA.n19 GNDA.t131 493.418
R859 GNDA.n26 GNDA.t119 493.418
R860 GNDA.n25 GNDA.t208 493.418
R861 GNDA.n2377 GNDA.n2375 489.601
R862 GNDA.n359 GNDA.n346 486.401
R863 GNDA.n2362 GNDA.n2333 476.8
R864 GNDA.n2474 GNDA.n47 476.8
R865 GNDA.n2361 GNDA.n2334 454.401
R866 GNDA.n2475 GNDA.n46 454.401
R867 GNDA.n1817 GNDA.n1803 453.007
R868 GNDA.n2206 GNDA.n2205 446.486
R869 GNDA.n1333 GNDA.n1329 444.8
R870 GNDA.n1333 GNDA.n1332 444.8
R871 GNDA.n1332 GNDA.n1331 441.601
R872 GNDA.n1330 GNDA.n1329 438.401
R873 GNDA.n347 GNDA.n343 435.2
R874 GNDA.n2437 GNDA.n2436 428.8
R875 GNDA.n1761 GNDA.n343 425.601
R876 GNDA.n17 GNDA.n16 422.401
R877 GNDA.n14 GNDA.n10 422.401
R878 GNDA.n28 GNDA.n27 422.401
R879 GNDA.n33 GNDA.n32 422.401
R880 GNDA.n1760 GNDA.n345 422.401
R881 GNDA.n1761 GNDA.n1760 419.2
R882 GNDA.n77 GNDA.t183 413.084
R883 GNDA.n79 GNDA.t122 413.084
R884 GNDA.n2190 GNDA.t162 413.084
R885 GNDA.n62 GNDA.t159 413.084
R886 GNDA.n2153 GNDA.t156 413.084
R887 GNDA.n81 GNDA.t186 413.084
R888 GNDA.n2332 GNDA.n2329 393.601
R889 GNDA.n2460 GNDA.n2259 393.601
R890 GNDA.n2368 GNDA.n2332 387.2
R891 GNDA.n2461 GNDA.n2460 387.2
R892 GNDA.n2205 GNDA.n66 376.262
R893 GNDA.n1172 GNDA.n373 370.214
R894 GNDA.n690 GNDA.n376 370.214
R895 GNDA.n1172 GNDA.n372 365.957
R896 GNDA.n690 GNDA.n375 365.957
R897 GNDA.n2438 GNDA.n2437 355.2
R898 GNDA.n1724 GNDA.n1723 352.627
R899 GNDA.n534 GNDA.n374 352.627
R900 GNDA.n534 GNDA.n521 352.627
R901 GNDA.n830 GNDA.n521 352.627
R902 GNDA.n831 GNDA.n830 352.627
R903 GNDA.n832 GNDA.n831 352.627
R904 GNDA.n768 GNDA.n361 343.452
R905 GNDA.n1734 GNDA.n362 343.452
R906 GNDA.t135 GNDA.n1722 342.784
R907 GNDA.n1773 GNDA.t137 342.784
R908 GNDA.t137 GNDA.n1831 342.784
R909 GNDA.n2366 GNDA.n2334 342.401
R910 GNDA.n2254 GNDA.n46 342.401
R911 GNDA.n2349 GNDA.n2345 332.8
R912 GNDA.n2469 GNDA.n2246 332.8
R913 GNDA.n2276 GNDA.t165 332.75
R914 GNDA.n2278 GNDA.t147 332.75
R915 GNDA.t135 GNDA.n372 327.661
R916 GNDA.t137 GNDA.n200 172.876
R917 GNDA.t135 GNDA.n375 327.661
R918 GNDA.t137 GNDA.n203 172.876
R919 GNDA.t135 GNDA.n373 323.404
R920 GNDA.t137 GNDA.n205 172.615
R921 GNDA.t135 GNDA.n376 323.404
R922 GNDA.n202 GNDA.t137 172.615
R923 GNDA.n87 GNDA.n86 323.2
R924 GNDA.n2348 GNDA.n2347 321.281
R925 GNDA.n2468 GNDA.n2467 321.281
R926 GNDA.n2349 GNDA.n2348 318.08
R927 GNDA.n2469 GNDA.n2468 318.08
R928 GNDA.n86 GNDA.n68 316.8
R929 GNDA.n2428 GNDA.n2315 310.401
R930 GNDA.n2376 GNDA.n2263 310.401
R931 GNDA.n763 GNDA.n562 304
R932 GNDA.n2373 GNDA.n2317 304
R933 GNDA.n2375 GNDA.n2261 304
R934 GNDA.n2152 GNDA.n2151 303.99
R935 GNDA.n371 GNDA.n362 301.474
R936 GNDA.n761 GNDA.n562 300.8
R937 GNDA.n763 GNDA.n762 300.8
R938 GNDA.n2297 GNDA.n2286 300.8
R939 GNDA.n2298 GNDA.n2297 300.8
R940 GNDA.n2345 GNDA.n2318 300.8
R941 GNDA.n2247 GNDA.n2246 300.8
R942 GNDA.n762 GNDA.n761 297.601
R943 GNDA.n1340 GNDA.n342 297.601
R944 GNDA.n1340 GNDA.n1339 297.601
R945 GNDA.n1338 GNDA.n1136 297.601
R946 GNDA.n1139 GNDA.n1136 297.601
R947 GNDA.n766 GNDA.n765 296.411
R948 GNDA.n2338 GNDA.n2337 296
R949 GNDA.n2479 GNDA.n2478 296
R950 GNDA.n88 GNDA.n87 294.401
R951 GNDA.n2180 GNDA.n2179 294.401
R952 GNDA.n2193 GNDA.n2180 294.401
R953 GNDA.n2299 GNDA.n2298 292.5
R954 GNDA.n2300 GNDA.n2299 292.5
R955 GNDA.n2297 GNDA.n2275 292.5
R956 GNDA.n2275 GNDA.n2274 292.5
R957 GNDA.n2286 GNDA.n2285 292.5
R958 GNDA.n2285 GNDA.n2284 292.5
R959 GNDA.n2279 GNDA.n2273 292.5
R960 GNDA.n2274 GNDA.n2273 292.5
R961 GNDA.n2499 GNDA.n2498 292.5
R962 GNDA.n2498 GNDA.n2497 292.5
R963 GNDA.n6 GNDA.n3 292.5
R964 GNDA.n2301 GNDA.n6 292.5
R965 GNDA.n2303 GNDA.n2302 292.5
R966 GNDA.n2304 GNDA.n2303 292.5
R967 GNDA.n5 GNDA.n4 292.5
R968 GNDA.n2301 GNDA.n5 292.5
R969 GNDA.n2444 GNDA.n2443 292.5
R970 GNDA.n2443 GNDA.n2442 292.5
R971 GNDA.n2446 GNDA.n2268 292.5
R972 GNDA.n2283 GNDA.n2268 292.5
R973 GNDA.n2449 GNDA.n2448 292.5
R974 GNDA.n2450 GNDA.n2449 292.5
R975 GNDA.n2269 GNDA.n2267 292.5
R976 GNDA.n2283 GNDA.n2267 292.5
R977 GNDA.n2435 GNDA.n2434 292.5
R978 GNDA.n2434 GNDA.n2433 292.5
R979 GNDA.n2437 GNDA.n2306 292.5
R980 GNDA.n2306 GNDA.n2305 292.5
R981 GNDA.n2440 GNDA.n2439 292.5
R982 GNDA.n2441 GNDA.n2440 292.5
R983 GNDA.n2307 GNDA.n2272 292.5
R984 GNDA.n2305 GNDA.n2272 292.5
R985 GNDA.n34 GNDA.n24 292.5
R986 GNDA.n2432 GNDA.n24 292.5
R987 GNDA.n36 GNDA.n35 292.5
R988 GNDA.n2490 GNDA.n36 292.5
R989 GNDA.n29 GNDA.n23 292.5
R990 GNDA.n2451 GNDA.n23 292.5
R991 GNDA.n2492 GNDA.n2491 292.5
R992 GNDA.n2491 GNDA.n2490 292.5
R993 GNDA.n2495 GNDA.n2494 292.5
R994 GNDA.n2496 GNDA.n2495 292.5
R995 GNDA.n2493 GNDA.n8 292.5
R996 GNDA.n2490 GNDA.n8 292.5
R997 GNDA.n2281 GNDA.n18 292.5
R998 GNDA.n2282 GNDA.n2281 292.5
R999 GNDA.n15 GNDA.n7 292.5
R1000 GNDA.n2490 GNDA.n7 292.5
R1001 GNDA.n2350 GNDA.n2349 292.5
R1002 GNDA.n2351 GNDA.n2350 292.5
R1003 GNDA.n2348 GNDA.n2344 292.5
R1004 GNDA.n2344 GNDA.n2343 292.5
R1005 GNDA.n2345 GNDA.n2341 292.5
R1006 GNDA.n2343 GNDA.n2341 292.5
R1007 GNDA.n2336 GNDA.n2334 292.5
R1008 GNDA.n2356 GNDA.n2336 292.5
R1009 GNDA.n2366 GNDA.n2365 292.5
R1010 GNDA.n2365 GNDA.n2364 292.5
R1011 GNDA.n2335 GNDA.n2333 292.5
R1012 GNDA.n2340 GNDA.n2335 292.5
R1013 GNDA.n2363 GNDA.n2362 292.5
R1014 GNDA.n2364 GNDA.n2363 292.5
R1015 GNDA.n2353 GNDA.n2337 292.5
R1016 GNDA.n2353 GNDA.n2352 292.5
R1017 GNDA.n2347 GNDA.n2346 292.5
R1018 GNDA.n2346 GNDA.n2319 292.5
R1019 GNDA.n2369 GNDA.n2368 292.5
R1020 GNDA.n2370 GNDA.n2369 292.5
R1021 GNDA.n2332 GNDA.n2322 292.5
R1022 GNDA.n2322 GNDA.t78 292.5
R1023 GNDA.n2329 GNDA.n2328 292.5
R1024 GNDA.n2328 GNDA.n2311 292.5
R1025 GNDA.n2326 GNDA.n2320 292.5
R1026 GNDA.t78 GNDA.n2320 292.5
R1027 GNDA.n2429 GNDA.n2428 292.5
R1028 GNDA.n2430 GNDA.n2429 292.5
R1029 GNDA.n2330 GNDA.n2312 292.5
R1030 GNDA.n2321 GNDA.n2312 292.5
R1031 GNDA.n2373 GNDA.n2372 292.5
R1032 GNDA.n2372 GNDA.n2371 292.5
R1033 GNDA.n2427 GNDA.n2313 292.5
R1034 GNDA.n2321 GNDA.n2313 292.5
R1035 GNDA.n2376 GNDA.n2265 292.5
R1036 GNDA.n2453 GNDA.n2265 292.5
R1037 GNDA.n2377 GNDA.n2266 292.5
R1038 GNDA.n2456 GNDA.n2266 292.5
R1039 GNDA.n2375 GNDA.n2264 292.5
R1040 GNDA.n2264 GNDA.n2249 292.5
R1041 GNDA.n2458 GNDA.n2457 292.5
R1042 GNDA.n2457 GNDA.n2456 292.5
R1043 GNDA.n2454 GNDA.n2259 292.5
R1044 GNDA.n2455 GNDA.n2454 292.5
R1045 GNDA.n2460 GNDA.n2251 292.5
R1046 GNDA.t52 GNDA.n2251 292.5
R1047 GNDA.n2462 GNDA.n2461 292.5
R1048 GNDA.n2463 GNDA.n2462 292.5
R1049 GNDA.n2257 GNDA.n2250 292.5
R1050 GNDA.t52 GNDA.n2250 292.5
R1051 GNDA.n2478 GNDA.n2477 292.5
R1052 GNDA.n2477 GNDA.n43 292.5
R1053 GNDA.n2178 GNDA.n2177 292.5
R1054 GNDA.n2177 GNDA.n2176 292.5
R1055 GNDA.n2156 GNDA.n2155 292.5
R1056 GNDA.n2157 GNDA.n2156 292.5
R1057 GNDA.n89 GNDA.n80 292.5
R1058 GNDA.n90 GNDA.n89 292.5
R1059 GNDA.n2193 GNDA.n76 292.5
R1060 GNDA.n2184 GNDA.n76 292.5
R1061 GNDA.n2196 GNDA.n2195 292.5
R1062 GNDA.n2199 GNDA.n2196 292.5
R1063 GNDA.n2179 GNDA.n75 292.5
R1064 GNDA.n2175 GNDA.n75 292.5
R1065 GNDA.n2180 GNDA.n74 292.5
R1066 GNDA.n2199 GNDA.n74 292.5
R1067 GNDA.n2467 GNDA.n2466 292.5
R1068 GNDA.n2466 GNDA.n2465 292.5
R1069 GNDA.n2468 GNDA.n2245 292.5
R1070 GNDA.n2464 GNDA.n2245 292.5
R1071 GNDA.n2470 GNDA.n2469 292.5
R1072 GNDA.n2471 GNDA.n2470 292.5
R1073 GNDA.n2246 GNDA.n2244 292.5
R1074 GNDA.n2464 GNDA.n2244 292.5
R1075 GNDA.n2210 GNDA.n2209 292.5
R1076 GNDA.n2209 GNDA.n2208 292.5
R1077 GNDA.n2192 GNDA.n2189 292.5
R1078 GNDA.n2189 GNDA.n2188 292.5
R1079 GNDA.n2185 GNDA.n61 292.5
R1080 GNDA.n2186 GNDA.n2185 292.5
R1081 GNDA.n72 GNDA.n70 292.5
R1082 GNDA.n72 GNDA.n53 292.5
R1083 GNDA.n2198 GNDA.n2197 292.5
R1084 GNDA.n2199 GNDA.n2198 292.5
R1085 GNDA.n71 GNDA.n69 292.5
R1086 GNDA.n2159 GNDA.n71 292.5
R1087 GNDA.n2201 GNDA.n2200 292.5
R1088 GNDA.n2200 GNDA.n2199 292.5
R1089 GNDA.n2168 GNDA.n2163 292.5
R1090 GNDA.n2163 GNDA.n2162 292.5
R1091 GNDA.n2167 GNDA.n91 292.5
R1092 GNDA.n2171 GNDA.n91 292.5
R1093 GNDA.n2164 GNDA.n2161 292.5
R1094 GNDA.n2161 GNDA.n2160 292.5
R1095 GNDA.n2170 GNDA.n2169 292.5
R1096 GNDA.n2171 GNDA.n2170 292.5
R1097 GNDA.n2238 GNDA.n2237 292.5
R1098 GNDA.n2239 GNDA.n2238 292.5
R1099 GNDA.n2236 GNDA.n55 292.5
R1100 GNDA.n2187 GNDA.n55 292.5
R1101 GNDA.n2181 GNDA.n57 292.5
R1102 GNDA.n2182 GNDA.n2181 292.5
R1103 GNDA.n56 GNDA.n54 292.5
R1104 GNDA.n2187 GNDA.n54 292.5
R1105 GNDA.n2173 GNDA.n68 292.5
R1106 GNDA.n2174 GNDA.n2173 292.5
R1107 GNDA.n2172 GNDA.n88 292.5
R1108 GNDA.n2172 GNDA.n2171 292.5
R1109 GNDA.n87 GNDA.n85 292.5
R1110 GNDA.n2158 GNDA.n85 292.5
R1111 GNDA.n86 GNDA.n84 292.5
R1112 GNDA.n2171 GNDA.n84 292.5
R1113 GNDA.n2474 GNDA.n2473 292.5
R1114 GNDA.n2473 GNDA.n2472 292.5
R1115 GNDA.n49 GNDA.n47 292.5
R1116 GNDA.n2243 GNDA.n49 292.5
R1117 GNDA.n2254 GNDA.n2242 292.5
R1118 GNDA.n2472 GNDA.n2242 292.5
R1119 GNDA.n48 GNDA.n46 292.5
R1120 GNDA.n2241 GNDA.n48 292.5
R1121 GNDA.n2207 GNDA.n2206 292.5
R1122 GNDA.n2204 GNDA.n67 292.5
R1123 GNDA.n2183 GNDA.n67 292.5
R1124 GNDA.n2187 GNDA.n66 292.5
R1125 GNDA.n1136 GNDA.n1131 292.5
R1126 GNDA.n1342 GNDA.n1131 292.5
R1127 GNDA.n1140 GNDA.n1139 292.5
R1128 GNDA.n1336 GNDA.n1140 292.5
R1129 GNDA.n1137 GNDA.n1135 292.5
R1130 GNDA.n1163 GNDA.n1137 292.5
R1131 GNDA.n1338 GNDA.n1337 292.5
R1132 GNDA.n1337 GNDA.n1336 292.5
R1133 GNDA.n764 GNDA.n763 292.5
R1134 GNDA.n765 GNDA.n764 292.5
R1135 GNDA.n762 GNDA.n561 292.5
R1136 GNDA.n729 GNDA.n561 292.5
R1137 GNDA.n761 GNDA.n760 292.5
R1138 GNDA.n760 GNDA.n759 292.5
R1139 GNDA.n562 GNDA.n560 292.5
R1140 GNDA.n729 GNDA.n560 292.5
R1141 GNDA.n1341 GNDA.n1340 292.5
R1142 GNDA.n1342 GNDA.n1341 292.5
R1143 GNDA.n1339 GNDA.n1133 292.5
R1144 GNDA.n1336 GNDA.n1133 292.5
R1145 GNDA.n1162 GNDA.n1134 292.5
R1146 GNDA.n1163 GNDA.n1162 292.5
R1147 GNDA.n1132 GNDA.n342 292.5
R1148 GNDA.n1336 GNDA.n1132 292.5
R1149 GNDA.n1332 GNDA.n1328 292.5
R1150 GNDA.n1328 GNDA.n350 292.5
R1151 GNDA.n1331 GNDA.n1141 292.5
R1152 GNDA.n1335 GNDA.n1141 292.5
R1153 GNDA.n1329 GNDA.n1327 292.5
R1154 GNDA.n1327 GNDA.n1326 292.5
R1155 GNDA.n1334 GNDA.n1333 292.5
R1156 GNDA.n1335 GNDA.n1334 292.5
R1157 GNDA.n1747 GNDA.n357 292.5
R1158 GNDA.n729 GNDA.n357 292.5
R1159 GNDA.n1746 GNDA.n1745 292.5
R1160 GNDA.n1745 GNDA.n1744 292.5
R1161 GNDA.n359 GNDA.n358 292.5
R1162 GNDA.n729 GNDA.n358 292.5
R1163 GNDA.n1749 GNDA.n1748 292.5
R1164 GNDA.n1750 GNDA.n1749 292.5
R1165 GNDA.n1760 GNDA.n1759 292.5
R1166 GNDA.n1759 GNDA.n1758 292.5
R1167 GNDA.n348 GNDA.n347 292.5
R1168 GNDA.n1336 GNDA.n348 292.5
R1169 GNDA.n1143 GNDA.n343 292.5
R1170 GNDA.n1326 GNDA.n1143 292.5
R1171 GNDA.n1761 GNDA.n344 292.5
R1172 GNDA.n1336 GNDA.n344 292.5
R1173 GNDA.n1134 GNDA.n342 291.2
R1174 GNDA.n1339 GNDA.n1134 291.2
R1175 GNDA.n1338 GNDA.n1135 291.2
R1176 GNDA.n1139 GNDA.n1135 291.2
R1177 GNDA.n88 GNDA.n68 288
R1178 GNDA.n2191 GNDA.n63 281.601
R1179 GNDA.n2154 GNDA.n82 281.601
R1180 GNDA.n2210 GNDA.n61 278.401
R1181 GNDA.n2155 GNDA.n80 278.401
R1182 GNDA.n1326 GNDA.n1142 276.707
R1183 GNDA.n2151 GNDA.n93 264.301
R1184 GNDA.n587 GNDA.n390 259.416
R1185 GNDA.n1845 GNDA.n1844 259.416
R1186 GNDA.n1199 GNDA.n396 259.416
R1187 GNDA.n1437 GNDA.n1436 259.416
R1188 GNDA.n2066 GNDA.n2065 259.416
R1189 GNDA.n989 GNDA.n988 259.416
R1190 GNDA.n458 GNDA.n99 259.416
R1191 GNDA.n2114 GNDA.n2113 259.416
R1192 GNDA.n833 GNDA.n403 259.416
R1193 GNDA.n2276 GNDA.t166 258.601
R1194 GNDA.n2278 GNDA.t149 258.601
R1195 GNDA.n190 GNDA.n189 254.442
R1196 GNDA.n923 GNDA.n205 254.34
R1197 GNDA.n920 GNDA.n205 254.34
R1198 GNDA.n902 GNDA.n205 254.34
R1199 GNDA.n913 GNDA.n205 254.34
R1200 GNDA.n905 GNDA.n205 254.34
R1201 GNDA.n906 GNDA.n205 254.34
R1202 GNDA.n695 GNDA.n376 254.34
R1203 GNDA.n718 GNDA.n376 254.34
R1204 GNDA.n698 GNDA.n376 254.34
R1205 GNDA.n711 GNDA.n376 254.34
R1206 GNDA.n701 GNDA.n376 254.34
R1207 GNDA.n704 GNDA.n376 254.34
R1208 GNDA.n2151 GNDA.n105 254.34
R1209 GNDA.n2151 GNDA.n104 254.34
R1210 GNDA.n2151 GNDA.n103 254.34
R1211 GNDA.n2151 GNDA.n102 254.34
R1212 GNDA.n2151 GNDA.n101 254.34
R1213 GNDA.n2151 GNDA.n100 254.34
R1214 GNDA.n2151 GNDA.n98 254.34
R1215 GNDA.n2151 GNDA.n97 254.34
R1216 GNDA.n2151 GNDA.n96 254.34
R1217 GNDA.n2151 GNDA.n95 254.34
R1218 GNDA.n2151 GNDA.n94 254.34
R1219 GNDA.n1965 GNDA.n264 254.34
R1220 GNDA.n1965 GNDA.n265 254.34
R1221 GNDA.n1965 GNDA.n266 254.34
R1222 GNDA.n1965 GNDA.n267 254.34
R1223 GNDA.n1965 GNDA.n1964 254.34
R1224 GNDA.n262 GNDA.n108 254.34
R1225 GNDA.n1965 GNDA.n263 254.34
R1226 GNDA.n1965 GNDA.n261 254.34
R1227 GNDA.n1965 GNDA.n260 254.34
R1228 GNDA.n1965 GNDA.n259 254.34
R1229 GNDA.n1965 GNDA.n258 254.34
R1230 GNDA.n284 GNDA.n273 254.34
R1231 GNDA.n1952 GNDA.n273 254.34
R1232 GNDA.n280 GNDA.n273 254.34
R1233 GNDA.n1959 GNDA.n273 254.34
R1234 GNDA.n273 GNDA.n272 254.34
R1235 GNDA.n1587 GNDA.n459 254.34
R1236 GNDA.n1583 GNDA.n273 254.34
R1237 GNDA.n1581 GNDA.n273 254.34
R1238 GNDA.n1573 GNDA.n273 254.34
R1239 GNDA.n1571 GNDA.n273 254.34
R1240 GNDA.n1563 GNDA.n273 254.34
R1241 GNDA.n1965 GNDA.n256 254.34
R1242 GNDA.n1965 GNDA.n255 254.34
R1243 GNDA.n1965 GNDA.n254 254.34
R1244 GNDA.n1965 GNDA.n253 254.34
R1245 GNDA.n1965 GNDA.n252 254.34
R1246 GNDA.n886 GNDA.n273 254.34
R1247 GNDA.n1428 GNDA.n273 254.34
R1248 GNDA.n1420 GNDA.n273 254.34
R1249 GNDA.n1418 GNDA.n273 254.34
R1250 GNDA.n1410 GNDA.n273 254.34
R1251 GNDA.n1386 GNDA.n928 254.34
R1252 GNDA.n1392 GNDA.n928 254.34
R1253 GNDA.n1394 GNDA.n928 254.34
R1254 GNDA.n1400 GNDA.n928 254.34
R1255 GNDA.n1402 GNDA.n928 254.34
R1256 GNDA.n1408 GNDA.n928 254.34
R1257 GNDA.n1538 GNDA.n504 254.34
R1258 GNDA.n1544 GNDA.n504 254.34
R1259 GNDA.n1546 GNDA.n504 254.34
R1260 GNDA.n1552 GNDA.n504 254.34
R1261 GNDA.n1554 GNDA.n504 254.34
R1262 GNDA.n1560 GNDA.n504 254.34
R1263 GNDA.n437 GNDA.n436 254.34
R1264 GNDA.n1686 GNDA.n435 254.34
R1265 GNDA.n1686 GNDA.n434 254.34
R1266 GNDA.n1686 GNDA.n433 254.34
R1267 GNDA.n1686 GNDA.n432 254.34
R1268 GNDA.n1686 GNDA.n431 254.34
R1269 GNDA.n836 GNDA.n835 254.34
R1270 GNDA.n1694 GNDA.n404 254.34
R1271 GNDA.n1694 GNDA.n405 254.34
R1272 GNDA.n1694 GNDA.n406 254.34
R1273 GNDA.n1694 GNDA.n407 254.34
R1274 GNDA.n1694 GNDA.n408 254.34
R1275 GNDA.n1686 GNDA.n429 254.34
R1276 GNDA.n1686 GNDA.n428 254.34
R1277 GNDA.n1686 GNDA.n427 254.34
R1278 GNDA.n1686 GNDA.n426 254.34
R1279 GNDA.n1686 GNDA.n425 254.34
R1280 GNDA.n1694 GNDA.n402 254.34
R1281 GNDA.n1694 GNDA.n401 254.34
R1282 GNDA.n1694 GNDA.n400 254.34
R1283 GNDA.n1694 GNDA.n399 254.34
R1284 GNDA.n1694 GNDA.n398 254.34
R1285 GNDA.n1965 GNDA.n251 254.34
R1286 GNDA.n312 GNDA.n200 254.34
R1287 GNDA.n1919 GNDA.n200 254.34
R1288 GNDA.n306 GNDA.n200 254.34
R1289 GNDA.n1930 GNDA.n200 254.34
R1290 GNDA.n297 GNDA.n200 254.34
R1291 GNDA.n1941 GNDA.n200 254.34
R1292 GNDA.n1686 GNDA.n424 254.34
R1293 GNDA.n985 GNDA.n962 254.34
R1294 GNDA.n1063 GNDA.n962 254.34
R1295 GNDA.n979 GNDA.n962 254.34
R1296 GNDA.n1074 GNDA.n962 254.34
R1297 GNDA.n970 GNDA.n962 254.34
R1298 GNDA.n1085 GNDA.n962 254.34
R1299 GNDA.n987 GNDA.n984 254.34
R1300 GNDA.n1198 GNDA.n372 254.34
R1301 GNDA.n1273 GNDA.n372 254.34
R1302 GNDA.n1191 GNDA.n372 254.34
R1303 GNDA.n1284 GNDA.n372 254.34
R1304 GNDA.n1178 GNDA.n372 254.34
R1305 GNDA.n1175 GNDA.n372 254.34
R1306 GNDA.n1197 GNDA.n1196 254.34
R1307 GNDA.n1686 GNDA.n423 254.34
R1308 GNDA.n1686 GNDA.n422 254.34
R1309 GNDA.n1686 GNDA.n421 254.34
R1310 GNDA.n1686 GNDA.n420 254.34
R1311 GNDA.n1686 GNDA.n419 254.34
R1312 GNDA.n1694 GNDA.n395 254.34
R1313 GNDA.n1694 GNDA.n394 254.34
R1314 GNDA.n1694 GNDA.n393 254.34
R1315 GNDA.n1694 GNDA.n392 254.34
R1316 GNDA.n1694 GNDA.n391 254.34
R1317 GNDA.n1363 GNDA.n373 254.34
R1318 GNDA.n1365 GNDA.n373 254.34
R1319 GNDA.n1371 GNDA.n373 254.34
R1320 GNDA.n1373 GNDA.n373 254.34
R1321 GNDA.n1379 GNDA.n373 254.34
R1322 GNDA.n1382 GNDA.n373 254.34
R1323 GNDA.n1966 GNDA.n1965 254.34
R1324 GNDA.n1687 GNDA.n1686 254.34
R1325 GNDA.n885 GNDA.n861 254.34
R1326 GNDA.n1511 GNDA.n861 254.34
R1327 GNDA.n879 GNDA.n861 254.34
R1328 GNDA.n1522 GNDA.n861 254.34
R1329 GNDA.n870 GNDA.n861 254.34
R1330 GNDA.n1533 GNDA.n861 254.34
R1331 GNDA.n1435 GNDA.n884 254.34
R1332 GNDA.n588 GNDA.n375 254.34
R1333 GNDA.n664 GNDA.n375 254.34
R1334 GNDA.n585 GNDA.n375 254.34
R1335 GNDA.n675 GNDA.n375 254.34
R1336 GNDA.n576 GNDA.n375 254.34
R1337 GNDA.n686 GNDA.n375 254.34
R1338 GNDA.n1692 GNDA.n1691 254.34
R1339 GNDA.n2064 GNDA.n203 254.34
R1340 GNDA.n2029 GNDA.n203 254.34
R1341 GNDA.n2042 GNDA.n203 254.34
R1342 GNDA.n2027 GNDA.n203 254.34
R1343 GNDA.n2052 GNDA.n203 254.34
R1344 GNDA.n2022 GNDA.n203 254.34
R1345 GNDA.n499 GNDA.n202 254.34
R1346 GNDA.n473 GNDA.n202 254.34
R1347 GNDA.n492 GNDA.n202 254.34
R1348 GNDA.n486 GNDA.n202 254.34
R1349 GNDA.n484 GNDA.n202 254.34
R1350 GNDA.n478 GNDA.n202 254.34
R1351 GNDA.n1843 GNDA.n311 254.34
R1352 GNDA.n2068 GNDA.n2067 254.34
R1353 GNDA.n1171 GNDA.n1170 254.34
R1354 GNDA.n564 GNDA.n353 254.34
R1355 GNDA.n732 GNDA.n731 254.34
R1356 GNDA.n1743 GNDA.n361 251.865
R1357 GNDA.n1769 GNDA.n336 250.349
R1358 GNDA.n826 GNDA.n825 250
R1359 GNDA.n1657 GNDA.n1656 250
R1360 GNDA.n187 GNDA.n122 250
R1361 GNDA.n1269 GNDA.n1268 250
R1362 GNDA.n1059 GNDA.n1058 250
R1363 GNDA.n1915 GNDA.n1914 250
R1364 GNDA.n660 GNDA.n659 250
R1365 GNDA.n1507 GNDA.n1506 250
R1366 GNDA.n2059 GNDA.n225 250
R1367 GNDA.n1383 GNDA.n1121 249.663
R1368 GNDA.n1818 GNDA.n1804 249.663
R1369 GNDA.n397 GNDA.n385 249.663
R1370 GNDA.n1411 GNDA.n1409 249.663
R1371 GNDA.n2087 GNDA.n208 249.663
R1372 GNDA.n1783 GNDA.n329 249.663
R1373 GNDA.n1562 GNDA.n1561 249.663
R1374 GNDA.n479 GNDA.n199 249.663
R1375 GNDA.n703 GNDA.n409 249.663
R1376 GNDA.n2367 GNDA.n2366 246.4
R1377 GNDA.n2255 GNDA.n2254 246.4
R1378 GNDA.n2360 GNDA.n2359 244.8
R1379 GNDA.n2476 GNDA.n45 244.8
R1380 GNDA.n1744 GNDA.n1743 242.96
R1381 GNDA.n2192 GNDA.n61 240
R1382 GNDA.n2178 GNDA.n80 240
R1383 GNDA.t135 GNDA.n374 239.004
R1384 GNDA.n2448 GNDA.n2269 233.601
R1385 GNDA.n2444 GNDA.n2269 233.601
R1386 GNDA.n2292 GNDA.n2290 227.096
R1387 GNDA.n2289 GNDA.n2287 227.096
R1388 GNDA.n2292 GNDA.n2291 226.534
R1389 GNDA.n2289 GNDA.n2288 226.534
R1390 GNDA.n2316 GNDA.t130 224.525
R1391 GNDA.n2314 GNDA.t146 224.525
R1392 GNDA.n2262 GNDA.t195 224.525
R1393 GNDA.n2260 GNDA.t201 224.525
R1394 GNDA.n1744 GNDA.n360 223.524
R1395 GNDA.n2295 GNDA.n2294 222.034
R1396 GNDA.n791 GNDA.n551 221.667
R1397 GNDA.n1622 GNDA.n1599 221.667
R1398 GNDA.n154 GNDA.n152 221.667
R1399 GNDA.n1234 GNDA.n1211 221.667
R1400 GNDA.n1024 GNDA.n1001 221.667
R1401 GNDA.n1880 GNDA.n1857 221.667
R1402 GNDA.n625 GNDA.n602 221.667
R1403 GNDA.n1472 GNDA.n1449 221.667
R1404 GNDA.n2002 GNDA.n2001 221.667
R1405 GNDA.n2499 GNDA.n4 217.601
R1406 GNDA.n2302 GNDA.n4 214.4
R1407 GNDA.n2280 GNDA.n2279 211.201
R1408 GNDA.n2279 GNDA.n2277 211.201
R1409 GNDA.n2327 GNDA.n2326 211.201
R1410 GNDA.n2326 GNDA.n2324 211.201
R1411 GNDA.n2257 GNDA.n2253 211.201
R1412 GNDA.n2258 GNDA.n2257 211.201
R1413 GNDA.n2485 GNDA.n40 209.183
R1414 GNDA.n2504 GNDA.n2502 206.177
R1415 GNDA.n2383 GNDA.n2381 206.052
R1416 GNDA.n2512 GNDA.n2511 205.488
R1417 GNDA.n2510 GNDA.n2509 205.488
R1418 GNDA.n2508 GNDA.n2507 205.488
R1419 GNDA.n2506 GNDA.n2505 205.488
R1420 GNDA.n2504 GNDA.n2503 205.488
R1421 GNDA.n2391 GNDA.n2390 205.488
R1422 GNDA.n2389 GNDA.n2388 205.488
R1423 GNDA.n2387 GNDA.n2386 205.488
R1424 GNDA.n2385 GNDA.n2384 205.488
R1425 GNDA.n2383 GNDA.n2382 205.488
R1426 GNDA.n2302 GNDA.n3 203.201
R1427 GNDA.n2500 GNDA.n2499 201.601
R1428 GNDA.n1768 GNDA.n337 197
R1429 GNDA.n688 GNDA.n565 197
R1430 GNDA.n1300 GNDA.n1299 197
R1431 GNDA.n1535 GNDA.n415 197
R1432 GNDA.n1685 GNDA.n1684 197
R1433 GNDA.n2150 GNDA.n107 197
R1434 GNDA.n767 GNDA.n558 197
R1435 GNDA.n1943 GNDA.n287 197
R1436 GNDA.n249 GNDA.n247 197
R1437 GNDA.n960 GNDA.n859 197
R1438 GNDA.n2359 GNDA.n2358 195
R1439 GNDA.n2358 GNDA.n2357 195
R1440 GNDA.n2339 GNDA.n2338 195
R1441 GNDA.n2342 GNDA.n2339 195
R1442 GNDA.n2480 GNDA.n2479 195
R1443 GNDA.n2481 GNDA.n2480 195
R1444 GNDA.n51 GNDA.n45 195
R1445 GNDA.n52 GNDA.n51 195
R1446 GNDA.n2330 GNDA.n2315 192
R1447 GNDA.n2458 GNDA.n2263 192
R1448 GNDA.n1326 GNDA.n1325 191.939
R1449 GNDA.t137 GNDA.n206 190.773
R1450 GNDA.t137 GNDA.n201 190.773
R1451 GNDA.n1358 GNDA.n1127 187.249
R1452 GNDA.n1324 GNDA.n1146 187.249
R1453 GNDA.n1095 GNDA.n858 187.249
R1454 GNDA.n1537 GNDA.n430 187.249
R1455 GNDA.n472 GNDA.n257 187.249
R1456 GNDA.n757 GNDA.n693 187.249
R1457 GNDA.n1787 GNDA.n268 187.249
R1458 GNDA.n898 GNDA.n896 187.249
R1459 GNDA.n1708 GNDA.n389 187.249
R1460 GNDA.t137 GNDA.n2088 186.691
R1461 GNDA.n2089 GNDA.t137 186.691
R1462 GNDA.n773 GNDA.n556 185
R1463 GNDA.n775 GNDA.n774 185
R1464 GNDA.n777 GNDA.n554 185
R1465 GNDA.n780 GNDA.n779 185
R1466 GNDA.n781 GNDA.n553 185
R1467 GNDA.n783 GNDA.n782 185
R1468 GNDA.n785 GNDA.n552 185
R1469 GNDA.n788 GNDA.n787 185
R1470 GNDA.n789 GNDA.n551 185
R1471 GNDA.n791 GNDA.n790 185
R1472 GNDA.n793 GNDA.n550 185
R1473 GNDA.n796 GNDA.n795 185
R1474 GNDA.n797 GNDA.n549 185
R1475 GNDA.n799 GNDA.n798 185
R1476 GNDA.n801 GNDA.n548 185
R1477 GNDA.n804 GNDA.n803 185
R1478 GNDA.n805 GNDA.n547 185
R1479 GNDA.n807 GNDA.n806 185
R1480 GNDA.n825 GNDA.n542 185
R1481 GNDA.n823 GNDA.n822 185
R1482 GNDA.n821 GNDA.n543 185
R1483 GNDA.n820 GNDA.n819 185
R1484 GNDA.n817 GNDA.n544 185
R1485 GNDA.n815 GNDA.n814 185
R1486 GNDA.n813 GNDA.n545 185
R1487 GNDA.n812 GNDA.n811 185
R1488 GNDA.n809 GNDA.n546 185
R1489 GNDA.n1604 GNDA.n1603 185
R1490 GNDA.n1606 GNDA.n1605 185
R1491 GNDA.n1608 GNDA.n1602 185
R1492 GNDA.n1611 GNDA.n1610 185
R1493 GNDA.n1612 GNDA.n1601 185
R1494 GNDA.n1614 GNDA.n1613 185
R1495 GNDA.n1616 GNDA.n1600 185
R1496 GNDA.n1619 GNDA.n1618 185
R1497 GNDA.n1620 GNDA.n1599 185
R1498 GNDA.n1622 GNDA.n1621 185
R1499 GNDA.n1624 GNDA.n1598 185
R1500 GNDA.n1627 GNDA.n1626 185
R1501 GNDA.n1628 GNDA.n1597 185
R1502 GNDA.n1630 GNDA.n1629 185
R1503 GNDA.n1632 GNDA.n1596 185
R1504 GNDA.n1635 GNDA.n1634 185
R1505 GNDA.n1636 GNDA.n1595 185
R1506 GNDA.n1638 GNDA.n1637 185
R1507 GNDA.n1656 GNDA.n1590 185
R1508 GNDA.n1654 GNDA.n1653 185
R1509 GNDA.n1652 GNDA.n1591 185
R1510 GNDA.n1651 GNDA.n1650 185
R1511 GNDA.n1648 GNDA.n1592 185
R1512 GNDA.n1646 GNDA.n1645 185
R1513 GNDA.n1644 GNDA.n1593 185
R1514 GNDA.n1643 GNDA.n1642 185
R1515 GNDA.n1640 GNDA.n1594 185
R1516 GNDA.n136 GNDA.n109 185
R1517 GNDA.n139 GNDA.n138 185
R1518 GNDA.n140 GNDA.n134 185
R1519 GNDA.n142 GNDA.n141 185
R1520 GNDA.n144 GNDA.n133 185
R1521 GNDA.n147 GNDA.n146 185
R1522 GNDA.n148 GNDA.n132 185
R1523 GNDA.n150 GNDA.n149 185
R1524 GNDA.n152 GNDA.n131 185
R1525 GNDA.n155 GNDA.n154 185
R1526 GNDA.n156 GNDA.n130 185
R1527 GNDA.n158 GNDA.n157 185
R1528 GNDA.n160 GNDA.n129 185
R1529 GNDA.n163 GNDA.n162 185
R1530 GNDA.n164 GNDA.n128 185
R1531 GNDA.n166 GNDA.n165 185
R1532 GNDA.n168 GNDA.n127 185
R1533 GNDA.n171 GNDA.n170 185
R1534 GNDA.n188 GNDA.n187 185
R1535 GNDA.n185 GNDA.n120 185
R1536 GNDA.n184 GNDA.n123 185
R1537 GNDA.n182 GNDA.n181 185
R1538 GNDA.n180 GNDA.n124 185
R1539 GNDA.n179 GNDA.n178 185
R1540 GNDA.n176 GNDA.n125 185
R1541 GNDA.n174 GNDA.n173 185
R1542 GNDA.n172 GNDA.n126 185
R1543 GNDA.n122 GNDA.n119 185
R1544 GNDA.n2121 GNDA.n118 185
R1545 GNDA.n2126 GNDA.n2125 185
R1546 GNDA.n2129 GNDA.n2128 185
R1547 GNDA.n117 GNDA.n114 185
R1548 GNDA.n2134 GNDA.n113 185
R1549 GNDA.n2139 GNDA.n2138 185
R1550 GNDA.n2142 GNDA.n2141 185
R1551 GNDA.n112 GNDA.n110 185
R1552 GNDA.n1658 GNDA.n1657 185
R1553 GNDA.n454 GNDA.n450 185
R1554 GNDA.n1664 GNDA.n1663 185
R1555 GNDA.n1666 GNDA.n449 185
R1556 GNDA.n1668 GNDA.n1667 185
R1557 GNDA.n446 GNDA.n442 185
R1558 GNDA.n1674 GNDA.n1673 185
R1559 GNDA.n1676 GNDA.n441 185
R1560 GNDA.n1678 GNDA.n1677 185
R1561 GNDA.n827 GNDA.n826 185
R1562 GNDA.n540 GNDA.n523 185
R1563 GNDA.n539 GNDA.n538 185
R1564 GNDA.n529 GNDA.n526 185
R1565 GNDA.n531 GNDA.n530 185
R1566 GNDA.n369 GNDA.n368 185
R1567 GNDA.n1728 GNDA.n1727 185
R1568 GNDA.n1731 GNDA.n1730 185
R1569 GNDA.n367 GNDA.n365 185
R1570 GNDA.n1216 GNDA.n1176 185
R1571 GNDA.n1218 GNDA.n1217 185
R1572 GNDA.n1220 GNDA.n1214 185
R1573 GNDA.n1223 GNDA.n1222 185
R1574 GNDA.n1224 GNDA.n1213 185
R1575 GNDA.n1226 GNDA.n1225 185
R1576 GNDA.n1228 GNDA.n1212 185
R1577 GNDA.n1231 GNDA.n1230 185
R1578 GNDA.n1232 GNDA.n1211 185
R1579 GNDA.n1234 GNDA.n1233 185
R1580 GNDA.n1236 GNDA.n1210 185
R1581 GNDA.n1239 GNDA.n1238 185
R1582 GNDA.n1240 GNDA.n1209 185
R1583 GNDA.n1242 GNDA.n1241 185
R1584 GNDA.n1244 GNDA.n1208 185
R1585 GNDA.n1247 GNDA.n1246 185
R1586 GNDA.n1248 GNDA.n1207 185
R1587 GNDA.n1250 GNDA.n1249 185
R1588 GNDA.n1268 GNDA.n1202 185
R1589 GNDA.n1266 GNDA.n1265 185
R1590 GNDA.n1264 GNDA.n1203 185
R1591 GNDA.n1263 GNDA.n1262 185
R1592 GNDA.n1260 GNDA.n1204 185
R1593 GNDA.n1258 GNDA.n1257 185
R1594 GNDA.n1256 GNDA.n1205 185
R1595 GNDA.n1255 GNDA.n1254 185
R1596 GNDA.n1252 GNDA.n1206 185
R1597 GNDA.n1006 GNDA.n1005 185
R1598 GNDA.n1008 GNDA.n1007 185
R1599 GNDA.n1010 GNDA.n1004 185
R1600 GNDA.n1013 GNDA.n1012 185
R1601 GNDA.n1014 GNDA.n1003 185
R1602 GNDA.n1016 GNDA.n1015 185
R1603 GNDA.n1018 GNDA.n1002 185
R1604 GNDA.n1021 GNDA.n1020 185
R1605 GNDA.n1022 GNDA.n1001 185
R1606 GNDA.n1024 GNDA.n1023 185
R1607 GNDA.n1026 GNDA.n1000 185
R1608 GNDA.n1029 GNDA.n1028 185
R1609 GNDA.n1030 GNDA.n999 185
R1610 GNDA.n1032 GNDA.n1031 185
R1611 GNDA.n1034 GNDA.n998 185
R1612 GNDA.n1037 GNDA.n1036 185
R1613 GNDA.n1038 GNDA.n997 185
R1614 GNDA.n1040 GNDA.n1039 185
R1615 GNDA.n1058 GNDA.n992 185
R1616 GNDA.n1056 GNDA.n1055 185
R1617 GNDA.n1054 GNDA.n993 185
R1618 GNDA.n1053 GNDA.n1052 185
R1619 GNDA.n1050 GNDA.n994 185
R1620 GNDA.n1048 GNDA.n1047 185
R1621 GNDA.n1046 GNDA.n995 185
R1622 GNDA.n1045 GNDA.n1044 185
R1623 GNDA.n1042 GNDA.n996 185
R1624 GNDA.n1862 GNDA.n1861 185
R1625 GNDA.n1864 GNDA.n1863 185
R1626 GNDA.n1866 GNDA.n1860 185
R1627 GNDA.n1869 GNDA.n1868 185
R1628 GNDA.n1870 GNDA.n1859 185
R1629 GNDA.n1872 GNDA.n1871 185
R1630 GNDA.n1874 GNDA.n1858 185
R1631 GNDA.n1877 GNDA.n1876 185
R1632 GNDA.n1878 GNDA.n1857 185
R1633 GNDA.n1880 GNDA.n1879 185
R1634 GNDA.n1882 GNDA.n1856 185
R1635 GNDA.n1885 GNDA.n1884 185
R1636 GNDA.n1886 GNDA.n1855 185
R1637 GNDA.n1888 GNDA.n1887 185
R1638 GNDA.n1890 GNDA.n1854 185
R1639 GNDA.n1893 GNDA.n1892 185
R1640 GNDA.n1894 GNDA.n1853 185
R1641 GNDA.n1896 GNDA.n1895 185
R1642 GNDA.n1914 GNDA.n1848 185
R1643 GNDA.n1912 GNDA.n1911 185
R1644 GNDA.n1910 GNDA.n1849 185
R1645 GNDA.n1909 GNDA.n1908 185
R1646 GNDA.n1906 GNDA.n1850 185
R1647 GNDA.n1904 GNDA.n1903 185
R1648 GNDA.n1902 GNDA.n1851 185
R1649 GNDA.n1901 GNDA.n1900 185
R1650 GNDA.n1898 GNDA.n1852 185
R1651 GNDA.n1916 GNDA.n1915 185
R1652 GNDA.n305 GNDA.n303 185
R1653 GNDA.n1923 GNDA.n1922 185
R1654 GNDA.n1925 GNDA.n302 185
R1655 GNDA.n1927 GNDA.n1926 185
R1656 GNDA.n296 GNDA.n294 185
R1657 GNDA.n1934 GNDA.n1933 185
R1658 GNDA.n1936 GNDA.n293 185
R1659 GNDA.n1938 GNDA.n1937 185
R1660 GNDA.n1060 GNDA.n1059 185
R1661 GNDA.n978 GNDA.n976 185
R1662 GNDA.n1067 GNDA.n1066 185
R1663 GNDA.n1069 GNDA.n975 185
R1664 GNDA.n1071 GNDA.n1070 185
R1665 GNDA.n969 GNDA.n967 185
R1666 GNDA.n1078 GNDA.n1077 185
R1667 GNDA.n1080 GNDA.n966 185
R1668 GNDA.n1082 GNDA.n1081 185
R1669 GNDA.n1270 GNDA.n1269 185
R1670 GNDA.n1190 GNDA.n1188 185
R1671 GNDA.n1277 GNDA.n1276 185
R1672 GNDA.n1279 GNDA.n1187 185
R1673 GNDA.n1281 GNDA.n1280 185
R1674 GNDA.n1182 GNDA.n1181 185
R1675 GNDA.n1288 GNDA.n1287 185
R1676 GNDA.n1291 GNDA.n1290 185
R1677 GNDA.n1180 GNDA.n1177 185
R1678 GNDA.n607 GNDA.n606 185
R1679 GNDA.n609 GNDA.n608 185
R1680 GNDA.n611 GNDA.n605 185
R1681 GNDA.n614 GNDA.n613 185
R1682 GNDA.n615 GNDA.n604 185
R1683 GNDA.n617 GNDA.n616 185
R1684 GNDA.n619 GNDA.n603 185
R1685 GNDA.n622 GNDA.n621 185
R1686 GNDA.n623 GNDA.n602 185
R1687 GNDA.n625 GNDA.n624 185
R1688 GNDA.n627 GNDA.n601 185
R1689 GNDA.n630 GNDA.n629 185
R1690 GNDA.n631 GNDA.n600 185
R1691 GNDA.n633 GNDA.n632 185
R1692 GNDA.n635 GNDA.n599 185
R1693 GNDA.n638 GNDA.n637 185
R1694 GNDA.n639 GNDA.n598 185
R1695 GNDA.n641 GNDA.n640 185
R1696 GNDA.n659 GNDA.n593 185
R1697 GNDA.n657 GNDA.n656 185
R1698 GNDA.n655 GNDA.n594 185
R1699 GNDA.n654 GNDA.n653 185
R1700 GNDA.n651 GNDA.n595 185
R1701 GNDA.n649 GNDA.n648 185
R1702 GNDA.n647 GNDA.n596 185
R1703 GNDA.n646 GNDA.n645 185
R1704 GNDA.n643 GNDA.n597 185
R1705 GNDA.n1454 GNDA.n1453 185
R1706 GNDA.n1456 GNDA.n1455 185
R1707 GNDA.n1458 GNDA.n1452 185
R1708 GNDA.n1461 GNDA.n1460 185
R1709 GNDA.n1462 GNDA.n1451 185
R1710 GNDA.n1464 GNDA.n1463 185
R1711 GNDA.n1466 GNDA.n1450 185
R1712 GNDA.n1469 GNDA.n1468 185
R1713 GNDA.n1470 GNDA.n1449 185
R1714 GNDA.n1472 GNDA.n1471 185
R1715 GNDA.n1474 GNDA.n1448 185
R1716 GNDA.n1477 GNDA.n1476 185
R1717 GNDA.n1478 GNDA.n1447 185
R1718 GNDA.n1480 GNDA.n1479 185
R1719 GNDA.n1482 GNDA.n1446 185
R1720 GNDA.n1485 GNDA.n1484 185
R1721 GNDA.n1486 GNDA.n1445 185
R1722 GNDA.n1488 GNDA.n1487 185
R1723 GNDA.n1506 GNDA.n1440 185
R1724 GNDA.n1504 GNDA.n1503 185
R1725 GNDA.n1502 GNDA.n1441 185
R1726 GNDA.n1501 GNDA.n1500 185
R1727 GNDA.n1498 GNDA.n1442 185
R1728 GNDA.n1496 GNDA.n1495 185
R1729 GNDA.n1494 GNDA.n1443 185
R1730 GNDA.n1493 GNDA.n1492 185
R1731 GNDA.n1490 GNDA.n1444 185
R1732 GNDA.n2018 GNDA.n243 185
R1733 GNDA.n2017 GNDA.n2016 185
R1734 GNDA.n2015 GNDA.n2014 185
R1735 GNDA.n2013 GNDA.n2012 185
R1736 GNDA.n2011 GNDA.n2010 185
R1737 GNDA.n2009 GNDA.n2008 185
R1738 GNDA.n2007 GNDA.n2006 185
R1739 GNDA.n2005 GNDA.n2004 185
R1740 GNDA.n2003 GNDA.n2002 185
R1741 GNDA.n2001 GNDA.n2000 185
R1742 GNDA.n1999 GNDA.n1998 185
R1743 GNDA.n1997 GNDA.n1996 185
R1744 GNDA.n1995 GNDA.n1994 185
R1745 GNDA.n1993 GNDA.n1992 185
R1746 GNDA.n1991 GNDA.n1990 185
R1747 GNDA.n1989 GNDA.n1988 185
R1748 GNDA.n1987 GNDA.n1986 185
R1749 GNDA.n1985 GNDA.n1984 185
R1750 GNDA.n2060 GNDA.n2059 185
R1751 GNDA.n226 GNDA.n224 185
R1752 GNDA.n1971 GNDA.n1970 185
R1753 GNDA.n1973 GNDA.n1972 185
R1754 GNDA.n1975 GNDA.n1974 185
R1755 GNDA.n1977 GNDA.n1976 185
R1756 GNDA.n1979 GNDA.n1978 185
R1757 GNDA.n1981 GNDA.n1980 185
R1758 GNDA.n1983 GNDA.n1982 185
R1759 GNDA.n225 GNDA.n223 185
R1760 GNDA.n2037 GNDA.n2036 185
R1761 GNDA.n2039 GNDA.n2038 185
R1762 GNDA.n2033 GNDA.n2032 185
R1763 GNDA.n2031 GNDA.n2026 185
R1764 GNDA.n2047 GNDA.n2046 185
R1765 GNDA.n2049 GNDA.n2048 185
R1766 GNDA.n246 GNDA.n244 185
R1767 GNDA.n2056 GNDA.n2055 185
R1768 GNDA.n1508 GNDA.n1507 185
R1769 GNDA.n878 GNDA.n876 185
R1770 GNDA.n1515 GNDA.n1514 185
R1771 GNDA.n1517 GNDA.n875 185
R1772 GNDA.n1519 GNDA.n1518 185
R1773 GNDA.n869 GNDA.n867 185
R1774 GNDA.n1526 GNDA.n1525 185
R1775 GNDA.n1528 GNDA.n866 185
R1776 GNDA.n1530 GNDA.n1529 185
R1777 GNDA.n661 GNDA.n660 185
R1778 GNDA.n584 GNDA.n582 185
R1779 GNDA.n668 GNDA.n667 185
R1780 GNDA.n670 GNDA.n581 185
R1781 GNDA.n672 GNDA.n671 185
R1782 GNDA.n575 GNDA.n573 185
R1783 GNDA.n679 GNDA.n678 185
R1784 GNDA.n681 GNDA.n572 185
R1785 GNDA.n683 GNDA.n682 185
R1786 GNDA.n2329 GNDA.n2327 182.4
R1787 GNDA.n2259 GNDA.n2258 182.4
R1788 GNDA.n2432 GNDA.n2431 179.363
R1789 GNDA.n2481 GNDA.n43 176.543
R1790 GNDA.n2482 GNDA.n2481 176.543
R1791 GNDA.n2195 GNDA.n78 176
R1792 GNDA.n2195 GNDA.n2194 176
R1793 GNDA.n2368 GNDA.n2324 176
R1794 GNDA.n2461 GNDA.n2253 176
R1795 GNDA.n52 GNDA.t350 175.864
R1796 GNDA.n1366 GNDA.n1364 175.546
R1797 GNDA.n1370 GNDA.n1125 175.546
R1798 GNDA.n1374 GNDA.n1372 175.546
R1799 GNDA.n1378 GNDA.n1123 175.546
R1800 GNDA.n1381 GNDA.n1380 175.546
R1801 GNDA.n1358 GNDA.n1129 175.546
R1802 GNDA.n1354 GNDA.n1129 175.546
R1803 GNDA.n1354 GNDA.n1343 175.546
R1804 GNDA.n1350 GNDA.n1343 175.546
R1805 GNDA.n1350 GNDA.n1346 175.546
R1806 GNDA.n1346 GNDA.n351 175.546
R1807 GNDA.n1756 GNDA.n351 175.546
R1808 GNDA.n1756 GNDA.n352 175.546
R1809 GNDA.n1752 GNDA.n352 175.546
R1810 GNDA.n1752 GNDA.n354 175.546
R1811 GNDA.n685 GNDA.n568 175.546
R1812 GNDA.n676 GNDA.n577 175.546
R1813 GNDA.n674 GNDA.n578 175.546
R1814 GNDA.n665 GNDA.n586 175.546
R1815 GNDA.n663 GNDA.n589 175.546
R1816 GNDA.n1118 GNDA.n1117 175.546
R1817 GNDA.n1114 GNDA.n1113 175.546
R1818 GNDA.n1110 GNDA.n1109 175.546
R1819 GNDA.n1106 GNDA.n1105 175.546
R1820 GNDA.n1693 GNDA.n411 175.546
R1821 GNDA.n1790 GNDA.n326 175.546
R1822 GNDA.n1794 GNDA.n326 175.546
R1823 GNDA.n1794 GNDA.n324 175.546
R1824 GNDA.n1798 GNDA.n324 175.546
R1825 GNDA.n1798 GNDA.n321 175.546
R1826 GNDA.n1830 GNDA.n321 175.546
R1827 GNDA.n1830 GNDA.n322 175.546
R1828 GNDA.n1826 GNDA.n322 175.546
R1829 GNDA.n1826 GNDA.n1802 175.546
R1830 GNDA.n1822 GNDA.n1802 175.546
R1831 GNDA.n1822 GNDA.n1804 175.546
R1832 GNDA.n1818 GNDA.n1806 175.546
R1833 GNDA.n1814 GNDA.n1806 175.546
R1834 GNDA.n1814 GNDA.n1808 175.546
R1835 GNDA.n1810 GNDA.n1808 175.546
R1836 GNDA.n1810 GNDA.n317 175.546
R1837 GNDA.n1833 GNDA.n317 175.546
R1838 GNDA.n1833 GNDA.n315 175.546
R1839 GNDA.n1838 GNDA.n315 175.546
R1840 GNDA.n1838 GNDA.n313 175.546
R1841 GNDA.n1842 GNDA.n313 175.546
R1842 GNDA.n1940 GNDA.n289 175.546
R1843 GNDA.n1931 GNDA.n298 175.546
R1844 GNDA.n1929 GNDA.n299 175.546
R1845 GNDA.n1920 GNDA.n307 175.546
R1846 GNDA.n1918 GNDA.n308 175.546
R1847 GNDA.n1157 GNDA.n1145 175.546
R1848 GNDA.n1157 GNDA.n1148 175.546
R1849 GNDA.n1153 GNDA.n1148 175.546
R1850 GNDA.n1153 GNDA.n1150 175.546
R1851 GNDA.n1150 GNDA.n379 175.546
R1852 GNDA.n1721 GNDA.n379 175.546
R1853 GNDA.n1721 GNDA.n380 175.546
R1854 GNDA.n1717 GNDA.n380 175.546
R1855 GNDA.n1717 GNDA.n383 175.546
R1856 GNDA.n1713 GNDA.n383 175.546
R1857 GNDA.n1713 GNDA.n385 175.546
R1858 GNDA.n1320 GNDA.n1146 175.546
R1859 GNDA.n1320 GNDA.n1161 175.546
R1860 GNDA.n1316 GNDA.n1161 175.546
R1861 GNDA.n1316 GNDA.n1165 175.546
R1862 GNDA.n1312 GNDA.n1165 175.546
R1863 GNDA.n1312 GNDA.n1167 175.546
R1864 GNDA.n1308 GNDA.n1167 175.546
R1865 GNDA.n1308 GNDA.n1169 175.546
R1866 GNDA.n1304 GNDA.n1169 175.546
R1867 GNDA.n1304 GNDA.n1303 175.546
R1868 GNDA.n1294 GNDA.n1293 175.546
R1869 GNDA.n1285 GNDA.n1183 175.546
R1870 GNDA.n1283 GNDA.n1184 175.546
R1871 GNDA.n1274 GNDA.n1192 175.546
R1872 GNDA.n1272 GNDA.n1193 175.546
R1873 GNDA.n938 GNDA.n937 175.546
R1874 GNDA.n944 GNDA.n943 175.546
R1875 GNDA.n950 GNDA.n949 175.546
R1876 GNDA.n956 GNDA.n955 175.546
R1877 GNDA.n958 GNDA.n410 175.546
R1878 GNDA.n1391 GNDA.n933 175.546
R1879 GNDA.n1395 GNDA.n1393 175.546
R1880 GNDA.n1399 GNDA.n931 175.546
R1881 GNDA.n1403 GNDA.n1401 175.546
R1882 GNDA.n1407 GNDA.n929 175.546
R1883 GNDA.n1097 GNDA.n1096 175.546
R1884 GNDA.n1099 GNDA.n1098 175.546
R1885 GNDA.n1101 GNDA.n1100 175.546
R1886 GNDA.n1103 GNDA.n1102 175.546
R1887 GNDA.n1688 GNDA.n417 175.546
R1888 GNDA.n1532 GNDA.n862 175.546
R1889 GNDA.n1523 GNDA.n871 175.546
R1890 GNDA.n1521 GNDA.n872 175.546
R1891 GNDA.n1512 GNDA.n880 175.546
R1892 GNDA.n1510 GNDA.n881 175.546
R1893 GNDA.n1417 GNDA.n894 175.546
R1894 GNDA.n1421 GNDA.n1419 175.546
R1895 GNDA.n1427 GNDA.n890 175.546
R1896 GNDA.n1430 GNDA.n1429 175.546
R1897 GNDA.n1434 GNDA.n1433 175.546
R1898 GNDA.n2053 GNDA.n2023 175.546
R1899 GNDA.n2051 GNDA.n2024 175.546
R1900 GNDA.n2044 GNDA.n2043 175.546
R1901 GNDA.n2041 GNDA.n2030 175.546
R1902 GNDA.n2063 GNDA.n222 175.546
R1903 GNDA.n2087 GNDA.n209 175.546
R1904 GNDA.n2083 GNDA.n209 175.546
R1905 GNDA.n2083 GNDA.n212 175.546
R1906 GNDA.n2079 GNDA.n212 175.546
R1907 GNDA.n2079 GNDA.n214 175.546
R1908 GNDA.n2075 GNDA.n214 175.546
R1909 GNDA.n2075 GNDA.n216 175.546
R1910 GNDA.n2071 GNDA.n216 175.546
R1911 GNDA.n2071 GNDA.n218 175.546
R1912 GNDA.n221 GNDA.n218 175.546
R1913 GNDA.n922 GNDA.n921 175.546
R1914 GNDA.n919 GNDA.n900 175.546
R1915 GNDA.n915 GNDA.n914 175.546
R1916 GNDA.n912 GNDA.n903 175.546
R1917 GNDA.n908 GNDA.n907 175.546
R1918 GNDA.n1704 GNDA.n388 175.546
R1919 GNDA.n1704 GNDA.n1697 175.546
R1920 GNDA.n1700 GNDA.n1697 175.546
R1921 GNDA.n1700 GNDA.n333 175.546
R1922 GNDA.n1771 GNDA.n333 175.546
R1923 GNDA.n1772 GNDA.n1771 175.546
R1924 GNDA.n1775 GNDA.n1772 175.546
R1925 GNDA.n1775 GNDA.n331 175.546
R1926 GNDA.n1779 GNDA.n331 175.546
R1927 GNDA.n1779 GNDA.n328 175.546
R1928 GNDA.n1783 GNDA.n328 175.546
R1929 GNDA.n1084 GNDA.n963 175.546
R1930 GNDA.n1075 GNDA.n971 175.546
R1931 GNDA.n1073 GNDA.n972 175.546
R1932 GNDA.n1064 GNDA.n980 175.546
R1933 GNDA.n1062 GNDA.n981 175.546
R1934 GNDA.n1961 GNDA.n1960 175.546
R1935 GNDA.n1958 GNDA.n274 175.546
R1936 GNDA.n1954 GNDA.n1953 175.546
R1937 GNDA.n1951 GNDA.n281 175.546
R1938 GNDA.n986 GNDA.n285 175.546
R1939 GNDA.n1543 GNDA.n509 175.546
R1940 GNDA.n1547 GNDA.n1545 175.546
R1941 GNDA.n1551 GNDA.n507 175.546
R1942 GNDA.n1555 GNDA.n1553 175.546
R1943 GNDA.n1559 GNDA.n505 175.546
R1944 GNDA.n1564 GNDA.n1562 175.546
R1945 GNDA.n1570 GNDA.n467 175.546
R1946 GNDA.n1574 GNDA.n1572 175.546
R1947 GNDA.n1580 GNDA.n463 175.546
R1948 GNDA.n1584 GNDA.n1582 175.546
R1949 GNDA.n1681 GNDA.n1680 175.546
R1950 GNDA.n444 GNDA.n443 175.546
R1951 GNDA.n1671 GNDA.n1670 175.546
R1952 GNDA.n452 GNDA.n451 175.546
R1953 GNDA.n1661 GNDA.n1660 175.546
R1954 GNDA.n455 GNDA.n99 175.546
R1955 GNDA.n510 GNDA.n430 175.546
R1956 GNDA.n512 GNDA.n511 175.546
R1957 GNDA.n514 GNDA.n513 175.546
R1958 GNDA.n516 GNDA.n515 175.546
R1959 GNDA.n518 GNDA.n517 175.546
R1960 GNDA.n498 GNDA.n497 175.546
R1961 GNDA.n494 GNDA.n493 175.546
R1962 GNDA.n491 GNDA.n475 175.546
R1963 GNDA.n487 GNDA.n485 175.546
R1964 GNDA.n483 GNDA.n477 175.546
R1965 GNDA.n2091 GNDA.n199 175.546
R1966 GNDA.n2091 GNDA.n197 175.546
R1967 GNDA.n2096 GNDA.n197 175.546
R1968 GNDA.n2096 GNDA.n194 175.546
R1969 GNDA.n2100 GNDA.n194 175.546
R1970 GNDA.n2101 GNDA.n2100 175.546
R1971 GNDA.n2105 GNDA.n2101 175.546
R1972 GNDA.n2105 GNDA.n192 175.546
R1973 GNDA.n2109 GNDA.n192 175.546
R1974 GNDA.n2110 GNDA.n2109 175.546
R1975 GNDA.n2145 GNDA.n2144 175.546
R1976 GNDA.n2136 GNDA.n2135 175.546
R1977 GNDA.n2132 GNDA.n2131 175.546
R1978 GNDA.n2123 GNDA.n2122 175.546
R1979 GNDA.n2119 GNDA.n2118 175.546
R1980 GNDA.n469 GNDA.n257 175.546
R1981 GNDA.n1568 GNDA.n1567 175.546
R1982 GNDA.n466 GNDA.n465 175.546
R1983 GNDA.n1578 GNDA.n1577 175.546
R1984 GNDA.n462 GNDA.n461 175.546
R1985 GNDA.n753 GNDA.n693 175.546
R1986 GNDA.n753 GNDA.n724 175.546
R1987 GNDA.n749 GNDA.n724 175.546
R1988 GNDA.n749 GNDA.n726 175.546
R1989 GNDA.n745 GNDA.n726 175.546
R1990 GNDA.n745 GNDA.n728 175.546
R1991 GNDA.n741 GNDA.n728 175.546
R1992 GNDA.n741 GNDA.n730 175.546
R1993 GNDA.n737 GNDA.n730 175.546
R1994 GNDA.n737 GNDA.n733 175.546
R1995 GNDA.n769 GNDA.n363 175.546
R1996 GNDA.n1733 GNDA.n363 175.546
R1997 GNDA.n1733 GNDA.n364 175.546
R1998 GNDA.n1725 GNDA.n364 175.546
R1999 GNDA.n1725 GNDA.n370 175.546
R2000 GNDA.n533 GNDA.n370 175.546
R2001 GNDA.n535 GNDA.n533 175.546
R2002 GNDA.n535 GNDA.n522 175.546
R2003 GNDA.n829 GNDA.n522 175.546
R2004 GNDA.n829 GNDA.n520 175.546
R2005 GNDA.n833 GNDA.n520 175.546
R2006 GNDA.n854 GNDA.n409 175.546
R2007 GNDA.n852 GNDA.n851 175.546
R2008 GNDA.n848 GNDA.n847 175.546
R2009 GNDA.n844 GNDA.n843 175.546
R2010 GNDA.n840 GNDA.n839 175.546
R2011 GNDA.n720 GNDA.n719 175.546
R2012 GNDA.n717 GNDA.n696 175.546
R2013 GNDA.n713 GNDA.n712 175.546
R2014 GNDA.n710 GNDA.n699 175.546
R2015 GNDA.n706 GNDA.n705 175.546
R2016 GNDA.n1963 GNDA.n269 175.546
R2017 GNDA.n276 GNDA.n275 175.546
R2018 GNDA.n278 GNDA.n277 175.546
R2019 GNDA.n283 GNDA.n282 175.546
R2020 GNDA.n1947 GNDA.n1946 175.546
R2021 GNDA.n1415 GNDA.n1414 175.546
R2022 GNDA.n893 GNDA.n892 175.546
R2023 GNDA.n1425 GNDA.n1424 175.546
R2024 GNDA.n889 GNDA.n888 175.546
R2025 GNDA.n1967 GNDA.n250 175.546
R2026 GNDA.n936 GNDA.n935 175.546
R2027 GNDA.n942 GNDA.n941 175.546
R2028 GNDA.n948 GNDA.n947 175.546
R2029 GNDA.n954 GNDA.n953 175.546
R2030 GNDA.n1090 GNDA.n1089 175.546
R2031 GNDA.n2159 GNDA.n2158 175.5
R2032 GNDA.n962 GNDA.t137 172.876
R2033 GNDA.n861 GNDA.t137 172.876
R2034 GNDA.n928 GNDA.t137 172.615
R2035 GNDA.n504 GNDA.t137 172.615
R2036 GNDA.n2431 GNDA.n2430 171.817
R2037 GNDA.n2207 GNDA.n53 169.232
R2038 GNDA.n2433 GNDA.n2432 164.906
R2039 GNDA.t135 GNDA.n377 162.964
R2040 GNDA.t137 GNDA.n319 162.964
R2041 GNDA.n77 GNDA.t185 160.725
R2042 GNDA.n79 GNDA.t124 160.725
R2043 GNDA.n2190 GNDA.t164 160.725
R2044 GNDA.n62 GNDA.t161 160.725
R2045 GNDA.n2153 GNDA.t158 160.725
R2046 GNDA.n81 GNDA.t188 160.725
R2047 GNDA.n18 GNDA.n17 160
R2048 GNDA.n2494 GNDA.n10 160
R2049 GNDA.n29 GNDA.n28 160
R2050 GNDA.n2331 GNDA.n2317 160
R2051 GNDA.n2459 GNDA.n2261 160
R2052 GNDA.n340 GNDA.t257 157.555
R2053 GNDA.n341 GNDA.t256 157.555
R2054 GNDA.n2448 GNDA.n2447 156.8
R2055 GNDA.n2439 GNDA.n2438 153.601
R2056 GNDA.n34 GNDA.n33 153.601
R2057 GNDA.n2232 GNDA.t32 153.294
R2058 GNDA.n2323 GNDA.t155 152.994
R2059 GNDA.n2325 GNDA.t143 152.994
R2060 GNDA.n2256 GNDA.t169 152.994
R2061 GNDA.n2252 GNDA.t152 152.994
R2062 GNDA.n1583 GNDA.n459 152.643
R2063 GNDA.n436 GNDA.n435 152.643
R2064 GNDA.n263 GNDA.n262 152.643
R2065 GNDA.n835 GNDA.n404 152.643
R2066 GNDA.n2205 GNDA.n2204 150.938
R2067 GNDA.n2436 GNDA.n2435 150.4
R2068 GNDA.n2445 GNDA.n2444 150.4
R2069 GNDA.n1730 GNDA.n367 150
R2070 GNDA.n1728 GNDA.n368 150
R2071 GNDA.n530 GNDA.n529 150
R2072 GNDA.n540 GNDA.n539 150
R2073 GNDA.n811 GNDA.n809 150
R2074 GNDA.n815 GNDA.n545 150
R2075 GNDA.n819 GNDA.n817 150
R2076 GNDA.n823 GNDA.n543 150
R2077 GNDA.n795 GNDA.n793 150
R2078 GNDA.n799 GNDA.n549 150
R2079 GNDA.n803 GNDA.n801 150
R2080 GNDA.n807 GNDA.n547 150
R2081 GNDA.n787 GNDA.n785 150
R2082 GNDA.n783 GNDA.n553 150
R2083 GNDA.n779 GNDA.n777 150
R2084 GNDA.n775 GNDA.n556 150
R2085 GNDA.n1677 GNDA.n1676 150
R2086 GNDA.n1674 GNDA.n442 150
R2087 GNDA.n1667 GNDA.n1666 150
R2088 GNDA.n1664 GNDA.n450 150
R2089 GNDA.n1642 GNDA.n1640 150
R2090 GNDA.n1646 GNDA.n1593 150
R2091 GNDA.n1650 GNDA.n1648 150
R2092 GNDA.n1654 GNDA.n1591 150
R2093 GNDA.n1626 GNDA.n1624 150
R2094 GNDA.n1630 GNDA.n1597 150
R2095 GNDA.n1634 GNDA.n1632 150
R2096 GNDA.n1638 GNDA.n1595 150
R2097 GNDA.n1618 GNDA.n1616 150
R2098 GNDA.n1614 GNDA.n1601 150
R2099 GNDA.n1610 GNDA.n1608 150
R2100 GNDA.n1606 GNDA.n1603 150
R2101 GNDA.n2141 GNDA.n112 150
R2102 GNDA.n2139 GNDA.n113 150
R2103 GNDA.n2128 GNDA.n117 150
R2104 GNDA.n2126 GNDA.n118 150
R2105 GNDA.n174 GNDA.n126 150
R2106 GNDA.n178 GNDA.n176 150
R2107 GNDA.n182 GNDA.n124 150
R2108 GNDA.n185 GNDA.n184 150
R2109 GNDA.n158 GNDA.n130 150
R2110 GNDA.n162 GNDA.n160 150
R2111 GNDA.n166 GNDA.n128 150
R2112 GNDA.n170 GNDA.n168 150
R2113 GNDA.n150 GNDA.n132 150
R2114 GNDA.n146 GNDA.n144 150
R2115 GNDA.n142 GNDA.n134 150
R2116 GNDA.n138 GNDA.n136 150
R2117 GNDA.n1290 GNDA.n1180 150
R2118 GNDA.n1288 GNDA.n1181 150
R2119 GNDA.n1280 GNDA.n1279 150
R2120 GNDA.n1277 GNDA.n1188 150
R2121 GNDA.n1254 GNDA.n1252 150
R2122 GNDA.n1258 GNDA.n1205 150
R2123 GNDA.n1262 GNDA.n1260 150
R2124 GNDA.n1266 GNDA.n1203 150
R2125 GNDA.n1238 GNDA.n1236 150
R2126 GNDA.n1242 GNDA.n1209 150
R2127 GNDA.n1246 GNDA.n1244 150
R2128 GNDA.n1250 GNDA.n1207 150
R2129 GNDA.n1230 GNDA.n1228 150
R2130 GNDA.n1226 GNDA.n1213 150
R2131 GNDA.n1222 GNDA.n1220 150
R2132 GNDA.n1218 GNDA.n1216 150
R2133 GNDA.n1081 GNDA.n1080 150
R2134 GNDA.n1078 GNDA.n967 150
R2135 GNDA.n1070 GNDA.n1069 150
R2136 GNDA.n1067 GNDA.n976 150
R2137 GNDA.n1044 GNDA.n1042 150
R2138 GNDA.n1048 GNDA.n995 150
R2139 GNDA.n1052 GNDA.n1050 150
R2140 GNDA.n1056 GNDA.n993 150
R2141 GNDA.n1028 GNDA.n1026 150
R2142 GNDA.n1032 GNDA.n999 150
R2143 GNDA.n1036 GNDA.n1034 150
R2144 GNDA.n1040 GNDA.n997 150
R2145 GNDA.n1020 GNDA.n1018 150
R2146 GNDA.n1016 GNDA.n1003 150
R2147 GNDA.n1012 GNDA.n1010 150
R2148 GNDA.n1008 GNDA.n1005 150
R2149 GNDA.n1937 GNDA.n1936 150
R2150 GNDA.n1934 GNDA.n294 150
R2151 GNDA.n1926 GNDA.n1925 150
R2152 GNDA.n1923 GNDA.n303 150
R2153 GNDA.n1900 GNDA.n1898 150
R2154 GNDA.n1904 GNDA.n1851 150
R2155 GNDA.n1908 GNDA.n1906 150
R2156 GNDA.n1912 GNDA.n1849 150
R2157 GNDA.n1884 GNDA.n1882 150
R2158 GNDA.n1888 GNDA.n1855 150
R2159 GNDA.n1892 GNDA.n1890 150
R2160 GNDA.n1896 GNDA.n1853 150
R2161 GNDA.n1876 GNDA.n1874 150
R2162 GNDA.n1872 GNDA.n1859 150
R2163 GNDA.n1868 GNDA.n1866 150
R2164 GNDA.n1864 GNDA.n1861 150
R2165 GNDA.n682 GNDA.n681 150
R2166 GNDA.n679 GNDA.n573 150
R2167 GNDA.n671 GNDA.n670 150
R2168 GNDA.n668 GNDA.n582 150
R2169 GNDA.n645 GNDA.n643 150
R2170 GNDA.n649 GNDA.n596 150
R2171 GNDA.n653 GNDA.n651 150
R2172 GNDA.n657 GNDA.n594 150
R2173 GNDA.n629 GNDA.n627 150
R2174 GNDA.n633 GNDA.n600 150
R2175 GNDA.n637 GNDA.n635 150
R2176 GNDA.n641 GNDA.n598 150
R2177 GNDA.n621 GNDA.n619 150
R2178 GNDA.n617 GNDA.n604 150
R2179 GNDA.n613 GNDA.n611 150
R2180 GNDA.n609 GNDA.n606 150
R2181 GNDA.n1529 GNDA.n1528 150
R2182 GNDA.n1526 GNDA.n867 150
R2183 GNDA.n1518 GNDA.n1517 150
R2184 GNDA.n1515 GNDA.n876 150
R2185 GNDA.n1492 GNDA.n1490 150
R2186 GNDA.n1496 GNDA.n1443 150
R2187 GNDA.n1500 GNDA.n1498 150
R2188 GNDA.n1504 GNDA.n1441 150
R2189 GNDA.n1476 GNDA.n1474 150
R2190 GNDA.n1480 GNDA.n1447 150
R2191 GNDA.n1484 GNDA.n1482 150
R2192 GNDA.n1488 GNDA.n1445 150
R2193 GNDA.n1468 GNDA.n1466 150
R2194 GNDA.n1464 GNDA.n1451 150
R2195 GNDA.n1460 GNDA.n1458 150
R2196 GNDA.n1456 GNDA.n1453 150
R2197 GNDA.n2056 GNDA.n244 150
R2198 GNDA.n2048 GNDA.n2047 150
R2199 GNDA.n2032 GNDA.n2031 150
R2200 GNDA.n2038 GNDA.n2037 150
R2201 GNDA.n1982 GNDA.n1981 150
R2202 GNDA.n1978 GNDA.n1977 150
R2203 GNDA.n1974 GNDA.n1973 150
R2204 GNDA.n1970 GNDA.n226 150
R2205 GNDA.n1998 GNDA.n1997 150
R2206 GNDA.n1994 GNDA.n1993 150
R2207 GNDA.n1990 GNDA.n1989 150
R2208 GNDA.n1986 GNDA.n1985 150
R2209 GNDA.n2006 GNDA.n2005 150
R2210 GNDA.n2010 GNDA.n2009 150
R2211 GNDA.n2014 GNDA.n2013 150
R2212 GNDA.n2016 GNDA.n243 150
R2213 GNDA.n338 GNDA.t251 148.906
R2214 GNDA.n338 GNDA.t242 148.653
R2215 GNDA.n768 GNDA.n360 145.013
R2216 GNDA.n2214 GNDA.n2212 139.639
R2217 GNDA.n2230 GNDA.n2229 139.077
R2218 GNDA.n2228 GNDA.n2227 139.077
R2219 GNDA.n2226 GNDA.n2225 139.077
R2220 GNDA.n2224 GNDA.n2223 139.077
R2221 GNDA.n2222 GNDA.n2221 139.077
R2222 GNDA.n2220 GNDA.n2219 139.077
R2223 GNDA.n2218 GNDA.n2217 139.077
R2224 GNDA.n2216 GNDA.n2215 139.077
R2225 GNDA.n2214 GNDA.n2213 139.077
R2226 GNDA.n2239 GNDA.n53 131.625
R2227 GNDA.t142 GNDA.n2311 130.731
R2228 GNDA.t168 GNDA.n2455 130.731
R2229 GNDA.n2452 GNDA.n2451 127.249
R2230 GNDA.n2160 GNDA.n2159 125.356
R2231 GNDA.n1362 GNDA.n1127 124.832
R2232 GNDA.n688 GNDA.n687 124.832
R2233 GNDA.n1790 GNDA.n1787 124.832
R2234 GNDA.n1943 GNDA.n1942 124.832
R2235 GNDA.n1324 GNDA.n1145 124.832
R2236 GNDA.n1299 GNDA.n1298 124.832
R2237 GNDA.n1387 GNDA.n858 124.832
R2238 GNDA.n1535 GNDA.n1534 124.832
R2239 GNDA.n2021 GNDA.n247 124.832
R2240 GNDA.n924 GNDA.n898 124.832
R2241 GNDA.n1708 GNDA.n388 124.832
R2242 GNDA.n1086 GNDA.n859 124.832
R2243 GNDA.n1539 GNDA.n1537 124.832
R2244 GNDA.n500 GNDA.n472 124.832
R2245 GNDA.n2150 GNDA.n106 124.832
R2246 GNDA.n769 GNDA.n767 124.832
R2247 GNDA.n757 GNDA.n692 124.832
R2248 GNDA.n2371 GNDA.n2370 119.525
R2249 GNDA.n2463 GNDA.n2249 119.525
R2250 GNDA.n2210 GNDA.n63 118.4
R2251 GNDA.n2192 GNDA.n2191 118.4
R2252 GNDA.n2194 GNDA.n2193 118.4
R2253 GNDA.n2179 GNDA.n78 118.4
R2254 GNDA.n2155 GNDA.n2154 118.4
R2255 GNDA.n2178 GNDA.n82 118.4
R2256 GNDA.n9 GNDA.t216 113.974
R2257 GNDA.n13 GNDA.t178 113.974
R2258 GNDA.n12 GNDA.t213 113.974
R2259 GNDA.n11 GNDA.t198 113.974
R2260 GNDA.n30 GNDA.t219 113.974
R2261 GNDA.n31 GNDA.t204 113.974
R2262 GNDA.n21 GNDA.t191 113.974
R2263 GNDA.n19 GNDA.t133 113.974
R2264 GNDA.n26 GNDA.t121 113.974
R2265 GNDA.n25 GNDA.t210 113.974
R2266 GNDA.n1723 GNDA.t135 113.624
R2267 GNDA.n1769 GNDA.t137 112.388
R2268 GNDA.n2286 GNDA.n2280 108.8
R2269 GNDA.n2298 GNDA.n2277 108.8
R2270 GNDA.n765 GNDA.n360 108.522
R2271 GNDA.n1965 GNDA.n0 14.555
R2272 GNDA.n2450 GNDA.t209 101.194
R2273 GNDA.n1695 GNDA.n1694 99.6276
R2274 GNDA.n2396 GNDA.n2395 99.0842
R2275 GNDA.n2400 GNDA.n2399 99.0842
R2276 GNDA.n2402 GNDA.n2401 99.0842
R2277 GNDA.n2404 GNDA.n2403 99.0842
R2278 GNDA.n2406 GNDA.n2405 99.0842
R2279 GNDA.n2408 GNDA.n2407 99.0842
R2280 GNDA.n2410 GNDA.n2409 99.0842
R2281 GNDA.n2412 GNDA.n2411 99.0842
R2282 GNDA.n2414 GNDA.n2413 99.0842
R2283 GNDA.n2416 GNDA.n2415 99.0842
R2284 GNDA.n2418 GNDA.n2417 99.0842
R2285 GNDA.n2420 GNDA.n2419 99.0842
R2286 GNDA.t270 GNDA.n2241 97.1515
R2287 GNDA.n2465 GNDA.t9 97.1515
R2288 GNDA.n2426 GNDA.n2425 95.101
R2289 GNDA.n2378 GNDA.n2374 95.101
R2290 GNDA.t207 GNDA.n2308 94.8842
R2291 GNDA.n2309 GNDA.t174 94.8842
R2292 GNDA.t140 GNDA.n2270 94.8842
R2293 GNDA.n2271 GNDA.t127 94.8842
R2294 GNDA.n2380 GNDA.n2379 94.601
R2295 GNDA.n2424 GNDA.n2423 94.601
R2296 GNDA.n2471 GNDA.n2243 94.0176
R2297 GNDA.n1817 GNDA.n1816 91.8159
R2298 GNDA.n1816 GNDA.n1815 91.8159
R2299 GNDA.n1815 GNDA.n1807 91.8159
R2300 GNDA.n1809 GNDA.n1807 91.8159
R2301 GNDA.n1809 GNDA.n318 91.8159
R2302 GNDA.n1832 GNDA.n314 91.8159
R2303 GNDA.n1839 GNDA.n314 91.8159
R2304 GNDA.n1840 GNDA.n1839 91.8159
R2305 GNDA.n1841 GNDA.n1840 91.8159
R2306 GNDA.n1841 GNDA.n206 91.8159
R2307 GNDA.n2088 GNDA.n207 91.8159
R2308 GNDA.n2082 GNDA.n207 91.8159
R2309 GNDA.n2082 GNDA.n2081 91.8159
R2310 GNDA.n2081 GNDA.n2080 91.8159
R2311 GNDA.n2080 GNDA.n213 91.8159
R2312 GNDA.n2074 GNDA.n2073 91.8159
R2313 GNDA.n2073 GNDA.n2072 91.8159
R2314 GNDA.n2072 GNDA.n217 91.8159
R2315 GNDA.n220 GNDA.n217 91.8159
R2316 GNDA.n220 GNDA.n201 91.8159
R2317 GNDA.n2090 GNDA.n2089 91.8159
R2318 GNDA.n2090 GNDA.n196 91.8159
R2319 GNDA.n2097 GNDA.n196 91.8159
R2320 GNDA.n2098 GNDA.n2097 91.8159
R2321 GNDA.n2099 GNDA.n2098 91.8159
R2322 GNDA.n2104 GNDA.n2102 91.8159
R2323 GNDA.n2104 GNDA.n2103 91.8159
R2324 GNDA.n2103 GNDA.n191 91.8159
R2325 GNDA.n2111 GNDA.n191 91.8159
R2326 GNDA.n2112 GNDA.n2111 91.8159
R2327 GNDA.n1743 GNDA.n1734 91.5877
R2328 GNDA.n2451 GNDA.n2450 89.9494
R2329 GNDA.n2367 GNDA.n2333 86.4005
R2330 GNDA.n2255 GNDA.n47 86.4005
R2331 GNDA.n2235 GNDA.n58 85.2842
R2332 GNDA.n2166 GNDA.n2165 85.2842
R2333 GNDA.n337 GNDA.n336 84.306
R2334 GNDA.n1694 GNDA.n92 83.2184
R2335 GNDA.t263 GNDA.t316 82.1737
R2336 GNDA.t66 GNDA.t93 82.1737
R2337 GNDA.t58 GNDA.t43 82.1737
R2338 GNDA.t285 GNDA.t154 82.1737
R2339 GNDA.t253 GNDA.t151 82.1737
R2340 GNDA.t348 GNDA.t272 82.1737
R2341 GNDA.t274 GNDA.t290 82.1737
R2342 GNDA.t347 GNDA.t273 82.1737
R2343 GNDA.n1301 GNDA.n1173 81.7969
R2344 GNDA.n689 GNDA.n563 81.7969
R2345 GNDA.n766 GNDA.n559 81.7969
R2346 GNDA.n2175 GNDA.n2174 81.482
R2347 GNDA.n2184 GNDA.n2183 81.482
R2348 GNDA.t271 GNDA.n2319 78.6626
R2349 GNDA.t254 GNDA.n2356 78.6626
R2350 GNDA.t262 GNDA.t145 78.4385
R2351 GNDA.t259 GNDA.t194 78.4385
R2352 GNDA.n1325 GNDA.n1144 77.7476
R2353 GNDA.n1357 GNDA.n1130 77.7476
R2354 GNDA.n758 GNDA.n691 77.7476
R2355 GNDA.n1363 GNDA.n1362 76.3222
R2356 GNDA.n1366 GNDA.n1365 76.3222
R2357 GNDA.n1371 GNDA.n1370 76.3222
R2358 GNDA.n1374 GNDA.n1373 76.3222
R2359 GNDA.n1379 GNDA.n1378 76.3222
R2360 GNDA.n1382 GNDA.n1381 76.3222
R2361 GNDA.n565 GNDA.n564 76.3222
R2362 GNDA.n686 GNDA.n685 76.3222
R2363 GNDA.n577 GNDA.n576 76.3222
R2364 GNDA.n675 GNDA.n674 76.3222
R2365 GNDA.n586 GNDA.n585 76.3222
R2366 GNDA.n664 GNDA.n663 76.3222
R2367 GNDA.n588 GNDA.n587 76.3222
R2368 GNDA.n1118 GNDA.n391 76.3222
R2369 GNDA.n1114 GNDA.n392 76.3222
R2370 GNDA.n1110 GNDA.n393 76.3222
R2371 GNDA.n1106 GNDA.n394 76.3222
R2372 GNDA.n411 GNDA.n395 76.3222
R2373 GNDA.n1692 GNDA.n390 76.3222
R2374 GNDA.n1844 GNDA.n1843 76.3222
R2375 GNDA.n1941 GNDA.n1940 76.3222
R2376 GNDA.n298 GNDA.n297 76.3222
R2377 GNDA.n1930 GNDA.n1929 76.3222
R2378 GNDA.n307 GNDA.n306 76.3222
R2379 GNDA.n1919 GNDA.n1918 76.3222
R2380 GNDA.n1845 GNDA.n312 76.3222
R2381 GNDA.n1300 GNDA.n1171 76.3222
R2382 GNDA.n1298 GNDA.n1175 76.3222
R2383 GNDA.n1293 GNDA.n1178 76.3222
R2384 GNDA.n1285 GNDA.n1284 76.3222
R2385 GNDA.n1191 GNDA.n1184 76.3222
R2386 GNDA.n1274 GNDA.n1273 76.3222
R2387 GNDA.n1198 GNDA.n1193 76.3222
R2388 GNDA.n937 GNDA.n398 76.3222
R2389 GNDA.n943 GNDA.n399 76.3222
R2390 GNDA.n949 GNDA.n400 76.3222
R2391 GNDA.n955 GNDA.n401 76.3222
R2392 GNDA.n958 GNDA.n402 76.3222
R2393 GNDA.n1196 GNDA.n396 76.3222
R2394 GNDA.n1387 GNDA.n1386 76.3222
R2395 GNDA.n1392 GNDA.n1391 76.3222
R2396 GNDA.n1395 GNDA.n1394 76.3222
R2397 GNDA.n1400 GNDA.n1399 76.3222
R2398 GNDA.n1403 GNDA.n1402 76.3222
R2399 GNDA.n1408 GNDA.n1407 76.3222
R2400 GNDA.n1095 GNDA.n419 76.3222
R2401 GNDA.n1097 GNDA.n420 76.3222
R2402 GNDA.n1099 GNDA.n421 76.3222
R2403 GNDA.n1101 GNDA.n422 76.3222
R2404 GNDA.n1103 GNDA.n423 76.3222
R2405 GNDA.n1688 GNDA.n1687 76.3222
R2406 GNDA.n1533 GNDA.n1532 76.3222
R2407 GNDA.n871 GNDA.n870 76.3222
R2408 GNDA.n1522 GNDA.n1521 76.3222
R2409 GNDA.n880 GNDA.n879 76.3222
R2410 GNDA.n1511 GNDA.n1510 76.3222
R2411 GNDA.n1437 GNDA.n885 76.3222
R2412 GNDA.n1410 GNDA.n894 76.3222
R2413 GNDA.n1419 GNDA.n1418 76.3222
R2414 GNDA.n1420 GNDA.n890 76.3222
R2415 GNDA.n1429 GNDA.n1428 76.3222
R2416 GNDA.n1433 GNDA.n886 76.3222
R2417 GNDA.n1436 GNDA.n1435 76.3222
R2418 GNDA.n2023 GNDA.n2022 76.3222
R2419 GNDA.n2052 GNDA.n2051 76.3222
R2420 GNDA.n2044 GNDA.n2027 76.3222
R2421 GNDA.n2042 GNDA.n2041 76.3222
R2422 GNDA.n2029 GNDA.n222 76.3222
R2423 GNDA.n2065 GNDA.n2064 76.3222
R2424 GNDA.n2067 GNDA.n2066 76.3222
R2425 GNDA.n923 GNDA.n922 76.3222
R2426 GNDA.n920 GNDA.n919 76.3222
R2427 GNDA.n915 GNDA.n902 76.3222
R2428 GNDA.n913 GNDA.n912 76.3222
R2429 GNDA.n908 GNDA.n905 76.3222
R2430 GNDA.n906 GNDA.n208 76.3222
R2431 GNDA.n924 GNDA.n923 76.3222
R2432 GNDA.n921 GNDA.n920 76.3222
R2433 GNDA.n902 GNDA.n900 76.3222
R2434 GNDA.n914 GNDA.n913 76.3222
R2435 GNDA.n905 GNDA.n903 76.3222
R2436 GNDA.n907 GNDA.n906 76.3222
R2437 GNDA.n1085 GNDA.n1084 76.3222
R2438 GNDA.n971 GNDA.n970 76.3222
R2439 GNDA.n1074 GNDA.n1073 76.3222
R2440 GNDA.n980 GNDA.n979 76.3222
R2441 GNDA.n1063 GNDA.n1062 76.3222
R2442 GNDA.n989 GNDA.n985 76.3222
R2443 GNDA.n1961 GNDA.n272 76.3222
R2444 GNDA.n1959 GNDA.n1958 76.3222
R2445 GNDA.n1954 GNDA.n280 76.3222
R2446 GNDA.n1952 GNDA.n1951 76.3222
R2447 GNDA.n285 GNDA.n284 76.3222
R2448 GNDA.n988 GNDA.n987 76.3222
R2449 GNDA.n1539 GNDA.n1538 76.3222
R2450 GNDA.n1544 GNDA.n1543 76.3222
R2451 GNDA.n1547 GNDA.n1546 76.3222
R2452 GNDA.n1552 GNDA.n1551 76.3222
R2453 GNDA.n1555 GNDA.n1554 76.3222
R2454 GNDA.n1560 GNDA.n1559 76.3222
R2455 GNDA.n1563 GNDA.n467 76.3222
R2456 GNDA.n1572 GNDA.n1571 76.3222
R2457 GNDA.n1573 GNDA.n463 76.3222
R2458 GNDA.n1582 GNDA.n1581 76.3222
R2459 GNDA.n459 GNDA.n458 76.3222
R2460 GNDA.n1680 GNDA.n94 76.3222
R2461 GNDA.n444 GNDA.n95 76.3222
R2462 GNDA.n1670 GNDA.n96 76.3222
R2463 GNDA.n452 GNDA.n97 76.3222
R2464 GNDA.n1660 GNDA.n98 76.3222
R2465 GNDA.n511 GNDA.n431 76.3222
R2466 GNDA.n513 GNDA.n432 76.3222
R2467 GNDA.n515 GNDA.n433 76.3222
R2468 GNDA.n517 GNDA.n434 76.3222
R2469 GNDA.n1685 GNDA.n436 76.3222
R2470 GNDA.n500 GNDA.n499 76.3222
R2471 GNDA.n497 GNDA.n473 76.3222
R2472 GNDA.n493 GNDA.n492 76.3222
R2473 GNDA.n486 GNDA.n475 76.3222
R2474 GNDA.n485 GNDA.n484 76.3222
R2475 GNDA.n478 GNDA.n477 76.3222
R2476 GNDA.n2113 GNDA.n190 76.3222
R2477 GNDA.n106 GNDA.n100 76.3222
R2478 GNDA.n2144 GNDA.n101 76.3222
R2479 GNDA.n2136 GNDA.n102 76.3222
R2480 GNDA.n2131 GNDA.n103 76.3222
R2481 GNDA.n2123 GNDA.n104 76.3222
R2482 GNDA.n2118 GNDA.n105 76.3222
R2483 GNDA.n1567 GNDA.n258 76.3222
R2484 GNDA.n465 GNDA.n259 76.3222
R2485 GNDA.n1577 GNDA.n260 76.3222
R2486 GNDA.n461 GNDA.n261 76.3222
R2487 GNDA.n732 GNDA.n558 76.3222
R2488 GNDA.n852 GNDA.n408 76.3222
R2489 GNDA.n848 GNDA.n407 76.3222
R2490 GNDA.n844 GNDA.n406 76.3222
R2491 GNDA.n840 GNDA.n405 76.3222
R2492 GNDA.n835 GNDA.n403 76.3222
R2493 GNDA.n720 GNDA.n695 76.3222
R2494 GNDA.n718 GNDA.n717 76.3222
R2495 GNDA.n713 GNDA.n698 76.3222
R2496 GNDA.n711 GNDA.n710 76.3222
R2497 GNDA.n706 GNDA.n701 76.3222
R2498 GNDA.n704 GNDA.n703 76.3222
R2499 GNDA.n695 GNDA.n692 76.3222
R2500 GNDA.n719 GNDA.n718 76.3222
R2501 GNDA.n698 GNDA.n696 76.3222
R2502 GNDA.n712 GNDA.n711 76.3222
R2503 GNDA.n701 GNDA.n699 76.3222
R2504 GNDA.n705 GNDA.n704 76.3222
R2505 GNDA.n2114 GNDA.n105 76.3222
R2506 GNDA.n2119 GNDA.n104 76.3222
R2507 GNDA.n2122 GNDA.n103 76.3222
R2508 GNDA.n2132 GNDA.n102 76.3222
R2509 GNDA.n2135 GNDA.n101 76.3222
R2510 GNDA.n2145 GNDA.n100 76.3222
R2511 GNDA.n455 GNDA.n98 76.3222
R2512 GNDA.n1661 GNDA.n97 76.3222
R2513 GNDA.n451 GNDA.n96 76.3222
R2514 GNDA.n1671 GNDA.n95 76.3222
R2515 GNDA.n443 GNDA.n94 76.3222
R2516 GNDA.n1964 GNDA.n1963 76.3222
R2517 GNDA.n275 GNDA.n267 76.3222
R2518 GNDA.n277 GNDA.n266 76.3222
R2519 GNDA.n282 GNDA.n265 76.3222
R2520 GNDA.n1947 GNDA.n264 76.3222
R2521 GNDA.n1946 GNDA.n251 76.3222
R2522 GNDA.n283 GNDA.n264 76.3222
R2523 GNDA.n278 GNDA.n265 76.3222
R2524 GNDA.n276 GNDA.n266 76.3222
R2525 GNDA.n269 GNDA.n267 76.3222
R2526 GNDA.n1964 GNDA.n268 76.3222
R2527 GNDA.n262 GNDA.n107 76.3222
R2528 GNDA.n462 GNDA.n263 76.3222
R2529 GNDA.n1578 GNDA.n261 76.3222
R2530 GNDA.n466 GNDA.n260 76.3222
R2531 GNDA.n1568 GNDA.n259 76.3222
R2532 GNDA.n469 GNDA.n258 76.3222
R2533 GNDA.n284 GNDA.n281 76.3222
R2534 GNDA.n1953 GNDA.n1952 76.3222
R2535 GNDA.n280 GNDA.n274 76.3222
R2536 GNDA.n1960 GNDA.n1959 76.3222
R2537 GNDA.n329 GNDA.n272 76.3222
R2538 GNDA.n1584 GNDA.n1583 76.3222
R2539 GNDA.n1581 GNDA.n1580 76.3222
R2540 GNDA.n1574 GNDA.n1573 76.3222
R2541 GNDA.n1571 GNDA.n1570 76.3222
R2542 GNDA.n1564 GNDA.n1563 76.3222
R2543 GNDA.n896 GNDA.n252 76.3222
R2544 GNDA.n1415 GNDA.n253 76.3222
R2545 GNDA.n893 GNDA.n254 76.3222
R2546 GNDA.n1425 GNDA.n255 76.3222
R2547 GNDA.n889 GNDA.n256 76.3222
R2548 GNDA.n1967 GNDA.n1966 76.3222
R2549 GNDA.n256 GNDA.n250 76.3222
R2550 GNDA.n888 GNDA.n255 76.3222
R2551 GNDA.n1424 GNDA.n254 76.3222
R2552 GNDA.n892 GNDA.n253 76.3222
R2553 GNDA.n1414 GNDA.n252 76.3222
R2554 GNDA.n1430 GNDA.n886 76.3222
R2555 GNDA.n1428 GNDA.n1427 76.3222
R2556 GNDA.n1421 GNDA.n1420 76.3222
R2557 GNDA.n1418 GNDA.n1417 76.3222
R2558 GNDA.n1411 GNDA.n1410 76.3222
R2559 GNDA.n1386 GNDA.n933 76.3222
R2560 GNDA.n1393 GNDA.n1392 76.3222
R2561 GNDA.n1394 GNDA.n931 76.3222
R2562 GNDA.n1401 GNDA.n1400 76.3222
R2563 GNDA.n1402 GNDA.n929 76.3222
R2564 GNDA.n1409 GNDA.n1408 76.3222
R2565 GNDA.n1538 GNDA.n509 76.3222
R2566 GNDA.n1545 GNDA.n1544 76.3222
R2567 GNDA.n1546 GNDA.n507 76.3222
R2568 GNDA.n1553 GNDA.n1552 76.3222
R2569 GNDA.n1554 GNDA.n505 76.3222
R2570 GNDA.n1561 GNDA.n1560 76.3222
R2571 GNDA.n518 GNDA.n435 76.3222
R2572 GNDA.n516 GNDA.n434 76.3222
R2573 GNDA.n514 GNDA.n433 76.3222
R2574 GNDA.n512 GNDA.n432 76.3222
R2575 GNDA.n510 GNDA.n431 76.3222
R2576 GNDA.n839 GNDA.n404 76.3222
R2577 GNDA.n843 GNDA.n405 76.3222
R2578 GNDA.n847 GNDA.n406 76.3222
R2579 GNDA.n851 GNDA.n407 76.3222
R2580 GNDA.n854 GNDA.n408 76.3222
R2581 GNDA.n425 GNDA.n389 76.3222
R2582 GNDA.n936 GNDA.n426 76.3222
R2583 GNDA.n942 GNDA.n427 76.3222
R2584 GNDA.n948 GNDA.n428 76.3222
R2585 GNDA.n954 GNDA.n429 76.3222
R2586 GNDA.n1090 GNDA.n424 76.3222
R2587 GNDA.n1089 GNDA.n429 76.3222
R2588 GNDA.n953 GNDA.n428 76.3222
R2589 GNDA.n947 GNDA.n427 76.3222
R2590 GNDA.n941 GNDA.n426 76.3222
R2591 GNDA.n935 GNDA.n425 76.3222
R2592 GNDA.n956 GNDA.n402 76.3222
R2593 GNDA.n950 GNDA.n401 76.3222
R2594 GNDA.n944 GNDA.n400 76.3222
R2595 GNDA.n938 GNDA.n399 76.3222
R2596 GNDA.n398 GNDA.n397 76.3222
R2597 GNDA.n287 GNDA.n251 76.3222
R2598 GNDA.n312 GNDA.n308 76.3222
R2599 GNDA.n1920 GNDA.n1919 76.3222
R2600 GNDA.n306 GNDA.n299 76.3222
R2601 GNDA.n1931 GNDA.n1930 76.3222
R2602 GNDA.n297 GNDA.n289 76.3222
R2603 GNDA.n1942 GNDA.n1941 76.3222
R2604 GNDA.n960 GNDA.n424 76.3222
R2605 GNDA.n985 GNDA.n981 76.3222
R2606 GNDA.n1064 GNDA.n1063 76.3222
R2607 GNDA.n979 GNDA.n972 76.3222
R2608 GNDA.n1075 GNDA.n1074 76.3222
R2609 GNDA.n970 GNDA.n963 76.3222
R2610 GNDA.n1086 GNDA.n1085 76.3222
R2611 GNDA.n987 GNDA.n986 76.3222
R2612 GNDA.n1199 GNDA.n1198 76.3222
R2613 GNDA.n1273 GNDA.n1272 76.3222
R2614 GNDA.n1192 GNDA.n1191 76.3222
R2615 GNDA.n1284 GNDA.n1283 76.3222
R2616 GNDA.n1183 GNDA.n1178 76.3222
R2617 GNDA.n1294 GNDA.n1175 76.3222
R2618 GNDA.n1196 GNDA.n410 76.3222
R2619 GNDA.n423 GNDA.n417 76.3222
R2620 GNDA.n1102 GNDA.n422 76.3222
R2621 GNDA.n1100 GNDA.n421 76.3222
R2622 GNDA.n1098 GNDA.n420 76.3222
R2623 GNDA.n1096 GNDA.n419 76.3222
R2624 GNDA.n1105 GNDA.n395 76.3222
R2625 GNDA.n1109 GNDA.n394 76.3222
R2626 GNDA.n1113 GNDA.n393 76.3222
R2627 GNDA.n1117 GNDA.n392 76.3222
R2628 GNDA.n1121 GNDA.n391 76.3222
R2629 GNDA.n1364 GNDA.n1363 76.3222
R2630 GNDA.n1365 GNDA.n1125 76.3222
R2631 GNDA.n1372 GNDA.n1371 76.3222
R2632 GNDA.n1373 GNDA.n1123 76.3222
R2633 GNDA.n1380 GNDA.n1379 76.3222
R2634 GNDA.n1383 GNDA.n1382 76.3222
R2635 GNDA.n1966 GNDA.n249 76.3222
R2636 GNDA.n1687 GNDA.n415 76.3222
R2637 GNDA.n885 GNDA.n881 76.3222
R2638 GNDA.n1512 GNDA.n1511 76.3222
R2639 GNDA.n879 GNDA.n872 76.3222
R2640 GNDA.n1523 GNDA.n1522 76.3222
R2641 GNDA.n870 GNDA.n862 76.3222
R2642 GNDA.n1534 GNDA.n1533 76.3222
R2643 GNDA.n1435 GNDA.n1434 76.3222
R2644 GNDA.n589 GNDA.n588 76.3222
R2645 GNDA.n665 GNDA.n664 76.3222
R2646 GNDA.n585 GNDA.n578 76.3222
R2647 GNDA.n676 GNDA.n675 76.3222
R2648 GNDA.n576 GNDA.n568 76.3222
R2649 GNDA.n687 GNDA.n686 76.3222
R2650 GNDA.n1693 GNDA.n1692 76.3222
R2651 GNDA.n2064 GNDA.n2063 76.3222
R2652 GNDA.n2030 GNDA.n2029 76.3222
R2653 GNDA.n2043 GNDA.n2042 76.3222
R2654 GNDA.n2027 GNDA.n2024 76.3222
R2655 GNDA.n2053 GNDA.n2052 76.3222
R2656 GNDA.n2022 GNDA.n2021 76.3222
R2657 GNDA.n499 GNDA.n498 76.3222
R2658 GNDA.n494 GNDA.n473 76.3222
R2659 GNDA.n492 GNDA.n491 76.3222
R2660 GNDA.n487 GNDA.n486 76.3222
R2661 GNDA.n484 GNDA.n483 76.3222
R2662 GNDA.n479 GNDA.n478 76.3222
R2663 GNDA.n1843 GNDA.n1842 76.3222
R2664 GNDA.n2067 GNDA.n221 76.3222
R2665 GNDA.n2110 GNDA.n190 76.3222
R2666 GNDA.n1303 GNDA.n1171 76.3222
R2667 GNDA.n564 GNDA.n354 76.3222
R2668 GNDA.n733 GNDA.n732 76.3222
R2669 GNDA.n2351 GNDA.n2340 76.1251
R2670 GNDA.n809 GNDA.n808 76.062
R2671 GNDA.n808 GNDA.n807 76.062
R2672 GNDA.n1640 GNDA.n1639 76.062
R2673 GNDA.n1639 GNDA.n1638 76.062
R2674 GNDA.n169 GNDA.n126 76.062
R2675 GNDA.n170 GNDA.n169 76.062
R2676 GNDA.n1252 GNDA.n1251 76.062
R2677 GNDA.n1251 GNDA.n1250 76.062
R2678 GNDA.n1042 GNDA.n1041 76.062
R2679 GNDA.n1041 GNDA.n1040 76.062
R2680 GNDA.n1898 GNDA.n1897 76.062
R2681 GNDA.n1897 GNDA.n1896 76.062
R2682 GNDA.n643 GNDA.n642 76.062
R2683 GNDA.n642 GNDA.n641 76.062
R2684 GNDA.n1490 GNDA.n1489 76.062
R2685 GNDA.n1489 GNDA.n1488 76.062
R2686 GNDA.n1982 GNDA.n227 76.062
R2687 GNDA.n1985 GNDA.n227 76.062
R2688 GNDA.t244 GNDA.t270 75.2142
R2689 GNDA.t323 GNDA.t96 75.2142
R2690 GNDA.n1319 GNDA.n1318 72.8884
R2691 GNDA.n1318 GNDA.n1317 72.8884
R2692 GNDA.n1317 GNDA.n1164 72.8884
R2693 GNDA.n1311 GNDA.n1164 72.8884
R2694 GNDA.n1310 GNDA.n1309 72.8884
R2695 GNDA.n1309 GNDA.n1168 72.8884
R2696 GNDA.n1168 GNDA.n1138 72.8884
R2697 GNDA.n1302 GNDA.n1301 72.8884
R2698 GNDA.n1357 GNDA.n1356 72.8884
R2699 GNDA.n1356 GNDA.n1355 72.8884
R2700 GNDA.n1349 GNDA.n1347 72.8884
R2701 GNDA.n1349 GNDA.n1348 72.8884
R2702 GNDA.n1751 GNDA.n355 72.8884
R2703 GNDA.n563 GNDA.n356 72.8884
R2704 GNDA.n752 GNDA.n691 72.8884
R2705 GNDA.n752 GNDA.n751 72.8884
R2706 GNDA.n751 GNDA.n750 72.8884
R2707 GNDA.n750 GNDA.n725 72.8884
R2708 GNDA.n744 GNDA.n725 72.8884
R2709 GNDA.n743 GNDA.n742 72.8884
R2710 GNDA.n736 GNDA.n734 72.8884
R2711 GNDA.n736 GNDA.n735 72.8884
R2712 GNDA.n735 GNDA.n559 72.8884
R2713 GNDA.t187 GNDA.t320 72.0803
R2714 GNDA.t275 GNDA.t163 72.0803
R2715 GNDA.t99 GNDA.t262 70.9682
R2716 GNDA.t129 GNDA.t285 70.9682
R2717 GNDA.t200 GNDA.t253 70.9682
R2718 GNDA.t97 GNDA.t259 70.9682
R2719 GNDA.n1172 GNDA.n1130 70.4588
R2720 GNDA.n1758 GNDA.n349 70.4588
R2721 GNDA.n2492 GNDA.n20 70.4005
R2722 GNDA.n2492 GNDA.n22 70.4005
R2723 GNDA.n1173 GNDA.n1172 69.6489
R2724 GNDA.n690 GNDA.n689 69.6489
R2725 GNDA.t351 GNDA.t184 68.9464
R2726 GNDA.t38 GNDA.t351 68.9464
R2727 GNDA.t328 GNDA.t38 68.9464
R2728 GNDA.t336 GNDA.t313 68.9464
R2729 GNDA.t14 GNDA.t336 68.9464
R2730 GNDA.t123 GNDA.t14 68.9464
R2731 GNDA.n776 GNDA.t134 65.8183
R2732 GNDA.n778 GNDA.t134 65.8183
R2733 GNDA.n784 GNDA.t134 65.8183
R2734 GNDA.n786 GNDA.t134 65.8183
R2735 GNDA.n792 GNDA.t134 65.8183
R2736 GNDA.n794 GNDA.t134 65.8183
R2737 GNDA.n800 GNDA.t134 65.8183
R2738 GNDA.n802 GNDA.t134 65.8183
R2739 GNDA.n824 GNDA.t134 65.8183
R2740 GNDA.n818 GNDA.t134 65.8183
R2741 GNDA.n816 GNDA.t134 65.8183
R2742 GNDA.n810 GNDA.t134 65.8183
R2743 GNDA.n1607 GNDA.t136 65.8183
R2744 GNDA.n1609 GNDA.t136 65.8183
R2745 GNDA.n1615 GNDA.t136 65.8183
R2746 GNDA.n1617 GNDA.t136 65.8183
R2747 GNDA.n1623 GNDA.t136 65.8183
R2748 GNDA.n1625 GNDA.t136 65.8183
R2749 GNDA.n1631 GNDA.t136 65.8183
R2750 GNDA.n1633 GNDA.t136 65.8183
R2751 GNDA.n1655 GNDA.t136 65.8183
R2752 GNDA.n1649 GNDA.t136 65.8183
R2753 GNDA.n1647 GNDA.t136 65.8183
R2754 GNDA.n1641 GNDA.t136 65.8183
R2755 GNDA.n137 GNDA.t170 65.8183
R2756 GNDA.n143 GNDA.t170 65.8183
R2757 GNDA.n145 GNDA.t170 65.8183
R2758 GNDA.n151 GNDA.t170 65.8183
R2759 GNDA.n153 GNDA.t170 65.8183
R2760 GNDA.n159 GNDA.t170 65.8183
R2761 GNDA.n161 GNDA.t170 65.8183
R2762 GNDA.n167 GNDA.t170 65.8183
R2763 GNDA.n186 GNDA.t170 65.8183
R2764 GNDA.n183 GNDA.t170 65.8183
R2765 GNDA.n177 GNDA.t170 65.8183
R2766 GNDA.n175 GNDA.t170 65.8183
R2767 GNDA.n121 GNDA.t170 65.8183
R2768 GNDA.n2127 GNDA.t170 65.8183
R2769 GNDA.n116 GNDA.t170 65.8183
R2770 GNDA.n2140 GNDA.t170 65.8183
R2771 GNDA.n457 GNDA.t136 65.8183
R2772 GNDA.n1665 GNDA.t136 65.8183
R2773 GNDA.n448 GNDA.t136 65.8183
R2774 GNDA.n1675 GNDA.t136 65.8183
R2775 GNDA.n541 GNDA.t134 65.8183
R2776 GNDA.n525 GNDA.t134 65.8183
R2777 GNDA.n528 GNDA.t134 65.8183
R2778 GNDA.n1729 GNDA.t134 65.8183
R2779 GNDA.n1219 GNDA.t180 65.8183
R2780 GNDA.n1221 GNDA.t180 65.8183
R2781 GNDA.n1227 GNDA.t180 65.8183
R2782 GNDA.n1229 GNDA.t180 65.8183
R2783 GNDA.n1235 GNDA.t180 65.8183
R2784 GNDA.n1237 GNDA.t180 65.8183
R2785 GNDA.n1243 GNDA.t180 65.8183
R2786 GNDA.n1245 GNDA.t180 65.8183
R2787 GNDA.n1267 GNDA.t180 65.8183
R2788 GNDA.n1261 GNDA.t180 65.8183
R2789 GNDA.n1259 GNDA.t180 65.8183
R2790 GNDA.n1253 GNDA.t180 65.8183
R2791 GNDA.n1009 GNDA.t182 65.8183
R2792 GNDA.n1011 GNDA.t182 65.8183
R2793 GNDA.n1017 GNDA.t182 65.8183
R2794 GNDA.n1019 GNDA.t182 65.8183
R2795 GNDA.n1025 GNDA.t182 65.8183
R2796 GNDA.n1027 GNDA.t182 65.8183
R2797 GNDA.n1033 GNDA.t182 65.8183
R2798 GNDA.n1035 GNDA.t182 65.8183
R2799 GNDA.n1057 GNDA.t182 65.8183
R2800 GNDA.n1051 GNDA.t182 65.8183
R2801 GNDA.n1049 GNDA.t182 65.8183
R2802 GNDA.n1043 GNDA.t182 65.8183
R2803 GNDA.n1865 GNDA.t192 65.8183
R2804 GNDA.n1867 GNDA.t192 65.8183
R2805 GNDA.n1873 GNDA.t192 65.8183
R2806 GNDA.n1875 GNDA.t192 65.8183
R2807 GNDA.n1881 GNDA.t192 65.8183
R2808 GNDA.n1883 GNDA.t192 65.8183
R2809 GNDA.n1889 GNDA.t192 65.8183
R2810 GNDA.n1891 GNDA.t192 65.8183
R2811 GNDA.n1913 GNDA.t192 65.8183
R2812 GNDA.n1907 GNDA.t192 65.8183
R2813 GNDA.n1905 GNDA.t192 65.8183
R2814 GNDA.n1899 GNDA.t192 65.8183
R2815 GNDA.n310 GNDA.t192 65.8183
R2816 GNDA.n1924 GNDA.t192 65.8183
R2817 GNDA.n301 GNDA.t192 65.8183
R2818 GNDA.n1935 GNDA.t192 65.8183
R2819 GNDA.n983 GNDA.t182 65.8183
R2820 GNDA.n1068 GNDA.t182 65.8183
R2821 GNDA.n974 GNDA.t182 65.8183
R2822 GNDA.n1079 GNDA.t182 65.8183
R2823 GNDA.n1195 GNDA.t180 65.8183
R2824 GNDA.n1278 GNDA.t180 65.8183
R2825 GNDA.n1186 GNDA.t180 65.8183
R2826 GNDA.n1289 GNDA.t180 65.8183
R2827 GNDA.n610 GNDA.t175 65.8183
R2828 GNDA.n612 GNDA.t175 65.8183
R2829 GNDA.n618 GNDA.t175 65.8183
R2830 GNDA.n620 GNDA.t175 65.8183
R2831 GNDA.n626 GNDA.t175 65.8183
R2832 GNDA.n628 GNDA.t175 65.8183
R2833 GNDA.n634 GNDA.t175 65.8183
R2834 GNDA.n636 GNDA.t175 65.8183
R2835 GNDA.n658 GNDA.t175 65.8183
R2836 GNDA.n652 GNDA.t175 65.8183
R2837 GNDA.n650 GNDA.t175 65.8183
R2838 GNDA.n644 GNDA.t175 65.8183
R2839 GNDA.n1457 GNDA.t179 65.8183
R2840 GNDA.n1459 GNDA.t179 65.8183
R2841 GNDA.n1465 GNDA.t179 65.8183
R2842 GNDA.n1467 GNDA.t179 65.8183
R2843 GNDA.n1473 GNDA.t179 65.8183
R2844 GNDA.n1475 GNDA.t179 65.8183
R2845 GNDA.n1481 GNDA.t179 65.8183
R2846 GNDA.n1483 GNDA.t179 65.8183
R2847 GNDA.n1505 GNDA.t179 65.8183
R2848 GNDA.n1499 GNDA.t179 65.8183
R2849 GNDA.n1497 GNDA.t179 65.8183
R2850 GNDA.n1491 GNDA.t179 65.8183
R2851 GNDA.t181 GNDA.n238 65.8183
R2852 GNDA.t181 GNDA.n236 65.8183
R2853 GNDA.t181 GNDA.n234 65.8183
R2854 GNDA.t181 GNDA.n228 65.8183
R2855 GNDA.t181 GNDA.n229 65.8183
R2856 GNDA.t181 GNDA.n230 65.8183
R2857 GNDA.t181 GNDA.n231 65.8183
R2858 GNDA.t181 GNDA.n232 65.8183
R2859 GNDA.n2058 GNDA.t181 65.8183
R2860 GNDA.t181 GNDA.n237 65.8183
R2861 GNDA.t181 GNDA.n235 65.8183
R2862 GNDA.t181 GNDA.n233 65.8183
R2863 GNDA.t181 GNDA.n239 65.8183
R2864 GNDA.t181 GNDA.n240 65.8183
R2865 GNDA.t181 GNDA.n241 65.8183
R2866 GNDA.t181 GNDA.n242 65.8183
R2867 GNDA.n883 GNDA.t179 65.8183
R2868 GNDA.n1516 GNDA.t179 65.8183
R2869 GNDA.n874 GNDA.t179 65.8183
R2870 GNDA.n1527 GNDA.t179 65.8183
R2871 GNDA.n591 GNDA.t175 65.8183
R2872 GNDA.n669 GNDA.t175 65.8183
R2873 GNDA.n580 GNDA.t175 65.8183
R2874 GNDA.n680 GNDA.t175 65.8183
R2875 GNDA.n2162 GNDA.t328 65.8125
R2876 GNDA.t313 GNDA.n2182 65.8125
R2877 GNDA.n135 GNDA.t170 64.1729
R2878 GNDA.t136 GNDA.n440 64.1729
R2879 GNDA.n555 GNDA.t134 64.1729
R2880 GNDA.t192 GNDA.n292 64.1729
R2881 GNDA.t182 GNDA.n965 64.1729
R2882 GNDA.n1215 GNDA.t180 64.1729
R2883 GNDA.t181 GNDA.n2057 64.1729
R2884 GNDA.t179 GNDA.n865 64.1729
R2885 GNDA.t175 GNDA.n571 64.1729
R2886 GNDA.n2157 GNDA.t226 62.6786
R2887 GNDA.n2208 GNDA.t319 62.6786
R2888 GNDA.n1355 GNDA.n1342 62.3602
R2889 GNDA.t137 GNDA.n0 32.9056
R2890 GNDA.n2446 GNDA.n2445 60.8005
R2891 GNDA.t116 GNDA.t247 59.5447
R2892 GNDA.t36 GNDA.t5 59.5447
R2893 GNDA.n555 GNDA.n367 56.6572
R2894 GNDA.n556 GNDA.n555 56.6572
R2895 GNDA.n1677 GNDA.n440 56.6572
R2896 GNDA.n1603 GNDA.n440 56.6572
R2897 GNDA.n135 GNDA.n112 56.6572
R2898 GNDA.n136 GNDA.n135 56.6572
R2899 GNDA.n1215 GNDA.n1180 56.6572
R2900 GNDA.n1216 GNDA.n1215 56.6572
R2901 GNDA.n1081 GNDA.n965 56.6572
R2902 GNDA.n1005 GNDA.n965 56.6572
R2903 GNDA.n1937 GNDA.n292 56.6572
R2904 GNDA.n1861 GNDA.n292 56.6572
R2905 GNDA.n682 GNDA.n571 56.6572
R2906 GNDA.n606 GNDA.n571 56.6572
R2907 GNDA.n1529 GNDA.n865 56.6572
R2908 GNDA.n1453 GNDA.n865 56.6572
R2909 GNDA.n2057 GNDA.n2056 56.6572
R2910 GNDA.n2057 GNDA.n243 56.6572
R2911 GNDA.n1684 GNDA.n93 56.3995
R2912 GNDA.n1681 GNDA.n93 56.3995
R2913 GNDA.t343 GNDA.t263 56.0277
R2914 GNDA.t245 GNDA.t58 56.0277
R2915 GNDA.t85 GNDA.t348 56.0277
R2916 GNDA.t308 GNDA.t347 56.0277
R2917 GNDA.n808 GNDA.t134 54.4705
R2918 GNDA.n1639 GNDA.t136 54.4705
R2919 GNDA.n169 GNDA.t170 54.4705
R2920 GNDA.n1251 GNDA.t180 54.4705
R2921 GNDA.n1041 GNDA.t182 54.4705
R2922 GNDA.n1897 GNDA.t192 54.4705
R2923 GNDA.n642 GNDA.t175 54.4705
R2924 GNDA.n1489 GNDA.t179 54.4705
R2925 GNDA.t181 GNDA.n227 54.4705
R2926 GNDA.n2447 GNDA.n2446 54.4005
R2927 GNDA.n1751 GNDA.n1750 54.2615
R2928 GNDA.n1729 GNDA.n1728 53.3664
R2929 GNDA.n530 GNDA.n528 53.3664
R2930 GNDA.n539 GNDA.n525 53.3664
R2931 GNDA.n826 GNDA.n541 53.3664
R2932 GNDA.n811 GNDA.n810 53.3664
R2933 GNDA.n816 GNDA.n815 53.3664
R2934 GNDA.n819 GNDA.n818 53.3664
R2935 GNDA.n824 GNDA.n823 53.3664
R2936 GNDA.n792 GNDA.n791 53.3664
R2937 GNDA.n795 GNDA.n794 53.3664
R2938 GNDA.n800 GNDA.n799 53.3664
R2939 GNDA.n803 GNDA.n802 53.3664
R2940 GNDA.n786 GNDA.n551 53.3664
R2941 GNDA.n785 GNDA.n784 53.3664
R2942 GNDA.n778 GNDA.n553 53.3664
R2943 GNDA.n777 GNDA.n776 53.3664
R2944 GNDA.n776 GNDA.n775 53.3664
R2945 GNDA.n779 GNDA.n778 53.3664
R2946 GNDA.n784 GNDA.n783 53.3664
R2947 GNDA.n787 GNDA.n786 53.3664
R2948 GNDA.n793 GNDA.n792 53.3664
R2949 GNDA.n794 GNDA.n549 53.3664
R2950 GNDA.n801 GNDA.n800 53.3664
R2951 GNDA.n802 GNDA.n547 53.3664
R2952 GNDA.n825 GNDA.n824 53.3664
R2953 GNDA.n818 GNDA.n543 53.3664
R2954 GNDA.n817 GNDA.n816 53.3664
R2955 GNDA.n810 GNDA.n545 53.3664
R2956 GNDA.n1675 GNDA.n1674 53.3664
R2957 GNDA.n1667 GNDA.n448 53.3664
R2958 GNDA.n1665 GNDA.n1664 53.3664
R2959 GNDA.n1657 GNDA.n457 53.3664
R2960 GNDA.n1642 GNDA.n1641 53.3664
R2961 GNDA.n1647 GNDA.n1646 53.3664
R2962 GNDA.n1650 GNDA.n1649 53.3664
R2963 GNDA.n1655 GNDA.n1654 53.3664
R2964 GNDA.n1623 GNDA.n1622 53.3664
R2965 GNDA.n1626 GNDA.n1625 53.3664
R2966 GNDA.n1631 GNDA.n1630 53.3664
R2967 GNDA.n1634 GNDA.n1633 53.3664
R2968 GNDA.n1617 GNDA.n1599 53.3664
R2969 GNDA.n1616 GNDA.n1615 53.3664
R2970 GNDA.n1609 GNDA.n1601 53.3664
R2971 GNDA.n1608 GNDA.n1607 53.3664
R2972 GNDA.n1607 GNDA.n1606 53.3664
R2973 GNDA.n1610 GNDA.n1609 53.3664
R2974 GNDA.n1615 GNDA.n1614 53.3664
R2975 GNDA.n1618 GNDA.n1617 53.3664
R2976 GNDA.n1624 GNDA.n1623 53.3664
R2977 GNDA.n1625 GNDA.n1597 53.3664
R2978 GNDA.n1632 GNDA.n1631 53.3664
R2979 GNDA.n1633 GNDA.n1595 53.3664
R2980 GNDA.n1656 GNDA.n1655 53.3664
R2981 GNDA.n1649 GNDA.n1591 53.3664
R2982 GNDA.n1648 GNDA.n1647 53.3664
R2983 GNDA.n1641 GNDA.n1593 53.3664
R2984 GNDA.n2140 GNDA.n2139 53.3664
R2985 GNDA.n117 GNDA.n116 53.3664
R2986 GNDA.n2127 GNDA.n2126 53.3664
R2987 GNDA.n122 GNDA.n121 53.3664
R2988 GNDA.n175 GNDA.n174 53.3664
R2989 GNDA.n178 GNDA.n177 53.3664
R2990 GNDA.n183 GNDA.n182 53.3664
R2991 GNDA.n186 GNDA.n185 53.3664
R2992 GNDA.n154 GNDA.n153 53.3664
R2993 GNDA.n159 GNDA.n158 53.3664
R2994 GNDA.n162 GNDA.n161 53.3664
R2995 GNDA.n167 GNDA.n166 53.3664
R2996 GNDA.n152 GNDA.n151 53.3664
R2997 GNDA.n145 GNDA.n132 53.3664
R2998 GNDA.n144 GNDA.n143 53.3664
R2999 GNDA.n137 GNDA.n134 53.3664
R3000 GNDA.n138 GNDA.n137 53.3664
R3001 GNDA.n143 GNDA.n142 53.3664
R3002 GNDA.n146 GNDA.n145 53.3664
R3003 GNDA.n151 GNDA.n150 53.3664
R3004 GNDA.n153 GNDA.n130 53.3664
R3005 GNDA.n160 GNDA.n159 53.3664
R3006 GNDA.n161 GNDA.n128 53.3664
R3007 GNDA.n168 GNDA.n167 53.3664
R3008 GNDA.n187 GNDA.n186 53.3664
R3009 GNDA.n184 GNDA.n183 53.3664
R3010 GNDA.n177 GNDA.n124 53.3664
R3011 GNDA.n176 GNDA.n175 53.3664
R3012 GNDA.n121 GNDA.n118 53.3664
R3013 GNDA.n2128 GNDA.n2127 53.3664
R3014 GNDA.n116 GNDA.n113 53.3664
R3015 GNDA.n2141 GNDA.n2140 53.3664
R3016 GNDA.n457 GNDA.n450 53.3664
R3017 GNDA.n1666 GNDA.n1665 53.3664
R3018 GNDA.n448 GNDA.n442 53.3664
R3019 GNDA.n1676 GNDA.n1675 53.3664
R3020 GNDA.n541 GNDA.n540 53.3664
R3021 GNDA.n529 GNDA.n525 53.3664
R3022 GNDA.n528 GNDA.n368 53.3664
R3023 GNDA.n1730 GNDA.n1729 53.3664
R3024 GNDA.n1289 GNDA.n1288 53.3664
R3025 GNDA.n1280 GNDA.n1186 53.3664
R3026 GNDA.n1278 GNDA.n1277 53.3664
R3027 GNDA.n1269 GNDA.n1195 53.3664
R3028 GNDA.n1254 GNDA.n1253 53.3664
R3029 GNDA.n1259 GNDA.n1258 53.3664
R3030 GNDA.n1262 GNDA.n1261 53.3664
R3031 GNDA.n1267 GNDA.n1266 53.3664
R3032 GNDA.n1235 GNDA.n1234 53.3664
R3033 GNDA.n1238 GNDA.n1237 53.3664
R3034 GNDA.n1243 GNDA.n1242 53.3664
R3035 GNDA.n1246 GNDA.n1245 53.3664
R3036 GNDA.n1229 GNDA.n1211 53.3664
R3037 GNDA.n1228 GNDA.n1227 53.3664
R3038 GNDA.n1221 GNDA.n1213 53.3664
R3039 GNDA.n1220 GNDA.n1219 53.3664
R3040 GNDA.n1219 GNDA.n1218 53.3664
R3041 GNDA.n1222 GNDA.n1221 53.3664
R3042 GNDA.n1227 GNDA.n1226 53.3664
R3043 GNDA.n1230 GNDA.n1229 53.3664
R3044 GNDA.n1236 GNDA.n1235 53.3664
R3045 GNDA.n1237 GNDA.n1209 53.3664
R3046 GNDA.n1244 GNDA.n1243 53.3664
R3047 GNDA.n1245 GNDA.n1207 53.3664
R3048 GNDA.n1268 GNDA.n1267 53.3664
R3049 GNDA.n1261 GNDA.n1203 53.3664
R3050 GNDA.n1260 GNDA.n1259 53.3664
R3051 GNDA.n1253 GNDA.n1205 53.3664
R3052 GNDA.n1079 GNDA.n1078 53.3664
R3053 GNDA.n1070 GNDA.n974 53.3664
R3054 GNDA.n1068 GNDA.n1067 53.3664
R3055 GNDA.n1059 GNDA.n983 53.3664
R3056 GNDA.n1044 GNDA.n1043 53.3664
R3057 GNDA.n1049 GNDA.n1048 53.3664
R3058 GNDA.n1052 GNDA.n1051 53.3664
R3059 GNDA.n1057 GNDA.n1056 53.3664
R3060 GNDA.n1025 GNDA.n1024 53.3664
R3061 GNDA.n1028 GNDA.n1027 53.3664
R3062 GNDA.n1033 GNDA.n1032 53.3664
R3063 GNDA.n1036 GNDA.n1035 53.3664
R3064 GNDA.n1019 GNDA.n1001 53.3664
R3065 GNDA.n1018 GNDA.n1017 53.3664
R3066 GNDA.n1011 GNDA.n1003 53.3664
R3067 GNDA.n1010 GNDA.n1009 53.3664
R3068 GNDA.n1009 GNDA.n1008 53.3664
R3069 GNDA.n1012 GNDA.n1011 53.3664
R3070 GNDA.n1017 GNDA.n1016 53.3664
R3071 GNDA.n1020 GNDA.n1019 53.3664
R3072 GNDA.n1026 GNDA.n1025 53.3664
R3073 GNDA.n1027 GNDA.n999 53.3664
R3074 GNDA.n1034 GNDA.n1033 53.3664
R3075 GNDA.n1035 GNDA.n997 53.3664
R3076 GNDA.n1058 GNDA.n1057 53.3664
R3077 GNDA.n1051 GNDA.n993 53.3664
R3078 GNDA.n1050 GNDA.n1049 53.3664
R3079 GNDA.n1043 GNDA.n995 53.3664
R3080 GNDA.n1935 GNDA.n1934 53.3664
R3081 GNDA.n1926 GNDA.n301 53.3664
R3082 GNDA.n1924 GNDA.n1923 53.3664
R3083 GNDA.n1915 GNDA.n310 53.3664
R3084 GNDA.n1900 GNDA.n1899 53.3664
R3085 GNDA.n1905 GNDA.n1904 53.3664
R3086 GNDA.n1908 GNDA.n1907 53.3664
R3087 GNDA.n1913 GNDA.n1912 53.3664
R3088 GNDA.n1881 GNDA.n1880 53.3664
R3089 GNDA.n1884 GNDA.n1883 53.3664
R3090 GNDA.n1889 GNDA.n1888 53.3664
R3091 GNDA.n1892 GNDA.n1891 53.3664
R3092 GNDA.n1875 GNDA.n1857 53.3664
R3093 GNDA.n1874 GNDA.n1873 53.3664
R3094 GNDA.n1867 GNDA.n1859 53.3664
R3095 GNDA.n1866 GNDA.n1865 53.3664
R3096 GNDA.n1865 GNDA.n1864 53.3664
R3097 GNDA.n1868 GNDA.n1867 53.3664
R3098 GNDA.n1873 GNDA.n1872 53.3664
R3099 GNDA.n1876 GNDA.n1875 53.3664
R3100 GNDA.n1882 GNDA.n1881 53.3664
R3101 GNDA.n1883 GNDA.n1855 53.3664
R3102 GNDA.n1890 GNDA.n1889 53.3664
R3103 GNDA.n1891 GNDA.n1853 53.3664
R3104 GNDA.n1914 GNDA.n1913 53.3664
R3105 GNDA.n1907 GNDA.n1849 53.3664
R3106 GNDA.n1906 GNDA.n1905 53.3664
R3107 GNDA.n1899 GNDA.n1851 53.3664
R3108 GNDA.n310 GNDA.n303 53.3664
R3109 GNDA.n1925 GNDA.n1924 53.3664
R3110 GNDA.n301 GNDA.n294 53.3664
R3111 GNDA.n1936 GNDA.n1935 53.3664
R3112 GNDA.n983 GNDA.n976 53.3664
R3113 GNDA.n1069 GNDA.n1068 53.3664
R3114 GNDA.n974 GNDA.n967 53.3664
R3115 GNDA.n1080 GNDA.n1079 53.3664
R3116 GNDA.n1195 GNDA.n1188 53.3664
R3117 GNDA.n1279 GNDA.n1278 53.3664
R3118 GNDA.n1186 GNDA.n1181 53.3664
R3119 GNDA.n1290 GNDA.n1289 53.3664
R3120 GNDA.n680 GNDA.n679 53.3664
R3121 GNDA.n671 GNDA.n580 53.3664
R3122 GNDA.n669 GNDA.n668 53.3664
R3123 GNDA.n660 GNDA.n591 53.3664
R3124 GNDA.n645 GNDA.n644 53.3664
R3125 GNDA.n650 GNDA.n649 53.3664
R3126 GNDA.n653 GNDA.n652 53.3664
R3127 GNDA.n658 GNDA.n657 53.3664
R3128 GNDA.n626 GNDA.n625 53.3664
R3129 GNDA.n629 GNDA.n628 53.3664
R3130 GNDA.n634 GNDA.n633 53.3664
R3131 GNDA.n637 GNDA.n636 53.3664
R3132 GNDA.n620 GNDA.n602 53.3664
R3133 GNDA.n619 GNDA.n618 53.3664
R3134 GNDA.n612 GNDA.n604 53.3664
R3135 GNDA.n611 GNDA.n610 53.3664
R3136 GNDA.n610 GNDA.n609 53.3664
R3137 GNDA.n613 GNDA.n612 53.3664
R3138 GNDA.n618 GNDA.n617 53.3664
R3139 GNDA.n621 GNDA.n620 53.3664
R3140 GNDA.n627 GNDA.n626 53.3664
R3141 GNDA.n628 GNDA.n600 53.3664
R3142 GNDA.n635 GNDA.n634 53.3664
R3143 GNDA.n636 GNDA.n598 53.3664
R3144 GNDA.n659 GNDA.n658 53.3664
R3145 GNDA.n652 GNDA.n594 53.3664
R3146 GNDA.n651 GNDA.n650 53.3664
R3147 GNDA.n644 GNDA.n596 53.3664
R3148 GNDA.n1527 GNDA.n1526 53.3664
R3149 GNDA.n1518 GNDA.n874 53.3664
R3150 GNDA.n1516 GNDA.n1515 53.3664
R3151 GNDA.n1507 GNDA.n883 53.3664
R3152 GNDA.n1492 GNDA.n1491 53.3664
R3153 GNDA.n1497 GNDA.n1496 53.3664
R3154 GNDA.n1500 GNDA.n1499 53.3664
R3155 GNDA.n1505 GNDA.n1504 53.3664
R3156 GNDA.n1473 GNDA.n1472 53.3664
R3157 GNDA.n1476 GNDA.n1475 53.3664
R3158 GNDA.n1481 GNDA.n1480 53.3664
R3159 GNDA.n1484 GNDA.n1483 53.3664
R3160 GNDA.n1467 GNDA.n1449 53.3664
R3161 GNDA.n1466 GNDA.n1465 53.3664
R3162 GNDA.n1459 GNDA.n1451 53.3664
R3163 GNDA.n1458 GNDA.n1457 53.3664
R3164 GNDA.n1457 GNDA.n1456 53.3664
R3165 GNDA.n1460 GNDA.n1459 53.3664
R3166 GNDA.n1465 GNDA.n1464 53.3664
R3167 GNDA.n1468 GNDA.n1467 53.3664
R3168 GNDA.n1474 GNDA.n1473 53.3664
R3169 GNDA.n1475 GNDA.n1447 53.3664
R3170 GNDA.n1482 GNDA.n1481 53.3664
R3171 GNDA.n1483 GNDA.n1445 53.3664
R3172 GNDA.n1506 GNDA.n1505 53.3664
R3173 GNDA.n1499 GNDA.n1441 53.3664
R3174 GNDA.n1498 GNDA.n1497 53.3664
R3175 GNDA.n1491 GNDA.n1443 53.3664
R3176 GNDA.n2048 GNDA.n242 53.3664
R3177 GNDA.n2031 GNDA.n241 53.3664
R3178 GNDA.n2038 GNDA.n240 53.3664
R3179 GNDA.n239 GNDA.n225 53.3664
R3180 GNDA.n1981 GNDA.n233 53.3664
R3181 GNDA.n1977 GNDA.n235 53.3664
R3182 GNDA.n1973 GNDA.n237 53.3664
R3183 GNDA.n2058 GNDA.n226 53.3664
R3184 GNDA.n2001 GNDA.n229 53.3664
R3185 GNDA.n1997 GNDA.n230 53.3664
R3186 GNDA.n1993 GNDA.n231 53.3664
R3187 GNDA.n1989 GNDA.n232 53.3664
R3188 GNDA.n2002 GNDA.n228 53.3664
R3189 GNDA.n2006 GNDA.n234 53.3664
R3190 GNDA.n2010 GNDA.n236 53.3664
R3191 GNDA.n2014 GNDA.n238 53.3664
R3192 GNDA.n2016 GNDA.n238 53.3664
R3193 GNDA.n2013 GNDA.n236 53.3664
R3194 GNDA.n2009 GNDA.n234 53.3664
R3195 GNDA.n2005 GNDA.n228 53.3664
R3196 GNDA.n1998 GNDA.n229 53.3664
R3197 GNDA.n1994 GNDA.n230 53.3664
R3198 GNDA.n1990 GNDA.n231 53.3664
R3199 GNDA.n1986 GNDA.n232 53.3664
R3200 GNDA.n2059 GNDA.n2058 53.3664
R3201 GNDA.n1970 GNDA.n237 53.3664
R3202 GNDA.n1974 GNDA.n235 53.3664
R3203 GNDA.n1978 GNDA.n233 53.3664
R3204 GNDA.n2037 GNDA.n239 53.3664
R3205 GNDA.n2032 GNDA.n240 53.3664
R3206 GNDA.n2047 GNDA.n241 53.3664
R3207 GNDA.n244 GNDA.n242 53.3664
R3208 GNDA.n883 GNDA.n876 53.3664
R3209 GNDA.n1517 GNDA.n1516 53.3664
R3210 GNDA.n874 GNDA.n867 53.3664
R3211 GNDA.n1528 GNDA.n1527 53.3664
R3212 GNDA.n591 GNDA.n582 53.3664
R3213 GNDA.n670 GNDA.n669 53.3664
R3214 GNDA.n580 GNDA.n573 53.3664
R3215 GNDA.n681 GNDA.n680 53.3664
R3216 GNDA.n2357 GNDA.t222 53.2877
R3217 GNDA.t335 GNDA.t268 52.4707
R3218 GNDA.t50 GNDA.t132 52.4707
R3219 GNDA.t212 GNDA.t25 52.4707
R3220 GNDA.n27 GNDA.n20 51.2005
R3221 GNDA.n32 GNDA.n22 51.2005
R3222 GNDA.n2360 GNDA.n2337 51.2005
R3223 GNDA.n2478 GNDA.n2476 51.2005
R3224 GNDA.n832 GNDA.n92 50.9355
R3225 GNDA.n1770 GNDA.n1769 50.5752
R3226 GNDA.n2158 GNDA.n2157 50.1429
R3227 GNDA.t260 GNDA.t312 50.1429
R3228 GNDA.t354 GNDA.t31 50.1429
R3229 GNDA.n2208 GNDA.n2207 50.1429
R3230 GNDA.n2497 GNDA.t172 48.7228
R3231 GNDA.n2321 GNDA.t317 48.5574
R3232 GNDA.n2456 GNDA.t287 48.5574
R3233 GNDA.n2151 GNDA.t137 48.2626
R3234 GNDA.n2294 GNDA.t81 48.0005
R3235 GNDA.n2294 GNDA.t311 48.0005
R3236 GNDA.n2291 GNDA.t45 48.0005
R3237 GNDA.n2291 GNDA.t325 48.0005
R3238 GNDA.n2290 GNDA.t269 48.0005
R3239 GNDA.n2290 GNDA.t295 48.0005
R3240 GNDA.n2288 GNDA.t65 48.0005
R3241 GNDA.n2288 GNDA.t265 48.0005
R3242 GNDA.n2287 GNDA.t342 48.0005
R3243 GNDA.n2287 GNDA.t249 48.0005
R3244 GNDA.t137 GNDA.n318 47.9486
R3245 GNDA.t137 GNDA.n213 47.9486
R3246 GNDA.n2099 GNDA.t137 47.9486
R3247 GNDA.n273 GNDA.t137 47.6748
R3248 GNDA.t226 GNDA.t157 47.009
R3249 GNDA.t40 GNDA.t327 47.009
R3250 GNDA.t318 GNDA.t10 47.009
R3251 GNDA.t160 GNDA.t319 47.009
R3252 GNDA.n1163 GNDA.n1144 46.1628
R3253 GNDA.n1757 GNDA.n350 46.1628
R3254 GNDA.n759 GNDA.n758 46.1628
R3255 GNDA.t321 GNDA.t238 44.9749
R3256 GNDA.t330 GNDA.t278 44.9749
R3257 GNDA.t54 GNDA.t3 44.9749
R3258 GNDA.t332 GNDA.t299 44.9749
R3259 GNDA.t234 GNDA.t230 44.9749
R3260 GNDA.t60 GNDA.t303 44.9749
R3261 GNDA.t233 GNDA.t112 44.9749
R3262 GNDA.t334 GNDA.t87 44.9749
R3263 GNDA.t63 GNDA.t282 44.9749
R3264 GNDA.t215 GNDA.t70 44.9749
R3265 GNDA.n2370 GNDA.n2319 44.8222
R3266 GNDA.n2465 GNDA.n2463 44.8222
R3267 GNDA.n1832 GNDA.t137 43.8679
R3268 GNDA.n2074 GNDA.t137 43.8679
R3269 GNDA.n2102 GNDA.t137 43.8679
R3270 GNDA.n2352 GNDA.t250 43.1378
R3271 GNDA.n1724 GNDA.n371 43.0993
R3272 GNDA.t105 GNDA.n2282 41.2271
R3273 GNDA.n2490 GNDA.t103 41.2271
R3274 GNDA.n2305 GNDA.t89 41.2271
R3275 GNDA.t23 GNDA.n2496 41.2271
R3276 GNDA.n2496 GNDA.t218 41.2271
R3277 GNDA.t78 GNDA.t16 41.0871
R3278 GNDA.t78 GNDA.t66 41.0871
R3279 GNDA.t52 GNDA.t274 41.0871
R3280 GNDA.t349 GNDA.t52 41.0871
R3281 GNDA.t240 GNDA.t34 40.7412
R3282 GNDA.t76 GNDA.t326 40.7412
R3283 GNDA.t296 GNDA.t12 40.7412
R3284 GNDA.t72 GNDA.t83 40.7412
R3285 GNDA.n2472 GNDA.t323 40.7412
R3286 GNDA.t9 GNDA.n2464 40.7412
R3287 GNDA.n1311 GNDA.t135 38.0642
R3288 GNDA.n1348 GNDA.t135 38.0642
R3289 GNDA.n744 GNDA.t135 38.0642
R3290 GNDA.n2171 GNDA.t74 37.6073
R3291 GNDA.n2176 GNDA.t320 37.6073
R3292 GNDA.n2176 GNDA.t223 37.6073
R3293 GNDA.n2188 GNDA.t118 37.6073
R3294 GNDA.n2188 GNDA.t275 37.6073
R3295 GNDA.t49 GNDA.n2187 37.6073
R3296 GNDA.t139 GNDA.t209 37.4792
R3297 GNDA.t28 GNDA.t126 37.4792
R3298 GNDA.t18 GNDA.t148 37.4792
R3299 GNDA.t111 GNDA.t248 37.4792
R3300 GNDA.t264 GNDA.t20 37.4792
R3301 GNDA.t80 GNDA.t108 37.4792
R3302 GNDA.t102 GNDA.t310 37.4792
R3303 GNDA.t24 GNDA.t44 37.4792
R3304 GNDA.t120 GNDA.t324 37.4792
R3305 GNDA.t235 GNDA.t236 37.4792
R3306 GNDA.t89 GNDA.t321 37.4792
R3307 GNDA.n2513 GNDA.n2512 37.0317
R3308 GNDA.n2392 GNDA.n2391 36.6567
R3309 GNDA.t135 GNDA.n1310 34.8247
R3310 GNDA.t135 GNDA.n349 34.8247
R3311 GNDA.t135 GNDA.n743 34.8247
R3312 GNDA.t34 GNDA.t37 34.4734
R3313 GNDA.t37 GNDA.t76 34.4734
R3314 GNDA.n2199 GNDA.t345 34.4734
R3315 GNDA.n2199 GNDA.t56 34.4734
R3316 GNDA.t12 GNDA.t82 34.4734
R3317 GNDA.t82 GNDA.t72 34.4734
R3318 GNDA.n2472 GNDA.t244 34.4734
R3319 GNDA.n2464 GNDA.t84 34.4734
R3320 GNDA.n2283 GNDA.t105 33.7313
R3321 GNDA.n2284 GNDA.t220 33.7313
R3322 GNDA.n2442 GNDA.t341 33.7313
R3323 GNDA.n2441 GNDA.t64 33.7313
R3324 GNDA.n2300 GNDA.t114 33.7313
R3325 GNDA.t16 GNDA.n2321 33.6168
R3326 GNDA.n2456 GNDA.t349 33.6168
R3327 GNDA.n2343 GNDA.t271 32.9878
R3328 GNDA.n2364 GNDA.t243 32.9878
R3329 GNDA.t8 GNDA.t241 32.3951
R3330 GNDA.n2331 GNDA.n2330 32.0005
R3331 GNDA.n2459 GNDA.n2458 32.0005
R3332 GNDA.n418 GNDA.t137 31.6472
R3333 GNDA.t223 GNDA.n2175 31.3395
R3334 GNDA.t118 GNDA.n2184 31.3395
R3335 GNDA.t126 GNDA.t197 29.9835
R3336 GNDA.t148 GNDA.t232 29.9835
R3337 GNDA.t341 GNDA.t51 29.9835
R3338 GNDA.t248 GNDA.t59 29.9835
R3339 GNDA.t322 GNDA.t64 29.9835
R3340 GNDA.t190 GNDA.t177 29.9835
R3341 GNDA.n2430 GNDA.n2311 29.8817
R3342 GNDA.n2455 GNDA.n2453 29.8817
R3343 GNDA.n2368 GNDA.n2367 28.413
R3344 GNDA.n2461 GNDA.n2255 28.413
R3345 GNDA.t157 GNDA.t240 28.2056
R3346 GNDA.t326 GNDA.t40 28.2056
R3347 GNDA.n2174 GNDA.t184 28.2056
R3348 GNDA.n2183 GNDA.t123 28.2056
R3349 GNDA.t10 GNDA.t296 28.2056
R3350 GNDA.t83 GNDA.t160 28.2056
R3351 GNDA.n1760 GNDA.n346 28.1318
R3352 GNDA.n2373 GNDA.n2318 28.038
R3353 GNDA.n2375 GNDA.n2247 28.038
R3354 GNDA.n2364 GNDA.t222 27.9128
R3355 GNDA.n2193 GNDA.n2192 27.8193
R3356 GNDA.n2179 GNDA.n2178 27.8193
R3357 GNDA.n806 GNDA.n546 27.5561
R3358 GNDA.n1637 GNDA.n1594 27.5561
R3359 GNDA.n172 GNDA.n171 27.5561
R3360 GNDA.n1249 GNDA.n1206 27.5561
R3361 GNDA.n1039 GNDA.n996 27.5561
R3362 GNDA.n1895 GNDA.n1852 27.5561
R3363 GNDA.n640 GNDA.n597 27.5561
R3364 GNDA.n1487 GNDA.n1444 27.5561
R3365 GNDA.n1984 GNDA.n1983 27.5561
R3366 GNDA.n0 GNDA.n204 8.60107
R3367 GNDA.n1319 GNDA.n1163 26.7261
R3368 GNDA.n355 GNDA.n350 26.7261
R3369 GNDA.n2490 GNDA.t68 26.2356
R3370 GNDA.n2433 GNDA.t218 26.2356
R3371 GNDA.t317 GNDA.t343 26.1465
R3372 GNDA.t93 GNDA.t245 26.1465
R3373 GNDA.t290 GNDA.t85 26.1465
R3374 GNDA.t287 GNDA.t308 26.1465
R3375 GNDA.n2112 GNDA.t137 24.4846
R3376 GNDA.n759 GNDA.n690 24.2965
R3377 GNDA.n2229 GNDA.t13 24.0005
R3378 GNDA.n2229 GNDA.t73 24.0005
R3379 GNDA.n2227 GNDA.t294 24.0005
R3380 GNDA.n2227 GNDA.t11 24.0005
R3381 GNDA.n2225 GNDA.t92 24.0005
R3382 GNDA.n2225 GNDA.t6 24.0005
R3383 GNDA.n2223 GNDA.t337 24.0005
R3384 GNDA.n2223 GNDA.t15 24.0005
R3385 GNDA.n2221 GNDA.t57 24.0005
R3386 GNDA.n2221 GNDA.t314 24.0005
R3387 GNDA.n2219 GNDA.t329 24.0005
R3388 GNDA.n2219 GNDA.t346 24.0005
R3389 GNDA.n2217 GNDA.t352 24.0005
R3390 GNDA.n2217 GNDA.t39 24.0005
R3391 GNDA.n2215 GNDA.t117 24.0005
R3392 GNDA.n2215 GNDA.t292 24.0005
R3393 GNDA.n2213 GNDA.t41 24.0005
R3394 GNDA.n2213 GNDA.t339 24.0005
R3395 GNDA.n2212 GNDA.t35 24.0005
R3396 GNDA.n2212 GNDA.t77 24.0005
R3397 GNDA.n790 GNDA.n789 23.6449
R3398 GNDA.n1621 GNDA.n1620 23.6449
R3399 GNDA.n155 GNDA.n131 23.6449
R3400 GNDA.n1233 GNDA.n1232 23.6449
R3401 GNDA.n1023 GNDA.n1022 23.6449
R3402 GNDA.n1879 GNDA.n1878 23.6449
R3403 GNDA.n624 GNDA.n623 23.6449
R3404 GNDA.n1471 GNDA.n1470 23.6449
R3405 GNDA.n2003 GNDA.n2000 23.6449
R3406 GNDA.n2152 GNDA.n92 23.509
R3407 GNDA.n34 GNDA.n1 23.488
R3408 GNDA.t238 GNDA.t203 22.4877
R3409 GNDA.t3 GNDA.t27 22.4877
R3410 GNDA.t299 GNDA.t21 22.4877
R3411 GNDA.t230 GNDA.t109 22.4877
R3412 GNDA.t112 GNDA.t26 22.4877
R3413 GNDA.t87 GNDA.t19 22.4877
R3414 GNDA.t282 GNDA.t107 22.4877
R3415 GNDA.t70 GNDA.t101 22.4877
R3416 GNDA.t172 GNDA.t23 22.4877
R3417 GNDA.n16 GNDA.n15 22.4005
R3418 GNDA.n15 GNDA.n14 22.4005
R3419 GNDA.n2438 GNDA.n2308 22.4005
R3420 GNDA.n2436 GNDA.n2309 22.4005
R3421 GNDA.n2447 GNDA.n2270 22.4005
R3422 GNDA.n2445 GNDA.n2271 22.4005
R3423 GNDA.n2347 GNDA.n2318 22.4005
R3424 GNDA.n2467 GNDA.n2247 22.4005
R3425 GNDA.t327 GNDA.t338 21.9378
R3426 GNDA.t293 GNDA.t318 21.9378
R3427 GNDA.n1302 GNDA.t0 21.8669
R3428 GNDA.n734 GNDA.t8 21.8669
R3429 GNDA.n1762 GNDA.n1761 21.4917
R3430 GNDA.n78 GNDA.n77 21.3338
R3431 GNDA.n2194 GNDA.n79 21.3338
R3432 GNDA.n2191 GNDA.n2190 21.3338
R3433 GNDA.n63 GNDA.n62 21.3338
R3434 GNDA.n2154 GNDA.n2153 21.3338
R3435 GNDA.n82 GNDA.n81 21.3338
R3436 GNDA.n2317 GNDA.n2316 21.3338
R3437 GNDA.n2315 GNDA.n2314 21.3338
R3438 GNDA.n10 GNDA.n9 21.3338
R3439 GNDA.n14 GNDA.n13 21.3338
R3440 GNDA.n16 GNDA.n12 21.3338
R3441 GNDA.n17 GNDA.n11 21.3338
R3442 GNDA.n33 GNDA.n30 21.3338
R3443 GNDA.n32 GNDA.n31 21.3338
R3444 GNDA.n22 GNDA.n21 21.3338
R3445 GNDA.n20 GNDA.n19 21.3338
R3446 GNDA.n27 GNDA.n26 21.3338
R3447 GNDA.n28 GNDA.n25 21.3338
R3448 GNDA.n2277 GNDA.n2276 21.3338
R3449 GNDA.n2280 GNDA.n2278 21.3338
R3450 GNDA.n2324 GNDA.n2323 21.3338
R3451 GNDA.n2327 GNDA.n2325 21.3338
R3452 GNDA.n2258 GNDA.n2256 21.3338
R3453 GNDA.n2253 GNDA.n2252 21.3338
R3454 GNDA.n2263 GNDA.n2262 21.3338
R3455 GNDA.n2261 GNDA.n2260 21.3338
R3456 GNDA.n2211 GNDA.n2210 21.1792
R3457 GNDA.n2343 GNDA.n2342 20.3004
R3458 GNDA.n2511 GNDA.t252 19.7005
R3459 GNDA.n2511 GNDA.t17 19.7005
R3460 GNDA.n2509 GNDA.t261 19.7005
R3461 GNDA.n2509 GNDA.t46 19.7005
R3462 GNDA.n2507 GNDA.t42 19.7005
R3463 GNDA.n2507 GNDA.t284 19.7005
R3464 GNDA.n2505 GNDA.t315 19.7005
R3465 GNDA.n2505 GNDA.t48 19.7005
R3466 GNDA.n2503 GNDA.t67 19.7005
R3467 GNDA.n2503 GNDA.t94 19.7005
R3468 GNDA.n2502 GNDA.t266 19.7005
R3469 GNDA.n2502 GNDA.t47 19.7005
R3470 GNDA.n2390 GNDA.t75 19.7005
R3471 GNDA.n2390 GNDA.t33 19.7005
R3472 GNDA.n2388 GNDA.t353 19.7005
R3473 GNDA.n2388 GNDA.t286 19.7005
R3474 GNDA.n2386 GNDA.t305 19.7005
R3475 GNDA.n2386 GNDA.t95 19.7005
R3476 GNDA.n2384 GNDA.t306 19.7005
R3477 GNDA.n2384 GNDA.t289 19.7005
R3478 GNDA.n2382 GNDA.t29 19.7005
R3479 GNDA.n2382 GNDA.t288 19.7005
R3480 GNDA.n2381 GNDA.t30 19.7005
R3481 GNDA.n2381 GNDA.t267 19.7005
R3482 GNDA.n339 GNDA.n338 19.4279
R3483 GNDA.n2361 GNDA.n2360 19.3505
R3484 GNDA.n2476 GNDA.n2475 19.3505
R3485 GNDA.n2493 GNDA.n2492 19.288
R3486 GNDA.n1330 GNDA.n345 19.2005
R3487 GNDA.n1761 GNDA.n342 19.2005
R3488 GNDA.n562 GNDA.n359 19.2005
R3489 GNDA.n1339 GNDA.n1338 19.2005
R3490 GNDA.n2236 GNDA.n2235 19.2005
R3491 GNDA.n2167 GNDA.n2166 19.2005
R3492 GNDA.n2362 GNDA.n2361 19.2005
R3493 GNDA.n2475 GNDA.n2474 19.2005
R3494 GNDA.n2332 GNDA.n2331 19.1005
R3495 GNDA.n2460 GNDA.n2459 19.1005
R3496 GNDA.t303 GNDA.n2301 18.7399
R3497 GNDA.n1750 GNDA.n356 18.6274
R3498 GNDA.n2355 GNDA.n40 18.0973
R3499 GNDA.n2166 GNDA.n59 17.613
R3500 GNDA.n2515 GNDA.n2514 17.508
R3501 GNDA.n1767 GNDA.n1763 17.4917
R3502 GNDA.t307 GNDA.t243 17.2554
R3503 GNDA.n1765 GNDA.n1764 16.9605
R3504 GNDA.n2086 GNDA.n210 16.9379
R3505 GNDA.n480 GNDA.n198 16.9379
R3506 GNDA.n1820 GNDA.n1819 16.9379
R3507 GNDA.n789 GNDA.n788 16.0005
R3508 GNDA.n788 GNDA.n552 16.0005
R3509 GNDA.n782 GNDA.n552 16.0005
R3510 GNDA.n782 GNDA.n781 16.0005
R3511 GNDA.n780 GNDA.n554 16.0005
R3512 GNDA.n774 GNDA.n554 16.0005
R3513 GNDA.n774 GNDA.n773 16.0005
R3514 GNDA.n790 GNDA.n550 16.0005
R3515 GNDA.n796 GNDA.n550 16.0005
R3516 GNDA.n797 GNDA.n796 16.0005
R3517 GNDA.n798 GNDA.n797 16.0005
R3518 GNDA.n798 GNDA.n548 16.0005
R3519 GNDA.n804 GNDA.n548 16.0005
R3520 GNDA.n805 GNDA.n804 16.0005
R3521 GNDA.n806 GNDA.n805 16.0005
R3522 GNDA.n812 GNDA.n546 16.0005
R3523 GNDA.n813 GNDA.n812 16.0005
R3524 GNDA.n814 GNDA.n813 16.0005
R3525 GNDA.n814 GNDA.n544 16.0005
R3526 GNDA.n820 GNDA.n544 16.0005
R3527 GNDA.n821 GNDA.n820 16.0005
R3528 GNDA.n822 GNDA.n821 16.0005
R3529 GNDA.n822 GNDA.n542 16.0005
R3530 GNDA.n1620 GNDA.n1619 16.0005
R3531 GNDA.n1619 GNDA.n1600 16.0005
R3532 GNDA.n1613 GNDA.n1600 16.0005
R3533 GNDA.n1613 GNDA.n1612 16.0005
R3534 GNDA.n1611 GNDA.n1602 16.0005
R3535 GNDA.n1605 GNDA.n1602 16.0005
R3536 GNDA.n1605 GNDA.n1604 16.0005
R3537 GNDA.n1621 GNDA.n1598 16.0005
R3538 GNDA.n1627 GNDA.n1598 16.0005
R3539 GNDA.n1628 GNDA.n1627 16.0005
R3540 GNDA.n1629 GNDA.n1628 16.0005
R3541 GNDA.n1629 GNDA.n1596 16.0005
R3542 GNDA.n1635 GNDA.n1596 16.0005
R3543 GNDA.n1636 GNDA.n1635 16.0005
R3544 GNDA.n1637 GNDA.n1636 16.0005
R3545 GNDA.n1643 GNDA.n1594 16.0005
R3546 GNDA.n1644 GNDA.n1643 16.0005
R3547 GNDA.n1645 GNDA.n1644 16.0005
R3548 GNDA.n1645 GNDA.n1592 16.0005
R3549 GNDA.n1651 GNDA.n1592 16.0005
R3550 GNDA.n1652 GNDA.n1651 16.0005
R3551 GNDA.n1653 GNDA.n1652 16.0005
R3552 GNDA.n1653 GNDA.n1590 16.0005
R3553 GNDA.n149 GNDA.n131 16.0005
R3554 GNDA.n149 GNDA.n148 16.0005
R3555 GNDA.n148 GNDA.n147 16.0005
R3556 GNDA.n147 GNDA.n133 16.0005
R3557 GNDA.n141 GNDA.n140 16.0005
R3558 GNDA.n140 GNDA.n139 16.0005
R3559 GNDA.n139 GNDA.n109 16.0005
R3560 GNDA.n156 GNDA.n155 16.0005
R3561 GNDA.n157 GNDA.n156 16.0005
R3562 GNDA.n157 GNDA.n129 16.0005
R3563 GNDA.n163 GNDA.n129 16.0005
R3564 GNDA.n164 GNDA.n163 16.0005
R3565 GNDA.n165 GNDA.n164 16.0005
R3566 GNDA.n165 GNDA.n127 16.0005
R3567 GNDA.n171 GNDA.n127 16.0005
R3568 GNDA.n173 GNDA.n172 16.0005
R3569 GNDA.n173 GNDA.n125 16.0005
R3570 GNDA.n179 GNDA.n125 16.0005
R3571 GNDA.n180 GNDA.n179 16.0005
R3572 GNDA.n181 GNDA.n180 16.0005
R3573 GNDA.n181 GNDA.n123 16.0005
R3574 GNDA.n123 GNDA.n120 16.0005
R3575 GNDA.n188 GNDA.n120 16.0005
R3576 GNDA.n1767 GNDA.n1766 16.0005
R3577 GNDA.n1766 GNDA.n1765 16.0005
R3578 GNDA.n1232 GNDA.n1231 16.0005
R3579 GNDA.n1231 GNDA.n1212 16.0005
R3580 GNDA.n1225 GNDA.n1212 16.0005
R3581 GNDA.n1225 GNDA.n1224 16.0005
R3582 GNDA.n1223 GNDA.n1214 16.0005
R3583 GNDA.n1217 GNDA.n1214 16.0005
R3584 GNDA.n1217 GNDA.n1176 16.0005
R3585 GNDA.n1233 GNDA.n1210 16.0005
R3586 GNDA.n1239 GNDA.n1210 16.0005
R3587 GNDA.n1240 GNDA.n1239 16.0005
R3588 GNDA.n1241 GNDA.n1240 16.0005
R3589 GNDA.n1241 GNDA.n1208 16.0005
R3590 GNDA.n1247 GNDA.n1208 16.0005
R3591 GNDA.n1248 GNDA.n1247 16.0005
R3592 GNDA.n1249 GNDA.n1248 16.0005
R3593 GNDA.n1255 GNDA.n1206 16.0005
R3594 GNDA.n1256 GNDA.n1255 16.0005
R3595 GNDA.n1257 GNDA.n1256 16.0005
R3596 GNDA.n1257 GNDA.n1204 16.0005
R3597 GNDA.n1263 GNDA.n1204 16.0005
R3598 GNDA.n1264 GNDA.n1263 16.0005
R3599 GNDA.n1265 GNDA.n1264 16.0005
R3600 GNDA.n1265 GNDA.n1202 16.0005
R3601 GNDA.n1022 GNDA.n1021 16.0005
R3602 GNDA.n1021 GNDA.n1002 16.0005
R3603 GNDA.n1015 GNDA.n1002 16.0005
R3604 GNDA.n1015 GNDA.n1014 16.0005
R3605 GNDA.n1013 GNDA.n1004 16.0005
R3606 GNDA.n1007 GNDA.n1004 16.0005
R3607 GNDA.n1007 GNDA.n1006 16.0005
R3608 GNDA.n1023 GNDA.n1000 16.0005
R3609 GNDA.n1029 GNDA.n1000 16.0005
R3610 GNDA.n1030 GNDA.n1029 16.0005
R3611 GNDA.n1031 GNDA.n1030 16.0005
R3612 GNDA.n1031 GNDA.n998 16.0005
R3613 GNDA.n1037 GNDA.n998 16.0005
R3614 GNDA.n1038 GNDA.n1037 16.0005
R3615 GNDA.n1039 GNDA.n1038 16.0005
R3616 GNDA.n1045 GNDA.n996 16.0005
R3617 GNDA.n1046 GNDA.n1045 16.0005
R3618 GNDA.n1047 GNDA.n1046 16.0005
R3619 GNDA.n1047 GNDA.n994 16.0005
R3620 GNDA.n1053 GNDA.n994 16.0005
R3621 GNDA.n1054 GNDA.n1053 16.0005
R3622 GNDA.n1055 GNDA.n1054 16.0005
R3623 GNDA.n1055 GNDA.n992 16.0005
R3624 GNDA.n1878 GNDA.n1877 16.0005
R3625 GNDA.n1877 GNDA.n1858 16.0005
R3626 GNDA.n1871 GNDA.n1858 16.0005
R3627 GNDA.n1871 GNDA.n1870 16.0005
R3628 GNDA.n1869 GNDA.n1860 16.0005
R3629 GNDA.n1863 GNDA.n1860 16.0005
R3630 GNDA.n1863 GNDA.n1862 16.0005
R3631 GNDA.n1879 GNDA.n1856 16.0005
R3632 GNDA.n1885 GNDA.n1856 16.0005
R3633 GNDA.n1886 GNDA.n1885 16.0005
R3634 GNDA.n1887 GNDA.n1886 16.0005
R3635 GNDA.n1887 GNDA.n1854 16.0005
R3636 GNDA.n1893 GNDA.n1854 16.0005
R3637 GNDA.n1894 GNDA.n1893 16.0005
R3638 GNDA.n1895 GNDA.n1894 16.0005
R3639 GNDA.n1901 GNDA.n1852 16.0005
R3640 GNDA.n1902 GNDA.n1901 16.0005
R3641 GNDA.n1903 GNDA.n1902 16.0005
R3642 GNDA.n1903 GNDA.n1850 16.0005
R3643 GNDA.n1909 GNDA.n1850 16.0005
R3644 GNDA.n1910 GNDA.n1909 16.0005
R3645 GNDA.n1911 GNDA.n1910 16.0005
R3646 GNDA.n1911 GNDA.n1848 16.0005
R3647 GNDA.n623 GNDA.n622 16.0005
R3648 GNDA.n622 GNDA.n603 16.0005
R3649 GNDA.n616 GNDA.n603 16.0005
R3650 GNDA.n616 GNDA.n615 16.0005
R3651 GNDA.n614 GNDA.n605 16.0005
R3652 GNDA.n608 GNDA.n605 16.0005
R3653 GNDA.n608 GNDA.n607 16.0005
R3654 GNDA.n624 GNDA.n601 16.0005
R3655 GNDA.n630 GNDA.n601 16.0005
R3656 GNDA.n631 GNDA.n630 16.0005
R3657 GNDA.n632 GNDA.n631 16.0005
R3658 GNDA.n632 GNDA.n599 16.0005
R3659 GNDA.n638 GNDA.n599 16.0005
R3660 GNDA.n639 GNDA.n638 16.0005
R3661 GNDA.n640 GNDA.n639 16.0005
R3662 GNDA.n646 GNDA.n597 16.0005
R3663 GNDA.n647 GNDA.n646 16.0005
R3664 GNDA.n648 GNDA.n647 16.0005
R3665 GNDA.n648 GNDA.n595 16.0005
R3666 GNDA.n654 GNDA.n595 16.0005
R3667 GNDA.n655 GNDA.n654 16.0005
R3668 GNDA.n656 GNDA.n655 16.0005
R3669 GNDA.n656 GNDA.n593 16.0005
R3670 GNDA.n1470 GNDA.n1469 16.0005
R3671 GNDA.n1469 GNDA.n1450 16.0005
R3672 GNDA.n1463 GNDA.n1450 16.0005
R3673 GNDA.n1463 GNDA.n1462 16.0005
R3674 GNDA.n1461 GNDA.n1452 16.0005
R3675 GNDA.n1455 GNDA.n1452 16.0005
R3676 GNDA.n1455 GNDA.n1454 16.0005
R3677 GNDA.n1471 GNDA.n1448 16.0005
R3678 GNDA.n1477 GNDA.n1448 16.0005
R3679 GNDA.n1478 GNDA.n1477 16.0005
R3680 GNDA.n1479 GNDA.n1478 16.0005
R3681 GNDA.n1479 GNDA.n1446 16.0005
R3682 GNDA.n1485 GNDA.n1446 16.0005
R3683 GNDA.n1486 GNDA.n1485 16.0005
R3684 GNDA.n1487 GNDA.n1486 16.0005
R3685 GNDA.n1493 GNDA.n1444 16.0005
R3686 GNDA.n1494 GNDA.n1493 16.0005
R3687 GNDA.n1495 GNDA.n1494 16.0005
R3688 GNDA.n1495 GNDA.n1442 16.0005
R3689 GNDA.n1501 GNDA.n1442 16.0005
R3690 GNDA.n1502 GNDA.n1501 16.0005
R3691 GNDA.n1503 GNDA.n1502 16.0005
R3692 GNDA.n1503 GNDA.n1440 16.0005
R3693 GNDA.n2004 GNDA.n2003 16.0005
R3694 GNDA.n2007 GNDA.n2004 16.0005
R3695 GNDA.n2008 GNDA.n2007 16.0005
R3696 GNDA.n2011 GNDA.n2008 16.0005
R3697 GNDA.n2015 GNDA.n2012 16.0005
R3698 GNDA.n2017 GNDA.n2015 16.0005
R3699 GNDA.n2018 GNDA.n2017 16.0005
R3700 GNDA.n2000 GNDA.n1999 16.0005
R3701 GNDA.n1999 GNDA.n1996 16.0005
R3702 GNDA.n1996 GNDA.n1995 16.0005
R3703 GNDA.n1995 GNDA.n1992 16.0005
R3704 GNDA.n1992 GNDA.n1991 16.0005
R3705 GNDA.n1991 GNDA.n1988 16.0005
R3706 GNDA.n1988 GNDA.n1987 16.0005
R3707 GNDA.n1987 GNDA.n1984 16.0005
R3708 GNDA.n1983 GNDA.n1980 16.0005
R3709 GNDA.n1980 GNDA.n1979 16.0005
R3710 GNDA.n1979 GNDA.n1976 16.0005
R3711 GNDA.n1976 GNDA.n1975 16.0005
R3712 GNDA.n1975 GNDA.n1972 16.0005
R3713 GNDA.n1972 GNDA.n1971 16.0005
R3714 GNDA.n1971 GNDA.n224 16.0005
R3715 GNDA.n2060 GNDA.n224 16.0005
R3716 GNDA.t74 GNDA.t116 15.67
R3717 GNDA.t291 GNDA.t260 15.67
R3718 GNDA.t31 GNDA.t91 15.67
R3719 GNDA.t5 GNDA.t49 15.67
R3720 GNDA.n2204 GNDA.n2203 15.363
R3721 GNDA.n2203 GNDA.n68 15.363
R3722 GNDA.t197 GNDA.t18 14.992
R3723 GNDA.t232 GNDA.t106 14.992
R3724 GNDA.t51 GNDA.t111 14.992
R3725 GNDA.t59 GNDA.t22 14.992
R3726 GNDA.t20 GNDA.t322 14.992
R3727 GNDA.t206 GNDA.t264 14.992
R3728 GNDA.t331 GNDA.t206 14.992
R3729 GNDA.t108 GNDA.t331 14.992
R3730 GNDA.t276 GNDA.t80 14.992
R3731 GNDA.t55 GNDA.t276 14.992
R3732 GNDA.t310 GNDA.t1 14.992
R3733 GNDA.t1 GNDA.t333 14.992
R3734 GNDA.t333 GNDA.t24 14.992
R3735 GNDA.t44 GNDA.t297 14.992
R3736 GNDA.t297 GNDA.t62 14.992
R3737 GNDA.t62 GNDA.t120 14.992
R3738 GNDA.t324 GNDA.t228 14.992
R3739 GNDA.t228 GNDA.t335 14.992
R3740 GNDA.t268 GNDA.t301 14.992
R3741 GNDA.t301 GNDA.t50 14.992
R3742 GNDA.t132 GNDA.t280 14.992
R3743 GNDA.t280 GNDA.t212 14.992
R3744 GNDA.t25 GNDA.t68 14.992
R3745 GNDA.t114 GNDA.t103 14.992
R3746 GNDA.t236 GNDA.t190 14.992
R3747 GNDA.t203 GNDA.t330 14.992
R3748 GNDA.t104 GNDA.t54 14.992
R3749 GNDA.t27 GNDA.t332 14.992
R3750 GNDA.t21 GNDA.t234 14.992
R3751 GNDA.t109 GNDA.t60 14.992
R3752 GNDA.t26 GNDA.t334 14.992
R3753 GNDA.t19 GNDA.t63 14.992
R3754 GNDA.t107 GNDA.t215 14.992
R3755 GNDA.n2453 GNDA.n2452 14.9411
R3756 GNDA.n339 GNDA 14.6989
R3757 GNDA.n2427 GNDA.n2426 14.0505
R3758 GNDA.n2378 GNDA.n2377 14.0505
R3759 GNDA GNDA.n780 14.0449
R3760 GNDA GNDA.n1611 14.0449
R3761 GNDA.n141 GNDA 14.0449
R3762 GNDA GNDA.n1223 14.0449
R3763 GNDA GNDA.n1013 14.0449
R3764 GNDA GNDA.n1869 14.0449
R3765 GNDA GNDA.n614 14.0449
R3766 GNDA GNDA.n1461 14.0449
R3767 GNDA.n2012 GNDA 14.0449
R3768 GNDA.n2501 GNDA.n2500 14.0193
R3769 GNDA.n1686 GNDA.n418 13.9984
R3770 GNDA.n2235 GNDA.n2234 13.8005
R3771 GNDA.n2421 GNDA.n2309 13.8005
R3772 GNDA.n2398 GNDA.n2308 13.8005
R3773 GNDA.n2397 GNDA.n2271 13.8005
R3774 GNDA.n2394 GNDA.n2270 13.8005
R3775 GNDA.n1336 GNDA.n1138 13.7682
R3776 GNDA.n742 GNDA.n729 13.7682
R3777 GNDA.n1763 GNDA.n60 13.4945
R3778 GNDA.n1335 GNDA.t0 12.9584
R3779 GNDA.n1690 GNDA.n413 12.9309
R3780 GNDA.n502 GNDA.n248 12.9309
R3781 GNDA.n926 GNDA.n286 12.9309
R3782 GNDA.n1385 GNDA.n1092 12.9309
R3783 GNDA.n2171 GNDA.n90 12.5361
R3784 GNDA.n2187 GNDA.n2186 12.5361
R3785 GNDA.n756 GNDA.n755 12.4126
R3786 GNDA.n1323 GNDA.n1322 12.4126
R3787 GNDA.n1360 GNDA.n1359 12.4126
R3788 GNDA.n2086 GNDA.n2085 11.6369
R3789 GNDA.n2085 GNDA.n2084 11.6369
R3790 GNDA.n2084 GNDA.n211 11.6369
R3791 GNDA.n2078 GNDA.n211 11.6369
R3792 GNDA.n2078 GNDA.n2077 11.6369
R3793 GNDA.n2077 GNDA.n2076 11.6369
R3794 GNDA.n2076 GNDA.n215 11.6369
R3795 GNDA.n2070 GNDA.n215 11.6369
R3796 GNDA.n2070 GNDA.n2069 11.6369
R3797 GNDA.n925 GNDA.n897 11.6369
R3798 GNDA.n899 GNDA.n897 11.6369
R3799 GNDA.n918 GNDA.n899 11.6369
R3800 GNDA.n918 GNDA.n917 11.6369
R3801 GNDA.n917 GNDA.n916 11.6369
R3802 GNDA.n916 GNDA.n901 11.6369
R3803 GNDA.n911 GNDA.n901 11.6369
R3804 GNDA.n911 GNDA.n910 11.6369
R3805 GNDA.n910 GNDA.n909 11.6369
R3806 GNDA.n909 GNDA.n904 11.6369
R3807 GNDA.n904 GNDA.n210 11.6369
R3808 GNDA.n755 GNDA.n754 11.6369
R3809 GNDA.n754 GNDA.n723 11.6369
R3810 GNDA.n748 GNDA.n723 11.6369
R3811 GNDA.n748 GNDA.n747 11.6369
R3812 GNDA.n747 GNDA.n746 11.6369
R3813 GNDA.n746 GNDA.n727 11.6369
R3814 GNDA.n740 GNDA.n739 11.6369
R3815 GNDA.n739 GNDA.n738 11.6369
R3816 GNDA.n722 GNDA.n721 11.6369
R3817 GNDA.n721 GNDA.n694 11.6369
R3818 GNDA.n716 GNDA.n694 11.6369
R3819 GNDA.n716 GNDA.n715 11.6369
R3820 GNDA.n715 GNDA.n714 11.6369
R3821 GNDA.n714 GNDA.n697 11.6369
R3822 GNDA.n709 GNDA.n697 11.6369
R3823 GNDA.n709 GNDA.n708 11.6369
R3824 GNDA.n708 GNDA.n707 11.6369
R3825 GNDA.n707 GNDA.n700 11.6369
R3826 GNDA.n702 GNDA.n700 11.6369
R3827 GNDA.n1541 GNDA.n1540 11.6369
R3828 GNDA.n1542 GNDA.n1541 11.6369
R3829 GNDA.n1542 GNDA.n508 11.6369
R3830 GNDA.n1548 GNDA.n508 11.6369
R3831 GNDA.n1549 GNDA.n1548 11.6369
R3832 GNDA.n1550 GNDA.n1549 11.6369
R3833 GNDA.n1550 GNDA.n506 11.6369
R3834 GNDA.n1556 GNDA.n506 11.6369
R3835 GNDA.n1557 GNDA.n1556 11.6369
R3836 GNDA.n1558 GNDA.n1557 11.6369
R3837 GNDA.n1558 GNDA.n503 11.6369
R3838 GNDA.n501 GNDA.n471 11.6369
R3839 GNDA.n496 GNDA.n471 11.6369
R3840 GNDA.n496 GNDA.n495 11.6369
R3841 GNDA.n495 GNDA.n474 11.6369
R3842 GNDA.n490 GNDA.n474 11.6369
R3843 GNDA.n490 GNDA.n489 11.6369
R3844 GNDA.n489 GNDA.n488 11.6369
R3845 GNDA.n488 GNDA.n476 11.6369
R3846 GNDA.n482 GNDA.n476 11.6369
R3847 GNDA.n482 GNDA.n481 11.6369
R3848 GNDA.n481 GNDA.n480 11.6369
R3849 GNDA.n2092 GNDA.n198 11.6369
R3850 GNDA.n2093 GNDA.n2092 11.6369
R3851 GNDA.n2095 GNDA.n2093 11.6369
R3852 GNDA.n2095 GNDA.n2094 11.6369
R3853 GNDA.n2094 GNDA.n195 11.6369
R3854 GNDA.n195 GNDA.n193 11.6369
R3855 GNDA.n2106 GNDA.n193 11.6369
R3856 GNDA.n2107 GNDA.n2106 11.6369
R3857 GNDA.n2108 GNDA.n2107 11.6369
R3858 GNDA.n1819 GNDA.n1805 11.6369
R3859 GNDA.n1813 GNDA.n1805 11.6369
R3860 GNDA.n1813 GNDA.n1812 11.6369
R3861 GNDA.n1812 GNDA.n1811 11.6369
R3862 GNDA.n1811 GNDA.n316 11.6369
R3863 GNDA.n1834 GNDA.n316 11.6369
R3864 GNDA.n1835 GNDA.n1834 11.6369
R3865 GNDA.n1837 GNDA.n1835 11.6369
R3866 GNDA.n1837 GNDA.n1836 11.6369
R3867 GNDA.n1703 GNDA.n386 11.6369
R3868 GNDA.n1703 GNDA.n1702 11.6369
R3869 GNDA.n1702 GNDA.n1701 11.6369
R3870 GNDA.n1701 GNDA.n1698 11.6369
R3871 GNDA.n1698 GNDA.n334 11.6369
R3872 GNDA.n1776 GNDA.n332 11.6369
R3873 GNDA.n1777 GNDA.n1776 11.6369
R3874 GNDA.n1778 GNDA.n1777 11.6369
R3875 GNDA.n1778 GNDA.n327 11.6369
R3876 GNDA.n1784 GNDA.n327 11.6369
R3877 GNDA.n1792 GNDA.n1791 11.6369
R3878 GNDA.n1793 GNDA.n1792 11.6369
R3879 GNDA.n1793 GNDA.n323 11.6369
R3880 GNDA.n1799 GNDA.n323 11.6369
R3881 GNDA.n1800 GNDA.n1799 11.6369
R3882 GNDA.n1829 GNDA.n1800 11.6369
R3883 GNDA.n1829 GNDA.n1828 11.6369
R3884 GNDA.n1828 GNDA.n1827 11.6369
R3885 GNDA.n1827 GNDA.n1801 11.6369
R3886 GNDA.n1821 GNDA.n1801 11.6369
R3887 GNDA.n1821 GNDA.n1820 11.6369
R3888 GNDA.n1389 GNDA.n1388 11.6369
R3889 GNDA.n1390 GNDA.n1389 11.6369
R3890 GNDA.n1390 GNDA.n932 11.6369
R3891 GNDA.n1396 GNDA.n932 11.6369
R3892 GNDA.n1397 GNDA.n1396 11.6369
R3893 GNDA.n1398 GNDA.n1397 11.6369
R3894 GNDA.n1398 GNDA.n930 11.6369
R3895 GNDA.n1404 GNDA.n930 11.6369
R3896 GNDA.n1405 GNDA.n1404 11.6369
R3897 GNDA.n1406 GNDA.n1405 11.6369
R3898 GNDA.n1406 GNDA.n927 11.6369
R3899 GNDA.n1159 GNDA.n1158 11.6369
R3900 GNDA.n1158 GNDA.n1147 11.6369
R3901 GNDA.n1152 GNDA.n1147 11.6369
R3902 GNDA.n1152 GNDA.n1151 11.6369
R3903 GNDA.n1151 GNDA.n381 11.6369
R3904 GNDA.n1720 GNDA.n381 11.6369
R3905 GNDA.n1720 GNDA.n1719 11.6369
R3906 GNDA.n1719 GNDA.n1718 11.6369
R3907 GNDA.n1718 GNDA.n382 11.6369
R3908 GNDA.n1712 GNDA.n382 11.6369
R3909 GNDA.n1712 GNDA.n1711 11.6369
R3910 GNDA.n1322 GNDA.n1321 11.6369
R3911 GNDA.n1321 GNDA.n1160 11.6369
R3912 GNDA.n1315 GNDA.n1160 11.6369
R3913 GNDA.n1315 GNDA.n1314 11.6369
R3914 GNDA.n1314 GNDA.n1313 11.6369
R3915 GNDA.n1313 GNDA.n1166 11.6369
R3916 GNDA.n1307 GNDA.n1306 11.6369
R3917 GNDA.n1306 GNDA.n1305 11.6369
R3918 GNDA.n1361 GNDA.n1126 11.6369
R3919 GNDA.n1367 GNDA.n1126 11.6369
R3920 GNDA.n1368 GNDA.n1367 11.6369
R3921 GNDA.n1369 GNDA.n1368 11.6369
R3922 GNDA.n1369 GNDA.n1124 11.6369
R3923 GNDA.n1375 GNDA.n1124 11.6369
R3924 GNDA.n1376 GNDA.n1375 11.6369
R3925 GNDA.n1377 GNDA.n1376 11.6369
R3926 GNDA.n1377 GNDA.n1122 11.6369
R3927 GNDA.n1122 GNDA.n1094 11.6369
R3928 GNDA.n1384 GNDA.n1094 11.6369
R3929 GNDA.n1359 GNDA.n1128 11.6369
R3930 GNDA.n1353 GNDA.n1128 11.6369
R3931 GNDA.n1353 GNDA.n1352 11.6369
R3932 GNDA.n1352 GNDA.n1351 11.6369
R3933 GNDA.n1351 GNDA.n1345 11.6369
R3934 GNDA.n1345 GNDA.n1344 11.6369
R3935 GNDA.n1755 GNDA.n1754 11.6369
R3936 GNDA.n1754 GNDA.n1753 11.6369
R3937 GNDA.n2393 GNDA.n2392 11.6255
R3938 GNDA.n740 GNDA 11.5076
R3939 GNDA.n1307 GNDA 11.5076
R3940 GNDA.n1755 GNDA 11.5076
R3941 GNDA.n738 GNDA.n731 11.3514
R3942 GNDA.n1305 GNDA.n1170 11.3514
R3943 GNDA.n1753 GNDA.n353 11.3514
R3944 GNDA.t255 GNDA.n1335 11.3386
R3945 GNDA.n2069 GNDA.n2068 11.249
R3946 GNDA.n2108 GNDA.n189 11.249
R3947 GNDA.n1836 GNDA.n311 11.249
R3948 GNDA.n2284 GNDA.t28 11.2441
R3949 GNDA.n2274 GNDA.t55 11.2441
R3950 GNDA.t278 GNDA.n2304 11.2441
R3951 GNDA.n2304 GNDA.t104 11.2441
R3952 GNDA.t61 GNDA.t233 11.2441
R3953 GNDA.n2497 GNDA.t101 11.2441
R3954 GNDA.t316 GNDA.t99 11.2059
R3955 GNDA.t43 GNDA.t129 11.2059
R3956 GNDA.n2371 GNDA.t154 11.2059
R3957 GNDA.t151 GNDA.n2249 11.2059
R3958 GNDA.t272 GNDA.t200 11.2059
R3959 GNDA.t273 GNDA.t97 11.2059
R3960 GNDA.n1347 GNDA.n1342 10.5288
R3961 GNDA.n1764 GNDA.n332 10.4732
R3962 GNDA.n2202 GNDA.n2201 9.78488
R3963 GNDA.n58 GNDA.t225 9.6005
R3964 GNDA.n58 GNDA.t340 9.6005
R3965 GNDA.n2165 GNDA.t227 9.6005
R3966 GNDA.n2165 GNDA.t224 9.6005
R3967 GNDA.n2395 GNDA.t140 9.6005
R3968 GNDA.n2395 GNDA.t221 9.6005
R3969 GNDA.n2399 GNDA.t207 9.6005
R3970 GNDA.n2399 GNDA.t277 9.6005
R3971 GNDA.n2401 GNDA.t2 9.6005
R3972 GNDA.n2401 GNDA.t298 9.6005
R3973 GNDA.n2403 GNDA.t229 9.6005
R3974 GNDA.n2403 GNDA.t302 9.6005
R3975 GNDA.n2405 GNDA.t281 9.6005
R3976 GNDA.n2405 GNDA.t69 9.6005
R3977 GNDA.n2407 GNDA.t115 9.6005
R3978 GNDA.n2407 GNDA.t237 9.6005
R3979 GNDA.n2409 GNDA.t90 9.6005
R3980 GNDA.n2409 GNDA.t239 9.6005
R3981 GNDA.n2411 GNDA.t279 9.6005
R3982 GNDA.n2411 GNDA.t4 9.6005
R3983 GNDA.n2413 GNDA.t300 9.6005
R3984 GNDA.n2413 GNDA.t231 9.6005
R3985 GNDA.n2415 GNDA.t304 9.6005
R3986 GNDA.n2415 GNDA.t113 9.6005
R3987 GNDA.n2417 GNDA.t88 9.6005
R3988 GNDA.n2417 GNDA.t283 9.6005
R3989 GNDA.n2419 GNDA.t71 9.6005
R3990 GNDA.n2419 GNDA.t173 9.6005
R3991 GNDA.t247 GNDA.t291 9.40221
R3992 GNDA.t91 GNDA.t36 9.40221
R3993 GNDA.n2234 GNDA.n2233 9.37925
R3994 GNDA.n2297 GNDA.n2296 9.3005
R3995 GNDA.n1536 GNDA.n418 8.98697
R3996 GNDA.n756 GNDA.n722 8.66313
R3997 GNDA.n1323 GNDA.n1159 8.66313
R3998 GNDA.n1361 GNDA.n1360 8.66313
R3999 GNDA.n926 GNDA.n925 8.53383
R4000 GNDA.n1540 GNDA.n413 8.53383
R4001 GNDA.n502 GNDA.n501 8.53383
R4002 GNDA.n1710 GNDA.n386 8.53383
R4003 GNDA.n1791 GNDA.n1785 8.53383
R4004 GNDA.n1388 GNDA.n1385 8.53383
R4005 GNDA.n2231 GNDA.n2230 8.44175
R4006 GNDA.n542 GNDA.n519 8.35606
R4007 GNDA.n1590 GNDA.n1589 8.35606
R4008 GNDA.n2116 GNDA.n188 8.35606
R4009 GNDA.n1202 GNDA.n1201 8.35606
R4010 GNDA.n992 GNDA.n991 8.35606
R4011 GNDA.n1848 GNDA.n1847 8.35606
R4012 GNDA.n593 GNDA.n592 8.35606
R4013 GNDA.n1440 GNDA.n1439 8.35606
R4014 GNDA.n2061 GNDA.n2060 8.35606
R4015 GNDA.t135 GNDA.n92 8.20508
R4016 GNDA.n1695 GNDA.t137 8.20508
R4017 GNDA.n2203 GNDA.n2202 7.71925
R4018 GNDA.n2342 GNDA.t258 7.61296
R4019 GNDA.n2357 GNDA.t254 7.61296
R4020 GNDA.n1336 GNDA.t7 7.28929
R4021 GNDA.n347 GNDA.n345 6.4005
R4022 GNDA.n60 GNDA 6.04837
R4023 GNDA.n2515 GNDA 5.6875
R4024 GNDA.t7 GNDA.t255 5.66956
R4025 GNDA.n2501 GNDA.n2 5.03175
R4026 GNDA.n2392 GNDA.n2 4.90675
R4027 GNDA.t241 GNDA.n729 4.85969
R4028 GNDA.n2296 GNDA.n2 4.7505
R4029 GNDA.n770 GNDA.n557 4.6085
R4030 GNDA.n1683 GNDA.n1682 4.6085
R4031 GNDA.n2149 GNDA.n2148 4.6085
R4032 GNDA.n1297 GNDA.n1174 4.6085
R4033 GNDA.n1088 GNDA.n1087 4.6085
R4034 GNDA.n1944 GNDA.n288 4.6085
R4035 GNDA.n567 GNDA.n566 4.6085
R4036 GNDA.n860 GNDA.n416 4.6085
R4037 GNDA.n2020 GNDA.n1969 4.6085
R4038 GNDA.n857 GNDA.n856 4.55161
R4039 GNDA.n470 GNDA.n468 4.55161
R4040 GNDA.n1786 GNDA.n270 4.55161
R4041 GNDA.n1412 GNDA.n895 4.55161
R4042 GNDA.n1709 GNDA.n387 4.55161
R4043 GNDA.n1120 GNDA.n1093 4.55161
R4044 GNDA.n837 GNDA.n437 4.5061
R4045 GNDA.n1586 GNDA.n108 4.5061
R4046 GNDA.n1092 GNDA.n1091 4.5061
R4047 GNDA.n1945 GNDA.n286 4.5061
R4048 GNDA.n1690 GNDA.n1689 4.5061
R4049 GNDA.n1968 GNDA.n248 4.5061
R4050 GNDA.n2202 GNDA.n59 4.5005
R4051 GNDA.n2295 GNDA.n2293 4.5005
R4052 GNDA.n2514 GNDA.n2513 4.5005
R4053 GNDA.n2422 GNDA.n1 4.5005
R4054 GNDA.n702 GNDA.n413 4.39646
R4055 GNDA.n503 GNDA.n502 4.39646
R4056 GNDA.n1785 GNDA.n1784 4.39646
R4057 GNDA.n927 GNDA.n926 4.39646
R4058 GNDA.n1711 GNDA.n1710 4.39646
R4059 GNDA.n1385 GNDA.n1384 4.39646
R4060 GNDA.n837 GNDA.n836 4.3525
R4061 GNDA.n1587 GNDA.n1586 4.3525
R4062 GNDA.n1197 GNDA.n1092 4.3525
R4063 GNDA.n984 GNDA.n286 4.3525
R4064 GNDA.n1691 GNDA.n1690 4.3525
R4065 GNDA.n884 GNDA.n248 4.3525
R4066 GNDA.n836 GNDA.n834 4.3013
R4067 GNDA.n1588 GNDA.n1587 4.3013
R4068 GNDA.n1200 GNDA.n1197 4.3013
R4069 GNDA.n990 GNDA.n984 4.3013
R4070 GNDA.n1846 GNDA.n311 4.3013
R4071 GNDA.n1691 GNDA.n412 4.3013
R4072 GNDA.n1438 GNDA.n884 4.3013
R4073 GNDA.n2068 GNDA.n219 4.3013
R4074 GNDA.n856 GNDA.n855 4.26717
R4075 GNDA.n855 GNDA.n853 4.26717
R4076 GNDA.n853 GNDA.n850 4.26717
R4077 GNDA.n850 GNDA.n849 4.26717
R4078 GNDA.n849 GNDA.n846 4.26717
R4079 GNDA.n846 GNDA.n845 4.26717
R4080 GNDA.n842 GNDA.n841 4.26717
R4081 GNDA.n841 GNDA.n838 4.26717
R4082 GNDA.n1565 GNDA.n468 4.26717
R4083 GNDA.n1566 GNDA.n1565 4.26717
R4084 GNDA.n1569 GNDA.n1566 4.26717
R4085 GNDA.n1569 GNDA.n464 4.26717
R4086 GNDA.n1575 GNDA.n464 4.26717
R4087 GNDA.n1576 GNDA.n1575 4.26717
R4088 GNDA.n1579 GNDA.n460 4.26717
R4089 GNDA.n1585 GNDA.n460 4.26717
R4090 GNDA.n1962 GNDA.n270 4.26717
R4091 GNDA.n1962 GNDA.n271 4.26717
R4092 GNDA.n1957 GNDA.n271 4.26717
R4093 GNDA.n1957 GNDA.n1956 4.26717
R4094 GNDA.n1956 GNDA.n1955 4.26717
R4095 GNDA.n1955 GNDA.n279 4.26717
R4096 GNDA.n1950 GNDA.n1949 4.26717
R4097 GNDA.n1949 GNDA.n1948 4.26717
R4098 GNDA.n1413 GNDA.n1412 4.26717
R4099 GNDA.n1416 GNDA.n1413 4.26717
R4100 GNDA.n1416 GNDA.n891 4.26717
R4101 GNDA.n1422 GNDA.n891 4.26717
R4102 GNDA.n1423 GNDA.n1422 4.26717
R4103 GNDA.n1426 GNDA.n1423 4.26717
R4104 GNDA.n1431 GNDA.n887 4.26717
R4105 GNDA.n1432 GNDA.n1431 4.26717
R4106 GNDA.n934 GNDA.n387 4.26717
R4107 GNDA.n939 GNDA.n934 4.26717
R4108 GNDA.n940 GNDA.n939 4.26717
R4109 GNDA.n945 GNDA.n940 4.26717
R4110 GNDA.n946 GNDA.n945 4.26717
R4111 GNDA.n951 GNDA.n946 4.26717
R4112 GNDA.n957 GNDA.n952 4.26717
R4113 GNDA.n959 GNDA.n957 4.26717
R4114 GNDA.n1120 GNDA.n1119 4.26717
R4115 GNDA.n1119 GNDA.n1116 4.26717
R4116 GNDA.n1116 GNDA.n1115 4.26717
R4117 GNDA.n1115 GNDA.n1112 4.26717
R4118 GNDA.n1112 GNDA.n1111 4.26717
R4119 GNDA.n1111 GNDA.n1108 4.26717
R4120 GNDA.n1107 GNDA.n1104 4.26717
R4121 GNDA.n1104 GNDA.n414 4.26717
R4122 GNDA.n842 GNDA 4.21976
R4123 GNDA.n1579 GNDA 4.21976
R4124 GNDA.n1950 GNDA 4.21976
R4125 GNDA GNDA.n887 4.21976
R4126 GNDA.n952 GNDA 4.21976
R4127 GNDA GNDA.n1107 4.21976
R4128 GNDA.n2115 GNDA.n189 4.1989
R4129 GNDA.n838 GNDA.n837 4.12494
R4130 GNDA.n1586 GNDA.n1585 4.12494
R4131 GNDA.n1948 GNDA.n286 4.12494
R4132 GNDA.n1432 GNDA.n248 4.12494
R4133 GNDA.n1092 GNDA.n959 4.12494
R4134 GNDA.n1690 GNDA.n414 4.12494
R4135 GNDA.n2234 GNDA.n59 3.813
R4136 GNDA.n2282 GNDA.t139 3.74837
R4137 GNDA.t220 GNDA.n2283 3.74837
R4138 GNDA.n2442 GNDA.t106 3.74837
R4139 GNDA.t22 GNDA.n2441 3.74837
R4140 GNDA.n2274 GNDA.t102 3.74837
R4141 GNDA.t177 GNDA.n2300 3.74837
R4142 GNDA.n2305 GNDA.t235 3.74837
R4143 GNDA.n2301 GNDA.t110 3.74837
R4144 GNDA.t110 GNDA.t61 3.74837
R4145 GNDA.t145 GNDA.t142 3.73564
R4146 GNDA.t194 GNDA.t168 3.73564
R4147 GNDA GNDA.n2515 3.7135
R4148 GNDA.n2233 GNDA 3.68412
R4149 GNDA.n2513 GNDA.n2501 3.6255
R4150 GNDA.n1732 GNDA.n365 3.5845
R4151 GNDA.n1731 GNDA.n366 3.5845
R4152 GNDA.n1727 GNDA.n1726 3.5845
R4153 GNDA.n527 GNDA.n369 3.5845
R4154 GNDA.n532 GNDA.n531 3.5845
R4155 GNDA.n536 GNDA.n526 3.5845
R4156 GNDA.n538 GNDA.n537 3.5845
R4157 GNDA.n828 GNDA.n523 3.5845
R4158 GNDA.n827 GNDA.n524 3.5845
R4159 GNDA.n1678 GNDA.n439 3.5845
R4160 GNDA.n445 GNDA.n441 3.5845
R4161 GNDA.n1673 GNDA.n1672 3.5845
R4162 GNDA.n1669 GNDA.n446 3.5845
R4163 GNDA.n1668 GNDA.n447 3.5845
R4164 GNDA.n453 GNDA.n449 3.5845
R4165 GNDA.n1663 GNDA.n1662 3.5845
R4166 GNDA.n1659 GNDA.n454 3.5845
R4167 GNDA.n1658 GNDA.n456 3.5845
R4168 GNDA.n2143 GNDA.n110 3.5845
R4169 GNDA.n2142 GNDA.n111 3.5845
R4170 GNDA.n2138 GNDA.n2137 3.5845
R4171 GNDA.n2134 GNDA.n2133 3.5845
R4172 GNDA.n2130 GNDA.n114 3.5845
R4173 GNDA.n2129 GNDA.n115 3.5845
R4174 GNDA.n2125 GNDA.n2124 3.5845
R4175 GNDA.n2121 GNDA.n2120 3.5845
R4176 GNDA.n2117 GNDA.n119 3.5845
R4177 GNDA.n1292 GNDA.n1177 3.5845
R4178 GNDA.n1291 GNDA.n1179 3.5845
R4179 GNDA.n1287 GNDA.n1286 3.5845
R4180 GNDA.n1282 GNDA.n1182 3.5845
R4181 GNDA.n1281 GNDA.n1185 3.5845
R4182 GNDA.n1189 GNDA.n1187 3.5845
R4183 GNDA.n1276 GNDA.n1275 3.5845
R4184 GNDA.n1271 GNDA.n1190 3.5845
R4185 GNDA.n1270 GNDA.n1194 3.5845
R4186 GNDA.n1082 GNDA.n964 3.5845
R4187 GNDA.n968 GNDA.n966 3.5845
R4188 GNDA.n1077 GNDA.n1076 3.5845
R4189 GNDA.n1072 GNDA.n969 3.5845
R4190 GNDA.n1071 GNDA.n973 3.5845
R4191 GNDA.n977 GNDA.n975 3.5845
R4192 GNDA.n1066 GNDA.n1065 3.5845
R4193 GNDA.n1061 GNDA.n978 3.5845
R4194 GNDA.n1060 GNDA.n982 3.5845
R4195 GNDA.n1938 GNDA.n291 3.5845
R4196 GNDA.n295 GNDA.n293 3.5845
R4197 GNDA.n1933 GNDA.n1932 3.5845
R4198 GNDA.n1928 GNDA.n296 3.5845
R4199 GNDA.n1927 GNDA.n300 3.5845
R4200 GNDA.n304 GNDA.n302 3.5845
R4201 GNDA.n1922 GNDA.n1921 3.5845
R4202 GNDA.n1917 GNDA.n305 3.5845
R4203 GNDA.n1916 GNDA.n309 3.5845
R4204 GNDA.n683 GNDA.n570 3.5845
R4205 GNDA.n574 GNDA.n572 3.5845
R4206 GNDA.n678 GNDA.n677 3.5845
R4207 GNDA.n673 GNDA.n575 3.5845
R4208 GNDA.n672 GNDA.n579 3.5845
R4209 GNDA.n583 GNDA.n581 3.5845
R4210 GNDA.n667 GNDA.n666 3.5845
R4211 GNDA.n662 GNDA.n584 3.5845
R4212 GNDA.n661 GNDA.n590 3.5845
R4213 GNDA.n1530 GNDA.n864 3.5845
R4214 GNDA.n868 GNDA.n866 3.5845
R4215 GNDA.n1525 GNDA.n1524 3.5845
R4216 GNDA.n1520 GNDA.n869 3.5845
R4217 GNDA.n1519 GNDA.n873 3.5845
R4218 GNDA.n877 GNDA.n875 3.5845
R4219 GNDA.n1514 GNDA.n1513 3.5845
R4220 GNDA.n1509 GNDA.n878 3.5845
R4221 GNDA.n1508 GNDA.n882 3.5845
R4222 GNDA.n2055 GNDA.n2054 3.5845
R4223 GNDA.n2050 GNDA.n246 3.5845
R4224 GNDA.n2049 GNDA.n2025 3.5845
R4225 GNDA.n2046 GNDA.n2045 3.5845
R4226 GNDA.n2028 GNDA.n2026 3.5845
R4227 GNDA.n2040 GNDA.n2033 3.5845
R4228 GNDA.n2039 GNDA.n2034 3.5845
R4229 GNDA.n2036 GNDA.n2035 3.5845
R4230 GNDA.n2062 GNDA.n223 3.5845
R4231 GNDA.n2379 GNDA.t309 3.42907
R4232 GNDA.n2379 GNDA.t98 3.42907
R4233 GNDA.n2423 GNDA.t100 3.42907
R4234 GNDA.n2423 GNDA.t344 3.42907
R4235 GNDA.n2425 GNDA.t79 3.42907
R4236 GNDA.n2425 GNDA.t246 3.42907
R4237 GNDA.n2374 GNDA.t86 3.42907
R4238 GNDA.n2374 GNDA.t53 3.42907
R4239 GNDA.n834 GNDA.n519 3.3797
R4240 GNDA.n1589 GNDA.n1588 3.3797
R4241 GNDA.n2116 GNDA.n2115 3.3797
R4242 GNDA.n1201 GNDA.n1200 3.3797
R4243 GNDA.n991 GNDA.n990 3.3797
R4244 GNDA.n1847 GNDA.n1846 3.3797
R4245 GNDA.n592 GNDA.n412 3.3797
R4246 GNDA.n1439 GNDA.n1438 3.3797
R4247 GNDA.n2061 GNDA.n219 3.3797
R4248 GNDA.n1331 GNDA.n1330 3.2005
R4249 GNDA.n1748 GNDA.n346 3.2005
R4250 GNDA.t338 GNDA.n90 3.1344
R4251 GNDA.t312 GNDA.t187 3.1344
R4252 GNDA.n2162 GNDA.t345 3.1344
R4253 GNDA.n2182 GNDA.t56 3.1344
R4254 GNDA.t163 GNDA.t354 3.1344
R4255 GNDA.n2186 GNDA.t293 3.1344
R4256 GNDA.t96 GNDA.n2471 3.1344
R4257 GNDA.t84 GNDA.n2243 3.1344
R4258 GNDA.n772 GNDA.n771 2.8677
R4259 GNDA.n1679 GNDA.n438 2.8677
R4260 GNDA.n2147 GNDA.n2146 2.8677
R4261 GNDA.n1296 GNDA.n1295 2.8677
R4262 GNDA.n1083 GNDA.n961 2.8677
R4263 GNDA.n1939 GNDA.n290 2.8677
R4264 GNDA.n684 GNDA.n569 2.8677
R4265 GNDA.n1531 GNDA.n863 2.8677
R4266 GNDA.n2019 GNDA.n245 2.8677
R4267 GNDA.t258 GNDA.n2340 2.53799
R4268 GNDA.t250 GNDA.n2351 2.53799
R4269 GNDA.n2514 GNDA.n1 2.5005
R4270 GNDA.n1758 GNDA.n1757 2.4301
R4271 GNDA.n2218 GNDA.n2216 2.34425
R4272 GNDA.n2226 GNDA.n2224 2.34425
R4273 GNDA.n773 GNDA.n772 2.31161
R4274 GNDA.n1604 GNDA.n438 2.31161
R4275 GNDA.n2147 GNDA.n109 2.31161
R4276 GNDA.n1296 GNDA.n1176 2.31161
R4277 GNDA.n1006 GNDA.n961 2.31161
R4278 GNDA.n1862 GNDA.n290 2.31161
R4279 GNDA.n607 GNDA.n569 2.31161
R4280 GNDA.n1454 GNDA.n863 2.31161
R4281 GNDA.n2019 GNDA.n2018 2.31161
R4282 GNDA.n2424 GNDA.n2422 2.063
R4283 GNDA.n781 GNDA 1.95606
R4284 GNDA.n1612 GNDA 1.95606
R4285 GNDA GNDA.n133 1.95606
R4286 GNDA.n1224 GNDA 1.95606
R4287 GNDA.n1014 GNDA 1.95606
R4288 GNDA.n1870 GNDA 1.95606
R4289 GNDA.n615 GNDA 1.95606
R4290 GNDA.n1462 GNDA 1.95606
R4291 GNDA GNDA.n2011 1.95606
R4292 GNDA.n2393 GNDA.n2380 1.813
R4293 GNDA.n2422 GNDA.n2421 1.78175
R4294 GNDA.n2394 GNDA.n2393 1.78175
R4295 GNDA.n772 GNDA.n770 1.7413
R4296 GNDA.n1682 GNDA.n438 1.7413
R4297 GNDA.n2148 GNDA.n2147 1.7413
R4298 GNDA.n1297 GNDA.n1296 1.7413
R4299 GNDA.n1087 GNDA.n961 1.7413
R4300 GNDA.n290 GNDA.n288 1.7413
R4301 GNDA.n569 GNDA.n567 1.7413
R4302 GNDA.n863 GNDA.n860 1.7413
R4303 GNDA.n2020 GNDA.n2019 1.7413
R4304 GNDA.n1763 GNDA.n1762 1.73362
R4305 GNDA.n2500 GNDA.n3 1.6005
R4306 GNDA.n524 GNDA.n519 1.2293
R4307 GNDA.n1589 GNDA.n456 1.2293
R4308 GNDA.n2117 GNDA.n2116 1.2293
R4309 GNDA.n1201 GNDA.n1194 1.2293
R4310 GNDA.n991 GNDA.n982 1.2293
R4311 GNDA.n1847 GNDA.n309 1.2293
R4312 GNDA.n592 GNDA.n590 1.2293
R4313 GNDA.n1439 GNDA.n882 1.2293
R4314 GNDA.n2062 GNDA.n2061 1.2293
R4315 GNDA.n2398 GNDA.n2397 1.21925
R4316 GNDA.n731 GNDA.n557 1.1781
R4317 GNDA.n1683 GNDA.n437 1.1781
R4318 GNDA.n2149 GNDA.n108 1.1781
R4319 GNDA.n1174 GNDA.n1170 1.1781
R4320 GNDA.n1091 GNDA.n1088 1.1781
R4321 GNDA.n1945 GNDA.n1944 1.1781
R4322 GNDA.n566 GNDA.n353 1.1781
R4323 GNDA.n1689 GNDA.n416 1.1781
R4324 GNDA.n1969 GNDA.n1968 1.1781
R4325 GNDA.n1764 GNDA.n334 1.16414
R4326 GNDA.n771 GNDA.n365 1.0245
R4327 GNDA.n1732 GNDA.n1731 1.0245
R4328 GNDA.n1727 GNDA.n366 1.0245
R4329 GNDA.n1726 GNDA.n369 1.0245
R4330 GNDA.n531 GNDA.n527 1.0245
R4331 GNDA.n532 GNDA.n526 1.0245
R4332 GNDA.n538 GNDA.n536 1.0245
R4333 GNDA.n537 GNDA.n523 1.0245
R4334 GNDA.n828 GNDA.n827 1.0245
R4335 GNDA.n1679 GNDA.n1678 1.0245
R4336 GNDA.n441 GNDA.n439 1.0245
R4337 GNDA.n1673 GNDA.n445 1.0245
R4338 GNDA.n1672 GNDA.n446 1.0245
R4339 GNDA.n1669 GNDA.n1668 1.0245
R4340 GNDA.n449 GNDA.n447 1.0245
R4341 GNDA.n1663 GNDA.n453 1.0245
R4342 GNDA.n1662 GNDA.n454 1.0245
R4343 GNDA.n1659 GNDA.n1658 1.0245
R4344 GNDA.n2146 GNDA.n110 1.0245
R4345 GNDA.n2143 GNDA.n2142 1.0245
R4346 GNDA.n2138 GNDA.n111 1.0245
R4347 GNDA.n2137 GNDA.n2134 1.0245
R4348 GNDA.n2133 GNDA.n114 1.0245
R4349 GNDA.n2130 GNDA.n2129 1.0245
R4350 GNDA.n2125 GNDA.n115 1.0245
R4351 GNDA.n2124 GNDA.n2121 1.0245
R4352 GNDA.n2120 GNDA.n119 1.0245
R4353 GNDA.n1295 GNDA.n1177 1.0245
R4354 GNDA.n1292 GNDA.n1291 1.0245
R4355 GNDA.n1287 GNDA.n1179 1.0245
R4356 GNDA.n1286 GNDA.n1182 1.0245
R4357 GNDA.n1282 GNDA.n1281 1.0245
R4358 GNDA.n1187 GNDA.n1185 1.0245
R4359 GNDA.n1276 GNDA.n1189 1.0245
R4360 GNDA.n1275 GNDA.n1190 1.0245
R4361 GNDA.n1271 GNDA.n1270 1.0245
R4362 GNDA.n1083 GNDA.n1082 1.0245
R4363 GNDA.n966 GNDA.n964 1.0245
R4364 GNDA.n1077 GNDA.n968 1.0245
R4365 GNDA.n1076 GNDA.n969 1.0245
R4366 GNDA.n1072 GNDA.n1071 1.0245
R4367 GNDA.n975 GNDA.n973 1.0245
R4368 GNDA.n1066 GNDA.n977 1.0245
R4369 GNDA.n1065 GNDA.n978 1.0245
R4370 GNDA.n1061 GNDA.n1060 1.0245
R4371 GNDA.n1939 GNDA.n1938 1.0245
R4372 GNDA.n293 GNDA.n291 1.0245
R4373 GNDA.n1933 GNDA.n295 1.0245
R4374 GNDA.n1932 GNDA.n296 1.0245
R4375 GNDA.n1928 GNDA.n1927 1.0245
R4376 GNDA.n302 GNDA.n300 1.0245
R4377 GNDA.n1922 GNDA.n304 1.0245
R4378 GNDA.n1921 GNDA.n305 1.0245
R4379 GNDA.n1917 GNDA.n1916 1.0245
R4380 GNDA.n684 GNDA.n683 1.0245
R4381 GNDA.n572 GNDA.n570 1.0245
R4382 GNDA.n678 GNDA.n574 1.0245
R4383 GNDA.n677 GNDA.n575 1.0245
R4384 GNDA.n673 GNDA.n672 1.0245
R4385 GNDA.n581 GNDA.n579 1.0245
R4386 GNDA.n667 GNDA.n583 1.0245
R4387 GNDA.n666 GNDA.n584 1.0245
R4388 GNDA.n662 GNDA.n661 1.0245
R4389 GNDA.n1531 GNDA.n1530 1.0245
R4390 GNDA.n866 GNDA.n864 1.0245
R4391 GNDA.n1525 GNDA.n868 1.0245
R4392 GNDA.n1524 GNDA.n869 1.0245
R4393 GNDA.n1520 GNDA.n1519 1.0245
R4394 GNDA.n875 GNDA.n873 1.0245
R4395 GNDA.n1514 GNDA.n877 1.0245
R4396 GNDA.n1513 GNDA.n878 1.0245
R4397 GNDA.n1509 GNDA.n1508 1.0245
R4398 GNDA.n2055 GNDA.n245 1.0245
R4399 GNDA.n2054 GNDA.n246 1.0245
R4400 GNDA.n2050 GNDA.n2049 1.0245
R4401 GNDA.n2046 GNDA.n2025 1.0245
R4402 GNDA.n2045 GNDA.n2026 1.0245
R4403 GNDA.n2033 GNDA.n2028 1.0245
R4404 GNDA.n2040 GNDA.n2039 1.0245
R4405 GNDA.n2036 GNDA.n2034 1.0245
R4406 GNDA.n2035 GNDA.n223 1.0245
R4407 GNDA.n2506 GNDA.n2504 0.688
R4408 GNDA.n2508 GNDA.n2506 0.688
R4409 GNDA.n2510 GNDA.n2508 0.688
R4410 GNDA.n2512 GNDA.n2510 0.688
R4411 GNDA.t350 GNDA.n43 0.679512
R4412 GNDA.n2397 GNDA.n2396 0.6255
R4413 GNDA.n2216 GNDA.n2214 0.563
R4414 GNDA.n2220 GNDA.n2218 0.563
R4415 GNDA.n2222 GNDA.n2220 0.563
R4416 GNDA.n2224 GNDA.n2222 0.563
R4417 GNDA.n2228 GNDA.n2226 0.563
R4418 GNDA.n2230 GNDA.n2228 0.563
R4419 GNDA.n2293 GNDA.n2292 0.563
R4420 GNDA.n2293 GNDA.n2289 0.563
R4421 GNDA.n2385 GNDA.n2383 0.563
R4422 GNDA.n2387 GNDA.n2385 0.563
R4423 GNDA.n2389 GNDA.n2387 0.563
R4424 GNDA.n2391 GNDA.n2389 0.563
R4425 GNDA.n2420 GNDA.n2418 0.563
R4426 GNDA.n2418 GNDA.n2416 0.563
R4427 GNDA.n2416 GNDA.n2414 0.563
R4428 GNDA.n2414 GNDA.n2412 0.563
R4429 GNDA.n2412 GNDA.n2410 0.563
R4430 GNDA.n2410 GNDA.n2408 0.563
R4431 GNDA.n2408 GNDA.n2406 0.563
R4432 GNDA.n2406 GNDA.n2404 0.563
R4433 GNDA.n2404 GNDA.n2402 0.563
R4434 GNDA.n2402 GNDA.n2400 0.563
R4435 GNDA.n2352 GNDA.t307 0.507997
R4436 GNDA.n2426 GNDA.n2424 0.5005
R4437 GNDA.n2380 GNDA.n2378 0.5005
R4438 GNDA.n340 GNDA.n339 0.41175
R4439 GNDA.n341 GNDA.n340 0.311875
R4440 GNDA.n2421 GNDA.n2420 0.28175
R4441 GNDA.n2233 GNDA.n2232 0.276625
R4442 GNDA.n2211 GNDA.n60 0.276625
R4443 GNDA.n2296 GNDA.n2295 0.2505
R4444 GNDA.n2400 GNDA.n2398 0.2505
R4445 GNDA.n2396 GNDA.n2394 0.2505
R4446 GNDA.n2232 GNDA.n2231 0.22375
R4447 GNDA GNDA.n727 0.129793
R4448 GNDA GNDA.n1166 0.129793
R4449 GNDA.n1344 GNDA 0.129793
R4450 GNDA.n2231 GNDA.n2211 0.100375
R4451 GNDA.n1762 GNDA.n341 0.076875
R4452 GNDA.n857 GNDA.n413 0.0479074
R4453 GNDA.n845 GNDA 0.0479074
R4454 GNDA.n502 GNDA.n470 0.0479074
R4455 GNDA.n1576 GNDA 0.0479074
R4456 GNDA.n1786 GNDA.n1785 0.0479074
R4457 GNDA GNDA.n279 0.0479074
R4458 GNDA.n926 GNDA.n895 0.0479074
R4459 GNDA.n1426 GNDA 0.0479074
R4460 GNDA.n1710 GNDA.n1709 0.0479074
R4461 GNDA GNDA.n951 0.0479074
R4462 GNDA.n1385 GNDA.n1093 0.0479074
R4463 GNDA.n1108 GNDA 0.0479074
R4464 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 114.719
R4465 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R4466 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R4467 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 114.156
R4468 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R4469 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R4470 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R4471 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R4472 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R4473 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R4474 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R4475 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R4476 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R4477 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R4478 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R4479 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R4480 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R4481 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R4482 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R4483 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R4484 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R4485 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R4486 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R4487 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R4488 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R4489 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R4490 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R4491 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R4492 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R4493 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R4494 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R4495 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R4496 two_stage_opamp_dummy_magic_0.VD2.t14 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R4497 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R4498 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R4499 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R4500 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R4501 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R4502 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R4503 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R4504 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n8 0.563
R4505 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n5 145.989
R4506 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n6 145.989
R4507 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n11 145.427
R4508 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n9 145.427
R4509 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n7 145.427
R4510 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n14 140.927
R4511 two_stage_opamp_dummy_magic_0.VOUT-.t16 two_stage_opamp_dummy_magic_0.VOUT-.n100 113.192
R4512 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n0 95.7303
R4513 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n3 94.6053
R4514 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n1 94.6053
R4515 two_stage_opamp_dummy_magic_0.VOUT-.n99 two_stage_opamp_dummy_magic_0.VOUT-.n15 20.5943
R4516 two_stage_opamp_dummy_magic_0.VOUT-.n99 two_stage_opamp_dummy_magic_0.VOUT-.n98 11.7059
R4517 two_stage_opamp_dummy_magic_0.VOUT-.n100 two_stage_opamp_dummy_magic_0.VOUT-.n99 10.6567
R4518 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t7 6.56717
R4519 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t6 6.56717
R4520 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t17 6.56717
R4521 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t3 6.56717
R4522 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t5 6.56717
R4523 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t4 6.56717
R4524 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t13 6.56717
R4525 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t0 6.56717
R4526 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t2 6.56717
R4527 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t15 6.56717
R4528 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t14 6.56717
R4529 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t1 6.56717
R4530 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.t83 4.8295
R4531 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.t90 4.8295
R4532 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t128 4.8295
R4533 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t26 4.8295
R4534 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t74 4.8295
R4535 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t39 4.8295
R4536 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t34 4.8295
R4537 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t136 4.8295
R4538 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t68 4.8295
R4539 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t36 4.8295
R4540 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t94 4.8295
R4541 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t64 4.8295
R4542 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t54 4.8295
R4543 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t29 4.8295
R4544 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t89 4.8295
R4545 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t57 4.8295
R4546 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t48 4.8295
R4547 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.t20 4.8295
R4548 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t148 4.8295
R4549 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.t121 4.8295
R4550 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t43 4.8295
R4551 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.t152 4.8295
R4552 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t107 4.8295
R4553 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t28 4.8295
R4554 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t24 4.8295
R4555 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t129 4.8295
R4556 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t59 4.8295
R4557 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t32 4.8295
R4558 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t99 4.8295
R4559 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t69 4.8295
R4560 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t67 4.8295
R4561 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t35 4.8295
R4562 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t104 4.8295
R4563 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.t76 4.8295
R4564 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.t115 4.8295
R4565 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t132 4.806
R4566 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t114 4.806
R4567 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t146 4.806
R4568 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t45 4.806
R4569 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t85 4.806
R4570 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t63 4.806
R4571 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t101 4.806
R4572 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t134 4.806
R4573 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t119 4.806
R4574 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t155 4.806
R4575 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t47 4.806
R4576 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t91 4.806
R4577 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t41 4.806
R4578 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t130 4.806
R4579 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t82 4.806
R4580 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t124 4.806
R4581 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t72 4.806
R4582 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t23 4.806
R4583 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t62 4.806
R4584 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t150 4.806
R4585 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t95 4.5005
R4586 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.t56 4.5005
R4587 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.t131 4.5005
R4588 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t103 4.5005
R4589 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t71 4.5005
R4590 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t31 4.5005
R4591 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t138 4.5005
R4592 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t106 4.5005
R4593 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t60 4.5005
R4594 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t40 4.5005
R4595 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t143 4.5005
R4596 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t113 4.5005
R4597 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t21 4.5005
R4598 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t125 4.5005
R4599 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t118 4.5005
R4600 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t80 4.5005
R4601 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t96 4.5005
R4602 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t61 4.5005
R4603 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t27 4.5005
R4604 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t44 4.5005
R4605 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t144 4.5005
R4606 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t111 4.5005
R4607 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t75 4.5005
R4608 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t92 4.5005
R4609 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t55 4.5005
R4610 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t19 4.5005
R4611 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t51 4.5005
R4612 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t156 4.5005
R4613 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t120 4.5005
R4614 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t87 4.5005
R4615 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t49 4.5005
R4616 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t151 4.5005
R4617 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t42 4.5005
R4618 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t145 4.5005
R4619 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t117 4.5005
R4620 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t141 4.5005
R4621 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t110 4.5005
R4622 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t79 4.5005
R4623 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t38 4.5005
R4624 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t139 4.5005
R4625 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t108 4.5005
R4626 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t135 4.5005
R4627 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t102 4.5005
R4628 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.t70 4.5005
R4629 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t98 4.5005
R4630 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t66 4.5005
R4631 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.t33 4.5005
R4632 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t133 4.5005
R4633 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.t97 4.5005
R4634 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.t65 4.5005
R4635 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.t100 4.5005
R4636 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t149 4.5005
R4637 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t86 4.5005
R4638 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t50 4.5005
R4639 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t137 4.5005
R4640 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t105 4.5005
R4641 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t73 4.5005
R4642 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t25 4.5005
R4643 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t127 4.5005
R4644 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t88 4.5005
R4645 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t53 4.5005
R4646 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t140 4.5005
R4647 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.t109 4.5005
R4648 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t78 4.5005
R4649 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t112 4.5005
R4650 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.t77 4.5005
R4651 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t37 4.5005
R4652 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t147 4.5005
R4653 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.t116 4.5005
R4654 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t81 4.5005
R4655 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t46 4.5005
R4656 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.t153 4.5005
R4657 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t122 4.5005
R4658 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t154 4.5005
R4659 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.t123 4.5005
R4660 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t84 4.5005
R4661 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t52 4.5005
R4662 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t22 4.5005
R4663 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.t126 4.5005
R4664 two_stage_opamp_dummy_magic_0.VOUT-.n98 two_stage_opamp_dummy_magic_0.VOUT-.t142 4.5005
R4665 two_stage_opamp_dummy_magic_0.VOUT-.n97 two_stage_opamp_dummy_magic_0.VOUT-.t93 4.5005
R4666 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.t58 4.5005
R4667 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.t30 4.5005
R4668 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n13 4.5005
R4669 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t12 3.42907
R4670 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t10 3.42907
R4671 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t18 3.42907
R4672 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t8 3.42907
R4673 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t11 3.42907
R4674 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t9 3.42907
R4675 two_stage_opamp_dummy_magic_0.VOUT-.n100 two_stage_opamp_dummy_magic_0.VOUT-.n4 2.03175
R4676 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n2 1.1255
R4677 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n8 0.563
R4678 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n10 0.563
R4679 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n12 0.563
R4680 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.n45 0.3295
R4681 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.n48 0.3295
R4682 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.n47 0.3295
R4683 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.n51 0.3295
R4684 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.n50 0.3295
R4685 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.n54 0.3295
R4686 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.n53 0.3295
R4687 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n57 0.3295
R4688 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n56 0.3295
R4689 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.n59 0.3295
R4690 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n60 0.3295
R4691 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.n61 0.3295
R4692 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n62 0.3295
R4693 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.n63 0.3295
R4694 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.n64 0.3295
R4695 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n65 0.3295
R4696 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.n66 0.3295
R4697 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.n67 0.3295
R4698 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n68 0.3295
R4699 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n69 0.3295
R4700 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n71 0.3295
R4701 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n72 0.3295
R4702 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n74 0.3295
R4703 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n75 0.3295
R4704 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n77 0.3295
R4705 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n78 0.3295
R4706 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n80 0.3295
R4707 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n81 0.3295
R4708 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n83 0.3295
R4709 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n84 0.3295
R4710 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.n86 0.3295
R4711 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.n87 0.3295
R4712 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.n89 0.3295
R4713 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.n90 0.3295
R4714 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.n92 0.3295
R4715 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.n93 0.3295
R4716 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.n16 0.3295
R4717 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.n18 0.3295
R4718 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.n19 0.3295
R4719 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.n20 0.3295
R4720 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.n21 0.3295
R4721 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.n22 0.3295
R4722 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n23 0.3295
R4723 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.n24 0.3295
R4724 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.n25 0.3295
R4725 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n26 0.3295
R4726 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n27 0.3295
R4727 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n28 0.3295
R4728 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n30 0.3295
R4729 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n31 0.3295
R4730 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n33 0.3295
R4731 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n34 0.3295
R4732 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n36 0.3295
R4733 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n37 0.3295
R4734 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n39 0.3295
R4735 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n40 0.3295
R4736 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.n42 0.3295
R4737 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.n43 0.3295
R4738 two_stage_opamp_dummy_magic_0.VOUT-.n98 two_stage_opamp_dummy_magic_0.VOUT-.n97 0.3295
R4739 two_stage_opamp_dummy_magic_0.VOUT-.n97 two_stage_opamp_dummy_magic_0.VOUT-.n96 0.3295
R4740 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n95 0.3295
R4741 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n49 0.306
R4742 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.n52 0.306
R4743 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.n55 0.306
R4744 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n58 0.306
R4745 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n46 0.2825
R4746 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n70 0.2825
R4747 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n73 0.2825
R4748 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n76 0.2825
R4749 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n79 0.2825
R4750 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n82 0.2825
R4751 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.n85 0.2825
R4752 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.n88 0.2825
R4753 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.n91 0.2825
R4754 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n17 0.2825
R4755 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n29 0.2825
R4756 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n32 0.2825
R4757 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n35 0.2825
R4758 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n38 0.2825
R4759 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.n41 0.2825
R4760 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n44 0.2825
R4761 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n94 0.2825
R4762 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R4763 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1603
R4764 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1603
R4765 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R4766 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R4767 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R4768 two_stage_opamp_dummy_magic_0.cap_res_X.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R4769 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R4770 two_stage_opamp_dummy_magic_0.cap_res_X.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1603
R4771 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R4772 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.1603
R4773 two_stage_opamp_dummy_magic_0.cap_res_X.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1603
R4774 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1603
R4775 two_stage_opamp_dummy_magic_0.cap_res_X.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R4776 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R4777 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R4778 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R4779 two_stage_opamp_dummy_magic_0.cap_res_X.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R4780 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R4781 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R4782 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R4783 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R4784 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R4785 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R4786 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R4787 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R4788 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R4789 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R4790 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R4791 two_stage_opamp_dummy_magic_0.cap_res_X.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R4792 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R4793 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R4794 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R4795 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R4796 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R4797 two_stage_opamp_dummy_magic_0.cap_res_X.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R4798 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R4799 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1603
R4800 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R4801 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R4802 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R4803 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1603
R4804 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R4805 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.1603
R4806 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R4807 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1603
R4808 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R4809 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R4810 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1603
R4811 two_stage_opamp_dummy_magic_0.cap_res_X.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R4812 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R4813 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R4814 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R4815 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R4816 two_stage_opamp_dummy_magic_0.cap_res_X.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R4817 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R4818 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R4819 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R4820 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.1603
R4821 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.159278
R4822 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R4823 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R4824 two_stage_opamp_dummy_magic_0.cap_res_X.t41 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R4825 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R4826 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R4827 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R4828 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R4829 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R4830 two_stage_opamp_dummy_magic_0.cap_res_X.t91 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R4831 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R4832 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R4833 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R4834 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R4835 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R4836 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R4837 two_stage_opamp_dummy_magic_0.cap_res_X.t102 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R4838 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R4839 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.159278
R4840 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R4841 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R4842 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.159278
R4843 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R4844 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.159278
R4845 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.159278
R4846 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.159278
R4847 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.159278
R4848 two_stage_opamp_dummy_magic_0.cap_res_X.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.137822
R4849 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R4850 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.1368
R4851 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.1368
R4852 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R4853 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1368
R4854 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1368
R4855 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1368
R4856 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R4857 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R4858 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1368
R4859 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R4860 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1368
R4861 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R4862 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R4863 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1368
R4864 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1368
R4865 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R4866 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R4867 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.1368
R4868 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R4869 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R4870 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1368
R4871 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R4872 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1368
R4873 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1368
R4874 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R4875 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R4876 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1368
R4877 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1368
R4878 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R4879 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R4880 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.118
R4881 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.114322
R4882 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R4883 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R4884 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R4885 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R4886 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R4887 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R4888 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R4889 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R4890 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R4891 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R4892 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R4893 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R4894 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R4895 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R4896 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R4897 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R4898 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R4899 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R4900 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R4901 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R4902 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R4903 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.00152174
R4904 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.00152174
R4905 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R4906 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R4907 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.00152174
R4908 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.00152174
R4909 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R4910 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.00152174
R4911 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.00152174
R4912 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R4913 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.00152174
R4914 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R4915 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.00152174
R4916 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R4917 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R4918 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R4919 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.00152174
R4920 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.00152174
R4921 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R4922 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R4923 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R4924 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.00152174
R4925 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R4926 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.00152174
R4927 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.00152174
R4928 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R4929 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R4930 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.00152174
R4931 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.00152174
R4932 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.00152174
R4933 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R4934 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R4935 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.00152174
R4936 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R4937 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t23 369.534
R4938 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t16 369.534
R4939 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t24 369.534
R4940 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t27 369.534
R4941 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R4942 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t29 369.534
R4943 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R4944 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R4945 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R4946 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R4947 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t20 238.322
R4948 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t11 238.322
R4949 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t0 194.895
R4950 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t17 192.8
R4951 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t28 192.8
R4952 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t14 192.8
R4953 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R4954 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t13 192.8
R4955 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t19 192.8
R4956 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t10 192.8
R4957 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t26 192.8
R4958 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t15 192.8
R4959 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t25 192.8
R4960 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t12 192.8
R4961 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t18 192.8
R4962 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R4963 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R4964 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R4965 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R4966 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R4967 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R4968 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R4969 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R4970 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R4971 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R4972 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t1 100.635
R4973 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R4974 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R4975 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R4976 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R4977 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R4978 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R4979 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t6 39.4005
R4980 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R4981 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t4 39.4005
R4982 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t8 39.4005
R4983 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t3 39.4005
R4984 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t7 39.4005
R4985 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t2 39.4005
R4986 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t5 39.4005
R4987 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R4988 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R4989 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R4990 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R4991 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R4992 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R4993 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R4994 VDDA.n121 VDDA.n89 6600
R4995 VDDA.n123 VDDA.n89 6600
R4996 VDDA.n121 VDDA.n88 6570
R4997 VDDA.n123 VDDA.n88 6570
R4998 VDDA.n78 VDDA.n11 4710
R4999 VDDA.n78 VDDA.n12 4710
R5000 VDDA.n76 VDDA.n12 4710
R5001 VDDA.n76 VDDA.n11 4710
R5002 VDDA.n30 VDDA.n23 4710
R5003 VDDA.n32 VDDA.n23 4710
R5004 VDDA.n30 VDDA.n29 4710
R5005 VDDA.n32 VDDA.n29 4710
R5006 VDDA.n356 VDDA.n352 4605
R5007 VDDA.n356 VDDA.n353 4605
R5008 VDDA.n257 VDDA.n243 4605
R5009 VDDA.n259 VDDA.n243 4605
R5010 VDDA.n421 VDDA.n397 4590
R5011 VDDA.n423 VDDA.n397 4590
R5012 VDDA.n423 VDDA.n398 4590
R5013 VDDA.n421 VDDA.n398 4590
R5014 VDDA.n358 VDDA.n352 4575
R5015 VDDA.n358 VDDA.n353 4575
R5016 VDDA.n257 VDDA.n244 4575
R5017 VDDA.n259 VDDA.n244 4575
R5018 VDDA.n316 VDDA.n309 4020
R5019 VDDA.n318 VDDA.n309 4020
R5020 VDDA.n316 VDDA.n315 4020
R5021 VDDA.n318 VDDA.n315 4020
R5022 VDDA.n292 VDDA.n285 4020
R5023 VDDA.n294 VDDA.n285 4020
R5024 VDDA.n292 VDDA.n291 4020
R5025 VDDA.n294 VDDA.n291 4020
R5026 VDDA.n187 VDDA.n155 3420
R5027 VDDA.n187 VDDA.n156 3420
R5028 VDDA.n336 VDDA.n329 3390
R5029 VDDA.n338 VDDA.n329 3390
R5030 VDDA.n336 VDDA.n335 3390
R5031 VDDA.n338 VDDA.n335 3390
R5032 VDDA.n236 VDDA.n229 3390
R5033 VDDA.n238 VDDA.n229 3390
R5034 VDDA.n236 VDDA.n235 3390
R5035 VDDA.n238 VDDA.n235 3390
R5036 VDDA.n378 VDDA.n372 2940
R5037 VDDA.n380 VDDA.n372 2940
R5038 VDDA.n380 VDDA.n377 2940
R5039 VDDA.n378 VDDA.n377 2940
R5040 VDDA.n386 VDDA.n367 2940
R5041 VDDA.n388 VDDA.n367 2940
R5042 VDDA.n388 VDDA.n385 2940
R5043 VDDA.n386 VDDA.n385 2940
R5044 VDDA.n189 VDDA.n155 2760
R5045 VDDA.n189 VDDA.n156 2760
R5046 VDDA.n450 VDDA.n439 2415
R5047 VDDA.n450 VDDA.n440 2370
R5048 VDDA.n447 VDDA.n440 2280
R5049 VDDA.n447 VDDA.n439 2235
R5050 VDDA.n203 VDDA.n150 2145
R5051 VDDA.n200 VDDA.n149 2100
R5052 VDDA.n203 VDDA.n149 2100
R5053 VDDA.n168 VDDA.n161 2100
R5054 VDDA.n170 VDDA.n161 2100
R5055 VDDA.n168 VDDA.n162 2100
R5056 VDDA.n170 VDDA.n162 2100
R5057 VDDA.n200 VDDA.n150 2055
R5058 VDDA.n135 VDDA.n130 1770
R5059 VDDA.n137 VDDA.n130 1770
R5060 VDDA.n135 VDDA.n133 1770
R5061 VDDA.n137 VDDA.n133 1770
R5062 VDDA.n97 VDDA.n92 1770
R5063 VDDA.n99 VDDA.n92 1770
R5064 VDDA.n97 VDDA.n95 1770
R5065 VDDA.n99 VDDA.n95 1770
R5066 VDDA.n462 VDDA.n435 1575
R5067 VDDA.n461 VDDA.n435 1575
R5068 VDDA.n461 VDDA.n434 1545
R5069 VDDA.n462 VDDA.n434 1545
R5070 VDDA.n350 VDDA.t48 1216.42
R5071 VDDA.n361 VDDA.t30 1216.42
R5072 VDDA.n254 VDDA.t42 1216.42
R5073 VDDA.n262 VDDA.t66 1216.42
R5074 VDDA.n124 VDDA.n87 704
R5075 VDDA.n120 VDDA.n87 704
R5076 VDDA.n374 VDDA.t29 689.4
R5077 VDDA.n373 VDDA.t41 689.4
R5078 VDDA.n369 VDDA.t114 689.4
R5079 VDDA.n368 VDDA.t11 689.4
R5080 VDDA.n417 VDDA.t93 663.801
R5081 VDDA.n427 VDDA.t90 663.801
R5082 VDDA.n312 VDDA.t100 660.109
R5083 VDDA.n310 VDDA.t18 660.109
R5084 VDDA.n288 VDDA.t3 660.109
R5085 VDDA.n286 VDDA.t76 660.109
R5086 VDDA.n457 VDDA.t38 647.54
R5087 VDDA.n466 VDDA.t72 647.54
R5088 VDDA.n431 VDDA.n430 633.361
R5089 VDDA.n394 VDDA.n393 626.534
R5090 VDDA.n400 VDDA.n399 626.534
R5091 VDDA.n402 VDDA.n401 626.534
R5092 VDDA.n404 VDDA.n403 626.534
R5093 VDDA.n406 VDDA.n405 626.534
R5094 VDDA.n408 VDDA.n407 626.534
R5095 VDDA.n410 VDDA.n409 626.534
R5096 VDDA.n412 VDDA.n411 626.534
R5097 VDDA.n414 VDDA.n413 626.534
R5098 VDDA.n416 VDDA.n415 626.534
R5099 VDDA.n444 VDDA.t6 623.958
R5100 VDDA.n453 VDDA.t21 623.958
R5101 VDDA.t6 VDDA.n443 615.926
R5102 VDDA.n332 VDDA.t33 573.75
R5103 VDDA.n330 VDDA.t57 573.75
R5104 VDDA.n232 VDDA.t54 573.75
R5105 VDDA.n230 VDDA.t73 573.75
R5106 VDDA.n119 VDDA.n86 518.4
R5107 VDDA.n125 VDDA.n86 518.4
R5108 VDDA.n34 VDDA.n33 496
R5109 VDDA.n34 VDDA.n22 496
R5110 VDDA.n355 VDDA.n327 491.2
R5111 VDDA.n355 VDDA.n354 491.2
R5112 VDDA.n260 VDDA.n242 491.2
R5113 VDDA.n256 VDDA.n242 491.2
R5114 VDDA.n420 VDDA.n396 489.601
R5115 VDDA.n424 VDDA.n396 489.601
R5116 VDDA.n320 VDDA.n319 428.8
R5117 VDDA.n320 VDDA.n308 428.8
R5118 VDDA.n296 VDDA.n295 428.8
R5119 VDDA.n296 VDDA.n284 428.8
R5120 VDDA.n128 VDDA.t97 419.108
R5121 VDDA.n131 VDDA.t109 419.108
R5122 VDDA.n90 VDDA.t106 413.084
R5123 VDDA.n93 VDDA.t24 413.084
R5124 VDDA.n197 VDDA.t15 409.067
R5125 VDDA.n206 VDDA.t94 409.067
R5126 VDDA.n184 VDDA.t82 409.067
R5127 VDDA.n192 VDDA.t63 409.067
R5128 VDDA.n165 VDDA.t79 409.067
R5129 VDDA.n173 VDDA.t103 390.322
R5130 VDDA.t92 VDDA.n421 389.375
R5131 VDDA.n423 VDDA.t89 389.375
R5132 VDDA.t113 VDDA.n385 389.375
R5133 VDDA.t10 VDDA.n367 389.375
R5134 VDDA.n128 VDDA.t99 389.185
R5135 VDDA.n131 VDDA.t111 389.185
R5136 VDDA.n419 VDDA.n395 387.2
R5137 VDDA.n425 VDDA.n395 387.2
R5138 VDDA.n192 VDDA.t65 387.051
R5139 VDDA.n184 VDDA.t84 387.051
R5140 VDDA.n90 VDDA.t108 384.918
R5141 VDDA.n93 VDDA.t26 384.918
R5142 VDDA.n72 VDDA.t117 384.918
R5143 VDDA.n9 VDDA.t87 384.918
R5144 VDDA.n26 VDDA.t53 384.918
R5145 VDDA.n24 VDDA.t14 384.918
R5146 VDDA.t28 VDDA.n377 384.168
R5147 VDDA.t40 VDDA.n372 384.168
R5148 VDDA.n74 VDDA.n73 384
R5149 VDDA.n73 VDDA.n10 384
R5150 VDDA.n28 VDDA.n27 384
R5151 VDDA.n28 VDDA.n25 384
R5152 VDDA.n173 VDDA.t105 370.728
R5153 VDDA.n165 VDDA.t81 370.728
R5154 VDDA.n206 VDDA.t96 370.3
R5155 VDDA.n197 VDDA.t17 370.3
R5156 VDDA.n186 VDDA.n154 364.8
R5157 VDDA.n118 VDDA.t60 360.868
R5158 VDDA.n126 VDDA.t45 360.868
R5159 VDDA.n72 VDDA.t115 358.858
R5160 VDDA.n9 VDDA.t85 358.858
R5161 VDDA.n26 VDDA.t51 358.858
R5162 VDDA.n24 VDDA.t12 358.858
R5163 VDDA.n340 VDDA.n339 355.2
R5164 VDDA.n340 VDDA.n328 355.2
R5165 VDDA.n240 VDDA.n239 355.2
R5166 VDDA.n240 VDDA.n228 355.2
R5167 VDDA.t116 VDDA.n76 351.591
R5168 VDDA.n78 VDDA.t86 351.591
R5169 VDDA.t52 VDDA.n30 351.591
R5170 VDDA.n32 VDDA.t13 351.591
R5171 VDDA.t37 VDDA.n461 346.668
R5172 VDDA.n462 VDDA.t70 346.668
R5173 VDDA.n158 VDDA.n157 345.127
R5174 VDDA.n164 VDDA.n163 345.127
R5175 VDDA.n146 VDDA.n145 344.7
R5176 VDDA.n195 VDDA.n194 344.7
R5177 VDDA.t16 VDDA.n200 344.394
R5178 VDDA.n203 VDDA.t95 344.394
R5179 VDDA.t98 VDDA.n135 344.394
R5180 VDDA.n137 VDDA.t110 344.394
R5181 VDDA.t107 VDDA.n97 344.394
R5182 VDDA.n99 VDDA.t25 344.394
R5183 VDDA.n17 VDDA.n15 342.301
R5184 VDDA.n45 VDDA.n44 341.676
R5185 VDDA.n43 VDDA.n42 341.676
R5186 VDDA.n41 VDDA.n40 341.676
R5187 VDDA.n39 VDDA.n38 341.676
R5188 VDDA.n21 VDDA.n20 341.676
R5189 VDDA.n19 VDDA.n18 341.676
R5190 VDDA.n17 VDDA.n16 341.676
R5191 VDDA.t83 VDDA.n187 340.635
R5192 VDDA.n189 VDDA.t64 340.635
R5193 VDDA.t80 VDDA.n168 340.635
R5194 VDDA.n170 VDDA.t104 340.635
R5195 VDDA.n152 VDDA.n151 339.272
R5196 VDDA.n176 VDDA.n175 339.272
R5197 VDDA.n178 VDDA.n177 339.272
R5198 VDDA.n180 VDDA.n179 339.272
R5199 VDDA.n182 VDDA.n181 339.272
R5200 VDDA.n81 VDDA.n5 337.176
R5201 VDDA.n7 VDDA.n6 337.176
R5202 VDDA.n53 VDDA.n52 337.176
R5203 VDDA.n57 VDDA.n56 337.176
R5204 VDDA.n49 VDDA.n48 337.176
R5205 VDDA.n61 VDDA.n60 337.176
R5206 VDDA.n64 VDDA.n47 337.176
R5207 VDDA.n67 VDDA.n66 337.176
R5208 VDDA.n70 VDDA.n14 337.176
R5209 VDDA.n36 VDDA.n35 337.176
R5210 VDDA.n142 VDDA.n141 335.022
R5211 VDDA.n418 VDDA.t91 332.75
R5212 VDDA.n426 VDDA.t88 332.75
R5213 VDDA.n374 VDDA.t27 332.75
R5214 VDDA.n373 VDDA.t39 332.75
R5215 VDDA.n369 VDDA.t112 332.75
R5216 VDDA.n368 VDDA.t9 332.75
R5217 VDDA.n458 VDDA.t36 314.274
R5218 VDDA.n465 VDDA.t69 314.274
R5219 VDDA.n376 VDDA.n371 313.601
R5220 VDDA.n383 VDDA.n371 307.2
R5221 VDDA.n391 VDDA.n366 307.2
R5222 VDDA.n384 VDDA.n366 307.2
R5223 VDDA.n190 VDDA.n154 294.401
R5224 VDDA.t34 VDDA.n336 285.815
R5225 VDDA.n338 VDDA.t58 285.815
R5226 VDDA.t55 VDDA.n236 285.815
R5227 VDDA.n238 VDDA.t74 285.815
R5228 VDDA.t61 VDDA.n121 278.95
R5229 VDDA.n123 VDDA.t46 278.95
R5230 VDDA.n332 VDDA.t35 277.916
R5231 VDDA.n330 VDDA.t59 277.916
R5232 VDDA.n232 VDDA.t56 277.916
R5233 VDDA.n230 VDDA.t75 277.916
R5234 VDDA.n360 VDDA.n327 276.8
R5235 VDDA.n354 VDDA.n351 276.8
R5236 VDDA.n261 VDDA.n260 276.8
R5237 VDDA.n256 VDDA.n255 276.8
R5238 VDDA.n126 VDDA.t47 270.705
R5239 VDDA.n118 VDDA.t62 270.705
R5240 VDDA.n451 VDDA.n438 257.601
R5241 VDDA.n185 VDDA.n153 246.4
R5242 VDDA.t101 VDDA.n316 239.915
R5243 VDDA.n318 VDDA.t19 239.915
R5244 VDDA.t4 VDDA.n292 239.915
R5245 VDDA.n294 VDDA.t77 239.915
R5246 VDDA.n446 VDDA.n438 238.4
R5247 VDDA.n314 VDDA.n313 230.4
R5248 VDDA.n314 VDDA.n311 230.4
R5249 VDDA.n290 VDDA.n289 230.4
R5250 VDDA.n290 VDDA.n287 230.4
R5251 VDDA.n204 VDDA.n148 228.8
R5252 VDDA.n171 VDDA.n160 224
R5253 VDDA.n167 VDDA.n160 224
R5254 VDDA.n199 VDDA.n148 219.201
R5255 VDDA.n381 VDDA.n375 211.201
R5256 VDDA.n382 VDDA.n381 211.201
R5257 VDDA.n390 VDDA.n389 211.201
R5258 VDDA.n334 VDDA.n333 211.201
R5259 VDDA.n334 VDDA.n331 211.201
R5260 VDDA.n234 VDDA.n233 211.201
R5261 VDDA.n234 VDDA.n231 211.201
R5262 VDDA.n360 VDDA.n359 204.8
R5263 VDDA.n359 VDDA.n351 204.8
R5264 VDDA.n255 VDDA.n241 204.8
R5265 VDDA.n261 VDDA.n241 204.8
R5266 VDDA.n389 VDDA.n370 202.971
R5267 VDDA.n319 VDDA.n311 198.4
R5268 VDDA.n313 VDDA.n308 198.4
R5269 VDDA.n295 VDDA.n287 198.4
R5270 VDDA.n289 VDDA.n284 198.4
R5271 VDDA.n446 VDDA.n445 192
R5272 VDDA.t329 VDDA.t37 190
R5273 VDDA.t70 VDDA.t329 190
R5274 VDDA.n452 VDDA.n451 188.8
R5275 VDDA.n138 VDDA.n132 188.8
R5276 VDDA.n134 VDDA.n132 188.8
R5277 VDDA.n100 VDDA.n94 188.8
R5278 VDDA.n96 VDDA.n94 188.8
R5279 VDDA.n80 VDDA.n79 188.8
R5280 VDDA.n75 VDDA.n71 188.8
R5281 VDDA.t219 VDDA.t92 186.607
R5282 VDDA.t351 VDDA.t219 186.607
R5283 VDDA.t191 VDDA.t351 186.607
R5284 VDDA.t357 VDDA.t191 186.607
R5285 VDDA.t264 VDDA.t357 186.607
R5286 VDDA.t347 VDDA.t264 186.607
R5287 VDDA.t166 VDDA.t347 186.607
R5288 VDDA.t363 VDDA.t166 186.607
R5289 VDDA.t276 VDDA.t363 186.607
R5290 VDDA.t217 VDDA.t276 186.607
R5291 VDDA.t365 VDDA.t355 186.607
R5292 VDDA.t359 VDDA.t365 186.607
R5293 VDDA.t262 VDDA.t359 186.607
R5294 VDDA.t353 VDDA.t262 186.607
R5295 VDDA.t164 VDDA.t353 186.607
R5296 VDDA.t349 VDDA.t164 186.607
R5297 VDDA.t318 VDDA.t349 186.607
R5298 VDDA.t193 VDDA.t318 186.607
R5299 VDDA.t361 VDDA.t193 186.607
R5300 VDDA.t89 VDDA.t361 186.607
R5301 VDDA.t227 VDDA.t113 186.607
R5302 VDDA.t433 VDDA.t227 186.607
R5303 VDDA.t436 VDDA.t433 186.607
R5304 VDDA.t229 VDDA.t436 186.607
R5305 VDDA.t215 VDDA.t229 186.607
R5306 VDDA.t186 VDDA.t372 186.607
R5307 VDDA.t372 VDDA.t190 186.607
R5308 VDDA.t190 VDDA.t258 186.607
R5309 VDDA.t258 VDDA.t337 186.607
R5310 VDDA.t337 VDDA.t10 186.607
R5311 VDDA.t216 VDDA.t28 183.333
R5312 VDDA.t373 VDDA.t216 183.333
R5313 VDDA.t371 VDDA.t373 183.333
R5314 VDDA.t259 VDDA.t371 183.333
R5315 VDDA.t228 VDDA.t259 183.333
R5316 VDDA.t305 VDDA.t2 183.333
R5317 VDDA.t2 VDDA.t155 183.333
R5318 VDDA.t155 VDDA.t189 183.333
R5319 VDDA.t189 VDDA.t340 183.333
R5320 VDDA.t340 VDDA.t40 183.333
R5321 VDDA.n125 VDDA.n124 182.4
R5322 VDDA.n120 VDDA.n119 182.4
R5323 VDDA.n349 VDDA.t50 178.124
R5324 VDDA.n362 VDDA.t32 178.124
R5325 VDDA.n253 VDDA.t44 178.124
R5326 VDDA.n263 VDDA.t68 178.124
R5327 VDDA.n191 VDDA.n153 176
R5328 VDDA.n441 VDDA.n436 174.393
R5329 VDDA.t441 VDDA.t116 172.727
R5330 VDDA.t134 VDDA.t441 172.727
R5331 VDDA.t343 VDDA.t134 172.727
R5332 VDDA.t120 VDDA.t343 172.727
R5333 VDDA.t422 VDDA.t120 172.727
R5334 VDDA.t254 VDDA.t422 172.727
R5335 VDDA.t439 VDDA.t254 172.727
R5336 VDDA.t132 VDDA.t439 172.727
R5337 VDDA.t341 VDDA.t132 172.727
R5338 VDDA.t236 VDDA.t118 172.727
R5339 VDDA.t252 VDDA.t236 172.727
R5340 VDDA.t437 VDDA.t252 172.727
R5341 VDDA.t345 VDDA.t437 172.727
R5342 VDDA.t338 VDDA.t345 172.727
R5343 VDDA.t234 VDDA.t338 172.727
R5344 VDDA.t242 VDDA.t234 172.727
R5345 VDDA.t250 VDDA.t242 172.727
R5346 VDDA.t86 VDDA.t250 172.727
R5347 VDDA.t268 VDDA.t52 172.727
R5348 VDDA.t312 VDDA.t268 172.727
R5349 VDDA.t314 VDDA.t312 172.727
R5350 VDDA.t448 VDDA.t314 172.727
R5351 VDDA.t296 VDDA.t448 172.727
R5352 VDDA.t205 VDDA.t296 172.727
R5353 VDDA.t270 VDDA.t205 172.727
R5354 VDDA.t199 VDDA.t270 172.727
R5355 VDDA.t260 VDDA.t199 172.727
R5356 VDDA.t431 VDDA.t290 172.727
R5357 VDDA.t238 VDDA.t431 172.727
R5358 VDDA.t203 VDDA.t238 172.727
R5359 VDDA.t461 VDDA.t203 172.727
R5360 VDDA.t429 VDDA.t461 172.727
R5361 VDDA.t279 VDDA.t429 172.727
R5362 VDDA.t248 VDDA.t279 172.727
R5363 VDDA.t272 VDDA.t248 172.727
R5364 VDDA.t13 VDDA.t272 172.727
R5365 VDDA.t7 VDDA.n447 172.554
R5366 VDDA.n450 VDDA.t22 172.554
R5367 VDDA.n85 VDDA.n84 168.435
R5368 VDDA.n104 VDDA.n103 168.435
R5369 VDDA.n106 VDDA.n105 168.435
R5370 VDDA.n108 VDDA.n107 168.435
R5371 VDDA.n110 VDDA.n109 168.435
R5372 VDDA.n112 VDDA.n111 168.435
R5373 VDDA.n114 VDDA.n113 168.435
R5374 VDDA.n116 VDDA.n115 168.435
R5375 VDDA.n460 VDDA.n433 164.8
R5376 VDDA.n463 VDDA.n433 164.8
R5377 VDDA.t31 VDDA.n352 161.817
R5378 VDDA.t49 VDDA.n353 161.817
R5379 VDDA.t43 VDDA.n257 161.817
R5380 VDDA.n259 VDDA.t67 161.817
R5381 VDDA.n306 VDDA.n304 160.428
R5382 VDDA.n303 VDDA.n301 160.428
R5383 VDDA.n282 VDDA.n280 160.428
R5384 VDDA.n279 VDDA.n277 160.428
R5385 VDDA.t195 VDDA.t61 159.814
R5386 VDDA.t294 VDDA.t195 159.814
R5387 VDDA.t244 VDDA.t294 159.814
R5388 VDDA.t450 VDDA.t244 159.814
R5389 VDDA.t208 VDDA.t450 159.814
R5390 VDDA.t240 VDDA.t208 159.814
R5391 VDDA.t181 VDDA.t240 159.814
R5392 VDDA.t307 VDDA.t181 159.814
R5393 VDDA.t178 VDDA.t141 159.814
R5394 VDDA.t221 VDDA.t178 159.814
R5395 VDDA.t224 VDDA.t221 159.814
R5396 VDDA.t443 VDDA.t224 159.814
R5397 VDDA.t197 VDDA.t443 159.814
R5398 VDDA.t299 VDDA.t197 159.814
R5399 VDDA.t292 VDDA.t299 159.814
R5400 VDDA.t46 VDDA.t292 159.814
R5401 VDDA.n306 VDDA.n305 159.803
R5402 VDDA.n303 VDDA.n302 159.803
R5403 VDDA.n282 VDDA.n281 159.803
R5404 VDDA.n279 VDDA.n278 159.803
R5405 VDDA.t404 VDDA.t16 158.333
R5406 VDDA.t380 VDDA.t404 158.333
R5407 VDDA.t390 VDDA.t402 158.333
R5408 VDDA.t95 VDDA.t390 158.333
R5409 VDDA.t414 VDDA.t98 158.333
R5410 VDDA.t110 VDDA.t396 158.333
R5411 VDDA.t282 VDDA.t107 158.333
R5412 VDDA.t25 VDDA.t281 158.333
R5413 VDDA.t382 VDDA.t83 155.97
R5414 VDDA.t386 VDDA.t382 155.97
R5415 VDDA.t406 VDDA.t386 155.97
R5416 VDDA.t384 VDDA.t406 155.97
R5417 VDDA.t416 VDDA.t384 155.97
R5418 VDDA.t398 VDDA.t416 155.97
R5419 VDDA.t392 VDDA.t410 155.97
R5420 VDDA.t408 VDDA.t392 155.97
R5421 VDDA.t388 VDDA.t408 155.97
R5422 VDDA.t64 VDDA.t388 155.97
R5423 VDDA.t378 VDDA.t80 155.97
R5424 VDDA.t400 VDDA.t378 155.97
R5425 VDDA.t394 VDDA.t412 155.97
R5426 VDDA.t104 VDDA.t394 155.97
R5427 VDDA.n312 VDDA.t102 155.125
R5428 VDDA.n310 VDDA.t20 155.125
R5429 VDDA.n288 VDDA.t5 155.125
R5430 VDDA.n286 VDDA.t78 155.125
R5431 VDDA.n349 VDDA.n348 151.882
R5432 VDDA.n253 VDDA.n252 151.882
R5433 VDDA.n363 VDDA.n362 151.321
R5434 VDDA.n264 VDDA.n263 151.321
R5435 VDDA.n339 VDDA.n331 150.4
R5436 VDDA.n333 VDDA.n328 150.4
R5437 VDDA.n239 VDDA.n231 150.4
R5438 VDDA.n233 VDDA.n228 150.4
R5439 VDDA.n322 VDDA.n321 146.002
R5440 VDDA.n298 VDDA.n297 146.002
R5441 VDDA.n326 VDDA.n325 145.429
R5442 VDDA.n342 VDDA.n341 145.429
R5443 VDDA.n344 VDDA.n343 145.429
R5444 VDDA.n346 VDDA.n345 145.429
R5445 VDDA.n348 VDDA.n347 145.429
R5446 VDDA.n227 VDDA.n226 145.429
R5447 VDDA.n246 VDDA.n245 145.429
R5448 VDDA.n248 VDDA.n247 145.429
R5449 VDDA.n250 VDDA.n249 145.429
R5450 VDDA.n252 VDDA.n251 145.429
R5451 VDDA.n362 VDDA.n361 135.387
R5452 VDDA.n350 VDDA.n349 135.387
R5453 VDDA.n263 VDDA.n262 135.387
R5454 VDDA.n254 VDDA.n253 135.387
R5455 VDDA.t169 VDDA.t34 121.513
R5456 VDDA.t177 VDDA.t169 121.513
R5457 VDDA.t202 VDDA.t177 121.513
R5458 VDDA.t424 VDDA.t202 121.513
R5459 VDDA.t170 VDDA.t424 121.513
R5460 VDDA.t316 VDDA.t156 121.513
R5461 VDDA.t283 VDDA.t316 121.513
R5462 VDDA.t168 VDDA.t283 121.513
R5463 VDDA.t266 VDDA.t168 121.513
R5464 VDDA.t58 VDDA.t266 121.513
R5465 VDDA.t146 VDDA.t55 121.513
R5466 VDDA.t466 VDDA.t146 121.513
R5467 VDDA.t324 VDDA.t466 121.513
R5468 VDDA.t367 VDDA.t324 121.513
R5469 VDDA.t210 VDDA.t367 121.513
R5470 VDDA.t327 VDDA.t368 121.513
R5471 VDDA.t144 VDDA.t327 121.513
R5472 VDDA.t326 VDDA.t144 121.513
R5473 VDDA.t145 VDDA.t326 121.513
R5474 VDDA.t74 VDDA.t145 121.513
R5475 VDDA.n205 VDDA.n204 118.4
R5476 VDDA.n199 VDDA.n198 118.4
R5477 VDDA.n191 VDDA.n190 118.4
R5478 VDDA.n186 VDDA.n185 118.4
R5479 VDDA.n172 VDDA.n171 118.4
R5480 VDDA.n167 VDDA.n166 118.4
R5481 VDDA.n139 VDDA.n138 118.4
R5482 VDDA.n134 VDDA.n129 118.4
R5483 VDDA.n101 VDDA.n100 118.4
R5484 VDDA.n96 VDDA.n91 118.4
R5485 VDDA.n79 VDDA.n10 118.4
R5486 VDDA.n75 VDDA.n74 118.4
R5487 VDDA.n33 VDDA.n25 118.4
R5488 VDDA.n27 VDDA.n22 118.4
R5489 VDDA.n460 VDDA.n459 110.4
R5490 VDDA.n464 VDDA.n463 110.4
R5491 VDDA.n198 VDDA.n147 105.6
R5492 VDDA.n205 VDDA.n147 105.6
R5493 VDDA.n166 VDDA.n159 105.6
R5494 VDDA.n172 VDDA.n159 105.6
R5495 VDDA.t22 VDDA.t331 102.704
R5496 VDDA.n420 VDDA.n419 102.4
R5497 VDDA.n425 VDDA.n424 102.4
R5498 VDDA.n376 VDDA.n375 102.4
R5499 VDDA.n455 VDDA.n454 101.267
R5500 VDDA.t147 VDDA.t101 98.2764
R5501 VDDA.t418 VDDA.t147 98.2764
R5502 VDDA.t420 VDDA.t418 98.2764
R5503 VDDA.t333 VDDA.t420 98.2764
R5504 VDDA.t130 VDDA.t333 98.2764
R5505 VDDA.t162 VDDA.t374 98.2764
R5506 VDDA.t171 VDDA.t162 98.2764
R5507 VDDA.t187 VDDA.t171 98.2764
R5508 VDDA.t446 VDDA.t187 98.2764
R5509 VDDA.t19 VDDA.t446 98.2764
R5510 VDDA.t369 VDDA.t4 98.2764
R5511 VDDA.t434 VDDA.t369 98.2764
R5512 VDDA.t153 VDDA.t434 98.2764
R5513 VDDA.t464 VDDA.t153 98.2764
R5514 VDDA.t213 VDDA.t464 98.2764
R5515 VDDA.t335 VDDA.t184 98.2764
R5516 VDDA.t376 VDDA.t335 98.2764
R5517 VDDA.t149 VDDA.t376 98.2764
R5518 VDDA.t151 VDDA.t149 98.2764
R5519 VDDA.t77 VDDA.t151 98.2764
R5520 VDDA.n267 VDDA.n265 97.4034
R5521 VDDA.n217 VDDA.n215 97.4034
R5522 VDDA.n275 VDDA.n274 96.8409
R5523 VDDA.n273 VDDA.n272 96.8409
R5524 VDDA.n271 VDDA.n270 96.8409
R5525 VDDA.n269 VDDA.n268 96.8409
R5526 VDDA.n267 VDDA.n266 96.8409
R5527 VDDA.n225 VDDA.n224 96.8409
R5528 VDDA.n223 VDDA.n222 96.8409
R5529 VDDA.n221 VDDA.n220 96.8409
R5530 VDDA.n219 VDDA.n218 96.8409
R5531 VDDA.n217 VDDA.n216 96.8409
R5532 VDDA.n383 VDDA.n382 96.0005
R5533 VDDA.n384 VDDA.n370 96.0005
R5534 VDDA.n391 VDDA.n390 96.0005
R5535 VDDA.n422 VDDA.t217 93.3041
R5536 VDDA.t355 VDDA.n422 93.3041
R5537 VDDA.n387 VDDA.t215 93.3041
R5538 VDDA.n387 VDDA.t186 93.3041
R5539 VDDA.n434 VDDA.n433 92.5005
R5540 VDDA.t329 VDDA.n434 92.5005
R5541 VDDA.n435 VDDA.n432 92.5005
R5542 VDDA.t329 VDDA.n435 92.5005
R5543 VDDA.n439 VDDA.n438 92.5005
R5544 VDDA.n448 VDDA.n439 92.5005
R5545 VDDA.n440 VDDA.n437 92.5005
R5546 VDDA.n449 VDDA.n440 92.5005
R5547 VDDA.n421 VDDA.n420 92.5005
R5548 VDDA.n397 VDDA.n396 92.5005
R5549 VDDA.n422 VDDA.n397 92.5005
R5550 VDDA.n424 VDDA.n423 92.5005
R5551 VDDA.n398 VDDA.n395 92.5005
R5552 VDDA.n422 VDDA.n398 92.5005
R5553 VDDA.n378 VDDA.n371 92.5005
R5554 VDDA.n379 VDDA.n378 92.5005
R5555 VDDA.n377 VDDA.n376 92.5005
R5556 VDDA.n381 VDDA.n380 92.5005
R5557 VDDA.n380 VDDA.n379 92.5005
R5558 VDDA.n383 VDDA.n372 92.5005
R5559 VDDA.n386 VDDA.n366 92.5005
R5560 VDDA.n387 VDDA.n386 92.5005
R5561 VDDA.n385 VDDA.n384 92.5005
R5562 VDDA.n389 VDDA.n388 92.5005
R5563 VDDA.n388 VDDA.n387 92.5005
R5564 VDDA.n391 VDDA.n367 92.5005
R5565 VDDA.n339 VDDA.n338 92.5005
R5566 VDDA.n335 VDDA.n334 92.5005
R5567 VDDA.n337 VDDA.n335 92.5005
R5568 VDDA.n336 VDDA.n328 92.5005
R5569 VDDA.n340 VDDA.n329 92.5005
R5570 VDDA.n337 VDDA.n329 92.5005
R5571 VDDA.n359 VDDA.n358 92.5005
R5572 VDDA.n358 VDDA.n357 92.5005
R5573 VDDA.n356 VDDA.n355 92.5005
R5574 VDDA.n357 VDDA.n356 92.5005
R5575 VDDA.n319 VDDA.n318 92.5005
R5576 VDDA.n315 VDDA.n314 92.5005
R5577 VDDA.n317 VDDA.n315 92.5005
R5578 VDDA.n316 VDDA.n308 92.5005
R5579 VDDA.n320 VDDA.n309 92.5005
R5580 VDDA.n317 VDDA.n309 92.5005
R5581 VDDA.n295 VDDA.n294 92.5005
R5582 VDDA.n291 VDDA.n290 92.5005
R5583 VDDA.n293 VDDA.n291 92.5005
R5584 VDDA.n292 VDDA.n284 92.5005
R5585 VDDA.n296 VDDA.n285 92.5005
R5586 VDDA.n293 VDDA.n285 92.5005
R5587 VDDA.n239 VDDA.n238 92.5005
R5588 VDDA.n235 VDDA.n234 92.5005
R5589 VDDA.n237 VDDA.n235 92.5005
R5590 VDDA.n236 VDDA.n228 92.5005
R5591 VDDA.n240 VDDA.n229 92.5005
R5592 VDDA.n237 VDDA.n229 92.5005
R5593 VDDA.n244 VDDA.n241 92.5005
R5594 VDDA.n258 VDDA.n244 92.5005
R5595 VDDA.n243 VDDA.n242 92.5005
R5596 VDDA.n258 VDDA.n243 92.5005
R5597 VDDA.n204 VDDA.n203 92.5005
R5598 VDDA.n150 VDDA.n148 92.5005
R5599 VDDA.n201 VDDA.n150 92.5005
R5600 VDDA.n200 VDDA.n199 92.5005
R5601 VDDA.n149 VDDA.n147 92.5005
R5602 VDDA.n202 VDDA.n149 92.5005
R5603 VDDA.n190 VDDA.n189 92.5005
R5604 VDDA.n156 VDDA.n154 92.5005
R5605 VDDA.n188 VDDA.n156 92.5005
R5606 VDDA.n187 VDDA.n186 92.5005
R5607 VDDA.n155 VDDA.n153 92.5005
R5608 VDDA.n188 VDDA.n155 92.5005
R5609 VDDA.n171 VDDA.n170 92.5005
R5610 VDDA.n162 VDDA.n160 92.5005
R5611 VDDA.n169 VDDA.n162 92.5005
R5612 VDDA.n168 VDDA.n167 92.5005
R5613 VDDA.n161 VDDA.n159 92.5005
R5614 VDDA.n169 VDDA.n161 92.5005
R5615 VDDA.n138 VDDA.n137 92.5005
R5616 VDDA.n133 VDDA.n132 92.5005
R5617 VDDA.n136 VDDA.n133 92.5005
R5618 VDDA.n135 VDDA.n134 92.5005
R5619 VDDA.n140 VDDA.n130 92.5005
R5620 VDDA.n136 VDDA.n130 92.5005
R5621 VDDA.n124 VDDA.n123 92.5005
R5622 VDDA.n89 VDDA.n87 92.5005
R5623 VDDA.n122 VDDA.n89 92.5005
R5624 VDDA.n121 VDDA.n120 92.5005
R5625 VDDA.n88 VDDA.n86 92.5005
R5626 VDDA.n122 VDDA.n88 92.5005
R5627 VDDA.n100 VDDA.n99 92.5005
R5628 VDDA.n95 VDDA.n94 92.5005
R5629 VDDA.n98 VDDA.n95 92.5005
R5630 VDDA.n97 VDDA.n96 92.5005
R5631 VDDA.n102 VDDA.n92 92.5005
R5632 VDDA.n98 VDDA.n92 92.5005
R5633 VDDA.n59 VDDA.n11 92.5005
R5634 VDDA.n77 VDDA.n11 92.5005
R5635 VDDA.n79 VDDA.n78 92.5005
R5636 VDDA.n73 VDDA.n12 92.5005
R5637 VDDA.n77 VDDA.n12 92.5005
R5638 VDDA.n76 VDDA.n75 92.5005
R5639 VDDA.n33 VDDA.n32 92.5005
R5640 VDDA.n29 VDDA.n28 92.5005
R5641 VDDA.n31 VDDA.n29 92.5005
R5642 VDDA.n30 VDDA.n22 92.5005
R5643 VDDA.n34 VDDA.n23 92.5005
R5644 VDDA.n31 VDDA.n23 92.5005
R5645 VDDA.n379 VDDA.t228 91.6672
R5646 VDDA.n379 VDDA.t305 91.6672
R5647 VDDA.n443 VDDA.n442 87.4672
R5648 VDDA.n77 VDDA.t341 86.3641
R5649 VDDA.t118 VDDA.n77 86.3641
R5650 VDDA.n31 VDDA.t260 86.3641
R5651 VDDA.t290 VDDA.n31 86.3641
R5652 VDDA.n442 VDDA.t8 85.438
R5653 VDDA.n454 VDDA.t23 85.438
R5654 VDDA.n448 VDDA.t7 81.3068
R5655 VDDA.n454 VDDA.n453 81.0672
R5656 VDDA.n444 VDDA.n442 81.0672
R5657 VDDA.n122 VDDA.t307 79.907
R5658 VDDA.t141 VDDA.n122 79.907
R5659 VDDA.t402 VDDA.n202 79.1672
R5660 VDDA.n136 VDDA.t414 79.1672
R5661 VDDA.t396 VDDA.n136 79.1672
R5662 VDDA.n98 VDDA.t282 79.1672
R5663 VDDA.t281 VDDA.n98 79.1672
R5664 VDDA.n393 VDDA.t194 78.8005
R5665 VDDA.n393 VDDA.t362 78.8005
R5666 VDDA.n399 VDDA.t350 78.8005
R5667 VDDA.n399 VDDA.t319 78.8005
R5668 VDDA.n401 VDDA.t354 78.8005
R5669 VDDA.n401 VDDA.t165 78.8005
R5670 VDDA.n403 VDDA.t360 78.8005
R5671 VDDA.n403 VDDA.t263 78.8005
R5672 VDDA.n405 VDDA.t356 78.8005
R5673 VDDA.n405 VDDA.t366 78.8005
R5674 VDDA.n407 VDDA.t277 78.8005
R5675 VDDA.n407 VDDA.t218 78.8005
R5676 VDDA.n409 VDDA.t167 78.8005
R5677 VDDA.n409 VDDA.t364 78.8005
R5678 VDDA.n411 VDDA.t265 78.8005
R5679 VDDA.n411 VDDA.t348 78.8005
R5680 VDDA.n413 VDDA.t192 78.8005
R5681 VDDA.n413 VDDA.t358 78.8005
R5682 VDDA.n415 VDDA.t220 78.8005
R5683 VDDA.n415 VDDA.t352 78.8005
R5684 VDDA.n188 VDDA.t398 77.9856
R5685 VDDA.t410 VDDA.n188 77.9856
R5686 VDDA.n169 VDDA.t400 77.9856
R5687 VDDA.t412 VDDA.n169 77.9856
R5688 VDDA.n452 VDDA.n437 64.0005
R5689 VDDA.n102 VDDA.n101 64.0005
R5690 VDDA.n102 VDDA.n91 64.0005
R5691 VDDA.n71 VDDA.n13 64.0005
R5692 VDDA.n63 VDDA.n13 64.0005
R5693 VDDA.n63 VDDA.n62 64.0005
R5694 VDDA.n62 VDDA.n59 64.0005
R5695 VDDA.n59 VDDA.n58 64.0005
R5696 VDDA.n58 VDDA.n50 64.0005
R5697 VDDA.n50 VDDA.n8 64.0005
R5698 VDDA.n80 VDDA.n8 64.0005
R5699 VDDA.t124 VDDA.t31 62.9523
R5700 VDDA.t173 VDDA.t124 62.9523
R5701 VDDA.t159 VDDA.t173 62.9523
R5702 VDDA.t425 VDDA.t159 62.9523
R5703 VDDA.t128 VDDA.t425 62.9523
R5704 VDDA.t157 VDDA.t136 62.9523
R5705 VDDA.t136 VDDA.t284 62.9523
R5706 VDDA.t284 VDDA.t122 62.9523
R5707 VDDA.t122 VDDA.t126 62.9523
R5708 VDDA.t126 VDDA.t49 62.9523
R5709 VDDA.t0 VDDA.t43 62.9523
R5710 VDDA.t303 VDDA.t0 62.9523
R5711 VDDA.t467 VDDA.t303 62.9523
R5712 VDDA.t457 VDDA.t467 62.9523
R5713 VDDA.t301 VDDA.t457 62.9523
R5714 VDDA.t320 VDDA.t454 62.9523
R5715 VDDA.t459 VDDA.t320 62.9523
R5716 VDDA.t322 VDDA.t459 62.9523
R5717 VDDA.t211 VDDA.t322 62.9523
R5718 VDDA.t67 VDDA.t211 62.9523
R5719 VDDA.n140 VDDA.n139 62.7205
R5720 VDDA.n140 VDDA.n129 62.7205
R5721 VDDA.n430 VDDA.t330 62.5402
R5722 VDDA.n430 VDDA.t71 62.5402
R5723 VDDA.n461 VDDA.n460 61.6672
R5724 VDDA.n463 VDDA.n462 61.6672
R5725 VDDA.n352 VDDA.n327 61.6672
R5726 VDDA.n354 VDDA.n353 61.6672
R5727 VDDA.n260 VDDA.n259 61.6672
R5728 VDDA.n257 VDDA.n256 61.6672
R5729 VDDA.n337 VDDA.t170 60.7563
R5730 VDDA.t156 VDDA.n337 60.7563
R5731 VDDA.n237 VDDA.t210 60.7563
R5732 VDDA.t368 VDDA.n237 60.7563
R5733 VDDA.n1 VDDA.t470 59.5681
R5734 VDDA.n0 VDDA.t469 59.5681
R5735 VDDA.n459 VDDA.n432 57.6005
R5736 VDDA.n464 VDDA.n432 57.6005
R5737 VDDA.n201 VDDA.t380 57.5763
R5738 VDDA.n0 VDDA.t471 51.8887
R5739 VDDA.n445 VDDA.n437 51.2005
R5740 VDDA.n317 VDDA.t130 49.1384
R5741 VDDA.t374 VDDA.n317 49.1384
R5742 VDDA.n293 VDDA.t213 49.1384
R5743 VDDA.t184 VDDA.n293 49.1384
R5744 VDDA.n2 VDDA.t472 48.9557
R5745 VDDA.n467 VDDA.n466 48.3605
R5746 VDDA.n457 VDDA.n456 43.8605
R5747 VDDA.n417 VDDA.n416 42.0963
R5748 VDDA.n428 VDDA.n427 41.5338
R5749 VDDA.n145 VDDA.t403 39.4005
R5750 VDDA.n145 VDDA.t391 39.4005
R5751 VDDA.n194 VDDA.t405 39.4005
R5752 VDDA.n194 VDDA.t381 39.4005
R5753 VDDA.n151 VDDA.t409 39.4005
R5754 VDDA.n151 VDDA.t389 39.4005
R5755 VDDA.n175 VDDA.t411 39.4005
R5756 VDDA.n175 VDDA.t393 39.4005
R5757 VDDA.n177 VDDA.t417 39.4005
R5758 VDDA.n177 VDDA.t399 39.4005
R5759 VDDA.n179 VDDA.t407 39.4005
R5760 VDDA.n179 VDDA.t385 39.4005
R5761 VDDA.n181 VDDA.t383 39.4005
R5762 VDDA.n181 VDDA.t387 39.4005
R5763 VDDA.n157 VDDA.t413 39.4005
R5764 VDDA.n157 VDDA.t395 39.4005
R5765 VDDA.n163 VDDA.t379 39.4005
R5766 VDDA.n163 VDDA.t401 39.4005
R5767 VDDA.n141 VDDA.t415 39.4005
R5768 VDDA.n141 VDDA.t397 39.4005
R5769 VDDA.n5 VDDA.t243 39.4005
R5770 VDDA.n5 VDDA.t251 39.4005
R5771 VDDA.n6 VDDA.t339 39.4005
R5772 VDDA.n6 VDDA.t235 39.4005
R5773 VDDA.n52 VDDA.t438 39.4005
R5774 VDDA.n52 VDDA.t346 39.4005
R5775 VDDA.n56 VDDA.t237 39.4005
R5776 VDDA.n56 VDDA.t253 39.4005
R5777 VDDA.n48 VDDA.t342 39.4005
R5778 VDDA.n48 VDDA.t119 39.4005
R5779 VDDA.n60 VDDA.t440 39.4005
R5780 VDDA.n60 VDDA.t133 39.4005
R5781 VDDA.n47 VDDA.t423 39.4005
R5782 VDDA.n47 VDDA.t255 39.4005
R5783 VDDA.n66 VDDA.t344 39.4005
R5784 VDDA.n66 VDDA.t121 39.4005
R5785 VDDA.n14 VDDA.t442 39.4005
R5786 VDDA.n14 VDDA.t135 39.4005
R5787 VDDA.n44 VDDA.t249 39.4005
R5788 VDDA.n44 VDDA.t273 39.4005
R5789 VDDA.n42 VDDA.t430 39.4005
R5790 VDDA.n42 VDDA.t280 39.4005
R5791 VDDA.n40 VDDA.t204 39.4005
R5792 VDDA.n40 VDDA.t462 39.4005
R5793 VDDA.n38 VDDA.t432 39.4005
R5794 VDDA.n38 VDDA.t239 39.4005
R5795 VDDA.n35 VDDA.t261 39.4005
R5796 VDDA.n35 VDDA.t291 39.4005
R5797 VDDA.n20 VDDA.t271 39.4005
R5798 VDDA.n20 VDDA.t200 39.4005
R5799 VDDA.n18 VDDA.t297 39.4005
R5800 VDDA.n18 VDDA.t206 39.4005
R5801 VDDA.n16 VDDA.t315 39.4005
R5802 VDDA.n16 VDDA.t449 39.4005
R5803 VDDA.n15 VDDA.t269 39.4005
R5804 VDDA.n15 VDDA.t313 39.4005
R5805 VDDA.n357 VDDA.t128 31.4764
R5806 VDDA.n357 VDDA.t157 31.4764
R5807 VDDA.n258 VDDA.t301 31.4764
R5808 VDDA.t454 VDDA.n258 31.4764
R5809 VDDA.n384 VDDA.n383 28.663
R5810 VDDA.n214 VDDA.n3 28.3337
R5811 VDDA.n466 VDDA.n465 25.6005
R5812 VDDA.n458 VDDA.n457 25.6005
R5813 VDDA.n427 VDDA.n426 25.6005
R5814 VDDA.n418 VDDA.n417 25.6005
R5815 VDDA.n465 VDDA.n464 24.5338
R5816 VDDA.n459 VDDA.n458 24.5338
R5817 VDDA.n453 VDDA.n452 24.5338
R5818 VDDA.n445 VDDA.n444 24.5338
R5819 VDDA.n202 VDDA.n201 21.5914
R5820 VDDA.n426 VDDA.n425 21.3338
R5821 VDDA.n419 VDDA.n418 21.3338
R5822 VDDA.n375 VDDA.n374 21.3338
R5823 VDDA.n382 VDDA.n373 21.3338
R5824 VDDA.n370 VDDA.n369 21.3338
R5825 VDDA.n390 VDDA.n368 21.3338
R5826 VDDA.n333 VDDA.n332 21.3338
R5827 VDDA.n331 VDDA.n330 21.3338
R5828 VDDA.n361 VDDA.n360 21.3338
R5829 VDDA.n351 VDDA.n350 21.3338
R5830 VDDA.n313 VDDA.n312 21.3338
R5831 VDDA.n311 VDDA.n310 21.3338
R5832 VDDA.n289 VDDA.n288 21.3338
R5833 VDDA.n287 VDDA.n286 21.3338
R5834 VDDA.n233 VDDA.n232 21.3338
R5835 VDDA.n231 VDDA.n230 21.3338
R5836 VDDA.n262 VDDA.n261 21.3338
R5837 VDDA.n255 VDDA.n254 21.3338
R5838 VDDA.n129 VDDA.n128 21.3338
R5839 VDDA.n139 VDDA.n131 21.3338
R5840 VDDA.n91 VDDA.n90 21.3338
R5841 VDDA.n101 VDDA.n93 21.3338
R5842 VDDA.n74 VDDA.n72 21.3338
R5843 VDDA.n10 VDDA.n9 21.3338
R5844 VDDA.n27 VDDA.n26 21.3338
R5845 VDDA.n25 VDDA.n24 21.3338
R5846 VDDA.n276 VDDA.n275 21.1567
R5847 VDDA.n392 VDDA.n391 19.5505
R5848 VDDA.n359 VDDA.n340 19.538
R5849 VDDA.n241 VDDA.n240 19.538
R5850 VDDA.n469 VDDA.n468 19.4142
R5851 VDDA.n322 VDDA.n320 19.2005
R5852 VDDA.n298 VDDA.n296 19.2005
R5853 VDDA.n206 VDDA.n205 19.2005
R5854 VDDA.n198 VDDA.n197 19.2005
R5855 VDDA.n192 VDDA.n191 19.2005
R5856 VDDA.n185 VDDA.n184 19.2005
R5857 VDDA.n173 VDDA.n172 19.2005
R5858 VDDA.n166 VDDA.n165 19.2005
R5859 VDDA.n126 VDDA.n125 19.2005
R5860 VDDA.n119 VDDA.n118 19.2005
R5861 VDDA.n447 VDDA.n446 18.5005
R5862 VDDA.n451 VDDA.n450 18.5005
R5863 VDDA.t331 VDDA.n449 17.1176
R5864 VDDA.n365 VDDA.n225 16.8443
R5865 VDDA.n117 VDDA.n102 16.363
R5866 VDDA.n213 VDDA.t226 15.0181
R5867 VDDA.n165 VDDA.n164 14.363
R5868 VDDA.n443 VDDA.n436 14.0505
R5869 VDDA.n197 VDDA.n196 13.8005
R5870 VDDA.n184 VDDA.n183 13.8005
R5871 VDDA.n174 VDDA.n173 13.8005
R5872 VDDA.n193 VDDA.n192 13.8005
R5873 VDDA.n207 VDDA.n206 13.8005
R5874 VDDA.n118 VDDA.n117 13.8005
R5875 VDDA.n127 VDDA.n126 13.8005
R5876 VDDA.n84 VDDA.t300 13.1338
R5877 VDDA.n84 VDDA.t293 13.1338
R5878 VDDA.n103 VDDA.t444 13.1338
R5879 VDDA.n103 VDDA.t198 13.1338
R5880 VDDA.n105 VDDA.t222 13.1338
R5881 VDDA.n105 VDDA.t225 13.1338
R5882 VDDA.n107 VDDA.t142 13.1338
R5883 VDDA.n107 VDDA.t179 13.1338
R5884 VDDA.n109 VDDA.t182 13.1338
R5885 VDDA.n109 VDDA.t308 13.1338
R5886 VDDA.n111 VDDA.t209 13.1338
R5887 VDDA.n111 VDDA.t241 13.1338
R5888 VDDA.n113 VDDA.t245 13.1338
R5889 VDDA.n113 VDDA.t451 13.1338
R5890 VDDA.n115 VDDA.t196 13.1338
R5891 VDDA.n115 VDDA.t295 13.1338
R5892 VDDA.t8 VDDA.n441 12.313
R5893 VDDA.n441 VDDA.t332 12.313
R5894 VDDA.n321 VDDA.t131 11.2576
R5895 VDDA.n321 VDDA.t375 11.2576
R5896 VDDA.n305 VDDA.t163 11.2576
R5897 VDDA.n305 VDDA.t172 11.2576
R5898 VDDA.n304 VDDA.t188 11.2576
R5899 VDDA.n304 VDDA.t447 11.2576
R5900 VDDA.n302 VDDA.t421 11.2576
R5901 VDDA.n302 VDDA.t334 11.2576
R5902 VDDA.n301 VDDA.t148 11.2576
R5903 VDDA.n301 VDDA.t419 11.2576
R5904 VDDA.n297 VDDA.t214 11.2576
R5905 VDDA.n297 VDDA.t185 11.2576
R5906 VDDA.n281 VDDA.t336 11.2576
R5907 VDDA.n281 VDDA.t377 11.2576
R5908 VDDA.n280 VDDA.t150 11.2576
R5909 VDDA.n280 VDDA.t152 11.2576
R5910 VDDA.n278 VDDA.t154 11.2576
R5911 VDDA.n278 VDDA.t465 11.2576
R5912 VDDA.n277 VDDA.t370 11.2576
R5913 VDDA.n277 VDDA.t435 11.2576
R5914 VDDA.n323 VDDA.n322 9.3005
R5915 VDDA.n299 VDDA.n298 9.3005
R5916 VDDA.n142 VDDA.n140 9.3005
R5917 VDDA.n67 VDDA.n13 9.3005
R5918 VDDA.n64 VDDA.n63 9.3005
R5919 VDDA.n62 VDDA.n61 9.3005
R5920 VDDA.n59 VDDA.n49 9.3005
R5921 VDDA.n58 VDDA.n57 9.3005
R5922 VDDA.n53 VDDA.n50 9.3005
R5923 VDDA.n8 VDDA.n7 9.3005
R5924 VDDA.n81 VDDA.n80 9.3005
R5925 VDDA.n71 VDDA.n70 9.3005
R5926 VDDA.n36 VDDA.n34 9.3005
R5927 VDDA.n456 VDDA.n455 8.53175
R5928 VDDA.n3 VDDA.n2 8.03219
R5929 VDDA.n274 VDDA.t278 8.0005
R5930 VDDA.n274 VDDA.t233 8.0005
R5931 VDDA.n272 VDDA.t453 8.0005
R5932 VDDA.n272 VDDA.t310 8.0005
R5933 VDDA.n270 VDDA.t463 8.0005
R5934 VDDA.n270 VDDA.t325 8.0005
R5935 VDDA.n268 VDDA.t328 8.0005
R5936 VDDA.n268 VDDA.t311 8.0005
R5937 VDDA.n266 VDDA.t309 8.0005
R5938 VDDA.n266 VDDA.t456 8.0005
R5939 VDDA.n265 VDDA.t231 8.0005
R5940 VDDA.n265 VDDA.t267 8.0005
R5941 VDDA.n224 VDDA.t230 8.0005
R5942 VDDA.n224 VDDA.t286 8.0005
R5943 VDDA.n222 VDDA.t427 8.0005
R5944 VDDA.n222 VDDA.t287 8.0005
R5945 VDDA.n220 VDDA.t428 8.0005
R5946 VDDA.n220 VDDA.t138 8.0005
R5947 VDDA.n218 VDDA.t176 8.0005
R5948 VDDA.n218 VDDA.t201 8.0005
R5949 VDDA.n216 VDDA.t175 8.0005
R5950 VDDA.n216 VDDA.t161 8.0005
R5951 VDDA.n215 VDDA.t317 8.0005
R5952 VDDA.n215 VDDA.t232 8.0005
R5953 VDDA.n208 VDDA.n207 7.44175
R5954 VDDA.n429 VDDA.n428 7.438
R5955 VDDA.n325 VDDA.t125 6.56717
R5956 VDDA.n325 VDDA.t174 6.56717
R5957 VDDA.n341 VDDA.t160 6.56717
R5958 VDDA.n341 VDDA.t426 6.56717
R5959 VDDA.n343 VDDA.t129 6.56717
R5960 VDDA.n343 VDDA.t158 6.56717
R5961 VDDA.n345 VDDA.t137 6.56717
R5962 VDDA.n345 VDDA.t285 6.56717
R5963 VDDA.n347 VDDA.t123 6.56717
R5964 VDDA.n347 VDDA.t127 6.56717
R5965 VDDA.n226 VDDA.t323 6.56717
R5966 VDDA.n226 VDDA.t212 6.56717
R5967 VDDA.n245 VDDA.t321 6.56717
R5968 VDDA.n245 VDDA.t460 6.56717
R5969 VDDA.n247 VDDA.t302 6.56717
R5970 VDDA.n247 VDDA.t455 6.56717
R5971 VDDA.n249 VDDA.t468 6.56717
R5972 VDDA.n249 VDDA.t458 6.56717
R5973 VDDA.n251 VDDA.t1 6.56717
R5974 VDDA.n251 VDDA.t304 6.56717
R5975 VDDA.n324 VDDA.n300 6.313
R5976 VDDA.n144 VDDA.n143 6.13371
R5977 VDDA.n83 VDDA.n82 6.098
R5978 VDDA.n468 VDDA.n467 6.0005
R5979 VDDA.n469 VDDA 5.6546
R5980 VDDA.n456 VDDA.n431 5.1255
R5981 VDDA.n324 VDDA.n323 5.063
R5982 VDDA.n300 VDDA.n299 5.063
R5983 VDDA.n323 VDDA.n307 4.5005
R5984 VDDA.n299 VDDA.n283 4.5005
R5985 VDDA.n365 VDDA.n364 4.5005
R5986 VDDA.n143 VDDA.n142 4.5005
R5987 VDDA.n37 VDDA.n36 4.5005
R5988 VDDA.n70 VDDA.n69 4.5005
R5989 VDDA.n68 VDDA.n67 4.5005
R5990 VDDA.n65 VDDA.n64 4.5005
R5991 VDDA.n61 VDDA.n46 4.5005
R5992 VDDA.n51 VDDA.n49 4.5005
R5993 VDDA.n57 VDDA.n55 4.5005
R5994 VDDA.n54 VDDA.n53 4.5005
R5995 VDDA.n7 VDDA.n4 4.5005
R5996 VDDA.n82 VDDA.n81 4.5005
R5997 VDDA.n449 VDDA.n448 4.27978
R5998 VDDA.n1 VDDA.n0 4.12334
R5999 VDDA.n214 VDDA 4.08025
R6000 VDDA VDDA.n469 3.7135
R6001 VDDA.n300 VDDA.n276 3.688
R6002 VDDA.n364 VDDA.n324 3.5005
R6003 VDDA.n69 VDDA.n45 3.3755
R6004 VDDA.n2 VDDA.n1 2.93377
R6005 VDDA.n429 VDDA.n392 2.813
R6006 VDDA.n468 VDDA.n429 2.563
R6007 VDDA.n196 VDDA.n193 2.5005
R6008 VDDA.n143 VDDA.n127 2.47371
R6009 VDDA.n183 VDDA.n174 1.813
R6010 VDDA.n392 VDDA.n365 1.46925
R6011 VDDA VDDA.n213 1.0815
R6012 VDDA.n117 VDDA.n116 1.0005
R6013 VDDA.n116 VDDA.n114 1.0005
R6014 VDDA.n114 VDDA.n112 1.0005
R6015 VDDA.n112 VDDA.n110 1.0005
R6016 VDDA.n110 VDDA.n108 1.0005
R6017 VDDA.n108 VDDA.n106 1.0005
R6018 VDDA.n106 VDDA.n104 1.0005
R6019 VDDA.n104 VDDA.n85 1.0005
R6020 VDDA.n127 VDDA.n85 1.0005
R6021 VDDA.n364 VDDA.n363 0.938
R6022 VDDA.n83 VDDA.n3 0.840625
R6023 VDDA.n276 VDDA.n264 0.7505
R6024 VDDA.n144 VDDA.n83 0.74075
R6025 VDDA.n455 VDDA.n436 0.6255
R6026 VDDA.n307 VDDA.n306 0.6255
R6027 VDDA.n307 VDDA.n303 0.6255
R6028 VDDA.n283 VDDA.n282 0.6255
R6029 VDDA.n283 VDDA.n279 0.6255
R6030 VDDA.n19 VDDA.n17 0.6255
R6031 VDDA.n21 VDDA.n19 0.6255
R6032 VDDA.n37 VDDA.n21 0.6255
R6033 VDDA.n39 VDDA.n37 0.6255
R6034 VDDA.n41 VDDA.n39 0.6255
R6035 VDDA.n43 VDDA.n41 0.6255
R6036 VDDA.n45 VDDA.n43 0.6255
R6037 VDDA.n69 VDDA.n68 0.6255
R6038 VDDA.n68 VDDA.n65 0.6255
R6039 VDDA.n65 VDDA.n46 0.6255
R6040 VDDA.n51 VDDA.n46 0.6255
R6041 VDDA.n55 VDDA.n51 0.6255
R6042 VDDA.n55 VDDA.n54 0.6255
R6043 VDDA.n54 VDDA.n4 0.6255
R6044 VDDA.n82 VDDA.n4 0.6255
R6045 VDDA.n416 VDDA.n414 0.563
R6046 VDDA.n414 VDDA.n412 0.563
R6047 VDDA.n412 VDDA.n410 0.563
R6048 VDDA.n410 VDDA.n408 0.563
R6049 VDDA.n408 VDDA.n406 0.563
R6050 VDDA.n406 VDDA.n404 0.563
R6051 VDDA.n404 VDDA.n402 0.563
R6052 VDDA.n402 VDDA.n400 0.563
R6053 VDDA.n400 VDDA.n394 0.563
R6054 VDDA.n428 VDDA.n394 0.563
R6055 VDDA.n348 VDDA.n346 0.563
R6056 VDDA.n346 VDDA.n344 0.563
R6057 VDDA.n344 VDDA.n342 0.563
R6058 VDDA.n342 VDDA.n326 0.563
R6059 VDDA.n363 VDDA.n326 0.563
R6060 VDDA.n269 VDDA.n267 0.563
R6061 VDDA.n271 VDDA.n269 0.563
R6062 VDDA.n273 VDDA.n271 0.563
R6063 VDDA.n275 VDDA.n273 0.563
R6064 VDDA.n252 VDDA.n250 0.563
R6065 VDDA.n250 VDDA.n248 0.563
R6066 VDDA.n248 VDDA.n246 0.563
R6067 VDDA.n246 VDDA.n227 0.563
R6068 VDDA.n264 VDDA.n227 0.563
R6069 VDDA.n219 VDDA.n217 0.563
R6070 VDDA.n221 VDDA.n219 0.563
R6071 VDDA.n223 VDDA.n221 0.563
R6072 VDDA.n225 VDDA.n223 0.563
R6073 VDDA.n164 VDDA.n158 0.563
R6074 VDDA.n174 VDDA.n158 0.563
R6075 VDDA.n183 VDDA.n182 0.563
R6076 VDDA.n182 VDDA.n180 0.563
R6077 VDDA.n180 VDDA.n178 0.563
R6078 VDDA.n178 VDDA.n176 0.563
R6079 VDDA.n176 VDDA.n152 0.563
R6080 VDDA.n193 VDDA.n152 0.563
R6081 VDDA.n196 VDDA.n195 0.563
R6082 VDDA.n195 VDDA.n146 0.563
R6083 VDDA.n207 VDDA.n146 0.563
R6084 VDDA.n208 VDDA.n144 0.546875
R6085 VDDA.n213 VDDA.n208 0.370625
R6086 VDDA.n467 VDDA.n431 0.2505
R6087 VDDA VDDA.n214 0.2355
R6088 VDDA.t183 VDDA.t289 0.1603
R6089 VDDA.t298 VDDA.t445 0.1603
R6090 VDDA.t180 VDDA.t139 0.1603
R6091 VDDA.t143 VDDA.t246 0.1603
R6092 VDDA.t452 VDDA.t274 0.1603
R6093 VDDA.t247 VDDA.t223 0.1603
R6094 VDDA.t275 VDDA.t140 0.1603
R6095 VDDA.t306 VDDA.t288 0.1603
R6096 VDDA.n210 VDDA.t257 0.159278
R6097 VDDA.n211 VDDA.t207 0.159278
R6098 VDDA.n212 VDDA.t256 0.159278
R6099 VDDA.n212 VDDA.t183 0.1368
R6100 VDDA.n212 VDDA.t298 0.1368
R6101 VDDA.n211 VDDA.t180 0.1368
R6102 VDDA.n211 VDDA.t143 0.1368
R6103 VDDA.n210 VDDA.t452 0.1368
R6104 VDDA.n210 VDDA.t247 0.1368
R6105 VDDA.n209 VDDA.t275 0.1368
R6106 VDDA.n209 VDDA.t306 0.1368
R6107 VDDA.t257 VDDA.n209 0.00152174
R6108 VDDA.t207 VDDA.n210 0.00152174
R6109 VDDA.t256 VDDA.n211 0.00152174
R6110 VDDA.t226 VDDA.n212 0.00152174
R6111 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 610.534
R6112 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 610.534
R6113 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R6114 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R6115 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R6116 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R6117 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R6118 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R6119 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R6120 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R6121 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R6122 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R6123 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R6124 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R6125 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R6126 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R6127 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R6128 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R6129 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R6130 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R6131 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 339.836
R6132 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.834
R6133 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R6134 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 334.772
R6135 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 221.293
R6136 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R6137 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R6138 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R6139 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R6140 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R6141 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R6142 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R6143 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R6144 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R6145 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R6146 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 176.733
R6147 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R6148 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R6149 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R6150 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R6151 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R6152 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 117.825
R6153 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n29 84.9693
R6154 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 65.2045
R6155 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 56.2338
R6156 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 56.2338
R6157 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 53.2453
R6158 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R6159 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 39.4005
R6160 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R6161 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 39.4005
R6162 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R6163 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 39.4005
R6164 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R6165 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 39.4005
R6166 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n6 18.3755
R6167 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 16.0005
R6168 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 16.0005
R6169 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 16.0005
R6170 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 16.0005
R6171 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 4.5005
R6172 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R6173 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6174 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6175 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 322.692
R6176 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6177 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 270.591
R6178 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 270.591
R6179 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 270.591
R6180 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 270.591
R6181 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6182 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6183 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6184 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6185 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6186 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6187 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 174.726
R6188 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 174.726
R6189 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 174.726
R6190 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 174.726
R6191 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.215
R6192 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.215
R6193 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.215
R6194 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 129.24
R6195 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6196 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 129.24
R6197 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6198 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6199 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6200 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 49.6255
R6201 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6202 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6203 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6204 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6205 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6206 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6207 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6208 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6209 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6210 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 3.688
R6211 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref 3.2505
R6212 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 3.1255
R6213 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 1.2755
R6214 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 1.2755
R6215 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 0.8005
R6216 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 0.8005
R6217 bgr_0.V_p_2.n5 bgr_0.V_p_2.n0 229.562
R6218 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R6219 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R6220 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 228.939
R6221 bgr_0.V_p_2.n0 bgr_0.V_p_2.n1 228.939
R6222 bgr_0.V_p_2.n0 bgr_0.V_p_2.t0 100.103
R6223 bgr_0.V_p_2.n4 bgr_0.V_p_2.t10 48.0005
R6224 bgr_0.V_p_2.n4 bgr_0.V_p_2.t5 48.0005
R6225 bgr_0.V_p_2.n3 bgr_0.V_p_2.t4 48.0005
R6226 bgr_0.V_p_2.n3 bgr_0.V_p_2.t8 48.0005
R6227 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R6228 bgr_0.V_p_2.n2 bgr_0.V_p_2.t7 48.0005
R6229 bgr_0.V_p_2.n1 bgr_0.V_p_2.t3 48.0005
R6230 bgr_0.V_p_2.n1 bgr_0.V_p_2.t9 48.0005
R6231 bgr_0.V_p_2.n5 bgr_0.V_p_2.t6 48.0005
R6232 bgr_0.V_p_2.t1 bgr_0.V_p_2.n5 48.0005
R6233 bgr_0.V_mir2.n4 bgr_0.V_mir2.n0 325.473
R6234 bgr_0.V_mir2.n9 bgr_0.V_mir2.n5 325.471
R6235 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.471
R6236 bgr_0.V_mir2.n16 bgr_0.V_mir2.t22 310.488
R6237 bgr_0.V_mir2.n6 bgr_0.V_mir2.t21 310.488
R6238 bgr_0.V_mir2.n1 bgr_0.V_mir2.t20 310.488
R6239 bgr_0.V_mir2.n12 bgr_0.V_mir2.t13 278.312
R6240 bgr_0.V_mir2.n12 bgr_0.V_mir2.n11 228.939
R6241 bgr_0.V_mir2.n13 bgr_0.V_mir2.n10 224.439
R6242 bgr_0.V_mir2.n18 bgr_0.V_mir2.t10 184.097
R6243 bgr_0.V_mir2.n8 bgr_0.V_mir2.t2 184.097
R6244 bgr_0.V_mir2.n3 bgr_0.V_mir2.t4 184.097
R6245 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6246 bgr_0.V_mir2.n7 bgr_0.V_mir2.n6 167.094
R6247 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 167.094
R6248 bgr_0.V_mir2.n9 bgr_0.V_mir2.n8 152
R6249 bgr_0.V_mir2.n4 bgr_0.V_mir2.n3 152
R6250 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6251 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R6252 bgr_0.V_mir2.n17 bgr_0.V_mir2.t8 120.501
R6253 bgr_0.V_mir2.n6 bgr_0.V_mir2.t18 120.501
R6254 bgr_0.V_mir2.n7 bgr_0.V_mir2.t6 120.501
R6255 bgr_0.V_mir2.n1 bgr_0.V_mir2.t17 120.501
R6256 bgr_0.V_mir2.n2 bgr_0.V_mir2.t0 120.501
R6257 bgr_0.V_mir2.n11 bgr_0.V_mir2.t12 48.0005
R6258 bgr_0.V_mir2.n11 bgr_0.V_mir2.t16 48.0005
R6259 bgr_0.V_mir2.n10 bgr_0.V_mir2.t14 48.0005
R6260 bgr_0.V_mir2.n10 bgr_0.V_mir2.t15 48.0005
R6261 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6262 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 40.7027
R6263 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 40.7027
R6264 bgr_0.V_mir2.n5 bgr_0.V_mir2.t7 39.4005
R6265 bgr_0.V_mir2.n5 bgr_0.V_mir2.t3 39.4005
R6266 bgr_0.V_mir2.n0 bgr_0.V_mir2.t1 39.4005
R6267 bgr_0.V_mir2.n0 bgr_0.V_mir2.t5 39.4005
R6268 bgr_0.V_mir2.n20 bgr_0.V_mir2.t9 39.4005
R6269 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R6270 bgr_0.V_mir2.n15 bgr_0.V_mir2.n4 15.8005
R6271 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 15.8005
R6272 bgr_0.V_mir2.n14 bgr_0.V_mir2.n9 9.3005
R6273 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 5.8755
R6274 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6275 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 0.78175
R6276 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R6277 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R6278 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t14 449.868
R6279 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t18 449.868
R6280 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.959
R6281 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R6282 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R6283 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R6284 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R6285 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R6286 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R6287 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R6288 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R6289 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R6290 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R6291 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R6292 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R6293 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R6294 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R6295 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R6296 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R6297 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R6298 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t3 184.625
R6299 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R6300 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R6301 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R6302 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R6303 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R6304 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R6305 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R6306 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R6307 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R6308 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R6309 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R6310 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R6311 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n11 170.269
R6312 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 165.8
R6313 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 73.0943
R6314 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t2 61.1914
R6315 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 56.2338
R6316 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n15 56.2338
R6317 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 56.2338
R6318 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 56.2338
R6319 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R6320 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R6321 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R6322 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R6323 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n21 17.8599
R6324 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 11.311
R6325 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 4.438
R6326 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t15 355.293
R6327 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t27 346.8
R6328 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R6329 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R6330 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n10 335.022
R6331 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t9 275.909
R6332 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n11 227.909
R6333 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.n13 222.034
R6334 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t12 184.097
R6335 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t18 184.097
R6336 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t13 184.097
R6337 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R6338 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R6339 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R6340 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R6341 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t8 48.0005
R6342 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t7 48.0005
R6343 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t6 48.0005
R6344 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t10 48.0005
R6345 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t1 39.4005
R6346 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t4 39.4005
R6347 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t0 39.4005
R6348 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t3 39.4005
R6349 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t2 39.4005
R6350 bgr_0.1st_Vout_2.t5 bgr_0.1st_Vout_2.n21 39.4005
R6351 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t16 4.8295
R6352 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t26 4.8295
R6353 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t23 4.8295
R6354 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t31 4.8295
R6355 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t14 4.8295
R6356 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t25 4.8295
R6357 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.8295
R6358 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R6359 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t11 4.5005
R6360 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t32 4.5005
R6361 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t28 4.5005
R6362 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R6363 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t36 4.5005
R6364 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t20 4.5005
R6365 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.5005
R6366 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.5005
R6367 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.5005
R6368 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R6369 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t24 4.5005
R6370 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t17 4.5005
R6371 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.n12 4.5005
R6372 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R6373 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R6374 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R6375 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R6376 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R6377 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R6378 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 0.78175
R6379 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R6380 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R6381 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R6382 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R6383 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R6384 bgr_0.cap_res2 bgr_0.cap_res2.t0 188.315
R6385 bgr_0.cap_res2 bgr_0.cap_res2.t8 0.259
R6386 bgr_0.cap_res2.t12 bgr_0.cap_res2.t17 0.1603
R6387 bgr_0.cap_res2.t3 bgr_0.cap_res2.t4 0.1603
R6388 bgr_0.cap_res2.t7 bgr_0.cap_res2.t11 0.1603
R6389 bgr_0.cap_res2.t16 bgr_0.cap_res2.t19 0.1603
R6390 bgr_0.cap_res2.t1 bgr_0.cap_res2.t6 0.1603
R6391 bgr_0.cap_res2.t9 bgr_0.cap_res2.t13 0.1603
R6392 bgr_0.cap_res2.t5 bgr_0.cap_res2.t10 0.1603
R6393 bgr_0.cap_res2.t14 bgr_0.cap_res2.t18 0.1603
R6394 bgr_0.cap_res2.n1 bgr_0.cap_res2.t20 0.159278
R6395 bgr_0.cap_res2.n2 bgr_0.cap_res2.t15 0.159278
R6396 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.159278
R6397 bgr_0.cap_res2.n3 bgr_0.cap_res2.t12 0.1368
R6398 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.1368
R6399 bgr_0.cap_res2.n2 bgr_0.cap_res2.t7 0.1368
R6400 bgr_0.cap_res2.n2 bgr_0.cap_res2.t16 0.1368
R6401 bgr_0.cap_res2.n1 bgr_0.cap_res2.t1 0.1368
R6402 bgr_0.cap_res2.n1 bgr_0.cap_res2.t9 0.1368
R6403 bgr_0.cap_res2.n0 bgr_0.cap_res2.t5 0.1368
R6404 bgr_0.cap_res2.n0 bgr_0.cap_res2.t14 0.1368
R6405 bgr_0.cap_res2.t20 bgr_0.cap_res2.n0 0.00152174
R6406 bgr_0.cap_res2.t15 bgr_0.cap_res2.n1 0.00152174
R6407 bgr_0.cap_res2.t2 bgr_0.cap_res2.n2 0.00152174
R6408 bgr_0.cap_res2.t8 bgr_0.cap_res2.n3 0.00152174
R6409 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 632.186
R6410 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6411 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6412 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 630.264
R6413 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 628.003
R6414 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 628.003
R6415 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 626.753
R6416 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 626.753
R6417 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 625.756
R6418 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 622.231
R6419 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6420 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6421 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6422 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6423 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6424 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6425 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6426 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6427 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6428 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6429 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6430 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6431 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6432 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6433 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6434 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6435 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6436 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6437 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6438 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6439 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 7.94147
R6440 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 6.188
R6441 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n22 630.264
R6442 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n24 627.316
R6443 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n26 626.784
R6444 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 626.784
R6445 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n23 626.784
R6446 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.n27 585
R6447 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6448 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6449 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n21 223.638
R6450 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6451 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.n2 176.733
R6452 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.n3 176.733
R6453 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.n4 176.733
R6454 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6455 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6456 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6457 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6458 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6459 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6460 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6461 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6462 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6463 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6464 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6465 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6466 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n20 162.214
R6467 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6468 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6469 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6470 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6471 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6472 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6473 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6474 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6475 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6476 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6477 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6478 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6479 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6480 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6481 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6482 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6483 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6484 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6485 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6486 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6487 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6488 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6489 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6490 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6491 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6492 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6493 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6494 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6495 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6496 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6497 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 49.8072
R6498 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n17 49.8072
R6499 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.n0 41.7838
R6500 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 39.8442
R6501 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t2 24.0005
R6502 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t13 24.0005
R6503 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n1 2.313
R6504 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t26 1172.87
R6505 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t35 1172.87
R6506 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.t45 996.134
R6507 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t34 996.134
R6508 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t48 996.134
R6509 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6510 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t51 996.134
R6511 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6512 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6513 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t30 996.134
R6514 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t29 690.867
R6515 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t40 690.867
R6516 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t54 530.201
R6517 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t33 530.201
R6518 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6519 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t49 514.134
R6520 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 514.134
R6521 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6522 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t31 514.134
R6523 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 514.134
R6524 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 514.134
R6525 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6526 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6527 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6528 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6529 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t42 353.467
R6530 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t28 353.467
R6531 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t44 353.467
R6532 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t32 353.467
R6533 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t47 353.467
R6534 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 176.733
R6535 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6536 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6537 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6538 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R6539 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.n47 176.733
R6540 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 176.733
R6541 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 176.733
R6542 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R6543 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6544 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6545 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6546 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 176.733
R6547 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6548 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6549 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6550 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6551 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6552 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 166.436
R6553 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n31 161.875
R6554 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 161.686
R6555 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n0 160.427
R6556 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 159.802
R6557 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 159.802
R6558 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 159.802
R6559 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n1 159.802
R6560 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 155.302
R6561 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n13 114.689
R6562 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n12 114.689
R6563 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 114.126
R6564 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 114.126
R6565 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 114.126
R6566 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n11 109.626
R6567 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 51.9494
R6568 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R6569 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 51.9494
R6570 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n23 51.9494
R6571 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R6572 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n32 51.9494
R6573 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.X.n52 49.3036
R6574 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R6575 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t13 16.0005
R6576 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R6577 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R6578 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6579 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R6580 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t18 16.0005
R6581 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t6 16.0005
R6582 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t5 16.0005
R6583 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R6584 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R6585 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R6586 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n42 15.7193
R6587 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R6588 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R6589 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t22 11.2576
R6590 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t3 11.2576
R6591 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R6592 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R6593 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t10 11.2576
R6594 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t8 11.2576
R6595 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R6596 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t11 11.2576
R6597 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t23 11.2576
R6598 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R6599 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n22 10.188
R6600 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 6.188
R6601 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n8 5.1255
R6602 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n20 4.5005
R6603 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 0.6255
R6604 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.6255
R6605 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.6255
R6606 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 0.563
R6607 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n17 0.563
R6608 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 0.563
R6609 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n10 0.5005
R6610 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 0.438
R6611 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R6612 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R6613 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R6614 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R6615 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R6616 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R6617 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R6618 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R6619 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 122.504
R6620 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 72.4688
R6621 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 60.5161
R6622 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R6623 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R6624 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R6625 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R6626 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R6627 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R6628 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 39.4005
R6629 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6630 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 19.7005
R6631 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R6632 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R6633 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R6634 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6635 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6636 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 19.7005
R6637 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6638 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R6639 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.09425
R6640 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R6641 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R6642 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R6643 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 0.09425
R6644 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t11 354.854
R6645 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t21 346.8
R6646 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R6647 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R6648 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n6 335.022
R6649 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t9 275.909
R6650 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.n7 227.909
R6651 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 222.034
R6652 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t26 184.097
R6653 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t34 184.097
R6654 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t18 184.097
R6655 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t24 184.097
R6656 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R6657 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R6658 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t7 48.0005
R6659 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t8 48.0005
R6660 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t4 48.0005
R6661 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t6 48.0005
R6662 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t2 39.4005
R6663 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t5 39.4005
R6664 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t10 39.4005
R6665 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t3 39.4005
R6666 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t1 39.4005
R6667 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t0 39.4005
R6668 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R6669 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R6670 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R6671 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t31 4.8295
R6672 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t22 4.8295
R6673 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R6674 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t30 4.8295
R6675 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.8295
R6676 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.8295
R6677 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t15 4.8295
R6678 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 4.5005
R6679 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.5005
R6680 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.5005
R6681 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R6682 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R6683 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t33 4.5005
R6684 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t36 4.5005
R6685 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t16 4.5005
R6686 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R6687 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t29 4.5005
R6688 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t12 4.5005
R6689 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.5005
R6690 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.5005
R6691 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R6692 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R6693 bgr_0.V_TOP.n0 bgr_0.V_TOP.t18 369.534
R6694 bgr_0.V_TOP.n10 bgr_0.V_TOP.n8 339.959
R6695 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R6696 bgr_0.V_TOP.n10 bgr_0.V_TOP.n9 339.272
R6697 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R6698 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6699 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 334.772
R6700 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R6701 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R6702 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R6703 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R6704 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R6705 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R6706 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R6707 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R6708 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R6709 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R6710 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R6711 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R6712 bgr_0.V_TOP bgr_0.V_TOP.t39 214.222
R6713 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R6714 bgr_0.V_TOP.n7 bgr_0.V_TOP.t13 176.114
R6715 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R6716 bgr_0.V_TOP.n27 bgr_0.V_TOP.t15 144.601
R6717 bgr_0.V_TOP.n26 bgr_0.V_TOP.t19 144.601
R6718 bgr_0.V_TOP.n25 bgr_0.V_TOP.t24 144.601
R6719 bgr_0.V_TOP.n24 bgr_0.V_TOP.t41 144.601
R6720 bgr_0.V_TOP.n23 bgr_0.V_TOP.t43 144.601
R6721 bgr_0.V_TOP.n22 bgr_0.V_TOP.t20 144.601
R6722 bgr_0.V_TOP.n21 bgr_0.V_TOP.t26 144.601
R6723 bgr_0.V_TOP.n20 bgr_0.V_TOP.t31 144.601
R6724 bgr_0.V_TOP.n0 bgr_0.V_TOP.t40 144.601
R6725 bgr_0.V_TOP.n1 bgr_0.V_TOP.t34 144.601
R6726 bgr_0.V_TOP.n2 bgr_0.V_TOP.t32 144.601
R6727 bgr_0.V_TOP.n3 bgr_0.V_TOP.t29 144.601
R6728 bgr_0.V_TOP.n4 bgr_0.V_TOP.t49 144.601
R6729 bgr_0.V_TOP.n5 bgr_0.V_TOP.t45 144.601
R6730 bgr_0.V_TOP.n18 bgr_0.V_TOP.t4 95.447
R6731 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R6732 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R6733 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R6734 bgr_0.V_TOP.n6 bgr_0.V_TOP.t2 39.4005
R6735 bgr_0.V_TOP.n6 bgr_0.V_TOP.t8 39.4005
R6736 bgr_0.V_TOP.n11 bgr_0.V_TOP.t7 39.4005
R6737 bgr_0.V_TOP.n11 bgr_0.V_TOP.t9 39.4005
R6738 bgr_0.V_TOP.n9 bgr_0.V_TOP.t11 39.4005
R6739 bgr_0.V_TOP.n9 bgr_0.V_TOP.t1 39.4005
R6740 bgr_0.V_TOP.n8 bgr_0.V_TOP.t3 39.4005
R6741 bgr_0.V_TOP.n8 bgr_0.V_TOP.t12 39.4005
R6742 bgr_0.V_TOP.n14 bgr_0.V_TOP.t5 39.4005
R6743 bgr_0.V_TOP.n14 bgr_0.V_TOP.t6 39.4005
R6744 bgr_0.V_TOP.n16 bgr_0.V_TOP.t10 39.4005
R6745 bgr_0.V_TOP.n16 bgr_0.V_TOP.t0 39.4005
R6746 bgr_0.V_TOP.n12 bgr_0.V_TOP.n10 8.313
R6747 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R6748 bgr_0.V_TOP.n28 bgr_0.V_TOP.t37 4.8295
R6749 bgr_0.V_TOP.n29 bgr_0.V_TOP.t48 4.8295
R6750 bgr_0.V_TOP.n31 bgr_0.V_TOP.t44 4.8295
R6751 bgr_0.V_TOP.n32 bgr_0.V_TOP.t22 4.8295
R6752 bgr_0.V_TOP.n34 bgr_0.V_TOP.t35 4.8295
R6753 bgr_0.V_TOP.n35 bgr_0.V_TOP.t47 4.8295
R6754 bgr_0.V_TOP.n37 bgr_0.V_TOP.t25 4.8295
R6755 bgr_0.V_TOP.n28 bgr_0.V_TOP.t30 4.5005
R6756 bgr_0.V_TOP.n30 bgr_0.V_TOP.t17 4.5005
R6757 bgr_0.V_TOP.n29 bgr_0.V_TOP.t23 4.5005
R6758 bgr_0.V_TOP.n31 bgr_0.V_TOP.t36 4.5005
R6759 bgr_0.V_TOP.n33 bgr_0.V_TOP.t28 4.5005
R6760 bgr_0.V_TOP.n32 bgr_0.V_TOP.t33 4.5005
R6761 bgr_0.V_TOP.n34 bgr_0.V_TOP.t27 4.5005
R6762 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R6763 bgr_0.V_TOP.n35 bgr_0.V_TOP.t21 4.5005
R6764 bgr_0.V_TOP.n37 bgr_0.V_TOP.t14 4.5005
R6765 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R6766 bgr_0.V_TOP.n39 bgr_0.V_TOP.t46 4.5005
R6767 bgr_0.V_TOP.n40 bgr_0.V_TOP.t38 4.5005
R6768 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R6769 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R6770 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R6771 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R6772 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R6773 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R6774 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R6775 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R6776 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R6777 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R6778 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R6779 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R6780 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R6781 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R6782 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R6783 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R6784 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t52 1172.87
R6785 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t27 1172.87
R6786 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t44 996.134
R6787 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6788 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R6789 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R6790 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6791 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R6792 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t42 996.134
R6793 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t29 996.134
R6794 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R6795 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t30 690.867
R6796 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t51 530.201
R6797 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t26 530.201
R6798 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t39 514.134
R6799 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t53 514.134
R6800 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R6801 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R6802 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t38 514.134
R6803 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t50 514.134
R6804 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R6805 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 514.134
R6806 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t34 353.467
R6807 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R6808 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t28 353.467
R6809 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t43 353.467
R6810 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R6811 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R6812 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R6813 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t46 353.467
R6814 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6815 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6816 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6817 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6818 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6819 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 176.733
R6820 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R6821 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6822 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6823 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6824 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6825 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6826 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R6827 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6828 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6829 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6830 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6831 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6832 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 166.375
R6833 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.875
R6834 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.686
R6835 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n0 160.427
R6836 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 159.802
R6837 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 159.802
R6838 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 159.802
R6839 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n1 159.802
R6840 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 155.302
R6841 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 114.689
R6842 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n12 114.689
R6843 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 114.126
R6844 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 114.126
R6845 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 114.126
R6846 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n11 109.626
R6847 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6848 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n42 51.9494
R6849 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6850 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R6851 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6852 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R6853 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t22 49.2412
R6854 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t18 16.0005
R6855 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R6856 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t16 16.0005
R6857 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t14 16.0005
R6858 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R6859 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t13 16.0005
R6860 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R6861 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6862 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R6863 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t17 16.0005
R6864 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R6865 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t19 16.0005
R6866 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 15.6567
R6867 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t8 11.2576
R6868 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t21 11.2576
R6869 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t3 11.2576
R6870 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t0 11.2576
R6871 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R6872 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R6873 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t9 11.2576
R6874 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t6 11.2576
R6875 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R6876 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t2 11.2576
R6877 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t24 11.2576
R6878 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t1 11.2576
R6879 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n51 10.313
R6880 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n40 6.063
R6881 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n8 5.1255
R6882 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 4.5005
R6883 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 0.6255
R6884 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.6255
R6885 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.6255
R6886 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n14 0.563
R6887 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n16 0.563
R6888 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n18 0.563
R6889 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n10 0.5005
R6890 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n21 0.438
R6891 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 144.827
R6892 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R6893 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 120.629
R6894 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 97.4009
R6895 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 96.8384
R6896 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 96.8384
R6897 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 96.8384
R6898 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 96.8384
R6899 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 53.2193
R6900 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 24.0005
R6901 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R6902 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 24.0005
R6903 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R6904 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 8.0005
R6905 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R6906 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 8.0005
R6907 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R6908 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R6909 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R6910 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R6911 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R6912 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R6913 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 8.0005
R6914 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 5.84425
R6915 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 1.438
R6916 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.563
R6917 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.563
R6918 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R6919 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n0 145.989
R6920 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n7 145.989
R6921 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n5 145.427
R6922 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n3 145.427
R6923 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n1 145.427
R6924 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n9 140.927
R6925 two_stage_opamp_dummy_magic_0.VOUT+.t0 two_stage_opamp_dummy_magic_0.VOUT+.n100 113.192
R6926 two_stage_opamp_dummy_magic_0.VOUT+.n97 two_stage_opamp_dummy_magic_0.VOUT+.n95 95.7303
R6927 two_stage_opamp_dummy_magic_0.VOUT+.n99 two_stage_opamp_dummy_magic_0.VOUT+.n98 94.6053
R6928 two_stage_opamp_dummy_magic_0.VOUT+.n97 two_stage_opamp_dummy_magic_0.VOUT+.n96 94.6053
R6929 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.n10 20.5943
R6930 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.n93 11.7059
R6931 two_stage_opamp_dummy_magic_0.VOUT+.n100 two_stage_opamp_dummy_magic_0.VOUT+.n94 10.6567
R6932 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t10 6.56717
R6933 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t14 6.56717
R6934 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t8 6.56717
R6935 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t2 6.56717
R6936 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t9 6.56717
R6937 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t13 6.56717
R6938 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t11 6.56717
R6939 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t15 6.56717
R6940 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t12 6.56717
R6941 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t16 6.56717
R6942 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t1 6.56717
R6943 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t17 6.56717
R6944 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t108 4.8295
R6945 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t25 4.8295
R6946 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t76 4.8295
R6947 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t113 4.8295
R6948 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.t145 4.8295
R6949 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t68 4.8295
R6950 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t28 4.8295
R6951 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t77 4.8295
R6952 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t63 4.8295
R6953 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t111 4.8295
R6954 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t114 4.8295
R6955 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t99 4.8295
R6956 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t74 4.8295
R6957 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t56 4.8295
R6958 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t109 4.8295
R6959 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t92 4.8295
R6960 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t69 4.8295
R6961 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t53 4.8295
R6962 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t30 4.8295
R6963 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t153 4.8295
R6964 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.t64 4.8295
R6965 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t47 4.8295
R6966 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t117 4.8295
R6967 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t72 4.8295
R6968 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t38 4.8295
R6969 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t20 4.8295
R6970 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t80 4.8295
R6971 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t61 4.8295
R6972 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t121 4.8295
R6973 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t104 4.8295
R6974 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t85 4.8295
R6975 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t67 4.8295
R6976 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t123 4.8295
R6977 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.t107 4.8295
R6978 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.t22 4.8295
R6979 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t33 4.806
R6980 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t150 4.806
R6981 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t51 4.806
R6982 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t88 4.806
R6983 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t125 4.806
R6984 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t105 4.806
R6985 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t140 4.806
R6986 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t37 4.806
R6987 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t156 4.806
R6988 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t54 4.806
R6989 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t73 4.806
R6990 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t116 4.806
R6991 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t65 4.806
R6992 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t154 4.806
R6993 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t106 4.806
R6994 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t143 4.806
R6995 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t96 4.806
R6996 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t43 4.806
R6997 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t87 4.806
R6998 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t35 4.806
R6999 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t70 4.5005
R7000 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.t91 4.5005
R7001 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t66 4.5005
R7002 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t81 4.5005
R7003 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t44 4.5005
R7004 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t118 4.5005
R7005 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t57 4.5005
R7006 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t21 4.5005
R7007 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t151 4.5005
R7008 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.t98 4.5005
R7009 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t60 4.5005
R7010 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.t45 4.5005
R7011 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t136 4.5005
R7012 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.t101 4.5005
R7013 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t31 4.5005
R7014 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t52 4.5005
R7015 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t155 4.5005
R7016 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t119 4.5005
R7017 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t139 4.5005
R7018 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t102 4.5005
R7019 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t62 4.5005
R7020 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t86 4.5005
R7021 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t46 4.5005
R7022 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t147 4.5005
R7023 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t110 4.5005
R7024 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t134 4.5005
R7025 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t130 4.5005
R7026 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t152 4.5005
R7027 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t115 4.5005
R7028 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t23 4.5005
R7029 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t48 4.5005
R7030 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t148 4.5005
R7031 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t79 4.5005
R7032 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t27 4.5005
R7033 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t132 4.5005
R7034 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t40 4.5005
R7035 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t128 4.5005
R7036 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t93 4.5005
R7037 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t71 4.5005
R7038 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t19 4.5005
R7039 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t126 4.5005
R7040 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t34 4.5005
R7041 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t122 4.5005
R7042 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t89 4.5005
R7043 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t135 4.5005
R7044 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t83 4.5005
R7045 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t49 4.5005
R7046 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.t29 4.5005
R7047 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.t120 4.5005
R7048 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t82 4.5005
R7049 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t26 4.5005
R7050 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.t124 4.5005
R7051 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t39 4.5005
R7052 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.t127 4.5005
R7053 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t95 4.5005
R7054 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t55 4.5005
R7055 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t144 4.5005
R7056 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t112 4.5005
R7057 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t75 4.5005
R7058 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t24 4.5005
R7059 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t131 4.5005
R7060 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t97 4.5005
R7061 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t59 4.5005
R7062 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t149 4.5005
R7063 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t142 4.5005
R7064 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.t94 4.5005
R7065 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t58 4.5005
R7066 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t42 4.5005
R7067 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.t133 4.5005
R7068 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t100 4.5005
R7069 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t84 4.5005
R7070 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.t32 4.5005
R7071 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t137 4.5005
R7072 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t50 4.5005
R7073 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.t138 4.5005
R7074 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t103 4.5005
R7075 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t90 4.5005
R7076 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t36 4.5005
R7077 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.t141 4.5005
R7078 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.t129 4.5005
R7079 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t78 4.5005
R7080 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t41 4.5005
R7081 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.t146 4.5005
R7082 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n8 4.5005
R7083 two_stage_opamp_dummy_magic_0.VOUT+.n98 two_stage_opamp_dummy_magic_0.VOUT+.t7 3.42907
R7084 two_stage_opamp_dummy_magic_0.VOUT+.n98 two_stage_opamp_dummy_magic_0.VOUT+.t4 3.42907
R7085 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.t3 3.42907
R7086 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.t18 3.42907
R7087 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.t5 3.42907
R7088 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.t6 3.42907
R7089 two_stage_opamp_dummy_magic_0.VOUT+.n100 two_stage_opamp_dummy_magic_0.VOUT+.n99 2.03175
R7090 two_stage_opamp_dummy_magic_0.VOUT+.n99 two_stage_opamp_dummy_magic_0.VOUT+.n97 1.1255
R7091 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n2 0.563
R7092 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n4 0.563
R7093 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n6 0.563
R7094 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n40 0.3295
R7095 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n53 0.3295
R7096 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n52 0.3295
R7097 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.n50 0.3295
R7098 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.n49 0.3295
R7099 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.n47 0.3295
R7100 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.n46 0.3295
R7101 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.n44 0.3295
R7102 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.n43 0.3295
R7103 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.n42 0.3295
R7104 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.n64 0.3295
R7105 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n63 0.3295
R7106 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.n62 0.3295
R7107 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.n61 0.3295
R7108 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n60 0.3295
R7109 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.n59 0.3295
R7110 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.n58 0.3295
R7111 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n57 0.3295
R7112 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.n56 0.3295
R7113 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.n55 0.3295
R7114 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.n66 0.3295
R7115 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.n67 0.3295
R7116 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.n69 0.3295
R7117 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.n70 0.3295
R7118 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.n72 0.3295
R7119 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.n73 0.3295
R7120 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.n75 0.3295
R7121 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.n76 0.3295
R7122 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.n78 0.3295
R7123 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.n79 0.3295
R7124 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.n81 0.3295
R7125 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.n82 0.3295
R7126 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.n84 0.3295
R7127 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.n85 0.3295
R7128 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.n87 0.3295
R7129 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.n88 0.3295
R7130 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.n11 0.3295
R7131 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n13 0.3295
R7132 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n23 0.3295
R7133 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.n22 0.3295
R7134 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.n21 0.3295
R7135 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.n20 0.3295
R7136 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.n19 0.3295
R7137 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.n18 0.3295
R7138 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.n17 0.3295
R7139 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.n16 0.3295
R7140 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.n15 0.3295
R7141 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.n14 0.3295
R7142 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n25 0.3295
R7143 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n26 0.3295
R7144 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n28 0.3295
R7145 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n29 0.3295
R7146 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n31 0.3295
R7147 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n32 0.3295
R7148 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n34 0.3295
R7149 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n35 0.3295
R7150 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.n37 0.3295
R7151 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.n38 0.3295
R7152 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.n90 0.3295
R7153 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.n91 0.3295
R7154 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n92 0.3295
R7155 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.n54 0.306
R7156 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.n51 0.306
R7157 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n48 0.306
R7158 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.n45 0.306
R7159 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.n41 0.2825
R7160 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.n65 0.2825
R7161 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.n68 0.2825
R7162 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.n71 0.2825
R7163 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.n74 0.2825
R7164 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.n77 0.2825
R7165 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.n80 0.2825
R7166 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.n83 0.2825
R7167 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.n86 0.2825
R7168 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n12 0.2825
R7169 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n24 0.2825
R7170 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n27 0.2825
R7171 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n30 0.2825
R7172 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n33 0.2825
R7173 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.n36 0.2825
R7174 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.n39 0.2825
R7175 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.n89 0.2825
R7176 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 49.2006
R7177 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1603
R7178 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R7179 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R7180 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R7181 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.1603
R7182 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R7183 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1603
R7184 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R7185 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R7186 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7187 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R7188 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1603
R7189 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.1603
R7190 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R7191 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7192 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R7193 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R7194 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7195 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R7196 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7197 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1603
R7198 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R7199 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R7200 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1603
R7201 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.1603
R7202 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7203 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7204 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7205 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7206 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R7207 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7208 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R7209 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R7210 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1603
R7211 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R7212 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1603
R7213 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R7214 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1603
R7215 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7216 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R7217 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7218 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7219 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R7220 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R7221 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R7222 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R7223 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.1603
R7224 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R7225 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R7226 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7227 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R7228 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R7229 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R7230 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R7231 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7232 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R7233 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.1603
R7234 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1603
R7235 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.159278
R7236 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.159278
R7237 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.159278
R7238 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.159278
R7239 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.159278
R7240 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.159278
R7241 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.159278
R7242 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7243 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7244 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7245 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7246 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7247 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7248 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7249 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7250 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7251 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7252 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7253 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7254 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7255 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7256 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7257 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7258 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.159278
R7259 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R7260 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.159278
R7261 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.159278
R7262 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.137822
R7263 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1368
R7264 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1368
R7265 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7266 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R7267 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1368
R7268 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1368
R7269 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1368
R7270 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1368
R7271 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7272 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1368
R7273 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1368
R7274 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R7275 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1368
R7276 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1368
R7277 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R7278 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1368
R7279 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1368
R7280 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7281 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1368
R7282 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R7283 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R7284 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1368
R7285 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1368
R7286 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1368
R7287 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1368
R7288 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R7289 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1368
R7290 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1368
R7291 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7292 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R7293 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1368
R7294 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.114322
R7295 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7296 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7297 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7298 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7299 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7300 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7301 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7302 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7303 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7304 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7305 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7306 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7307 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7308 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7309 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7310 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7311 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7312 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7313 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7314 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7315 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.00152174
R7316 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.00152174
R7317 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.00152174
R7318 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.00152174
R7319 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.00152174
R7320 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.00152174
R7321 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R7322 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.00152174
R7323 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.00152174
R7324 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R7325 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R7326 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.00152174
R7327 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.00152174
R7328 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.00152174
R7329 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R7330 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.00152174
R7331 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R7332 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.00152174
R7333 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.00152174
R7334 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R7335 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.00152174
R7336 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.00152174
R7337 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7338 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.00152174
R7339 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.00152174
R7340 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.00152174
R7341 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7342 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.00152174
R7343 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.00152174
R7344 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.00152174
R7345 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.00152174
R7346 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.00152174
R7347 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R7348 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7349 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7350 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 525.38
R7351 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 525.38
R7352 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 366.856
R7353 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 366.856
R7354 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7355 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 281.168
R7356 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7357 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R7358 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7359 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7360 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7361 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7362 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7363 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7364 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7365 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7366 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 39.5005
R7367 a_5750_2946.t0 a_5750_2946.t1 169.905
R7368 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7369 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7370 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7371 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7372 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t6 660.109
R7373 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t3 660.109
R7374 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n14 428.8
R7375 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n15 428.8
R7376 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.VD3.n16 239.915
R7377 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.n17 239.915
R7378 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n19 230.4
R7379 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 230.4
R7380 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n14 198.4
R7381 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n15 198.4
R7382 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n11 160.428
R7383 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 160.427
R7384 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.427
R7385 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 160.053
R7386 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 159.803
R7387 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 159.803
R7388 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 159.802
R7389 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 159.802
R7390 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.802
R7391 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 155.302
R7392 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t5 155.125
R7393 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t8 155.125
R7394 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 146.002
R7395 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.t7 98.2764
R7396 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.VD3.t36 98.2764
R7397 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t31 98.2764
R7398 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t16 98.2764
R7399 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.t10 98.2764
R7400 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.VD3.t21 98.2764
R7401 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.VD3.t12 98.2764
R7402 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t27 98.2764
R7403 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t33 98.2764
R7404 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t4 98.2764
R7405 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.n14 92.5005
R7406 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n25 92.5005
R7407 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 92.5005
R7408 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 92.5005
R7409 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 92.5005
R7410 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n23 92.5005
R7411 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t19 49.1384
R7412 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t24 49.1384
R7413 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 21.3338
R7414 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 21.3338
R7415 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n26 19.2005
R7416 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 13.8005
R7417 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R7418 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R7419 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R7420 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R7421 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R7422 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R7423 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R7424 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t14 11.2576
R7425 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R7426 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R7427 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R7428 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R7429 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R7430 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R7431 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t28 11.2576
R7432 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t34 11.2576
R7433 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R7434 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R7435 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R7436 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t32 11.2576
R7437 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R7438 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R7439 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 5.40675
R7440 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n8 4.5005
R7441 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n10 0.78175
R7442 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7443 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7444 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.6255
R7445 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.6255
R7446 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n13 0.6255
R7447 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.2505
R7448 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 628.034
R7449 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 626.784
R7450 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 626.784
R7451 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 289.2
R7452 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 289.2
R7453 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 228.252
R7454 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 212.733
R7455 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 212.733
R7456 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R7457 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R7458 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R7459 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 176.733
R7460 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 176.733
R7461 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 152
R7462 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 152
R7463 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R7464 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R7465 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 112.468
R7466 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 112.468
R7467 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R7468 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R7469 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 112.468
R7470 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 112.468
R7471 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R7472 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 78.8005
R7473 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 78.8005
R7474 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R7475 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 78.8005
R7476 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R7477 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 48.0005
R7478 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 48.0005
R7479 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 48.0005
R7480 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 48.0005
R7481 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R7482 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R7483 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R7484 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 45.5227
R7485 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R7486 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R7487 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 33.8443
R7488 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 14.2693
R7489 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 14.2693
R7490 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 1.2505
R7491 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 1.2505
R7492 bgr_0.START_UP.n3 bgr_0.START_UP.t6 238.322
R7493 bgr_0.START_UP.n3 bgr_0.START_UP.t7 238.322
R7494 bgr_0.START_UP.n2 bgr_0.START_UP.n0 175.56
R7495 bgr_0.START_UP.n2 bgr_0.START_UP.n1 168.935
R7496 bgr_0.START_UP.n4 bgr_0.START_UP.n3 166.925
R7497 bgr_0.START_UP.n5 bgr_0.START_UP.t5 130.001
R7498 bgr_0.START_UP.n5 bgr_0.START_UP.t4 81.7084
R7499 bgr_0.START_UP bgr_0.START_UP.n5 38.2614
R7500 bgr_0.START_UP bgr_0.START_UP.n4 14.7817
R7501 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R7502 bgr_0.START_UP.n1 bgr_0.START_UP.t1 13.1338
R7503 bgr_0.START_UP.n0 bgr_0.START_UP.t2 13.1338
R7504 bgr_0.START_UP.n0 bgr_0.START_UP.t3 13.1338
R7505 bgr_0.START_UP.n4 bgr_0.START_UP.n2 4.21925
R7506 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t16 623.701
R7507 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t23 611.739
R7508 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R7509 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t17 611.739
R7510 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t26 611.739
R7511 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R7512 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R7513 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R7514 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R7515 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R7516 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R7517 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R7518 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R7519 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R7520 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t20 421.75
R7521 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t25 421.75
R7522 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t12 421.75
R7523 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R7524 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R7525 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R7526 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R7527 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 172.667
R7528 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n13 172.436
R7529 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R7530 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R7531 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R7532 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R7533 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R7534 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R7535 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R7536 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R7537 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R7538 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R7539 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R7540 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R7541 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 166.25
R7542 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n1 139.638
R7543 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n0 139.638
R7544 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 134.577
R7545 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 84.4536
R7546 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 47.1294
R7547 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n17 47.1294
R7548 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 47.1294
R7549 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n8 47.1294
R7550 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 27.9067
R7551 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R7552 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R7553 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R7554 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R7555 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R7556 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R7557 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t4 10.9449
R7558 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R7559 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n2 4.5005
R7560 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n24 4.29738
R7561 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 1.2505
R7562 bgr_0.cap_res1.t20 bgr_0.cap_res1.t17 178.633
R7563 bgr_0.cap_res1.t14 bgr_0.cap_res1.t18 0.1603
R7564 bgr_0.cap_res1.t19 bgr_0.cap_res1.t16 0.1603
R7565 bgr_0.cap_res1.t6 bgr_0.cap_res1.t13 0.1603
R7566 bgr_0.cap_res1.t15 bgr_0.cap_res1.t8 0.1603
R7567 bgr_0.cap_res1.t0 bgr_0.cap_res1.t5 0.1603
R7568 bgr_0.cap_res1.t7 bgr_0.cap_res1.t1 0.1603
R7569 bgr_0.cap_res1.t3 bgr_0.cap_res1.t11 0.1603
R7570 bgr_0.cap_res1.t12 bgr_0.cap_res1.t4 0.1603
R7571 bgr_0.cap_res1.n1 bgr_0.cap_res1.t9 0.159278
R7572 bgr_0.cap_res1.n2 bgr_0.cap_res1.t2 0.159278
R7573 bgr_0.cap_res1.n3 bgr_0.cap_res1.t10 0.159278
R7574 bgr_0.cap_res1.n3 bgr_0.cap_res1.t14 0.1368
R7575 bgr_0.cap_res1.n3 bgr_0.cap_res1.t19 0.1368
R7576 bgr_0.cap_res1.n2 bgr_0.cap_res1.t6 0.1368
R7577 bgr_0.cap_res1.n2 bgr_0.cap_res1.t15 0.1368
R7578 bgr_0.cap_res1.n1 bgr_0.cap_res1.t0 0.1368
R7579 bgr_0.cap_res1.n1 bgr_0.cap_res1.t7 0.1368
R7580 bgr_0.cap_res1.n0 bgr_0.cap_res1.t3 0.1368
R7581 bgr_0.cap_res1.n0 bgr_0.cap_res1.t12 0.1368
R7582 bgr_0.cap_res1.t9 bgr_0.cap_res1.n0 0.00152174
R7583 bgr_0.cap_res1.t2 bgr_0.cap_res1.n1 0.00152174
R7584 bgr_0.cap_res1.t10 bgr_0.cap_res1.n2 0.00152174
R7585 bgr_0.cap_res1.t17 bgr_0.cap_res1.n3 0.00152174
R7586 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n7 114.719
R7587 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7588 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 114.156
R7589 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7590 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7591 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7592 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7593 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7594 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7595 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7596 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7597 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7598 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7599 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7600 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7601 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7602 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7603 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7604 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7605 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7606 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7607 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7608 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7609 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7610 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7611 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7612 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7613 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7614 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7615 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7616 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7617 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7618 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7619 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7620 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7621 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7622 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7623 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7624 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7625 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 0.563
R7626 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7627 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7628 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7629 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7630 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7631 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7632 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7633 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7634 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7635 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7636 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7637 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7638 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7639 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7640 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7641 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7642 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7643 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7644 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7645 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7646 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7647 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7648 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7649 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7650 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7651 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7652 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7653 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7654 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7655 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7656 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7657 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7658 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7659 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7660 two_stage_opamp_dummy_magic_0.V_err_p.t12 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7661 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7662 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7663 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.3272
R7664 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7665 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7666 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7667 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7668 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7669 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7670 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7671 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7672 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7673 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7674 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7675 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7676 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.n0 165.8
R7677 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7678 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7679 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7680 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7681 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7682 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7683 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t1 117.591
R7684 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R7685 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t2 108.424
R7686 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R7687 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 42.6121
R7688 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 21.2996
R7689 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n8 17.0005
R7690 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 3.31612
R7691 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 1.26612
R7692 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.2505
R7693 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n4 1.15363
R7694 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R7695 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R7696 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t5 303.259
R7697 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R7698 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R7699 bgr_0.V_CUR_REF_REG.t2 bgr_0.V_CUR_REF_REG.n5 245.284
R7700 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 174.726
R7701 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t7 174.726
R7702 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R7703 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R7704 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R7705 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t1 39.4005
R7706 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t0 39.4005
R7707 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t40 202.595
R7708 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n9 118.168
R7709 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.n2 117.831
R7710 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n16 117.269
R7711 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.n14 117.269
R7712 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.n12 117.269
R7713 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n10 117.269
R7714 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.n7 117.269
R7715 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.n5 117.269
R7716 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.n3 117.269
R7717 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.n1 113.136
R7718 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.n0 101.335
R7719 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.n29 99.647
R7720 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 99.0857
R7721 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n32 99.0845
R7722 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.n30 99.0845
R7723 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n27 99.0845
R7724 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.n25 99.0845
R7725 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.n23 99.0845
R7726 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n34 94.5845
R7727 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 94.5845
R7728 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.t30 16.0005
R7729 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.t8 16.0005
R7730 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t3 16.0005
R7731 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t35 16.0005
R7732 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t36 16.0005
R7733 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t7 16.0005
R7734 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t1 16.0005
R7735 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t33 16.0005
R7736 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t28 16.0005
R7737 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t5 16.0005
R7738 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.t2 16.0005
R7739 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.t34 16.0005
R7740 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.t37 16.0005
R7741 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.t4 16.0005
R7742 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t0 16.0005
R7743 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t32 16.0005
R7744 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.t31 16.0005
R7745 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.t9 16.0005
R7746 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t29 16.0005
R7747 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t6 16.0005
R7748 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.t26 9.6005
R7749 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.t15 9.6005
R7750 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.t24 9.6005
R7751 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.t13 9.6005
R7752 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.t22 9.6005
R7753 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.t11 9.6005
R7754 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t20 9.6005
R7755 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t18 9.6005
R7756 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t10 9.6005
R7757 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t19 9.6005
R7758 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.t12 9.6005
R7759 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.t21 9.6005
R7760 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.t14 9.6005
R7761 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.t23 9.6005
R7762 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t16 9.6005
R7763 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t25 9.6005
R7764 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t39 9.6005
R7765 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t38 9.6005
R7766 two_stage_opamp_dummy_magic_0.V_p.t27 two_stage_opamp_dummy_magic_0.V_p.n38 9.6005
R7767 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t17 9.6005
R7768 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 4.5005
R7769 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.n18 4.5005
R7770 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.n21 4.5005
R7771 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n17 3.65675
R7772 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n19 1.28175
R7773 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n31 0.563
R7774 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n33 0.563
R7775 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 0.563
R7776 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.n11 0.563
R7777 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.n13 0.563
R7778 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n15 0.563
R7779 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.n4 0.563
R7780 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.n6 0.563
R7781 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.n22 0.563
R7782 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.n24 0.563
R7783 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n26 0.563
R7784 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n28 0.563
R7785 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n8 0.53175
R7786 bgr_0.V_mir1.n4 bgr_0.V_mir1.n0 325.473
R7787 bgr_0.V_mir1.n9 bgr_0.V_mir1.n5 325.471
R7788 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.471
R7789 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R7790 bgr_0.V_mir1.n6 bgr_0.V_mir1.t22 310.488
R7791 bgr_0.V_mir1.n1 bgr_0.V_mir1.t21 310.488
R7792 bgr_0.V_mir1.n12 bgr_0.V_mir1.t16 278.312
R7793 bgr_0.V_mir1.n12 bgr_0.V_mir1.n11 228.939
R7794 bgr_0.V_mir1.n13 bgr_0.V_mir1.n10 224.439
R7795 bgr_0.V_mir1.n18 bgr_0.V_mir1.t14 184.097
R7796 bgr_0.V_mir1.n8 bgr_0.V_mir1.t4 184.097
R7797 bgr_0.V_mir1.n3 bgr_0.V_mir1.t6 184.097
R7798 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7799 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 167.094
R7800 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 167.094
R7801 bgr_0.V_mir1.n9 bgr_0.V_mir1.n8 152
R7802 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 152
R7803 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7804 bgr_0.V_mir1.n16 bgr_0.V_mir1.t20 120.501
R7805 bgr_0.V_mir1.n17 bgr_0.V_mir1.t8 120.501
R7806 bgr_0.V_mir1.n6 bgr_0.V_mir1.t18 120.501
R7807 bgr_0.V_mir1.n7 bgr_0.V_mir1.t10 120.501
R7808 bgr_0.V_mir1.n1 bgr_0.V_mir1.t17 120.501
R7809 bgr_0.V_mir1.n2 bgr_0.V_mir1.t12 120.501
R7810 bgr_0.V_mir1.n11 bgr_0.V_mir1.t1 48.0005
R7811 bgr_0.V_mir1.n11 bgr_0.V_mir1.t3 48.0005
R7812 bgr_0.V_mir1.n10 bgr_0.V_mir1.t2 48.0005
R7813 bgr_0.V_mir1.n10 bgr_0.V_mir1.t0 48.0005
R7814 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7815 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 40.7027
R7816 bgr_0.V_mir1.n3 bgr_0.V_mir1.n2 40.7027
R7817 bgr_0.V_mir1.n5 bgr_0.V_mir1.t5 39.4005
R7818 bgr_0.V_mir1.n5 bgr_0.V_mir1.t11 39.4005
R7819 bgr_0.V_mir1.n0 bgr_0.V_mir1.t7 39.4005
R7820 bgr_0.V_mir1.n0 bgr_0.V_mir1.t13 39.4005
R7821 bgr_0.V_mir1.t15 bgr_0.V_mir1.n20 39.4005
R7822 bgr_0.V_mir1.n20 bgr_0.V_mir1.t9 39.4005
R7823 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7824 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7825 bgr_0.V_mir1.n14 bgr_0.V_mir1.n9 9.3005
R7826 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 5.8755
R7827 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7828 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 0.78175
R7829 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t2 384.967
R7830 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t6 369.534
R7831 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t7 369.534
R7832 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.t22 369.534
R7833 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 369.534
R7834 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t13 369.534
R7835 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.n19 369.534
R7836 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n0 365.491
R7837 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t16 192.8
R7838 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t21 192.8
R7839 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.t10 192.8
R7840 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t18 192.8
R7841 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.t11 192.8
R7842 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t5 192.8
R7843 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R7844 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t19 192.8
R7845 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t23 192.8
R7846 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t12 192.8
R7847 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t20 192.8
R7848 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t9 192.8
R7849 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t17 192.8
R7850 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t14 192.8
R7851 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 176.733
R7852 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R7853 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R7854 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.n6 176.733
R7855 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.n3 176.733
R7856 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R7857 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n18 176.733
R7858 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R7859 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 169.852
R7860 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n9 169.852
R7861 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 166.133
R7862 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.n1 126.876
R7863 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 56.2338
R7864 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n10 56.2338
R7865 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.n8 56.2338
R7866 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.n7 56.2338
R7867 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n4 56.2338
R7868 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 56.2338
R7869 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t0 39.4005
R7870 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 39.4005
R7871 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 28.6755
R7872 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t1 24.0005
R7873 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t3 24.0005
R7874 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.t16 673.346
R7875 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 619.134
R7876 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t24 611.739
R7877 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t12 611.739
R7878 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t18 611.739
R7879 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t27 611.739
R7880 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t28 421.75
R7881 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R7882 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R7883 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R7884 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t31 421.75
R7885 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R7886 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R7887 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R7888 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R7889 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R7890 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R7891 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R7892 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t22 421.75
R7893 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R7894 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R7895 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R7896 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t9 288.166
R7897 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 169.125
R7898 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n15 169.125
R7899 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 167.094
R7900 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 167.094
R7901 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.n22 167.094
R7902 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R7903 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R7904 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 167.094
R7905 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R7906 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R7907 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R7908 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R7909 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R7910 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 167.094
R7911 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n3 140.546
R7912 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n0 140.546
R7913 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 139.296
R7914 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n1 139.296
R7915 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 86.188
R7916 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t0 62.5402
R7917 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t10 62.5402
R7918 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 47.1294
R7919 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n19 47.1294
R7920 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n14 47.1294
R7921 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n10 47.1294
R7922 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n25 38.7817
R7923 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R7924 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R7925 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R7926 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R7927 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t1 24.0005
R7928 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R7929 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R7930 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R7931 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 14.6443
R7932 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 7.78175
R7933 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n6 5.6255
R7934 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 3.71925
R7935 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n2 3.71925
R7936 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7937 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7938 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R7939 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R7940 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R7941 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R7942 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R7943 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R7944 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R7945 bgr_0.Vin+.t0 bgr_0.Vin+.n8 158.796
R7946 bgr_0.Vin+.n8 bgr_0.Vin+.t1 147.981
R7947 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7948 bgr_0.Vin+.n3 bgr_0.Vin+.t10 96.4005
R7949 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R7950 bgr_0.Vin+.n5 bgr_0.Vin+.t2 13.1338
R7951 bgr_0.Vin+.n5 bgr_0.Vin+.t3 13.1338
R7952 bgr_0.Vin+.n4 bgr_0.Vin+.t5 13.1338
R7953 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R7954 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R7955 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 229.562
R7956 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R7957 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R7958 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R7959 bgr_0.V_p_1.n6 bgr_0.V_p_1.n0 228.938
R7960 bgr_0.V_p_1.n0 bgr_0.V_p_1.t0 98.2282
R7961 bgr_0.V_p_1.n5 bgr_0.V_p_1.t4 48.0005
R7962 bgr_0.V_p_1.n5 bgr_0.V_p_1.t6 48.0005
R7963 bgr_0.V_p_1.n4 bgr_0.V_p_1.t7 48.0005
R7964 bgr_0.V_p_1.n4 bgr_0.V_p_1.t10 48.0005
R7965 bgr_0.V_p_1.n3 bgr_0.V_p_1.t1 48.0005
R7966 bgr_0.V_p_1.n3 bgr_0.V_p_1.t8 48.0005
R7967 bgr_0.V_p_1.n2 bgr_0.V_p_1.t5 48.0005
R7968 bgr_0.V_p_1.n2 bgr_0.V_p_1.t3 48.0005
R7969 bgr_0.V_p_1.t9 bgr_0.V_p_1.n6 48.0005
R7970 bgr_0.V_p_1.n6 bgr_0.V_p_1.t2 48.0005
R7971 bgr_0.V_p_1.n0 bgr_0.V_p_1.n1 1.8755
R7972 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 144.827
R7973 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 134.577
R7974 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 120.66
R7975 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 108.281
R7976 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 97.4009
R7977 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 96.8384
R7978 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 96.8384
R7979 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 96.8384
R7980 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 96.8384
R7981 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 24.0005
R7982 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R7983 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R7984 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 24.0005
R7985 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R7986 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R7987 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R7988 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R7989 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R7990 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R7991 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R7992 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R7993 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R7994 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R7995 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 5.813
R7996 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 1.46925
R7997 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.563
R7998 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.563
R7999 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R8000 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8001 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8002 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8003 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8004 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t12 660.109
R8005 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t15 660.109
R8006 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 428.8
R8007 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n0 428.8
R8008 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.n8 239.915
R8009 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t16 239.915
R8010 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 230.4
R8011 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n3 230.4
R8012 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R8013 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n0 198.4
R8014 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n28 160.428
R8015 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 160.427
R8016 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n14 160.427
R8017 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n13 160.053
R8018 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n29 159.803
R8019 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.803
R8020 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 159.802
R8021 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.802
R8022 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 159.802
R8023 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n23 155.302
R8024 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t14 155.125
R8025 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t17 155.125
R8026 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 146.004
R8027 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t13 98.2764
R8028 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t18 98.2764
R8029 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.VD4.t24 98.2764
R8030 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.VD4.t32 98.2764
R8031 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.VD4.t28 98.2764
R8032 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t36 98.2764
R8033 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t20 98.2764
R8034 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t26 98.2764
R8035 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.VD4.t22 98.2764
R8036 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t30 98.2764
R8037 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R8038 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.n6 92.5005
R8039 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n7 92.5005
R8040 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n0 92.5005
R8041 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8042 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8043 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t34 49.1384
R8044 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.n9 49.1384
R8045 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n4 21.3338
R8046 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.n2 21.3338
R8047 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n12 19.2005
R8048 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 13.8005
R8049 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R8050 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R8051 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R8052 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R8053 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R8054 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8055 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R8056 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8057 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8058 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8059 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8060 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R8061 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8062 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R8063 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8064 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R8065 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R8066 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R8067 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R8068 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R8069 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R8070 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.VD4.n33 11.2576
R8071 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 6.188
R8072 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n22 4.5005
R8073 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 0.6255
R8074 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n17 0.6255
R8075 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n19 0.6255
R8076 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 0.6255
R8077 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R8078 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.2505
R8079 bgr_0.Vin-.n14 bgr_0.Vin-.t8 688.859
R8080 bgr_0.Vin-.n16 bgr_0.Vin-.n15 514.134
R8081 bgr_0.Vin-.n12 bgr_0.Vin-.n11 345.116
R8082 bgr_0.Vin-.n18 bgr_0.Vin-.n17 214.713
R8083 bgr_0.Vin-.n14 bgr_0.Vin-.t11 174.726
R8084 bgr_0.Vin-.n15 bgr_0.Vin-.t12 174.726
R8085 bgr_0.Vin-.n16 bgr_0.Vin-.t9 174.726
R8086 bgr_0.Vin-.n17 bgr_0.Vin-.t10 174.726
R8087 bgr_0.Vin-.n10 bgr_0.Vin-.n8 173.029
R8088 bgr_0.Vin-.n10 bgr_0.Vin-.n9 168.654
R8089 bgr_0.Vin-.n12 bgr_0.Vin-.t0 162.921
R8090 bgr_0.Vin-.n15 bgr_0.Vin-.n14 128.534
R8091 bgr_0.Vin-.n17 bgr_0.Vin-.n16 128.534
R8092 bgr_0.Vin-.n3 bgr_0.Vin-.n0 83.5719
R8093 bgr_0.Vin-.n5 bgr_0.Vin-.n4 83.5719
R8094 bgr_0.Vin-.n3 bgr_0.Vin-.n1 73.3165
R8095 bgr_0.Vin-.t1 bgr_0.Vin-.n2 65.0299
R8096 bgr_0.Vin-.n11 bgr_0.Vin-.t6 39.4005
R8097 bgr_0.Vin-.n11 bgr_0.Vin-.t7 39.4005
R8098 bgr_0.Vin-.n4 bgr_0.Vin-.n3 26.074
R8099 bgr_0.Vin-.n19 bgr_0.Vin-.n18 17.526
R8100 bgr_0.Vin-.n9 bgr_0.Vin-.t3 13.1338
R8101 bgr_0.Vin-.n9 bgr_0.Vin-.t4 13.1338
R8102 bgr_0.Vin-.n8 bgr_0.Vin-.t2 13.1338
R8103 bgr_0.Vin-.n8 bgr_0.Vin-.t5 13.1338
R8104 bgr_0.Vin-.n18 bgr_0.Vin-.n13 12.5317
R8105 bgr_0.Vin-.n13 bgr_0.Vin-.n12 6.40675
R8106 bgr_0.Vin-.n13 bgr_0.Vin-.n10 3.8755
R8107 bgr_0.Vin-.n19 bgr_0.Vin-.n1 2.19742
R8108 bgr_0.Vin-.n5 bgr_0.Vin-.n2 1.56363
R8109 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1.5505
R8110 bgr_0.Vin-.n7 bgr_0.Vin-.n6 1.5505
R8111 bgr_0.Vin-.n21 bgr_0.Vin-.n1 1.19225
R8112 bgr_0.Vin-.n6 bgr_0.Vin-.n0 0.885803
R8113 bgr_0.Vin-.n6 bgr_0.Vin-.n5 0.77514
R8114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R8115 bgr_0.Vin-.n7 bgr_0.Vin-.n2 0.537712
R8116 bgr_0.Vin-.n4 bgr_0.Vin-.t1 0.290206
R8117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n21 0.203382
R8118 bgr_0.Vin-.n20 bgr_0.Vin-.n7 0.0183571
R8119 bgr_0.Vin-.n20 bgr_0.Vin-.n19 0.0183571
R8120 a_29640_9790.t0 a_29640_9790.t1 258.591
R8121 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 413.99
R8122 bgr_0.Vbe2.n95 bgr_0.Vbe2.t8 162.458
R8123 bgr_0.Vbe2.n146 bgr_0.Vbe2.n145 84.0884
R8124 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 83.5719
R8125 bgr_0.Vbe2.n56 bgr_0.Vbe2.n49 83.5719
R8126 bgr_0.Vbe2.n55 bgr_0.Vbe2.n54 83.5719
R8127 bgr_0.Vbe2.n128 bgr_0.Vbe2.n6 83.5719
R8128 bgr_0.Vbe2.n123 bgr_0.Vbe2.n7 83.5719
R8129 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 83.5719
R8130 bgr_0.Vbe2.n72 bgr_0.Vbe2.n71 83.5719
R8131 bgr_0.Vbe2.n70 bgr_0.Vbe2.n69 83.5719
R8132 bgr_0.Vbe2.n38 bgr_0.Vbe2.n37 83.5719
R8133 bgr_0.Vbe2.n33 bgr_0.Vbe2.n31 83.5719
R8134 bgr_0.Vbe2.n84 bgr_0.Vbe2.n30 83.5719
R8135 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 83.5719
R8136 bgr_0.Vbe2.n28 bgr_0.Vbe2.n26 83.5719
R8137 bgr_0.Vbe2.n98 bgr_0.Vbe2.n25 83.5719
R8138 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 83.5719
R8139 bgr_0.Vbe2.n23 bgr_0.Vbe2.n22 83.5719
R8140 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 83.5719
R8141 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 83.5719
R8142 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 83.5719
R8143 bgr_0.Vbe2.n143 bgr_0.Vbe2.n1 83.5719
R8144 bgr_0.Vbe2.n142 bgr_0.Vbe2.n0 83.5719
R8145 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 83.5719
R8146 bgr_0.Vbe2.n133 bgr_0.Vbe2.n4 83.5719
R8147 bgr_0.Vbe2.n57 bgr_0.Vbe2.n48 73.8495
R8148 bgr_0.Vbe2.n130 bgr_0.Vbe2.n6 73.3165
R8149 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 73.3165
R8150 bgr_0.Vbe2.n37 bgr_0.Vbe2.n36 73.3165
R8151 bgr_0.Vbe2.n91 bgr_0.Vbe2.n90 73.3165
R8152 bgr_0.Vbe2.n105 bgr_0.Vbe2.n104 73.3165
R8153 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 73.3165
R8154 bgr_0.Vbe2.n55 bgr_0.Vbe2.n50 73.19
R8155 bgr_0.Vbe2.n70 bgr_0.Vbe2.n46 73.19
R8156 bgr_0.Vbe2.n86 bgr_0.Vbe2.n30 73.19
R8157 bgr_0.Vbe2.n100 bgr_0.Vbe2.n25 73.19
R8158 bgr_0.Vbe2.n112 bgr_0.Vbe2.n13 73.19
R8159 bgr_0.Vbe2.n134 bgr_0.Vbe2.n133 73.19
R8160 bgr_0.Vbe2.n124 bgr_0.Vbe2.t6 65.0299
R8161 bgr_0.Vbe2.t3 bgr_0.Vbe2.n20 65.0299
R8162 bgr_0.Vbe2.n57 bgr_0.Vbe2.n56 26.074
R8163 bgr_0.Vbe2.n123 bgr_0.Vbe2.n6 26.074
R8164 bgr_0.Vbe2.n74 bgr_0.Vbe2.n72 26.074
R8165 bgr_0.Vbe2.n37 bgr_0.Vbe2.n33 26.074
R8166 bgr_0.Vbe2.n91 bgr_0.Vbe2.n28 26.074
R8167 bgr_0.Vbe2.n105 bgr_0.Vbe2.n23 26.074
R8168 bgr_0.Vbe2.n116 bgr_0.Vbe2.n114 26.074
R8169 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 26.074
R8170 bgr_0.Vbe2.n143 bgr_0.Vbe2.n142 26.074
R8171 bgr_0.Vbe2.n145 bgr_0.Vbe2.n143 26.074
R8172 bgr_0.Vbe2.t2 bgr_0.Vbe2.n55 25.7843
R8173 bgr_0.Vbe2.t1 bgr_0.Vbe2.n70 25.7843
R8174 bgr_0.Vbe2.t0 bgr_0.Vbe2.n30 25.7843
R8175 bgr_0.Vbe2.t5 bgr_0.Vbe2.n25 25.7843
R8176 bgr_0.Vbe2.t4 bgr_0.Vbe2.n112 25.7843
R8177 bgr_0.Vbe2.n133 bgr_0.Vbe2.t7 25.7843
R8178 bgr_0.Vbe2.n15 bgr_0.Vbe2.n11 9.3005
R8179 bgr_0.Vbe2.n15 bgr_0.Vbe2.n10 9.3005
R8180 bgr_0.Vbe2.n15 bgr_0.Vbe2.n12 9.3005
R8181 bgr_0.Vbe2.n121 bgr_0.Vbe2.n15 9.3005
R8182 bgr_0.Vbe2.n17 bgr_0.Vbe2.n11 9.3005
R8183 bgr_0.Vbe2.n17 bgr_0.Vbe2.n10 9.3005
R8184 bgr_0.Vbe2.n17 bgr_0.Vbe2.n12 9.3005
R8185 bgr_0.Vbe2.n121 bgr_0.Vbe2.n17 9.3005
R8186 bgr_0.Vbe2.n14 bgr_0.Vbe2.n11 9.3005
R8187 bgr_0.Vbe2.n14 bgr_0.Vbe2.n10 9.3005
R8188 bgr_0.Vbe2.n14 bgr_0.Vbe2.n12 9.3005
R8189 bgr_0.Vbe2.n121 bgr_0.Vbe2.n14 9.3005
R8190 bgr_0.Vbe2.n19 bgr_0.Vbe2.n11 9.3005
R8191 bgr_0.Vbe2.n19 bgr_0.Vbe2.n10 9.3005
R8192 bgr_0.Vbe2.n19 bgr_0.Vbe2.n12 9.3005
R8193 bgr_0.Vbe2.n121 bgr_0.Vbe2.n19 9.3005
R8194 bgr_0.Vbe2.n122 bgr_0.Vbe2.n11 9.3005
R8195 bgr_0.Vbe2.n122 bgr_0.Vbe2.n10 9.3005
R8196 bgr_0.Vbe2.n122 bgr_0.Vbe2.n12 9.3005
R8197 bgr_0.Vbe2.n122 bgr_0.Vbe2.n9 9.3005
R8198 bgr_0.Vbe2.n122 bgr_0.Vbe2.n121 9.3005
R8199 bgr_0.Vbe2.n120 bgr_0.Vbe2.n11 9.3005
R8200 bgr_0.Vbe2.n120 bgr_0.Vbe2.n10 9.3005
R8201 bgr_0.Vbe2.n120 bgr_0.Vbe2.n12 9.3005
R8202 bgr_0.Vbe2.n120 bgr_0.Vbe2.n9 9.3005
R8203 bgr_0.Vbe2.n121 bgr_0.Vbe2.n120 9.3005
R8204 bgr_0.Vbe2.n64 bgr_0.Vbe2.n44 9.3005
R8205 bgr_0.Vbe2.n64 bgr_0.Vbe2.n42 9.3005
R8206 bgr_0.Vbe2.n64 bgr_0.Vbe2.n45 9.3005
R8207 bgr_0.Vbe2.n79 bgr_0.Vbe2.n64 9.3005
R8208 bgr_0.Vbe2.n66 bgr_0.Vbe2.n44 9.3005
R8209 bgr_0.Vbe2.n66 bgr_0.Vbe2.n42 9.3005
R8210 bgr_0.Vbe2.n66 bgr_0.Vbe2.n45 9.3005
R8211 bgr_0.Vbe2.n79 bgr_0.Vbe2.n66 9.3005
R8212 bgr_0.Vbe2.n63 bgr_0.Vbe2.n44 9.3005
R8213 bgr_0.Vbe2.n63 bgr_0.Vbe2.n42 9.3005
R8214 bgr_0.Vbe2.n63 bgr_0.Vbe2.n45 9.3005
R8215 bgr_0.Vbe2.n79 bgr_0.Vbe2.n63 9.3005
R8216 bgr_0.Vbe2.n78 bgr_0.Vbe2.n44 9.3005
R8217 bgr_0.Vbe2.n78 bgr_0.Vbe2.n42 9.3005
R8218 bgr_0.Vbe2.n78 bgr_0.Vbe2.n45 9.3005
R8219 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 9.3005
R8220 bgr_0.Vbe2.n62 bgr_0.Vbe2.n44 9.3005
R8221 bgr_0.Vbe2.n62 bgr_0.Vbe2.n42 9.3005
R8222 bgr_0.Vbe2.n62 bgr_0.Vbe2.n45 9.3005
R8223 bgr_0.Vbe2.n62 bgr_0.Vbe2.n41 9.3005
R8224 bgr_0.Vbe2.n79 bgr_0.Vbe2.n62 9.3005
R8225 bgr_0.Vbe2.n80 bgr_0.Vbe2.n44 9.3005
R8226 bgr_0.Vbe2.n80 bgr_0.Vbe2.n42 9.3005
R8227 bgr_0.Vbe2.n80 bgr_0.Vbe2.n45 9.3005
R8228 bgr_0.Vbe2.n80 bgr_0.Vbe2.n41 9.3005
R8229 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 9.3005
R8230 bgr_0.Vbe2.n16 bgr_0.Vbe2.n9 4.64654
R8231 bgr_0.Vbe2.n118 bgr_0.Vbe2.n110 4.64654
R8232 bgr_0.Vbe2.n18 bgr_0.Vbe2.n9 4.64654
R8233 bgr_0.Vbe2.n118 bgr_0.Vbe2.n8 4.64654
R8234 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 4.64654
R8235 bgr_0.Vbe2.n65 bgr_0.Vbe2.n41 4.64654
R8236 bgr_0.Vbe2.n76 bgr_0.Vbe2.n68 4.64654
R8237 bgr_0.Vbe2.n67 bgr_0.Vbe2.n41 4.64654
R8238 bgr_0.Vbe2.n77 bgr_0.Vbe2.n76 4.64654
R8239 bgr_0.Vbe2.n76 bgr_0.Vbe2.n43 4.64654
R8240 bgr_0.Vbe2.n50 bgr_0.Vbe2.n3 2.36206
R8241 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 2.36206
R8242 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 2.36206
R8243 bgr_0.Vbe2.n134 bgr_0.Vbe2.n132 2.36206
R8244 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 2.19742
R8245 bgr_0.Vbe2.n36 bgr_0.Vbe2.n34 2.19742
R8246 bgr_0.Vbe2.n90 bgr_0.Vbe2.n88 2.19742
R8247 bgr_0.Vbe2.n104 bgr_0.Vbe2.n102 2.19742
R8248 bgr_0.Vbe2.n124 bgr_0.Vbe2.n7 1.56363
R8249 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 1.56363
R8250 bgr_0.Vbe2.n103 bgr_0.Vbe2.n21 1.5505
R8251 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 1.5505
R8252 bgr_0.Vbe2.n89 bgr_0.Vbe2.n27 1.5505
R8253 bgr_0.Vbe2.n94 bgr_0.Vbe2.n93 1.5505
R8254 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 1.5505
R8255 bgr_0.Vbe2.n99 bgr_0.Vbe2.n24 1.5505
R8256 bgr_0.Vbe2.n35 bgr_0.Vbe2.n32 1.5505
R8257 bgr_0.Vbe2.n40 bgr_0.Vbe2.n39 1.5505
R8258 bgr_0.Vbe2.n83 bgr_0.Vbe2.n82 1.5505
R8259 bgr_0.Vbe2.n85 bgr_0.Vbe2.n29 1.5505
R8260 bgr_0.Vbe2.n129 bgr_0.Vbe2.n5 1.5505
R8261 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 1.5505
R8262 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 1.5505
R8263 bgr_0.Vbe2.n53 bgr_0.Vbe2.n47 1.5505
R8264 bgr_0.Vbe2.n52 bgr_0.Vbe2.n51 1.5505
R8265 bgr_0.Vbe2.n147 bgr_0.Vbe2.n146 1.5505
R8266 bgr_0.Vbe2.n149 bgr_0.Vbe2.n148 1.5505
R8267 bgr_0.Vbe2.n139 bgr_0.Vbe2.n2 1.5505
R8268 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R8269 bgr_0.Vbe2.n136 bgr_0.Vbe2.n135 1.5505
R8270 bgr_0.Vbe2.n54 bgr_0.Vbe2.n52 1.25468
R8271 bgr_0.Vbe2.n69 bgr_0.Vbe2.n41 1.25468
R8272 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 1.25468
R8273 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 1.25468
R8274 bgr_0.Vbe2.n111 bgr_0.Vbe2.n9 1.25468
R8275 bgr_0.Vbe2.n135 bgr_0.Vbe2.n4 1.25468
R8276 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 1.19225
R8277 bgr_0.Vbe2.n75 bgr_0.Vbe2.n44 1.19225
R8278 bgr_0.Vbe2.n36 bgr_0.Vbe2.n35 1.19225
R8279 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 1.19225
R8280 bgr_0.Vbe2.n104 bgr_0.Vbe2.n103 1.19225
R8281 bgr_0.Vbe2.n117 bgr_0.Vbe2.n11 1.19225
R8282 bgr_0.Vbe2.n146 bgr_0.Vbe2.n1 1.14402
R8283 bgr_0.Vbe2.n53 bgr_0.Vbe2.n49 1.07024
R8284 bgr_0.Vbe2.n71 bgr_0.Vbe2.n45 1.07024
R8285 bgr_0.Vbe2.n83 bgr_0.Vbe2.n31 1.07024
R8286 bgr_0.Vbe2.n97 bgr_0.Vbe2.n26 1.07024
R8287 bgr_0.Vbe2.n113 bgr_0.Vbe2.n12 1.07024
R8288 bgr_0.Vbe2.n140 bgr_0.Vbe2.n138 1.07024
R8289 bgr_0.Vbe2.n52 bgr_0.Vbe2.n50 1.0237
R8290 bgr_0.Vbe2.n46 bgr_0.Vbe2.n41 1.0237
R8291 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 1.0237
R8292 bgr_0.Vbe2.n100 bgr_0.Vbe2.n99 1.0237
R8293 bgr_0.Vbe2.n13 bgr_0.Vbe2.n9 1.0237
R8294 bgr_0.Vbe2.n135 bgr_0.Vbe2.n134 1.0237
R8295 bgr_0.Vbe2.n59 bgr_0.Vbe2.n58 0.885803
R8296 bgr_0.Vbe2.n128 bgr_0.Vbe2.n127 0.885803
R8297 bgr_0.Vbe2.n73 bgr_0.Vbe2.n42 0.885803
R8298 bgr_0.Vbe2.n39 bgr_0.Vbe2.n38 0.885803
R8299 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 0.885803
R8300 bgr_0.Vbe2.n107 bgr_0.Vbe2.n106 0.885803
R8301 bgr_0.Vbe2.n115 bgr_0.Vbe2.n10 0.885803
R8302 bgr_0.Vbe2.n139 bgr_0.Vbe2.n0 0.885803
R8303 bgr_0.Vbe2.n79 bgr_0.Vbe2.n46 0.812055
R8304 bgr_0.Vbe2.n121 bgr_0.Vbe2.n13 0.812055
R8305 bgr_0.Vbe2.n59 bgr_0.Vbe2.n49 0.77514
R8306 bgr_0.Vbe2.n127 bgr_0.Vbe2.n7 0.77514
R8307 bgr_0.Vbe2.n71 bgr_0.Vbe2.n42 0.77514
R8308 bgr_0.Vbe2.n39 bgr_0.Vbe2.n31 0.77514
R8309 bgr_0.Vbe2.n93 bgr_0.Vbe2.n26 0.77514
R8310 bgr_0.Vbe2.n107 bgr_0.Vbe2.n22 0.77514
R8311 bgr_0.Vbe2.n113 bgr_0.Vbe2.n10 0.77514
R8312 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.77514
R8313 bgr_0.Vbe2.n58 bgr_0.Vbe2 0.756696
R8314 bgr_0.Vbe2 bgr_0.Vbe2.n128 0.756696
R8315 bgr_0.Vbe2.n73 bgr_0.Vbe2 0.756696
R8316 bgr_0.Vbe2.n38 bgr_0.Vbe2 0.756696
R8317 bgr_0.Vbe2.n92 bgr_0.Vbe2 0.756696
R8318 bgr_0.Vbe2.n106 bgr_0.Vbe2 0.756696
R8319 bgr_0.Vbe2.n115 bgr_0.Vbe2 0.756696
R8320 bgr_0.Vbe2 bgr_0.Vbe2.n0 0.756696
R8321 bgr_0.Vbe2.n60 bgr_0.Vbe2.n48 0.711459
R8322 bgr_0.Vbe2.n149 bgr_0.Vbe2.n1 0.701365
R8323 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 0.647417
R8324 bgr_0.Vbe2.n118 bgr_0.Vbe2.n117 0.647417
R8325 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 0.590702
R8326 bgr_0.Vbe2.n69 bgr_0.Vbe2.n45 0.590702
R8327 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 0.590702
R8328 bgr_0.Vbe2.n98 bgr_0.Vbe2.n97 0.590702
R8329 bgr_0.Vbe2.n111 bgr_0.Vbe2.n12 0.590702
R8330 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.590702
R8331 bgr_0.Vbe2 bgr_0.Vbe2.n48 0.576566
R8332 bgr_0.Vbe2.n109 bgr_0.Vbe2.n20 0.530034
R8333 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.530034
R8334 bgr_0.Vbe2.n56 bgr_0.Vbe2.t2 0.290206
R8335 bgr_0.Vbe2.t6 bgr_0.Vbe2.n123 0.290206
R8336 bgr_0.Vbe2.n72 bgr_0.Vbe2.t1 0.290206
R8337 bgr_0.Vbe2.n33 bgr_0.Vbe2.t0 0.290206
R8338 bgr_0.Vbe2.n28 bgr_0.Vbe2.t5 0.290206
R8339 bgr_0.Vbe2.n23 bgr_0.Vbe2.t3 0.290206
R8340 bgr_0.Vbe2.n114 bgr_0.Vbe2.t4 0.290206
R8341 bgr_0.Vbe2.n141 bgr_0.Vbe2.t7 0.290206
R8342 bgr_0.Vbe2.n129 bgr_0.Vbe2 0.203382
R8343 bgr_0.Vbe2 bgr_0.Vbe2.n44 0.203382
R8344 bgr_0.Vbe2.n35 bgr_0.Vbe2 0.203382
R8345 bgr_0.Vbe2.n89 bgr_0.Vbe2 0.203382
R8346 bgr_0.Vbe2.n103 bgr_0.Vbe2 0.203382
R8347 bgr_0.Vbe2 bgr_0.Vbe2.n11 0.203382
R8348 bgr_0.Vbe2 bgr_0.Vbe2.n149 0.203382
R8349 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 0.154071
R8350 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 0.154071
R8351 bgr_0.Vbe2.n132 bgr_0.Vbe2.n131 0.154071
R8352 bgr_0.Vbe2.n147 bgr_0.Vbe2.n3 0.154071
R8353 bgr_0.Vbe2.n120 bgr_0.Vbe2.n109 0.137464
R8354 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 0.137464
R8355 bgr_0.Vbe2.n125 bgr_0.Vbe2.n122 0.134964
R8356 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 0.134964
R8357 bgr_0.Vbe2.n34 bgr_0.Vbe2 0.0196071
R8358 bgr_0.Vbe2.n108 bgr_0.Vbe2.n21 0.0183571
R8359 bgr_0.Vbe2.n102 bgr_0.Vbe2.n21 0.0183571
R8360 bgr_0.Vbe2.n101 bgr_0.Vbe2.n24 0.0183571
R8361 bgr_0.Vbe2.n96 bgr_0.Vbe2.n24 0.0183571
R8362 bgr_0.Vbe2.n94 bgr_0.Vbe2.n27 0.0183571
R8363 bgr_0.Vbe2.n88 bgr_0.Vbe2.n27 0.0183571
R8364 bgr_0.Vbe2.n87 bgr_0.Vbe2.n29 0.0183571
R8365 bgr_0.Vbe2.n82 bgr_0.Vbe2.n29 0.0183571
R8366 bgr_0.Vbe2.n40 bgr_0.Vbe2.n32 0.0183571
R8367 bgr_0.Vbe2.n34 bgr_0.Vbe2.n32 0.0183571
R8368 bgr_0.Vbe2.n126 bgr_0.Vbe2.n5 0.0183571
R8369 bgr_0.Vbe2.n131 bgr_0.Vbe2.n5 0.0183571
R8370 bgr_0.Vbe2.n136 bgr_0.Vbe2.n132 0.0183571
R8371 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.0183571
R8372 bgr_0.Vbe2.n137 bgr_0.Vbe2.n2 0.0183571
R8373 bgr_0.Vbe2.n148 bgr_0.Vbe2.n2 0.0183571
R8374 bgr_0.Vbe2.n148 bgr_0.Vbe2.n147 0.0183571
R8375 bgr_0.Vbe2.n51 bgr_0.Vbe2.n3 0.0183571
R8376 bgr_0.Vbe2.n51 bgr_0.Vbe2.n47 0.0183571
R8377 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.0106786
R8378 bgr_0.Vbe2.n61 bgr_0.Vbe2.n47 0.0106786
R8379 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.00996429
R8380 bgr_0.Vbe2.n120 bgr_0.Vbe2.n119 0.00992001
R8381 bgr_0.Vbe2.n17 bgr_0.Vbe2.n16 0.00992001
R8382 bgr_0.Vbe2.n110 bgr_0.Vbe2.n14 0.00992001
R8383 bgr_0.Vbe2.n19 bgr_0.Vbe2.n18 0.00992001
R8384 bgr_0.Vbe2.n122 bgr_0.Vbe2.n8 0.00992001
R8385 bgr_0.Vbe2.n119 bgr_0.Vbe2.n15 0.00992001
R8386 bgr_0.Vbe2.n16 bgr_0.Vbe2.n15 0.00992001
R8387 bgr_0.Vbe2.n110 bgr_0.Vbe2.n17 0.00992001
R8388 bgr_0.Vbe2.n18 bgr_0.Vbe2.n14 0.00992001
R8389 bgr_0.Vbe2.n19 bgr_0.Vbe2.n8 0.00992001
R8390 bgr_0.Vbe2.n80 bgr_0.Vbe2.n43 0.00992001
R8391 bgr_0.Vbe2.n66 bgr_0.Vbe2.n65 0.00992001
R8392 bgr_0.Vbe2.n68 bgr_0.Vbe2.n63 0.00992001
R8393 bgr_0.Vbe2.n78 bgr_0.Vbe2.n67 0.00992001
R8394 bgr_0.Vbe2.n77 bgr_0.Vbe2.n62 0.00992001
R8395 bgr_0.Vbe2.n64 bgr_0.Vbe2.n43 0.00992001
R8396 bgr_0.Vbe2.n65 bgr_0.Vbe2.n64 0.00992001
R8397 bgr_0.Vbe2.n68 bgr_0.Vbe2.n66 0.00992001
R8398 bgr_0.Vbe2.n67 bgr_0.Vbe2.n63 0.00992001
R8399 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 0.00992001
R8400 bgr_0.Vbe2.n96 bgr_0.Vbe2.n95 0.00889286
R8401 bgr_0.Vbe2.n109 bgr_0.Vbe2.n108 0.00817857
R8402 bgr_0.Vbe2.n81 bgr_0.Vbe2.n40 0.00817857
R8403 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 0.00817857
R8404 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 0.00817857
R8405 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t12 650.729
R8406 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n6 630.607
R8407 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 627.128
R8408 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n10 627.128
R8409 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 227.784
R8410 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 226.534
R8411 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n3 226.534
R8412 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8413 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t11 78.8005
R8414 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t8 78.8005
R8415 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t10 78.8005
R8416 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t7 78.8005
R8417 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t9 78.8005
R8418 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t2 48.0005
R8419 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t4 48.0005
R8420 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t1 48.0005
R8421 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t3 48.0005
R8422 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8423 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R8424 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n5 21.1255
R8425 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n4 10.8755
R8426 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n7 1.3755
R8427 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.2505
R8428 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 1.2505
R8429 a_5230_5758.t0 a_5230_5758.t1 294.339
R8430 a_14520_5738.t0 a_14520_5738.t1 294.339
R8431 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8432 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8433 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8434 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8435 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 672.159
R8436 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 672.159
R8437 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8438 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8439 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8440 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8441 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8442 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8443 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8444 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 160.517
R8445 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8446 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8447 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 95.7988
R8448 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8449 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8450 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8451 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8452 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8453 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8454 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8455 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 75.9449
R8456 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 75.9449
R8457 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 47.8997
R8458 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8459 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8460 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8461 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8462 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8463 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8464 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 12.313
R8465 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 12.313
R8466 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 10.9449
R8467 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 10.9449
R8468 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8469 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8470 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 220.678
R8471 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R8472 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R8473 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R8474 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t1 9.6005
R8475 a_5350_5758.t0 a_5350_5758.t1 169.905
R8476 a_27130_9400.t0 a_27130_9400.t1 258.591
R8477 a_28738_9040.t0 a_28738_9040.t1 376.99
R8478 a_14240_2946.t0 a_14240_2946.t1 169.905
R8479 a_28738_9160.t0 a_28738_9160.t1 258.591
R8480 a_27130_9280.t0 a_27130_9280.t1 376.99
R8481 a_29700_9260.t0 a_29700_9260.t1 258.591
R8482 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
C0 VDDA bgr_0.START_UP 1.39151f
C1 two_stage_opamp_dummy_magic_0.V_err_gate bgr_0.NFET_GATE_10uA 0.134659f
C2 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47368f
C3 bgr_0.Vbe2 bgr_0.V_TOP 0.285619f
C4 m2_24450_7140# bgr_0.V_TOP 0.012f
C5 VDDA m2_23090_7140# 0.010446f
C6 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.559544f
C7 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 3.88146f
C8 bgr_0.1st_Vout_1 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.477103f
C9 bgr_0.PFET_GATE_10uA bgr_0.START_UP 0.166283f
C10 bgr_0.Vbe2 bgr_0.START_UP 0.193132f
C11 VDDA two_stage_opamp_dummy_magic_0.cap_res_X 0.720924f
C12 VDDA two_stage_opamp_dummy_magic_0.V_err_amp_ref 4.25984f
C13 VDDA two_stage_opamp_dummy_magic_0.VD3 3.78008f
C14 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.err_amp_out 0.040365f
C15 VDDA two_stage_opamp_dummy_magic_0.err_amp_out 1.00936f
C16 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.953371f
C17 bgr_0.START_UP_NFET1 bgr_0.NFET_GATE_10uA 0.308028f
C18 m2_23090_7140# bgr_0.PFET_GATE_10uA 0.012f
C19 VDDA bgr_0.START_UP_NFET1 0.135132f
C20 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.46515f
C21 bgr_0.1st_Vout_1 bgr_0.NFET_GATE_10uA 1.02268f
C22 bgr_0.Vbe2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.014154f
C23 two_stage_opamp_dummy_magic_0.VIN- two_stage_opamp_dummy_magic_0.VIN+ 0.555219f
C24 VDDA bgr_0.NFET_GATE_10uA 1.08124f
C25 VDDA bgr_0.1st_Vout_1 2.06087f
C26 bgr_0.V_TOP bgr_0.START_UP 0.815644f
C27 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.551434f
C28 VDDA two_stage_opamp_dummy_magic_0.Y 4.15025f
C29 bgr_0.PFET_GATE_10uA bgr_0.NFET_GATE_10uA 0.050552f
C30 bgr_0.1st_Vout_1 bgr_0.PFET_GATE_10uA 0.035393f
C31 bgr_0.Vbe2 bgr_0.NFET_GATE_10uA 0.021455f
C32 bgr_0.1st_Vout_1 m2_24450_7140# 0.075543f
C33 VDDA bgr_0.PFET_GATE_10uA 10.3925f
C34 VDDA bgr_0.Vbe2 0.02318f
C35 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13886f
C36 VDDA m2_24450_7140# 0.010446f
C37 bgr_0.cap_res2 bgr_0.1st_Vout_1 0.822981f
C38 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.09763f
C39 bgr_0.Vbe2 bgr_0.PFET_GATE_10uA 0.242909f
C40 VDDA bgr_0.cap_res2 0.551012f
C41 bgr_0.cap_res2 li_26520_10220# 0.020538f
C42 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C43 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.04259f
C44 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_err_gate 0.011317f
C45 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.080353f
C46 bgr_0.1st_Vout_1 bgr_0.V_TOP 0.925484f
C47 bgr_0.cap_res2 bgr_0.PFET_GATE_10uA 0.018633f
C48 li_21620_10330# bgr_0.V_TOP 0.020062f
C49 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VIN+ 0.057219f
C50 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VIN- 0.856672f
C51 bgr_0.1st_Vout_1 li_28620_10330# 0.020439f
C52 VDDA li_23020_10430# 0.021911f
C53 VDDA bgr_0.V_TOP 16.1322f
C54 bgr_0.START_UP bgr_0.NFET_GATE_10uA 0.529424f
C55 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.err_amp_out 0.4371f
C56 bgr_0.1st_Vout_1 bgr_0.START_UP 0.030647f
C57 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.cap_res_X 0.04831f
C58 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.Y 1.06369f
C59 VDDA GNDA 0.15623p
C60 li_26520_10220# GNDA 0.049096f $ **FLOATING
C61 li_25120_10220# GNDA 0.043891f $ **FLOATING
C62 li_30020_10330# GNDA 0.050514f $ **FLOATING
C63 li_28620_10330# GNDA 0.049721f $ **FLOATING
C64 li_21620_10330# GNDA 0.047034f $ **FLOATING
C65 li_23020_10430# GNDA 0.050654f $ **FLOATING
C66 two_stage_opamp_dummy_magic_0.VIN+ GNDA 2.04185f
C67 two_stage_opamp_dummy_magic_0.VIN- GNDA 2.11372f
C68 bgr_0.START_UP_NFET1 GNDA 5.30912f
C69 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.37246f
C70 bgr_0.1st_Vout_1 GNDA 4.988921f
C71 bgr_0.cap_res2 GNDA 8.276167f
C72 bgr_0.Vbe2 GNDA 17.2131f
C73 bgr_0.START_UP GNDA 7.199363f
C74 bgr_0.V_TOP GNDA 6.820207f
C75 two_stage_opamp_dummy_magic_0.Y GNDA 4.956086f
C76 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 33.49125f
C77 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.661512f
C78 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 8.773118f
C79 bgr_0.NFET_GATE_10uA GNDA 7.5446f
C80 bgr_0.PFET_GATE_10uA GNDA 5.1321f
C81 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 5.42546f
C82 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.547144f
C83 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.61532f
C84 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA 0.01309f
C85 two_stage_opamp_dummy_magic_0.err_amp_out.t3 GNDA 0.01309f
C86 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.037674f
C87 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA 0.01309f
C88 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA 0.01309f
C89 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.036553f
C90 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.4546f
C91 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA 0.01309f
C92 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA 0.01309f
C93 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.036553f
C94 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.485293f
C95 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.093535f
C96 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 1.57366f
C97 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA 0.01309f
C98 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA 0.01309f
C99 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 0.030403f
C100 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.898277f
C101 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA 0.01309f
C102 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA 0.01309f
C103 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.030646f
C104 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.343721f
C105 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA 0.01309f
C106 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA 0.01309f
C107 two_stage_opamp_dummy_magic_0.err_amp_out.n10 GNDA 0.030646f
C108 bgr_0.Vin-.n0 GNDA 0.073641f
C109 bgr_0.Vin-.n1 GNDA 0.338978f
C110 bgr_0.Vin-.n2 GNDA 0.510829f
C111 bgr_0.Vin-.t1 GNDA 0.276208f
C112 bgr_0.Vin-.n3 GNDA 0.331333f
C113 bgr_0.Vin-.n4 GNDA 0.073776f
C114 bgr_0.Vin-.n5 GNDA 0.126176f
C115 bgr_0.Vin-.n6 GNDA 0.074468f
C116 bgr_0.Vin-.n7 GNDA 0.998979f
C117 bgr_0.Vin-.t2 GNDA 0.028614f
C118 bgr_0.Vin-.t5 GNDA 0.028614f
C119 bgr_0.Vin-.n8 GNDA 0.099613f
C120 bgr_0.Vin-.t3 GNDA 0.028614f
C121 bgr_0.Vin-.t4 GNDA 0.028614f
C122 bgr_0.Vin-.n9 GNDA 0.095121f
C123 bgr_0.Vin-.n10 GNDA 0.408067f
C124 bgr_0.Vin-.t0 GNDA 0.098662f
C125 bgr_0.Vin-.n11 GNDA 0.025702f
C126 bgr_0.Vin-.n12 GNDA 0.469862f
C127 bgr_0.Vin-.n13 GNDA 0.222852f
C128 bgr_0.Vin-.t8 GNDA 0.023594f
C129 bgr_0.Vin-.n14 GNDA 0.027673f
C130 bgr_0.Vin-.n15 GNDA 0.022653f
C131 bgr_0.Vin-.n16 GNDA 0.022653f
C132 bgr_0.Vin-.n17 GNDA 0.040466f
C133 bgr_0.Vin-.n18 GNDA 0.524007f
C134 bgr_0.Vin-.n19 GNDA 0.461298f
C135 bgr_0.Vin-.n20 GNDA 0.166915f
C136 bgr_0.Vin-.n21 GNDA 0.074625f
C137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C138 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.024416f
C139 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.069509f
C140 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.094519f
C141 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.120449f
C142 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.042516f
C143 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.078578f
C144 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.050655f
C145 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.120449f
C146 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.042516f
C147 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.078578f
C148 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.050655f
C149 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.050227f
C150 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.094519f
C151 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.281683f
C152 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.420453f
C153 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.242764f
C154 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.242764f
C155 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.242764f
C156 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.242764f
C157 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.182073f
C158 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.121382f
C159 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.182073f
C160 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.242764f
C161 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.242764f
C162 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.242764f
C163 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.242764f
C164 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.420453f
C165 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.281683f
C166 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.069509f
C167 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.097309f
C168 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.024416f
C169 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.024416f
C170 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.084727f
C171 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.024416f
C172 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.024416f
C173 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.084913f
C174 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.024416f
C175 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.024416f
C176 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.084913f
C177 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.024416f
C178 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.024416f
C179 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.084613f
C180 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.15974f
C181 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.024416f
C182 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.024416f
C183 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.084613f
C184 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.082811f
C185 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.024416f
C186 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.024416f
C187 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.084613f
C188 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.082811f
C189 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.099252f
C190 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.024416f
C191 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.024416f
C192 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.08286f
C193 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.100481f
C194 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.094683f
C195 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.024416f
C196 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.024416f
C197 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.084612f
C198 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.078625f
C199 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.024416f
C200 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.024416f
C201 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.084913f
C202 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.024416f
C203 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.024416f
C204 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.084612f
C205 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.15974f
C206 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.029845f
C207 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.057972f
C208 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.079606f
C209 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.024416f
C210 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.015587f
C211 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.015587f
C212 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.056655f
C213 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.015587f
C214 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.015587f
C215 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.04708f
C216 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.294319f
C217 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.19407f
C218 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.046762f
C219 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.046762f
C220 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.193378f
C221 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.046762f
C222 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.046762f
C223 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.192636f
C224 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.267091f
C225 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.046762f
C226 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.046762f
C227 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.192636f
C228 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.139372f
C229 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.046762f
C230 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.046762f
C231 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.192636f
C232 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.139372f
C233 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.046762f
C234 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.046762f
C235 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.192636f
C236 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.200313f
C237 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 2.57755f
C238 bgr_0.V_CMFB_S2 GNDA 2.49029f
C239 bgr_0.Vin+.t1 GNDA 0.125873f
C240 bgr_0.Vin+.t8 GNDA 0.020459f
C241 bgr_0.Vin+.t9 GNDA 0.013299f
C242 bgr_0.Vin+.n0 GNDA 0.04388f
C243 bgr_0.Vin+.t6 GNDA 0.013299f
C244 bgr_0.Vin+.n1 GNDA 0.034146f
C245 bgr_0.Vin+.t7 GNDA 0.013299f
C246 bgr_0.Vin+.n2 GNDA 0.034607f
C247 bgr_0.Vin+.n3 GNDA 0.074523f
C248 bgr_0.Vin+.t5 GNDA 0.043132f
C249 bgr_0.Vin+.t4 GNDA 0.043132f
C250 bgr_0.Vin+.n4 GNDA 0.144858f
C251 bgr_0.Vin+.t2 GNDA 0.043132f
C252 bgr_0.Vin+.t3 GNDA 0.043132f
C253 bgr_0.Vin+.n5 GNDA 0.142496f
C254 bgr_0.Vin+.n6 GNDA 0.656763f
C255 bgr_0.Vin+.n7 GNDA 0.71769f
C256 bgr_0.Vin+.n8 GNDA 0.446219f
C257 bgr_0.Vin+.t0 GNDA 0.137433f
C258 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.024686f
C259 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.024686f
C260 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.082767f
C261 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.024686f
C262 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.024686f
C263 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.080497f
C264 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.650124f
C265 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.024686f
C266 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.024686f
C267 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.082767f
C268 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.024686f
C269 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.024686f
C270 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.080497f
C271 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.650123f
C272 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.339096f
C273 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.122193f
C274 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.122193f
C275 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.122193f
C276 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.122193f
C277 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.14101f
C278 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.114485f
C279 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.070354f
C280 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.070354f
C281 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.065877f
C282 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.122193f
C283 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.122193f
C284 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.122193f
C285 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.122193f
C286 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.14101f
C287 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.114485f
C288 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.070354f
C289 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.070354f
C290 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.065877f
C291 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.044064f
C292 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.122193f
C293 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.122193f
C294 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.122193f
C295 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.122193f
C296 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.14101f
C297 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.114485f
C298 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.070354f
C299 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.070354f
C300 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.065877f
C301 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.122193f
C302 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.122193f
C303 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.122193f
C304 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.122193f
C305 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.14101f
C306 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.114485f
C307 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.070354f
C308 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.070354f
C309 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.065877f
C310 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.044064f
C311 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 1.65653f
C312 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.015552f
C313 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.015552f
C314 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.033701f
C315 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.048299f
C316 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.163832f
C317 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 1.44981f
C318 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.147668f
C319 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 3.20916f
C320 bgr_0.VB2_CUR_BIAS GNDA 2.805f
C321 bgr_0.V_mir1.t9 GNDA 0.03537f
C322 bgr_0.V_mir1.t7 GNDA 0.03537f
C323 bgr_0.V_mir1.t13 GNDA 0.03537f
C324 bgr_0.V_mir1.n0 GNDA 0.08097f
C325 bgr_0.V_mir1.t6 GNDA 0.053881f
C326 bgr_0.V_mir1.t12 GNDA 0.042444f
C327 bgr_0.V_mir1.t17 GNDA 0.042444f
C328 bgr_0.V_mir1.t21 GNDA 0.06851f
C329 bgr_0.V_mir1.n1 GNDA 0.076506f
C330 bgr_0.V_mir1.n2 GNDA 0.052264f
C331 bgr_0.V_mir1.n3 GNDA 0.081315f
C332 bgr_0.V_mir1.n4 GNDA 0.201563f
C333 bgr_0.V_mir1.t5 GNDA 0.03537f
C334 bgr_0.V_mir1.t11 GNDA 0.03537f
C335 bgr_0.V_mir1.n5 GNDA 0.08097f
C336 bgr_0.V_mir1.t4 GNDA 0.053881f
C337 bgr_0.V_mir1.t10 GNDA 0.042444f
C338 bgr_0.V_mir1.t18 GNDA 0.042444f
C339 bgr_0.V_mir1.t22 GNDA 0.06851f
C340 bgr_0.V_mir1.n6 GNDA 0.076506f
C341 bgr_0.V_mir1.n7 GNDA 0.052264f
C342 bgr_0.V_mir1.n8 GNDA 0.081315f
C343 bgr_0.V_mir1.n9 GNDA 0.156007f
C344 bgr_0.V_mir1.t2 GNDA 0.017685f
C345 bgr_0.V_mir1.t0 GNDA 0.017685f
C346 bgr_0.V_mir1.n10 GNDA 0.046242f
C347 bgr_0.V_mir1.t16 GNDA 0.075466f
C348 bgr_0.V_mir1.t1 GNDA 0.017685f
C349 bgr_0.V_mir1.t3 GNDA 0.017685f
C350 bgr_0.V_mir1.n11 GNDA 0.050199f
C351 bgr_0.V_mir1.n12 GNDA 0.827814f
C352 bgr_0.V_mir1.n13 GNDA 0.268286f
C353 bgr_0.V_mir1.n14 GNDA 0.09373f
C354 bgr_0.V_mir1.n15 GNDA 0.699157f
C355 bgr_0.V_mir1.t14 GNDA 0.053881f
C356 bgr_0.V_mir1.t8 GNDA 0.042444f
C357 bgr_0.V_mir1.t20 GNDA 0.042444f
C358 bgr_0.V_mir1.t19 GNDA 0.06851f
C359 bgr_0.V_mir1.n16 GNDA 0.076506f
C360 bgr_0.V_mir1.n17 GNDA 0.052264f
C361 bgr_0.V_mir1.n18 GNDA 0.081315f
C362 bgr_0.V_mir1.n19 GNDA 0.203577f
C363 bgr_0.V_mir1.n20 GNDA 0.08097f
C364 bgr_0.V_mir1.t15 GNDA 0.03537f
C365 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.024373f
C366 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.024373f
C367 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.024373f
C368 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.099127f
C369 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA 0.014624f
C370 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.014624f
C371 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.049685f
C372 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.014624f
C373 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.014624f
C374 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.052539f
C375 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.014624f
C376 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.014624f
C377 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.052133f
C378 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.176305f
C379 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.014624f
C380 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.014624f
C381 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.052133f
C382 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.091767f
C383 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.014624f
C384 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.014624f
C385 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.052133f
C386 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.09128f
C387 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.014624f
C388 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.014624f
C389 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.052516f
C390 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.014624f
C391 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.014624f
C392 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.052133f
C393 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.174572f
C394 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.014624f
C395 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.014624f
C396 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.052133f
C397 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.091767f
C398 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.014624f
C399 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.014624f
C400 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.052133f
C401 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.091767f
C402 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.014624f
C403 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.014624f
C404 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.052133f
C405 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.140027f
C406 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.07702f
C407 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.082224f
C408 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.024373f
C409 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.024373f
C410 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.094049f
C411 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.078027f
C412 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.159231f
C413 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.024373f
C414 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.024373f
C415 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.096773f
C416 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.086515f
C417 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.024373f
C418 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.024373f
C419 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.096773f
C420 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.086515f
C421 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.024373f
C422 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.024373f
C423 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.096773f
C424 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.086515f
C425 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.024373f
C426 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.024373f
C427 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.097223f
C428 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.024373f
C429 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.024373f
C430 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.096773f
C431 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.165755f
C432 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.024373f
C433 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.024373f
C434 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.096773f
C435 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.086515f
C436 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.085877f
C437 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.024373f
C438 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.024373f
C439 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.094049f
C440 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.56785f
C441 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.029248f
C442 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.086515f
C443 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.096773f
C444 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA 0.024373f
C445 bgr_0.V_CUR_REF_REG.t5 GNDA 0.014208f
C446 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C447 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C448 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C449 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C450 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C451 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C452 bgr_0.V_CUR_REF_REG.t2 GNDA 0.42777f
C453 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.092891f
C454 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.011218f
C455 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.018267f
C456 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.106822f
C457 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.021464f
C458 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.095301f
C459 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.011144f
C460 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.091464f
C461 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.021464f
C462 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.066547f
C463 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.021464f
C464 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.204094f
C465 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.098951f
C466 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.092891f
C467 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.321853f
C468 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 0.772935f
C469 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.513063f
C470 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.098962f
C471 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.02127f
C472 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020358f
C473 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020407f
C474 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021244f
C475 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.021116f
C476 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.299998f
C477 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.021116f
C478 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.156484f
C479 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.021116f
C480 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.190977f
C481 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.153542f
C482 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.133374f
C483 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.242929f
C484 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.02127f
C485 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020976f
C486 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.328367f
C487 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020976f
C488 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.180843f
C489 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.180843f
C490 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020976f
C491 bgr_0.cap_res1.t16 GNDA 0.417173f
C492 bgr_0.cap_res1.t19 GNDA 0.418684f
C493 bgr_0.cap_res1.t18 GNDA 0.417173f
C494 bgr_0.cap_res1.t14 GNDA 0.418684f
C495 bgr_0.cap_res1.t8 GNDA 0.417173f
C496 bgr_0.cap_res1.t15 GNDA 0.418684f
C497 bgr_0.cap_res1.t13 GNDA 0.417173f
C498 bgr_0.cap_res1.t6 GNDA 0.418684f
C499 bgr_0.cap_res1.t1 GNDA 0.417173f
C500 bgr_0.cap_res1.t7 GNDA 0.418684f
C501 bgr_0.cap_res1.t5 GNDA 0.417173f
C502 bgr_0.cap_res1.t0 GNDA 0.418684f
C503 bgr_0.cap_res1.t4 GNDA 0.417173f
C504 bgr_0.cap_res1.t12 GNDA 0.418684f
C505 bgr_0.cap_res1.t11 GNDA 0.417173f
C506 bgr_0.cap_res1.t3 GNDA 0.418684f
C507 bgr_0.cap_res1.n0 GNDA 0.279631f
C508 bgr_0.cap_res1.t9 GNDA 0.222685f
C509 bgr_0.cap_res1.n1 GNDA 0.303406f
C510 bgr_0.cap_res1.t2 GNDA 0.222685f
C511 bgr_0.cap_res1.n2 GNDA 0.303406f
C512 bgr_0.cap_res1.t10 GNDA 0.222685f
C513 bgr_0.cap_res1.n3 GNDA 0.303406f
C514 bgr_0.cap_res1.t17 GNDA 0.649059f
C515 bgr_0.cap_res1.t20 GNDA 0.10618f
C516 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.037347f
C517 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.037347f
C518 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.120297f
C519 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.037347f
C520 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.037347f
C521 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.120297f
C522 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.663191f
C523 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.037347f
C524 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.037347f
C525 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.112802f
C526 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.263837f
C527 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.184865f
C528 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.184865f
C529 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.184865f
C530 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.184865f
C531 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.213333f
C532 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.173203f
C533 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.106437f
C534 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.106437f
C535 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.099664f
C536 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.184865f
C537 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.184865f
C538 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.184865f
C539 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.184865f
C540 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.213333f
C541 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.173203f
C542 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.106437f
C543 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.106437f
C544 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.099664f
C545 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.08188f
C546 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.184865f
C547 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.184865f
C548 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.184865f
C549 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.184865f
C550 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.213333f
C551 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.173203f
C552 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.106437f
C553 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.106437f
C554 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.099664f
C555 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.184865f
C556 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.184865f
C557 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.184865f
C558 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.184865f
C559 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.213333f
C560 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.173203f
C561 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.106437f
C562 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.106437f
C563 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.099664f
C564 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.060182f
C565 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 2.37764f
C566 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.214211f
C567 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 1.78048f
C568 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.134447f
C569 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.134447f
C570 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.481197f
C571 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 4.507339f
C572 bgr_0.VB3_CUR_BIAS GNDA 4.06955f
C573 bgr_0.START_UP.t2 GNDA 0.041701f
C574 bgr_0.START_UP.t3 GNDA 0.041701f
C575 bgr_0.START_UP.n0 GNDA 0.151283f
C576 bgr_0.START_UP.t0 GNDA 0.041701f
C577 bgr_0.START_UP.t1 GNDA 0.041701f
C578 bgr_0.START_UP.n1 GNDA 0.139173f
C579 bgr_0.START_UP.n2 GNDA 0.720787f
C580 bgr_0.START_UP.t7 GNDA 0.01567f
C581 bgr_0.START_UP.t6 GNDA 0.01567f
C582 bgr_0.START_UP.n3 GNDA 0.044238f
C583 bgr_0.START_UP.n4 GNDA 0.445182f
C584 bgr_0.START_UP.t4 GNDA 1.66229f
C585 bgr_0.START_UP.t5 GNDA 0.043697f
C586 bgr_0.START_UP.n5 GNDA 1.12863f
C587 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA 0.019956f
C588 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA 0.019956f
C589 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA 0.019956f
C590 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.047077f
C591 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA 0.019956f
C592 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 GNDA 0.019956f
C593 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.04628f
C594 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.872497f
C595 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA 0.019956f
C596 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA 0.019956f
C597 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.04628f
C598 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 2.07772f
C599 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 1.95387f
C600 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA 0.019956f
C601 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA 0.019956f
C602 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.047116f
C603 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA 0.016463f
C604 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA 0.016463f
C605 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA 0.016463f
C606 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA 0.016463f
C607 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA 0.016463f
C608 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA 0.035671f
C609 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.050916f
C610 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA 0.019956f
C611 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA 0.019956f
C612 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.047116f
C613 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.177455f
C614 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.057314f
C615 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.038693f
C616 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.043403f
C617 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.043403f
C618 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.038693f
C619 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.016463f
C620 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA 0.016463f
C621 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA 0.016463f
C622 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA 0.035671f
C623 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.055626f
C624 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.043403f
C625 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.038693f
C626 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.057314f
C627 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.177455f
C628 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.736607f
C629 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.060552f
C630 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA 0.019956f
C631 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.032109f
C632 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.032109f
C633 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.111667f
C634 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.032109f
C635 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.032109f
C636 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.111271f
C637 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.210069f
C638 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.032109f
C639 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.032109f
C640 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.111271f
C641 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.108902f
C642 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.032109f
C643 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.032109f
C644 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.111271f
C645 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.108902f
C646 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.032109f
C647 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.032109f
C648 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.111667f
C649 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.130524f
C650 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.032109f
C651 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.032109f
C652 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.108966f
C653 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.091263f
C654 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.032109f
C655 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.032109f
C656 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.111667f
C657 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.032109f
C658 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.032109f
C659 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.111271f
C660 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.210069f
C661 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.091409f
C662 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.091409f
C663 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.370433f
C664 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.370433f
C665 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.552925f
C666 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.319251f
C667 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.319251f
C668 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.319251f
C669 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.319251f
C670 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.239438f
C671 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.158399f
C672 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.055912f
C673 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.103335f
C674 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.066614f
C675 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.158399f
C676 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.055912f
C677 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.103335f
C678 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.066614f
C679 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.066052f
C680 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.124299f
C681 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.552925f
C682 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.319251f
C683 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.319251f
C684 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.319251f
C685 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.319251f
C686 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.239438f
C687 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.159625f
C688 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.124299f
C689 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.127969f
C690 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.032109f
C691 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.032109f
C692 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.104687f
C693 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.076237f
C694 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.039248f
C695 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.032109f
C696 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.032109f
C697 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.111271f
C698 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.103398f
C699 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.032109f
C700 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.032109f
C701 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.111421f
C702 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.118607f
C703 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.163765f
C704 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.446073f
C705 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.409099f
C706 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.409099f
C707 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.485537f
C708 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.256457f
C709 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.162306f
C710 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.149996f
C711 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.917423f
C712 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.409099f
C713 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.409099f
C714 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.485537f
C715 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.256457f
C716 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.162306f
C717 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.446073f
C718 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.149996f
C719 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.917914f
C720 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.163765f
C721 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.345114f
C722 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.346365f
C723 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.345114f
C724 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.34782f
C725 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.378304f
C726 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.345114f
C727 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.346365f
C728 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.345114f
C729 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.346365f
C730 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.345114f
C731 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.346365f
C732 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.345114f
C733 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.346365f
C734 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.345114f
C735 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.346365f
C736 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.345114f
C737 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.346365f
C738 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.345114f
C739 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.346365f
C740 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.345114f
C741 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.346365f
C742 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345114f
C743 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.346365f
C744 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.345114f
C745 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.346365f
C746 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.345114f
C747 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.346365f
C748 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.345114f
C749 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.346365f
C750 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345114f
C751 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.346365f
C752 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.345114f
C753 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.346365f
C754 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.345114f
C755 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.346365f
C756 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.345114f
C757 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.346365f
C758 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.345114f
C759 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.346365f
C760 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.345114f
C761 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.346365f
C762 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.345114f
C763 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.346365f
C764 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.345114f
C765 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.346365f
C766 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.345114f
C767 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.346365f
C768 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.345114f
C769 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.346365f
C770 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.345114f
C771 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.346365f
C772 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.345114f
C773 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.346365f
C774 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.345114f
C775 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.346365f
C776 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.345114f
C777 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.346365f
C778 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345114f
C779 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.346365f
C780 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.345114f
C781 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.346365f
C782 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.345114f
C783 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.346365f
C784 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.345114f
C785 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.362035f
C786 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.345114f
C787 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.185368f
C788 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198389f
C789 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.345114f
C790 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185368f
C791 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196789f
C792 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345114f
C793 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.185368f
C794 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196789f
C795 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.345114f
C796 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.185368f
C797 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196789f
C798 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.345114f
C799 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185368f
C800 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196789f
C801 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.345114f
C802 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.185368f
C803 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196789f
C804 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.345114f
C805 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185368f
C806 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196789f
C807 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.345114f
C808 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.185368f
C809 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196789f
C810 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.345114f
C811 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.185368f
C812 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196789f
C813 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.345114f
C814 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.346365f
C815 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.166846f
C816 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.215207f
C817 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.18422f
C818 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.233728f
C819 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.18422f
C820 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250999f
C821 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.18422f
C822 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250999f
C823 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.18422f
C824 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250999f
C825 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.18422f
C826 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250999f
C827 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.18422f
C828 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250999f
C829 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.18422f
C830 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250999f
C831 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.18422f
C832 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250999f
C833 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.18422f
C834 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250999f
C835 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.18422f
C836 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250999f
C837 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.18422f
C838 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250999f
C839 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18422f
C840 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250999f
C841 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.18422f
C842 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250999f
C843 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.18422f
C844 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250999f
C845 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.18422f
C846 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250999f
C847 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.18422f
C848 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.233728f
C849 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.343967f
C850 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.166846f
C851 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216458f
C852 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.343967f
C853 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.166846f
C854 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216458f
C855 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.343967f
C856 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.345114f
C857 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.363635f
C858 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.363635f
C859 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.363635f
C860 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.185368f
C861 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216458f
C862 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.343967f
C863 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.166846f
C864 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197936f
C865 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.343967f
C866 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.166846f
C867 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216458f
C868 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.343967f
C869 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.166846f
C870 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216458f
C871 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.343967f
C872 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.166846f
C873 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216458f
C874 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.343967f
C875 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.345114f
C876 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.363635f
C877 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.363635f
C878 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.363635f
C879 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.185368f
C880 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216458f
C881 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.343967f
C882 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.345114f
C883 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.363635f
C884 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.363635f
C885 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363635f
C886 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.185368f
C887 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216458f
C888 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.343967f
C889 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216458f
C890 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.185368f
C891 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.363635f
C892 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.363635f
C893 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.363635f
C894 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.602274f
C895 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.298233f
C896 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA 0.043577f
C897 two_stage_opamp_dummy_magic_0.VOUT+.t17 GNDA 0.043577f
C898 two_stage_opamp_dummy_magic_0.VOUT+.n0 GNDA 0.175148f
C899 two_stage_opamp_dummy_magic_0.VOUT+.t12 GNDA 0.043577f
C900 two_stage_opamp_dummy_magic_0.VOUT+.t16 GNDA 0.043577f
C901 two_stage_opamp_dummy_magic_0.VOUT+.n1 GNDA 0.174825f
C902 two_stage_opamp_dummy_magic_0.VOUT+.n2 GNDA 0.172223f
C903 two_stage_opamp_dummy_magic_0.VOUT+.t11 GNDA 0.043577f
C904 two_stage_opamp_dummy_magic_0.VOUT+.t15 GNDA 0.043577f
C905 two_stage_opamp_dummy_magic_0.VOUT+.n3 GNDA 0.174825f
C906 two_stage_opamp_dummy_magic_0.VOUT+.n4 GNDA 0.088815f
C907 two_stage_opamp_dummy_magic_0.VOUT+.t9 GNDA 0.043577f
C908 two_stage_opamp_dummy_magic_0.VOUT+.t13 GNDA 0.043577f
C909 two_stage_opamp_dummy_magic_0.VOUT+.n5 GNDA 0.174825f
C910 two_stage_opamp_dummy_magic_0.VOUT+.n6 GNDA 0.088815f
C911 two_stage_opamp_dummy_magic_0.VOUT+.t8 GNDA 0.043577f
C912 two_stage_opamp_dummy_magic_0.VOUT+.t2 GNDA 0.043577f
C913 two_stage_opamp_dummy_magic_0.VOUT+.n7 GNDA 0.175148f
C914 two_stage_opamp_dummy_magic_0.VOUT+.n8 GNDA 0.105197f
C915 two_stage_opamp_dummy_magic_0.VOUT+.t10 GNDA 0.043577f
C916 two_stage_opamp_dummy_magic_0.VOUT+.t14 GNDA 0.043577f
C917 two_stage_opamp_dummy_magic_0.VOUT+.n9 GNDA 0.172685f
C918 two_stage_opamp_dummy_magic_0.VOUT+.n10 GNDA 0.210763f
C919 two_stage_opamp_dummy_magic_0.VOUT+.t117 GNDA 0.295461f
C920 two_stage_opamp_dummy_magic_0.VOUT+.t26 GNDA 0.290513f
C921 two_stage_opamp_dummy_magic_0.VOUT+.n11 GNDA 0.194779f
C922 two_stage_opamp_dummy_magic_0.VOUT+.t124 GNDA 0.290513f
C923 two_stage_opamp_dummy_magic_0.VOUT+.n12 GNDA 0.127099f
C924 two_stage_opamp_dummy_magic_0.VOUT+.t72 GNDA 0.295461f
C925 two_stage_opamp_dummy_magic_0.VOUT+.t39 GNDA 0.290513f
C926 two_stage_opamp_dummy_magic_0.VOUT+.n13 GNDA 0.194779f
C927 two_stage_opamp_dummy_magic_0.VOUT+.t127 GNDA 0.290513f
C928 two_stage_opamp_dummy_magic_0.VOUT+.t35 GNDA 0.294841f
C929 two_stage_opamp_dummy_magic_0.VOUT+.t87 GNDA 0.294841f
C930 two_stage_opamp_dummy_magic_0.VOUT+.t43 GNDA 0.294841f
C931 two_stage_opamp_dummy_magic_0.VOUT+.t96 GNDA 0.294841f
C932 two_stage_opamp_dummy_magic_0.VOUT+.t143 GNDA 0.294841f
C933 two_stage_opamp_dummy_magic_0.VOUT+.t106 GNDA 0.294841f
C934 two_stage_opamp_dummy_magic_0.VOUT+.t154 GNDA 0.294841f
C935 two_stage_opamp_dummy_magic_0.VOUT+.t65 GNDA 0.294841f
C936 two_stage_opamp_dummy_magic_0.VOUT+.t116 GNDA 0.294841f
C937 two_stage_opamp_dummy_magic_0.VOUT+.t73 GNDA 0.294841f
C938 two_stage_opamp_dummy_magic_0.VOUT+.t149 GNDA 0.290513f
C939 two_stage_opamp_dummy_magic_0.VOUT+.n14 GNDA 0.195399f
C940 two_stage_opamp_dummy_magic_0.VOUT+.t59 GNDA 0.290513f
C941 two_stage_opamp_dummy_magic_0.VOUT+.n15 GNDA 0.24987f
C942 two_stage_opamp_dummy_magic_0.VOUT+.t97 GNDA 0.290513f
C943 two_stage_opamp_dummy_magic_0.VOUT+.n16 GNDA 0.24987f
C944 two_stage_opamp_dummy_magic_0.VOUT+.t131 GNDA 0.290513f
C945 two_stage_opamp_dummy_magic_0.VOUT+.n17 GNDA 0.24987f
C946 two_stage_opamp_dummy_magic_0.VOUT+.t24 GNDA 0.290513f
C947 two_stage_opamp_dummy_magic_0.VOUT+.n18 GNDA 0.24987f
C948 two_stage_opamp_dummy_magic_0.VOUT+.t75 GNDA 0.290513f
C949 two_stage_opamp_dummy_magic_0.VOUT+.n19 GNDA 0.24987f
C950 two_stage_opamp_dummy_magic_0.VOUT+.t112 GNDA 0.290513f
C951 two_stage_opamp_dummy_magic_0.VOUT+.n20 GNDA 0.24987f
C952 two_stage_opamp_dummy_magic_0.VOUT+.t144 GNDA 0.290513f
C953 two_stage_opamp_dummy_magic_0.VOUT+.n21 GNDA 0.24987f
C954 two_stage_opamp_dummy_magic_0.VOUT+.t55 GNDA 0.290513f
C955 two_stage_opamp_dummy_magic_0.VOUT+.n22 GNDA 0.24987f
C956 two_stage_opamp_dummy_magic_0.VOUT+.t95 GNDA 0.290513f
C957 two_stage_opamp_dummy_magic_0.VOUT+.n23 GNDA 0.24987f
C958 two_stage_opamp_dummy_magic_0.VOUT+.n24 GNDA 0.236042f
C959 two_stage_opamp_dummy_magic_0.VOUT+.t38 GNDA 0.295461f
C960 two_stage_opamp_dummy_magic_0.VOUT+.t142 GNDA 0.290513f
C961 two_stage_opamp_dummy_magic_0.VOUT+.n25 GNDA 0.194779f
C962 two_stage_opamp_dummy_magic_0.VOUT+.t94 GNDA 0.290513f
C963 two_stage_opamp_dummy_magic_0.VOUT+.t20 GNDA 0.295461f
C964 two_stage_opamp_dummy_magic_0.VOUT+.t58 GNDA 0.290513f
C965 two_stage_opamp_dummy_magic_0.VOUT+.n26 GNDA 0.194779f
C966 two_stage_opamp_dummy_magic_0.VOUT+.n27 GNDA 0.236042f
C967 two_stage_opamp_dummy_magic_0.VOUT+.t80 GNDA 0.295461f
C968 two_stage_opamp_dummy_magic_0.VOUT+.t42 GNDA 0.290513f
C969 two_stage_opamp_dummy_magic_0.VOUT+.n28 GNDA 0.194779f
C970 two_stage_opamp_dummy_magic_0.VOUT+.t133 GNDA 0.290513f
C971 two_stage_opamp_dummy_magic_0.VOUT+.t61 GNDA 0.295461f
C972 two_stage_opamp_dummy_magic_0.VOUT+.t100 GNDA 0.290513f
C973 two_stage_opamp_dummy_magic_0.VOUT+.n29 GNDA 0.194779f
C974 two_stage_opamp_dummy_magic_0.VOUT+.n30 GNDA 0.236042f
C975 two_stage_opamp_dummy_magic_0.VOUT+.t121 GNDA 0.295461f
C976 two_stage_opamp_dummy_magic_0.VOUT+.t84 GNDA 0.290513f
C977 two_stage_opamp_dummy_magic_0.VOUT+.n31 GNDA 0.194779f
C978 two_stage_opamp_dummy_magic_0.VOUT+.t32 GNDA 0.290513f
C979 two_stage_opamp_dummy_magic_0.VOUT+.t104 GNDA 0.295461f
C980 two_stage_opamp_dummy_magic_0.VOUT+.t137 GNDA 0.290513f
C981 two_stage_opamp_dummy_magic_0.VOUT+.n32 GNDA 0.194779f
C982 two_stage_opamp_dummy_magic_0.VOUT+.n33 GNDA 0.236042f
C983 two_stage_opamp_dummy_magic_0.VOUT+.t85 GNDA 0.295461f
C984 two_stage_opamp_dummy_magic_0.VOUT+.t50 GNDA 0.290513f
C985 two_stage_opamp_dummy_magic_0.VOUT+.n34 GNDA 0.194779f
C986 two_stage_opamp_dummy_magic_0.VOUT+.t138 GNDA 0.290513f
C987 two_stage_opamp_dummy_magic_0.VOUT+.t67 GNDA 0.295461f
C988 two_stage_opamp_dummy_magic_0.VOUT+.t103 GNDA 0.290513f
C989 two_stage_opamp_dummy_magic_0.VOUT+.n35 GNDA 0.194779f
C990 two_stage_opamp_dummy_magic_0.VOUT+.n36 GNDA 0.236042f
C991 two_stage_opamp_dummy_magic_0.VOUT+.t123 GNDA 0.295461f
C992 two_stage_opamp_dummy_magic_0.VOUT+.t90 GNDA 0.290513f
C993 two_stage_opamp_dummy_magic_0.VOUT+.n37 GNDA 0.194779f
C994 two_stage_opamp_dummy_magic_0.VOUT+.t36 GNDA 0.290513f
C995 two_stage_opamp_dummy_magic_0.VOUT+.t107 GNDA 0.295337f
C996 two_stage_opamp_dummy_magic_0.VOUT+.t141 GNDA 0.290513f
C997 two_stage_opamp_dummy_magic_0.VOUT+.n38 GNDA 0.193087f
C998 two_stage_opamp_dummy_magic_0.VOUT+.n39 GNDA 0.236042f
C999 two_stage_opamp_dummy_magic_0.VOUT+.t108 GNDA 0.295461f
C1000 two_stage_opamp_dummy_magic_0.VOUT+.t70 GNDA 0.290513f
C1001 two_stage_opamp_dummy_magic_0.VOUT+.n40 GNDA 0.194779f
C1002 two_stage_opamp_dummy_magic_0.VOUT+.t91 GNDA 0.290513f
C1003 two_stage_opamp_dummy_magic_0.VOUT+.n41 GNDA 0.127099f
C1004 two_stage_opamp_dummy_magic_0.VOUT+.t68 GNDA 0.295461f
C1005 two_stage_opamp_dummy_magic_0.VOUT+.t31 GNDA 0.290513f
C1006 two_stage_opamp_dummy_magic_0.VOUT+.n42 GNDA 0.194779f
C1007 two_stage_opamp_dummy_magic_0.VOUT+.t52 GNDA 0.290513f
C1008 two_stage_opamp_dummy_magic_0.VOUT+.t54 GNDA 0.294841f
C1009 two_stage_opamp_dummy_magic_0.VOUT+.t156 GNDA 0.294841f
C1010 two_stage_opamp_dummy_magic_0.VOUT+.t145 GNDA 0.295461f
C1011 two_stage_opamp_dummy_magic_0.VOUT+.t45 GNDA 0.290513f
C1012 two_stage_opamp_dummy_magic_0.VOUT+.n43 GNDA 0.194779f
C1013 two_stage_opamp_dummy_magic_0.VOUT+.t136 GNDA 0.290513f
C1014 two_stage_opamp_dummy_magic_0.VOUT+.n44 GNDA 0.127099f
C1015 two_stage_opamp_dummy_magic_0.VOUT+.t101 GNDA 0.290513f
C1016 two_stage_opamp_dummy_magic_0.VOUT+.n45 GNDA 0.12256f
C1017 two_stage_opamp_dummy_magic_0.VOUT+.t37 GNDA 0.294841f
C1018 two_stage_opamp_dummy_magic_0.VOUT+.t113 GNDA 0.295461f
C1019 two_stage_opamp_dummy_magic_0.VOUT+.t151 GNDA 0.290513f
C1020 two_stage_opamp_dummy_magic_0.VOUT+.n46 GNDA 0.194779f
C1021 two_stage_opamp_dummy_magic_0.VOUT+.t98 GNDA 0.290513f
C1022 two_stage_opamp_dummy_magic_0.VOUT+.n47 GNDA 0.127099f
C1023 two_stage_opamp_dummy_magic_0.VOUT+.t60 GNDA 0.290513f
C1024 two_stage_opamp_dummy_magic_0.VOUT+.n48 GNDA 0.12256f
C1025 two_stage_opamp_dummy_magic_0.VOUT+.t140 GNDA 0.294841f
C1026 two_stage_opamp_dummy_magic_0.VOUT+.t76 GNDA 0.295461f
C1027 two_stage_opamp_dummy_magic_0.VOUT+.t118 GNDA 0.290513f
C1028 two_stage_opamp_dummy_magic_0.VOUT+.n49 GNDA 0.194779f
C1029 two_stage_opamp_dummy_magic_0.VOUT+.t57 GNDA 0.290513f
C1030 two_stage_opamp_dummy_magic_0.VOUT+.n50 GNDA 0.127099f
C1031 two_stage_opamp_dummy_magic_0.VOUT+.t21 GNDA 0.290513f
C1032 two_stage_opamp_dummy_magic_0.VOUT+.n51 GNDA 0.12256f
C1033 two_stage_opamp_dummy_magic_0.VOUT+.t105 GNDA 0.294841f
C1034 two_stage_opamp_dummy_magic_0.VOUT+.t25 GNDA 0.295461f
C1035 two_stage_opamp_dummy_magic_0.VOUT+.t66 GNDA 0.290513f
C1036 two_stage_opamp_dummy_magic_0.VOUT+.n52 GNDA 0.194779f
C1037 two_stage_opamp_dummy_magic_0.VOUT+.t81 GNDA 0.290513f
C1038 two_stage_opamp_dummy_magic_0.VOUT+.n53 GNDA 0.127099f
C1039 two_stage_opamp_dummy_magic_0.VOUT+.t44 GNDA 0.290513f
C1040 two_stage_opamp_dummy_magic_0.VOUT+.n54 GNDA 0.12256f
C1041 two_stage_opamp_dummy_magic_0.VOUT+.t125 GNDA 0.294841f
C1042 two_stage_opamp_dummy_magic_0.VOUT+.t88 GNDA 0.294841f
C1043 two_stage_opamp_dummy_magic_0.VOUT+.t51 GNDA 0.294841f
C1044 two_stage_opamp_dummy_magic_0.VOUT+.t150 GNDA 0.294841f
C1045 two_stage_opamp_dummy_magic_0.VOUT+.t33 GNDA 0.294841f
C1046 two_stage_opamp_dummy_magic_0.VOUT+.t134 GNDA 0.290513f
C1047 two_stage_opamp_dummy_magic_0.VOUT+.n55 GNDA 0.195399f
C1048 two_stage_opamp_dummy_magic_0.VOUT+.t110 GNDA 0.290513f
C1049 two_stage_opamp_dummy_magic_0.VOUT+.n56 GNDA 0.24987f
C1050 two_stage_opamp_dummy_magic_0.VOUT+.t147 GNDA 0.290513f
C1051 two_stage_opamp_dummy_magic_0.VOUT+.n57 GNDA 0.24987f
C1052 two_stage_opamp_dummy_magic_0.VOUT+.t46 GNDA 0.290513f
C1053 two_stage_opamp_dummy_magic_0.VOUT+.n58 GNDA 0.24987f
C1054 two_stage_opamp_dummy_magic_0.VOUT+.t86 GNDA 0.290513f
C1055 two_stage_opamp_dummy_magic_0.VOUT+.n59 GNDA 0.30888f
C1056 two_stage_opamp_dummy_magic_0.VOUT+.t62 GNDA 0.290513f
C1057 two_stage_opamp_dummy_magic_0.VOUT+.n60 GNDA 0.30888f
C1058 two_stage_opamp_dummy_magic_0.VOUT+.t102 GNDA 0.290513f
C1059 two_stage_opamp_dummy_magic_0.VOUT+.n61 GNDA 0.30888f
C1060 two_stage_opamp_dummy_magic_0.VOUT+.t139 GNDA 0.290513f
C1061 two_stage_opamp_dummy_magic_0.VOUT+.n62 GNDA 0.30888f
C1062 two_stage_opamp_dummy_magic_0.VOUT+.t119 GNDA 0.290513f
C1063 two_stage_opamp_dummy_magic_0.VOUT+.n63 GNDA 0.24987f
C1064 two_stage_opamp_dummy_magic_0.VOUT+.t155 GNDA 0.290513f
C1065 two_stage_opamp_dummy_magic_0.VOUT+.n64 GNDA 0.24987f
C1066 two_stage_opamp_dummy_magic_0.VOUT+.n65 GNDA 0.236042f
C1067 two_stage_opamp_dummy_magic_0.VOUT+.t28 GNDA 0.295461f
C1068 two_stage_opamp_dummy_magic_0.VOUT+.t130 GNDA 0.290513f
C1069 two_stage_opamp_dummy_magic_0.VOUT+.n66 GNDA 0.194779f
C1070 two_stage_opamp_dummy_magic_0.VOUT+.t152 GNDA 0.290513f
C1071 two_stage_opamp_dummy_magic_0.VOUT+.t77 GNDA 0.295461f
C1072 two_stage_opamp_dummy_magic_0.VOUT+.t115 GNDA 0.290513f
C1073 two_stage_opamp_dummy_magic_0.VOUT+.n67 GNDA 0.194779f
C1074 two_stage_opamp_dummy_magic_0.VOUT+.n68 GNDA 0.236042f
C1075 two_stage_opamp_dummy_magic_0.VOUT+.t63 GNDA 0.295461f
C1076 two_stage_opamp_dummy_magic_0.VOUT+.t23 GNDA 0.290513f
C1077 two_stage_opamp_dummy_magic_0.VOUT+.n69 GNDA 0.194779f
C1078 two_stage_opamp_dummy_magic_0.VOUT+.t48 GNDA 0.290513f
C1079 two_stage_opamp_dummy_magic_0.VOUT+.t111 GNDA 0.295461f
C1080 two_stage_opamp_dummy_magic_0.VOUT+.t148 GNDA 0.290513f
C1081 two_stage_opamp_dummy_magic_0.VOUT+.n70 GNDA 0.194779f
C1082 two_stage_opamp_dummy_magic_0.VOUT+.n71 GNDA 0.236042f
C1083 two_stage_opamp_dummy_magic_0.VOUT+.t114 GNDA 0.295461f
C1084 two_stage_opamp_dummy_magic_0.VOUT+.t79 GNDA 0.290513f
C1085 two_stage_opamp_dummy_magic_0.VOUT+.n72 GNDA 0.194779f
C1086 two_stage_opamp_dummy_magic_0.VOUT+.t27 GNDA 0.290513f
C1087 two_stage_opamp_dummy_magic_0.VOUT+.t99 GNDA 0.295461f
C1088 two_stage_opamp_dummy_magic_0.VOUT+.t132 GNDA 0.290513f
C1089 two_stage_opamp_dummy_magic_0.VOUT+.n73 GNDA 0.194779f
C1090 two_stage_opamp_dummy_magic_0.VOUT+.n74 GNDA 0.236042f
C1091 two_stage_opamp_dummy_magic_0.VOUT+.t74 GNDA 0.295461f
C1092 two_stage_opamp_dummy_magic_0.VOUT+.t40 GNDA 0.290513f
C1093 two_stage_opamp_dummy_magic_0.VOUT+.n75 GNDA 0.194779f
C1094 two_stage_opamp_dummy_magic_0.VOUT+.t128 GNDA 0.290513f
C1095 two_stage_opamp_dummy_magic_0.VOUT+.t56 GNDA 0.295461f
C1096 two_stage_opamp_dummy_magic_0.VOUT+.t93 GNDA 0.290513f
C1097 two_stage_opamp_dummy_magic_0.VOUT+.n76 GNDA 0.194779f
C1098 two_stage_opamp_dummy_magic_0.VOUT+.n77 GNDA 0.236042f
C1099 two_stage_opamp_dummy_magic_0.VOUT+.t109 GNDA 0.295461f
C1100 two_stage_opamp_dummy_magic_0.VOUT+.t71 GNDA 0.290513f
C1101 two_stage_opamp_dummy_magic_0.VOUT+.n78 GNDA 0.194779f
C1102 two_stage_opamp_dummy_magic_0.VOUT+.t19 GNDA 0.290513f
C1103 two_stage_opamp_dummy_magic_0.VOUT+.t92 GNDA 0.295461f
C1104 two_stage_opamp_dummy_magic_0.VOUT+.t126 GNDA 0.290513f
C1105 two_stage_opamp_dummy_magic_0.VOUT+.n79 GNDA 0.194779f
C1106 two_stage_opamp_dummy_magic_0.VOUT+.n80 GNDA 0.236042f
C1107 two_stage_opamp_dummy_magic_0.VOUT+.t69 GNDA 0.295461f
C1108 two_stage_opamp_dummy_magic_0.VOUT+.t34 GNDA 0.290513f
C1109 two_stage_opamp_dummy_magic_0.VOUT+.n81 GNDA 0.194779f
C1110 two_stage_opamp_dummy_magic_0.VOUT+.t122 GNDA 0.290513f
C1111 two_stage_opamp_dummy_magic_0.VOUT+.t53 GNDA 0.295461f
C1112 two_stage_opamp_dummy_magic_0.VOUT+.t89 GNDA 0.290513f
C1113 two_stage_opamp_dummy_magic_0.VOUT+.n82 GNDA 0.194779f
C1114 two_stage_opamp_dummy_magic_0.VOUT+.n83 GNDA 0.236042f
C1115 two_stage_opamp_dummy_magic_0.VOUT+.t30 GNDA 0.295461f
C1116 two_stage_opamp_dummy_magic_0.VOUT+.t135 GNDA 0.290513f
C1117 two_stage_opamp_dummy_magic_0.VOUT+.n84 GNDA 0.194779f
C1118 two_stage_opamp_dummy_magic_0.VOUT+.t83 GNDA 0.290513f
C1119 two_stage_opamp_dummy_magic_0.VOUT+.t153 GNDA 0.295461f
C1120 two_stage_opamp_dummy_magic_0.VOUT+.t49 GNDA 0.290513f
C1121 two_stage_opamp_dummy_magic_0.VOUT+.n85 GNDA 0.194779f
C1122 two_stage_opamp_dummy_magic_0.VOUT+.n86 GNDA 0.236042f
C1123 two_stage_opamp_dummy_magic_0.VOUT+.t64 GNDA 0.295461f
C1124 two_stage_opamp_dummy_magic_0.VOUT+.t29 GNDA 0.290513f
C1125 two_stage_opamp_dummy_magic_0.VOUT+.n87 GNDA 0.194779f
C1126 two_stage_opamp_dummy_magic_0.VOUT+.t120 GNDA 0.290513f
C1127 two_stage_opamp_dummy_magic_0.VOUT+.t47 GNDA 0.295461f
C1128 two_stage_opamp_dummy_magic_0.VOUT+.t82 GNDA 0.290513f
C1129 two_stage_opamp_dummy_magic_0.VOUT+.n88 GNDA 0.194779f
C1130 two_stage_opamp_dummy_magic_0.VOUT+.n89 GNDA 0.236042f
C1131 two_stage_opamp_dummy_magic_0.VOUT+.t22 GNDA 0.295461f
C1132 two_stage_opamp_dummy_magic_0.VOUT+.t129 GNDA 0.290513f
C1133 two_stage_opamp_dummy_magic_0.VOUT+.n90 GNDA 0.194779f
C1134 two_stage_opamp_dummy_magic_0.VOUT+.t78 GNDA 0.290513f
C1135 two_stage_opamp_dummy_magic_0.VOUT+.n91 GNDA 0.236042f
C1136 two_stage_opamp_dummy_magic_0.VOUT+.t41 GNDA 0.290513f
C1137 two_stage_opamp_dummy_magic_0.VOUT+.n92 GNDA 0.127099f
C1138 two_stage_opamp_dummy_magic_0.VOUT+.t146 GNDA 0.290513f
C1139 two_stage_opamp_dummy_magic_0.VOUT+.n93 GNDA 0.238016f
C1140 two_stage_opamp_dummy_magic_0.VOUT+.n94 GNDA 0.28569f
C1141 two_stage_opamp_dummy_magic_0.VOUT+.t5 GNDA 0.05084f
C1142 two_stage_opamp_dummy_magic_0.VOUT+.t6 GNDA 0.05084f
C1143 two_stage_opamp_dummy_magic_0.VOUT+.n95 GNDA 0.235187f
C1144 two_stage_opamp_dummy_magic_0.VOUT+.t3 GNDA 0.05084f
C1145 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA 0.05084f
C1146 two_stage_opamp_dummy_magic_0.VOUT+.n96 GNDA 0.2344f
C1147 two_stage_opamp_dummy_magic_0.VOUT+.n97 GNDA 0.144847f
C1148 two_stage_opamp_dummy_magic_0.VOUT+.t7 GNDA 0.05084f
C1149 two_stage_opamp_dummy_magic_0.VOUT+.t4 GNDA 0.05084f
C1150 two_stage_opamp_dummy_magic_0.VOUT+.n98 GNDA 0.2344f
C1151 two_stage_opamp_dummy_magic_0.VOUT+.n99 GNDA 0.089159f
C1152 two_stage_opamp_dummy_magic_0.VOUT+.n100 GNDA 0.165939f
C1153 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA 0.084056f
C1154 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.027492f
C1155 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.022846f
C1156 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.142463f
C1157 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.09411f
C1158 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.022691f
C1159 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.022691f
C1160 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.093837f
C1161 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.022691f
C1162 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.022691f
C1163 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.093477f
C1164 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.129606f
C1165 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.022691f
C1166 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.022691f
C1167 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.093477f
C1168 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.06763f
C1169 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.022691f
C1170 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.022691f
C1171 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.093477f
C1172 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.06763f
C1173 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.022691f
C1174 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.022691f
C1175 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.093477f
C1176 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.097762f
C1177 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.61699f
C1178 bgr_0.V_CMFB_S4 GNDA 0.50856f
C1179 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.053187f
C1180 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.053187f
C1181 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.184972f
C1182 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.053187f
C1183 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.053187f
C1184 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.184316f
C1185 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.347971f
C1186 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.053187f
C1187 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.053187f
C1188 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.184316f
C1189 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.180392f
C1190 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.053187f
C1191 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.053187f
C1192 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.184316f
C1193 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.180392f
C1194 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.053187f
C1195 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.053187f
C1196 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.184316f
C1197 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.212415f
C1198 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.053187f
C1199 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.053187f
C1200 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.180498f
C1201 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.149147f
C1202 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.022794f
C1203 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.022794f
C1204 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.076959f
C1205 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.022794f
C1206 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.022794f
C1207 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.082252f
C1208 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.022794f
C1209 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.022794f
C1210 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.081534f
C1211 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.302737f
C1212 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.022794f
C1213 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.022794f
C1214 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.081534f
C1215 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.157046f
C1216 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.022794f
C1217 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.022794f
C1218 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.081534f
C1219 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.157046f
C1220 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.022794f
C1221 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.022794f
C1222 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.082252f
C1223 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.191279f
C1224 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.123631f
C1225 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.031912f
C1226 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.031912f
C1227 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.031912f
C1228 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.031912f
C1229 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.031912f
C1230 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.031912f
C1231 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.031912f
C1232 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.03875f
C1233 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.03875f
C1234 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.025074f
C1235 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.025074f
C1236 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.025074f
C1237 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.025074f
C1238 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.025074f
C1239 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.022459f
C1240 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.031912f
C1241 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.03875f
C1242 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.036135f
C1243 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.022101f
C1244 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.049008f
C1245 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.049008f
C1246 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.049008f
C1247 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.049008f
C1248 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.049008f
C1249 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.049008f
C1250 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.049008f
C1251 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.055713f
C1252 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.05028f
C1253 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.030772f
C1254 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.030772f
C1255 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.030772f
C1256 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.030772f
C1257 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.030772f
C1258 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.028157f
C1259 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.049008f
C1260 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.055713f
C1261 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.047665f
C1262 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.022031f
C1263 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.153015f
C1264 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.741299f
C1265 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.100295f
C1266 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.100295f
C1267 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.106821f
C1268 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.084651f
C1269 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.045253f
C1270 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.100295f
C1271 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.100295f
C1272 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.100295f
C1273 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.100295f
C1274 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.100295f
C1275 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.100295f
C1276 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.106821f
C1277 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.084651f
C1278 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.047868f
C1279 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.047868f
C1280 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.047868f
C1281 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.047868f
C1282 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.045253f
C1283 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.024415f
C1284 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 1.03694f
C1285 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.458663f
C1286 bgr_0.V_TOP.t15 GNDA 0.115045f
C1287 bgr_0.V_TOP.t19 GNDA 0.115045f
C1288 bgr_0.V_TOP.t24 GNDA 0.115045f
C1289 bgr_0.V_TOP.t41 GNDA 0.115045f
C1290 bgr_0.V_TOP.t43 GNDA 0.115045f
C1291 bgr_0.V_TOP.t20 GNDA 0.115045f
C1292 bgr_0.V_TOP.t26 GNDA 0.115045f
C1293 bgr_0.V_TOP.t31 GNDA 0.115045f
C1294 bgr_0.V_TOP.t45 GNDA 0.115045f
C1295 bgr_0.V_TOP.t49 GNDA 0.115045f
C1296 bgr_0.V_TOP.t29 GNDA 0.115045f
C1297 bgr_0.V_TOP.t32 GNDA 0.115045f
C1298 bgr_0.V_TOP.t34 GNDA 0.115045f
C1299 bgr_0.V_TOP.t40 GNDA 0.115045f
C1300 bgr_0.V_TOP.t18 GNDA 0.150392f
C1301 bgr_0.V_TOP.n0 GNDA 0.084081f
C1302 bgr_0.V_TOP.n1 GNDA 0.061357f
C1303 bgr_0.V_TOP.n2 GNDA 0.061357f
C1304 bgr_0.V_TOP.n3 GNDA 0.061357f
C1305 bgr_0.V_TOP.n4 GNDA 0.061357f
C1306 bgr_0.V_TOP.n5 GNDA 0.057217f
C1307 bgr_0.V_TOP.t4 GNDA 0.147947f
C1308 bgr_0.V_TOP.t13 GNDA 0.155772f
C1309 bgr_0.V_TOP.t2 GNDA 0.010957f
C1310 bgr_0.V_TOP.t8 GNDA 0.010957f
C1311 bgr_0.V_TOP.n6 GNDA 0.027281f
C1312 bgr_0.V_TOP.n7 GNDA 0.726844f
C1313 bgr_0.V_TOP.t3 GNDA 0.010957f
C1314 bgr_0.V_TOP.t12 GNDA 0.010957f
C1315 bgr_0.V_TOP.n8 GNDA 0.027465f
C1316 bgr_0.V_TOP.t11 GNDA 0.010957f
C1317 bgr_0.V_TOP.t1 GNDA 0.010957f
C1318 bgr_0.V_TOP.n9 GNDA 0.027281f
C1319 bgr_0.V_TOP.n10 GNDA 0.252824f
C1320 bgr_0.V_TOP.t7 GNDA 0.010957f
C1321 bgr_0.V_TOP.t9 GNDA 0.010957f
C1322 bgr_0.V_TOP.n11 GNDA 0.026425f
C1323 bgr_0.V_TOP.n12 GNDA 0.153577f
C1324 bgr_0.V_TOP.n13 GNDA 0.087653f
C1325 bgr_0.V_TOP.t5 GNDA 0.010957f
C1326 bgr_0.V_TOP.t6 GNDA 0.010957f
C1327 bgr_0.V_TOP.n14 GNDA 0.027281f
C1328 bgr_0.V_TOP.n15 GNDA 0.151313f
C1329 bgr_0.V_TOP.t10 GNDA 0.010957f
C1330 bgr_0.V_TOP.t0 GNDA 0.010957f
C1331 bgr_0.V_TOP.n16 GNDA 0.027281f
C1332 bgr_0.V_TOP.n17 GNDA 0.149874f
C1333 bgr_0.V_TOP.n18 GNDA 0.329448f
C1334 bgr_0.V_TOP.n19 GNDA 0.023183f
C1335 bgr_0.V_TOP.n20 GNDA 0.057217f
C1336 bgr_0.V_TOP.n21 GNDA 0.061357f
C1337 bgr_0.V_TOP.n22 GNDA 0.061357f
C1338 bgr_0.V_TOP.n23 GNDA 0.061357f
C1339 bgr_0.V_TOP.n24 GNDA 0.061357f
C1340 bgr_0.V_TOP.n25 GNDA 0.061357f
C1341 bgr_0.V_TOP.n26 GNDA 0.061357f
C1342 bgr_0.V_TOP.n27 GNDA 0.057217f
C1343 bgr_0.V_TOP.t39 GNDA 0.132572f
C1344 bgr_0.V_TOP.t37 GNDA 0.445732f
C1345 bgr_0.V_TOP.t30 GNDA 0.438267f
C1346 bgr_0.V_TOP.n28 GNDA 0.293844f
C1347 bgr_0.V_TOP.t17 GNDA 0.438267f
C1348 bgr_0.V_TOP.t48 GNDA 0.445732f
C1349 bgr_0.V_TOP.t23 GNDA 0.438267f
C1350 bgr_0.V_TOP.n29 GNDA 0.293844f
C1351 bgr_0.V_TOP.n30 GNDA 0.273917f
C1352 bgr_0.V_TOP.t44 GNDA 0.445732f
C1353 bgr_0.V_TOP.t36 GNDA 0.438267f
C1354 bgr_0.V_TOP.n31 GNDA 0.293844f
C1355 bgr_0.V_TOP.t28 GNDA 0.438267f
C1356 bgr_0.V_TOP.t22 GNDA 0.445732f
C1357 bgr_0.V_TOP.t33 GNDA 0.438267f
C1358 bgr_0.V_TOP.n32 GNDA 0.293844f
C1359 bgr_0.V_TOP.n33 GNDA 0.356092f
C1360 bgr_0.V_TOP.t35 GNDA 0.445732f
C1361 bgr_0.V_TOP.t27 GNDA 0.438267f
C1362 bgr_0.V_TOP.n34 GNDA 0.293844f
C1363 bgr_0.V_TOP.t16 GNDA 0.438267f
C1364 bgr_0.V_TOP.t47 GNDA 0.445732f
C1365 bgr_0.V_TOP.t21 GNDA 0.438267f
C1366 bgr_0.V_TOP.n35 GNDA 0.293844f
C1367 bgr_0.V_TOP.n36 GNDA 0.356092f
C1368 bgr_0.V_TOP.t25 GNDA 0.445732f
C1369 bgr_0.V_TOP.t14 GNDA 0.438267f
C1370 bgr_0.V_TOP.n37 GNDA 0.293844f
C1371 bgr_0.V_TOP.t42 GNDA 0.438267f
C1372 bgr_0.V_TOP.n38 GNDA 0.273917f
C1373 bgr_0.V_TOP.t46 GNDA 0.438267f
C1374 bgr_0.V_TOP.n39 GNDA 0.191742f
C1375 bgr_0.V_TOP.t38 GNDA 0.438267f
C1376 bgr_0.V_TOP.n40 GNDA 0.893239f
C1377 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C1378 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C1379 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C1380 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C1381 bgr_0.1st_Vout_1.t31 GNDA 0.352846f
C1382 bgr_0.1st_Vout_1.t20 GNDA 0.346937f
C1383 bgr_0.1st_Vout_1.t25 GNDA 0.346937f
C1384 bgr_0.1st_Vout_1.t22 GNDA 0.352846f
C1385 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C1386 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C1387 bgr_0.1st_Vout_1.t28 GNDA 0.346937f
C1388 bgr_0.1st_Vout_1.t33 GNDA 0.346937f
C1389 bgr_0.1st_Vout_1.t30 GNDA 0.352846f
C1390 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C1391 bgr_0.1st_Vout_1.t27 GNDA 0.352846f
C1392 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C1393 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C1394 bgr_0.1st_Vout_1.t19 GNDA 0.352846f
C1395 bgr_0.1st_Vout_1.t29 GNDA 0.346937f
C1396 bgr_0.1st_Vout_1.t15 GNDA 0.352846f
C1397 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C1398 bgr_0.1st_Vout_1.t14 GNDA 0.346937f
C1399 bgr_0.1st_Vout_1.t17 GNDA 0.346937f
C1400 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C1401 bgr_0.1st_Vout_1.t21 GNDA 0.022665f
C1402 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C1403 bgr_0.1st_Vout_1.t24 GNDA 0.013213f
C1404 bgr_0.1st_Vout_1.t18 GNDA 0.013213f
C1405 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C1406 bgr_0.1st_Vout_1.n6 GNDA 0.020958f
C1407 bgr_0.1st_Vout_1.t9 GNDA 0.018268f
C1408 bgr_0.1st_Vout_1.n7 GNDA 0.012529f
C1409 bgr_0.1st_Vout_1.n8 GNDA 0.189508f
C1410 bgr_0.1st_Vout_1.n9 GNDA 0.011336f
C1411 bgr_0.1st_Vout_1.t34 GNDA 0.013213f
C1412 bgr_0.1st_Vout_1.t26 GNDA 0.013213f
C1413 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C1414 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C1415 bgr_0.1st_Vout_1.t11 GNDA 0.020738f
C1416 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.013658f
C1417 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.013658f
C1418 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.034236f
C1419 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.013658f
C1420 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.013658f
C1421 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.034056f
C1422 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.302687f
C1423 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.013658f
C1424 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.013658f
C1425 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.027316f
C1426 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.164359f
C1427 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.174921f
C1428 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.027316f
C1429 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.027316f
C1430 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.080145f
C1431 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.027316f
C1432 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.027316f
C1433 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.079781f
C1434 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.27577f
C1435 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.027316f
C1436 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.027316f
C1437 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.079781f
C1438 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.142847f
C1439 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.027316f
C1440 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.027316f
C1441 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.079781f
C1442 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.142847f
C1443 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.027316f
C1444 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.027316f
C1445 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.079781f
C1446 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.205223f
C1447 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 1.58562f
C1448 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 2.05369f
C1449 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.052601f
C1450 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.052601f
C1451 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.182935f
C1452 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.052601f
C1453 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.052601f
C1454 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.182287f
C1455 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.344139f
C1456 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.052601f
C1457 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.052601f
C1458 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.182287f
C1459 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.178405f
C1460 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.052601f
C1461 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.052601f
C1462 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.182287f
C1463 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.178405f
C1464 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.052601f
C1465 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.052601f
C1466 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.182287f
C1467 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.210076f
C1468 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.052601f
C1469 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.052601f
C1470 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.178511f
C1471 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.147505f
C1472 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.022543f
C1473 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.022543f
C1474 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.076111f
C1475 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.022543f
C1476 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.022543f
C1477 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.081346f
C1478 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.022543f
C1479 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.022543f
C1480 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.081346f
C1481 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.022543f
C1482 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.022543f
C1483 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.080636f
C1484 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.299403f
C1485 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.022543f
C1486 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.022543f
C1487 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.080636f
C1488 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.155317f
C1489 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.022543f
C1490 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.022543f
C1491 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.080636f
C1492 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.155317f
C1493 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.189173f
C1494 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.122269f
C1495 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.128676f
C1496 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.03156f
C1497 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.038324f
C1498 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.035737f
C1499 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.03156f
C1500 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.03156f
C1501 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.03156f
C1502 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.03156f
C1503 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.03156f
C1504 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.03156f
C1505 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.03156f
C1506 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.038324f
C1507 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.038324f
C1508 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.024798f
C1509 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.024798f
C1510 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.024798f
C1511 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.024798f
C1512 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.024798f
C1513 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.022211f
C1514 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.021857f
C1515 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.048468f
C1516 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.0551f
C1517 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.04714f
C1518 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.048468f
C1519 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.048468f
C1520 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.048468f
C1521 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.048468f
C1522 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.048468f
C1523 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.048468f
C1524 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.048468f
C1525 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.0551f
C1526 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.049726f
C1527 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.030433f
C1528 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.030433f
C1529 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.030433f
C1530 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.030433f
C1531 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.030433f
C1532 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.027847f
C1533 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.021789f
C1534 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.153028f
C1535 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.454714f
C1536 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.09919f
C1537 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.09919f
C1538 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.09919f
C1539 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.09919f
C1540 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.09919f
C1541 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.09919f
C1542 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.105644f
C1543 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.083719f
C1544 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.047341f
C1545 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.047341f
C1546 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.047341f
C1547 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.047341f
C1548 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.044755f
C1549 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.09919f
C1550 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.09919f
C1551 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.105644f
C1552 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.083719f
C1553 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.044755f
C1554 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.024251f
C1555 two_stage_opamp_dummy_magic_0.X.n52 GNDA 1.03308f
C1556 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.734227f
C1557 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.29369f
C1558 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 7.33588f
C1559 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.015003f
C1560 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.015003f
C1561 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.015003f
C1562 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.015003f
C1563 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.015003f
C1564 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.015003f
C1565 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.015003f
C1566 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.015003f
C1567 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.015003f
C1568 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.015003f
C1569 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.015003f
C1570 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.015003f
C1571 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.015003f
C1572 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.015003f
C1573 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.015003f
C1574 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.015003f
C1575 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.032506f
C1576 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.050691f
C1577 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.039552f
C1578 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.039552f
C1579 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.039552f
C1580 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.039552f
C1581 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.039552f
C1582 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.039552f
C1583 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.039552f
C1584 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.039552f
C1585 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.039552f
C1586 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.039552f
C1587 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.039552f
C1588 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.039552f
C1589 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.039552f
C1590 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.039552f
C1591 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.033846f
C1592 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.015003f
C1593 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.015003f
C1594 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.032506f
C1595 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.050691f
C1596 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.033846f
C1597 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.054538f
C1598 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.03637f
C1599 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.03637f
C1600 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 1.84824f
C1601 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.018185f
C1602 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.018185f
C1603 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.041859f
C1604 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.018185f
C1605 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.018185f
C1606 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.042173f
C1607 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.018185f
C1608 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.018185f
C1609 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.042447f
C1610 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.018185f
C1611 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.018185f
C1612 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.042173f
C1613 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.018185f
C1614 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.018185f
C1615 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.042173f
C1616 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.018185f
C1617 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.018185f
C1618 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.03637f
C1619 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.108338f
C1620 bgr_0.cap_res2.t4 GNDA 0.406156f
C1621 bgr_0.cap_res2.t3 GNDA 0.407628f
C1622 bgr_0.cap_res2.t17 GNDA 0.406156f
C1623 bgr_0.cap_res2.t12 GNDA 0.407628f
C1624 bgr_0.cap_res2.t19 GNDA 0.406156f
C1625 bgr_0.cap_res2.t16 GNDA 0.407628f
C1626 bgr_0.cap_res2.t11 GNDA 0.406156f
C1627 bgr_0.cap_res2.t7 GNDA 0.407628f
C1628 bgr_0.cap_res2.t13 GNDA 0.406156f
C1629 bgr_0.cap_res2.t9 GNDA 0.407628f
C1630 bgr_0.cap_res2.t6 GNDA 0.406156f
C1631 bgr_0.cap_res2.t1 GNDA 0.407628f
C1632 bgr_0.cap_res2.t18 GNDA 0.406156f
C1633 bgr_0.cap_res2.t14 GNDA 0.407628f
C1634 bgr_0.cap_res2.t10 GNDA 0.406156f
C1635 bgr_0.cap_res2.t5 GNDA 0.407628f
C1636 bgr_0.cap_res2.n0 GNDA 0.272247f
C1637 bgr_0.cap_res2.t20 GNDA 0.216805f
C1638 bgr_0.cap_res2.n1 GNDA 0.295394f
C1639 bgr_0.cap_res2.t15 GNDA 0.216805f
C1640 bgr_0.cap_res2.n2 GNDA 0.295394f
C1641 bgr_0.cap_res2.t2 GNDA 0.216805f
C1642 bgr_0.cap_res2.n3 GNDA 0.295394f
C1643 bgr_0.cap_res2.t8 GNDA 0.214043f
C1644 bgr_0.cap_res2.t0 GNDA 0.133038f
C1645 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C1646 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C1647 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C1648 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C1649 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C1650 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C1651 bgr_0.1st_Vout_2.t15 GNDA 0.021508f
C1652 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C1653 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C1654 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C1655 bgr_0.1st_Vout_2.t13 GNDA 0.013652f
C1656 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C1657 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C1658 bgr_0.1st_Vout_2.n10 GNDA 0.021654f
C1659 bgr_0.1st_Vout_2.n11 GNDA 0.012945f
C1660 bgr_0.1st_Vout_2.t9 GNDA 0.018875f
C1661 bgr_0.1st_Vout_2.n12 GNDA 0.195802f
C1662 bgr_0.1st_Vout_2.n13 GNDA 0.011712f
C1663 bgr_0.1st_Vout_2.n14 GNDA 0.049674f
C1664 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C1665 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C1666 bgr_0.1st_Vout_2.t18 GNDA 0.013652f
C1667 bgr_0.1st_Vout_2.t12 GNDA 0.013652f
C1668 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C1669 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C1670 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C1671 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C1672 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C1673 bgr_0.1st_Vout_2.t26 GNDA 0.364565f
C1674 bgr_0.1st_Vout_2.t32 GNDA 0.358459f
C1675 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C1676 bgr_0.1st_Vout_2.t28 GNDA 0.358459f
C1677 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C1678 bgr_0.1st_Vout_2.t31 GNDA 0.364565f
C1679 bgr_0.1st_Vout_2.t36 GNDA 0.358459f
C1680 bgr_0.1st_Vout_2.t14 GNDA 0.364565f
C1681 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C1682 bgr_0.1st_Vout_2.t35 GNDA 0.358459f
C1683 bgr_0.1st_Vout_2.t25 GNDA 0.364565f
C1684 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C1685 bgr_0.1st_Vout_2.t33 GNDA 0.364565f
C1686 bgr_0.1st_Vout_2.t34 GNDA 0.358459f
C1687 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C1688 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C1689 bgr_0.1st_Vout_2.t17 GNDA 0.358459f
C1690 bgr_0.1st_Vout_2.t27 GNDA 0.023417f
C1691 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C1692 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C1693 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C1694 two_stage_opamp_dummy_magic_0.Vb1.t0 GNDA 0.012623f
C1695 two_stage_opamp_dummy_magic_0.Vb1.t5 GNDA 0.012623f
C1696 two_stage_opamp_dummy_magic_0.Vb1.n0 GNDA 0.031643f
C1697 two_stage_opamp_dummy_magic_0.Vb1.t4 GNDA 0.012623f
C1698 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA 0.012623f
C1699 two_stage_opamp_dummy_magic_0.Vb1.n1 GNDA 0.031431f
C1700 two_stage_opamp_dummy_magic_0.Vb1.n2 GNDA 0.296652f
C1701 two_stage_opamp_dummy_magic_0.Vb1.t21 GNDA 0.019408f
C1702 two_stage_opamp_dummy_magic_0.Vb1.t9 GNDA 0.019408f
C1703 two_stage_opamp_dummy_magic_0.Vb1.t6 GNDA 0.019408f
C1704 two_stage_opamp_dummy_magic_0.Vb1.t15 GNDA 0.019408f
C1705 two_stage_opamp_dummy_magic_0.Vb1.t18 GNDA 0.025174f
C1706 two_stage_opamp_dummy_magic_0.Vb1.n3 GNDA 0.027371f
C1707 two_stage_opamp_dummy_magic_0.Vb1.n4 GNDA 0.018462f
C1708 two_stage_opamp_dummy_magic_0.Vb1.n5 GNDA 0.018462f
C1709 two_stage_opamp_dummy_magic_0.Vb1.n6 GNDA 0.015993f
C1710 two_stage_opamp_dummy_magic_0.Vb1.t11 GNDA 0.019408f
C1711 two_stage_opamp_dummy_magic_0.Vb1.t23 GNDA 0.019408f
C1712 two_stage_opamp_dummy_magic_0.Vb1.t12 GNDA 0.019408f
C1713 two_stage_opamp_dummy_magic_0.Vb1.t25 GNDA 0.019408f
C1714 two_stage_opamp_dummy_magic_0.Vb1.t14 GNDA 0.025174f
C1715 two_stage_opamp_dummy_magic_0.Vb1.n7 GNDA 0.027371f
C1716 two_stage_opamp_dummy_magic_0.Vb1.n8 GNDA 0.018462f
C1717 two_stage_opamp_dummy_magic_0.Vb1.n9 GNDA 0.018462f
C1718 two_stage_opamp_dummy_magic_0.Vb1.n10 GNDA 0.015993f
C1719 two_stage_opamp_dummy_magic_0.Vb1.n11 GNDA 0.021438f
C1720 two_stage_opamp_dummy_magic_0.Vb1.t22 GNDA 0.019408f
C1721 two_stage_opamp_dummy_magic_0.Vb1.t10 GNDA 0.019408f
C1722 two_stage_opamp_dummy_magic_0.Vb1.t20 GNDA 0.019408f
C1723 two_stage_opamp_dummy_magic_0.Vb1.t8 GNDA 0.019408f
C1724 two_stage_opamp_dummy_magic_0.Vb1.t17 GNDA 0.025174f
C1725 two_stage_opamp_dummy_magic_0.Vb1.n12 GNDA 0.027371f
C1726 two_stage_opamp_dummy_magic_0.Vb1.n13 GNDA 0.018462f
C1727 two_stage_opamp_dummy_magic_0.Vb1.n14 GNDA 0.018462f
C1728 two_stage_opamp_dummy_magic_0.Vb1.n15 GNDA 0.015993f
C1729 two_stage_opamp_dummy_magic_0.Vb1.t16 GNDA 0.019408f
C1730 two_stage_opamp_dummy_magic_0.Vb1.t7 GNDA 0.019408f
C1731 two_stage_opamp_dummy_magic_0.Vb1.t19 GNDA 0.019408f
C1732 two_stage_opamp_dummy_magic_0.Vb1.t24 GNDA 0.019408f
C1733 two_stage_opamp_dummy_magic_0.Vb1.t13 GNDA 0.025174f
C1734 two_stage_opamp_dummy_magic_0.Vb1.n16 GNDA 0.027371f
C1735 two_stage_opamp_dummy_magic_0.Vb1.n17 GNDA 0.018462f
C1736 two_stage_opamp_dummy_magic_0.Vb1.n18 GNDA 0.018462f
C1737 two_stage_opamp_dummy_magic_0.Vb1.n19 GNDA 0.015993f
C1738 two_stage_opamp_dummy_magic_0.Vb1.n20 GNDA 0.01797f
C1739 two_stage_opamp_dummy_magic_0.Vb1.n21 GNDA 0.525851f
C1740 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA 0.057793f
C1741 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA 0.365115f
C1742 two_stage_opamp_dummy_magic_0.Vb1.n22 GNDA 0.299393f
C1743 two_stage_opamp_dummy_magic_0.Vb1.n23 GNDA 1.74677f
C1744 bgr_0.VB1_CUR_BIAS GNDA 1.32307f
C1745 bgr_0.V_mir2.t9 GNDA 0.03537f
C1746 bgr_0.V_mir2.t1 GNDA 0.03537f
C1747 bgr_0.V_mir2.t5 GNDA 0.03537f
C1748 bgr_0.V_mir2.n0 GNDA 0.08097f
C1749 bgr_0.V_mir2.t0 GNDA 0.042444f
C1750 bgr_0.V_mir2.t17 GNDA 0.042444f
C1751 bgr_0.V_mir2.t20 GNDA 0.06851f
C1752 bgr_0.V_mir2.n1 GNDA 0.076506f
C1753 bgr_0.V_mir2.n2 GNDA 0.052264f
C1754 bgr_0.V_mir2.t4 GNDA 0.053881f
C1755 bgr_0.V_mir2.n3 GNDA 0.081315f
C1756 bgr_0.V_mir2.n4 GNDA 0.203577f
C1757 bgr_0.V_mir2.t7 GNDA 0.03537f
C1758 bgr_0.V_mir2.t3 GNDA 0.03537f
C1759 bgr_0.V_mir2.n5 GNDA 0.08097f
C1760 bgr_0.V_mir2.t6 GNDA 0.042444f
C1761 bgr_0.V_mir2.t18 GNDA 0.042444f
C1762 bgr_0.V_mir2.t21 GNDA 0.06851f
C1763 bgr_0.V_mir2.n6 GNDA 0.076506f
C1764 bgr_0.V_mir2.n7 GNDA 0.052264f
C1765 bgr_0.V_mir2.t2 GNDA 0.053881f
C1766 bgr_0.V_mir2.n8 GNDA 0.081315f
C1767 bgr_0.V_mir2.n9 GNDA 0.156007f
C1768 bgr_0.V_mir2.t14 GNDA 0.017685f
C1769 bgr_0.V_mir2.t15 GNDA 0.017685f
C1770 bgr_0.V_mir2.n10 GNDA 0.046242f
C1771 bgr_0.V_mir2.t13 GNDA 0.075466f
C1772 bgr_0.V_mir2.t12 GNDA 0.017685f
C1773 bgr_0.V_mir2.t16 GNDA 0.017685f
C1774 bgr_0.V_mir2.n11 GNDA 0.050199f
C1775 bgr_0.V_mir2.n12 GNDA 0.827814f
C1776 bgr_0.V_mir2.n13 GNDA 0.268286f
C1777 bgr_0.V_mir2.n14 GNDA 0.09373f
C1778 bgr_0.V_mir2.n15 GNDA 0.699157f
C1779 bgr_0.V_mir2.t8 GNDA 0.042444f
C1780 bgr_0.V_mir2.t19 GNDA 0.042444f
C1781 bgr_0.V_mir2.t22 GNDA 0.06851f
C1782 bgr_0.V_mir2.n16 GNDA 0.076506f
C1783 bgr_0.V_mir2.n17 GNDA 0.052264f
C1784 bgr_0.V_mir2.t10 GNDA 0.053881f
C1785 bgr_0.V_mir2.n18 GNDA 0.081315f
C1786 bgr_0.V_mir2.n19 GNDA 0.201563f
C1787 bgr_0.V_mir2.n20 GNDA 0.08097f
C1788 bgr_0.V_mir2.t11 GNDA 0.03537f
C1789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.065996f
C1790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.024678f
C1791 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.077404f
C1792 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.024678f
C1793 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.063363f
C1794 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.024678f
C1795 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.063363f
C1796 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.024678f
C1797 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.09721f
C1798 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.630211f
C1799 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.080037f
C1800 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.080037f
C1801 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.268206f
C1802 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 3.02207f
C1803 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.080037f
C1804 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.080037f
C1805 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.268206f
C1806 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.724255f
C1807 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.080037f
C1808 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.080037f
C1809 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.268206f
C1810 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.03545f
C1811 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.900713f
C1812 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.012115f
C1813 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.022607f
C1814 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.053973f
C1815 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.292984f
C1816 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.012115f
C1817 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.022607f
C1818 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.053973f
C1819 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.1885f
C1820 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.038199f
C1821 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.30356f
C1822 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.012115f
C1823 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.022607f
C1824 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.053973f
C1825 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.311758f
C1826 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.012115f
C1827 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.022607f
C1828 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.053973f
C1829 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.1885f
C1830 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.038199f
C1831 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 GNDA 1.63304f
C1832 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.016017f
C1833 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.016625f
C1834 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.016536f
C1835 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.112284f
C1836 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.016625f
C1837 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.073697f
C1838 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.171055f
C1839 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.017683f
C1840 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.017683f
C1841 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.017683f
C1842 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.017683f
C1843 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.017683f
C1844 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.017683f
C1845 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.017683f
C1846 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.020638f
C1847 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.019459f
C1848 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.012203f
C1849 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.012203f
C1850 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.012203f
C1851 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.012203f
C1852 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.012203f
C1853 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.010905f
C1854 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.017683f
C1855 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.017683f
C1856 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.017683f
C1857 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.017683f
C1858 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.017683f
C1859 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.017683f
C1860 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.017683f
C1861 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.017683f
C1862 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.017683f
C1863 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.017683f
C1864 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.017683f
C1865 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.020638f
C1866 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.019459f
C1867 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.012203f
C1868 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.012203f
C1869 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.012203f
C1870 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.012203f
C1871 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.012203f
C1872 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.012203f
C1873 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.012203f
C1874 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.012203f
C1875 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.012203f
C1876 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.010905f
C1877 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.027252f
C1878 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.019924f
C1879 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.077697f
C1880 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.035725f
C1881 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.806182f
C1882 bgr_0.TAIL_CUR_MIR_BIAS GNDA 0.826265f
C1883 VDDA.t472 GNDA 0.70711f
C1884 VDDA.t470 GNDA 0.753644f
C1885 VDDA.t469 GNDA 0.753644f
C1886 VDDA.t471 GNDA 0.722682f
C1887 VDDA.n0 GNDA 0.505164f
C1888 VDDA.n1 GNDA 0.245259f
C1889 VDDA.n2 GNDA 0.314438f
C1890 VDDA.n3 GNDA 2.53346f
C1891 VDDA.n4 GNDA 0.020467f
C1892 VDDA.n5 GNDA 0.015491f
C1893 VDDA.n6 GNDA 0.015491f
C1894 VDDA.n7 GNDA 0.045271f
C1895 VDDA.n8 GNDA 0.020467f
C1896 VDDA.t87 GNDA 0.024027f
C1897 VDDA.t85 GNDA 0.015833f
C1898 VDDA.n9 GNDA 0.037692f
C1899 VDDA.n10 GNDA 0.053632f
C1900 VDDA.n11 GNDA 0.100825f
C1901 VDDA.n12 GNDA 0.100825f
C1902 VDDA.n13 GNDA 0.020467f
C1903 VDDA.n14 GNDA 0.015491f
C1904 VDDA.n15 GNDA 0.016197f
C1905 VDDA.n16 GNDA 0.016087f
C1906 VDDA.n17 GNDA 0.125058f
C1907 VDDA.n18 GNDA 0.016087f
C1908 VDDA.n19 GNDA 0.065142f
C1909 VDDA.n20 GNDA 0.016087f
C1910 VDDA.n21 GNDA 0.065142f
C1911 VDDA.n22 GNDA 0.062915f
C1912 VDDA.n23 GNDA 0.100825f
C1913 VDDA.t14 GNDA 0.024027f
C1914 VDDA.t12 GNDA 0.015833f
C1915 VDDA.n24 GNDA 0.037692f
C1916 VDDA.n25 GNDA 0.053632f
C1917 VDDA.t53 GNDA 0.024027f
C1918 VDDA.t51 GNDA 0.015833f
C1919 VDDA.n26 GNDA 0.037692f
C1920 VDDA.n27 GNDA 0.053632f
C1921 VDDA.n28 GNDA 0.076753f
C1922 VDDA.n29 GNDA 0.100825f
C1923 VDDA.n30 GNDA 0.219223f
C1924 VDDA.t52 GNDA 0.19995f
C1925 VDDA.t268 GNDA 0.126642f
C1926 VDDA.t312 GNDA 0.126642f
C1927 VDDA.t314 GNDA 0.126642f
C1928 VDDA.t448 GNDA 0.126642f
C1929 VDDA.t296 GNDA 0.126642f
C1930 VDDA.t205 GNDA 0.126642f
C1931 VDDA.t270 GNDA 0.126642f
C1932 VDDA.t199 GNDA 0.126642f
C1933 VDDA.t260 GNDA 0.094981f
C1934 VDDA.n31 GNDA 0.063321f
C1935 VDDA.t290 GNDA 0.094981f
C1936 VDDA.t431 GNDA 0.126642f
C1937 VDDA.t238 GNDA 0.126642f
C1938 VDDA.t203 GNDA 0.126642f
C1939 VDDA.t461 GNDA 0.126642f
C1940 VDDA.t429 GNDA 0.126642f
C1941 VDDA.t279 GNDA 0.126642f
C1942 VDDA.t248 GNDA 0.126642f
C1943 VDDA.t272 GNDA 0.126642f
C1944 VDDA.t13 GNDA 0.19995f
C1945 VDDA.n32 GNDA 0.219223f
C1946 VDDA.n33 GNDA 0.062915f
C1947 VDDA.n34 GNDA 0.107177f
C1948 VDDA.n35 GNDA 0.015491f
C1949 VDDA.n36 GNDA 0.045271f
C1950 VDDA.n37 GNDA 0.020467f
C1951 VDDA.n38 GNDA 0.016087f
C1952 VDDA.n39 GNDA 0.065142f
C1953 VDDA.n40 GNDA 0.016087f
C1954 VDDA.n41 GNDA 0.065142f
C1955 VDDA.n42 GNDA 0.016087f
C1956 VDDA.n43 GNDA 0.065142f
C1957 VDDA.n44 GNDA 0.016087f
C1958 VDDA.n45 GNDA 0.093285f
C1959 VDDA.n46 GNDA 0.020467f
C1960 VDDA.n47 GNDA 0.015491f
C1961 VDDA.n48 GNDA 0.015491f
C1962 VDDA.n49 GNDA 0.045271f
C1963 VDDA.n50 GNDA 0.020467f
C1964 VDDA.n51 GNDA 0.020467f
C1965 VDDA.n52 GNDA 0.015491f
C1966 VDDA.n53 GNDA 0.045271f
C1967 VDDA.n54 GNDA 0.020467f
C1968 VDDA.n55 GNDA 0.020467f
C1969 VDDA.n56 GNDA 0.015491f
C1970 VDDA.n57 GNDA 0.045271f
C1971 VDDA.n58 GNDA 0.020467f
C1972 VDDA.n59 GNDA 0.020467f
C1973 VDDA.n60 GNDA 0.015491f
C1974 VDDA.n61 GNDA 0.045271f
C1975 VDDA.n62 GNDA 0.020467f
C1976 VDDA.n63 GNDA 0.020467f
C1977 VDDA.n64 GNDA 0.045271f
C1978 VDDA.n65 GNDA 0.020467f
C1979 VDDA.n66 GNDA 0.015491f
C1980 VDDA.n67 GNDA 0.045271f
C1981 VDDA.n68 GNDA 0.020467f
C1982 VDDA.n69 GNDA 0.04861f
C1983 VDDA.n70 GNDA 0.045271f
C1984 VDDA.n71 GNDA 0.033417f
C1985 VDDA.t117 GNDA 0.024027f
C1986 VDDA.t115 GNDA 0.015833f
C1987 VDDA.n72 GNDA 0.037692f
C1988 VDDA.n73 GNDA 0.076753f
C1989 VDDA.n74 GNDA 0.053632f
C1990 VDDA.n75 GNDA 0.031918f
C1991 VDDA.n76 GNDA 0.219223f
C1992 VDDA.t116 GNDA 0.19995f
C1993 VDDA.t441 GNDA 0.126642f
C1994 VDDA.t134 GNDA 0.126642f
C1995 VDDA.t343 GNDA 0.126642f
C1996 VDDA.t120 GNDA 0.126642f
C1997 VDDA.t422 GNDA 0.126642f
C1998 VDDA.t254 GNDA 0.126642f
C1999 VDDA.t439 GNDA 0.126642f
C2000 VDDA.t132 GNDA 0.126642f
C2001 VDDA.t341 GNDA 0.094981f
C2002 VDDA.n77 GNDA 0.063321f
C2003 VDDA.t118 GNDA 0.094981f
C2004 VDDA.t236 GNDA 0.126642f
C2005 VDDA.t252 GNDA 0.126642f
C2006 VDDA.t437 GNDA 0.126642f
C2007 VDDA.t345 GNDA 0.126642f
C2008 VDDA.t338 GNDA 0.126642f
C2009 VDDA.t234 GNDA 0.126642f
C2010 VDDA.t242 GNDA 0.126642f
C2011 VDDA.t250 GNDA 0.126642f
C2012 VDDA.t86 GNDA 0.19995f
C2013 VDDA.n78 GNDA 0.219223f
C2014 VDDA.n79 GNDA 0.031918f
C2015 VDDA.n80 GNDA 0.033417f
C2016 VDDA.n81 GNDA 0.045271f
C2017 VDDA.n82 GNDA 0.061963f
C2018 VDDA.n83 GNDA 0.188123f
C2019 VDDA.t300 GNDA 0.019188f
C2020 VDDA.t293 GNDA 0.019188f
C2021 VDDA.n84 GNDA 0.063392f
C2022 VDDA.n85 GNDA 0.081799f
C2023 VDDA.n86 GNDA 0.103616f
C2024 VDDA.n87 GNDA 0.141248f
C2025 VDDA.n88 GNDA 0.140599f
C2026 VDDA.n89 GNDA 0.141248f
C2027 VDDA.t60 GNDA 0.091497f
C2028 VDDA.t62 GNDA 0.058804f
C2029 VDDA.t108 GNDA 0.024027f
C2030 VDDA.t106 GNDA 0.012125f
C2031 VDDA.n90 GNDA 0.037882f
C2032 VDDA.n91 GNDA 0.021843f
C2033 VDDA.n92 GNDA 0.038821f
C2034 VDDA.t26 GNDA 0.024027f
C2035 VDDA.t24 GNDA 0.012125f
C2036 VDDA.n93 GNDA 0.037882f
C2037 VDDA.n94 GNDA 0.038821f
C2038 VDDA.n95 GNDA 0.038821f
C2039 VDDA.n96 GNDA 0.031853f
C2040 VDDA.n97 GNDA 0.153065f
C2041 VDDA.t107 GNDA 0.192197f
C2042 VDDA.t282 GNDA 0.087066f
C2043 VDDA.n98 GNDA 0.058044f
C2044 VDDA.t281 GNDA 0.087066f
C2045 VDDA.t25 GNDA 0.195031f
C2046 VDDA.n99 GNDA 0.160784f
C2047 VDDA.n100 GNDA 0.031853f
C2048 VDDA.n101 GNDA 0.021843f
C2049 VDDA.n102 GNDA 0.030687f
C2050 VDDA.t444 GNDA 0.019188f
C2051 VDDA.t198 GNDA 0.019188f
C2052 VDDA.n103 GNDA 0.063392f
C2053 VDDA.n104 GNDA 0.081799f
C2054 VDDA.t222 GNDA 0.019188f
C2055 VDDA.t225 GNDA 0.019188f
C2056 VDDA.n105 GNDA 0.063392f
C2057 VDDA.n106 GNDA 0.081799f
C2058 VDDA.t142 GNDA 0.019188f
C2059 VDDA.t179 GNDA 0.019188f
C2060 VDDA.n107 GNDA 0.063392f
C2061 VDDA.n108 GNDA 0.081799f
C2062 VDDA.t182 GNDA 0.019188f
C2063 VDDA.t308 GNDA 0.019188f
C2064 VDDA.n109 GNDA 0.063392f
C2065 VDDA.n110 GNDA 0.081799f
C2066 VDDA.t209 GNDA 0.019188f
C2067 VDDA.t241 GNDA 0.019188f
C2068 VDDA.n111 GNDA 0.063392f
C2069 VDDA.n112 GNDA 0.081799f
C2070 VDDA.t245 GNDA 0.019188f
C2071 VDDA.t451 GNDA 0.019188f
C2072 VDDA.n113 GNDA 0.063392f
C2073 VDDA.n114 GNDA 0.081799f
C2074 VDDA.t196 GNDA 0.019188f
C2075 VDDA.t295 GNDA 0.019188f
C2076 VDDA.n115 GNDA 0.063392f
C2077 VDDA.n116 GNDA 0.081799f
C2078 VDDA.n117 GNDA 0.090315f
C2079 VDDA.n118 GNDA 0.109198f
C2080 VDDA.n119 GNDA 0.073605f
C2081 VDDA.n120 GNDA 0.089866f
C2082 VDDA.n121 GNDA 0.331114f
C2083 VDDA.t61 GNDA 0.427247f
C2084 VDDA.t195 GNDA 0.30797f
C2085 VDDA.t294 GNDA 0.30797f
C2086 VDDA.t244 GNDA 0.30797f
C2087 VDDA.t450 GNDA 0.30797f
C2088 VDDA.t208 GNDA 0.30797f
C2089 VDDA.t240 GNDA 0.30797f
C2090 VDDA.t181 GNDA 0.30797f
C2091 VDDA.t307 GNDA 0.230977f
C2092 VDDA.n122 GNDA 0.153985f
C2093 VDDA.t141 GNDA 0.230977f
C2094 VDDA.t178 GNDA 0.30797f
C2095 VDDA.t221 GNDA 0.30797f
C2096 VDDA.t224 GNDA 0.30797f
C2097 VDDA.t443 GNDA 0.30797f
C2098 VDDA.t197 GNDA 0.30797f
C2099 VDDA.t299 GNDA 0.30797f
C2100 VDDA.t292 GNDA 0.30797f
C2101 VDDA.t46 GNDA 0.427247f
C2102 VDDA.n123 GNDA 0.331114f
C2103 VDDA.n124 GNDA 0.089866f
C2104 VDDA.n125 GNDA 0.073605f
C2105 VDDA.t47 GNDA 0.058804f
C2106 VDDA.t45 GNDA 0.091497f
C2107 VDDA.n126 GNDA 0.109198f
C2108 VDDA.n127 GNDA 0.050127f
C2109 VDDA.t99 GNDA 0.024206f
C2110 VDDA.t97 GNDA 0.011812f
C2111 VDDA.n128 GNDA 0.036258f
C2112 VDDA.n129 GNDA 0.021743f
C2113 VDDA.n130 GNDA 0.038821f
C2114 VDDA.t111 GNDA 0.024206f
C2115 VDDA.t109 GNDA 0.011812f
C2116 VDDA.n131 GNDA 0.036258f
C2117 VDDA.n132 GNDA 0.038821f
C2118 VDDA.n133 GNDA 0.038821f
C2119 VDDA.n134 GNDA 0.031853f
C2120 VDDA.n135 GNDA 0.153065f
C2121 VDDA.t98 GNDA 0.192197f
C2122 VDDA.t414 GNDA 0.087066f
C2123 VDDA.n136 GNDA 0.058044f
C2124 VDDA.t396 GNDA 0.087066f
C2125 VDDA.t110 GNDA 0.192197f
C2126 VDDA.n137 GNDA 0.153065f
C2127 VDDA.n138 GNDA 0.031853f
C2128 VDDA.n139 GNDA 0.021743f
C2129 VDDA.n140 GNDA 0.022843f
C2130 VDDA.n141 GNDA 0.015447f
C2131 VDDA.n142 GNDA 0.042757f
C2132 VDDA.n143 GNDA 0.090084f
C2133 VDDA.n144 GNDA 0.156428f
C2134 VDDA.n145 GNDA 0.015955f
C2135 VDDA.n146 GNDA 0.05632f
C2136 VDDA.n147 GNDA 0.021107f
C2137 VDDA.n148 GNDA 0.045687f
C2138 VDDA.n149 GNDA 0.045686f
C2139 VDDA.n150 GNDA 0.045687f
C2140 VDDA.t15 GNDA 0.012596f
C2141 VDDA.t17 GNDA 0.025242f
C2142 VDDA.n151 GNDA 0.015925f
C2143 VDDA.n152 GNDA 0.05635f
C2144 VDDA.n153 GNDA 0.042214f
C2145 VDDA.n154 GNDA 0.066507f
C2146 VDDA.n155 GNDA 0.066507f
C2147 VDDA.n156 GNDA 0.066507f
C2148 VDDA.t82 GNDA 0.012596f
C2149 VDDA.t84 GNDA 0.024089f
C2150 VDDA.n157 GNDA 0.015962f
C2151 VDDA.n158 GNDA 0.056314f
C2152 VDDA.n159 GNDA 0.021107f
C2153 VDDA.n160 GNDA 0.045686f
C2154 VDDA.n161 GNDA 0.045686f
C2155 VDDA.n162 GNDA 0.045686f
C2156 VDDA.t79 GNDA 0.012596f
C2157 VDDA.t81 GNDA 0.025252f
C2158 VDDA.n163 GNDA 0.015962f
C2159 VDDA.n164 GNDA 0.077075f
C2160 VDDA.n165 GNDA 0.043247f
C2161 VDDA.n166 GNDA 0.025809f
C2162 VDDA.n167 GNDA 0.035456f
C2163 VDDA.n168 GNDA 0.161528f
C2164 VDDA.t80 GNDA 0.195577f
C2165 VDDA.t378 GNDA 0.117847f
C2166 VDDA.t400 GNDA 0.088385f
C2167 VDDA.n169 GNDA 0.058924f
C2168 VDDA.t412 GNDA 0.088385f
C2169 VDDA.t394 GNDA 0.117847f
C2170 VDDA.t104 GNDA 0.195577f
C2171 VDDA.n170 GNDA 0.161528f
C2172 VDDA.n171 GNDA 0.035456f
C2173 VDDA.n172 GNDA 0.025809f
C2174 VDDA.t105 GNDA 0.025252f
C2175 VDDA.t103 GNDA 0.012996f
C2176 VDDA.n173 GNDA 0.042801f
C2177 VDDA.n174 GNDA 0.038877f
C2178 VDDA.n175 GNDA 0.015925f
C2179 VDDA.n176 GNDA 0.05635f
C2180 VDDA.n177 GNDA 0.015925f
C2181 VDDA.n178 GNDA 0.05635f
C2182 VDDA.n179 GNDA 0.015925f
C2183 VDDA.n180 GNDA 0.05635f
C2184 VDDA.n181 GNDA 0.015925f
C2185 VDDA.n182 GNDA 0.05635f
C2186 VDDA.n183 GNDA 0.038877f
C2187 VDDA.n184 GNDA 0.043565f
C2188 VDDA.n185 GNDA 0.03988f
C2189 VDDA.n186 GNDA 0.049704f
C2190 VDDA.n187 GNDA 0.190023f
C2191 VDDA.t83 GNDA 0.195577f
C2192 VDDA.t382 GNDA 0.117847f
C2193 VDDA.t386 GNDA 0.117847f
C2194 VDDA.t406 GNDA 0.117847f
C2195 VDDA.t384 GNDA 0.117847f
C2196 VDDA.t416 GNDA 0.117847f
C2197 VDDA.t398 GNDA 0.088385f
C2198 VDDA.n188 GNDA 0.058924f
C2199 VDDA.t410 GNDA 0.088385f
C2200 VDDA.t392 GNDA 0.117847f
C2201 VDDA.t408 GNDA 0.117847f
C2202 VDDA.t388 GNDA 0.117847f
C2203 VDDA.t64 GNDA 0.195577f
C2204 VDDA.n189 GNDA 0.175818f
C2205 VDDA.n190 GNDA 0.042601f
C2206 VDDA.n191 GNDA 0.032845f
C2207 VDDA.t65 GNDA 0.024089f
C2208 VDDA.t63 GNDA 0.012596f
C2209 VDDA.n192 GNDA 0.043565f
C2210 VDDA.n193 GNDA 0.045912f
C2211 VDDA.n194 GNDA 0.015955f
C2212 VDDA.n195 GNDA 0.05632f
C2213 VDDA.n196 GNDA 0.045912f
C2214 VDDA.n197 GNDA 0.042411f
C2215 VDDA.n198 GNDA 0.025809f
C2216 VDDA.n199 GNDA 0.034966f
C2217 VDDA.n200 GNDA 0.159782f
C2218 VDDA.t16 GNDA 0.192197f
C2219 VDDA.t404 GNDA 0.116088f
C2220 VDDA.t380 GNDA 0.079151f
C2221 VDDA.n201 GNDA 0.029022f
C2222 VDDA.n202 GNDA 0.036937f
C2223 VDDA.t402 GNDA 0.087066f
C2224 VDDA.t390 GNDA 0.116088f
C2225 VDDA.t95 GNDA 0.192197f
C2226 VDDA.n203 GNDA 0.160761f
C2227 VDDA.n204 GNDA 0.035945f
C2228 VDDA.n205 GNDA 0.025809f
C2229 VDDA.t96 GNDA 0.025242f
C2230 VDDA.t94 GNDA 0.012596f
C2231 VDDA.n206 GNDA 0.042411f
C2232 VDDA.n207 GNDA 0.084591f
C2233 VDDA.n208 GNDA 0.126979f
C2234 VDDA.t445 GNDA 0.357539f
C2235 VDDA.t298 GNDA 0.358835f
C2236 VDDA.t289 GNDA 0.357539f
C2237 VDDA.t183 GNDA 0.358835f
C2238 VDDA.t246 GNDA 0.357539f
C2239 VDDA.t143 GNDA 0.358835f
C2240 VDDA.t139 GNDA 0.357539f
C2241 VDDA.t180 GNDA 0.358835f
C2242 VDDA.t223 GNDA 0.357539f
C2243 VDDA.t247 GNDA 0.358835f
C2244 VDDA.t274 GNDA 0.357539f
C2245 VDDA.t452 GNDA 0.358835f
C2246 VDDA.t288 GNDA 0.357539f
C2247 VDDA.t306 GNDA 0.358835f
C2248 VDDA.t140 GNDA 0.357539f
C2249 VDDA.t275 GNDA 0.358835f
C2250 VDDA.n209 GNDA 0.239659f
C2251 VDDA.t257 GNDA 0.190853f
C2252 VDDA.n210 GNDA 0.260035f
C2253 VDDA.t207 GNDA 0.190853f
C2254 VDDA.n211 GNDA 0.260035f
C2255 VDDA.t256 GNDA 0.190853f
C2256 VDDA.n212 GNDA 0.260035f
C2257 VDDA.t226 GNDA 0.284791f
C2258 VDDA.n213 GNDA 0.24816f
C2259 VDDA.n214 GNDA 3.00103f
C2260 VDDA.t317 GNDA 0.019188f
C2261 VDDA.t232 GNDA 0.019188f
C2262 VDDA.n215 GNDA 0.079352f
C2263 VDDA.t175 GNDA 0.019188f
C2264 VDDA.t161 GNDA 0.019188f
C2265 VDDA.n216 GNDA 0.079048f
C2266 VDDA.n217 GNDA 0.109595f
C2267 VDDA.t176 GNDA 0.019188f
C2268 VDDA.t201 GNDA 0.019188f
C2269 VDDA.n218 GNDA 0.079048f
C2270 VDDA.n219 GNDA 0.057188f
C2271 VDDA.t428 GNDA 0.019188f
C2272 VDDA.t138 GNDA 0.019188f
C2273 VDDA.n220 GNDA 0.079048f
C2274 VDDA.n221 GNDA 0.057188f
C2275 VDDA.t427 GNDA 0.019188f
C2276 VDDA.t287 GNDA 0.019188f
C2277 VDDA.n222 GNDA 0.079048f
C2278 VDDA.n223 GNDA 0.057188f
C2279 VDDA.t230 GNDA 0.019188f
C2280 VDDA.t286 GNDA 0.019188f
C2281 VDDA.n224 GNDA 0.079048f
C2282 VDDA.n225 GNDA 0.165166f
C2283 VDDA.t323 GNDA 0.038376f
C2284 VDDA.t212 GNDA 0.038376f
C2285 VDDA.n226 GNDA 0.153961f
C2286 VDDA.n227 GNDA 0.078216f
C2287 VDDA.t68 GNDA 0.038229f
C2288 VDDA.n228 GNDA 0.051766f
C2289 VDDA.n229 GNDA 0.073068f
C2290 VDDA.t75 GNDA 0.042458f
C2291 VDDA.t73 GNDA 0.018593f
C2292 VDDA.n230 GNDA 0.06735f
C2293 VDDA.n231 GNDA 0.039649f
C2294 VDDA.t56 GNDA 0.042458f
C2295 VDDA.t54 GNDA 0.018593f
C2296 VDDA.n232 GNDA 0.06735f
C2297 VDDA.n233 GNDA 0.039649f
C2298 VDDA.n234 GNDA 0.042214f
C2299 VDDA.n235 GNDA 0.073068f
C2300 VDDA.n236 GNDA 0.211231f
C2301 VDDA.t55 GNDA 0.261604f
C2302 VDDA.t146 GNDA 0.151267f
C2303 VDDA.t466 GNDA 0.151267f
C2304 VDDA.t324 GNDA 0.151267f
C2305 VDDA.t367 GNDA 0.151267f
C2306 VDDA.t210 GNDA 0.11345f
C2307 VDDA.n237 GNDA 0.075633f
C2308 VDDA.t368 GNDA 0.11345f
C2309 VDDA.t327 GNDA 0.151267f
C2310 VDDA.t144 GNDA 0.151267f
C2311 VDDA.t326 GNDA 0.151267f
C2312 VDDA.t145 GNDA 0.151267f
C2313 VDDA.t74 GNDA 0.261604f
C2314 VDDA.n238 GNDA 0.211231f
C2315 VDDA.n239 GNDA 0.051766f
C2316 VDDA.n240 GNDA 0.097957f
C2317 VDDA.n241 GNDA 0.067039f
C2318 VDDA.n242 GNDA 0.099438f
C2319 VDDA.n243 GNDA 0.099438f
C2320 VDDA.n244 GNDA 0.09879f
C2321 VDDA.t44 GNDA 0.038229f
C2322 VDDA.t321 GNDA 0.038376f
C2323 VDDA.t460 GNDA 0.038376f
C2324 VDDA.n245 GNDA 0.153961f
C2325 VDDA.n246 GNDA 0.078216f
C2326 VDDA.t302 GNDA 0.038376f
C2327 VDDA.t455 GNDA 0.038376f
C2328 VDDA.n247 GNDA 0.153961f
C2329 VDDA.n248 GNDA 0.078216f
C2330 VDDA.t468 GNDA 0.038376f
C2331 VDDA.t458 GNDA 0.038376f
C2332 VDDA.n249 GNDA 0.153961f
C2333 VDDA.n250 GNDA 0.078216f
C2334 VDDA.t1 GNDA 0.038376f
C2335 VDDA.t304 GNDA 0.038376f
C2336 VDDA.n251 GNDA 0.153961f
C2337 VDDA.n252 GNDA 0.164359f
C2338 VDDA.n253 GNDA 0.124094f
C2339 VDDA.t42 GNDA 0.046386f
C2340 VDDA.n254 GNDA 0.08875f
C2341 VDDA.n255 GNDA 0.05185f
C2342 VDDA.n256 GNDA 0.07758f
C2343 VDDA.n257 GNDA 0.341479f
C2344 VDDA.t43 GNDA 0.527449f
C2345 VDDA.t0 GNDA 0.29198f
C2346 VDDA.t303 GNDA 0.29198f
C2347 VDDA.t467 GNDA 0.29198f
C2348 VDDA.t457 GNDA 0.29198f
C2349 VDDA.t301 GNDA 0.218985f
C2350 VDDA.n258 GNDA 0.14599f
C2351 VDDA.t454 GNDA 0.218985f
C2352 VDDA.t320 GNDA 0.29198f
C2353 VDDA.t459 GNDA 0.29198f
C2354 VDDA.t322 GNDA 0.29198f
C2355 VDDA.t211 GNDA 0.29198f
C2356 VDDA.t67 GNDA 0.527449f
C2357 VDDA.n259 GNDA 0.341479f
C2358 VDDA.n260 GNDA 0.07758f
C2359 VDDA.n261 GNDA 0.05185f
C2360 VDDA.t66 GNDA 0.046386f
C2361 VDDA.n262 GNDA 0.08875f
C2362 VDDA.n263 GNDA 0.123774f
C2363 VDDA.n264 GNDA 0.09286f
C2364 VDDA.t231 GNDA 0.019188f
C2365 VDDA.t267 GNDA 0.019188f
C2366 VDDA.n265 GNDA 0.079352f
C2367 VDDA.t309 GNDA 0.019188f
C2368 VDDA.t456 GNDA 0.019188f
C2369 VDDA.n266 GNDA 0.079048f
C2370 VDDA.n267 GNDA 0.109595f
C2371 VDDA.t328 GNDA 0.019188f
C2372 VDDA.t311 GNDA 0.019188f
C2373 VDDA.n268 GNDA 0.079048f
C2374 VDDA.n269 GNDA 0.057188f
C2375 VDDA.t463 GNDA 0.019188f
C2376 VDDA.t325 GNDA 0.019188f
C2377 VDDA.n270 GNDA 0.079048f
C2378 VDDA.n271 GNDA 0.057188f
C2379 VDDA.t453 GNDA 0.019188f
C2380 VDDA.t310 GNDA 0.019188f
C2381 VDDA.n272 GNDA 0.079048f
C2382 VDDA.n273 GNDA 0.057188f
C2383 VDDA.t278 GNDA 0.019188f
C2384 VDDA.t233 GNDA 0.019188f
C2385 VDDA.n274 GNDA 0.079048f
C2386 VDDA.n275 GNDA 0.19758f
C2387 VDDA.n276 GNDA 0.182609f
C2388 VDDA.t370 GNDA 0.022386f
C2389 VDDA.t435 GNDA 0.022386f
C2390 VDDA.n277 GNDA 0.077854f
C2391 VDDA.t154 GNDA 0.022386f
C2392 VDDA.t465 GNDA 0.022386f
C2393 VDDA.n278 GNDA 0.077578f
C2394 VDDA.n279 GNDA 0.146461f
C2395 VDDA.t150 GNDA 0.022386f
C2396 VDDA.t152 GNDA 0.022386f
C2397 VDDA.n280 GNDA 0.077854f
C2398 VDDA.t336 GNDA 0.022386f
C2399 VDDA.t377 GNDA 0.022386f
C2400 VDDA.n281 GNDA 0.077578f
C2401 VDDA.n282 GNDA 0.146461f
C2402 VDDA.n283 GNDA 0.020467f
C2403 VDDA.n284 GNDA 0.063731f
C2404 VDDA.n285 GNDA 0.086662f
C2405 VDDA.t78 GNDA 0.110436f
C2406 VDDA.t76 GNDA 0.038982f
C2407 VDDA.n286 GNDA 0.072045f
C2408 VDDA.n287 GNDA 0.046444f
C2409 VDDA.t5 GNDA 0.110436f
C2410 VDDA.t3 GNDA 0.038982f
C2411 VDDA.n288 GNDA 0.072045f
C2412 VDDA.n289 GNDA 0.046444f
C2413 VDDA.n290 GNDA 0.046052f
C2414 VDDA.n291 GNDA 0.086662f
C2415 VDDA.n292 GNDA 0.258267f
C2416 VDDA.t4 GNDA 0.3855f
C2417 VDDA.t369 GNDA 0.222583f
C2418 VDDA.t434 GNDA 0.222583f
C2419 VDDA.t153 GNDA 0.222583f
C2420 VDDA.t464 GNDA 0.222583f
C2421 VDDA.t213 GNDA 0.166937f
C2422 VDDA.n293 GNDA 0.111291f
C2423 VDDA.t184 GNDA 0.166937f
C2424 VDDA.t335 GNDA 0.222583f
C2425 VDDA.t376 GNDA 0.222583f
C2426 VDDA.t149 GNDA 0.222583f
C2427 VDDA.t151 GNDA 0.222583f
C2428 VDDA.t77 GNDA 0.3855f
C2429 VDDA.n294 GNDA 0.258267f
C2430 VDDA.n295 GNDA 0.063731f
C2431 VDDA.n296 GNDA 0.08922f
C2432 VDDA.t214 GNDA 0.022386f
C2433 VDDA.t185 GNDA 0.022386f
C2434 VDDA.n297 GNDA 0.072988f
C2435 VDDA.n298 GNDA 0.049816f
C2436 VDDA.n299 GNDA 0.027787f
C2437 VDDA.n300 GNDA 0.111647f
C2438 VDDA.t148 GNDA 0.022386f
C2439 VDDA.t419 GNDA 0.022386f
C2440 VDDA.n301 GNDA 0.077854f
C2441 VDDA.t421 GNDA 0.022386f
C2442 VDDA.t334 GNDA 0.022386f
C2443 VDDA.n302 GNDA 0.077578f
C2444 VDDA.n303 GNDA 0.146461f
C2445 VDDA.t188 GNDA 0.022386f
C2446 VDDA.t447 GNDA 0.022386f
C2447 VDDA.n304 GNDA 0.077854f
C2448 VDDA.t163 GNDA 0.022386f
C2449 VDDA.t172 GNDA 0.022386f
C2450 VDDA.n305 GNDA 0.077578f
C2451 VDDA.n306 GNDA 0.146461f
C2452 VDDA.n307 GNDA 0.020467f
C2453 VDDA.n308 GNDA 0.063731f
C2454 VDDA.n309 GNDA 0.086662f
C2455 VDDA.t20 GNDA 0.110436f
C2456 VDDA.t18 GNDA 0.038982f
C2457 VDDA.n310 GNDA 0.072045f
C2458 VDDA.n311 GNDA 0.046444f
C2459 VDDA.t102 GNDA 0.110436f
C2460 VDDA.t100 GNDA 0.038982f
C2461 VDDA.n312 GNDA 0.072045f
C2462 VDDA.n313 GNDA 0.046444f
C2463 VDDA.n314 GNDA 0.046052f
C2464 VDDA.n315 GNDA 0.086662f
C2465 VDDA.n316 GNDA 0.258267f
C2466 VDDA.t101 GNDA 0.3855f
C2467 VDDA.t147 GNDA 0.222583f
C2468 VDDA.t418 GNDA 0.222583f
C2469 VDDA.t420 GNDA 0.222583f
C2470 VDDA.t333 GNDA 0.222583f
C2471 VDDA.t130 GNDA 0.166937f
C2472 VDDA.n317 GNDA 0.111291f
C2473 VDDA.t374 GNDA 0.166937f
C2474 VDDA.t162 GNDA 0.222583f
C2475 VDDA.t171 GNDA 0.222583f
C2476 VDDA.t187 GNDA 0.222583f
C2477 VDDA.t446 GNDA 0.222583f
C2478 VDDA.t19 GNDA 0.3855f
C2479 VDDA.n318 GNDA 0.258267f
C2480 VDDA.n319 GNDA 0.063731f
C2481 VDDA.n320 GNDA 0.08922f
C2482 VDDA.t131 GNDA 0.022386f
C2483 VDDA.t375 GNDA 0.022386f
C2484 VDDA.n321 GNDA 0.072988f
C2485 VDDA.n322 GNDA 0.049816f
C2486 VDDA.n323 GNDA 0.027787f
C2487 VDDA.n324 GNDA 0.109728f
C2488 VDDA.t125 GNDA 0.038376f
C2489 VDDA.t174 GNDA 0.038376f
C2490 VDDA.n325 GNDA 0.153961f
C2491 VDDA.n326 GNDA 0.078216f
C2492 VDDA.t32 GNDA 0.038229f
C2493 VDDA.n327 GNDA 0.07758f
C2494 VDDA.n328 GNDA 0.051766f
C2495 VDDA.n329 GNDA 0.073068f
C2496 VDDA.t59 GNDA 0.042458f
C2497 VDDA.t57 GNDA 0.018593f
C2498 VDDA.n330 GNDA 0.06735f
C2499 VDDA.n331 GNDA 0.039649f
C2500 VDDA.t35 GNDA 0.042458f
C2501 VDDA.t33 GNDA 0.018593f
C2502 VDDA.n332 GNDA 0.06735f
C2503 VDDA.n333 GNDA 0.039649f
C2504 VDDA.n334 GNDA 0.042214f
C2505 VDDA.n335 GNDA 0.073068f
C2506 VDDA.n336 GNDA 0.211231f
C2507 VDDA.t34 GNDA 0.261604f
C2508 VDDA.t169 GNDA 0.151267f
C2509 VDDA.t177 GNDA 0.151267f
C2510 VDDA.t202 GNDA 0.151267f
C2511 VDDA.t424 GNDA 0.151267f
C2512 VDDA.t170 GNDA 0.11345f
C2513 VDDA.n337 GNDA 0.075633f
C2514 VDDA.t156 GNDA 0.11345f
C2515 VDDA.t316 GNDA 0.151267f
C2516 VDDA.t283 GNDA 0.151267f
C2517 VDDA.t168 GNDA 0.151267f
C2518 VDDA.t266 GNDA 0.151267f
C2519 VDDA.t58 GNDA 0.261604f
C2520 VDDA.n338 GNDA 0.211231f
C2521 VDDA.n339 GNDA 0.051766f
C2522 VDDA.n340 GNDA 0.097957f
C2523 VDDA.t50 GNDA 0.038229f
C2524 VDDA.t160 GNDA 0.038376f
C2525 VDDA.t426 GNDA 0.038376f
C2526 VDDA.n341 GNDA 0.153961f
C2527 VDDA.n342 GNDA 0.078216f
C2528 VDDA.t129 GNDA 0.038376f
C2529 VDDA.t158 GNDA 0.038376f
C2530 VDDA.n343 GNDA 0.153961f
C2531 VDDA.n344 GNDA 0.078216f
C2532 VDDA.t137 GNDA 0.038376f
C2533 VDDA.t285 GNDA 0.038376f
C2534 VDDA.n345 GNDA 0.153961f
C2535 VDDA.n346 GNDA 0.078216f
C2536 VDDA.t123 GNDA 0.038376f
C2537 VDDA.t127 GNDA 0.038376f
C2538 VDDA.n347 GNDA 0.153961f
C2539 VDDA.n348 GNDA 0.164359f
C2540 VDDA.n349 GNDA 0.124094f
C2541 VDDA.t48 GNDA 0.046386f
C2542 VDDA.n350 GNDA 0.08875f
C2543 VDDA.n351 GNDA 0.05185f
C2544 VDDA.n352 GNDA 0.341479f
C2545 VDDA.n353 GNDA 0.341479f
C2546 VDDA.t31 GNDA 0.527449f
C2547 VDDA.t124 GNDA 0.29198f
C2548 VDDA.t173 GNDA 0.29198f
C2549 VDDA.t159 GNDA 0.29198f
C2550 VDDA.t425 GNDA 0.29198f
C2551 VDDA.t128 GNDA 0.218985f
C2552 VDDA.n354 GNDA 0.07758f
C2553 VDDA.n355 GNDA 0.099438f
C2554 VDDA.n356 GNDA 0.099438f
C2555 VDDA.t49 GNDA 0.527449f
C2556 VDDA.t126 GNDA 0.29198f
C2557 VDDA.t122 GNDA 0.29198f
C2558 VDDA.t284 GNDA 0.29198f
C2559 VDDA.t136 GNDA 0.29198f
C2560 VDDA.t157 GNDA 0.218985f
C2561 VDDA.n357 GNDA 0.14599f
C2562 VDDA.n358 GNDA 0.09879f
C2563 VDDA.n359 GNDA 0.067039f
C2564 VDDA.n360 GNDA 0.05185f
C2565 VDDA.t30 GNDA 0.046386f
C2566 VDDA.n361 GNDA 0.08875f
C2567 VDDA.n362 GNDA 0.123774f
C2568 VDDA.n363 GNDA 0.094779f
C2569 VDDA.n364 GNDA 0.053087f
C2570 VDDA.n365 GNDA 0.179525f
C2571 VDDA.n366 GNDA 0.061962f
C2572 VDDA.n367 GNDA 0.165419f
C2573 VDDA.t11 GNDA 0.012052f
C2574 VDDA.n368 GNDA 0.025644f
C2575 VDDA.t114 GNDA 0.012052f
C2576 VDDA.n369 GNDA 0.025644f
C2577 VDDA.n370 GNDA 0.037234f
C2578 VDDA.n371 GNDA 0.062583f
C2579 VDDA.n372 GNDA 0.166785f
C2580 VDDA.t41 GNDA 0.012052f
C2581 VDDA.n373 GNDA 0.025644f
C2582 VDDA.t29 GNDA 0.012052f
C2583 VDDA.n374 GNDA 0.025644f
C2584 VDDA.n375 GNDA 0.034699f
C2585 VDDA.n376 GNDA 0.043072f
C2586 VDDA.n377 GNDA 0.166785f
C2587 VDDA.t28 GNDA 0.16225f
C2588 VDDA.t216 GNDA 0.100258f
C2589 VDDA.t373 GNDA 0.100258f
C2590 VDDA.t371 GNDA 0.100258f
C2591 VDDA.t259 GNDA 0.100258f
C2592 VDDA.t228 GNDA 0.075194f
C2593 VDDA.t40 GNDA 0.16225f
C2594 VDDA.t340 GNDA 0.100258f
C2595 VDDA.t189 GNDA 0.100258f
C2596 VDDA.t155 GNDA 0.100258f
C2597 VDDA.t2 GNDA 0.100258f
C2598 VDDA.t305 GNDA 0.075194f
C2599 VDDA.n378 GNDA 0.063203f
C2600 VDDA.n379 GNDA 0.050129f
C2601 VDDA.n380 GNDA 0.063203f
C2602 VDDA.n381 GNDA 0.042214f
C2603 VDDA.n382 GNDA 0.034155f
C2604 VDDA.n383 GNDA 0.079415f
C2605 VDDA.n384 GNDA 0.079415f
C2606 VDDA.n385 GNDA 0.165419f
C2607 VDDA.t113 GNDA 0.158978f
C2608 VDDA.t227 GNDA 0.098499f
C2609 VDDA.t433 GNDA 0.098499f
C2610 VDDA.t436 GNDA 0.098499f
C2611 VDDA.t229 GNDA 0.098499f
C2612 VDDA.t215 GNDA 0.073874f
C2613 VDDA.t10 GNDA 0.158978f
C2614 VDDA.t337 GNDA 0.098499f
C2615 VDDA.t258 GNDA 0.098499f
C2616 VDDA.t190 GNDA 0.098499f
C2617 VDDA.t372 GNDA 0.098499f
C2618 VDDA.t186 GNDA 0.073874f
C2619 VDDA.n386 GNDA 0.063203f
C2620 VDDA.n387 GNDA 0.04925f
C2621 VDDA.n388 GNDA 0.063203f
C2622 VDDA.n389 GNDA 0.042013f
C2623 VDDA.n390 GNDA 0.034155f
C2624 VDDA.n391 GNDA 0.066121f
C2625 VDDA.n392 GNDA 0.088448f
C2626 VDDA.n394 GNDA 0.048973f
C2627 VDDA.n395 GNDA 0.077392f
C2628 VDDA.n396 GNDA 0.098194f
C2629 VDDA.n397 GNDA 0.098194f
C2630 VDDA.n398 GNDA 0.098194f
C2631 VDDA.n400 GNDA 0.048973f
C2632 VDDA.n402 GNDA 0.048973f
C2633 VDDA.n404 GNDA 0.048973f
C2634 VDDA.n406 GNDA 0.048973f
C2635 VDDA.n408 GNDA 0.048973f
C2636 VDDA.n410 GNDA 0.048973f
C2637 VDDA.n412 GNDA 0.048973f
C2638 VDDA.n414 GNDA 0.048973f
C2639 VDDA.n416 GNDA 0.08014f
C2640 VDDA.t93 GNDA 0.011653f
C2641 VDDA.n417 GNDA 0.017303f
C2642 VDDA.n418 GNDA 0.015309f
C2643 VDDA.n419 GNDA 0.052288f
C2644 VDDA.n420 GNDA 0.060755f
C2645 VDDA.n421 GNDA 0.200785f
C2646 VDDA.t92 GNDA 0.158978f
C2647 VDDA.t219 GNDA 0.098499f
C2648 VDDA.t351 GNDA 0.098499f
C2649 VDDA.t191 GNDA 0.098499f
C2650 VDDA.t357 GNDA 0.098499f
C2651 VDDA.t264 GNDA 0.098499f
C2652 VDDA.t347 GNDA 0.098499f
C2653 VDDA.t166 GNDA 0.098499f
C2654 VDDA.t363 GNDA 0.098499f
C2655 VDDA.t276 GNDA 0.098499f
C2656 VDDA.t217 GNDA 0.073874f
C2657 VDDA.n422 GNDA 0.04925f
C2658 VDDA.t355 GNDA 0.073874f
C2659 VDDA.t365 GNDA 0.098499f
C2660 VDDA.t359 GNDA 0.098499f
C2661 VDDA.t262 GNDA 0.098499f
C2662 VDDA.t353 GNDA 0.098499f
C2663 VDDA.t164 GNDA 0.098499f
C2664 VDDA.t349 GNDA 0.098499f
C2665 VDDA.t318 GNDA 0.098499f
C2666 VDDA.t193 GNDA 0.098499f
C2667 VDDA.t361 GNDA 0.098499f
C2668 VDDA.t89 GNDA 0.158978f
C2669 VDDA.n423 GNDA 0.200785f
C2670 VDDA.n424 GNDA 0.060755f
C2671 VDDA.n425 GNDA 0.052288f
C2672 VDDA.n426 GNDA 0.015309f
C2673 VDDA.t90 GNDA 0.011653f
C2674 VDDA.n427 GNDA 0.016881f
C2675 VDDA.n428 GNDA 0.083978f
C2676 VDDA.n429 GNDA 0.078091f
C2677 VDDA.n431 GNDA 0.062411f
C2678 VDDA.n432 GNDA 0.011513f
C2679 VDDA.n433 GNDA 0.034008f
C2680 VDDA.n434 GNDA 0.034008f
C2681 VDDA.n435 GNDA 0.034676f
C2682 VDDA.n436 GNDA 0.087131f
C2683 VDDA.n437 GNDA 0.011513f
C2684 VDDA.n438 GNDA 0.051139f
C2685 VDDA.n439 GNDA 0.051139f
C2686 VDDA.n440 GNDA 0.051138f
C2687 VDDA.t332 GNDA 0.020467f
C2688 VDDA.n441 GNDA 0.071025f
C2689 VDDA.t8 GNDA 0.093488f
C2690 VDDA.n442 GNDA 0.046359f
C2691 VDDA.n443 GNDA 0.044505f
C2692 VDDA.t6 GNDA 0.035523f
C2693 VDDA.n444 GNDA 0.037609f
C2694 VDDA.n445 GNDA 0.028151f
C2695 VDDA.n446 GNDA 0.043741f
C2696 VDDA.n447 GNDA 0.286765f
C2697 VDDA.t7 GNDA 0.272593f
C2698 VDDA.n448 GNDA 0.088745f
C2699 VDDA.n449 GNDA 0.022186f
C2700 VDDA.t331 GNDA 0.124243f
C2701 VDDA.t22 GNDA 0.294779f
C2702 VDDA.n450 GNDA 0.289735f
C2703 VDDA.n451 GNDA 0.045389f
C2704 VDDA.n452 GNDA 0.029106f
C2705 VDDA.t21 GNDA 0.036161f
C2706 VDDA.n453 GNDA 0.037609f
C2707 VDDA.t23 GNDA 0.073021f
C2708 VDDA.n454 GNDA 0.050113f
C2709 VDDA.n455 GNDA 0.099727f
C2710 VDDA.n456 GNDA 0.066341f
C2711 VDDA.t38 GNDA 0.01495f
C2712 VDDA.n457 GNDA 0.016242f
C2713 VDDA.t36 GNDA 0.012542f
C2714 VDDA.n458 GNDA 0.01588f
C2715 VDDA.n459 GNDA 0.020446f
C2716 VDDA.n460 GNDA 0.028693f
C2717 VDDA.n461 GNDA 0.153047f
C2718 VDDA.t37 GNDA 0.169511f
C2719 VDDA.t329 GNDA 0.115129f
C2720 VDDA.t70 GNDA 0.169511f
C2721 VDDA.n462 GNDA 0.153047f
C2722 VDDA.n463 GNDA 0.028693f
C2723 VDDA.n464 GNDA 0.020446f
C2724 VDDA.t69 GNDA 0.012542f
C2725 VDDA.n465 GNDA 0.01588f
C2726 VDDA.t72 GNDA 0.01495f
C2727 VDDA.n466 GNDA 0.018131f
C2728 VDDA.n467 GNDA 0.06222f
C2729 VDDA.n468 GNDA 0.182726f
C2730 VDDA.n469 GNDA 1.6515f
C2731 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039179f
C2732 bgr_0.PFET_GATE_10uA.t29 GNDA 0.057916f
C2733 bgr_0.PFET_GATE_10uA.n0 GNDA 0.063817f
C2734 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039179f
C2735 bgr_0.PFET_GATE_10uA.t21 GNDA 0.057916f
C2736 bgr_0.PFET_GATE_10uA.n1 GNDA 0.063817f
C2737 bgr_0.PFET_GATE_10uA.n2 GNDA 0.076791f
C2738 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039179f
C2739 bgr_0.PFET_GATE_10uA.t16 GNDA 0.057916f
C2740 bgr_0.PFET_GATE_10uA.n3 GNDA 0.063817f
C2741 bgr_0.PFET_GATE_10uA.t17 GNDA 0.039179f
C2742 bgr_0.PFET_GATE_10uA.t23 GNDA 0.057916f
C2743 bgr_0.PFET_GATE_10uA.n4 GNDA 0.063817f
C2744 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064022f
C2745 bgr_0.PFET_GATE_10uA.t0 GNDA 0.781422f
C2746 bgr_0.PFET_GATE_10uA.t1 GNDA 0.586977f
C2747 bgr_0.PFET_GATE_10uA.t2 GNDA 0.040183f
C2748 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040183f
C2749 bgr_0.PFET_GATE_10uA.n6 GNDA 0.102705f
C2750 bgr_0.PFET_GATE_10uA.t3 GNDA 0.040183f
C2751 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040183f
C2752 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100051f
C2753 bgr_0.PFET_GATE_10uA.n8 GNDA 0.978629f
C2754 bgr_0.PFET_GATE_10uA.t4 GNDA 0.040183f
C2755 bgr_0.PFET_GATE_10uA.t8 GNDA 0.040183f
C2756 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100051f
C2757 bgr_0.PFET_GATE_10uA.n10 GNDA 0.554934f
C2758 bgr_0.PFET_GATE_10uA.n11 GNDA 1.13286f
C2759 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040183f
C2760 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040183f
C2761 bgr_0.PFET_GATE_10uA.n12 GNDA 0.096913f
C2762 bgr_0.PFET_GATE_10uA.n13 GNDA 0.356682f
C2763 bgr_0.PFET_GATE_10uA.n14 GNDA 3.84996f
C2764 bgr_0.PFET_GATE_10uA.t11 GNDA 0.045299f
C2765 bgr_0.PFET_GATE_10uA.t20 GNDA 0.045299f
C2766 bgr_0.PFET_GATE_10uA.n15 GNDA 0.137138f
C2767 bgr_0.PFET_GATE_10uA.n16 GNDA 1.78858f
C2768 bgr_0.PFET_GATE_10uA.n17 GNDA 1.41725f
C2769 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039179f
C2770 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039179f
C2771 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039179f
C2772 bgr_0.PFET_GATE_10uA.t15 GNDA 0.039179f
C2773 bgr_0.PFET_GATE_10uA.t25 GNDA 0.039179f
C2774 bgr_0.PFET_GATE_10uA.t27 GNDA 0.057916f
C2775 bgr_0.PFET_GATE_10uA.n18 GNDA 0.071675f
C2776 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051234f
C2777 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051234f
C2778 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051234f
C2779 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043376f
C2780 bgr_0.PFET_GATE_10uA.t13 GNDA 0.039179f
C2781 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039179f
C2782 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039179f
C2783 bgr_0.PFET_GATE_10uA.t24 GNDA 0.057916f
C2784 bgr_0.PFET_GATE_10uA.n23 GNDA 0.071675f
C2785 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051234f
C2786 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043376f
C2787 bgr_0.PFET_GATE_10uA.n26 GNDA 0.05954f
C2788 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.344645f
C2789 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.167175f
C2790 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198327f
C2791 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.344645f
C2792 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.167175f
C2793 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216884f
C2794 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.344645f
C2795 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.167175f
C2796 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216884f
C2797 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.344645f
C2798 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.167175f
C2799 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216884f
C2800 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C2801 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.345795f
C2802 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.364353f
C2803 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.364353f
C2804 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.364353f
C2805 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185733f
C2806 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216884f
C2807 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C2808 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.345795f
C2809 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.364353f
C2810 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.364353f
C2811 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.364353f
C2812 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.185733f
C2813 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216884f
C2814 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345795f
C2815 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.347048f
C2816 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345795f
C2817 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.348506f
C2818 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.37905f
C2819 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.345795f
C2820 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.347048f
C2821 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.345795f
C2822 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.347048f
C2823 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.345795f
C2824 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.347048f
C2825 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.345795f
C2826 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.347048f
C2827 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345795f
C2828 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.347048f
C2829 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.345795f
C2830 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.347048f
C2831 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.345795f
C2832 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.347048f
C2833 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.345795f
C2834 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.347048f
C2835 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345795f
C2836 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.347048f
C2837 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345795f
C2838 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.347048f
C2839 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345795f
C2840 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.347048f
C2841 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.345795f
C2842 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.347048f
C2843 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345795f
C2844 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.347048f
C2845 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345795f
C2846 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.347048f
C2847 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345795f
C2848 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.347048f
C2849 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.345795f
C2850 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.347048f
C2851 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345795f
C2852 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.347048f
C2853 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345795f
C2854 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.347048f
C2855 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.345795f
C2856 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.347048f
C2857 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.345795f
C2858 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.347048f
C2859 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345795f
C2860 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.347048f
C2861 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.345795f
C2862 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.347048f
C2863 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345795f
C2864 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.347048f
C2865 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.345795f
C2866 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.347048f
C2867 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.345795f
C2868 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.347048f
C2869 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.345795f
C2870 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.347048f
C2871 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.345795f
C2872 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.347048f
C2873 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345795f
C2874 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.347048f
C2875 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.345795f
C2876 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.362749f
C2877 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.345795f
C2878 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.185733f
C2879 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.198781f
C2880 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345795f
C2881 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185733f
C2882 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197177f
C2883 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345795f
C2884 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.185733f
C2885 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197177f
C2886 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.345795f
C2887 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.185733f
C2888 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.197177f
C2889 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.345795f
C2890 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185733f
C2891 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.197177f
C2892 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345795f
C2893 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.185733f
C2894 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.197177f
C2895 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345795f
C2896 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.185733f
C2897 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.197177f
C2898 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.345795f
C2899 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.185733f
C2900 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.197177f
C2901 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345795f
C2902 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185733f
C2903 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.197177f
C2904 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345795f
C2905 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.347048f
C2906 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.345795f
C2907 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.347048f
C2908 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.167175f
C2909 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.215631f
C2910 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.184584f
C2911 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.234189f
C2912 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.184584f
C2913 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251494f
C2914 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.184584f
C2915 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251494f
C2916 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.184584f
C2917 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251494f
C2918 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.184584f
C2919 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251494f
C2920 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.184584f
C2921 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251494f
C2922 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.184584f
C2923 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251494f
C2924 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.184584f
C2925 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251494f
C2926 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.184584f
C2927 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251494f
C2928 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.184584f
C2929 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.251494f
C2930 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.184584f
C2931 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.251494f
C2932 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.184584f
C2933 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.251494f
C2934 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.184584f
C2935 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.251494f
C2936 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.184584f
C2937 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.251494f
C2938 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.184584f
C2939 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.251494f
C2940 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.184584f
C2941 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.234189f
C2942 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.344645f
C2943 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.167175f
C2944 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216884f
C2945 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C2946 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.167175f
C2947 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216884f
C2948 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C2949 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.345795f
C2950 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.364353f
C2951 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.364353f
C2952 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.364353f
C2953 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185733f
C2954 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216884f
C2955 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.344645f
C2956 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216884f
C2957 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185733f
C2958 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.364353f
C2959 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.364353f
C2960 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.364353f
C2961 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.337351f
C2962 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.298183f
C2963 two_stage_opamp_dummy_magic_0.VOUT-.t11 GNDA 0.051003f
C2964 two_stage_opamp_dummy_magic_0.VOUT-.t9 GNDA 0.051003f
C2965 two_stage_opamp_dummy_magic_0.VOUT-.n0 GNDA 0.235943f
C2966 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA 0.051003f
C2967 two_stage_opamp_dummy_magic_0.VOUT-.t8 GNDA 0.051003f
C2968 two_stage_opamp_dummy_magic_0.VOUT-.n1 GNDA 0.235153f
C2969 two_stage_opamp_dummy_magic_0.VOUT-.n2 GNDA 0.145313f
C2970 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA 0.051003f
C2971 two_stage_opamp_dummy_magic_0.VOUT-.t10 GNDA 0.051003f
C2972 two_stage_opamp_dummy_magic_0.VOUT-.n3 GNDA 0.235153f
C2973 two_stage_opamp_dummy_magic_0.VOUT-.n4 GNDA 0.089445f
C2974 two_stage_opamp_dummy_magic_0.VOUT-.t14 GNDA 0.043717f
C2975 two_stage_opamp_dummy_magic_0.VOUT-.t1 GNDA 0.043717f
C2976 two_stage_opamp_dummy_magic_0.VOUT-.n5 GNDA 0.175711f
C2977 two_stage_opamp_dummy_magic_0.VOUT-.t2 GNDA 0.043717f
C2978 two_stage_opamp_dummy_magic_0.VOUT-.t15 GNDA 0.043717f
C2979 two_stage_opamp_dummy_magic_0.VOUT-.n6 GNDA 0.17571f
C2980 two_stage_opamp_dummy_magic_0.VOUT-.t13 GNDA 0.043717f
C2981 two_stage_opamp_dummy_magic_0.VOUT-.t0 GNDA 0.043717f
C2982 two_stage_opamp_dummy_magic_0.VOUT-.n7 GNDA 0.175387f
C2983 two_stage_opamp_dummy_magic_0.VOUT-.n8 GNDA 0.172777f
C2984 two_stage_opamp_dummy_magic_0.VOUT-.t5 GNDA 0.043717f
C2985 two_stage_opamp_dummy_magic_0.VOUT-.t4 GNDA 0.043717f
C2986 two_stage_opamp_dummy_magic_0.VOUT-.n9 GNDA 0.175387f
C2987 two_stage_opamp_dummy_magic_0.VOUT-.n10 GNDA 0.0891f
C2988 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA 0.043717f
C2989 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA 0.043717f
C2990 two_stage_opamp_dummy_magic_0.VOUT-.n11 GNDA 0.175387f
C2991 two_stage_opamp_dummy_magic_0.VOUT-.n12 GNDA 0.0891f
C2992 two_stage_opamp_dummy_magic_0.VOUT-.n13 GNDA 0.105535f
C2993 two_stage_opamp_dummy_magic_0.VOUT-.t7 GNDA 0.043717f
C2994 two_stage_opamp_dummy_magic_0.VOUT-.t6 GNDA 0.043717f
C2995 two_stage_opamp_dummy_magic_0.VOUT-.n14 GNDA 0.17324f
C2996 two_stage_opamp_dummy_magic_0.VOUT-.n15 GNDA 0.211953f
C2997 two_stage_opamp_dummy_magic_0.VOUT-.t100 GNDA 0.291446f
C2998 two_stage_opamp_dummy_magic_0.VOUT-.t107 GNDA 0.29641f
C2999 two_stage_opamp_dummy_magic_0.VOUT-.t149 GNDA 0.291446f
C3000 two_stage_opamp_dummy_magic_0.VOUT-.n16 GNDA 0.195405f
C3001 two_stage_opamp_dummy_magic_0.VOUT-.n17 GNDA 0.127508f
C3002 two_stage_opamp_dummy_magic_0.VOUT-.t47 GNDA 0.295788f
C3003 two_stage_opamp_dummy_magic_0.VOUT-.t91 GNDA 0.295788f
C3004 two_stage_opamp_dummy_magic_0.VOUT-.t41 GNDA 0.295788f
C3005 two_stage_opamp_dummy_magic_0.VOUT-.t130 GNDA 0.295788f
C3006 two_stage_opamp_dummy_magic_0.VOUT-.t82 GNDA 0.295788f
C3007 two_stage_opamp_dummy_magic_0.VOUT-.t124 GNDA 0.295788f
C3008 two_stage_opamp_dummy_magic_0.VOUT-.t72 GNDA 0.295788f
C3009 two_stage_opamp_dummy_magic_0.VOUT-.t23 GNDA 0.295788f
C3010 two_stage_opamp_dummy_magic_0.VOUT-.t62 GNDA 0.295788f
C3011 two_stage_opamp_dummy_magic_0.VOUT-.t150 GNDA 0.295788f
C3012 two_stage_opamp_dummy_magic_0.VOUT-.t86 GNDA 0.291446f
C3013 two_stage_opamp_dummy_magic_0.VOUT-.n18 GNDA 0.196026f
C3014 two_stage_opamp_dummy_magic_0.VOUT-.t50 GNDA 0.291446f
C3015 two_stage_opamp_dummy_magic_0.VOUT-.n19 GNDA 0.250673f
C3016 two_stage_opamp_dummy_magic_0.VOUT-.t137 GNDA 0.291446f
C3017 two_stage_opamp_dummy_magic_0.VOUT-.n20 GNDA 0.250673f
C3018 two_stage_opamp_dummy_magic_0.VOUT-.t105 GNDA 0.291446f
C3019 two_stage_opamp_dummy_magic_0.VOUT-.n21 GNDA 0.250673f
C3020 two_stage_opamp_dummy_magic_0.VOUT-.t73 GNDA 0.291446f
C3021 two_stage_opamp_dummy_magic_0.VOUT-.n22 GNDA 0.250673f
C3022 two_stage_opamp_dummy_magic_0.VOUT-.t25 GNDA 0.291446f
C3023 two_stage_opamp_dummy_magic_0.VOUT-.n23 GNDA 0.250673f
C3024 two_stage_opamp_dummy_magic_0.VOUT-.t127 GNDA 0.291446f
C3025 two_stage_opamp_dummy_magic_0.VOUT-.n24 GNDA 0.250673f
C3026 two_stage_opamp_dummy_magic_0.VOUT-.t88 GNDA 0.291446f
C3027 two_stage_opamp_dummy_magic_0.VOUT-.n25 GNDA 0.250673f
C3028 two_stage_opamp_dummy_magic_0.VOUT-.t53 GNDA 0.291446f
C3029 two_stage_opamp_dummy_magic_0.VOUT-.n26 GNDA 0.250673f
C3030 two_stage_opamp_dummy_magic_0.VOUT-.t140 GNDA 0.291446f
C3031 two_stage_opamp_dummy_magic_0.VOUT-.n27 GNDA 0.250673f
C3032 two_stage_opamp_dummy_magic_0.VOUT-.t109 GNDA 0.291446f
C3033 two_stage_opamp_dummy_magic_0.VOUT-.t28 GNDA 0.29641f
C3034 two_stage_opamp_dummy_magic_0.VOUT-.t78 GNDA 0.291446f
C3035 two_stage_opamp_dummy_magic_0.VOUT-.n28 GNDA 0.195405f
C3036 two_stage_opamp_dummy_magic_0.VOUT-.n29 GNDA 0.2368f
C3037 two_stage_opamp_dummy_magic_0.VOUT-.t24 GNDA 0.29641f
C3038 two_stage_opamp_dummy_magic_0.VOUT-.t112 GNDA 0.291446f
C3039 two_stage_opamp_dummy_magic_0.VOUT-.n30 GNDA 0.195405f
C3040 two_stage_opamp_dummy_magic_0.VOUT-.t77 GNDA 0.291446f
C3041 two_stage_opamp_dummy_magic_0.VOUT-.t129 GNDA 0.29641f
C3042 two_stage_opamp_dummy_magic_0.VOUT-.t37 GNDA 0.291446f
C3043 two_stage_opamp_dummy_magic_0.VOUT-.n31 GNDA 0.195405f
C3044 two_stage_opamp_dummy_magic_0.VOUT-.n32 GNDA 0.2368f
C3045 two_stage_opamp_dummy_magic_0.VOUT-.t59 GNDA 0.29641f
C3046 two_stage_opamp_dummy_magic_0.VOUT-.t147 GNDA 0.291446f
C3047 two_stage_opamp_dummy_magic_0.VOUT-.n33 GNDA 0.195405f
C3048 two_stage_opamp_dummy_magic_0.VOUT-.t116 GNDA 0.291446f
C3049 two_stage_opamp_dummy_magic_0.VOUT-.t32 GNDA 0.29641f
C3050 two_stage_opamp_dummy_magic_0.VOUT-.t81 GNDA 0.291446f
C3051 two_stage_opamp_dummy_magic_0.VOUT-.n34 GNDA 0.195405f
C3052 two_stage_opamp_dummy_magic_0.VOUT-.n35 GNDA 0.2368f
C3053 two_stage_opamp_dummy_magic_0.VOUT-.t99 GNDA 0.29641f
C3054 two_stage_opamp_dummy_magic_0.VOUT-.t46 GNDA 0.291446f
C3055 two_stage_opamp_dummy_magic_0.VOUT-.n36 GNDA 0.195405f
C3056 two_stage_opamp_dummy_magic_0.VOUT-.t153 GNDA 0.291446f
C3057 two_stage_opamp_dummy_magic_0.VOUT-.t69 GNDA 0.29641f
C3058 two_stage_opamp_dummy_magic_0.VOUT-.t122 GNDA 0.291446f
C3059 two_stage_opamp_dummy_magic_0.VOUT-.n37 GNDA 0.195405f
C3060 two_stage_opamp_dummy_magic_0.VOUT-.n38 GNDA 0.2368f
C3061 two_stage_opamp_dummy_magic_0.VOUT-.t67 GNDA 0.29641f
C3062 two_stage_opamp_dummy_magic_0.VOUT-.t154 GNDA 0.291446f
C3063 two_stage_opamp_dummy_magic_0.VOUT-.n39 GNDA 0.195405f
C3064 two_stage_opamp_dummy_magic_0.VOUT-.t123 GNDA 0.291446f
C3065 two_stage_opamp_dummy_magic_0.VOUT-.t35 GNDA 0.29641f
C3066 two_stage_opamp_dummy_magic_0.VOUT-.t84 GNDA 0.291446f
C3067 two_stage_opamp_dummy_magic_0.VOUT-.n40 GNDA 0.195405f
C3068 two_stage_opamp_dummy_magic_0.VOUT-.n41 GNDA 0.2368f
C3069 two_stage_opamp_dummy_magic_0.VOUT-.t104 GNDA 0.29641f
C3070 two_stage_opamp_dummy_magic_0.VOUT-.t52 GNDA 0.291446f
C3071 two_stage_opamp_dummy_magic_0.VOUT-.n42 GNDA 0.195405f
C3072 two_stage_opamp_dummy_magic_0.VOUT-.t22 GNDA 0.291446f
C3073 two_stage_opamp_dummy_magic_0.VOUT-.t76 GNDA 0.29641f
C3074 two_stage_opamp_dummy_magic_0.VOUT-.t126 GNDA 0.291446f
C3075 two_stage_opamp_dummy_magic_0.VOUT-.n43 GNDA 0.195405f
C3076 two_stage_opamp_dummy_magic_0.VOUT-.n44 GNDA 0.2368f
C3077 two_stage_opamp_dummy_magic_0.VOUT-.t95 GNDA 0.291446f
C3078 two_stage_opamp_dummy_magic_0.VOUT-.t83 GNDA 0.29641f
C3079 two_stage_opamp_dummy_magic_0.VOUT-.t56 GNDA 0.291446f
C3080 two_stage_opamp_dummy_magic_0.VOUT-.n45 GNDA 0.195405f
C3081 two_stage_opamp_dummy_magic_0.VOUT-.n46 GNDA 0.127508f
C3082 two_stage_opamp_dummy_magic_0.VOUT-.t132 GNDA 0.295788f
C3083 two_stage_opamp_dummy_magic_0.VOUT-.t114 GNDA 0.295788f
C3084 two_stage_opamp_dummy_magic_0.VOUT-.t90 GNDA 0.29641f
C3085 two_stage_opamp_dummy_magic_0.VOUT-.t131 GNDA 0.291446f
C3086 two_stage_opamp_dummy_magic_0.VOUT-.n47 GNDA 0.195405f
C3087 two_stage_opamp_dummy_magic_0.VOUT-.t103 GNDA 0.291446f
C3088 two_stage_opamp_dummy_magic_0.VOUT-.n48 GNDA 0.127508f
C3089 two_stage_opamp_dummy_magic_0.VOUT-.t71 GNDA 0.291446f
C3090 two_stage_opamp_dummy_magic_0.VOUT-.n49 GNDA 0.122954f
C3091 two_stage_opamp_dummy_magic_0.VOUT-.t146 GNDA 0.295788f
C3092 two_stage_opamp_dummy_magic_0.VOUT-.t128 GNDA 0.29641f
C3093 two_stage_opamp_dummy_magic_0.VOUT-.t31 GNDA 0.291446f
C3094 two_stage_opamp_dummy_magic_0.VOUT-.n50 GNDA 0.195405f
C3095 two_stage_opamp_dummy_magic_0.VOUT-.t138 GNDA 0.291446f
C3096 two_stage_opamp_dummy_magic_0.VOUT-.n51 GNDA 0.127508f
C3097 two_stage_opamp_dummy_magic_0.VOUT-.t106 GNDA 0.291446f
C3098 two_stage_opamp_dummy_magic_0.VOUT-.n52 GNDA 0.122954f
C3099 two_stage_opamp_dummy_magic_0.VOUT-.t45 GNDA 0.295788f
C3100 two_stage_opamp_dummy_magic_0.VOUT-.t26 GNDA 0.29641f
C3101 two_stage_opamp_dummy_magic_0.VOUT-.t60 GNDA 0.291446f
C3102 two_stage_opamp_dummy_magic_0.VOUT-.n53 GNDA 0.195405f
C3103 two_stage_opamp_dummy_magic_0.VOUT-.t40 GNDA 0.291446f
C3104 two_stage_opamp_dummy_magic_0.VOUT-.n54 GNDA 0.127508f
C3105 two_stage_opamp_dummy_magic_0.VOUT-.t143 GNDA 0.291446f
C3106 two_stage_opamp_dummy_magic_0.VOUT-.n55 GNDA 0.122954f
C3107 two_stage_opamp_dummy_magic_0.VOUT-.t85 GNDA 0.295788f
C3108 two_stage_opamp_dummy_magic_0.VOUT-.t74 GNDA 0.29641f
C3109 two_stage_opamp_dummy_magic_0.VOUT-.t113 GNDA 0.291446f
C3110 two_stage_opamp_dummy_magic_0.VOUT-.n56 GNDA 0.195405f
C3111 two_stage_opamp_dummy_magic_0.VOUT-.t21 GNDA 0.291446f
C3112 two_stage_opamp_dummy_magic_0.VOUT-.n57 GNDA 0.127508f
C3113 two_stage_opamp_dummy_magic_0.VOUT-.t125 GNDA 0.291446f
C3114 two_stage_opamp_dummy_magic_0.VOUT-.n58 GNDA 0.122954f
C3115 two_stage_opamp_dummy_magic_0.VOUT-.t63 GNDA 0.295788f
C3116 two_stage_opamp_dummy_magic_0.VOUT-.t101 GNDA 0.295788f
C3117 two_stage_opamp_dummy_magic_0.VOUT-.t134 GNDA 0.295788f
C3118 two_stage_opamp_dummy_magic_0.VOUT-.t119 GNDA 0.295788f
C3119 two_stage_opamp_dummy_magic_0.VOUT-.t155 GNDA 0.295788f
C3120 two_stage_opamp_dummy_magic_0.VOUT-.t118 GNDA 0.291446f
C3121 two_stage_opamp_dummy_magic_0.VOUT-.n59 GNDA 0.196026f
C3122 two_stage_opamp_dummy_magic_0.VOUT-.t80 GNDA 0.291446f
C3123 two_stage_opamp_dummy_magic_0.VOUT-.n60 GNDA 0.250673f
C3124 two_stage_opamp_dummy_magic_0.VOUT-.t96 GNDA 0.291446f
C3125 two_stage_opamp_dummy_magic_0.VOUT-.n61 GNDA 0.250673f
C3126 two_stage_opamp_dummy_magic_0.VOUT-.t61 GNDA 0.291446f
C3127 two_stage_opamp_dummy_magic_0.VOUT-.n62 GNDA 0.250673f
C3128 two_stage_opamp_dummy_magic_0.VOUT-.t27 GNDA 0.291446f
C3129 two_stage_opamp_dummy_magic_0.VOUT-.n63 GNDA 0.309872f
C3130 two_stage_opamp_dummy_magic_0.VOUT-.t44 GNDA 0.291446f
C3131 two_stage_opamp_dummy_magic_0.VOUT-.n64 GNDA 0.309872f
C3132 two_stage_opamp_dummy_magic_0.VOUT-.t144 GNDA 0.291446f
C3133 two_stage_opamp_dummy_magic_0.VOUT-.n65 GNDA 0.309872f
C3134 two_stage_opamp_dummy_magic_0.VOUT-.t111 GNDA 0.291446f
C3135 two_stage_opamp_dummy_magic_0.VOUT-.n66 GNDA 0.309872f
C3136 two_stage_opamp_dummy_magic_0.VOUT-.t75 GNDA 0.291446f
C3137 two_stage_opamp_dummy_magic_0.VOUT-.n67 GNDA 0.250673f
C3138 two_stage_opamp_dummy_magic_0.VOUT-.t92 GNDA 0.291446f
C3139 two_stage_opamp_dummy_magic_0.VOUT-.n68 GNDA 0.250673f
C3140 two_stage_opamp_dummy_magic_0.VOUT-.t55 GNDA 0.291446f
C3141 two_stage_opamp_dummy_magic_0.VOUT-.t39 GNDA 0.29641f
C3142 two_stage_opamp_dummy_magic_0.VOUT-.t19 GNDA 0.291446f
C3143 two_stage_opamp_dummy_magic_0.VOUT-.n69 GNDA 0.195405f
C3144 two_stage_opamp_dummy_magic_0.VOUT-.n70 GNDA 0.2368f
C3145 two_stage_opamp_dummy_magic_0.VOUT-.t34 GNDA 0.29641f
C3146 two_stage_opamp_dummy_magic_0.VOUT-.t51 GNDA 0.291446f
C3147 two_stage_opamp_dummy_magic_0.VOUT-.n71 GNDA 0.195405f
C3148 two_stage_opamp_dummy_magic_0.VOUT-.t156 GNDA 0.291446f
C3149 two_stage_opamp_dummy_magic_0.VOUT-.t136 GNDA 0.29641f
C3150 two_stage_opamp_dummy_magic_0.VOUT-.t120 GNDA 0.291446f
C3151 two_stage_opamp_dummy_magic_0.VOUT-.n72 GNDA 0.195405f
C3152 two_stage_opamp_dummy_magic_0.VOUT-.n73 GNDA 0.2368f
C3153 two_stage_opamp_dummy_magic_0.VOUT-.t68 GNDA 0.29641f
C3154 two_stage_opamp_dummy_magic_0.VOUT-.t87 GNDA 0.291446f
C3155 two_stage_opamp_dummy_magic_0.VOUT-.n74 GNDA 0.195405f
C3156 two_stage_opamp_dummy_magic_0.VOUT-.t49 GNDA 0.291446f
C3157 two_stage_opamp_dummy_magic_0.VOUT-.t36 GNDA 0.29641f
C3158 two_stage_opamp_dummy_magic_0.VOUT-.t151 GNDA 0.291446f
C3159 two_stage_opamp_dummy_magic_0.VOUT-.n75 GNDA 0.195405f
C3160 two_stage_opamp_dummy_magic_0.VOUT-.n76 GNDA 0.2368f
C3161 two_stage_opamp_dummy_magic_0.VOUT-.t94 GNDA 0.29641f
C3162 two_stage_opamp_dummy_magic_0.VOUT-.t42 GNDA 0.291446f
C3163 two_stage_opamp_dummy_magic_0.VOUT-.n77 GNDA 0.195405f
C3164 two_stage_opamp_dummy_magic_0.VOUT-.t145 GNDA 0.291446f
C3165 two_stage_opamp_dummy_magic_0.VOUT-.t64 GNDA 0.29641f
C3166 two_stage_opamp_dummy_magic_0.VOUT-.t117 GNDA 0.291446f
C3167 two_stage_opamp_dummy_magic_0.VOUT-.n78 GNDA 0.195405f
C3168 two_stage_opamp_dummy_magic_0.VOUT-.n79 GNDA 0.2368f
C3169 two_stage_opamp_dummy_magic_0.VOUT-.t54 GNDA 0.29641f
C3170 two_stage_opamp_dummy_magic_0.VOUT-.t141 GNDA 0.291446f
C3171 two_stage_opamp_dummy_magic_0.VOUT-.n80 GNDA 0.195405f
C3172 two_stage_opamp_dummy_magic_0.VOUT-.t110 GNDA 0.291446f
C3173 two_stage_opamp_dummy_magic_0.VOUT-.t29 GNDA 0.29641f
C3174 two_stage_opamp_dummy_magic_0.VOUT-.t79 GNDA 0.291446f
C3175 two_stage_opamp_dummy_magic_0.VOUT-.n81 GNDA 0.195405f
C3176 two_stage_opamp_dummy_magic_0.VOUT-.n82 GNDA 0.2368f
C3177 two_stage_opamp_dummy_magic_0.VOUT-.t89 GNDA 0.29641f
C3178 two_stage_opamp_dummy_magic_0.VOUT-.t38 GNDA 0.291446f
C3179 two_stage_opamp_dummy_magic_0.VOUT-.n83 GNDA 0.195405f
C3180 two_stage_opamp_dummy_magic_0.VOUT-.t139 GNDA 0.291446f
C3181 two_stage_opamp_dummy_magic_0.VOUT-.t57 GNDA 0.29641f
C3182 two_stage_opamp_dummy_magic_0.VOUT-.t108 GNDA 0.291446f
C3183 two_stage_opamp_dummy_magic_0.VOUT-.n84 GNDA 0.195405f
C3184 two_stage_opamp_dummy_magic_0.VOUT-.n85 GNDA 0.2368f
C3185 two_stage_opamp_dummy_magic_0.VOUT-.t48 GNDA 0.29641f
C3186 two_stage_opamp_dummy_magic_0.VOUT-.t135 GNDA 0.291446f
C3187 two_stage_opamp_dummy_magic_0.VOUT-.n86 GNDA 0.195405f
C3188 two_stage_opamp_dummy_magic_0.VOUT-.t102 GNDA 0.291446f
C3189 two_stage_opamp_dummy_magic_0.VOUT-.t20 GNDA 0.29641f
C3190 two_stage_opamp_dummy_magic_0.VOUT-.t70 GNDA 0.291446f
C3191 two_stage_opamp_dummy_magic_0.VOUT-.n87 GNDA 0.195405f
C3192 two_stage_opamp_dummy_magic_0.VOUT-.n88 GNDA 0.2368f
C3193 two_stage_opamp_dummy_magic_0.VOUT-.t148 GNDA 0.29641f
C3194 two_stage_opamp_dummy_magic_0.VOUT-.t98 GNDA 0.291446f
C3195 two_stage_opamp_dummy_magic_0.VOUT-.n89 GNDA 0.195405f
C3196 two_stage_opamp_dummy_magic_0.VOUT-.t66 GNDA 0.291446f
C3197 two_stage_opamp_dummy_magic_0.VOUT-.t121 GNDA 0.29641f
C3198 two_stage_opamp_dummy_magic_0.VOUT-.t33 GNDA 0.291446f
C3199 two_stage_opamp_dummy_magic_0.VOUT-.n90 GNDA 0.195405f
C3200 two_stage_opamp_dummy_magic_0.VOUT-.n91 GNDA 0.2368f
C3201 two_stage_opamp_dummy_magic_0.VOUT-.t43 GNDA 0.29641f
C3202 two_stage_opamp_dummy_magic_0.VOUT-.t133 GNDA 0.291446f
C3203 two_stage_opamp_dummy_magic_0.VOUT-.n92 GNDA 0.195405f
C3204 two_stage_opamp_dummy_magic_0.VOUT-.t97 GNDA 0.291446f
C3205 two_stage_opamp_dummy_magic_0.VOUT-.t152 GNDA 0.29641f
C3206 two_stage_opamp_dummy_magic_0.VOUT-.t65 GNDA 0.291446f
C3207 two_stage_opamp_dummy_magic_0.VOUT-.n93 GNDA 0.195405f
C3208 two_stage_opamp_dummy_magic_0.VOUT-.n94 GNDA 0.2368f
C3209 two_stage_opamp_dummy_magic_0.VOUT-.t115 GNDA 0.29641f
C3210 two_stage_opamp_dummy_magic_0.VOUT-.t30 GNDA 0.291446f
C3211 two_stage_opamp_dummy_magic_0.VOUT-.n95 GNDA 0.195405f
C3212 two_stage_opamp_dummy_magic_0.VOUT-.t58 GNDA 0.291446f
C3213 two_stage_opamp_dummy_magic_0.VOUT-.n96 GNDA 0.2368f
C3214 two_stage_opamp_dummy_magic_0.VOUT-.t93 GNDA 0.291446f
C3215 two_stage_opamp_dummy_magic_0.VOUT-.n97 GNDA 0.127508f
C3216 two_stage_opamp_dummy_magic_0.VOUT-.t142 GNDA 0.291446f
C3217 two_stage_opamp_dummy_magic_0.VOUT-.n98 GNDA 0.23878f
C3218 two_stage_opamp_dummy_magic_0.VOUT-.n99 GNDA 0.286094f
C3219 two_stage_opamp_dummy_magic_0.VOUT-.n100 GNDA 0.166472f
C3220 two_stage_opamp_dummy_magic_0.VOUT-.t16 GNDA 0.084326f
C3221 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C3222 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C3223 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C3224 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C3225 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C3226 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C3227 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C3228 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C3229 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C3230 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C3231 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C3232 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C3233 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C3234 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C3235 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C3236 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C3237 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C3238 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C3239 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C3240 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C3241 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.04969f
C3242 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.186051f
C3243 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C3244 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C3245 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.050131f
C3246 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C3247 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C3248 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C3249 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.186051f
C3250 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.027755f
C3251 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C3252 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C3253 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C3254 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C3255 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C3256 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C3257 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C3258 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C3259 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C3260 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C3261 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C3262 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C3263 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.02366f
C3264 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.023535f
C3265 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.159426f
C3266 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.023535f
C3267 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.172681f
C3268 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.120742f
C3269 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.018869f
C3270 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.018869f
C3271 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.055362f
C3272 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.018869f
C3273 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.018869f
C3274 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.055111f
C3275 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.190495f
C3276 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.018869f
C3277 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.018869f
C3278 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.055111f
C3279 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.098676f
C3280 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.018869f
C3281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.018869f
C3282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.055111f
C3283 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.098676f
C3284 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.018869f
C3285 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.018869f
C3286 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.055111f
C3287 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.142441f
C3288 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 0.684243f
C3289 bgr_0.V_CMFB_S3 GNDA 0.540781f
.ends

