* NGSPICE file created from vco2_2_flat.ext - technology: sky130A

.subckt vco2_2_flat
X0 a_82_186# a_38_n62# V_OSC VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X1 a_636_n552# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X2 a_1190_n552# V_OSC a_592_n62# GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X3 a_82_186# GNDA VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X4 GNDA V_CONT a_n746_764.t2 GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X5 VDDA.t14 a_n746_764.t0 a_n746_764.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X6 a_82_n552# a_38_n62# V_OSC GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X7 a_1190_n552# VDDA.t17 GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X8 a_1190_n552# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X9 a_636_186# a_592_n62# a_38_n62# VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X10 a_82_n552# VDDA.t18 GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X11 a_82_n552# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X12 a_636_186# a_n746_764.t3 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X13 a_636_n552# a_592_n62# a_38_n62# GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X14 a_82_186# a_n746_764.t4 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X15 a_1190_186# V_OSC a_592_n62# VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X16 a_1190_186# a_n746_764.t5 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X17 a_636_186# GNDA VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X18 a_1190_186# GNDA VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X19 a_636_n552# VDDA.t19 GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
R0 VDDA.n1 VDDA.t17 1007.38
R1 VDDA.n2 VDDA.t18 618.567
R2 VDDA.t9 VDDA.t13 488.219
R3 VDDA.t2 VDDA.t15 480.288
R4 VDDA.n3 VDDA.n2 357.406
R5 VDDA VDDA.t1 354.445
R6 VDDA VDDA.t5 354.418
R7 VDDA.n3 VDDA.t3 349.767
R8 VDDA.n0 VDDA.t4 341.048
R9 VDDA.n2 VDDA.n1 308.481
R10 VDDA.n3 VDDA.n0 185
R11 VDDA VDDA.t14 143.486
R12 VDDA VDDA.t10 143.486
R13 VDDA VDDA.t12 143.486
R14 VDDA VDDA.t16 143.486
R15 VDDA.n0 VDDA.t11 139.239
R16 VDDA.n1 VDDA.t19 117.287
R17 VDDA.t7 VDDA.t0 6.16933
R18 VDDA.t6 VDDA.t2 6.16933
R19 VDDA.t4 VDDA.t8 6.16933
R20 VDDA VDDA.n3 2.50857
R21 VDDA.t15 VDDA.t7 1.76302
R22 VDDA.t11 VDDA.t6 1.76302
R23 VDDA.t8 VDDA.t9 1.76302
R24 a_n746_764.t2 a_n746_764.n2 466.82
R25 a_n746_764.n2 a_n746_764.t0 225.869
R26 a_n746_764.n2 a_n746_764.t1 225.786
R27 a_n746_764.t0 a_n746_764.n1 188.501
R28 a_n746_764.n0 a_n746_764.t5 188.501
R29 a_n746_764.n1 a_n746_764.n0 107.442
R30 a_n746_764.n1 a_n746_764.t4 81.0592
R31 a_n746_764.n0 a_n746_764.t3 81.0592
C0 a_1190_n552# V_OSC 0.302653f
C1 V_OSC a_592_n62# 0.077754f
C2 a_636_n552# a_636_186# 0.003006f
C3 a_1190_186# VDDA 0.529355f
C4 a_38_n62# VDDA 0.393692f
C5 VDDA a_636_186# 0.729489f
C6 V_CONT a_82_186# 0.002777f
C7 V_CONT a_82_n552# 0.041598f
C8 a_82_186# a_592_n62# 9.21e-20
C9 V_CONT a_636_n552# 0.041369f
C10 a_82_n552# a_592_n62# 6.76e-20
C11 a_636_n552# a_1190_n552# 0.005181f
C12 a_636_n552# a_592_n62# 0.040416f
C13 V_OSC a_82_186# 0.046372f
C14 a_82_n552# V_OSC 0.02745f
C15 a_1190_186# a_636_186# 0.006705f
C16 V_CONT VDDA 0.063762f
C17 a_636_n552# V_OSC 4.78e-19
C18 a_38_n62# a_636_186# 0.046372f
C19 VDDA a_1190_n552# 0.017309f
C20 VDDA a_592_n62# 0.251636f
C21 VDDA V_OSC 0.26411f
C22 a_82_n552# a_82_186# 0.001731f
C23 a_38_n62# V_CONT 0.002755f
C24 a_1190_186# a_592_n62# 0.046372f
C25 a_38_n62# a_592_n62# 0.073513f
C26 a_636_n552# a_82_n552# 0.007761f
C27 V_CONT a_636_186# 0.002777f
C28 a_1190_186# V_OSC 0.05908f
C29 a_38_n62# V_OSC 0.055458f
C30 VDDA a_82_186# 0.761173f
C31 a_592_n62# a_636_186# 0.045359f
C32 VDDA a_82_n552# 0.059058f
C33 VDDA a_636_n552# 0.053801f
C34 V_OSC a_636_186# 6.76e-20
C35 V_CONT a_1190_n552# 0.01611f
C36 V_CONT a_592_n62# 0.00118f
C37 a_38_n62# a_82_186# 0.048257f
C38 a_38_n62# a_82_n552# 0.043485f
C39 a_1190_n552# a_592_n62# 0.025048f
C40 a_38_n62# a_636_n552# 0.025048f
C41 V_CONT V_OSC 0.453326f
C42 a_82_186# a_636_186# 0.00532f
C43 a_1190_n552# GNDA 0.297521f
C44 a_636_n552# GNDA 0.418948f
C45 a_82_n552# GNDA 0.405917f
C46 V_CONT GNDA 1.51311f
C47 V_OSC GNDA 1.89306f
C48 a_592_n62# GNDA 0.484689f
C49 a_38_n62# GNDA 0.380768f
C50 a_1190_186# GNDA 0.204232f
C51 a_636_186# GNDA 0.088562f
C52 a_82_186# GNDA 0.05245f
C53 VDDA GNDA 10.900789f
C54 a_n746_764.t1 GNDA 0.153998f
C55 a_n746_764.t5 GNDA 0.465957f
C56 a_n746_764.t3 GNDA 0.365904f
C57 a_n746_764.n0 GNDA 0.27731f
C58 a_n746_764.t4 GNDA 0.365904f
C59 a_n746_764.n1 GNDA 0.276948f
C60 a_n746_764.t0 GNDA 0.518928f
C61 a_n746_764.n2 GNDA 0.237652f
C62 a_n746_764.t2 GNDA 0.137401f
C63 VDDA.t1 GNDA 0.009925f
C64 VDDA.t16 GNDA 0.022852f
C65 VDDA.t0 GNDA 0.195936f
C66 VDDA.t7 GNDA 0.003143f
C67 VDDA.t15 GNDA 0.191046f
C68 VDDA.t2 GNDA 0.192792f
C69 VDDA.t6 GNDA 0.003143f
C70 VDDA.t11 GNDA 0.055882f
C71 VDDA.t13 GNDA 0.444959f
C72 VDDA.t9 GNDA 0.194189f
C73 VDDA.t8 GNDA 0.003143f
C74 VDDA.t4 GNDA 0.137609f
C75 VDDA.n0 GNDA 0.184775f
C76 VDDA.t19 GNDA 9.62e-19
C77 VDDA.t17 GNDA 0.006605f
C78 VDDA.n1 GNDA 0.008774f
C79 VDDA.t18 GNDA 0.004266f
C80 VDDA.n2 GNDA 0.015998f
C81 VDDA.t3 GNDA 0.009777f
C82 VDDA.n3 GNDA 0.023552f
C83 VDDA.t12 GNDA 0.022852f
C84 VDDA.t5 GNDA 0.009803f
C85 VDDA.t10 GNDA 0.022852f
C86 VDDA.t14 GNDA 0.022852f
.ends

