magic
tech sky130A
timestamp 1737638164
<< nmos >>
rect -216 160 -194 203
rect -144 160 -122 203
rect -72 160 -50 203
rect 0 160 22 203
rect 72 160 94 203
rect 144 160 166 203
rect 0 0 22 43
rect 72 0 94 43
rect 144 0 166 43
<< ndiff >>
rect -266 195 -216 203
rect -266 170 -251 195
rect -231 170 -216 195
rect -266 160 -216 170
rect -194 195 -144 203
rect -194 170 -179 195
rect -159 170 -144 195
rect -194 160 -144 170
rect -122 195 -72 203
rect -122 170 -107 195
rect -87 170 -72 195
rect -122 160 -72 170
rect -50 195 0 203
rect -50 170 -35 195
rect -15 170 0 195
rect -50 160 0 170
rect 22 195 72 203
rect 22 170 37 195
rect 57 170 72 195
rect 22 160 72 170
rect 94 195 144 203
rect 94 170 109 195
rect 129 170 144 195
rect 94 160 144 170
rect 166 195 216 203
rect 166 170 181 195
rect 201 170 216 195
rect 166 160 216 170
rect -50 35 0 43
rect -50 10 -35 35
rect -15 10 0 35
rect -50 0 0 10
rect 22 35 72 43
rect 22 10 37 35
rect 57 10 72 35
rect 22 0 72 10
rect 94 35 144 43
rect 94 10 109 35
rect 129 10 144 35
rect 94 0 144 10
rect 166 35 216 43
rect 166 10 181 35
rect 201 10 216 35
rect 166 0 216 10
<< ndiffc >>
rect -251 170 -231 195
rect -179 170 -159 195
rect -107 170 -87 195
rect -35 170 -15 195
rect 37 170 57 195
rect 109 170 129 195
rect 181 170 201 195
rect -35 10 -15 35
rect 37 10 57 35
rect 109 10 129 35
rect 181 10 201 35
<< poly >>
rect -216 203 -194 218
rect -144 203 -122 218
rect -72 203 -50 218
rect 0 203 22 218
rect 72 203 94 218
rect 144 203 166 218
rect -216 145 -194 160
rect -144 145 -122 160
rect -72 145 -50 160
rect 0 145 22 160
rect 72 145 94 160
rect 144 145 166 160
rect 0 43 22 58
rect 72 43 94 58
rect 144 43 166 58
rect 0 -15 22 0
rect 72 -15 94 0
rect 144 -15 166 0
<< locali >>
rect -261 223 211 243
rect -261 195 -221 223
rect -261 170 -251 195
rect -231 170 -221 195
rect -261 160 -221 170
rect -189 195 -149 203
rect -189 170 -179 195
rect -159 170 -149 195
rect -189 140 -149 170
rect -117 195 -77 203
rect -117 170 -107 195
rect -87 170 -77 195
rect -117 160 -77 170
rect -45 195 -5 203
rect -45 170 -35 195
rect -15 170 -5 195
rect -45 160 -5 170
rect 27 195 67 203
rect 27 170 37 195
rect 57 170 67 195
rect 27 160 67 170
rect 99 195 139 203
rect 99 170 109 195
rect 129 170 139 195
rect 99 140 139 170
rect 171 195 211 223
rect 171 170 181 195
rect 201 170 211 195
rect 171 160 211 170
rect -189 120 139 140
rect -45 35 -5 43
rect -45 10 -35 35
rect -15 10 -5 35
rect -45 0 -5 10
rect 27 35 67 43
rect 27 10 37 35
rect 57 10 67 35
rect 27 0 67 10
rect 99 35 139 43
rect 99 10 109 35
rect 129 10 139 35
rect 99 0 139 10
rect 171 35 211 43
rect 171 10 181 35
rect 201 10 211 35
rect 171 0 211 10
<< end >>
