magic
tech sky130A
timestamp 1738412368
<< nwell >>
rect 605 105 1145 210
<< nmos >>
rect 665 -35 680 15
rect 720 -35 735 15
rect 775 -35 790 15
rect 940 -35 955 15
rect 995 -35 1010 15
rect 1050 -35 1065 15
rect 1105 -35 1120 15
<< pmos >>
rect 665 125 680 175
rect 720 125 735 175
rect 845 125 860 175
rect 900 125 915 175
rect 1070 125 1085 175
<< ndiff >>
rect 625 0 665 15
rect 625 -20 635 0
rect 655 -20 665 0
rect 625 -35 665 -20
rect 680 0 720 15
rect 680 -20 690 0
rect 710 -20 720 0
rect 680 -35 720 -20
rect 735 0 775 15
rect 735 -20 745 0
rect 765 -20 775 0
rect 735 -35 775 -20
rect 790 0 830 15
rect 790 -20 800 0
rect 820 -20 830 0
rect 790 -35 830 -20
rect 900 0 940 15
rect 900 -20 910 0
rect 930 -20 940 0
rect 900 -35 940 -20
rect 955 0 995 15
rect 955 -20 965 0
rect 985 -20 995 0
rect 955 -35 995 -20
rect 1010 0 1050 15
rect 1010 -20 1020 0
rect 1040 -20 1050 0
rect 1010 -35 1050 -20
rect 1065 0 1105 15
rect 1065 -20 1075 0
rect 1095 -20 1105 0
rect 1065 -35 1105 -20
rect 1120 0 1160 15
rect 1120 -20 1130 0
rect 1150 -20 1160 0
rect 1120 -35 1160 -20
<< pdiff >>
rect 625 160 665 175
rect 625 140 635 160
rect 655 140 665 160
rect 625 125 665 140
rect 680 160 720 175
rect 680 140 690 160
rect 710 140 720 160
rect 680 125 720 140
rect 735 160 775 175
rect 735 140 745 160
rect 765 140 775 160
rect 735 125 775 140
rect 805 160 845 175
rect 805 140 815 160
rect 835 140 845 160
rect 805 125 845 140
rect 860 160 900 175
rect 860 140 870 160
rect 890 140 900 160
rect 860 125 900 140
rect 915 160 955 175
rect 915 140 925 160
rect 945 140 955 160
rect 915 125 955 140
rect 1030 160 1070 175
rect 1030 140 1040 160
rect 1060 140 1070 160
rect 1030 125 1070 140
rect 1085 160 1125 175
rect 1085 140 1095 160
rect 1115 140 1125 160
rect 1085 125 1125 140
<< ndiffc >>
rect 635 -20 655 0
rect 690 -20 710 0
rect 745 -20 765 0
rect 800 -20 820 0
rect 910 -20 930 0
rect 965 -20 985 0
rect 1020 -20 1040 0
rect 1075 -20 1095 0
rect 1130 -20 1150 0
<< pdiffc >>
rect 635 140 655 160
rect 690 140 710 160
rect 745 140 765 160
rect 815 140 835 160
rect 870 140 890 160
rect 925 140 945 160
rect 1040 140 1060 160
rect 1095 140 1115 160
<< psubdiff >>
rect 1190 0 1230 15
rect 1190 -20 1200 0
rect 1220 -20 1230 0
rect 1190 -35 1230 -20
<< nsubdiff >>
rect 990 160 1030 175
rect 990 140 1000 160
rect 1020 140 1030 160
rect 990 125 1030 140
<< psubdiffcont >>
rect 1200 -20 1220 0
<< nsubdiffcont >>
rect 1000 140 1020 160
<< poly >>
rect 820 220 860 230
rect 820 200 830 220
rect 850 200 860 220
rect 665 185 735 200
rect 820 190 860 200
rect 665 175 680 185
rect 720 175 735 185
rect 845 175 860 190
rect 900 175 915 190
rect 1070 175 1085 190
rect 665 70 680 125
rect 720 110 735 125
rect 845 115 860 125
rect 760 100 860 115
rect 900 110 915 125
rect 1070 110 1085 125
rect 885 100 925 110
rect 760 85 775 100
rect 605 55 680 70
rect 665 15 680 55
rect 720 70 775 85
rect 885 80 895 100
rect 915 80 925 100
rect 885 70 925 80
rect 1050 95 1085 110
rect 720 15 735 70
rect 800 60 840 70
rect 800 40 810 60
rect 830 40 840 60
rect 1050 40 1065 95
rect 775 25 1065 40
rect 1090 60 1130 70
rect 1090 40 1100 60
rect 1120 40 1130 60
rect 1090 30 1130 40
rect 775 15 790 25
rect 940 15 955 25
rect 995 15 1010 25
rect 1050 15 1065 25
rect 1105 15 1120 30
rect 665 -50 680 -35
rect 720 -50 735 -35
rect 775 -50 790 -35
rect 940 -50 955 -35
rect 995 -50 1010 -35
rect 1050 -50 1065 -35
rect 1105 -50 1120 -35
<< polycont >>
rect 830 200 850 220
rect 895 80 915 100
rect 810 40 830 60
rect 1100 40 1120 60
<< locali >>
rect 820 220 860 230
rect 820 200 830 220
rect 850 210 860 220
rect 850 200 1115 210
rect 820 190 1115 200
rect 1095 170 1115 190
rect 630 160 660 170
rect 630 140 635 160
rect 655 140 660 160
rect 630 130 660 140
rect 685 160 715 170
rect 685 140 690 160
rect 710 140 715 160
rect 685 130 715 140
rect 740 160 770 170
rect 740 140 745 160
rect 765 140 770 160
rect 740 130 770 140
rect 810 160 840 170
rect 810 140 815 160
rect 835 140 840 160
rect 810 130 840 140
rect 865 160 895 170
rect 865 140 870 160
rect 890 140 895 160
rect 865 130 895 140
rect 920 160 965 170
rect 920 140 925 160
rect 945 140 965 160
rect 920 130 965 140
rect 995 160 1065 170
rect 995 140 1000 160
rect 1020 140 1040 160
rect 1060 140 1065 160
rect 995 130 1065 140
rect 1090 160 1120 170
rect 1090 140 1095 160
rect 1115 140 1175 160
rect 1090 130 1120 140
rect 635 50 655 130
rect 745 50 765 130
rect 815 110 835 130
rect 815 100 925 110
rect 815 90 895 100
rect 865 80 895 90
rect 915 80 925 100
rect 865 70 925 80
rect 800 60 840 70
rect 800 50 810 60
rect 635 40 810 50
rect 830 40 840 60
rect 635 30 840 40
rect 635 10 655 30
rect 865 10 885 70
rect 945 50 965 130
rect 1155 80 1175 140
rect 1090 60 1130 70
rect 1090 50 1100 60
rect 910 40 1100 50
rect 1120 40 1130 60
rect 910 30 1130 40
rect 1155 60 1230 80
rect 910 10 930 30
rect 1020 10 1040 30
rect 1155 10 1175 60
rect 630 0 660 10
rect 630 -20 635 0
rect 655 -20 660 0
rect 630 -30 660 -20
rect 685 0 715 10
rect 685 -20 690 0
rect 710 -20 715 0
rect 685 -30 715 -20
rect 740 0 770 10
rect 740 -20 745 0
rect 765 -20 770 0
rect 740 -30 770 -20
rect 795 0 885 10
rect 795 -20 800 0
rect 820 -10 885 0
rect 905 0 935 10
rect 820 -20 825 -10
rect 795 -30 825 -20
rect 905 -20 910 0
rect 930 -20 935 0
rect 905 -30 935 -20
rect 960 0 990 10
rect 960 -20 965 0
rect 985 -20 990 0
rect 960 -30 990 -20
rect 1015 0 1045 10
rect 1015 -20 1020 0
rect 1040 -20 1045 0
rect 1015 -30 1045 -20
rect 1070 0 1100 10
rect 1070 -20 1075 0
rect 1095 -20 1100 0
rect 1070 -30 1100 -20
rect 1125 0 1175 10
rect 1125 -20 1130 0
rect 1150 -20 1175 0
rect 1195 0 1225 10
rect 1195 -20 1200 0
rect 1220 -20 1225 0
rect 1125 -30 1155 -20
rect 1195 -30 1225 -20
<< viali >>
rect 690 140 710 160
rect 870 140 890 160
rect 1000 140 1020 160
rect 1040 140 1060 160
rect 690 -20 710 0
rect 965 -20 985 0
rect 1075 -20 1095 0
rect 1200 -20 1220 0
<< metal1 >>
rect 605 160 1145 175
rect 605 140 690 160
rect 710 140 870 160
rect 890 140 1000 160
rect 1020 140 1040 160
rect 1060 140 1145 160
rect 605 125 1145 140
rect 605 0 1230 15
rect 605 -20 690 0
rect 710 -20 965 0
rect 985 -20 1075 0
rect 1095 -20 1200 0
rect 1220 -20 1230 0
rect 605 -35 1230 -20
<< labels >>
flabel metal1 605 150 605 150 7 FreeSans 160 0 -80 0 VDDA
flabel metal1 605 -10 605 -10 7 FreeSans 160 0 -80 0 GNDA
flabel poly 605 60 605 60 7 FreeSans 160 0 -80 0 VIN
flabel locali 965 80 965 80 3 FreeSans 160 0 80 0 C
flabel locali 1230 70 1230 70 3 FreeSans 160 0 80 0 VOUT
flabel locali 700 50 700 50 1 FreeSans 160 0 0 80 CLK
flabel locali 755 -30 755 -30 5 FreeSans 160 0 0 -80 B
flabel locali 885 55 885 55 3 FreeSans 160 0 80 0 A
<< end >>
