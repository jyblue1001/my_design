magic
tech sky130A
timestamp 1738233458
<< nwell >>
rect 990 130 2040 650
<< nmos >>
rect 1060 -175 1075 -125
rect 1125 -175 1140 -125
rect 1190 -175 1205 -125
rect 1255 -175 1270 -125
rect 1420 -175 1435 -125
rect 1485 -175 1500 -125
rect 1550 -175 1565 -125
rect 1615 -175 1630 -125
rect 1760 -175 1775 -125
rect 1825 -175 1840 -125
rect 1890 -175 1905 -125
rect 1955 -175 1970 -125
rect 1570 -555 1620 -305
rect 1670 -555 1720 -305
rect 1770 -555 1820 -305
rect 1870 -555 1920 -305
<< pmos >>
rect 1075 345 1125 595
rect 1175 345 1225 595
rect 1275 345 1325 595
rect 1375 345 1425 595
rect 1475 345 1525 595
rect 1575 345 1625 595
rect 1675 345 1725 595
rect 1775 345 1825 595
rect 1060 155 1075 255
rect 1125 155 1140 255
rect 1190 155 1205 255
rect 1255 155 1270 255
rect 1420 155 1435 255
rect 1485 155 1500 255
rect 1550 155 1565 255
rect 1615 155 1630 255
rect 1760 155 1775 255
rect 1825 155 1840 255
rect 1890 155 1905 255
rect 1955 155 1970 255
<< ndiff >>
rect 1010 -140 1060 -125
rect 1010 -160 1025 -140
rect 1045 -160 1060 -140
rect 1010 -175 1060 -160
rect 1075 -140 1125 -125
rect 1075 -160 1090 -140
rect 1110 -160 1125 -140
rect 1075 -175 1125 -160
rect 1140 -140 1190 -125
rect 1140 -160 1155 -140
rect 1175 -160 1190 -140
rect 1140 -175 1190 -160
rect 1205 -140 1255 -125
rect 1205 -160 1220 -140
rect 1240 -160 1255 -140
rect 1205 -175 1255 -160
rect 1270 -140 1320 -125
rect 1270 -160 1285 -140
rect 1305 -160 1320 -140
rect 1270 -175 1320 -160
rect 1370 -140 1420 -125
rect 1370 -160 1385 -140
rect 1405 -160 1420 -140
rect 1370 -175 1420 -160
rect 1435 -140 1485 -125
rect 1435 -160 1450 -140
rect 1470 -160 1485 -140
rect 1435 -175 1485 -160
rect 1500 -140 1550 -125
rect 1500 -160 1515 -140
rect 1535 -160 1550 -140
rect 1500 -175 1550 -160
rect 1565 -140 1615 -125
rect 1565 -160 1580 -140
rect 1600 -160 1615 -140
rect 1565 -175 1615 -160
rect 1630 -140 1680 -125
rect 1630 -160 1645 -140
rect 1665 -160 1680 -140
rect 1630 -175 1680 -160
rect 1710 -140 1760 -125
rect 1710 -160 1725 -140
rect 1745 -160 1760 -140
rect 1710 -175 1760 -160
rect 1775 -140 1825 -125
rect 1775 -160 1790 -140
rect 1810 -160 1825 -140
rect 1775 -175 1825 -160
rect 1840 -140 1890 -125
rect 1840 -160 1855 -140
rect 1875 -160 1890 -140
rect 1840 -175 1890 -160
rect 1905 -140 1955 -125
rect 1905 -160 1920 -140
rect 1940 -160 1955 -140
rect 1905 -175 1955 -160
rect 1970 -140 2020 -125
rect 1970 -160 1985 -140
rect 2005 -160 2020 -140
rect 1970 -175 2020 -160
rect 1520 -320 1570 -305
rect 1520 -540 1535 -320
rect 1555 -540 1570 -320
rect 1520 -555 1570 -540
rect 1620 -320 1670 -305
rect 1620 -540 1635 -320
rect 1655 -540 1670 -320
rect 1620 -555 1670 -540
rect 1720 -320 1770 -305
rect 1720 -540 1735 -320
rect 1755 -540 1770 -320
rect 1720 -555 1770 -540
rect 1820 -320 1870 -305
rect 1820 -540 1835 -320
rect 1855 -540 1870 -320
rect 1820 -555 1870 -540
rect 1920 -320 1970 -305
rect 1920 -540 1935 -320
rect 1955 -540 1970 -320
rect 1920 -555 1970 -540
<< pdiff >>
rect 1025 580 1075 595
rect 1025 360 1040 580
rect 1060 360 1075 580
rect 1025 345 1075 360
rect 1125 580 1175 595
rect 1125 360 1140 580
rect 1160 360 1175 580
rect 1125 345 1175 360
rect 1225 580 1275 595
rect 1225 360 1240 580
rect 1260 360 1275 580
rect 1225 345 1275 360
rect 1325 580 1375 595
rect 1325 360 1340 580
rect 1360 360 1375 580
rect 1325 345 1375 360
rect 1425 580 1475 595
rect 1425 360 1440 580
rect 1460 360 1475 580
rect 1425 345 1475 360
rect 1525 580 1575 595
rect 1525 360 1540 580
rect 1560 360 1575 580
rect 1525 345 1575 360
rect 1625 580 1675 595
rect 1625 360 1640 580
rect 1660 360 1675 580
rect 1625 345 1675 360
rect 1725 580 1775 595
rect 1725 360 1740 580
rect 1760 360 1775 580
rect 1725 345 1775 360
rect 1825 580 1875 595
rect 1825 360 1840 580
rect 1860 360 1875 580
rect 1825 345 1875 360
rect 1010 240 1060 255
rect 1010 170 1025 240
rect 1045 170 1060 240
rect 1010 155 1060 170
rect 1075 240 1125 255
rect 1075 170 1090 240
rect 1110 170 1125 240
rect 1075 155 1125 170
rect 1140 240 1190 255
rect 1140 170 1155 240
rect 1175 170 1190 240
rect 1140 155 1190 170
rect 1205 240 1255 255
rect 1205 170 1220 240
rect 1240 170 1255 240
rect 1205 155 1255 170
rect 1270 240 1320 255
rect 1270 170 1285 240
rect 1305 170 1320 240
rect 1270 155 1320 170
rect 1370 240 1420 255
rect 1370 170 1385 240
rect 1405 170 1420 240
rect 1370 155 1420 170
rect 1435 240 1485 255
rect 1435 170 1450 240
rect 1470 170 1485 240
rect 1435 155 1485 170
rect 1500 240 1550 255
rect 1500 170 1515 240
rect 1535 170 1550 240
rect 1500 155 1550 170
rect 1565 240 1615 255
rect 1565 170 1580 240
rect 1600 170 1615 240
rect 1565 155 1615 170
rect 1630 240 1680 255
rect 1630 170 1645 240
rect 1665 170 1680 240
rect 1630 155 1680 170
rect 1710 240 1760 255
rect 1710 170 1725 240
rect 1745 170 1760 240
rect 1710 155 1760 170
rect 1775 240 1825 255
rect 1775 170 1790 240
rect 1810 170 1825 240
rect 1775 155 1825 170
rect 1840 240 1890 255
rect 1840 170 1855 240
rect 1875 170 1890 240
rect 1840 155 1890 170
rect 1905 240 1955 255
rect 1905 170 1920 240
rect 1940 170 1955 240
rect 1905 155 1955 170
rect 1970 240 2020 255
rect 1970 170 1985 240
rect 2005 170 2020 240
rect 1970 155 2020 170
<< ndiffc >>
rect 1025 -160 1045 -140
rect 1090 -160 1110 -140
rect 1155 -160 1175 -140
rect 1220 -160 1240 -140
rect 1285 -160 1305 -140
rect 1385 -160 1405 -140
rect 1450 -160 1470 -140
rect 1515 -160 1535 -140
rect 1580 -160 1600 -140
rect 1645 -160 1665 -140
rect 1725 -160 1745 -140
rect 1790 -160 1810 -140
rect 1855 -160 1875 -140
rect 1920 -160 1940 -140
rect 1985 -160 2005 -140
rect 1535 -540 1555 -320
rect 1635 -540 1655 -320
rect 1735 -540 1755 -320
rect 1835 -540 1855 -320
rect 1935 -540 1955 -320
<< pdiffc >>
rect 1040 360 1060 580
rect 1140 360 1160 580
rect 1240 360 1260 580
rect 1340 360 1360 580
rect 1440 360 1460 580
rect 1540 360 1560 580
rect 1640 360 1660 580
rect 1740 360 1760 580
rect 1840 360 1860 580
rect 1025 170 1045 240
rect 1090 170 1110 240
rect 1155 170 1175 240
rect 1220 170 1240 240
rect 1285 170 1305 240
rect 1385 170 1405 240
rect 1450 170 1470 240
rect 1515 170 1535 240
rect 1580 170 1600 240
rect 1645 170 1665 240
rect 1725 170 1745 240
rect 1790 170 1810 240
rect 1855 170 1875 240
rect 1920 170 1940 240
rect 1985 170 2005 240
<< psubdiff >>
rect 1140 -220 1190 -205
rect 1140 -240 1155 -220
rect 1175 -240 1190 -220
rect 1140 -255 1190 -240
rect 1200 -690 1250 -640
rect 1970 -705 2020 -655
<< nsubdiff >>
rect 1920 580 1970 595
rect 1920 360 1935 580
rect 1955 360 1970 580
rect 1920 345 1970 360
<< psubdiffcont >>
rect 1155 -240 1175 -220
<< nsubdiffcont >>
rect 1935 360 1955 580
<< poly >>
rect 1055 640 1095 650
rect 1055 620 1065 640
rect 1085 620 1095 640
rect 1430 640 1470 650
rect 1430 620 1440 640
rect 1460 620 1470 640
rect 1810 640 1850 650
rect 1810 620 1820 640
rect 1840 620 1850 640
rect 1055 610 1850 620
rect 1075 605 1825 610
rect 1075 595 1125 605
rect 1175 595 1225 605
rect 1275 595 1325 605
rect 1375 595 1425 605
rect 1475 595 1525 605
rect 1575 595 1625 605
rect 1675 595 1725 605
rect 1775 595 1825 605
rect 1075 330 1125 345
rect 1175 330 1225 345
rect 1275 330 1325 345
rect 1375 330 1425 345
rect 1475 330 1525 345
rect 1575 330 1625 345
rect 1675 330 1725 345
rect 1775 330 1825 345
rect 735 265 1140 280
rect 750 -30 765 265
rect 1060 255 1075 265
rect 1125 255 1140 265
rect 1190 255 1205 270
rect 1255 255 1270 270
rect 1420 255 1435 270
rect 1485 255 1500 270
rect 1550 255 1565 270
rect 1615 255 1630 270
rect 1760 255 1775 270
rect 1825 255 1840 270
rect 1890 255 1905 270
rect 1955 255 1970 270
rect 2065 155 2105 165
rect 1060 140 1075 155
rect 1125 140 1140 155
rect 1190 115 1205 155
rect 1255 115 1270 155
rect 1420 145 1435 155
rect 1485 145 1500 155
rect 1550 145 1565 155
rect 1615 145 1630 155
rect 1420 140 1630 145
rect 1760 145 1775 155
rect 1825 145 1840 155
rect 1890 145 1905 155
rect 1955 145 1970 155
rect 2065 145 2075 155
rect 1390 130 1665 140
rect 815 105 1365 115
rect 815 100 1335 105
rect 1325 85 1335 100
rect 1355 85 1365 105
rect 1390 110 1400 130
rect 1420 125 1635 130
rect 1420 110 1430 125
rect 1390 100 1430 110
rect 1625 110 1635 125
rect 1655 110 1665 130
rect 1625 100 1665 110
rect 1760 135 2075 145
rect 2095 135 2105 155
rect 1760 130 2105 135
rect 1760 110 1770 130
rect 1790 110 1800 130
rect 2065 125 2105 130
rect 1760 100 1800 110
rect 1325 75 1365 85
rect 1155 25 1195 35
rect 1155 5 1165 25
rect 1185 10 1195 25
rect 1185 5 1775 10
rect 1155 -5 1775 5
rect 750 -45 1500 -30
rect 1025 -80 1065 -70
rect 1025 -100 1035 -80
rect 1055 -95 1065 -80
rect 1265 -80 1305 -70
rect 1265 -95 1275 -80
rect 1055 -100 1275 -95
rect 1295 -100 1305 -80
rect 1025 -110 1305 -100
rect 1060 -115 1270 -110
rect 1060 -125 1075 -115
rect 1125 -125 1140 -115
rect 1190 -125 1205 -115
rect 1255 -125 1270 -115
rect 1420 -125 1435 -45
rect 1485 -125 1500 -45
rect 1760 -100 1775 -5
rect 1550 -125 1565 -110
rect 1615 -125 1630 -110
rect 1760 -115 2105 -100
rect 1760 -125 1775 -115
rect 1825 -125 1840 -115
rect 1890 -125 1905 -115
rect 1955 -125 1970 -115
rect 1060 -190 1075 -175
rect 1125 -190 1140 -175
rect 1190 -190 1205 -175
rect 1255 -190 1270 -175
rect 1420 -190 1435 -175
rect 1485 -190 1500 -175
rect 1315 -210 1355 -200
rect 1315 -230 1325 -210
rect 1345 -215 1355 -210
rect 1550 -215 1565 -175
rect 1615 -215 1630 -175
rect 1760 -190 1775 -175
rect 1825 -190 1840 -175
rect 1890 -190 1905 -175
rect 1955 -190 1970 -175
rect 1345 -230 1630 -215
rect 1315 -240 1355 -230
rect 2090 -265 2105 -115
rect 2065 -275 2105 -265
rect 1570 -305 1620 -290
rect 1670 -305 1720 -290
rect 1770 -305 1820 -290
rect 1870 -305 1920 -290
rect 2065 -295 2075 -275
rect 2095 -295 2105 -275
rect 2065 -305 2105 -295
rect 1570 -565 1620 -555
rect 1670 -565 1720 -555
rect 1770 -565 1820 -555
rect 1870 -565 1920 -555
rect 1570 -575 1920 -565
rect 1570 -580 1585 -575
rect 1575 -595 1585 -580
rect 1605 -580 1885 -575
rect 1605 -595 1615 -580
rect 1575 -605 1615 -595
rect 1875 -595 1885 -580
rect 1905 -580 1920 -575
rect 1905 -595 1915 -580
rect 1875 -605 1915 -595
<< polycont >>
rect 1065 620 1085 640
rect 1440 620 1460 640
rect 1820 620 1840 640
rect 1335 85 1355 105
rect 1400 110 1420 130
rect 1635 110 1655 130
rect 2075 135 2095 155
rect 1770 110 1790 130
rect 1165 5 1185 25
rect 1035 -100 1055 -80
rect 1275 -100 1295 -80
rect 1325 -230 1345 -210
rect 2075 -295 2095 -275
rect 1585 -595 1605 -575
rect 1885 -595 1905 -575
<< xpolycontact >>
rect 2070 533 2105 753
rect 2070 215 2105 435
rect 990 -590 1210 -305
rect 1245 -590 1465 -305
rect 2070 -640 2105 -420
rect 2070 -930 2105 -710
<< xpolyres >>
rect 2070 435 2105 533
rect 1210 -590 1245 -305
rect 2070 -710 2105 -640
<< locali >>
rect 2125 1080 2175 1090
rect 2125 1070 2135 1080
rect 2085 1050 2135 1070
rect 2165 1050 2175 1080
rect 2085 753 2105 1050
rect 2125 1040 2175 1050
rect 1055 640 1095 650
rect 1055 635 1065 640
rect 920 620 1065 635
rect 1085 635 1095 640
rect 1430 640 1470 650
rect 1430 635 1440 640
rect 1085 620 1440 635
rect 1460 635 1470 640
rect 1810 640 1850 650
rect 1810 635 1820 640
rect 1460 620 1820 635
rect 1840 635 1850 640
rect 1840 620 1860 635
rect 920 615 1860 620
rect 920 -305 940 615
rect 1040 610 1095 615
rect 1430 610 1470 615
rect 1810 610 1860 615
rect 1040 590 1060 610
rect 1440 590 1460 610
rect 1840 590 1860 610
rect 1025 580 1070 590
rect 1025 360 1040 580
rect 1060 360 1070 580
rect 1025 350 1070 360
rect 1130 580 1170 590
rect 1130 360 1140 580
rect 1160 360 1170 580
rect 1130 350 1170 360
rect 1230 580 1270 590
rect 1230 360 1240 580
rect 1260 360 1270 580
rect 1230 350 1270 360
rect 1330 580 1370 590
rect 1330 360 1340 580
rect 1360 360 1370 580
rect 1330 350 1370 360
rect 1430 580 1470 590
rect 1430 360 1440 580
rect 1460 360 1470 580
rect 1430 350 1470 360
rect 1530 580 1570 590
rect 1530 360 1540 580
rect 1560 360 1570 580
rect 1530 350 1570 360
rect 1630 580 1670 590
rect 1630 360 1640 580
rect 1660 360 1670 580
rect 1630 350 1670 360
rect 1730 580 1770 590
rect 1730 360 1740 580
rect 1760 360 1770 580
rect 1730 350 1770 360
rect 1830 580 1870 590
rect 1830 360 1840 580
rect 1860 360 1870 580
rect 1830 350 1870 360
rect 1925 580 1965 590
rect 1925 360 1935 580
rect 1955 360 1965 580
rect 1925 350 1965 360
rect 1240 330 1260 350
rect 1640 330 1660 350
rect 1105 310 1660 330
rect 1105 290 1125 310
rect 1025 270 1305 290
rect 1025 250 1045 270
rect 1155 250 1175 270
rect 1285 250 1305 270
rect 1725 270 2005 290
rect 1725 250 1745 270
rect 1855 250 1875 270
rect 1985 250 2005 270
rect 1015 240 1055 250
rect 1015 170 1025 240
rect 1045 170 1055 240
rect 1015 160 1055 170
rect 1080 240 1120 250
rect 1080 170 1090 240
rect 1110 170 1120 240
rect 1080 160 1120 170
rect 1145 240 1185 250
rect 1145 170 1155 240
rect 1175 170 1185 240
rect 1145 160 1185 170
rect 1210 240 1250 250
rect 1210 170 1220 240
rect 1240 170 1250 240
rect 1210 160 1250 170
rect 1275 240 1320 250
rect 1275 170 1285 240
rect 1305 170 1320 240
rect 1275 160 1320 170
rect 1375 240 1415 250
rect 1375 170 1385 240
rect 1405 170 1415 240
rect 1375 160 1415 170
rect 1440 240 1480 250
rect 1440 170 1450 240
rect 1470 170 1480 240
rect 1440 160 1480 170
rect 1505 240 1545 250
rect 1505 170 1515 240
rect 1535 170 1545 240
rect 1505 160 1545 170
rect 1570 240 1615 250
rect 1570 170 1580 240
rect 1600 170 1615 240
rect 1570 160 1615 170
rect 1635 240 1675 250
rect 1635 170 1645 240
rect 1665 170 1675 240
rect 1635 160 1675 170
rect 1715 240 1755 250
rect 1715 170 1725 240
rect 1745 170 1755 240
rect 1715 160 1755 170
rect 1780 240 1820 250
rect 1780 170 1790 240
rect 1810 170 1820 240
rect 1780 160 1820 170
rect 1845 240 1885 250
rect 1845 170 1855 240
rect 1875 170 1885 240
rect 1845 160 1885 170
rect 1910 240 1950 250
rect 1910 170 1920 240
rect 1940 170 1950 240
rect 1910 160 1950 170
rect 1975 240 2015 250
rect 1975 170 1985 240
rect 2005 170 2015 240
rect 1975 160 2015 170
rect 2070 165 2090 215
rect 1090 75 1110 160
rect 1220 75 1240 160
rect 1385 140 1410 160
rect 1390 130 1430 140
rect 1325 105 1365 115
rect 1325 85 1335 105
rect 1355 85 1365 105
rect 1390 110 1400 130
rect 1420 110 1430 130
rect 1390 100 1430 110
rect 1325 75 1365 85
rect 1395 75 1415 100
rect 1035 50 1110 75
rect 1165 55 1240 75
rect 1035 -70 1055 50
rect 1165 35 1185 55
rect 1155 25 1195 35
rect 1155 5 1165 25
rect 1185 5 1195 25
rect 1155 -5 1195 5
rect 1025 -80 1065 -70
rect 1025 -100 1035 -80
rect 1055 -100 1065 -80
rect 1025 -110 1065 -100
rect 1025 -130 1045 -110
rect 1155 -130 1175 -5
rect 1265 -80 1305 -70
rect 1265 -100 1275 -80
rect 1295 -100 1305 -80
rect 1265 -110 1305 -100
rect 1285 -130 1305 -110
rect 1015 -140 1055 -130
rect 1015 -160 1025 -140
rect 1045 -160 1055 -140
rect 1015 -170 1055 -160
rect 1080 -140 1120 -130
rect 1080 -160 1090 -140
rect 1110 -160 1120 -140
rect 1080 -170 1120 -160
rect 1145 -140 1185 -130
rect 1145 -160 1155 -140
rect 1175 -160 1185 -140
rect 1145 -170 1185 -160
rect 1210 -140 1250 -130
rect 1210 -160 1220 -140
rect 1240 -160 1250 -140
rect 1210 -170 1250 -160
rect 1275 -140 1315 -130
rect 1275 -160 1285 -140
rect 1305 -160 1315 -140
rect 1275 -170 1315 -160
rect 1090 -220 1110 -170
rect 1145 -220 1185 -210
rect 1220 -220 1240 -170
rect 1335 -200 1355 75
rect 1395 55 1470 75
rect 1450 -130 1470 55
rect 1515 65 1535 160
rect 1645 140 1665 160
rect 1625 130 1665 140
rect 1625 110 1635 130
rect 1655 110 1665 130
rect 1625 100 1665 110
rect 1760 130 1800 140
rect 1760 110 1770 130
rect 1790 110 1800 130
rect 1760 100 1800 110
rect 1760 65 1780 100
rect 1515 45 1780 65
rect 1580 -130 1600 45
rect 1985 30 2005 160
rect 2065 155 2105 165
rect 2065 135 2075 155
rect 2095 135 2105 155
rect 2065 125 2105 135
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 30 2145 70
rect 1985 10 2285 30
rect 2265 -10 2285 10
rect 2265 -30 3385 -10
rect 2265 -50 2285 -30
rect 1985 -70 2285 -50
rect 1985 -130 2005 -70
rect 2125 -125 2145 -70
rect 1375 -140 1415 -130
rect 1375 -160 1385 -140
rect 1405 -160 1415 -140
rect 1375 -170 1415 -160
rect 1440 -140 1480 -130
rect 1440 -160 1450 -140
rect 1470 -160 1480 -140
rect 1440 -170 1480 -160
rect 1505 -140 1545 -130
rect 1505 -160 1515 -140
rect 1535 -160 1545 -140
rect 1505 -170 1545 -160
rect 1570 -140 1610 -130
rect 1570 -160 1580 -140
rect 1600 -160 1610 -140
rect 1570 -170 1610 -160
rect 1635 -140 1675 -130
rect 1635 -160 1645 -140
rect 1665 -160 1675 -140
rect 1635 -170 1675 -160
rect 1715 -140 1755 -130
rect 1715 -160 1725 -140
rect 1745 -160 1755 -140
rect 1715 -170 1755 -160
rect 1780 -140 1820 -130
rect 1780 -160 1790 -140
rect 1810 -160 1820 -140
rect 1780 -170 1820 -160
rect 1845 -140 1885 -130
rect 1845 -160 1855 -140
rect 1875 -160 1885 -140
rect 1845 -170 1885 -160
rect 1910 -140 1950 -130
rect 1910 -160 1920 -140
rect 1940 -160 1950 -140
rect 1910 -170 1950 -160
rect 1975 -140 2015 -130
rect 1975 -160 1985 -140
rect 2005 -160 2015 -140
rect 1975 -170 2015 -160
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 1090 -240 1155 -220
rect 1175 -240 1240 -220
rect 1315 -210 1355 -200
rect 1385 -190 1405 -170
rect 1515 -190 1535 -170
rect 1645 -190 1665 -170
rect 1385 -210 1665 -190
rect 1725 -190 1745 -170
rect 1855 -190 1875 -170
rect 1985 -190 2005 -170
rect 2125 -180 2180 -170
rect 1315 -230 1325 -210
rect 1345 -230 1355 -210
rect 1315 -240 1355 -230
rect 1145 -250 1185 -240
rect 1515 -270 1535 -210
rect 1725 -215 2005 -190
rect 1515 -290 1755 -270
rect 920 -325 990 -305
rect 1735 -310 1755 -290
rect 2065 -275 2105 -265
rect 2065 -295 2075 -275
rect 2095 -295 2105 -275
rect 2065 -305 2105 -295
rect 1525 -320 1565 -310
rect 1525 -540 1535 -320
rect 1555 -540 1565 -320
rect 1525 -550 1565 -540
rect 1625 -320 1665 -310
rect 1625 -540 1635 -320
rect 1655 -540 1665 -320
rect 1625 -550 1665 -540
rect 1725 -320 1765 -310
rect 1725 -540 1735 -320
rect 1755 -540 1765 -320
rect 1725 -550 1765 -540
rect 1825 -320 1865 -310
rect 1825 -540 1835 -320
rect 1855 -540 1865 -320
rect 1825 -550 1865 -540
rect 1925 -320 1965 -310
rect 1925 -540 1935 -320
rect 1955 -540 1965 -320
rect 2085 -420 2105 -305
rect 1925 -550 1965 -540
rect 1535 -570 1555 -550
rect 1575 -570 1615 -565
rect 1875 -570 1915 -565
rect 1935 -570 1955 -550
rect 1465 -575 1955 -570
rect 1465 -590 1585 -575
rect 1575 -595 1585 -590
rect 1605 -590 1885 -575
rect 1605 -595 1615 -590
rect 1575 -605 1615 -595
rect 1875 -595 1885 -590
rect 1905 -590 1955 -575
rect 1905 -595 1915 -590
rect 1875 -605 1915 -595
rect 1205 -655 1245 -645
rect 1205 -675 1215 -655
rect 1235 -675 1245 -655
rect 1205 -685 1245 -675
rect 1975 -670 2015 -660
rect 1975 -690 1985 -670
rect 2005 -690 2015 -670
rect 1975 -700 2015 -690
rect 2085 -1105 2105 -930
rect 2125 -1105 2175 -1095
rect 2085 -1125 2135 -1105
rect 2125 -1135 2135 -1125
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< viali >>
rect 2135 1050 2165 1080
rect 1140 360 1160 580
rect 1340 360 1360 580
rect 1540 360 1560 580
rect 1740 360 1760 580
rect 1935 360 1955 580
rect 1450 170 1470 240
rect 1580 170 1600 240
rect 1790 170 1810 240
rect 1920 170 1940 240
rect 1090 -160 1110 -140
rect 1220 -160 1240 -140
rect 2135 80 2170 115
rect 1790 -160 1810 -140
rect 1920 -160 1940 -140
rect 2135 -170 2170 -135
rect 1155 -240 1175 -220
rect 1635 -540 1655 -320
rect 1835 -540 1855 -320
rect 1215 -675 1235 -655
rect 1985 -690 2005 -670
rect 2135 -1135 2165 -1105
<< metal1 >>
rect 2125 1080 2175 1090
rect 2125 1050 2135 1080
rect 2165 1050 2175 1080
rect 2125 1040 2175 1050
rect 960 580 2040 650
rect 960 360 1140 580
rect 1160 360 1340 580
rect 1360 360 1540 580
rect 1560 360 1740 580
rect 1760 360 1935 580
rect 1955 360 2040 580
rect 960 240 2040 360
rect 960 170 1450 240
rect 1470 170 1580 240
rect 1600 170 1790 240
rect 1810 170 1920 240
rect 1940 170 2040 240
rect 960 130 2040 170
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 970 -140 2040 -85
rect 970 -160 1090 -140
rect 1110 -160 1220 -140
rect 1240 -160 1790 -140
rect 1810 -160 1920 -140
rect 1940 -160 2040 -140
rect 970 -220 2040 -160
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 970 -240 1155 -220
rect 1175 -240 2040 -220
rect 970 -320 2040 -240
rect 970 -540 1635 -320
rect 1655 -540 1835 -320
rect 1855 -540 2040 -320
rect 970 -655 2040 -540
rect 970 -675 1215 -655
rect 1235 -670 2040 -655
rect 1235 -675 1985 -670
rect 970 -690 1985 -675
rect 2005 -690 2040 -670
rect 970 -715 2040 -690
rect 2125 -1105 2175 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< via1 >>
rect 2135 1050 2165 1080
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -1135 2165 -1105
<< metal2 >>
rect 2125 1080 2175 1090
rect 2125 1050 2135 1080
rect 2165 1050 2175 1080
rect 2125 1040 2175 1050
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2125 -1105 2175 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< via2 >>
rect 2135 1050 2165 1080
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -1135 2165 -1105
<< metal3 >>
rect 2125 1085 2175 1090
rect 2125 1080 3330 1085
rect 2125 1050 2135 1080
rect 2165 1050 3330 1080
rect 2125 1040 3330 1050
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2300 55 3330 1040
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2300 -1095 3330 -110
rect 2125 -1105 3330 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 3330 -1105
rect 2125 -1140 3330 -1135
rect 2125 -1145 2175 -1140
<< via3 >>
rect 2135 80 2170 115
rect 2135 -170 2170 -135
<< mimcap >>
rect 2315 115 3315 1070
rect 2315 80 2325 115
rect 2360 80 3315 115
rect 2315 70 3315 80
rect 2315 -135 3315 -125
rect 2315 -170 2325 -135
rect 2360 -170 3315 -135
rect 2315 -1125 3315 -170
<< mimcapcontact >>
rect 2325 80 2360 115
rect 2325 -170 2360 -135
<< metal4 >>
rect 2125 115 2365 125
rect 2125 80 2135 115
rect 2170 80 2325 115
rect 2360 80 2365 115
rect 2125 70 2365 80
rect 2125 -135 2365 -125
rect 2125 -170 2135 -135
rect 2170 -170 2325 -135
rect 2360 -170 2365 -135
rect 2125 -180 2365 -170
<< labels >>
flabel metal1 960 355 960 355 7 FreeSans 400 0 0 0 VDDA
flabel metal1 970 -330 970 -330 7 FreeSans 400 0 0 0 GNDA
flabel locali 920 495 920 495 7 FreeSans 160 0 -80 0 p_bias
flabel locali 1500 -590 1500 -590 5 FreeSans 160 0 0 -80 n_bias
flabel locali 1755 -270 1755 -270 2 FreeSans 160 0 80 80 v_common_n
flabel locali 1660 310 1660 310 4 FreeSans 160 0 80 -80 v_common_p
flabel locali 1780 45 1780 45 3 FreeSans 160 0 160 80 n_right
flabel poly 1775 10 1775 10 3 FreeSans 160 0 160 -80 p_right
flabel locali 1035 40 1035 40 7 FreeSans 160 0 -80 0 p_left
flabel locali 1450 40 1450 40 7 FreeSans 160 0 -80 0 n_left
flabel locali 3385 -21 3385 -21 3 FreeSans 80 0 40 0 VOUT
flabel poly 735 270 735 270 7 FreeSans 400 0 -200 0 VIN+
flabel poly 815 105 815 105 7 FreeSans 400 0 -200 0 VIN-
<< end >>
