** sch_path: /foss/designs/my_design/projects/pll/full_pll/magic/tb_pll_bgr_magic.sch
**.subckt tb_pll_bgr_magic
V1 VDD GND 1.8
V2 F_REF GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
x1 V_OSC VDD GND F_REF pll_bgr_magic
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.include /foss/designs/my_design/projects/pll/full_pll/magic/pll_bgr_magic.spice

.option method=gear
* .option method=trap
.option wnflag=1
* .option savecurrents

.save
+v(x1.v_cont.n0)
+v(x1.f_vco.t0)
+v(x1.pfd_8_0.qa.n0)
+v(x1.pfd_8_0.qb.n0)
+v(x1.pfd_8_0.up_input.n0)
+v(x1.pfd_8_0.down_input.n0)
+v(x1.charge_pump_cell_6_0.x.n0)
+v(x1.vco_fd_magic_0.div120_2_0.div2.n0)
+v(x1.vco_fd_magic_0.div120_2_0.div4.n0)
+v(x1.vco_fd_magic_0.div120_2_0.div8.n0)
+v(x1.vco_fd_magic_0.div120_2_0.div24.n0)
+@m.x1.x58.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x124.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x160.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x161.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x214.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x255.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x382.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x424.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x430.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x463.msky130_fd_pr__pfet_01v8[id]

* V_out initial voltage

.ic v(x1.v_cont.n0) = 0.0


.control
  save v(v_osc)

  * timestep for exact simulation results
  tran 100ps 2us

  remzerovec
  * write tb_pll_bgr_magic.raw
  write tb_pll_bgr_magic_2.raw
  wrdata /foss/designs/my_design/projects/pll/full_pll/magic/tb_pll_bgr_magic_v_osc.txt v(v_osc)
  set appendwrite

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
