magic
tech sky130A
timestamp 1738244200
<< poly >>
rect 6050 -100 8405 -85
rect 6050 -560 6065 -100
rect 6090 -545 6130 -535
rect 6090 -560 6100 -545
rect 6050 -565 6100 -560
rect 6120 -565 6130 -545
rect 8390 -560 8405 -100
rect 6050 -575 6130 -565
rect 8160 -570 8200 -560
rect 8325 -570 8365 -560
rect 8160 -590 8170 -570
rect 8190 -585 8335 -570
rect 8190 -590 8200 -585
rect 8160 -600 8200 -590
rect 8325 -590 8335 -585
rect 8355 -590 8365 -570
rect 8390 -570 8610 -560
rect 8390 -580 8580 -570
rect 8325 -600 8365 -590
rect 8570 -590 8580 -580
rect 8600 -590 8610 -570
rect 8570 -600 8610 -590
rect 8390 -865 8405 -690
rect 8570 -850 8610 -840
rect 8430 -860 8470 -850
rect 8430 -865 8440 -860
rect 8340 -880 8440 -865
rect 8460 -880 8470 -860
rect 8570 -870 8580 -850
rect 8600 -870 8610 -850
rect 8570 -880 8610 -870
rect 8430 -890 8470 -880
<< polycont >>
rect 6100 -565 6120 -545
rect 8170 -590 8190 -570
rect 8335 -590 8355 -570
rect 8580 -590 8600 -570
rect 8440 -880 8460 -860
rect 8580 -870 8600 -850
<< locali >>
rect 8440 -35 9195 -15
rect 6090 -545 6130 -535
rect 6090 -565 6100 -545
rect 6120 -555 6130 -545
rect 6120 -565 6190 -555
rect 6090 -575 6190 -565
rect 8160 -570 8200 -560
rect 6885 -590 8170 -570
rect 8190 -590 8200 -570
rect 8160 -600 8200 -590
rect 8325 -570 8365 -560
rect 8325 -590 8335 -570
rect 8355 -590 8365 -570
rect 8325 -600 8365 -590
rect 8335 -1950 8355 -600
rect 8440 -850 8460 -35
rect 8570 -570 8610 -560
rect 8570 -590 8580 -570
rect 8600 -590 8610 -570
rect 8570 -600 8610 -590
rect 8580 -840 8600 -600
rect 8570 -850 8610 -840
rect 8430 -860 8470 -850
rect 8430 -880 8440 -860
rect 8460 -880 8470 -860
rect 8570 -870 8580 -850
rect 8600 -870 8610 -850
rect 8570 -880 8610 -870
rect 8430 -890 8470 -880
rect 8335 -1970 9470 -1950
<< metal1 >>
rect 6080 -890 6235 -255
rect 8345 -560 8720 -255
rect 8160 -600 8200 -560
rect 8325 -600 8720 -560
rect 8345 -890 8720 -600
rect 6085 -1375 6235 -1020
rect 8345 -1375 8720 -1020
use charge_pump_cell  charge_pump_cell_0
timestamp 1738241744
transform 1 0 -2540 0 1 -2680
box 8630 -35 10885 2425
use opamp_cell  opamp_cell_0
timestamp 1738242334
transform 1 0 4730 0 1 -3070
box 3660 -1 5900 2750
<< labels >>
flabel locali 9195 -25 9195 -25 3 FreeSans 400 0 200 0 VOUT
flabel metal1 6080 -655 6080 -655 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 6085 -1210 6085 -1210 7 FreeSans 400 0 -200 0 GNDA
flabel space 6190 -505 6190 -505 7 FreeSans 400 0 -200 0 x
<< end >>
