magic
tech sky130A
timestamp 1738167417
<< nwell >>
rect -5 190 315 430
<< pwell >>
rect -5 -15 315 95
<< nmos >>
rect 150 -10 165 90
<< pmos >>
rect 150 210 165 410
<< ndiff >>
rect 100 75 150 90
rect 100 5 115 75
rect 135 5 150 75
rect 100 -10 150 5
rect 165 75 215 90
rect 165 5 180 75
rect 200 5 215 75
rect 165 -10 215 5
<< pdiff >>
rect 100 395 150 410
rect 100 225 115 395
rect 135 225 150 395
rect 100 210 150 225
rect 165 395 215 410
rect 165 225 180 395
rect 200 225 215 395
rect 165 210 215 225
<< ndiffc >>
rect 115 5 135 75
rect 180 5 200 75
<< pdiffc >>
rect 115 225 135 395
rect 180 225 200 395
<< psubdiff >>
rect 245 75 295 90
rect 245 5 260 75
rect 280 5 295 75
rect 245 -10 295 5
<< nsubdiff >>
rect 20 395 70 410
rect 20 225 35 395
rect 55 225 70 395
rect 20 210 70 225
<< psubdiffcont >>
rect 260 5 280 75
<< nsubdiffcont >>
rect 35 225 55 395
<< poly >>
rect 150 490 190 500
rect 150 470 160 490
rect 180 470 190 490
rect 150 460 190 470
rect 150 410 165 460
rect 150 195 165 210
rect 105 160 145 170
rect 105 155 115 160
rect 10 140 115 155
rect 135 140 145 160
rect 105 130 145 140
rect 170 160 210 170
rect 170 140 180 160
rect 200 155 210 160
rect 200 140 310 155
rect 170 130 210 140
rect 150 90 165 105
rect 150 -60 165 -10
rect 150 -70 190 -60
rect 150 -90 160 -70
rect 180 -90 190 -70
rect 150 -100 190 -90
<< polycont >>
rect 160 470 180 490
rect 115 140 135 160
rect 180 140 200 160
rect 160 -90 180 -70
<< locali >>
rect -180 500 405 520
rect -180 480 -45 500
rect -25 480 0 500
rect 20 480 150 500
rect 170 490 295 500
rect 180 480 295 490
rect 315 480 350 500
rect 370 480 405 500
rect -180 470 160 480
rect 180 470 405 480
rect -180 460 405 470
rect 25 395 65 405
rect 25 225 35 395
rect 55 225 65 395
rect 25 215 65 225
rect 100 395 145 405
rect 100 225 115 395
rect 135 225 145 395
rect 100 215 145 225
rect 170 395 210 405
rect 170 225 180 395
rect 200 225 210 395
rect 170 215 210 225
rect 35 -60 55 215
rect 115 170 135 215
rect 180 170 200 215
rect 105 160 145 170
rect 105 140 115 160
rect 135 140 145 160
rect 105 130 145 140
rect 170 160 210 170
rect 170 140 180 160
rect 200 140 210 160
rect 170 130 210 140
rect 115 85 135 130
rect 180 85 200 130
rect 260 85 280 460
rect 105 75 145 85
rect 105 5 115 75
rect 135 5 145 75
rect 105 -5 145 5
rect 170 75 210 85
rect 170 5 180 75
rect 200 5 210 75
rect 170 -5 210 5
rect 250 75 290 85
rect 250 5 260 75
rect 280 5 290 75
rect 250 -5 290 5
rect -185 -70 405 -60
rect -185 -80 160 -70
rect 180 -80 405 -70
rect -185 -100 -100 -80
rect -80 -100 -35 -80
rect -15 -100 5 -80
rect 25 -100 150 -80
rect 180 -90 250 -80
rect 170 -100 250 -90
rect 270 -100 295 -80
rect 315 -100 350 -80
rect 370 -100 405 -80
rect -185 -120 405 -100
<< viali >>
rect -45 480 -25 500
rect 0 480 20 500
rect 150 490 170 500
rect 150 480 160 490
rect 160 480 170 490
rect 295 480 315 500
rect 350 480 370 500
rect -100 -100 -80 -80
rect -35 -100 -15 -80
rect 5 -100 25 -80
rect 150 -90 160 -80
rect 160 -90 170 -80
rect 150 -100 170 -90
rect 250 -100 270 -80
rect 295 -100 315 -80
rect 350 -100 370 -80
<< metal1 >>
rect -180 500 405 530
rect -180 480 -45 500
rect -25 480 0 500
rect 20 480 150 500
rect 170 480 295 500
rect 315 480 350 500
rect 370 480 405 500
rect -180 450 405 480
rect -185 -80 405 -50
rect -185 -100 -100 -80
rect -80 -100 -35 -80
rect -15 -100 5 -80
rect 25 -100 150 -80
rect 170 -100 250 -80
rect 270 -100 295 -80
rect 315 -100 350 -80
rect 370 -100 405 -80
rect -185 -130 405 -100
<< labels >>
flabel metal1 -185 -90 -185 -90 7 FreeSans 400 0 -80 0 GNDA
flabel metal1 -180 490 -180 490 7 FreeSans 400 0 -80 0 VDDA
flabel poly 10 150 10 150 7 FreeSans 400 0 -80 0 A
flabel poly 310 150 310 150 3 FreeSans 400 0 80 0 B
<< end >>
