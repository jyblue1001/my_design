magic
tech sky130A
timestamp 1749581722
<< nwell >>
rect 26185 4675 26975 4990
rect 27155 4675 27825 4965
rect 16145 4270 16995 4390
rect 17125 4265 17765 4365
rect 26180 4265 27570 4545
rect 16190 4035 17560 4125
rect 26130 3850 27715 4135
rect 16135 3730 17695 3820
rect 14945 2965 15765 3605
rect 16160 3105 17640 3545
rect 18085 2965 18905 3605
rect 24945 2965 25765 3605
rect 26150 3090 27650 3720
rect 2545 1880 5285 2950
rect 16655 2865 16755 2870
rect 17665 2865 17765 2870
rect 26655 2865 26755 2870
rect 14945 2435 15765 2675
rect 15955 2470 16835 2865
rect 16965 2470 17845 2865
rect 16180 2465 16290 2470
rect 17190 2465 17300 2470
rect 18085 2435 18905 2675
rect 24945 2435 25765 2675
rect 25955 2470 26835 2865
rect 26180 2465 26290 2470
rect 26965 2380 27865 2960
rect 28075 2950 28915 3780
rect 28075 2390 28915 2820
<< pwell >>
rect 29030 3700 29320 3705
rect 29030 3680 29135 3700
rect 29215 3680 29320 3700
rect 29030 2955 29320 3680
rect 15005 1965 15705 2265
rect 16275 1980 17525 2130
rect 18145 1965 18845 2265
rect 25005 1965 25705 2265
rect 26220 1880 27580 2230
rect 28090 1845 28900 2345
rect 28990 1900 29355 2690
rect -45 1685 130 1725
rect 3165 1615 3805 1665
rect 4205 1615 4845 1665
rect 2835 1205 3955 1455
rect 4055 1205 5175 1455
rect 2945 975 5065 1075
rect 15005 955 15645 1655
rect 16030 1515 16730 1665
rect 16770 1515 17030 1665
rect 17070 1515 17770 1665
rect 25935 1660 27865 1825
rect 16205 935 17620 1185
rect 18205 955 18845 1655
rect 25005 955 25645 1655
rect 25935 1520 27770 1660
rect 27775 1520 27865 1660
rect 25935 1355 27865 1520
rect 2995 780 5015 880
rect 16260 650 16530 750
rect 16880 700 17580 750
rect 26135 715 27695 1215
rect 28150 845 28900 1765
rect 28985 825 29230 1720
rect 26200 385 26595 655
rect 26810 400 27640 660
<< nmos >>
rect 15045 1965 15060 2265
rect 15100 1965 15115 2265
rect 15155 1965 15170 2265
rect 15210 1965 15225 2265
rect 15265 1965 15280 2265
rect 15320 1965 15335 2265
rect 15375 1965 15390 2265
rect 15430 1965 15445 2265
rect 15485 1965 15500 2265
rect 15540 1965 15555 2265
rect 15595 1965 15610 2265
rect 15650 1965 15665 2265
rect 16315 1980 16330 2130
rect 16370 1980 16385 2130
rect 16425 1980 16440 2130
rect 16480 1980 16495 2130
rect 16535 1980 16550 2130
rect 16590 1980 16605 2130
rect 16645 1980 16660 2130
rect 16700 1980 16715 2130
rect 16755 1980 16770 2130
rect 16810 1980 16825 2130
rect 16865 1980 16880 2130
rect 16920 1980 16935 2130
rect 16975 1980 16990 2130
rect 17030 1980 17045 2130
rect 17085 1980 17100 2130
rect 17140 1980 17155 2130
rect 17195 1980 17210 2130
rect 17250 1980 17265 2130
rect 17305 1980 17320 2130
rect 17360 1980 17375 2130
rect 17415 1980 17430 2130
rect 17470 1980 17485 2130
rect 18185 1965 18200 2265
rect 18240 1965 18255 2265
rect 18295 1965 18310 2265
rect 18350 1965 18365 2265
rect 18405 1965 18420 2265
rect 18460 1965 18475 2265
rect 18515 1965 18530 2265
rect 18570 1965 18585 2265
rect 18625 1965 18640 2265
rect 18680 1965 18695 2265
rect 18735 1965 18750 2265
rect 18790 1965 18805 2265
rect 25045 1965 25060 2265
rect 25100 1965 25115 2265
rect 25155 1965 25170 2265
rect 25210 1965 25225 2265
rect 25265 1965 25280 2265
rect 25320 1965 25335 2265
rect 25375 1965 25390 2265
rect 25430 1965 25445 2265
rect 25485 1965 25500 2265
rect 25540 1965 25555 2265
rect 25595 1965 25610 2265
rect 25650 1965 25665 2265
rect 26315 1980 26330 2130
rect 26370 1980 26385 2130
rect 26425 1980 26440 2130
rect 26480 1980 26495 2130
rect 26535 1980 26550 2130
rect 26590 1980 26605 2130
rect 26645 1980 26660 2130
rect 26700 1980 26715 2130
rect 26755 1980 26770 2130
rect 26810 1980 26825 2130
rect 26865 1980 26880 2130
rect 26920 1980 26935 2130
rect 26975 1980 26990 2130
rect 27030 1980 27045 2130
rect 27085 1980 27100 2130
rect 27140 1980 27155 2130
rect 27195 1980 27210 2130
rect 27250 1980 27265 2130
rect 27305 1980 27320 2130
rect 27360 1980 27375 2130
rect 27415 1980 27430 2130
rect 27470 1980 27485 2130
rect 28185 1945 28200 2245
rect 28240 1945 28255 2245
rect 28295 1945 28310 2245
rect 28350 1945 28365 2245
rect 28405 1945 28420 2245
rect 28460 1945 28475 2245
rect 28515 1945 28530 2245
rect 28570 1945 28585 2245
rect 28625 1945 28640 2245
rect 28680 1945 28695 2245
rect 28735 1945 28750 2245
rect 28790 1945 28805 2245
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 4785 1615 4805 1665
rect 2875 1205 3375 1455
rect 3415 1205 3915 1455
rect 4095 1205 4595 1455
rect 4635 1205 5135 1455
rect 2985 975 3985 1075
rect 4025 975 5025 1075
rect 15045 955 15105 1655
rect 15145 955 15205 1655
rect 15245 955 15305 1655
rect 15345 955 15405 1655
rect 15445 955 15505 1655
rect 15545 955 15605 1655
rect 16070 1515 16085 1665
rect 16125 1515 16140 1665
rect 16180 1515 16195 1665
rect 16235 1515 16250 1665
rect 16290 1515 16305 1665
rect 16345 1515 16360 1665
rect 16400 1515 16415 1665
rect 16455 1515 16470 1665
rect 16510 1515 16525 1665
rect 16565 1515 16580 1665
rect 16620 1515 16635 1665
rect 16675 1515 16690 1665
rect 16810 1515 16825 1665
rect 16865 1515 16880 1665
rect 16920 1515 16935 1665
rect 16975 1515 16990 1665
rect 17110 1515 17125 1665
rect 17165 1515 17180 1665
rect 17220 1515 17235 1665
rect 17275 1515 17290 1665
rect 17330 1515 17345 1665
rect 17385 1515 17400 1665
rect 17440 1515 17455 1665
rect 17495 1515 17510 1665
rect 17550 1515 17565 1665
rect 17605 1515 17620 1665
rect 17660 1515 17675 1665
rect 17715 1515 17730 1665
rect 16245 935 16260 1185
rect 16300 935 16315 1185
rect 16355 935 16370 1185
rect 16410 935 16425 1185
rect 16465 935 16480 1185
rect 16520 935 16535 1185
rect 16575 935 16590 1185
rect 16630 935 16645 1185
rect 16685 935 16700 1185
rect 16740 935 16755 1185
rect 16795 935 16810 1185
rect 16850 935 16865 1185
rect 16905 935 16920 1185
rect 16960 935 16975 1185
rect 17015 935 17030 1185
rect 17070 935 17085 1185
rect 17125 935 17140 1185
rect 17180 935 17195 1185
rect 17235 935 17250 1185
rect 17290 935 17305 1185
rect 17345 935 17360 1185
rect 17400 935 17415 1185
rect 17455 935 17470 1185
rect 17510 935 17525 1185
rect 17565 935 17580 1185
rect 18245 955 18305 1655
rect 18345 955 18405 1655
rect 18445 955 18505 1655
rect 18545 955 18605 1655
rect 18645 955 18705 1655
rect 18745 955 18805 1655
rect 25045 955 25105 1655
rect 25145 955 25205 1655
rect 25245 955 25305 1655
rect 25345 955 25405 1655
rect 25445 955 25505 1655
rect 25545 955 25605 1655
rect 26070 1515 26085 1665
rect 26125 1515 26140 1665
rect 26180 1515 26195 1665
rect 26235 1515 26250 1665
rect 26290 1515 26305 1665
rect 26345 1515 26360 1665
rect 26400 1515 26415 1665
rect 26455 1515 26470 1665
rect 26510 1515 26525 1665
rect 26565 1515 26580 1665
rect 26620 1515 26635 1665
rect 26675 1515 26690 1665
rect 26810 1515 26825 1665
rect 26865 1515 26880 1665
rect 26920 1515 26935 1665
rect 26975 1515 26990 1665
rect 27110 1515 27125 1665
rect 27165 1515 27180 1665
rect 27220 1515 27235 1665
rect 27275 1515 27290 1665
rect 27330 1515 27345 1665
rect 27385 1515 27400 1665
rect 27440 1515 27455 1665
rect 27495 1515 27510 1665
rect 27550 1515 27565 1665
rect 27605 1515 27620 1665
rect 27660 1515 27675 1665
rect 27715 1515 27730 1665
rect 3035 780 3085 880
rect 3125 780 3175 880
rect 3215 780 3265 880
rect 3305 780 3355 880
rect 3395 780 3445 880
rect 3485 780 3535 880
rect 3575 780 3625 880
rect 3665 780 3715 880
rect 3755 780 3805 880
rect 3845 780 3895 880
rect 3935 780 3985 880
rect 4025 780 4075 880
rect 4115 780 4165 880
rect 4205 780 4255 880
rect 4295 780 4345 880
rect 4385 780 4435 880
rect 4475 780 4525 880
rect 4565 780 4615 880
rect 4655 780 4705 880
rect 4745 780 4795 880
rect 4835 780 4885 880
rect 4925 780 4975 880
rect 26245 835 26260 1085
rect 26300 835 26315 1085
rect 26355 835 26370 1085
rect 26410 835 26425 1085
rect 26465 835 26480 1085
rect 26520 835 26535 1085
rect 26575 835 26590 1085
rect 26630 835 26645 1085
rect 26685 835 26700 1085
rect 26740 835 26755 1085
rect 26795 835 26810 1085
rect 26850 835 26865 1085
rect 26905 835 26920 1085
rect 26960 835 26975 1085
rect 27015 835 27030 1085
rect 27070 835 27085 1085
rect 27125 835 27140 1085
rect 27180 835 27195 1085
rect 27235 835 27250 1085
rect 27290 835 27305 1085
rect 27345 835 27360 1085
rect 27400 835 27415 1085
rect 27455 835 27470 1085
rect 27510 835 27525 1085
rect 27565 835 27580 1085
rect 28245 955 28305 1655
rect 28345 955 28405 1655
rect 28445 955 28505 1655
rect 28545 955 28605 1655
rect 28645 955 28705 1655
rect 28745 955 28805 1655
rect 16300 650 16490 750
rect 16920 700 16935 750
rect 16975 700 16990 750
rect 17030 700 17045 750
rect 17085 700 17100 750
rect 17140 700 17155 750
rect 17195 700 17210 750
rect 17250 700 17265 750
rect 17305 700 17320 750
rect 17360 700 17375 750
rect 17415 700 17430 750
rect 17470 700 17485 750
rect 17525 700 17540 750
rect 26300 450 26490 550
rect 26920 500 26935 550
rect 26975 500 26990 550
rect 27030 500 27045 550
rect 27085 500 27100 550
rect 27140 500 27155 550
rect 27195 500 27210 550
rect 27250 500 27265 550
rect 27305 500 27320 550
rect 27360 500 27375 550
rect 27415 500 27430 550
rect 27470 500 27485 550
rect 27525 500 27540 550
<< pmos >>
rect 26295 4795 26315 4858
rect 26355 4795 26375 4858
rect 26415 4795 26435 4858
rect 26545 4795 26565 4875
rect 26605 4795 26625 4875
rect 26665 4795 26685 4875
rect 26725 4795 26745 4875
rect 26785 4795 26805 4875
rect 26845 4795 26865 4875
rect 27275 4790 27295 4850
rect 27335 4790 27355 4850
rect 27395 4790 27415 4850
rect 27455 4790 27475 4850
rect 27515 4790 27535 4850
rect 27575 4790 27595 4850
rect 27635 4790 27655 4850
rect 27695 4790 27715 4850
rect 16245 4290 16265 4353
rect 16305 4290 16325 4353
rect 16365 4290 16385 4353
rect 16575 4290 16595 4370
rect 16635 4290 16655 4370
rect 16695 4290 16715 4370
rect 16755 4290 16775 4370
rect 16815 4290 16835 4370
rect 16875 4290 16895 4370
rect 26290 4380 26305 4430
rect 26345 4380 26360 4430
rect 26400 4380 26415 4430
rect 26455 4380 26470 4430
rect 26510 4380 26525 4430
rect 26565 4380 26580 4430
rect 26620 4380 26635 4430
rect 26675 4380 26690 4430
rect 26730 4380 26745 4430
rect 26785 4380 26800 4430
rect 26840 4380 26855 4430
rect 26895 4380 26910 4430
rect 26950 4380 26965 4430
rect 27005 4380 27020 4430
rect 27060 4380 27075 4430
rect 27115 4380 27130 4430
rect 27170 4380 27185 4430
rect 27225 4380 27240 4430
rect 27280 4380 27295 4430
rect 27335 4380 27350 4430
rect 27390 4380 27405 4430
rect 27445 4380 27460 4430
rect 17225 4285 17245 4345
rect 17285 4285 17305 4345
rect 17345 4285 17365 4345
rect 17405 4285 17425 4345
rect 17465 4285 17485 4345
rect 17525 4285 17545 4345
rect 17585 4285 17605 4345
rect 17645 4285 17665 4345
rect 16290 4055 16305 4105
rect 16345 4055 16360 4105
rect 16400 4055 16415 4105
rect 16455 4055 16470 4105
rect 16510 4055 16525 4105
rect 16565 4055 16580 4105
rect 16620 4055 16635 4105
rect 16675 4055 16690 4105
rect 16730 4055 16745 4105
rect 16785 4055 16800 4105
rect 16840 4055 16855 4105
rect 16895 4055 16910 4105
rect 16950 4055 16965 4105
rect 17005 4055 17020 4105
rect 17060 4055 17075 4105
rect 17115 4055 17130 4105
rect 17170 4055 17185 4105
rect 17225 4055 17240 4105
rect 17280 4055 17295 4105
rect 17335 4055 17350 4105
rect 17390 4055 17405 4105
rect 17445 4055 17460 4105
rect 26240 3970 26255 4020
rect 26295 3970 26310 4020
rect 26350 3970 26365 4020
rect 26405 3970 26420 4020
rect 26460 3970 26475 4020
rect 26515 3970 26530 4020
rect 26570 3970 26585 4020
rect 26625 3970 26640 4020
rect 26680 3970 26695 4020
rect 26735 3970 26750 4020
rect 26790 3970 26805 4020
rect 26845 3970 26860 4020
rect 26970 3970 26985 4020
rect 27025 3970 27040 4020
rect 27080 3970 27095 4020
rect 27135 3970 27150 4020
rect 27190 3970 27205 4020
rect 27245 3970 27260 4020
rect 27300 3970 27315 4020
rect 27355 3970 27370 4020
rect 27410 3970 27425 4020
rect 27465 3970 27480 4020
rect 27520 3970 27535 4020
rect 27575 3970 27590 4020
rect 16235 3750 16250 3800
rect 16290 3750 16305 3800
rect 16345 3750 16360 3800
rect 16400 3750 16415 3800
rect 16455 3750 16470 3800
rect 16510 3750 16525 3800
rect 16565 3750 16580 3800
rect 16620 3750 16635 3800
rect 16675 3750 16690 3800
rect 16730 3750 16745 3800
rect 16785 3750 16800 3800
rect 16840 3750 16855 3800
rect 16975 3750 16990 3800
rect 17030 3750 17045 3800
rect 17085 3750 17100 3800
rect 17140 3750 17155 3800
rect 17195 3750 17210 3800
rect 17250 3750 17265 3800
rect 17305 3750 17320 3800
rect 17360 3750 17375 3800
rect 17415 3750 17430 3800
rect 17470 3750 17485 3800
rect 17525 3750 17540 3800
rect 17580 3750 17595 3800
rect 15045 2985 15060 3585
rect 15100 2985 15115 3585
rect 15155 2985 15170 3585
rect 15210 2985 15225 3585
rect 15265 2985 15280 3585
rect 15320 2985 15335 3585
rect 15375 2985 15390 3585
rect 15430 2985 15445 3585
rect 15485 2985 15500 3585
rect 15540 2985 15555 3585
rect 15595 2985 15610 3585
rect 15650 2985 15665 3585
rect 16260 3125 16280 3525
rect 16320 3125 16340 3525
rect 16380 3125 16400 3525
rect 16440 3125 16460 3525
rect 16500 3125 16520 3525
rect 16560 3125 16580 3525
rect 16620 3125 16640 3525
rect 16680 3125 16700 3525
rect 16740 3125 16760 3525
rect 16800 3125 16820 3525
rect 16860 3125 16880 3525
rect 16920 3125 16940 3525
rect 16980 3125 17000 3525
rect 17040 3125 17060 3525
rect 17100 3125 17120 3525
rect 17160 3125 17180 3525
rect 17220 3125 17240 3525
rect 17280 3125 17300 3525
rect 17340 3125 17360 3525
rect 17400 3125 17420 3525
rect 17460 3125 17480 3525
rect 17520 3125 17540 3525
rect 18185 2985 18200 3585
rect 18240 2985 18255 3585
rect 18295 2985 18310 3585
rect 18350 2985 18365 3585
rect 18405 2985 18420 3585
rect 18460 2985 18475 3585
rect 18515 2985 18530 3585
rect 18570 2985 18585 3585
rect 18625 2985 18640 3585
rect 18680 2985 18695 3585
rect 18735 2985 18750 3585
rect 18790 2985 18805 3585
rect 25045 2985 25060 3585
rect 25100 2985 25115 3585
rect 25155 2985 25170 3585
rect 25210 2985 25225 3585
rect 25265 2985 25280 3585
rect 25320 2985 25335 3585
rect 25375 2985 25390 3585
rect 25430 2985 25445 3585
rect 25485 2985 25500 3585
rect 25540 2985 25555 3585
rect 25595 2985 25610 3585
rect 25650 2985 25665 3585
rect 26260 3205 26280 3605
rect 26320 3205 26340 3605
rect 26380 3205 26400 3605
rect 26440 3205 26460 3605
rect 26500 3205 26520 3605
rect 26560 3205 26580 3605
rect 26620 3205 26640 3605
rect 26680 3205 26700 3605
rect 26740 3205 26760 3605
rect 26800 3205 26820 3605
rect 26860 3205 26880 3605
rect 26920 3205 26940 3605
rect 26980 3205 27000 3605
rect 27040 3205 27060 3605
rect 27100 3205 27120 3605
rect 27160 3205 27180 3605
rect 27220 3205 27240 3605
rect 27280 3205 27300 3605
rect 27340 3205 27360 3605
rect 27400 3205 27420 3605
rect 27460 3205 27480 3605
rect 27520 3205 27540 3605
rect 28185 3065 28200 3665
rect 28240 3065 28255 3665
rect 28295 3065 28310 3665
rect 28350 3065 28365 3665
rect 28405 3065 28420 3665
rect 28460 3065 28475 3665
rect 28515 3065 28530 3665
rect 28570 3065 28585 3665
rect 28625 3065 28640 3665
rect 28680 3065 28695 3665
rect 28735 3065 28750 3665
rect 28790 3065 28805 3665
rect 3035 2830 3085 2930
rect 3125 2830 3175 2930
rect 3215 2830 3265 2930
rect 3305 2830 3355 2930
rect 3395 2830 3445 2930
rect 3485 2830 3535 2930
rect 3575 2830 3625 2930
rect 3665 2830 3715 2930
rect 3755 2830 3805 2930
rect 3845 2830 3895 2930
rect 3935 2830 3985 2930
rect 4025 2830 4075 2930
rect 4115 2830 4165 2930
rect 4205 2830 4255 2930
rect 4295 2830 4345 2930
rect 4385 2830 4435 2930
rect 4475 2830 4525 2930
rect 4565 2830 4615 2930
rect 4655 2830 4705 2930
rect 4745 2830 4795 2930
rect 4835 2830 4885 2930
rect 4925 2830 4975 2930
rect 3215 2400 3265 2700
rect 3305 2400 3355 2700
rect 3395 2400 3445 2700
rect 3485 2400 3535 2700
rect 3575 2400 3625 2700
rect 3665 2400 3715 2700
rect 3755 2400 3805 2700
rect 3845 2400 3895 2700
rect 3935 2400 3985 2700
rect 4025 2400 4075 2700
rect 4115 2400 4165 2700
rect 4205 2400 4255 2700
rect 4295 2400 4345 2700
rect 4385 2400 4435 2700
rect 4475 2400 4525 2700
rect 4565 2400 4615 2700
rect 4655 2400 4705 2700
rect 4745 2400 4795 2700
rect 15045 2455 15060 2655
rect 15100 2455 15115 2655
rect 15155 2455 15170 2655
rect 15210 2455 15225 2655
rect 15265 2455 15280 2655
rect 15320 2455 15335 2655
rect 15375 2455 15390 2655
rect 15430 2455 15445 2655
rect 15485 2455 15500 2655
rect 15540 2455 15555 2655
rect 15595 2455 15610 2655
rect 15650 2455 15665 2655
rect 16055 2495 16075 2845
rect 16115 2495 16135 2845
rect 16175 2495 16195 2845
rect 16235 2495 16255 2845
rect 16295 2495 16315 2845
rect 16355 2495 16375 2845
rect 16415 2495 16435 2845
rect 16475 2495 16495 2845
rect 16535 2495 16555 2845
rect 16595 2495 16615 2845
rect 16655 2495 16675 2845
rect 16715 2495 16735 2845
rect 17065 2495 17085 2845
rect 17125 2495 17145 2845
rect 17185 2495 17205 2845
rect 17245 2495 17265 2845
rect 17305 2495 17325 2845
rect 17365 2495 17385 2845
rect 17425 2495 17445 2845
rect 17485 2495 17505 2845
rect 17545 2495 17565 2845
rect 17605 2495 17625 2845
rect 17665 2495 17685 2845
rect 17725 2495 17745 2845
rect 18185 2455 18200 2655
rect 18240 2455 18255 2655
rect 18295 2455 18310 2655
rect 18350 2455 18365 2655
rect 18405 2455 18420 2655
rect 18460 2455 18475 2655
rect 18515 2455 18530 2655
rect 18570 2455 18585 2655
rect 18625 2455 18640 2655
rect 18680 2455 18695 2655
rect 18735 2455 18750 2655
rect 18790 2455 18805 2655
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 5205 1900 5225 2000
rect 25045 2455 25060 2655
rect 25100 2455 25115 2655
rect 25155 2455 25170 2655
rect 25210 2455 25225 2655
rect 25265 2455 25280 2655
rect 25320 2455 25335 2655
rect 25375 2455 25390 2655
rect 25430 2455 25445 2655
rect 25485 2455 25500 2655
rect 25540 2455 25555 2655
rect 25595 2455 25610 2655
rect 25650 2455 25665 2655
rect 26055 2495 26075 2845
rect 26115 2495 26135 2845
rect 26175 2495 26195 2845
rect 26235 2495 26255 2845
rect 26295 2495 26315 2845
rect 26355 2495 26375 2845
rect 26415 2495 26435 2845
rect 26475 2495 26495 2845
rect 26535 2495 26555 2845
rect 26595 2495 26615 2845
rect 26655 2495 26675 2845
rect 26715 2495 26735 2845
rect 27075 2495 27095 2845
rect 27135 2495 27155 2845
rect 27195 2495 27215 2845
rect 27255 2495 27275 2845
rect 27315 2495 27335 2845
rect 27375 2495 27395 2845
rect 27435 2495 27455 2845
rect 27495 2495 27515 2845
rect 27555 2495 27575 2845
rect 27615 2495 27635 2845
rect 27675 2495 27695 2845
rect 27735 2495 27755 2845
rect 28185 2505 28200 2705
rect 28240 2505 28255 2705
rect 28295 2505 28310 2705
rect 28350 2505 28365 2705
rect 28405 2505 28420 2705
rect 28460 2505 28475 2705
rect 28515 2505 28530 2705
rect 28570 2505 28585 2705
rect 28625 2505 28640 2705
rect 28680 2505 28695 2705
rect 28735 2505 28750 2705
rect 28790 2505 28805 2705
<< ndiff >>
rect 15005 2250 15045 2265
rect 15005 2230 15015 2250
rect 15035 2230 15045 2250
rect 15005 2200 15045 2230
rect 15005 2180 15015 2200
rect 15035 2180 15045 2200
rect 15005 2150 15045 2180
rect 15005 2130 15015 2150
rect 15035 2130 15045 2150
rect 15005 2100 15045 2130
rect 15005 2080 15015 2100
rect 15035 2080 15045 2100
rect 15005 2050 15045 2080
rect 15005 2030 15015 2050
rect 15035 2030 15045 2050
rect 15005 2000 15045 2030
rect 15005 1980 15015 2000
rect 15035 1980 15045 2000
rect 15005 1965 15045 1980
rect 15060 2250 15100 2265
rect 15060 2230 15070 2250
rect 15090 2230 15100 2250
rect 15060 2200 15100 2230
rect 15060 2180 15070 2200
rect 15090 2180 15100 2200
rect 15060 2150 15100 2180
rect 15060 2130 15070 2150
rect 15090 2130 15100 2150
rect 15060 2100 15100 2130
rect 15060 2080 15070 2100
rect 15090 2080 15100 2100
rect 15060 2050 15100 2080
rect 15060 2030 15070 2050
rect 15090 2030 15100 2050
rect 15060 2000 15100 2030
rect 15060 1980 15070 2000
rect 15090 1980 15100 2000
rect 15060 1965 15100 1980
rect 15115 2250 15155 2265
rect 15115 2230 15125 2250
rect 15145 2230 15155 2250
rect 15115 2200 15155 2230
rect 15115 2180 15125 2200
rect 15145 2180 15155 2200
rect 15115 2150 15155 2180
rect 15115 2130 15125 2150
rect 15145 2130 15155 2150
rect 15115 2100 15155 2130
rect 15115 2080 15125 2100
rect 15145 2080 15155 2100
rect 15115 2050 15155 2080
rect 15115 2030 15125 2050
rect 15145 2030 15155 2050
rect 15115 2000 15155 2030
rect 15115 1980 15125 2000
rect 15145 1980 15155 2000
rect 15115 1965 15155 1980
rect 15170 2250 15210 2265
rect 15170 2230 15180 2250
rect 15200 2230 15210 2250
rect 15170 2200 15210 2230
rect 15170 2180 15180 2200
rect 15200 2180 15210 2200
rect 15170 2150 15210 2180
rect 15170 2130 15180 2150
rect 15200 2130 15210 2150
rect 15170 2100 15210 2130
rect 15170 2080 15180 2100
rect 15200 2080 15210 2100
rect 15170 2050 15210 2080
rect 15170 2030 15180 2050
rect 15200 2030 15210 2050
rect 15170 2000 15210 2030
rect 15170 1980 15180 2000
rect 15200 1980 15210 2000
rect 15170 1965 15210 1980
rect 15225 2250 15265 2265
rect 15225 2230 15235 2250
rect 15255 2230 15265 2250
rect 15225 2200 15265 2230
rect 15225 2180 15235 2200
rect 15255 2180 15265 2200
rect 15225 2150 15265 2180
rect 15225 2130 15235 2150
rect 15255 2130 15265 2150
rect 15225 2100 15265 2130
rect 15225 2080 15235 2100
rect 15255 2080 15265 2100
rect 15225 2050 15265 2080
rect 15225 2030 15235 2050
rect 15255 2030 15265 2050
rect 15225 2000 15265 2030
rect 15225 1980 15235 2000
rect 15255 1980 15265 2000
rect 15225 1965 15265 1980
rect 15280 2250 15320 2265
rect 15280 2230 15290 2250
rect 15310 2230 15320 2250
rect 15280 2200 15320 2230
rect 15280 2180 15290 2200
rect 15310 2180 15320 2200
rect 15280 2150 15320 2180
rect 15280 2130 15290 2150
rect 15310 2130 15320 2150
rect 15280 2100 15320 2130
rect 15280 2080 15290 2100
rect 15310 2080 15320 2100
rect 15280 2050 15320 2080
rect 15280 2030 15290 2050
rect 15310 2030 15320 2050
rect 15280 2000 15320 2030
rect 15280 1980 15290 2000
rect 15310 1980 15320 2000
rect 15280 1965 15320 1980
rect 15335 2250 15375 2265
rect 15335 2230 15345 2250
rect 15365 2230 15375 2250
rect 15335 2200 15375 2230
rect 15335 2180 15345 2200
rect 15365 2180 15375 2200
rect 15335 2150 15375 2180
rect 15335 2130 15345 2150
rect 15365 2130 15375 2150
rect 15335 2100 15375 2130
rect 15335 2080 15345 2100
rect 15365 2080 15375 2100
rect 15335 2050 15375 2080
rect 15335 2030 15345 2050
rect 15365 2030 15375 2050
rect 15335 2000 15375 2030
rect 15335 1980 15345 2000
rect 15365 1980 15375 2000
rect 15335 1965 15375 1980
rect 15390 2250 15430 2265
rect 15390 2230 15400 2250
rect 15420 2230 15430 2250
rect 15390 2200 15430 2230
rect 15390 2180 15400 2200
rect 15420 2180 15430 2200
rect 15390 2150 15430 2180
rect 15390 2130 15400 2150
rect 15420 2130 15430 2150
rect 15390 2100 15430 2130
rect 15390 2080 15400 2100
rect 15420 2080 15430 2100
rect 15390 2050 15430 2080
rect 15390 2030 15400 2050
rect 15420 2030 15430 2050
rect 15390 2000 15430 2030
rect 15390 1980 15400 2000
rect 15420 1980 15430 2000
rect 15390 1965 15430 1980
rect 15445 2250 15485 2265
rect 15445 2230 15455 2250
rect 15475 2230 15485 2250
rect 15445 2200 15485 2230
rect 15445 2180 15455 2200
rect 15475 2180 15485 2200
rect 15445 2150 15485 2180
rect 15445 2130 15455 2150
rect 15475 2130 15485 2150
rect 15445 2100 15485 2130
rect 15445 2080 15455 2100
rect 15475 2080 15485 2100
rect 15445 2050 15485 2080
rect 15445 2030 15455 2050
rect 15475 2030 15485 2050
rect 15445 2000 15485 2030
rect 15445 1980 15455 2000
rect 15475 1980 15485 2000
rect 15445 1965 15485 1980
rect 15500 2250 15540 2265
rect 15500 2230 15510 2250
rect 15530 2230 15540 2250
rect 15500 2200 15540 2230
rect 15500 2180 15510 2200
rect 15530 2180 15540 2200
rect 15500 2150 15540 2180
rect 15500 2130 15510 2150
rect 15530 2130 15540 2150
rect 15500 2100 15540 2130
rect 15500 2080 15510 2100
rect 15530 2080 15540 2100
rect 15500 2050 15540 2080
rect 15500 2030 15510 2050
rect 15530 2030 15540 2050
rect 15500 2000 15540 2030
rect 15500 1980 15510 2000
rect 15530 1980 15540 2000
rect 15500 1965 15540 1980
rect 15555 2250 15595 2265
rect 15555 2230 15565 2250
rect 15585 2230 15595 2250
rect 15555 2200 15595 2230
rect 15555 2180 15565 2200
rect 15585 2180 15595 2200
rect 15555 2150 15595 2180
rect 15555 2130 15565 2150
rect 15585 2130 15595 2150
rect 15555 2100 15595 2130
rect 15555 2080 15565 2100
rect 15585 2080 15595 2100
rect 15555 2050 15595 2080
rect 15555 2030 15565 2050
rect 15585 2030 15595 2050
rect 15555 2000 15595 2030
rect 15555 1980 15565 2000
rect 15585 1980 15595 2000
rect 15555 1965 15595 1980
rect 15610 2250 15650 2265
rect 15610 2230 15620 2250
rect 15640 2230 15650 2250
rect 15610 2200 15650 2230
rect 15610 2180 15620 2200
rect 15640 2180 15650 2200
rect 15610 2150 15650 2180
rect 15610 2130 15620 2150
rect 15640 2130 15650 2150
rect 15610 2100 15650 2130
rect 15610 2080 15620 2100
rect 15640 2080 15650 2100
rect 15610 2050 15650 2080
rect 15610 2030 15620 2050
rect 15640 2030 15650 2050
rect 15610 2000 15650 2030
rect 15610 1980 15620 2000
rect 15640 1980 15650 2000
rect 15610 1965 15650 1980
rect 15665 2250 15705 2265
rect 15665 2230 15675 2250
rect 15695 2230 15705 2250
rect 15665 2200 15705 2230
rect 15665 2180 15675 2200
rect 15695 2180 15705 2200
rect 18145 2250 18185 2265
rect 18145 2230 18155 2250
rect 18175 2230 18185 2250
rect 18145 2200 18185 2230
rect 15665 2150 15705 2180
rect 18145 2180 18155 2200
rect 18175 2180 18185 2200
rect 15665 2130 15675 2150
rect 15695 2130 15705 2150
rect 18145 2150 18185 2180
rect 18145 2130 18155 2150
rect 18175 2130 18185 2150
rect 15665 2100 15705 2130
rect 15665 2080 15675 2100
rect 15695 2080 15705 2100
rect 15665 2050 15705 2080
rect 15665 2030 15675 2050
rect 15695 2030 15705 2050
rect 15665 2000 15705 2030
rect 15665 1980 15675 2000
rect 15695 1980 15705 2000
rect 16275 2115 16315 2130
rect 16275 2095 16285 2115
rect 16305 2095 16315 2115
rect 16275 2065 16315 2095
rect 16275 2045 16285 2065
rect 16305 2045 16315 2065
rect 16275 2015 16315 2045
rect 16275 1995 16285 2015
rect 16305 1995 16315 2015
rect 16275 1980 16315 1995
rect 16330 2115 16370 2130
rect 16330 2095 16340 2115
rect 16360 2095 16370 2115
rect 16330 2065 16370 2095
rect 16330 2045 16340 2065
rect 16360 2045 16370 2065
rect 16330 2015 16370 2045
rect 16330 1995 16340 2015
rect 16360 1995 16370 2015
rect 16330 1980 16370 1995
rect 16385 2115 16425 2130
rect 16385 2095 16395 2115
rect 16415 2095 16425 2115
rect 16385 2065 16425 2095
rect 16385 2045 16395 2065
rect 16415 2045 16425 2065
rect 16385 2015 16425 2045
rect 16385 1995 16395 2015
rect 16415 1995 16425 2015
rect 16385 1980 16425 1995
rect 16440 2115 16480 2130
rect 16440 2095 16450 2115
rect 16470 2095 16480 2115
rect 16440 2065 16480 2095
rect 16440 2045 16450 2065
rect 16470 2045 16480 2065
rect 16440 2015 16480 2045
rect 16440 1995 16450 2015
rect 16470 1995 16480 2015
rect 16440 1980 16480 1995
rect 16495 2115 16535 2130
rect 16495 2095 16505 2115
rect 16525 2095 16535 2115
rect 16495 2065 16535 2095
rect 16495 2045 16505 2065
rect 16525 2045 16535 2065
rect 16495 2015 16535 2045
rect 16495 1995 16505 2015
rect 16525 1995 16535 2015
rect 16495 1980 16535 1995
rect 16550 2115 16590 2130
rect 16550 2095 16560 2115
rect 16580 2095 16590 2115
rect 16550 2065 16590 2095
rect 16550 2045 16560 2065
rect 16580 2045 16590 2065
rect 16550 2015 16590 2045
rect 16550 1995 16560 2015
rect 16580 1995 16590 2015
rect 16550 1980 16590 1995
rect 16605 2115 16645 2130
rect 16605 2095 16615 2115
rect 16635 2095 16645 2115
rect 16605 2065 16645 2095
rect 16605 2045 16615 2065
rect 16635 2045 16645 2065
rect 16605 2015 16645 2045
rect 16605 1995 16615 2015
rect 16635 1995 16645 2015
rect 16605 1980 16645 1995
rect 16660 2115 16700 2130
rect 16660 2095 16670 2115
rect 16690 2095 16700 2115
rect 16660 2065 16700 2095
rect 16660 2045 16670 2065
rect 16690 2045 16700 2065
rect 16660 2015 16700 2045
rect 16660 1995 16670 2015
rect 16690 1995 16700 2015
rect 16660 1980 16700 1995
rect 16715 2115 16755 2130
rect 16715 2095 16725 2115
rect 16745 2095 16755 2115
rect 16715 2065 16755 2095
rect 16715 2045 16725 2065
rect 16745 2045 16755 2065
rect 16715 2015 16755 2045
rect 16715 1995 16725 2015
rect 16745 1995 16755 2015
rect 16715 1980 16755 1995
rect 16770 2115 16810 2130
rect 16770 2095 16780 2115
rect 16800 2095 16810 2115
rect 16770 2065 16810 2095
rect 16770 2045 16780 2065
rect 16800 2045 16810 2065
rect 16770 2015 16810 2045
rect 16770 1995 16780 2015
rect 16800 1995 16810 2015
rect 16770 1980 16810 1995
rect 16825 2115 16865 2130
rect 16825 2095 16835 2115
rect 16855 2095 16865 2115
rect 16825 2065 16865 2095
rect 16825 2045 16835 2065
rect 16855 2045 16865 2065
rect 16825 2015 16865 2045
rect 16825 1995 16835 2015
rect 16855 1995 16865 2015
rect 16825 1980 16865 1995
rect 16880 2115 16920 2130
rect 16880 2095 16890 2115
rect 16910 2095 16920 2115
rect 16880 2065 16920 2095
rect 16880 2045 16890 2065
rect 16910 2045 16920 2065
rect 16880 2015 16920 2045
rect 16880 1995 16890 2015
rect 16910 1995 16920 2015
rect 16880 1980 16920 1995
rect 16935 2115 16975 2130
rect 16935 2095 16945 2115
rect 16965 2095 16975 2115
rect 16935 2065 16975 2095
rect 16935 2045 16945 2065
rect 16965 2045 16975 2065
rect 16935 2015 16975 2045
rect 16935 1995 16945 2015
rect 16965 1995 16975 2015
rect 16935 1980 16975 1995
rect 16990 2115 17030 2130
rect 16990 2095 17000 2115
rect 17020 2095 17030 2115
rect 16990 2065 17030 2095
rect 16990 2045 17000 2065
rect 17020 2045 17030 2065
rect 16990 2015 17030 2045
rect 16990 1995 17000 2015
rect 17020 1995 17030 2015
rect 16990 1980 17030 1995
rect 17045 2115 17085 2130
rect 17045 2095 17055 2115
rect 17075 2095 17085 2115
rect 17045 2065 17085 2095
rect 17045 2045 17055 2065
rect 17075 2045 17085 2065
rect 17045 2015 17085 2045
rect 17045 1995 17055 2015
rect 17075 1995 17085 2015
rect 17045 1980 17085 1995
rect 17100 2115 17140 2130
rect 17100 2095 17110 2115
rect 17130 2095 17140 2115
rect 17100 2065 17140 2095
rect 17100 2045 17110 2065
rect 17130 2045 17140 2065
rect 17100 2015 17140 2045
rect 17100 1995 17110 2015
rect 17130 1995 17140 2015
rect 17100 1980 17140 1995
rect 17155 2115 17195 2130
rect 17155 2095 17165 2115
rect 17185 2095 17195 2115
rect 17155 2065 17195 2095
rect 17155 2045 17165 2065
rect 17185 2045 17195 2065
rect 17155 2015 17195 2045
rect 17155 1995 17165 2015
rect 17185 1995 17195 2015
rect 17155 1980 17195 1995
rect 17210 2115 17250 2130
rect 17210 2095 17220 2115
rect 17240 2095 17250 2115
rect 17210 2065 17250 2095
rect 17210 2045 17220 2065
rect 17240 2045 17250 2065
rect 17210 2015 17250 2045
rect 17210 1995 17220 2015
rect 17240 1995 17250 2015
rect 17210 1980 17250 1995
rect 17265 2115 17305 2130
rect 17265 2095 17275 2115
rect 17295 2095 17305 2115
rect 17265 2065 17305 2095
rect 17265 2045 17275 2065
rect 17295 2045 17305 2065
rect 17265 2015 17305 2045
rect 17265 1995 17275 2015
rect 17295 1995 17305 2015
rect 17265 1980 17305 1995
rect 17320 2115 17360 2130
rect 17320 2095 17330 2115
rect 17350 2095 17360 2115
rect 17320 2065 17360 2095
rect 17320 2045 17330 2065
rect 17350 2045 17360 2065
rect 17320 2015 17360 2045
rect 17320 1995 17330 2015
rect 17350 1995 17360 2015
rect 17320 1980 17360 1995
rect 17375 2115 17415 2130
rect 17375 2095 17385 2115
rect 17405 2095 17415 2115
rect 17375 2065 17415 2095
rect 17375 2045 17385 2065
rect 17405 2045 17415 2065
rect 17375 2015 17415 2045
rect 17375 1995 17385 2015
rect 17405 1995 17415 2015
rect 17375 1980 17415 1995
rect 17430 2115 17470 2130
rect 17430 2095 17440 2115
rect 17460 2095 17470 2115
rect 17430 2065 17470 2095
rect 17430 2045 17440 2065
rect 17460 2045 17470 2065
rect 17430 2015 17470 2045
rect 17430 1995 17440 2015
rect 17460 1995 17470 2015
rect 17430 1980 17470 1995
rect 17485 2115 17525 2130
rect 17485 2095 17495 2115
rect 17515 2095 17525 2115
rect 17485 2065 17525 2095
rect 17485 2045 17495 2065
rect 17515 2045 17525 2065
rect 17485 2015 17525 2045
rect 17485 1995 17495 2015
rect 17515 1995 17525 2015
rect 17485 1980 17525 1995
rect 18145 2100 18185 2130
rect 18145 2080 18155 2100
rect 18175 2080 18185 2100
rect 18145 2050 18185 2080
rect 18145 2030 18155 2050
rect 18175 2030 18185 2050
rect 18145 2000 18185 2030
rect 18145 1980 18155 2000
rect 18175 1980 18185 2000
rect 15665 1965 15705 1980
rect 18145 1965 18185 1980
rect 18200 2250 18240 2265
rect 18200 2230 18210 2250
rect 18230 2230 18240 2250
rect 18200 2200 18240 2230
rect 18200 2180 18210 2200
rect 18230 2180 18240 2200
rect 18200 2150 18240 2180
rect 18200 2130 18210 2150
rect 18230 2130 18240 2150
rect 18200 2100 18240 2130
rect 18200 2080 18210 2100
rect 18230 2080 18240 2100
rect 18200 2050 18240 2080
rect 18200 2030 18210 2050
rect 18230 2030 18240 2050
rect 18200 2000 18240 2030
rect 18200 1980 18210 2000
rect 18230 1980 18240 2000
rect 18200 1965 18240 1980
rect 18255 2250 18295 2265
rect 18255 2230 18265 2250
rect 18285 2230 18295 2250
rect 18255 2200 18295 2230
rect 18255 2180 18265 2200
rect 18285 2180 18295 2200
rect 18255 2150 18295 2180
rect 18255 2130 18265 2150
rect 18285 2130 18295 2150
rect 18255 2100 18295 2130
rect 18255 2080 18265 2100
rect 18285 2080 18295 2100
rect 18255 2050 18295 2080
rect 18255 2030 18265 2050
rect 18285 2030 18295 2050
rect 18255 2000 18295 2030
rect 18255 1980 18265 2000
rect 18285 1980 18295 2000
rect 18255 1965 18295 1980
rect 18310 2250 18350 2265
rect 18310 2230 18320 2250
rect 18340 2230 18350 2250
rect 18310 2200 18350 2230
rect 18310 2180 18320 2200
rect 18340 2180 18350 2200
rect 18310 2150 18350 2180
rect 18310 2130 18320 2150
rect 18340 2130 18350 2150
rect 18310 2100 18350 2130
rect 18310 2080 18320 2100
rect 18340 2080 18350 2100
rect 18310 2050 18350 2080
rect 18310 2030 18320 2050
rect 18340 2030 18350 2050
rect 18310 2000 18350 2030
rect 18310 1980 18320 2000
rect 18340 1980 18350 2000
rect 18310 1965 18350 1980
rect 18365 2250 18405 2265
rect 18365 2230 18375 2250
rect 18395 2230 18405 2250
rect 18365 2200 18405 2230
rect 18365 2180 18375 2200
rect 18395 2180 18405 2200
rect 18365 2150 18405 2180
rect 18365 2130 18375 2150
rect 18395 2130 18405 2150
rect 18365 2100 18405 2130
rect 18365 2080 18375 2100
rect 18395 2080 18405 2100
rect 18365 2050 18405 2080
rect 18365 2030 18375 2050
rect 18395 2030 18405 2050
rect 18365 2000 18405 2030
rect 18365 1980 18375 2000
rect 18395 1980 18405 2000
rect 18365 1965 18405 1980
rect 18420 2250 18460 2265
rect 18420 2230 18430 2250
rect 18450 2230 18460 2250
rect 18420 2200 18460 2230
rect 18420 2180 18430 2200
rect 18450 2180 18460 2200
rect 18420 2150 18460 2180
rect 18420 2130 18430 2150
rect 18450 2130 18460 2150
rect 18420 2100 18460 2130
rect 18420 2080 18430 2100
rect 18450 2080 18460 2100
rect 18420 2050 18460 2080
rect 18420 2030 18430 2050
rect 18450 2030 18460 2050
rect 18420 2000 18460 2030
rect 18420 1980 18430 2000
rect 18450 1980 18460 2000
rect 18420 1965 18460 1980
rect 18475 2250 18515 2265
rect 18475 2230 18485 2250
rect 18505 2230 18515 2250
rect 18475 2200 18515 2230
rect 18475 2180 18485 2200
rect 18505 2180 18515 2200
rect 18475 2150 18515 2180
rect 18475 2130 18485 2150
rect 18505 2130 18515 2150
rect 18475 2100 18515 2130
rect 18475 2080 18485 2100
rect 18505 2080 18515 2100
rect 18475 2050 18515 2080
rect 18475 2030 18485 2050
rect 18505 2030 18515 2050
rect 18475 2000 18515 2030
rect 18475 1980 18485 2000
rect 18505 1980 18515 2000
rect 18475 1965 18515 1980
rect 18530 2250 18570 2265
rect 18530 2230 18540 2250
rect 18560 2230 18570 2250
rect 18530 2200 18570 2230
rect 18530 2180 18540 2200
rect 18560 2180 18570 2200
rect 18530 2150 18570 2180
rect 18530 2130 18540 2150
rect 18560 2130 18570 2150
rect 18530 2100 18570 2130
rect 18530 2080 18540 2100
rect 18560 2080 18570 2100
rect 18530 2050 18570 2080
rect 18530 2030 18540 2050
rect 18560 2030 18570 2050
rect 18530 2000 18570 2030
rect 18530 1980 18540 2000
rect 18560 1980 18570 2000
rect 18530 1965 18570 1980
rect 18585 2250 18625 2265
rect 18585 2230 18595 2250
rect 18615 2230 18625 2250
rect 18585 2200 18625 2230
rect 18585 2180 18595 2200
rect 18615 2180 18625 2200
rect 18585 2150 18625 2180
rect 18585 2130 18595 2150
rect 18615 2130 18625 2150
rect 18585 2100 18625 2130
rect 18585 2080 18595 2100
rect 18615 2080 18625 2100
rect 18585 2050 18625 2080
rect 18585 2030 18595 2050
rect 18615 2030 18625 2050
rect 18585 2000 18625 2030
rect 18585 1980 18595 2000
rect 18615 1980 18625 2000
rect 18585 1965 18625 1980
rect 18640 2250 18680 2265
rect 18640 2230 18650 2250
rect 18670 2230 18680 2250
rect 18640 2200 18680 2230
rect 18640 2180 18650 2200
rect 18670 2180 18680 2200
rect 18640 2150 18680 2180
rect 18640 2130 18650 2150
rect 18670 2130 18680 2150
rect 18640 2100 18680 2130
rect 18640 2080 18650 2100
rect 18670 2080 18680 2100
rect 18640 2050 18680 2080
rect 18640 2030 18650 2050
rect 18670 2030 18680 2050
rect 18640 2000 18680 2030
rect 18640 1980 18650 2000
rect 18670 1980 18680 2000
rect 18640 1965 18680 1980
rect 18695 2250 18735 2265
rect 18695 2230 18705 2250
rect 18725 2230 18735 2250
rect 18695 2200 18735 2230
rect 18695 2180 18705 2200
rect 18725 2180 18735 2200
rect 18695 2150 18735 2180
rect 18695 2130 18705 2150
rect 18725 2130 18735 2150
rect 18695 2100 18735 2130
rect 18695 2080 18705 2100
rect 18725 2080 18735 2100
rect 18695 2050 18735 2080
rect 18695 2030 18705 2050
rect 18725 2030 18735 2050
rect 18695 2000 18735 2030
rect 18695 1980 18705 2000
rect 18725 1980 18735 2000
rect 18695 1965 18735 1980
rect 18750 2250 18790 2265
rect 18750 2230 18760 2250
rect 18780 2230 18790 2250
rect 18750 2200 18790 2230
rect 18750 2180 18760 2200
rect 18780 2180 18790 2200
rect 18750 2150 18790 2180
rect 18750 2130 18760 2150
rect 18780 2130 18790 2150
rect 18750 2100 18790 2130
rect 18750 2080 18760 2100
rect 18780 2080 18790 2100
rect 18750 2050 18790 2080
rect 18750 2030 18760 2050
rect 18780 2030 18790 2050
rect 18750 2000 18790 2030
rect 18750 1980 18760 2000
rect 18780 1980 18790 2000
rect 18750 1965 18790 1980
rect 18805 2250 18845 2265
rect 18805 2230 18815 2250
rect 18835 2230 18845 2250
rect 18805 2200 18845 2230
rect 18805 2180 18815 2200
rect 18835 2180 18845 2200
rect 18805 2150 18845 2180
rect 18805 2130 18815 2150
rect 18835 2130 18845 2150
rect 18805 2100 18845 2130
rect 18805 2080 18815 2100
rect 18835 2080 18845 2100
rect 18805 2050 18845 2080
rect 18805 2030 18815 2050
rect 18835 2030 18845 2050
rect 18805 2000 18845 2030
rect 25005 2250 25045 2265
rect 25005 2230 25015 2250
rect 25035 2230 25045 2250
rect 25005 2200 25045 2230
rect 25005 2180 25015 2200
rect 25035 2180 25045 2200
rect 25005 2150 25045 2180
rect 25005 2130 25015 2150
rect 25035 2130 25045 2150
rect 25005 2100 25045 2130
rect 25005 2080 25015 2100
rect 25035 2080 25045 2100
rect 25005 2050 25045 2080
rect 25005 2030 25015 2050
rect 25035 2030 25045 2050
rect 18805 1980 18815 2000
rect 18835 1980 18845 2000
rect 18805 1965 18845 1980
rect 25005 2000 25045 2030
rect 25005 1980 25015 2000
rect 25035 1980 25045 2000
rect 25005 1965 25045 1980
rect 25060 2250 25100 2265
rect 25060 2230 25070 2250
rect 25090 2230 25100 2250
rect 25060 2200 25100 2230
rect 25060 2180 25070 2200
rect 25090 2180 25100 2200
rect 25060 2150 25100 2180
rect 25060 2130 25070 2150
rect 25090 2130 25100 2150
rect 25060 2100 25100 2130
rect 25060 2080 25070 2100
rect 25090 2080 25100 2100
rect 25060 2050 25100 2080
rect 25060 2030 25070 2050
rect 25090 2030 25100 2050
rect 25060 2000 25100 2030
rect 25060 1980 25070 2000
rect 25090 1980 25100 2000
rect 25060 1965 25100 1980
rect 25115 2250 25155 2265
rect 25115 2230 25125 2250
rect 25145 2230 25155 2250
rect 25115 2200 25155 2230
rect 25115 2180 25125 2200
rect 25145 2180 25155 2200
rect 25115 2150 25155 2180
rect 25115 2130 25125 2150
rect 25145 2130 25155 2150
rect 25115 2100 25155 2130
rect 25115 2080 25125 2100
rect 25145 2080 25155 2100
rect 25115 2050 25155 2080
rect 25115 2030 25125 2050
rect 25145 2030 25155 2050
rect 25115 2000 25155 2030
rect 25115 1980 25125 2000
rect 25145 1980 25155 2000
rect 25115 1965 25155 1980
rect 25170 2250 25210 2265
rect 25170 2230 25180 2250
rect 25200 2230 25210 2250
rect 25170 2200 25210 2230
rect 25170 2180 25180 2200
rect 25200 2180 25210 2200
rect 25170 2150 25210 2180
rect 25170 2130 25180 2150
rect 25200 2130 25210 2150
rect 25170 2100 25210 2130
rect 25170 2080 25180 2100
rect 25200 2080 25210 2100
rect 25170 2050 25210 2080
rect 25170 2030 25180 2050
rect 25200 2030 25210 2050
rect 25170 2000 25210 2030
rect 25170 1980 25180 2000
rect 25200 1980 25210 2000
rect 25170 1965 25210 1980
rect 25225 2250 25265 2265
rect 25225 2230 25235 2250
rect 25255 2230 25265 2250
rect 25225 2200 25265 2230
rect 25225 2180 25235 2200
rect 25255 2180 25265 2200
rect 25225 2150 25265 2180
rect 25225 2130 25235 2150
rect 25255 2130 25265 2150
rect 25225 2100 25265 2130
rect 25225 2080 25235 2100
rect 25255 2080 25265 2100
rect 25225 2050 25265 2080
rect 25225 2030 25235 2050
rect 25255 2030 25265 2050
rect 25225 2000 25265 2030
rect 25225 1980 25235 2000
rect 25255 1980 25265 2000
rect 25225 1965 25265 1980
rect 25280 2250 25320 2265
rect 25280 2230 25290 2250
rect 25310 2230 25320 2250
rect 25280 2200 25320 2230
rect 25280 2180 25290 2200
rect 25310 2180 25320 2200
rect 25280 2150 25320 2180
rect 25280 2130 25290 2150
rect 25310 2130 25320 2150
rect 25280 2100 25320 2130
rect 25280 2080 25290 2100
rect 25310 2080 25320 2100
rect 25280 2050 25320 2080
rect 25280 2030 25290 2050
rect 25310 2030 25320 2050
rect 25280 2000 25320 2030
rect 25280 1980 25290 2000
rect 25310 1980 25320 2000
rect 25280 1965 25320 1980
rect 25335 2250 25375 2265
rect 25335 2230 25345 2250
rect 25365 2230 25375 2250
rect 25335 2200 25375 2230
rect 25335 2180 25345 2200
rect 25365 2180 25375 2200
rect 25335 2150 25375 2180
rect 25335 2130 25345 2150
rect 25365 2130 25375 2150
rect 25335 2100 25375 2130
rect 25335 2080 25345 2100
rect 25365 2080 25375 2100
rect 25335 2050 25375 2080
rect 25335 2030 25345 2050
rect 25365 2030 25375 2050
rect 25335 2000 25375 2030
rect 25335 1980 25345 2000
rect 25365 1980 25375 2000
rect 25335 1965 25375 1980
rect 25390 2250 25430 2265
rect 25390 2230 25400 2250
rect 25420 2230 25430 2250
rect 25390 2200 25430 2230
rect 25390 2180 25400 2200
rect 25420 2180 25430 2200
rect 25390 2150 25430 2180
rect 25390 2130 25400 2150
rect 25420 2130 25430 2150
rect 25390 2100 25430 2130
rect 25390 2080 25400 2100
rect 25420 2080 25430 2100
rect 25390 2050 25430 2080
rect 25390 2030 25400 2050
rect 25420 2030 25430 2050
rect 25390 2000 25430 2030
rect 25390 1980 25400 2000
rect 25420 1980 25430 2000
rect 25390 1965 25430 1980
rect 25445 2250 25485 2265
rect 25445 2230 25455 2250
rect 25475 2230 25485 2250
rect 25445 2200 25485 2230
rect 25445 2180 25455 2200
rect 25475 2180 25485 2200
rect 25445 2150 25485 2180
rect 25445 2130 25455 2150
rect 25475 2130 25485 2150
rect 25445 2100 25485 2130
rect 25445 2080 25455 2100
rect 25475 2080 25485 2100
rect 25445 2050 25485 2080
rect 25445 2030 25455 2050
rect 25475 2030 25485 2050
rect 25445 2000 25485 2030
rect 25445 1980 25455 2000
rect 25475 1980 25485 2000
rect 25445 1965 25485 1980
rect 25500 2250 25540 2265
rect 25500 2230 25510 2250
rect 25530 2230 25540 2250
rect 25500 2200 25540 2230
rect 25500 2180 25510 2200
rect 25530 2180 25540 2200
rect 25500 2150 25540 2180
rect 25500 2130 25510 2150
rect 25530 2130 25540 2150
rect 25500 2100 25540 2130
rect 25500 2080 25510 2100
rect 25530 2080 25540 2100
rect 25500 2050 25540 2080
rect 25500 2030 25510 2050
rect 25530 2030 25540 2050
rect 25500 2000 25540 2030
rect 25500 1980 25510 2000
rect 25530 1980 25540 2000
rect 25500 1965 25540 1980
rect 25555 2250 25595 2265
rect 25555 2230 25565 2250
rect 25585 2230 25595 2250
rect 25555 2200 25595 2230
rect 25555 2180 25565 2200
rect 25585 2180 25595 2200
rect 25555 2150 25595 2180
rect 25555 2130 25565 2150
rect 25585 2130 25595 2150
rect 25555 2100 25595 2130
rect 25555 2080 25565 2100
rect 25585 2080 25595 2100
rect 25555 2050 25595 2080
rect 25555 2030 25565 2050
rect 25585 2030 25595 2050
rect 25555 2000 25595 2030
rect 25555 1980 25565 2000
rect 25585 1980 25595 2000
rect 25555 1965 25595 1980
rect 25610 2250 25650 2265
rect 25610 2230 25620 2250
rect 25640 2230 25650 2250
rect 25610 2200 25650 2230
rect 25610 2180 25620 2200
rect 25640 2180 25650 2200
rect 25610 2150 25650 2180
rect 25610 2130 25620 2150
rect 25640 2130 25650 2150
rect 25610 2100 25650 2130
rect 25610 2080 25620 2100
rect 25640 2080 25650 2100
rect 25610 2050 25650 2080
rect 25610 2030 25620 2050
rect 25640 2030 25650 2050
rect 25610 2000 25650 2030
rect 25610 1980 25620 2000
rect 25640 1980 25650 2000
rect 25610 1965 25650 1980
rect 25665 2250 25705 2265
rect 25665 2230 25675 2250
rect 25695 2230 25705 2250
rect 25665 2200 25705 2230
rect 25665 2180 25675 2200
rect 25695 2180 25705 2200
rect 25665 2150 25705 2180
rect 25665 2130 25675 2150
rect 25695 2130 25705 2150
rect 25665 2100 25705 2130
rect 25665 2080 25675 2100
rect 25695 2080 25705 2100
rect 25665 2050 25705 2080
rect 25665 2030 25675 2050
rect 25695 2030 25705 2050
rect 25665 2000 25705 2030
rect 25665 1980 25675 2000
rect 25695 1980 25705 2000
rect 25665 1965 25705 1980
rect 26275 2115 26315 2130
rect 26275 2095 26285 2115
rect 26305 2095 26315 2115
rect 26275 2065 26315 2095
rect 26275 2045 26285 2065
rect 26305 2045 26315 2065
rect 26275 2015 26315 2045
rect 26275 1995 26285 2015
rect 26305 1995 26315 2015
rect 26275 1980 26315 1995
rect 26330 2115 26370 2130
rect 26330 2095 26340 2115
rect 26360 2095 26370 2115
rect 26330 2065 26370 2095
rect 26330 2045 26340 2065
rect 26360 2045 26370 2065
rect 26330 2015 26370 2045
rect 26330 1995 26340 2015
rect 26360 1995 26370 2015
rect 26330 1980 26370 1995
rect 26385 2115 26425 2130
rect 26385 2095 26395 2115
rect 26415 2095 26425 2115
rect 26385 2065 26425 2095
rect 26385 2045 26395 2065
rect 26415 2045 26425 2065
rect 26385 2015 26425 2045
rect 26385 1995 26395 2015
rect 26415 1995 26425 2015
rect 26385 1980 26425 1995
rect 26440 2115 26480 2130
rect 26440 2095 26450 2115
rect 26470 2095 26480 2115
rect 26440 2065 26480 2095
rect 26440 2045 26450 2065
rect 26470 2045 26480 2065
rect 26440 2015 26480 2045
rect 26440 1995 26450 2015
rect 26470 1995 26480 2015
rect 26440 1980 26480 1995
rect 26495 2115 26535 2130
rect 26495 2095 26505 2115
rect 26525 2095 26535 2115
rect 26495 2065 26535 2095
rect 26495 2045 26505 2065
rect 26525 2045 26535 2065
rect 26495 2015 26535 2045
rect 26495 1995 26505 2015
rect 26525 1995 26535 2015
rect 26495 1980 26535 1995
rect 26550 2115 26590 2130
rect 26550 2095 26560 2115
rect 26580 2095 26590 2115
rect 26550 2065 26590 2095
rect 26550 2045 26560 2065
rect 26580 2045 26590 2065
rect 26550 2015 26590 2045
rect 26550 1995 26560 2015
rect 26580 1995 26590 2015
rect 26550 1980 26590 1995
rect 26605 2115 26645 2130
rect 26605 2095 26615 2115
rect 26635 2095 26645 2115
rect 26605 2065 26645 2095
rect 26605 2045 26615 2065
rect 26635 2045 26645 2065
rect 26605 2015 26645 2045
rect 26605 1995 26615 2015
rect 26635 1995 26645 2015
rect 26605 1980 26645 1995
rect 26660 2115 26700 2130
rect 26660 2095 26670 2115
rect 26690 2095 26700 2115
rect 26660 2065 26700 2095
rect 26660 2045 26670 2065
rect 26690 2045 26700 2065
rect 26660 2015 26700 2045
rect 26660 1995 26670 2015
rect 26690 1995 26700 2015
rect 26660 1980 26700 1995
rect 26715 2115 26755 2130
rect 26715 2095 26725 2115
rect 26745 2095 26755 2115
rect 26715 2065 26755 2095
rect 26715 2045 26725 2065
rect 26745 2045 26755 2065
rect 26715 2015 26755 2045
rect 26715 1995 26725 2015
rect 26745 1995 26755 2015
rect 26715 1980 26755 1995
rect 26770 2115 26810 2130
rect 26770 2095 26780 2115
rect 26800 2095 26810 2115
rect 26770 2065 26810 2095
rect 26770 2045 26780 2065
rect 26800 2045 26810 2065
rect 26770 2015 26810 2045
rect 26770 1995 26780 2015
rect 26800 1995 26810 2015
rect 26770 1980 26810 1995
rect 26825 2115 26865 2130
rect 26825 2095 26835 2115
rect 26855 2095 26865 2115
rect 26825 2065 26865 2095
rect 26825 2045 26835 2065
rect 26855 2045 26865 2065
rect 26825 2015 26865 2045
rect 26825 1995 26835 2015
rect 26855 1995 26865 2015
rect 26825 1980 26865 1995
rect 26880 2115 26920 2130
rect 26880 2095 26890 2115
rect 26910 2095 26920 2115
rect 26880 2065 26920 2095
rect 26880 2045 26890 2065
rect 26910 2045 26920 2065
rect 26880 2015 26920 2045
rect 26880 1995 26890 2015
rect 26910 1995 26920 2015
rect 26880 1980 26920 1995
rect 26935 2115 26975 2130
rect 26935 2095 26945 2115
rect 26965 2095 26975 2115
rect 26935 2065 26975 2095
rect 26935 2045 26945 2065
rect 26965 2045 26975 2065
rect 26935 2015 26975 2045
rect 26935 1995 26945 2015
rect 26965 1995 26975 2015
rect 26935 1980 26975 1995
rect 26990 2115 27030 2130
rect 26990 2095 27000 2115
rect 27020 2095 27030 2115
rect 26990 2065 27030 2095
rect 26990 2045 27000 2065
rect 27020 2045 27030 2065
rect 26990 2015 27030 2045
rect 26990 1995 27000 2015
rect 27020 1995 27030 2015
rect 26990 1980 27030 1995
rect 27045 2115 27085 2130
rect 27045 2095 27055 2115
rect 27075 2095 27085 2115
rect 27045 2065 27085 2095
rect 27045 2045 27055 2065
rect 27075 2045 27085 2065
rect 27045 2015 27085 2045
rect 27045 1995 27055 2015
rect 27075 1995 27085 2015
rect 27045 1980 27085 1995
rect 27100 2115 27140 2130
rect 27100 2095 27110 2115
rect 27130 2095 27140 2115
rect 27100 2065 27140 2095
rect 27100 2045 27110 2065
rect 27130 2045 27140 2065
rect 27100 2015 27140 2045
rect 27100 1995 27110 2015
rect 27130 1995 27140 2015
rect 27100 1980 27140 1995
rect 27155 2115 27195 2130
rect 27155 2095 27165 2115
rect 27185 2095 27195 2115
rect 27155 2065 27195 2095
rect 27155 2045 27165 2065
rect 27185 2045 27195 2065
rect 27155 2015 27195 2045
rect 27155 1995 27165 2015
rect 27185 1995 27195 2015
rect 27155 1980 27195 1995
rect 27210 2115 27250 2130
rect 27210 2095 27220 2115
rect 27240 2095 27250 2115
rect 27210 2065 27250 2095
rect 27210 2045 27220 2065
rect 27240 2045 27250 2065
rect 27210 2015 27250 2045
rect 27210 1995 27220 2015
rect 27240 1995 27250 2015
rect 27210 1980 27250 1995
rect 27265 2115 27305 2130
rect 27265 2095 27275 2115
rect 27295 2095 27305 2115
rect 27265 2065 27305 2095
rect 27265 2045 27275 2065
rect 27295 2045 27305 2065
rect 27265 2015 27305 2045
rect 27265 1995 27275 2015
rect 27295 1995 27305 2015
rect 27265 1980 27305 1995
rect 27320 2115 27360 2130
rect 27320 2095 27330 2115
rect 27350 2095 27360 2115
rect 27320 2065 27360 2095
rect 27320 2045 27330 2065
rect 27350 2045 27360 2065
rect 27320 2015 27360 2045
rect 27320 1995 27330 2015
rect 27350 1995 27360 2015
rect 27320 1980 27360 1995
rect 27375 2115 27415 2130
rect 27375 2095 27385 2115
rect 27405 2095 27415 2115
rect 27375 2065 27415 2095
rect 27375 2045 27385 2065
rect 27405 2045 27415 2065
rect 27375 2015 27415 2045
rect 27375 1995 27385 2015
rect 27405 1995 27415 2015
rect 27375 1980 27415 1995
rect 27430 2115 27470 2130
rect 27430 2095 27440 2115
rect 27460 2095 27470 2115
rect 27430 2065 27470 2095
rect 27430 2045 27440 2065
rect 27460 2045 27470 2065
rect 27430 2015 27470 2045
rect 27430 1995 27440 2015
rect 27460 1995 27470 2015
rect 27430 1980 27470 1995
rect 27485 2115 27525 2130
rect 27485 2095 27495 2115
rect 27515 2095 27525 2115
rect 27485 2065 27525 2095
rect 27485 2045 27495 2065
rect 27515 2045 27525 2065
rect 27485 2015 27525 2045
rect 27485 1995 27495 2015
rect 27515 1995 27525 2015
rect 27485 1980 27525 1995
rect 28145 2230 28185 2245
rect 28145 2210 28155 2230
rect 28175 2210 28185 2230
rect 28145 2180 28185 2210
rect 28145 2160 28155 2180
rect 28175 2160 28185 2180
rect 28145 2130 28185 2160
rect 28145 2110 28155 2130
rect 28175 2110 28185 2130
rect 28145 2080 28185 2110
rect 28145 2060 28155 2080
rect 28175 2060 28185 2080
rect 28145 2030 28185 2060
rect 28145 2010 28155 2030
rect 28175 2010 28185 2030
rect 28145 1980 28185 2010
rect 28145 1960 28155 1980
rect 28175 1960 28185 1980
rect 28145 1945 28185 1960
rect 28200 2230 28240 2245
rect 28200 2210 28210 2230
rect 28230 2210 28240 2230
rect 28200 2180 28240 2210
rect 28200 2160 28210 2180
rect 28230 2160 28240 2180
rect 28200 2130 28240 2160
rect 28200 2110 28210 2130
rect 28230 2110 28240 2130
rect 28200 2080 28240 2110
rect 28200 2060 28210 2080
rect 28230 2060 28240 2080
rect 28200 2030 28240 2060
rect 28200 2010 28210 2030
rect 28230 2010 28240 2030
rect 28200 1980 28240 2010
rect 28200 1960 28210 1980
rect 28230 1960 28240 1980
rect 28200 1945 28240 1960
rect 28255 2230 28295 2245
rect 28255 2210 28265 2230
rect 28285 2210 28295 2230
rect 28255 2180 28295 2210
rect 28255 2160 28265 2180
rect 28285 2160 28295 2180
rect 28255 2130 28295 2160
rect 28255 2110 28265 2130
rect 28285 2110 28295 2130
rect 28255 2080 28295 2110
rect 28255 2060 28265 2080
rect 28285 2060 28295 2080
rect 28255 2030 28295 2060
rect 28255 2010 28265 2030
rect 28285 2010 28295 2030
rect 28255 1980 28295 2010
rect 28255 1960 28265 1980
rect 28285 1960 28295 1980
rect 28255 1945 28295 1960
rect 28310 2230 28350 2245
rect 28310 2210 28320 2230
rect 28340 2210 28350 2230
rect 28310 2180 28350 2210
rect 28310 2160 28320 2180
rect 28340 2160 28350 2180
rect 28310 2130 28350 2160
rect 28310 2110 28320 2130
rect 28340 2110 28350 2130
rect 28310 2080 28350 2110
rect 28310 2060 28320 2080
rect 28340 2060 28350 2080
rect 28310 2030 28350 2060
rect 28310 2010 28320 2030
rect 28340 2010 28350 2030
rect 28310 1980 28350 2010
rect 28310 1960 28320 1980
rect 28340 1960 28350 1980
rect 28310 1945 28350 1960
rect 28365 2230 28405 2245
rect 28365 2210 28375 2230
rect 28395 2210 28405 2230
rect 28365 2180 28405 2210
rect 28365 2160 28375 2180
rect 28395 2160 28405 2180
rect 28365 2130 28405 2160
rect 28365 2110 28375 2130
rect 28395 2110 28405 2130
rect 28365 2080 28405 2110
rect 28365 2060 28375 2080
rect 28395 2060 28405 2080
rect 28365 2030 28405 2060
rect 28365 2010 28375 2030
rect 28395 2010 28405 2030
rect 28365 1980 28405 2010
rect 28365 1960 28375 1980
rect 28395 1960 28405 1980
rect 28365 1945 28405 1960
rect 28420 2230 28460 2245
rect 28420 2210 28430 2230
rect 28450 2210 28460 2230
rect 28420 2180 28460 2210
rect 28420 2160 28430 2180
rect 28450 2160 28460 2180
rect 28420 2130 28460 2160
rect 28420 2110 28430 2130
rect 28450 2110 28460 2130
rect 28420 2080 28460 2110
rect 28420 2060 28430 2080
rect 28450 2060 28460 2080
rect 28420 2030 28460 2060
rect 28420 2010 28430 2030
rect 28450 2010 28460 2030
rect 28420 1980 28460 2010
rect 28420 1960 28430 1980
rect 28450 1960 28460 1980
rect 28420 1945 28460 1960
rect 28475 2230 28515 2245
rect 28475 2210 28485 2230
rect 28505 2210 28515 2230
rect 28475 2180 28515 2210
rect 28475 2160 28485 2180
rect 28505 2160 28515 2180
rect 28475 2130 28515 2160
rect 28475 2110 28485 2130
rect 28505 2110 28515 2130
rect 28475 2080 28515 2110
rect 28475 2060 28485 2080
rect 28505 2060 28515 2080
rect 28475 2030 28515 2060
rect 28475 2010 28485 2030
rect 28505 2010 28515 2030
rect 28475 1980 28515 2010
rect 28475 1960 28485 1980
rect 28505 1960 28515 1980
rect 28475 1945 28515 1960
rect 28530 2230 28570 2245
rect 28530 2210 28540 2230
rect 28560 2210 28570 2230
rect 28530 2180 28570 2210
rect 28530 2160 28540 2180
rect 28560 2160 28570 2180
rect 28530 2130 28570 2160
rect 28530 2110 28540 2130
rect 28560 2110 28570 2130
rect 28530 2080 28570 2110
rect 28530 2060 28540 2080
rect 28560 2060 28570 2080
rect 28530 2030 28570 2060
rect 28530 2010 28540 2030
rect 28560 2010 28570 2030
rect 28530 1980 28570 2010
rect 28530 1960 28540 1980
rect 28560 1960 28570 1980
rect 28530 1945 28570 1960
rect 28585 2230 28625 2245
rect 28585 2210 28595 2230
rect 28615 2210 28625 2230
rect 28585 2180 28625 2210
rect 28585 2160 28595 2180
rect 28615 2160 28625 2180
rect 28585 2130 28625 2160
rect 28585 2110 28595 2130
rect 28615 2110 28625 2130
rect 28585 2080 28625 2110
rect 28585 2060 28595 2080
rect 28615 2060 28625 2080
rect 28585 2030 28625 2060
rect 28585 2010 28595 2030
rect 28615 2010 28625 2030
rect 28585 1980 28625 2010
rect 28585 1960 28595 1980
rect 28615 1960 28625 1980
rect 28585 1945 28625 1960
rect 28640 2230 28680 2245
rect 28640 2210 28650 2230
rect 28670 2210 28680 2230
rect 28640 2180 28680 2210
rect 28640 2160 28650 2180
rect 28670 2160 28680 2180
rect 28640 2130 28680 2160
rect 28640 2110 28650 2130
rect 28670 2110 28680 2130
rect 28640 2080 28680 2110
rect 28640 2060 28650 2080
rect 28670 2060 28680 2080
rect 28640 2030 28680 2060
rect 28640 2010 28650 2030
rect 28670 2010 28680 2030
rect 28640 1980 28680 2010
rect 28640 1960 28650 1980
rect 28670 1960 28680 1980
rect 28640 1945 28680 1960
rect 28695 2230 28735 2245
rect 28695 2210 28705 2230
rect 28725 2210 28735 2230
rect 28695 2180 28735 2210
rect 28695 2160 28705 2180
rect 28725 2160 28735 2180
rect 28695 2130 28735 2160
rect 28695 2110 28705 2130
rect 28725 2110 28735 2130
rect 28695 2080 28735 2110
rect 28695 2060 28705 2080
rect 28725 2060 28735 2080
rect 28695 2030 28735 2060
rect 28695 2010 28705 2030
rect 28725 2010 28735 2030
rect 28695 1980 28735 2010
rect 28695 1960 28705 1980
rect 28725 1960 28735 1980
rect 28695 1945 28735 1960
rect 28750 2230 28790 2245
rect 28750 2210 28760 2230
rect 28780 2210 28790 2230
rect 28750 2180 28790 2210
rect 28750 2160 28760 2180
rect 28780 2160 28790 2180
rect 28750 2130 28790 2160
rect 28750 2110 28760 2130
rect 28780 2110 28790 2130
rect 28750 2080 28790 2110
rect 28750 2060 28760 2080
rect 28780 2060 28790 2080
rect 28750 2030 28790 2060
rect 28750 2010 28760 2030
rect 28780 2010 28790 2030
rect 28750 1980 28790 2010
rect 28750 1960 28760 1980
rect 28780 1960 28790 1980
rect 28750 1945 28790 1960
rect 28805 2230 28845 2245
rect 28805 2210 28815 2230
rect 28835 2210 28845 2230
rect 28805 2180 28845 2210
rect 28805 2160 28815 2180
rect 28835 2160 28845 2180
rect 28805 2130 28845 2160
rect 28805 2110 28815 2130
rect 28835 2110 28845 2130
rect 28805 2080 28845 2110
rect 28805 2060 28815 2080
rect 28835 2060 28845 2080
rect 28805 2030 28845 2060
rect 28805 2010 28815 2030
rect 28835 2010 28845 2030
rect 28805 1980 28845 2010
rect 28805 1960 28815 1980
rect 28835 1960 28845 1980
rect 28805 1945 28845 1960
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 4805 1650 4845 1665
rect 4805 1630 4815 1650
rect 4835 1630 4845 1650
rect 4805 1615 4845 1630
rect 15005 1640 15045 1655
rect 15005 1620 15015 1640
rect 15035 1620 15045 1640
rect 2835 1440 2875 1455
rect 2835 1420 2845 1440
rect 2865 1420 2875 1440
rect 2835 1390 2875 1420
rect 2835 1370 2845 1390
rect 2865 1370 2875 1390
rect 2835 1340 2875 1370
rect 2835 1320 2845 1340
rect 2865 1320 2875 1340
rect 2835 1290 2875 1320
rect 2835 1270 2845 1290
rect 2865 1270 2875 1290
rect 2835 1240 2875 1270
rect 2835 1220 2845 1240
rect 2865 1220 2875 1240
rect 2835 1205 2875 1220
rect 3375 1440 3415 1455
rect 3375 1420 3385 1440
rect 3405 1420 3415 1440
rect 3375 1390 3415 1420
rect 3375 1370 3385 1390
rect 3405 1370 3415 1390
rect 3375 1340 3415 1370
rect 3375 1320 3385 1340
rect 3405 1320 3415 1340
rect 3375 1290 3415 1320
rect 3375 1270 3385 1290
rect 3405 1270 3415 1290
rect 3375 1240 3415 1270
rect 3375 1220 3385 1240
rect 3405 1220 3415 1240
rect 3375 1205 3415 1220
rect 3915 1440 3955 1455
rect 3915 1420 3925 1440
rect 3945 1420 3955 1440
rect 3915 1390 3955 1420
rect 3915 1370 3925 1390
rect 3945 1370 3955 1390
rect 3915 1340 3955 1370
rect 3915 1320 3925 1340
rect 3945 1320 3955 1340
rect 3915 1290 3955 1320
rect 3915 1270 3925 1290
rect 3945 1270 3955 1290
rect 3915 1240 3955 1270
rect 3915 1220 3925 1240
rect 3945 1220 3955 1240
rect 3915 1205 3955 1220
rect 4055 1440 4095 1455
rect 4055 1420 4065 1440
rect 4085 1420 4095 1440
rect 4055 1390 4095 1420
rect 4055 1370 4065 1390
rect 4085 1370 4095 1390
rect 4055 1340 4095 1370
rect 4055 1320 4065 1340
rect 4085 1320 4095 1340
rect 4055 1290 4095 1320
rect 4055 1270 4065 1290
rect 4085 1270 4095 1290
rect 4055 1240 4095 1270
rect 4055 1220 4065 1240
rect 4085 1220 4095 1240
rect 4055 1205 4095 1220
rect 4595 1440 4635 1455
rect 4595 1420 4605 1440
rect 4625 1420 4635 1440
rect 4595 1390 4635 1420
rect 4595 1370 4605 1390
rect 4625 1370 4635 1390
rect 4595 1340 4635 1370
rect 4595 1320 4605 1340
rect 4625 1320 4635 1340
rect 4595 1290 4635 1320
rect 4595 1270 4605 1290
rect 4625 1270 4635 1290
rect 4595 1240 4635 1270
rect 4595 1220 4605 1240
rect 4625 1220 4635 1240
rect 4595 1205 4635 1220
rect 5135 1440 5175 1455
rect 5135 1420 5145 1440
rect 5165 1420 5175 1440
rect 5135 1390 5175 1420
rect 5135 1370 5145 1390
rect 5165 1370 5175 1390
rect 5135 1340 5175 1370
rect 5135 1320 5145 1340
rect 5165 1320 5175 1340
rect 5135 1290 5175 1320
rect 5135 1270 5145 1290
rect 5165 1270 5175 1290
rect 5135 1240 5175 1270
rect 5135 1220 5145 1240
rect 5165 1220 5175 1240
rect 5135 1205 5175 1220
rect 2945 1060 2985 1075
rect 2945 1040 2955 1060
rect 2975 1040 2985 1060
rect 2945 1010 2985 1040
rect 2945 990 2955 1010
rect 2975 990 2985 1010
rect 2945 975 2985 990
rect 3985 1060 4025 1075
rect 3985 1040 3995 1060
rect 4015 1040 4025 1060
rect 3985 1010 4025 1040
rect 3985 990 3995 1010
rect 4015 990 4025 1010
rect 3985 975 4025 990
rect 5025 1060 5065 1075
rect 5025 1040 5035 1060
rect 5055 1040 5065 1060
rect 5025 1010 5065 1040
rect 5025 990 5035 1010
rect 5055 990 5065 1010
rect 5025 975 5065 990
rect 15005 1590 15045 1620
rect 15005 1570 15015 1590
rect 15035 1570 15045 1590
rect 15005 1540 15045 1570
rect 15005 1520 15015 1540
rect 15035 1520 15045 1540
rect 15005 1490 15045 1520
rect 15005 1470 15015 1490
rect 15035 1470 15045 1490
rect 15005 1440 15045 1470
rect 15005 1420 15015 1440
rect 15035 1420 15045 1440
rect 15005 1390 15045 1420
rect 15005 1370 15015 1390
rect 15035 1370 15045 1390
rect 15005 1340 15045 1370
rect 15005 1320 15015 1340
rect 15035 1320 15045 1340
rect 15005 1290 15045 1320
rect 15005 1270 15015 1290
rect 15035 1270 15045 1290
rect 15005 1240 15045 1270
rect 15005 1220 15015 1240
rect 15035 1220 15045 1240
rect 15005 1190 15045 1220
rect 15005 1170 15015 1190
rect 15035 1170 15045 1190
rect 15005 1140 15045 1170
rect 15005 1120 15015 1140
rect 15035 1120 15045 1140
rect 15005 1090 15045 1120
rect 15005 1070 15015 1090
rect 15035 1070 15045 1090
rect 15005 1040 15045 1070
rect 15005 1020 15015 1040
rect 15035 1020 15045 1040
rect 15005 990 15045 1020
rect 15005 970 15015 990
rect 15035 970 15045 990
rect 15005 955 15045 970
rect 15105 1640 15145 1655
rect 15105 1620 15115 1640
rect 15135 1620 15145 1640
rect 15105 1590 15145 1620
rect 15105 1570 15115 1590
rect 15135 1570 15145 1590
rect 15105 1540 15145 1570
rect 15105 1520 15115 1540
rect 15135 1520 15145 1540
rect 15105 1490 15145 1520
rect 15105 1470 15115 1490
rect 15135 1470 15145 1490
rect 15105 1440 15145 1470
rect 15105 1420 15115 1440
rect 15135 1420 15145 1440
rect 15105 1390 15145 1420
rect 15105 1370 15115 1390
rect 15135 1370 15145 1390
rect 15105 1340 15145 1370
rect 15105 1320 15115 1340
rect 15135 1320 15145 1340
rect 15105 1290 15145 1320
rect 15105 1270 15115 1290
rect 15135 1270 15145 1290
rect 15105 1240 15145 1270
rect 15105 1220 15115 1240
rect 15135 1220 15145 1240
rect 15105 1190 15145 1220
rect 15105 1170 15115 1190
rect 15135 1170 15145 1190
rect 15105 1140 15145 1170
rect 15105 1120 15115 1140
rect 15135 1120 15145 1140
rect 15105 1090 15145 1120
rect 15105 1070 15115 1090
rect 15135 1070 15145 1090
rect 15105 1040 15145 1070
rect 15105 1020 15115 1040
rect 15135 1020 15145 1040
rect 15105 990 15145 1020
rect 15105 970 15115 990
rect 15135 970 15145 990
rect 15105 955 15145 970
rect 15205 1640 15245 1655
rect 15205 1620 15215 1640
rect 15235 1620 15245 1640
rect 15205 1590 15245 1620
rect 15205 1570 15215 1590
rect 15235 1570 15245 1590
rect 15205 1540 15245 1570
rect 15205 1520 15215 1540
rect 15235 1520 15245 1540
rect 15205 1490 15245 1520
rect 15205 1470 15215 1490
rect 15235 1470 15245 1490
rect 15205 1440 15245 1470
rect 15205 1420 15215 1440
rect 15235 1420 15245 1440
rect 15205 1390 15245 1420
rect 15205 1370 15215 1390
rect 15235 1370 15245 1390
rect 15205 1340 15245 1370
rect 15205 1320 15215 1340
rect 15235 1320 15245 1340
rect 15205 1290 15245 1320
rect 15205 1270 15215 1290
rect 15235 1270 15245 1290
rect 15205 1240 15245 1270
rect 15205 1220 15215 1240
rect 15235 1220 15245 1240
rect 15205 1190 15245 1220
rect 15205 1170 15215 1190
rect 15235 1170 15245 1190
rect 15205 1140 15245 1170
rect 15205 1120 15215 1140
rect 15235 1120 15245 1140
rect 15205 1090 15245 1120
rect 15205 1070 15215 1090
rect 15235 1070 15245 1090
rect 15205 1040 15245 1070
rect 15205 1020 15215 1040
rect 15235 1020 15245 1040
rect 15205 990 15245 1020
rect 15205 970 15215 990
rect 15235 970 15245 990
rect 15205 955 15245 970
rect 15305 1640 15345 1655
rect 15305 1620 15315 1640
rect 15335 1620 15345 1640
rect 15305 1590 15345 1620
rect 15305 1570 15315 1590
rect 15335 1570 15345 1590
rect 15305 1540 15345 1570
rect 15305 1520 15315 1540
rect 15335 1520 15345 1540
rect 15305 1490 15345 1520
rect 15305 1470 15315 1490
rect 15335 1470 15345 1490
rect 15305 1440 15345 1470
rect 15305 1420 15315 1440
rect 15335 1420 15345 1440
rect 15305 1390 15345 1420
rect 15305 1370 15315 1390
rect 15335 1370 15345 1390
rect 15305 1340 15345 1370
rect 15305 1320 15315 1340
rect 15335 1320 15345 1340
rect 15305 1290 15345 1320
rect 15305 1270 15315 1290
rect 15335 1270 15345 1290
rect 15305 1240 15345 1270
rect 15305 1220 15315 1240
rect 15335 1220 15345 1240
rect 15305 1190 15345 1220
rect 15305 1170 15315 1190
rect 15335 1170 15345 1190
rect 15305 1140 15345 1170
rect 15305 1120 15315 1140
rect 15335 1120 15345 1140
rect 15305 1090 15345 1120
rect 15305 1070 15315 1090
rect 15335 1070 15345 1090
rect 15305 1040 15345 1070
rect 15305 1020 15315 1040
rect 15335 1020 15345 1040
rect 15305 990 15345 1020
rect 15305 970 15315 990
rect 15335 970 15345 990
rect 15305 955 15345 970
rect 15405 1640 15445 1655
rect 15405 1620 15415 1640
rect 15435 1620 15445 1640
rect 15405 1590 15445 1620
rect 15405 1570 15415 1590
rect 15435 1570 15445 1590
rect 15405 1540 15445 1570
rect 15405 1520 15415 1540
rect 15435 1520 15445 1540
rect 15405 1490 15445 1520
rect 15405 1470 15415 1490
rect 15435 1470 15445 1490
rect 15405 1440 15445 1470
rect 15405 1420 15415 1440
rect 15435 1420 15445 1440
rect 15405 1390 15445 1420
rect 15405 1370 15415 1390
rect 15435 1370 15445 1390
rect 15405 1340 15445 1370
rect 15405 1320 15415 1340
rect 15435 1320 15445 1340
rect 15405 1290 15445 1320
rect 15405 1270 15415 1290
rect 15435 1270 15445 1290
rect 15405 1240 15445 1270
rect 15405 1220 15415 1240
rect 15435 1220 15445 1240
rect 15405 1190 15445 1220
rect 15405 1170 15415 1190
rect 15435 1170 15445 1190
rect 15405 1140 15445 1170
rect 15405 1120 15415 1140
rect 15435 1120 15445 1140
rect 15405 1090 15445 1120
rect 15405 1070 15415 1090
rect 15435 1070 15445 1090
rect 15405 1040 15445 1070
rect 15405 1020 15415 1040
rect 15435 1020 15445 1040
rect 15405 990 15445 1020
rect 15405 970 15415 990
rect 15435 970 15445 990
rect 15405 955 15445 970
rect 15505 1640 15545 1655
rect 15505 1620 15515 1640
rect 15535 1620 15545 1640
rect 15505 1590 15545 1620
rect 15505 1570 15515 1590
rect 15535 1570 15545 1590
rect 15505 1540 15545 1570
rect 15505 1520 15515 1540
rect 15535 1520 15545 1540
rect 15505 1490 15545 1520
rect 15505 1470 15515 1490
rect 15535 1470 15545 1490
rect 15505 1440 15545 1470
rect 15505 1420 15515 1440
rect 15535 1420 15545 1440
rect 15505 1390 15545 1420
rect 15505 1370 15515 1390
rect 15535 1370 15545 1390
rect 15505 1340 15545 1370
rect 15505 1320 15515 1340
rect 15535 1320 15545 1340
rect 15505 1290 15545 1320
rect 15505 1270 15515 1290
rect 15535 1270 15545 1290
rect 15505 1240 15545 1270
rect 15505 1220 15515 1240
rect 15535 1220 15545 1240
rect 15505 1190 15545 1220
rect 15505 1170 15515 1190
rect 15535 1170 15545 1190
rect 15505 1140 15545 1170
rect 15505 1120 15515 1140
rect 15535 1120 15545 1140
rect 15505 1090 15545 1120
rect 15505 1070 15515 1090
rect 15535 1070 15545 1090
rect 15505 1040 15545 1070
rect 15505 1020 15515 1040
rect 15535 1020 15545 1040
rect 15505 990 15545 1020
rect 15505 970 15515 990
rect 15535 970 15545 990
rect 15505 955 15545 970
rect 15605 1640 15645 1655
rect 15605 1620 15615 1640
rect 15635 1620 15645 1640
rect 15605 1590 15645 1620
rect 15605 1570 15615 1590
rect 15635 1570 15645 1590
rect 15605 1540 15645 1570
rect 15605 1520 15615 1540
rect 15635 1520 15645 1540
rect 15605 1490 15645 1520
rect 16030 1650 16070 1665
rect 16030 1630 16040 1650
rect 16060 1630 16070 1650
rect 16030 1600 16070 1630
rect 16030 1580 16040 1600
rect 16060 1580 16070 1600
rect 16030 1550 16070 1580
rect 16030 1530 16040 1550
rect 16060 1530 16070 1550
rect 16030 1515 16070 1530
rect 16085 1650 16125 1665
rect 16085 1630 16095 1650
rect 16115 1630 16125 1650
rect 16085 1600 16125 1630
rect 16085 1580 16095 1600
rect 16115 1580 16125 1600
rect 16085 1550 16125 1580
rect 16085 1530 16095 1550
rect 16115 1530 16125 1550
rect 16085 1515 16125 1530
rect 16140 1650 16180 1665
rect 16140 1630 16150 1650
rect 16170 1630 16180 1650
rect 16140 1600 16180 1630
rect 16140 1580 16150 1600
rect 16170 1580 16180 1600
rect 16140 1550 16180 1580
rect 16140 1530 16150 1550
rect 16170 1530 16180 1550
rect 16140 1515 16180 1530
rect 16195 1650 16235 1665
rect 16195 1630 16205 1650
rect 16225 1630 16235 1650
rect 16195 1600 16235 1630
rect 16195 1580 16205 1600
rect 16225 1580 16235 1600
rect 16195 1550 16235 1580
rect 16195 1530 16205 1550
rect 16225 1530 16235 1550
rect 16195 1515 16235 1530
rect 16250 1650 16290 1665
rect 16250 1630 16260 1650
rect 16280 1630 16290 1650
rect 16250 1600 16290 1630
rect 16250 1580 16260 1600
rect 16280 1580 16290 1600
rect 16250 1550 16290 1580
rect 16250 1530 16260 1550
rect 16280 1530 16290 1550
rect 16250 1515 16290 1530
rect 16305 1650 16345 1665
rect 16305 1630 16315 1650
rect 16335 1630 16345 1650
rect 16305 1600 16345 1630
rect 16305 1580 16315 1600
rect 16335 1580 16345 1600
rect 16305 1550 16345 1580
rect 16305 1530 16315 1550
rect 16335 1530 16345 1550
rect 16305 1515 16345 1530
rect 16360 1650 16400 1665
rect 16360 1630 16370 1650
rect 16390 1630 16400 1650
rect 16360 1600 16400 1630
rect 16360 1580 16370 1600
rect 16390 1580 16400 1600
rect 16360 1550 16400 1580
rect 16360 1530 16370 1550
rect 16390 1530 16400 1550
rect 16360 1515 16400 1530
rect 16415 1650 16455 1665
rect 16415 1630 16425 1650
rect 16445 1630 16455 1650
rect 16415 1600 16455 1630
rect 16415 1580 16425 1600
rect 16445 1580 16455 1600
rect 16415 1550 16455 1580
rect 16415 1530 16425 1550
rect 16445 1530 16455 1550
rect 16415 1515 16455 1530
rect 16470 1650 16510 1665
rect 16470 1630 16480 1650
rect 16500 1630 16510 1650
rect 16470 1600 16510 1630
rect 16470 1580 16480 1600
rect 16500 1580 16510 1600
rect 16470 1550 16510 1580
rect 16470 1530 16480 1550
rect 16500 1530 16510 1550
rect 16470 1515 16510 1530
rect 16525 1650 16565 1665
rect 16525 1630 16535 1650
rect 16555 1630 16565 1650
rect 16525 1600 16565 1630
rect 16525 1580 16535 1600
rect 16555 1580 16565 1600
rect 16525 1550 16565 1580
rect 16525 1530 16535 1550
rect 16555 1530 16565 1550
rect 16525 1515 16565 1530
rect 16580 1650 16620 1665
rect 16580 1630 16590 1650
rect 16610 1630 16620 1650
rect 16580 1600 16620 1630
rect 16580 1580 16590 1600
rect 16610 1580 16620 1600
rect 16580 1550 16620 1580
rect 16580 1530 16590 1550
rect 16610 1530 16620 1550
rect 16580 1515 16620 1530
rect 16635 1650 16675 1665
rect 16635 1630 16645 1650
rect 16665 1630 16675 1650
rect 16635 1600 16675 1630
rect 16635 1580 16645 1600
rect 16665 1580 16675 1600
rect 16635 1550 16675 1580
rect 16635 1530 16645 1550
rect 16665 1530 16675 1550
rect 16635 1515 16675 1530
rect 16690 1650 16730 1665
rect 16770 1650 16810 1665
rect 16690 1630 16700 1650
rect 16720 1630 16730 1650
rect 16770 1630 16780 1650
rect 16800 1630 16810 1650
rect 16690 1600 16730 1630
rect 16770 1600 16810 1630
rect 16690 1580 16700 1600
rect 16720 1580 16730 1600
rect 16770 1580 16780 1600
rect 16800 1580 16810 1600
rect 16690 1550 16730 1580
rect 16770 1550 16810 1580
rect 16690 1530 16700 1550
rect 16720 1530 16730 1550
rect 16770 1530 16780 1550
rect 16800 1530 16810 1550
rect 16690 1515 16730 1530
rect 16770 1515 16810 1530
rect 16825 1650 16865 1665
rect 16825 1630 16835 1650
rect 16855 1630 16865 1650
rect 16825 1600 16865 1630
rect 16825 1580 16835 1600
rect 16855 1580 16865 1600
rect 16825 1550 16865 1580
rect 16825 1530 16835 1550
rect 16855 1530 16865 1550
rect 16825 1515 16865 1530
rect 16880 1650 16920 1665
rect 16880 1630 16890 1650
rect 16910 1630 16920 1650
rect 16880 1600 16920 1630
rect 16880 1580 16890 1600
rect 16910 1580 16920 1600
rect 16880 1550 16920 1580
rect 16880 1530 16890 1550
rect 16910 1530 16920 1550
rect 16880 1515 16920 1530
rect 16935 1650 16975 1665
rect 16935 1630 16945 1650
rect 16965 1630 16975 1650
rect 16935 1600 16975 1630
rect 16935 1580 16945 1600
rect 16965 1580 16975 1600
rect 16935 1550 16975 1580
rect 16935 1530 16945 1550
rect 16965 1530 16975 1550
rect 16935 1515 16975 1530
rect 16990 1650 17030 1665
rect 17070 1650 17110 1665
rect 16990 1630 17000 1650
rect 17020 1630 17030 1650
rect 17070 1630 17080 1650
rect 17100 1630 17110 1650
rect 16990 1600 17030 1630
rect 17070 1600 17110 1630
rect 16990 1580 17000 1600
rect 17020 1580 17030 1600
rect 17070 1580 17080 1600
rect 17100 1580 17110 1600
rect 16990 1550 17030 1580
rect 17070 1550 17110 1580
rect 16990 1530 17000 1550
rect 17020 1530 17030 1550
rect 17070 1530 17080 1550
rect 17100 1530 17110 1550
rect 16990 1515 17030 1530
rect 17070 1515 17110 1530
rect 17125 1650 17165 1665
rect 17125 1630 17135 1650
rect 17155 1630 17165 1650
rect 17125 1600 17165 1630
rect 17125 1580 17135 1600
rect 17155 1580 17165 1600
rect 17125 1550 17165 1580
rect 17125 1530 17135 1550
rect 17155 1530 17165 1550
rect 17125 1515 17165 1530
rect 17180 1650 17220 1665
rect 17180 1630 17190 1650
rect 17210 1630 17220 1650
rect 17180 1600 17220 1630
rect 17180 1580 17190 1600
rect 17210 1580 17220 1600
rect 17180 1550 17220 1580
rect 17180 1530 17190 1550
rect 17210 1530 17220 1550
rect 17180 1515 17220 1530
rect 17235 1650 17275 1665
rect 17235 1630 17245 1650
rect 17265 1630 17275 1650
rect 17235 1600 17275 1630
rect 17235 1580 17245 1600
rect 17265 1580 17275 1600
rect 17235 1550 17275 1580
rect 17235 1530 17245 1550
rect 17265 1530 17275 1550
rect 17235 1515 17275 1530
rect 17290 1650 17330 1665
rect 17290 1630 17300 1650
rect 17320 1630 17330 1650
rect 17290 1600 17330 1630
rect 17290 1580 17300 1600
rect 17320 1580 17330 1600
rect 17290 1550 17330 1580
rect 17290 1530 17300 1550
rect 17320 1530 17330 1550
rect 17290 1515 17330 1530
rect 17345 1650 17385 1665
rect 17345 1630 17355 1650
rect 17375 1630 17385 1650
rect 17345 1600 17385 1630
rect 17345 1580 17355 1600
rect 17375 1580 17385 1600
rect 17345 1550 17385 1580
rect 17345 1530 17355 1550
rect 17375 1530 17385 1550
rect 17345 1515 17385 1530
rect 17400 1650 17440 1665
rect 17400 1630 17410 1650
rect 17430 1630 17440 1650
rect 17400 1600 17440 1630
rect 17400 1580 17410 1600
rect 17430 1580 17440 1600
rect 17400 1550 17440 1580
rect 17400 1530 17410 1550
rect 17430 1530 17440 1550
rect 17400 1515 17440 1530
rect 17455 1650 17495 1665
rect 17455 1630 17465 1650
rect 17485 1630 17495 1650
rect 17455 1600 17495 1630
rect 17455 1580 17465 1600
rect 17485 1580 17495 1600
rect 17455 1550 17495 1580
rect 17455 1530 17465 1550
rect 17485 1530 17495 1550
rect 17455 1515 17495 1530
rect 17510 1650 17550 1665
rect 17510 1630 17520 1650
rect 17540 1630 17550 1650
rect 17510 1600 17550 1630
rect 17510 1580 17520 1600
rect 17540 1580 17550 1600
rect 17510 1550 17550 1580
rect 17510 1530 17520 1550
rect 17540 1530 17550 1550
rect 17510 1515 17550 1530
rect 17565 1650 17605 1665
rect 17565 1630 17575 1650
rect 17595 1630 17605 1650
rect 17565 1600 17605 1630
rect 17565 1580 17575 1600
rect 17595 1580 17605 1600
rect 17565 1550 17605 1580
rect 17565 1530 17575 1550
rect 17595 1530 17605 1550
rect 17565 1515 17605 1530
rect 17620 1650 17660 1665
rect 17620 1630 17630 1650
rect 17650 1630 17660 1650
rect 17620 1600 17660 1630
rect 17620 1580 17630 1600
rect 17650 1580 17660 1600
rect 17620 1550 17660 1580
rect 17620 1530 17630 1550
rect 17650 1530 17660 1550
rect 17620 1515 17660 1530
rect 17675 1650 17715 1665
rect 17675 1630 17685 1650
rect 17705 1630 17715 1650
rect 17675 1600 17715 1630
rect 17675 1580 17685 1600
rect 17705 1580 17715 1600
rect 17675 1550 17715 1580
rect 17675 1530 17685 1550
rect 17705 1530 17715 1550
rect 17675 1515 17715 1530
rect 17730 1650 17770 1665
rect 17730 1630 17740 1650
rect 17760 1630 17770 1650
rect 17730 1600 17770 1630
rect 17730 1580 17740 1600
rect 17760 1580 17770 1600
rect 17730 1550 17770 1580
rect 17730 1530 17740 1550
rect 17760 1530 17770 1550
rect 17730 1515 17770 1530
rect 18205 1640 18245 1655
rect 18205 1620 18215 1640
rect 18235 1620 18245 1640
rect 18205 1590 18245 1620
rect 18205 1570 18215 1590
rect 18235 1570 18245 1590
rect 18205 1540 18245 1570
rect 18205 1520 18215 1540
rect 18235 1520 18245 1540
rect 15605 1470 15615 1490
rect 15635 1470 15645 1490
rect 15605 1440 15645 1470
rect 18205 1490 18245 1520
rect 18205 1470 18215 1490
rect 18235 1470 18245 1490
rect 15605 1420 15615 1440
rect 15635 1420 15645 1440
rect 15605 1390 15645 1420
rect 15605 1370 15615 1390
rect 15635 1370 15645 1390
rect 15605 1340 15645 1370
rect 15605 1320 15615 1340
rect 15635 1320 15645 1340
rect 15605 1290 15645 1320
rect 15605 1270 15615 1290
rect 15635 1270 15645 1290
rect 15605 1240 15645 1270
rect 18205 1440 18245 1470
rect 18205 1420 18215 1440
rect 18235 1420 18245 1440
rect 18205 1390 18245 1420
rect 18205 1370 18215 1390
rect 18235 1370 18245 1390
rect 18205 1340 18245 1370
rect 18205 1320 18215 1340
rect 18235 1320 18245 1340
rect 18205 1290 18245 1320
rect 18205 1270 18215 1290
rect 18235 1270 18245 1290
rect 15605 1220 15615 1240
rect 15635 1220 15645 1240
rect 15605 1190 15645 1220
rect 15605 1170 15615 1190
rect 15635 1170 15645 1190
rect 18205 1240 18245 1270
rect 18205 1220 18215 1240
rect 18235 1220 18245 1240
rect 18205 1190 18245 1220
rect 15605 1140 15645 1170
rect 15605 1120 15615 1140
rect 15635 1120 15645 1140
rect 15605 1090 15645 1120
rect 15605 1070 15615 1090
rect 15635 1070 15645 1090
rect 15605 1040 15645 1070
rect 15605 1020 15615 1040
rect 15635 1020 15645 1040
rect 15605 990 15645 1020
rect 15605 970 15615 990
rect 15635 970 15645 990
rect 15605 955 15645 970
rect 16205 1170 16245 1185
rect 16205 1150 16215 1170
rect 16235 1150 16245 1170
rect 16205 1120 16245 1150
rect 16205 1100 16215 1120
rect 16235 1100 16245 1120
rect 16205 1070 16245 1100
rect 16205 1050 16215 1070
rect 16235 1050 16245 1070
rect 16205 1020 16245 1050
rect 16205 1000 16215 1020
rect 16235 1000 16245 1020
rect 16205 970 16245 1000
rect 16205 950 16215 970
rect 16235 950 16245 970
rect 16205 935 16245 950
rect 16260 1170 16300 1185
rect 16260 1150 16270 1170
rect 16290 1150 16300 1170
rect 16260 1120 16300 1150
rect 16260 1100 16270 1120
rect 16290 1100 16300 1120
rect 16260 1070 16300 1100
rect 16260 1050 16270 1070
rect 16290 1050 16300 1070
rect 16260 1020 16300 1050
rect 16260 1000 16270 1020
rect 16290 1000 16300 1020
rect 16260 970 16300 1000
rect 16260 950 16270 970
rect 16290 950 16300 970
rect 16260 935 16300 950
rect 16315 1170 16355 1185
rect 16315 1150 16325 1170
rect 16345 1150 16355 1170
rect 16315 1120 16355 1150
rect 16315 1100 16325 1120
rect 16345 1100 16355 1120
rect 16315 1070 16355 1100
rect 16315 1050 16325 1070
rect 16345 1050 16355 1070
rect 16315 1020 16355 1050
rect 16315 1000 16325 1020
rect 16345 1000 16355 1020
rect 16315 970 16355 1000
rect 16315 950 16325 970
rect 16345 950 16355 970
rect 16315 935 16355 950
rect 16370 1170 16410 1185
rect 16370 1150 16380 1170
rect 16400 1150 16410 1170
rect 16370 1120 16410 1150
rect 16370 1100 16380 1120
rect 16400 1100 16410 1120
rect 16370 1070 16410 1100
rect 16370 1050 16380 1070
rect 16400 1050 16410 1070
rect 16370 1020 16410 1050
rect 16370 1000 16380 1020
rect 16400 1000 16410 1020
rect 16370 970 16410 1000
rect 16370 950 16380 970
rect 16400 950 16410 970
rect 16370 935 16410 950
rect 16425 1170 16465 1185
rect 16425 1150 16435 1170
rect 16455 1150 16465 1170
rect 16425 1120 16465 1150
rect 16425 1100 16435 1120
rect 16455 1100 16465 1120
rect 16425 1070 16465 1100
rect 16425 1050 16435 1070
rect 16455 1050 16465 1070
rect 16425 1020 16465 1050
rect 16425 1000 16435 1020
rect 16455 1000 16465 1020
rect 16425 970 16465 1000
rect 16425 950 16435 970
rect 16455 950 16465 970
rect 16425 935 16465 950
rect 16480 1170 16520 1185
rect 16480 1150 16490 1170
rect 16510 1150 16520 1170
rect 16480 1120 16520 1150
rect 16480 1100 16490 1120
rect 16510 1100 16520 1120
rect 16480 1070 16520 1100
rect 16480 1050 16490 1070
rect 16510 1050 16520 1070
rect 16480 1020 16520 1050
rect 16480 1000 16490 1020
rect 16510 1000 16520 1020
rect 16480 970 16520 1000
rect 16480 950 16490 970
rect 16510 950 16520 970
rect 16480 935 16520 950
rect 16535 1170 16575 1185
rect 16535 1150 16545 1170
rect 16565 1150 16575 1170
rect 16535 1120 16575 1150
rect 16535 1100 16545 1120
rect 16565 1100 16575 1120
rect 16535 1070 16575 1100
rect 16535 1050 16545 1070
rect 16565 1050 16575 1070
rect 16535 1020 16575 1050
rect 16535 1000 16545 1020
rect 16565 1000 16575 1020
rect 16535 970 16575 1000
rect 16535 950 16545 970
rect 16565 950 16575 970
rect 16535 935 16575 950
rect 16590 1170 16630 1185
rect 16590 1150 16600 1170
rect 16620 1150 16630 1170
rect 16590 1120 16630 1150
rect 16590 1100 16600 1120
rect 16620 1100 16630 1120
rect 16590 1070 16630 1100
rect 16590 1050 16600 1070
rect 16620 1050 16630 1070
rect 16590 1020 16630 1050
rect 16590 1000 16600 1020
rect 16620 1000 16630 1020
rect 16590 970 16630 1000
rect 16590 950 16600 970
rect 16620 950 16630 970
rect 16590 935 16630 950
rect 16645 1170 16685 1185
rect 16645 1150 16655 1170
rect 16675 1150 16685 1170
rect 16645 1120 16685 1150
rect 16645 1100 16655 1120
rect 16675 1100 16685 1120
rect 16645 1070 16685 1100
rect 16645 1050 16655 1070
rect 16675 1050 16685 1070
rect 16645 1020 16685 1050
rect 16645 1000 16655 1020
rect 16675 1000 16685 1020
rect 16645 970 16685 1000
rect 16645 950 16655 970
rect 16675 950 16685 970
rect 16645 935 16685 950
rect 16700 1170 16740 1185
rect 16700 1150 16710 1170
rect 16730 1150 16740 1170
rect 16700 1120 16740 1150
rect 16700 1100 16710 1120
rect 16730 1100 16740 1120
rect 16700 1070 16740 1100
rect 16700 1050 16710 1070
rect 16730 1050 16740 1070
rect 16700 1020 16740 1050
rect 16700 1000 16710 1020
rect 16730 1000 16740 1020
rect 16700 970 16740 1000
rect 16700 950 16710 970
rect 16730 950 16740 970
rect 16700 935 16740 950
rect 16755 1170 16795 1185
rect 16755 1150 16765 1170
rect 16785 1150 16795 1170
rect 16755 1120 16795 1150
rect 16755 1100 16765 1120
rect 16785 1100 16795 1120
rect 16755 1070 16795 1100
rect 16755 1050 16765 1070
rect 16785 1050 16795 1070
rect 16755 1020 16795 1050
rect 16755 1000 16765 1020
rect 16785 1000 16795 1020
rect 16755 970 16795 1000
rect 16755 950 16765 970
rect 16785 950 16795 970
rect 16755 935 16795 950
rect 16810 1170 16850 1185
rect 16810 1150 16820 1170
rect 16840 1150 16850 1170
rect 16810 1120 16850 1150
rect 16810 1100 16820 1120
rect 16840 1100 16850 1120
rect 16810 1070 16850 1100
rect 16810 1050 16820 1070
rect 16840 1050 16850 1070
rect 16810 1020 16850 1050
rect 16810 1000 16820 1020
rect 16840 1000 16850 1020
rect 16810 970 16850 1000
rect 16810 950 16820 970
rect 16840 950 16850 970
rect 16810 935 16850 950
rect 16865 1170 16905 1185
rect 16865 1150 16875 1170
rect 16895 1150 16905 1170
rect 16865 1120 16905 1150
rect 16865 1100 16875 1120
rect 16895 1100 16905 1120
rect 16865 1070 16905 1100
rect 16865 1050 16875 1070
rect 16895 1050 16905 1070
rect 16865 1020 16905 1050
rect 16865 1000 16875 1020
rect 16895 1000 16905 1020
rect 16865 970 16905 1000
rect 16865 950 16875 970
rect 16895 950 16905 970
rect 16865 935 16905 950
rect 16920 1170 16960 1185
rect 16920 1150 16930 1170
rect 16950 1150 16960 1170
rect 16920 1120 16960 1150
rect 16920 1100 16930 1120
rect 16950 1100 16960 1120
rect 16920 1070 16960 1100
rect 16920 1050 16930 1070
rect 16950 1050 16960 1070
rect 16920 1020 16960 1050
rect 16920 1000 16930 1020
rect 16950 1000 16960 1020
rect 16920 970 16960 1000
rect 16920 950 16930 970
rect 16950 950 16960 970
rect 16920 935 16960 950
rect 16975 1170 17015 1185
rect 16975 1150 16985 1170
rect 17005 1150 17015 1170
rect 16975 1120 17015 1150
rect 16975 1100 16985 1120
rect 17005 1100 17015 1120
rect 16975 1070 17015 1100
rect 16975 1050 16985 1070
rect 17005 1050 17015 1070
rect 16975 1020 17015 1050
rect 16975 1000 16985 1020
rect 17005 1000 17015 1020
rect 16975 970 17015 1000
rect 16975 950 16985 970
rect 17005 950 17015 970
rect 16975 935 17015 950
rect 17030 1170 17070 1185
rect 17030 1150 17040 1170
rect 17060 1150 17070 1170
rect 17030 1120 17070 1150
rect 17030 1100 17040 1120
rect 17060 1100 17070 1120
rect 17030 1070 17070 1100
rect 17030 1050 17040 1070
rect 17060 1050 17070 1070
rect 17030 1020 17070 1050
rect 17030 1000 17040 1020
rect 17060 1000 17070 1020
rect 17030 970 17070 1000
rect 17030 950 17040 970
rect 17060 950 17070 970
rect 17030 935 17070 950
rect 17085 1170 17125 1185
rect 17085 1150 17095 1170
rect 17115 1150 17125 1170
rect 17085 1120 17125 1150
rect 17085 1100 17095 1120
rect 17115 1100 17125 1120
rect 17085 1070 17125 1100
rect 17085 1050 17095 1070
rect 17115 1050 17125 1070
rect 17085 1020 17125 1050
rect 17085 1000 17095 1020
rect 17115 1000 17125 1020
rect 17085 970 17125 1000
rect 17085 950 17095 970
rect 17115 950 17125 970
rect 17085 935 17125 950
rect 17140 1170 17180 1185
rect 17140 1150 17150 1170
rect 17170 1150 17180 1170
rect 17140 1120 17180 1150
rect 17140 1100 17150 1120
rect 17170 1100 17180 1120
rect 17140 1070 17180 1100
rect 17140 1050 17150 1070
rect 17170 1050 17180 1070
rect 17140 1020 17180 1050
rect 17140 1000 17150 1020
rect 17170 1000 17180 1020
rect 17140 970 17180 1000
rect 17140 950 17150 970
rect 17170 950 17180 970
rect 17140 935 17180 950
rect 17195 1170 17235 1185
rect 17195 1150 17205 1170
rect 17225 1150 17235 1170
rect 17195 1120 17235 1150
rect 17195 1100 17205 1120
rect 17225 1100 17235 1120
rect 17195 1070 17235 1100
rect 17195 1050 17205 1070
rect 17225 1050 17235 1070
rect 17195 1020 17235 1050
rect 17195 1000 17205 1020
rect 17225 1000 17235 1020
rect 17195 970 17235 1000
rect 17195 950 17205 970
rect 17225 950 17235 970
rect 17195 935 17235 950
rect 17250 1170 17290 1185
rect 17250 1150 17260 1170
rect 17280 1150 17290 1170
rect 17250 1120 17290 1150
rect 17250 1100 17260 1120
rect 17280 1100 17290 1120
rect 17250 1070 17290 1100
rect 17250 1050 17260 1070
rect 17280 1050 17290 1070
rect 17250 1020 17290 1050
rect 17250 1000 17260 1020
rect 17280 1000 17290 1020
rect 17250 970 17290 1000
rect 17250 950 17260 970
rect 17280 950 17290 970
rect 17250 935 17290 950
rect 17305 1170 17345 1185
rect 17305 1150 17315 1170
rect 17335 1150 17345 1170
rect 17305 1120 17345 1150
rect 17305 1100 17315 1120
rect 17335 1100 17345 1120
rect 17305 1070 17345 1100
rect 17305 1050 17315 1070
rect 17335 1050 17345 1070
rect 17305 1020 17345 1050
rect 17305 1000 17315 1020
rect 17335 1000 17345 1020
rect 17305 970 17345 1000
rect 17305 950 17315 970
rect 17335 950 17345 970
rect 17305 935 17345 950
rect 17360 1170 17400 1185
rect 17360 1150 17370 1170
rect 17390 1150 17400 1170
rect 17360 1120 17400 1150
rect 17360 1100 17370 1120
rect 17390 1100 17400 1120
rect 17360 1070 17400 1100
rect 17360 1050 17370 1070
rect 17390 1050 17400 1070
rect 17360 1020 17400 1050
rect 17360 1000 17370 1020
rect 17390 1000 17400 1020
rect 17360 970 17400 1000
rect 17360 950 17370 970
rect 17390 950 17400 970
rect 17360 935 17400 950
rect 17415 1170 17455 1185
rect 17415 1150 17425 1170
rect 17445 1150 17455 1170
rect 17415 1120 17455 1150
rect 17415 1100 17425 1120
rect 17445 1100 17455 1120
rect 17415 1070 17455 1100
rect 17415 1050 17425 1070
rect 17445 1050 17455 1070
rect 17415 1020 17455 1050
rect 17415 1000 17425 1020
rect 17445 1000 17455 1020
rect 17415 970 17455 1000
rect 17415 950 17425 970
rect 17445 950 17455 970
rect 17415 935 17455 950
rect 17470 1170 17510 1185
rect 17470 1150 17480 1170
rect 17500 1150 17510 1170
rect 17470 1120 17510 1150
rect 17470 1100 17480 1120
rect 17500 1100 17510 1120
rect 17470 1070 17510 1100
rect 17470 1050 17480 1070
rect 17500 1050 17510 1070
rect 17470 1020 17510 1050
rect 17470 1000 17480 1020
rect 17500 1000 17510 1020
rect 17470 970 17510 1000
rect 17470 950 17480 970
rect 17500 950 17510 970
rect 17470 935 17510 950
rect 17525 1170 17565 1185
rect 17525 1150 17535 1170
rect 17555 1150 17565 1170
rect 17525 1120 17565 1150
rect 17525 1100 17535 1120
rect 17555 1100 17565 1120
rect 17525 1070 17565 1100
rect 17525 1050 17535 1070
rect 17555 1050 17565 1070
rect 17525 1020 17565 1050
rect 17525 1000 17535 1020
rect 17555 1000 17565 1020
rect 17525 970 17565 1000
rect 17525 950 17535 970
rect 17555 950 17565 970
rect 17525 935 17565 950
rect 17580 1170 17620 1185
rect 17580 1150 17590 1170
rect 17610 1150 17620 1170
rect 17580 1120 17620 1150
rect 17580 1100 17590 1120
rect 17610 1100 17620 1120
rect 17580 1070 17620 1100
rect 17580 1050 17590 1070
rect 17610 1050 17620 1070
rect 17580 1020 17620 1050
rect 17580 1000 17590 1020
rect 17610 1000 17620 1020
rect 17580 970 17620 1000
rect 17580 950 17590 970
rect 17610 950 17620 970
rect 18205 1170 18215 1190
rect 18235 1170 18245 1190
rect 18205 1140 18245 1170
rect 18205 1120 18215 1140
rect 18235 1120 18245 1140
rect 18205 1090 18245 1120
rect 18205 1070 18215 1090
rect 18235 1070 18245 1090
rect 18205 1040 18245 1070
rect 18205 1020 18215 1040
rect 18235 1020 18245 1040
rect 18205 990 18245 1020
rect 18205 970 18215 990
rect 18235 970 18245 990
rect 18205 955 18245 970
rect 18305 1640 18345 1655
rect 18305 1620 18315 1640
rect 18335 1620 18345 1640
rect 18305 1590 18345 1620
rect 18305 1570 18315 1590
rect 18335 1570 18345 1590
rect 18305 1540 18345 1570
rect 18305 1520 18315 1540
rect 18335 1520 18345 1540
rect 18305 1490 18345 1520
rect 18305 1470 18315 1490
rect 18335 1470 18345 1490
rect 18305 1440 18345 1470
rect 18305 1420 18315 1440
rect 18335 1420 18345 1440
rect 18305 1390 18345 1420
rect 18305 1370 18315 1390
rect 18335 1370 18345 1390
rect 18305 1340 18345 1370
rect 18305 1320 18315 1340
rect 18335 1320 18345 1340
rect 18305 1290 18345 1320
rect 18305 1270 18315 1290
rect 18335 1270 18345 1290
rect 18305 1240 18345 1270
rect 18305 1220 18315 1240
rect 18335 1220 18345 1240
rect 18305 1190 18345 1220
rect 18305 1170 18315 1190
rect 18335 1170 18345 1190
rect 18305 1140 18345 1170
rect 18305 1120 18315 1140
rect 18335 1120 18345 1140
rect 18305 1090 18345 1120
rect 18305 1070 18315 1090
rect 18335 1070 18345 1090
rect 18305 1040 18345 1070
rect 18305 1020 18315 1040
rect 18335 1020 18345 1040
rect 18305 990 18345 1020
rect 18305 970 18315 990
rect 18335 970 18345 990
rect 18305 955 18345 970
rect 18405 1640 18445 1655
rect 18405 1620 18415 1640
rect 18435 1620 18445 1640
rect 18405 1590 18445 1620
rect 18405 1570 18415 1590
rect 18435 1570 18445 1590
rect 18405 1540 18445 1570
rect 18405 1520 18415 1540
rect 18435 1520 18445 1540
rect 18405 1490 18445 1520
rect 18405 1470 18415 1490
rect 18435 1470 18445 1490
rect 18405 1440 18445 1470
rect 18405 1420 18415 1440
rect 18435 1420 18445 1440
rect 18405 1390 18445 1420
rect 18405 1370 18415 1390
rect 18435 1370 18445 1390
rect 18405 1340 18445 1370
rect 18405 1320 18415 1340
rect 18435 1320 18445 1340
rect 18405 1290 18445 1320
rect 18405 1270 18415 1290
rect 18435 1270 18445 1290
rect 18405 1240 18445 1270
rect 18405 1220 18415 1240
rect 18435 1220 18445 1240
rect 18405 1190 18445 1220
rect 18405 1170 18415 1190
rect 18435 1170 18445 1190
rect 18405 1140 18445 1170
rect 18405 1120 18415 1140
rect 18435 1120 18445 1140
rect 18405 1090 18445 1120
rect 18405 1070 18415 1090
rect 18435 1070 18445 1090
rect 18405 1040 18445 1070
rect 18405 1020 18415 1040
rect 18435 1020 18445 1040
rect 18405 990 18445 1020
rect 18405 970 18415 990
rect 18435 970 18445 990
rect 18405 955 18445 970
rect 18505 1640 18545 1655
rect 18505 1620 18515 1640
rect 18535 1620 18545 1640
rect 18505 1590 18545 1620
rect 18505 1570 18515 1590
rect 18535 1570 18545 1590
rect 18505 1540 18545 1570
rect 18505 1520 18515 1540
rect 18535 1520 18545 1540
rect 18505 1490 18545 1520
rect 18505 1470 18515 1490
rect 18535 1470 18545 1490
rect 18505 1440 18545 1470
rect 18505 1420 18515 1440
rect 18535 1420 18545 1440
rect 18505 1390 18545 1420
rect 18505 1370 18515 1390
rect 18535 1370 18545 1390
rect 18505 1340 18545 1370
rect 18505 1320 18515 1340
rect 18535 1320 18545 1340
rect 18505 1290 18545 1320
rect 18505 1270 18515 1290
rect 18535 1270 18545 1290
rect 18505 1240 18545 1270
rect 18505 1220 18515 1240
rect 18535 1220 18545 1240
rect 18505 1190 18545 1220
rect 18505 1170 18515 1190
rect 18535 1170 18545 1190
rect 18505 1140 18545 1170
rect 18505 1120 18515 1140
rect 18535 1120 18545 1140
rect 18505 1090 18545 1120
rect 18505 1070 18515 1090
rect 18535 1070 18545 1090
rect 18505 1040 18545 1070
rect 18505 1020 18515 1040
rect 18535 1020 18545 1040
rect 18505 990 18545 1020
rect 18505 970 18515 990
rect 18535 970 18545 990
rect 18505 955 18545 970
rect 18605 1640 18645 1655
rect 18605 1620 18615 1640
rect 18635 1620 18645 1640
rect 18605 1590 18645 1620
rect 18605 1570 18615 1590
rect 18635 1570 18645 1590
rect 18605 1540 18645 1570
rect 18605 1520 18615 1540
rect 18635 1520 18645 1540
rect 18605 1490 18645 1520
rect 18605 1470 18615 1490
rect 18635 1470 18645 1490
rect 18605 1440 18645 1470
rect 18605 1420 18615 1440
rect 18635 1420 18645 1440
rect 18605 1390 18645 1420
rect 18605 1370 18615 1390
rect 18635 1370 18645 1390
rect 18605 1340 18645 1370
rect 18605 1320 18615 1340
rect 18635 1320 18645 1340
rect 18605 1290 18645 1320
rect 18605 1270 18615 1290
rect 18635 1270 18645 1290
rect 18605 1240 18645 1270
rect 18605 1220 18615 1240
rect 18635 1220 18645 1240
rect 18605 1190 18645 1220
rect 18605 1170 18615 1190
rect 18635 1170 18645 1190
rect 18605 1140 18645 1170
rect 18605 1120 18615 1140
rect 18635 1120 18645 1140
rect 18605 1090 18645 1120
rect 18605 1070 18615 1090
rect 18635 1070 18645 1090
rect 18605 1040 18645 1070
rect 18605 1020 18615 1040
rect 18635 1020 18645 1040
rect 18605 990 18645 1020
rect 18605 970 18615 990
rect 18635 970 18645 990
rect 18605 955 18645 970
rect 18705 1640 18745 1655
rect 18705 1620 18715 1640
rect 18735 1620 18745 1640
rect 18705 1590 18745 1620
rect 18705 1570 18715 1590
rect 18735 1570 18745 1590
rect 18705 1540 18745 1570
rect 18705 1520 18715 1540
rect 18735 1520 18745 1540
rect 18705 1490 18745 1520
rect 18705 1470 18715 1490
rect 18735 1470 18745 1490
rect 18705 1440 18745 1470
rect 18705 1420 18715 1440
rect 18735 1420 18745 1440
rect 18705 1390 18745 1420
rect 18705 1370 18715 1390
rect 18735 1370 18745 1390
rect 18705 1340 18745 1370
rect 18705 1320 18715 1340
rect 18735 1320 18745 1340
rect 18705 1290 18745 1320
rect 18705 1270 18715 1290
rect 18735 1270 18745 1290
rect 18705 1240 18745 1270
rect 18705 1220 18715 1240
rect 18735 1220 18745 1240
rect 18705 1190 18745 1220
rect 18705 1170 18715 1190
rect 18735 1170 18745 1190
rect 18705 1140 18745 1170
rect 18705 1120 18715 1140
rect 18735 1120 18745 1140
rect 18705 1090 18745 1120
rect 18705 1070 18715 1090
rect 18735 1070 18745 1090
rect 18705 1040 18745 1070
rect 18705 1020 18715 1040
rect 18735 1020 18745 1040
rect 18705 990 18745 1020
rect 18705 970 18715 990
rect 18735 970 18745 990
rect 18705 955 18745 970
rect 18805 1640 18845 1655
rect 18805 1620 18815 1640
rect 18835 1620 18845 1640
rect 18805 1590 18845 1620
rect 25005 1640 25045 1655
rect 25005 1620 25015 1640
rect 25035 1620 25045 1640
rect 18805 1570 18815 1590
rect 18835 1570 18845 1590
rect 18805 1540 18845 1570
rect 18805 1520 18815 1540
rect 18835 1520 18845 1540
rect 18805 1490 18845 1520
rect 18805 1470 18815 1490
rect 18835 1470 18845 1490
rect 18805 1440 18845 1470
rect 18805 1420 18815 1440
rect 18835 1420 18845 1440
rect 18805 1390 18845 1420
rect 18805 1370 18815 1390
rect 18835 1370 18845 1390
rect 18805 1340 18845 1370
rect 18805 1320 18815 1340
rect 18835 1320 18845 1340
rect 18805 1290 18845 1320
rect 18805 1270 18815 1290
rect 18835 1270 18845 1290
rect 18805 1240 18845 1270
rect 18805 1220 18815 1240
rect 18835 1220 18845 1240
rect 18805 1190 18845 1220
rect 18805 1170 18815 1190
rect 18835 1170 18845 1190
rect 18805 1140 18845 1170
rect 18805 1120 18815 1140
rect 18835 1120 18845 1140
rect 18805 1090 18845 1120
rect 18805 1070 18815 1090
rect 18835 1070 18845 1090
rect 18805 1040 18845 1070
rect 18805 1020 18815 1040
rect 18835 1020 18845 1040
rect 18805 990 18845 1020
rect 18805 970 18815 990
rect 18835 970 18845 990
rect 18805 955 18845 970
rect 17580 935 17620 950
rect 25005 1590 25045 1620
rect 25005 1570 25015 1590
rect 25035 1570 25045 1590
rect 25005 1540 25045 1570
rect 25005 1520 25015 1540
rect 25035 1520 25045 1540
rect 25005 1490 25045 1520
rect 25005 1470 25015 1490
rect 25035 1470 25045 1490
rect 25005 1440 25045 1470
rect 25005 1420 25015 1440
rect 25035 1420 25045 1440
rect 25005 1390 25045 1420
rect 25005 1370 25015 1390
rect 25035 1370 25045 1390
rect 25005 1340 25045 1370
rect 25005 1320 25015 1340
rect 25035 1320 25045 1340
rect 25005 1290 25045 1320
rect 25005 1270 25015 1290
rect 25035 1270 25045 1290
rect 25005 1240 25045 1270
rect 25005 1220 25015 1240
rect 25035 1220 25045 1240
rect 25005 1190 25045 1220
rect 25005 1170 25015 1190
rect 25035 1170 25045 1190
rect 25005 1140 25045 1170
rect 25005 1120 25015 1140
rect 25035 1120 25045 1140
rect 25005 1090 25045 1120
rect 25005 1070 25015 1090
rect 25035 1070 25045 1090
rect 25005 1040 25045 1070
rect 25005 1020 25015 1040
rect 25035 1020 25045 1040
rect 25005 990 25045 1020
rect 25005 970 25015 990
rect 25035 970 25045 990
rect 25005 955 25045 970
rect 25105 1640 25145 1655
rect 25105 1620 25115 1640
rect 25135 1620 25145 1640
rect 25105 1590 25145 1620
rect 25105 1570 25115 1590
rect 25135 1570 25145 1590
rect 25105 1540 25145 1570
rect 25105 1520 25115 1540
rect 25135 1520 25145 1540
rect 25105 1490 25145 1520
rect 25105 1470 25115 1490
rect 25135 1470 25145 1490
rect 25105 1440 25145 1470
rect 25105 1420 25115 1440
rect 25135 1420 25145 1440
rect 25105 1390 25145 1420
rect 25105 1370 25115 1390
rect 25135 1370 25145 1390
rect 25105 1340 25145 1370
rect 25105 1320 25115 1340
rect 25135 1320 25145 1340
rect 25105 1290 25145 1320
rect 25105 1270 25115 1290
rect 25135 1270 25145 1290
rect 25105 1240 25145 1270
rect 25105 1220 25115 1240
rect 25135 1220 25145 1240
rect 25105 1190 25145 1220
rect 25105 1170 25115 1190
rect 25135 1170 25145 1190
rect 25105 1140 25145 1170
rect 25105 1120 25115 1140
rect 25135 1120 25145 1140
rect 25105 1090 25145 1120
rect 25105 1070 25115 1090
rect 25135 1070 25145 1090
rect 25105 1040 25145 1070
rect 25105 1020 25115 1040
rect 25135 1020 25145 1040
rect 25105 990 25145 1020
rect 25105 970 25115 990
rect 25135 970 25145 990
rect 25105 955 25145 970
rect 25205 1640 25245 1655
rect 25205 1620 25215 1640
rect 25235 1620 25245 1640
rect 25205 1590 25245 1620
rect 25205 1570 25215 1590
rect 25235 1570 25245 1590
rect 25205 1540 25245 1570
rect 25205 1520 25215 1540
rect 25235 1520 25245 1540
rect 25205 1490 25245 1520
rect 25205 1470 25215 1490
rect 25235 1470 25245 1490
rect 25205 1440 25245 1470
rect 25205 1420 25215 1440
rect 25235 1420 25245 1440
rect 25205 1390 25245 1420
rect 25205 1370 25215 1390
rect 25235 1370 25245 1390
rect 25205 1340 25245 1370
rect 25205 1320 25215 1340
rect 25235 1320 25245 1340
rect 25205 1290 25245 1320
rect 25205 1270 25215 1290
rect 25235 1270 25245 1290
rect 25205 1240 25245 1270
rect 25205 1220 25215 1240
rect 25235 1220 25245 1240
rect 25205 1190 25245 1220
rect 25205 1170 25215 1190
rect 25235 1170 25245 1190
rect 25205 1140 25245 1170
rect 25205 1120 25215 1140
rect 25235 1120 25245 1140
rect 25205 1090 25245 1120
rect 25205 1070 25215 1090
rect 25235 1070 25245 1090
rect 25205 1040 25245 1070
rect 25205 1020 25215 1040
rect 25235 1020 25245 1040
rect 25205 990 25245 1020
rect 25205 970 25215 990
rect 25235 970 25245 990
rect 25205 955 25245 970
rect 25305 1640 25345 1655
rect 25305 1620 25315 1640
rect 25335 1620 25345 1640
rect 25305 1590 25345 1620
rect 25305 1570 25315 1590
rect 25335 1570 25345 1590
rect 25305 1540 25345 1570
rect 25305 1520 25315 1540
rect 25335 1520 25345 1540
rect 25305 1490 25345 1520
rect 25305 1470 25315 1490
rect 25335 1470 25345 1490
rect 25305 1440 25345 1470
rect 25305 1420 25315 1440
rect 25335 1420 25345 1440
rect 25305 1390 25345 1420
rect 25305 1370 25315 1390
rect 25335 1370 25345 1390
rect 25305 1340 25345 1370
rect 25305 1320 25315 1340
rect 25335 1320 25345 1340
rect 25305 1290 25345 1320
rect 25305 1270 25315 1290
rect 25335 1270 25345 1290
rect 25305 1240 25345 1270
rect 25305 1220 25315 1240
rect 25335 1220 25345 1240
rect 25305 1190 25345 1220
rect 25305 1170 25315 1190
rect 25335 1170 25345 1190
rect 25305 1140 25345 1170
rect 25305 1120 25315 1140
rect 25335 1120 25345 1140
rect 25305 1090 25345 1120
rect 25305 1070 25315 1090
rect 25335 1070 25345 1090
rect 25305 1040 25345 1070
rect 25305 1020 25315 1040
rect 25335 1020 25345 1040
rect 25305 990 25345 1020
rect 25305 970 25315 990
rect 25335 970 25345 990
rect 25305 955 25345 970
rect 25405 1640 25445 1655
rect 25405 1620 25415 1640
rect 25435 1620 25445 1640
rect 25405 1590 25445 1620
rect 25405 1570 25415 1590
rect 25435 1570 25445 1590
rect 25405 1540 25445 1570
rect 25405 1520 25415 1540
rect 25435 1520 25445 1540
rect 25405 1490 25445 1520
rect 25405 1470 25415 1490
rect 25435 1470 25445 1490
rect 25405 1440 25445 1470
rect 25405 1420 25415 1440
rect 25435 1420 25445 1440
rect 25405 1390 25445 1420
rect 25405 1370 25415 1390
rect 25435 1370 25445 1390
rect 25405 1340 25445 1370
rect 25405 1320 25415 1340
rect 25435 1320 25445 1340
rect 25405 1290 25445 1320
rect 25405 1270 25415 1290
rect 25435 1270 25445 1290
rect 25405 1240 25445 1270
rect 25405 1220 25415 1240
rect 25435 1220 25445 1240
rect 25405 1190 25445 1220
rect 25405 1170 25415 1190
rect 25435 1170 25445 1190
rect 25405 1140 25445 1170
rect 25405 1120 25415 1140
rect 25435 1120 25445 1140
rect 25405 1090 25445 1120
rect 25405 1070 25415 1090
rect 25435 1070 25445 1090
rect 25405 1040 25445 1070
rect 25405 1020 25415 1040
rect 25435 1020 25445 1040
rect 25405 990 25445 1020
rect 25405 970 25415 990
rect 25435 970 25445 990
rect 25405 955 25445 970
rect 25505 1640 25545 1655
rect 25505 1620 25515 1640
rect 25535 1620 25545 1640
rect 25505 1590 25545 1620
rect 25505 1570 25515 1590
rect 25535 1570 25545 1590
rect 25505 1540 25545 1570
rect 25505 1520 25515 1540
rect 25535 1520 25545 1540
rect 25505 1490 25545 1520
rect 25505 1470 25515 1490
rect 25535 1470 25545 1490
rect 25505 1440 25545 1470
rect 25505 1420 25515 1440
rect 25535 1420 25545 1440
rect 25505 1390 25545 1420
rect 25505 1370 25515 1390
rect 25535 1370 25545 1390
rect 25505 1340 25545 1370
rect 25505 1320 25515 1340
rect 25535 1320 25545 1340
rect 25505 1290 25545 1320
rect 25505 1270 25515 1290
rect 25535 1270 25545 1290
rect 25505 1240 25545 1270
rect 25505 1220 25515 1240
rect 25535 1220 25545 1240
rect 25505 1190 25545 1220
rect 25505 1170 25515 1190
rect 25535 1170 25545 1190
rect 25505 1140 25545 1170
rect 25505 1120 25515 1140
rect 25535 1120 25545 1140
rect 25505 1090 25545 1120
rect 25505 1070 25515 1090
rect 25535 1070 25545 1090
rect 25505 1040 25545 1070
rect 25505 1020 25515 1040
rect 25535 1020 25545 1040
rect 25505 990 25545 1020
rect 25505 970 25515 990
rect 25535 970 25545 990
rect 25505 955 25545 970
rect 25605 1640 25645 1655
rect 25605 1620 25615 1640
rect 25635 1620 25645 1640
rect 25605 1590 25645 1620
rect 25605 1570 25615 1590
rect 25635 1570 25645 1590
rect 25605 1540 25645 1570
rect 25605 1520 25615 1540
rect 25635 1520 25645 1540
rect 25605 1490 25645 1520
rect 25605 1470 25615 1490
rect 25635 1470 25645 1490
rect 25605 1440 25645 1470
rect 25605 1420 25615 1440
rect 25635 1420 25645 1440
rect 25605 1390 25645 1420
rect 25605 1370 25615 1390
rect 25635 1370 25645 1390
rect 25605 1340 25645 1370
rect 26030 1650 26070 1665
rect 26030 1630 26040 1650
rect 26060 1630 26070 1650
rect 26030 1600 26070 1630
rect 26030 1580 26040 1600
rect 26060 1580 26070 1600
rect 26030 1550 26070 1580
rect 26030 1530 26040 1550
rect 26060 1530 26070 1550
rect 26030 1515 26070 1530
rect 26085 1650 26125 1665
rect 26085 1630 26095 1650
rect 26115 1630 26125 1650
rect 26085 1600 26125 1630
rect 26085 1580 26095 1600
rect 26115 1580 26125 1600
rect 26085 1550 26125 1580
rect 26085 1530 26095 1550
rect 26115 1530 26125 1550
rect 26085 1515 26125 1530
rect 26140 1650 26180 1665
rect 26140 1630 26150 1650
rect 26170 1630 26180 1650
rect 26140 1600 26180 1630
rect 26140 1580 26150 1600
rect 26170 1580 26180 1600
rect 26140 1550 26180 1580
rect 26140 1530 26150 1550
rect 26170 1530 26180 1550
rect 26140 1515 26180 1530
rect 26195 1650 26235 1665
rect 26195 1630 26205 1650
rect 26225 1630 26235 1650
rect 26195 1600 26235 1630
rect 26195 1580 26205 1600
rect 26225 1580 26235 1600
rect 26195 1550 26235 1580
rect 26195 1530 26205 1550
rect 26225 1530 26235 1550
rect 26195 1515 26235 1530
rect 26250 1650 26290 1665
rect 26250 1630 26260 1650
rect 26280 1630 26290 1650
rect 26250 1600 26290 1630
rect 26250 1580 26260 1600
rect 26280 1580 26290 1600
rect 26250 1550 26290 1580
rect 26250 1530 26260 1550
rect 26280 1530 26290 1550
rect 26250 1515 26290 1530
rect 26305 1650 26345 1665
rect 26305 1630 26315 1650
rect 26335 1630 26345 1650
rect 26305 1600 26345 1630
rect 26305 1580 26315 1600
rect 26335 1580 26345 1600
rect 26305 1550 26345 1580
rect 26305 1530 26315 1550
rect 26335 1530 26345 1550
rect 26305 1515 26345 1530
rect 26360 1650 26400 1665
rect 26360 1630 26370 1650
rect 26390 1630 26400 1650
rect 26360 1600 26400 1630
rect 26360 1580 26370 1600
rect 26390 1580 26400 1600
rect 26360 1550 26400 1580
rect 26360 1530 26370 1550
rect 26390 1530 26400 1550
rect 26360 1515 26400 1530
rect 26415 1650 26455 1665
rect 26415 1630 26425 1650
rect 26445 1630 26455 1650
rect 26415 1600 26455 1630
rect 26415 1580 26425 1600
rect 26445 1580 26455 1600
rect 26415 1550 26455 1580
rect 26415 1530 26425 1550
rect 26445 1530 26455 1550
rect 26415 1515 26455 1530
rect 26470 1650 26510 1665
rect 26470 1630 26480 1650
rect 26500 1630 26510 1650
rect 26470 1600 26510 1630
rect 26470 1580 26480 1600
rect 26500 1580 26510 1600
rect 26470 1550 26510 1580
rect 26470 1530 26480 1550
rect 26500 1530 26510 1550
rect 26470 1515 26510 1530
rect 26525 1650 26565 1665
rect 26525 1630 26535 1650
rect 26555 1630 26565 1650
rect 26525 1600 26565 1630
rect 26525 1580 26535 1600
rect 26555 1580 26565 1600
rect 26525 1550 26565 1580
rect 26525 1530 26535 1550
rect 26555 1530 26565 1550
rect 26525 1515 26565 1530
rect 26580 1650 26620 1665
rect 26580 1630 26590 1650
rect 26610 1630 26620 1650
rect 26580 1600 26620 1630
rect 26580 1580 26590 1600
rect 26610 1580 26620 1600
rect 26580 1550 26620 1580
rect 26580 1530 26590 1550
rect 26610 1530 26620 1550
rect 26580 1515 26620 1530
rect 26635 1650 26675 1665
rect 26635 1630 26645 1650
rect 26665 1630 26675 1650
rect 26635 1600 26675 1630
rect 26635 1580 26645 1600
rect 26665 1580 26675 1600
rect 26635 1550 26675 1580
rect 26635 1530 26645 1550
rect 26665 1530 26675 1550
rect 26635 1515 26675 1530
rect 26690 1650 26730 1665
rect 26770 1650 26810 1665
rect 26690 1630 26700 1650
rect 26720 1630 26730 1650
rect 26770 1630 26780 1650
rect 26800 1630 26810 1650
rect 26690 1600 26730 1630
rect 26770 1600 26810 1630
rect 26690 1580 26700 1600
rect 26720 1580 26730 1600
rect 26770 1580 26780 1600
rect 26800 1580 26810 1600
rect 26690 1550 26730 1580
rect 26770 1550 26810 1580
rect 26690 1530 26700 1550
rect 26720 1530 26730 1550
rect 26770 1530 26780 1550
rect 26800 1530 26810 1550
rect 26690 1515 26730 1530
rect 26770 1515 26810 1530
rect 26825 1650 26865 1665
rect 26825 1630 26835 1650
rect 26855 1630 26865 1650
rect 26825 1600 26865 1630
rect 26825 1580 26835 1600
rect 26855 1580 26865 1600
rect 26825 1550 26865 1580
rect 26825 1530 26835 1550
rect 26855 1530 26865 1550
rect 26825 1515 26865 1530
rect 26880 1650 26920 1665
rect 26880 1630 26890 1650
rect 26910 1630 26920 1650
rect 26880 1600 26920 1630
rect 26880 1580 26890 1600
rect 26910 1580 26920 1600
rect 26880 1550 26920 1580
rect 26880 1530 26890 1550
rect 26910 1530 26920 1550
rect 26880 1515 26920 1530
rect 26935 1650 26975 1665
rect 26935 1630 26945 1650
rect 26965 1630 26975 1650
rect 26935 1600 26975 1630
rect 26935 1580 26945 1600
rect 26965 1580 26975 1600
rect 26935 1550 26975 1580
rect 26935 1530 26945 1550
rect 26965 1530 26975 1550
rect 26935 1515 26975 1530
rect 26990 1650 27030 1665
rect 27070 1650 27110 1665
rect 26990 1630 27000 1650
rect 27020 1630 27030 1650
rect 27070 1630 27080 1650
rect 27100 1630 27110 1650
rect 26990 1600 27030 1630
rect 27070 1600 27110 1630
rect 26990 1580 27000 1600
rect 27020 1580 27030 1600
rect 27070 1580 27080 1600
rect 27100 1580 27110 1600
rect 26990 1550 27030 1580
rect 27070 1550 27110 1580
rect 26990 1530 27000 1550
rect 27020 1530 27030 1550
rect 27070 1530 27080 1550
rect 27100 1530 27110 1550
rect 26990 1515 27030 1530
rect 27070 1515 27110 1530
rect 27125 1650 27165 1665
rect 27125 1630 27135 1650
rect 27155 1630 27165 1650
rect 27125 1600 27165 1630
rect 27125 1580 27135 1600
rect 27155 1580 27165 1600
rect 27125 1550 27165 1580
rect 27125 1530 27135 1550
rect 27155 1530 27165 1550
rect 27125 1515 27165 1530
rect 27180 1650 27220 1665
rect 27180 1630 27190 1650
rect 27210 1630 27220 1650
rect 27180 1600 27220 1630
rect 27180 1580 27190 1600
rect 27210 1580 27220 1600
rect 27180 1550 27220 1580
rect 27180 1530 27190 1550
rect 27210 1530 27220 1550
rect 27180 1515 27220 1530
rect 27235 1650 27275 1665
rect 27235 1630 27245 1650
rect 27265 1630 27275 1650
rect 27235 1600 27275 1630
rect 27235 1580 27245 1600
rect 27265 1580 27275 1600
rect 27235 1550 27275 1580
rect 27235 1530 27245 1550
rect 27265 1530 27275 1550
rect 27235 1515 27275 1530
rect 27290 1650 27330 1665
rect 27290 1630 27300 1650
rect 27320 1630 27330 1650
rect 27290 1600 27330 1630
rect 27290 1580 27300 1600
rect 27320 1580 27330 1600
rect 27290 1550 27330 1580
rect 27290 1530 27300 1550
rect 27320 1530 27330 1550
rect 27290 1515 27330 1530
rect 27345 1650 27385 1665
rect 27345 1630 27355 1650
rect 27375 1630 27385 1650
rect 27345 1600 27385 1630
rect 27345 1580 27355 1600
rect 27375 1580 27385 1600
rect 27345 1550 27385 1580
rect 27345 1530 27355 1550
rect 27375 1530 27385 1550
rect 27345 1515 27385 1530
rect 27400 1650 27440 1665
rect 27400 1630 27410 1650
rect 27430 1630 27440 1650
rect 27400 1600 27440 1630
rect 27400 1580 27410 1600
rect 27430 1580 27440 1600
rect 27400 1550 27440 1580
rect 27400 1530 27410 1550
rect 27430 1530 27440 1550
rect 27400 1515 27440 1530
rect 27455 1650 27495 1665
rect 27455 1630 27465 1650
rect 27485 1630 27495 1650
rect 27455 1600 27495 1630
rect 27455 1580 27465 1600
rect 27485 1580 27495 1600
rect 27455 1550 27495 1580
rect 27455 1530 27465 1550
rect 27485 1530 27495 1550
rect 27455 1515 27495 1530
rect 27510 1650 27550 1665
rect 27510 1630 27520 1650
rect 27540 1630 27550 1650
rect 27510 1600 27550 1630
rect 27510 1580 27520 1600
rect 27540 1580 27550 1600
rect 27510 1550 27550 1580
rect 27510 1530 27520 1550
rect 27540 1530 27550 1550
rect 27510 1515 27550 1530
rect 27565 1650 27605 1665
rect 27565 1630 27575 1650
rect 27595 1630 27605 1650
rect 27565 1600 27605 1630
rect 27565 1580 27575 1600
rect 27595 1580 27605 1600
rect 27565 1550 27605 1580
rect 27565 1530 27575 1550
rect 27595 1530 27605 1550
rect 27565 1515 27605 1530
rect 27620 1650 27660 1665
rect 27620 1630 27630 1650
rect 27650 1630 27660 1650
rect 27620 1600 27660 1630
rect 27620 1580 27630 1600
rect 27650 1580 27660 1600
rect 27620 1550 27660 1580
rect 27620 1530 27630 1550
rect 27650 1530 27660 1550
rect 27620 1515 27660 1530
rect 27675 1650 27715 1665
rect 27675 1630 27685 1650
rect 27705 1630 27715 1650
rect 27675 1600 27715 1630
rect 27675 1580 27685 1600
rect 27705 1580 27715 1600
rect 27675 1550 27715 1580
rect 27675 1530 27685 1550
rect 27705 1530 27715 1550
rect 27675 1515 27715 1530
rect 27730 1650 27770 1665
rect 27730 1630 27740 1650
rect 27760 1630 27770 1650
rect 27730 1600 27770 1630
rect 27730 1580 27740 1600
rect 27760 1580 27770 1600
rect 27730 1550 27770 1580
rect 27730 1530 27740 1550
rect 27760 1530 27770 1550
rect 27730 1515 27770 1530
rect 25605 1320 25615 1340
rect 25635 1320 25645 1340
rect 25605 1290 25645 1320
rect 25605 1270 25615 1290
rect 25635 1270 25645 1290
rect 25605 1240 25645 1270
rect 25605 1220 25615 1240
rect 25635 1220 25645 1240
rect 25605 1190 25645 1220
rect 25605 1170 25615 1190
rect 25635 1170 25645 1190
rect 25605 1140 25645 1170
rect 25605 1120 25615 1140
rect 25635 1120 25645 1140
rect 25605 1090 25645 1120
rect 25605 1070 25615 1090
rect 25635 1070 25645 1090
rect 25605 1040 25645 1070
rect 25605 1020 25615 1040
rect 25635 1020 25645 1040
rect 25605 990 25645 1020
rect 25605 970 25615 990
rect 25635 970 25645 990
rect 25605 955 25645 970
rect 2995 865 3035 880
rect 2995 845 3005 865
rect 3025 845 3035 865
rect 2995 815 3035 845
rect 2995 795 3005 815
rect 3025 795 3035 815
rect 2995 780 3035 795
rect 3085 865 3125 880
rect 3085 845 3095 865
rect 3115 845 3125 865
rect 3085 815 3125 845
rect 3085 795 3095 815
rect 3115 795 3125 815
rect 3085 780 3125 795
rect 3175 865 3215 880
rect 3175 845 3185 865
rect 3205 845 3215 865
rect 3175 815 3215 845
rect 3175 795 3185 815
rect 3205 795 3215 815
rect 3175 780 3215 795
rect 3265 865 3305 880
rect 3265 845 3275 865
rect 3295 845 3305 865
rect 3265 815 3305 845
rect 3265 795 3275 815
rect 3295 795 3305 815
rect 3265 780 3305 795
rect 3355 865 3395 880
rect 3355 845 3365 865
rect 3385 845 3395 865
rect 3355 815 3395 845
rect 3355 795 3365 815
rect 3385 795 3395 815
rect 3355 780 3395 795
rect 3445 865 3485 880
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 815 3485 845
rect 3445 795 3455 815
rect 3475 795 3485 815
rect 3445 780 3485 795
rect 3535 865 3575 880
rect 3535 845 3545 865
rect 3565 845 3575 865
rect 3535 815 3575 845
rect 3535 795 3545 815
rect 3565 795 3575 815
rect 3535 780 3575 795
rect 3625 865 3665 880
rect 3625 845 3635 865
rect 3655 845 3665 865
rect 3625 815 3665 845
rect 3625 795 3635 815
rect 3655 795 3665 815
rect 3625 780 3665 795
rect 3715 865 3755 880
rect 3715 845 3725 865
rect 3745 845 3755 865
rect 3715 815 3755 845
rect 3715 795 3725 815
rect 3745 795 3755 815
rect 3715 780 3755 795
rect 3805 865 3845 880
rect 3805 845 3815 865
rect 3835 845 3845 865
rect 3805 815 3845 845
rect 3805 795 3815 815
rect 3835 795 3845 815
rect 3805 780 3845 795
rect 3895 865 3935 880
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 815 3935 845
rect 3895 795 3905 815
rect 3925 795 3935 815
rect 3895 780 3935 795
rect 3985 865 4025 880
rect 3985 845 3995 865
rect 4015 845 4025 865
rect 3985 815 4025 845
rect 3985 795 3995 815
rect 4015 795 4025 815
rect 3985 780 4025 795
rect 4075 865 4115 880
rect 4075 845 4085 865
rect 4105 845 4115 865
rect 4075 815 4115 845
rect 4075 795 4085 815
rect 4105 795 4115 815
rect 4075 780 4115 795
rect 4165 865 4205 880
rect 4165 845 4175 865
rect 4195 845 4205 865
rect 4165 815 4205 845
rect 4165 795 4175 815
rect 4195 795 4205 815
rect 4165 780 4205 795
rect 4255 865 4295 880
rect 4255 845 4265 865
rect 4285 845 4295 865
rect 4255 815 4295 845
rect 4255 795 4265 815
rect 4285 795 4295 815
rect 4255 780 4295 795
rect 4345 865 4385 880
rect 4345 845 4355 865
rect 4375 845 4385 865
rect 4345 815 4385 845
rect 4345 795 4355 815
rect 4375 795 4385 815
rect 4345 780 4385 795
rect 4435 865 4475 880
rect 4435 845 4445 865
rect 4465 845 4475 865
rect 4435 815 4475 845
rect 4435 795 4445 815
rect 4465 795 4475 815
rect 4435 780 4475 795
rect 4525 865 4565 880
rect 4525 845 4535 865
rect 4555 845 4565 865
rect 4525 815 4565 845
rect 4525 795 4535 815
rect 4555 795 4565 815
rect 4525 780 4565 795
rect 4615 865 4655 880
rect 4615 845 4625 865
rect 4645 845 4655 865
rect 4615 815 4655 845
rect 4615 795 4625 815
rect 4645 795 4655 815
rect 4615 780 4655 795
rect 4705 865 4745 880
rect 4705 845 4715 865
rect 4735 845 4745 865
rect 4705 815 4745 845
rect 4705 795 4715 815
rect 4735 795 4745 815
rect 4705 780 4745 795
rect 4795 865 4835 880
rect 4795 845 4805 865
rect 4825 845 4835 865
rect 4795 815 4835 845
rect 4795 795 4805 815
rect 4825 795 4835 815
rect 4795 780 4835 795
rect 4885 865 4925 880
rect 4885 845 4895 865
rect 4915 845 4925 865
rect 4885 815 4925 845
rect 4885 795 4895 815
rect 4915 795 4925 815
rect 4885 780 4925 795
rect 4975 865 5015 880
rect 4975 845 4985 865
rect 5005 845 5015 865
rect 4975 815 5015 845
rect 4975 795 4985 815
rect 5005 795 5015 815
rect 4975 780 5015 795
rect 26205 1070 26245 1085
rect 26205 1050 26215 1070
rect 26235 1050 26245 1070
rect 26205 1020 26245 1050
rect 26205 1000 26215 1020
rect 26235 1000 26245 1020
rect 26205 970 26245 1000
rect 26205 950 26215 970
rect 26235 950 26245 970
rect 26205 920 26245 950
rect 26205 900 26215 920
rect 26235 900 26245 920
rect 26205 870 26245 900
rect 26205 850 26215 870
rect 26235 850 26245 870
rect 26205 835 26245 850
rect 26260 1070 26300 1085
rect 26260 1050 26270 1070
rect 26290 1050 26300 1070
rect 26260 1020 26300 1050
rect 26260 1000 26270 1020
rect 26290 1000 26300 1020
rect 26260 970 26300 1000
rect 26260 950 26270 970
rect 26290 950 26300 970
rect 26260 920 26300 950
rect 26260 900 26270 920
rect 26290 900 26300 920
rect 26260 870 26300 900
rect 26260 850 26270 870
rect 26290 850 26300 870
rect 26260 835 26300 850
rect 26315 1070 26355 1085
rect 26315 1050 26325 1070
rect 26345 1050 26355 1070
rect 26315 1020 26355 1050
rect 26315 1000 26325 1020
rect 26345 1000 26355 1020
rect 26315 970 26355 1000
rect 26315 950 26325 970
rect 26345 950 26355 970
rect 26315 920 26355 950
rect 26315 900 26325 920
rect 26345 900 26355 920
rect 26315 870 26355 900
rect 26315 850 26325 870
rect 26345 850 26355 870
rect 26315 835 26355 850
rect 26370 1070 26410 1085
rect 26370 1050 26380 1070
rect 26400 1050 26410 1070
rect 26370 1020 26410 1050
rect 26370 1000 26380 1020
rect 26400 1000 26410 1020
rect 26370 970 26410 1000
rect 26370 950 26380 970
rect 26400 950 26410 970
rect 26370 920 26410 950
rect 26370 900 26380 920
rect 26400 900 26410 920
rect 26370 870 26410 900
rect 26370 850 26380 870
rect 26400 850 26410 870
rect 26370 835 26410 850
rect 26425 1070 26465 1085
rect 26425 1050 26435 1070
rect 26455 1050 26465 1070
rect 26425 1020 26465 1050
rect 26425 1000 26435 1020
rect 26455 1000 26465 1020
rect 26425 970 26465 1000
rect 26425 950 26435 970
rect 26455 950 26465 970
rect 26425 920 26465 950
rect 26425 900 26435 920
rect 26455 900 26465 920
rect 26425 870 26465 900
rect 26425 850 26435 870
rect 26455 850 26465 870
rect 26425 835 26465 850
rect 26480 1070 26520 1085
rect 26480 1050 26490 1070
rect 26510 1050 26520 1070
rect 26480 1020 26520 1050
rect 26480 1000 26490 1020
rect 26510 1000 26520 1020
rect 26480 970 26520 1000
rect 26480 950 26490 970
rect 26510 950 26520 970
rect 26480 920 26520 950
rect 26480 900 26490 920
rect 26510 900 26520 920
rect 26480 870 26520 900
rect 26480 850 26490 870
rect 26510 850 26520 870
rect 26480 835 26520 850
rect 26535 1070 26575 1085
rect 26535 1050 26545 1070
rect 26565 1050 26575 1070
rect 26535 1020 26575 1050
rect 26535 1000 26545 1020
rect 26565 1000 26575 1020
rect 26535 970 26575 1000
rect 26535 950 26545 970
rect 26565 950 26575 970
rect 26535 920 26575 950
rect 26535 900 26545 920
rect 26565 900 26575 920
rect 26535 870 26575 900
rect 26535 850 26545 870
rect 26565 850 26575 870
rect 26535 835 26575 850
rect 26590 1070 26630 1085
rect 26590 1050 26600 1070
rect 26620 1050 26630 1070
rect 26590 1020 26630 1050
rect 26590 1000 26600 1020
rect 26620 1000 26630 1020
rect 26590 970 26630 1000
rect 26590 950 26600 970
rect 26620 950 26630 970
rect 26590 920 26630 950
rect 26590 900 26600 920
rect 26620 900 26630 920
rect 26590 870 26630 900
rect 26590 850 26600 870
rect 26620 850 26630 870
rect 26590 835 26630 850
rect 26645 1070 26685 1085
rect 26645 1050 26655 1070
rect 26675 1050 26685 1070
rect 26645 1020 26685 1050
rect 26645 1000 26655 1020
rect 26675 1000 26685 1020
rect 26645 970 26685 1000
rect 26645 950 26655 970
rect 26675 950 26685 970
rect 26645 920 26685 950
rect 26645 900 26655 920
rect 26675 900 26685 920
rect 26645 870 26685 900
rect 26645 850 26655 870
rect 26675 850 26685 870
rect 26645 835 26685 850
rect 26700 1070 26740 1085
rect 26700 1050 26710 1070
rect 26730 1050 26740 1070
rect 26700 1020 26740 1050
rect 26700 1000 26710 1020
rect 26730 1000 26740 1020
rect 26700 970 26740 1000
rect 26700 950 26710 970
rect 26730 950 26740 970
rect 26700 920 26740 950
rect 26700 900 26710 920
rect 26730 900 26740 920
rect 26700 870 26740 900
rect 26700 850 26710 870
rect 26730 850 26740 870
rect 26700 835 26740 850
rect 26755 1070 26795 1085
rect 26755 1050 26765 1070
rect 26785 1050 26795 1070
rect 26755 1020 26795 1050
rect 26755 1000 26765 1020
rect 26785 1000 26795 1020
rect 26755 970 26795 1000
rect 26755 950 26765 970
rect 26785 950 26795 970
rect 26755 920 26795 950
rect 26755 900 26765 920
rect 26785 900 26795 920
rect 26755 870 26795 900
rect 26755 850 26765 870
rect 26785 850 26795 870
rect 26755 835 26795 850
rect 26810 1070 26850 1085
rect 26810 1050 26820 1070
rect 26840 1050 26850 1070
rect 26810 1020 26850 1050
rect 26810 1000 26820 1020
rect 26840 1000 26850 1020
rect 26810 970 26850 1000
rect 26810 950 26820 970
rect 26840 950 26850 970
rect 26810 920 26850 950
rect 26810 900 26820 920
rect 26840 900 26850 920
rect 26810 870 26850 900
rect 26810 850 26820 870
rect 26840 850 26850 870
rect 26810 835 26850 850
rect 26865 1070 26905 1085
rect 26865 1050 26875 1070
rect 26895 1050 26905 1070
rect 26865 1020 26905 1050
rect 26865 1000 26875 1020
rect 26895 1000 26905 1020
rect 26865 970 26905 1000
rect 26865 950 26875 970
rect 26895 950 26905 970
rect 26865 920 26905 950
rect 26865 900 26875 920
rect 26895 900 26905 920
rect 26865 870 26905 900
rect 26865 850 26875 870
rect 26895 850 26905 870
rect 26865 835 26905 850
rect 26920 1070 26960 1085
rect 26920 1050 26930 1070
rect 26950 1050 26960 1070
rect 26920 1020 26960 1050
rect 26920 1000 26930 1020
rect 26950 1000 26960 1020
rect 26920 970 26960 1000
rect 26920 950 26930 970
rect 26950 950 26960 970
rect 26920 920 26960 950
rect 26920 900 26930 920
rect 26950 900 26960 920
rect 26920 870 26960 900
rect 26920 850 26930 870
rect 26950 850 26960 870
rect 26920 835 26960 850
rect 26975 1070 27015 1085
rect 26975 1050 26985 1070
rect 27005 1050 27015 1070
rect 26975 1020 27015 1050
rect 26975 1000 26985 1020
rect 27005 1000 27015 1020
rect 26975 970 27015 1000
rect 26975 950 26985 970
rect 27005 950 27015 970
rect 26975 920 27015 950
rect 26975 900 26985 920
rect 27005 900 27015 920
rect 26975 870 27015 900
rect 26975 850 26985 870
rect 27005 850 27015 870
rect 26975 835 27015 850
rect 27030 1070 27070 1085
rect 27030 1050 27040 1070
rect 27060 1050 27070 1070
rect 27030 1020 27070 1050
rect 27030 1000 27040 1020
rect 27060 1000 27070 1020
rect 27030 970 27070 1000
rect 27030 950 27040 970
rect 27060 950 27070 970
rect 27030 920 27070 950
rect 27030 900 27040 920
rect 27060 900 27070 920
rect 27030 870 27070 900
rect 27030 850 27040 870
rect 27060 850 27070 870
rect 27030 835 27070 850
rect 27085 1070 27125 1085
rect 27085 1050 27095 1070
rect 27115 1050 27125 1070
rect 27085 1020 27125 1050
rect 27085 1000 27095 1020
rect 27115 1000 27125 1020
rect 27085 970 27125 1000
rect 27085 950 27095 970
rect 27115 950 27125 970
rect 27085 920 27125 950
rect 27085 900 27095 920
rect 27115 900 27125 920
rect 27085 870 27125 900
rect 27085 850 27095 870
rect 27115 850 27125 870
rect 27085 835 27125 850
rect 27140 1070 27180 1085
rect 27140 1050 27150 1070
rect 27170 1050 27180 1070
rect 27140 1020 27180 1050
rect 27140 1000 27150 1020
rect 27170 1000 27180 1020
rect 27140 970 27180 1000
rect 27140 950 27150 970
rect 27170 950 27180 970
rect 27140 920 27180 950
rect 27140 900 27150 920
rect 27170 900 27180 920
rect 27140 870 27180 900
rect 27140 850 27150 870
rect 27170 850 27180 870
rect 27140 835 27180 850
rect 27195 1070 27235 1085
rect 27195 1050 27205 1070
rect 27225 1050 27235 1070
rect 27195 1020 27235 1050
rect 27195 1000 27205 1020
rect 27225 1000 27235 1020
rect 27195 970 27235 1000
rect 27195 950 27205 970
rect 27225 950 27235 970
rect 27195 920 27235 950
rect 27195 900 27205 920
rect 27225 900 27235 920
rect 27195 870 27235 900
rect 27195 850 27205 870
rect 27225 850 27235 870
rect 27195 835 27235 850
rect 27250 1070 27290 1085
rect 27250 1050 27260 1070
rect 27280 1050 27290 1070
rect 27250 1020 27290 1050
rect 27250 1000 27260 1020
rect 27280 1000 27290 1020
rect 27250 970 27290 1000
rect 27250 950 27260 970
rect 27280 950 27290 970
rect 27250 920 27290 950
rect 27250 900 27260 920
rect 27280 900 27290 920
rect 27250 870 27290 900
rect 27250 850 27260 870
rect 27280 850 27290 870
rect 27250 835 27290 850
rect 27305 1070 27345 1085
rect 27305 1050 27315 1070
rect 27335 1050 27345 1070
rect 27305 1020 27345 1050
rect 27305 1000 27315 1020
rect 27335 1000 27345 1020
rect 27305 970 27345 1000
rect 27305 950 27315 970
rect 27335 950 27345 970
rect 27305 920 27345 950
rect 27305 900 27315 920
rect 27335 900 27345 920
rect 27305 870 27345 900
rect 27305 850 27315 870
rect 27335 850 27345 870
rect 27305 835 27345 850
rect 27360 1070 27400 1085
rect 27360 1050 27370 1070
rect 27390 1050 27400 1070
rect 27360 1020 27400 1050
rect 27360 1000 27370 1020
rect 27390 1000 27400 1020
rect 27360 970 27400 1000
rect 27360 950 27370 970
rect 27390 950 27400 970
rect 27360 920 27400 950
rect 27360 900 27370 920
rect 27390 900 27400 920
rect 27360 870 27400 900
rect 27360 850 27370 870
rect 27390 850 27400 870
rect 27360 835 27400 850
rect 27415 1070 27455 1085
rect 27415 1050 27425 1070
rect 27445 1050 27455 1070
rect 27415 1020 27455 1050
rect 27415 1000 27425 1020
rect 27445 1000 27455 1020
rect 27415 970 27455 1000
rect 27415 950 27425 970
rect 27445 950 27455 970
rect 27415 920 27455 950
rect 27415 900 27425 920
rect 27445 900 27455 920
rect 27415 870 27455 900
rect 27415 850 27425 870
rect 27445 850 27455 870
rect 27415 835 27455 850
rect 27470 1070 27510 1085
rect 27470 1050 27480 1070
rect 27500 1050 27510 1070
rect 27470 1020 27510 1050
rect 27470 1000 27480 1020
rect 27500 1000 27510 1020
rect 27470 970 27510 1000
rect 27470 950 27480 970
rect 27500 950 27510 970
rect 27470 920 27510 950
rect 27470 900 27480 920
rect 27500 900 27510 920
rect 27470 870 27510 900
rect 27470 850 27480 870
rect 27500 850 27510 870
rect 27470 835 27510 850
rect 27525 1070 27565 1085
rect 27525 1050 27535 1070
rect 27555 1050 27565 1070
rect 27525 1020 27565 1050
rect 27525 1000 27535 1020
rect 27555 1000 27565 1020
rect 27525 970 27565 1000
rect 27525 950 27535 970
rect 27555 950 27565 970
rect 27525 920 27565 950
rect 27525 900 27535 920
rect 27555 900 27565 920
rect 27525 870 27565 900
rect 27525 850 27535 870
rect 27555 850 27565 870
rect 27525 835 27565 850
rect 27580 1070 27620 1085
rect 27580 1050 27590 1070
rect 27610 1050 27620 1070
rect 27580 1020 27620 1050
rect 27580 1000 27590 1020
rect 27610 1000 27620 1020
rect 27580 970 27620 1000
rect 27580 950 27590 970
rect 27610 950 27620 970
rect 27580 920 27620 950
rect 27580 900 27590 920
rect 27610 900 27620 920
rect 27580 870 27620 900
rect 27580 850 27590 870
rect 27610 850 27620 870
rect 27580 835 27620 850
rect 28205 1640 28245 1655
rect 28205 1620 28215 1640
rect 28235 1620 28245 1640
rect 28205 1590 28245 1620
rect 28205 1570 28215 1590
rect 28235 1570 28245 1590
rect 28205 1540 28245 1570
rect 28205 1520 28215 1540
rect 28235 1520 28245 1540
rect 28205 1490 28245 1520
rect 28205 1470 28215 1490
rect 28235 1470 28245 1490
rect 28205 1440 28245 1470
rect 28205 1420 28215 1440
rect 28235 1420 28245 1440
rect 28205 1390 28245 1420
rect 28205 1370 28215 1390
rect 28235 1370 28245 1390
rect 28205 1340 28245 1370
rect 28205 1320 28215 1340
rect 28235 1320 28245 1340
rect 28205 1290 28245 1320
rect 28205 1270 28215 1290
rect 28235 1270 28245 1290
rect 28205 1240 28245 1270
rect 28205 1220 28215 1240
rect 28235 1220 28245 1240
rect 28205 1190 28245 1220
rect 28205 1170 28215 1190
rect 28235 1170 28245 1190
rect 28205 1140 28245 1170
rect 28205 1120 28215 1140
rect 28235 1120 28245 1140
rect 28205 1090 28245 1120
rect 28205 1070 28215 1090
rect 28235 1070 28245 1090
rect 28205 1040 28245 1070
rect 28205 1020 28215 1040
rect 28235 1020 28245 1040
rect 28205 990 28245 1020
rect 28205 970 28215 990
rect 28235 970 28245 990
rect 28205 955 28245 970
rect 28305 1640 28345 1655
rect 28305 1620 28315 1640
rect 28335 1620 28345 1640
rect 28305 1590 28345 1620
rect 28305 1570 28315 1590
rect 28335 1570 28345 1590
rect 28305 1540 28345 1570
rect 28305 1520 28315 1540
rect 28335 1520 28345 1540
rect 28305 1490 28345 1520
rect 28305 1470 28315 1490
rect 28335 1470 28345 1490
rect 28305 1440 28345 1470
rect 28305 1420 28315 1440
rect 28335 1420 28345 1440
rect 28305 1390 28345 1420
rect 28305 1370 28315 1390
rect 28335 1370 28345 1390
rect 28305 1340 28345 1370
rect 28305 1320 28315 1340
rect 28335 1320 28345 1340
rect 28305 1290 28345 1320
rect 28305 1270 28315 1290
rect 28335 1270 28345 1290
rect 28305 1240 28345 1270
rect 28305 1220 28315 1240
rect 28335 1220 28345 1240
rect 28305 1190 28345 1220
rect 28305 1170 28315 1190
rect 28335 1170 28345 1190
rect 28305 1140 28345 1170
rect 28305 1120 28315 1140
rect 28335 1120 28345 1140
rect 28305 1090 28345 1120
rect 28305 1070 28315 1090
rect 28335 1070 28345 1090
rect 28305 1040 28345 1070
rect 28305 1020 28315 1040
rect 28335 1020 28345 1040
rect 28305 990 28345 1020
rect 28305 970 28315 990
rect 28335 970 28345 990
rect 28305 955 28345 970
rect 28405 1640 28445 1655
rect 28405 1620 28415 1640
rect 28435 1620 28445 1640
rect 28405 1590 28445 1620
rect 28405 1570 28415 1590
rect 28435 1570 28445 1590
rect 28405 1540 28445 1570
rect 28405 1520 28415 1540
rect 28435 1520 28445 1540
rect 28405 1490 28445 1520
rect 28405 1470 28415 1490
rect 28435 1470 28445 1490
rect 28405 1440 28445 1470
rect 28405 1420 28415 1440
rect 28435 1420 28445 1440
rect 28405 1390 28445 1420
rect 28405 1370 28415 1390
rect 28435 1370 28445 1390
rect 28405 1340 28445 1370
rect 28405 1320 28415 1340
rect 28435 1320 28445 1340
rect 28405 1290 28445 1320
rect 28405 1270 28415 1290
rect 28435 1270 28445 1290
rect 28405 1240 28445 1270
rect 28405 1220 28415 1240
rect 28435 1220 28445 1240
rect 28405 1190 28445 1220
rect 28405 1170 28415 1190
rect 28435 1170 28445 1190
rect 28405 1140 28445 1170
rect 28405 1120 28415 1140
rect 28435 1120 28445 1140
rect 28405 1090 28445 1120
rect 28405 1070 28415 1090
rect 28435 1070 28445 1090
rect 28405 1040 28445 1070
rect 28405 1020 28415 1040
rect 28435 1020 28445 1040
rect 28405 990 28445 1020
rect 28405 970 28415 990
rect 28435 970 28445 990
rect 28405 955 28445 970
rect 28505 1640 28545 1655
rect 28505 1620 28515 1640
rect 28535 1620 28545 1640
rect 28505 1590 28545 1620
rect 28505 1570 28515 1590
rect 28535 1570 28545 1590
rect 28505 1540 28545 1570
rect 28505 1520 28515 1540
rect 28535 1520 28545 1540
rect 28505 1490 28545 1520
rect 28505 1470 28515 1490
rect 28535 1470 28545 1490
rect 28505 1440 28545 1470
rect 28505 1420 28515 1440
rect 28535 1420 28545 1440
rect 28505 1390 28545 1420
rect 28505 1370 28515 1390
rect 28535 1370 28545 1390
rect 28505 1340 28545 1370
rect 28505 1320 28515 1340
rect 28535 1320 28545 1340
rect 28505 1290 28545 1320
rect 28505 1270 28515 1290
rect 28535 1270 28545 1290
rect 28505 1240 28545 1270
rect 28505 1220 28515 1240
rect 28535 1220 28545 1240
rect 28505 1190 28545 1220
rect 28505 1170 28515 1190
rect 28535 1170 28545 1190
rect 28505 1140 28545 1170
rect 28505 1120 28515 1140
rect 28535 1120 28545 1140
rect 28505 1090 28545 1120
rect 28505 1070 28515 1090
rect 28535 1070 28545 1090
rect 28505 1040 28545 1070
rect 28505 1020 28515 1040
rect 28535 1020 28545 1040
rect 28505 990 28545 1020
rect 28505 970 28515 990
rect 28535 970 28545 990
rect 28505 955 28545 970
rect 28605 1640 28645 1655
rect 28605 1620 28615 1640
rect 28635 1620 28645 1640
rect 28605 1590 28645 1620
rect 28605 1570 28615 1590
rect 28635 1570 28645 1590
rect 28605 1540 28645 1570
rect 28605 1520 28615 1540
rect 28635 1520 28645 1540
rect 28605 1490 28645 1520
rect 28605 1470 28615 1490
rect 28635 1470 28645 1490
rect 28605 1440 28645 1470
rect 28605 1420 28615 1440
rect 28635 1420 28645 1440
rect 28605 1390 28645 1420
rect 28605 1370 28615 1390
rect 28635 1370 28645 1390
rect 28605 1340 28645 1370
rect 28605 1320 28615 1340
rect 28635 1320 28645 1340
rect 28605 1290 28645 1320
rect 28605 1270 28615 1290
rect 28635 1270 28645 1290
rect 28605 1240 28645 1270
rect 28605 1220 28615 1240
rect 28635 1220 28645 1240
rect 28605 1190 28645 1220
rect 28605 1170 28615 1190
rect 28635 1170 28645 1190
rect 28605 1140 28645 1170
rect 28605 1120 28615 1140
rect 28635 1120 28645 1140
rect 28605 1090 28645 1120
rect 28605 1070 28615 1090
rect 28635 1070 28645 1090
rect 28605 1040 28645 1070
rect 28605 1020 28615 1040
rect 28635 1020 28645 1040
rect 28605 990 28645 1020
rect 28605 970 28615 990
rect 28635 970 28645 990
rect 28605 955 28645 970
rect 28705 1640 28745 1655
rect 28705 1620 28715 1640
rect 28735 1620 28745 1640
rect 28705 1590 28745 1620
rect 28705 1570 28715 1590
rect 28735 1570 28745 1590
rect 28705 1540 28745 1570
rect 28705 1520 28715 1540
rect 28735 1520 28745 1540
rect 28705 1490 28745 1520
rect 28705 1470 28715 1490
rect 28735 1470 28745 1490
rect 28705 1440 28745 1470
rect 28705 1420 28715 1440
rect 28735 1420 28745 1440
rect 28705 1390 28745 1420
rect 28705 1370 28715 1390
rect 28735 1370 28745 1390
rect 28705 1340 28745 1370
rect 28705 1320 28715 1340
rect 28735 1320 28745 1340
rect 28705 1290 28745 1320
rect 28705 1270 28715 1290
rect 28735 1270 28745 1290
rect 28705 1240 28745 1270
rect 28705 1220 28715 1240
rect 28735 1220 28745 1240
rect 28705 1190 28745 1220
rect 28705 1170 28715 1190
rect 28735 1170 28745 1190
rect 28705 1140 28745 1170
rect 28705 1120 28715 1140
rect 28735 1120 28745 1140
rect 28705 1090 28745 1120
rect 28705 1070 28715 1090
rect 28735 1070 28745 1090
rect 28705 1040 28745 1070
rect 28705 1020 28715 1040
rect 28735 1020 28745 1040
rect 28705 990 28745 1020
rect 28705 970 28715 990
rect 28735 970 28745 990
rect 28705 955 28745 970
rect 28805 1640 28845 1655
rect 28805 1620 28815 1640
rect 28835 1620 28845 1640
rect 28805 1590 28845 1620
rect 28805 1570 28815 1590
rect 28835 1570 28845 1590
rect 28805 1540 28845 1570
rect 28805 1520 28815 1540
rect 28835 1520 28845 1540
rect 28805 1490 28845 1520
rect 28805 1470 28815 1490
rect 28835 1470 28845 1490
rect 28805 1440 28845 1470
rect 28805 1420 28815 1440
rect 28835 1420 28845 1440
rect 28805 1390 28845 1420
rect 28805 1370 28815 1390
rect 28835 1370 28845 1390
rect 28805 1340 28845 1370
rect 28805 1320 28815 1340
rect 28835 1320 28845 1340
rect 28805 1290 28845 1320
rect 28805 1270 28815 1290
rect 28835 1270 28845 1290
rect 28805 1240 28845 1270
rect 28805 1220 28815 1240
rect 28835 1220 28845 1240
rect 28805 1190 28845 1220
rect 28805 1170 28815 1190
rect 28835 1170 28845 1190
rect 28805 1140 28845 1170
rect 28805 1120 28815 1140
rect 28835 1120 28845 1140
rect 28805 1090 28845 1120
rect 28805 1070 28815 1090
rect 28835 1070 28845 1090
rect 28805 1040 28845 1070
rect 28805 1020 28815 1040
rect 28835 1020 28845 1040
rect 28805 990 28845 1020
rect 28805 970 28815 990
rect 28835 970 28845 990
rect 28805 955 28845 970
rect 16260 735 16300 750
rect 16260 715 16270 735
rect 16290 715 16300 735
rect 16260 685 16300 715
rect 16260 665 16270 685
rect 16290 665 16300 685
rect 16260 650 16300 665
rect 16490 735 16530 750
rect 16490 715 16500 735
rect 16520 715 16530 735
rect 16490 685 16530 715
rect 16880 735 16920 750
rect 16880 715 16890 735
rect 16910 715 16920 735
rect 16880 700 16920 715
rect 16935 735 16975 750
rect 16935 715 16945 735
rect 16965 715 16975 735
rect 16935 700 16975 715
rect 16990 735 17030 750
rect 16990 715 17000 735
rect 17020 715 17030 735
rect 16990 700 17030 715
rect 17045 735 17085 750
rect 17045 715 17055 735
rect 17075 715 17085 735
rect 17045 700 17085 715
rect 17100 735 17140 750
rect 17100 715 17110 735
rect 17130 715 17140 735
rect 17100 700 17140 715
rect 17155 735 17195 750
rect 17155 715 17165 735
rect 17185 715 17195 735
rect 17155 700 17195 715
rect 17210 735 17250 750
rect 17210 715 17220 735
rect 17240 715 17250 735
rect 17210 700 17250 715
rect 17265 735 17305 750
rect 17265 715 17275 735
rect 17295 715 17305 735
rect 17265 700 17305 715
rect 17320 735 17360 750
rect 17320 715 17330 735
rect 17350 715 17360 735
rect 17320 700 17360 715
rect 17375 735 17415 750
rect 17375 715 17385 735
rect 17405 715 17415 735
rect 17375 700 17415 715
rect 17430 735 17470 750
rect 17430 715 17440 735
rect 17460 715 17470 735
rect 17430 700 17470 715
rect 17485 735 17525 750
rect 17485 715 17495 735
rect 17515 715 17525 735
rect 17485 700 17525 715
rect 17540 735 17580 750
rect 17540 715 17550 735
rect 17570 715 17580 735
rect 17540 700 17580 715
rect 16490 665 16500 685
rect 16520 665 16530 685
rect 16490 650 16530 665
rect 26260 535 26300 550
rect 26260 515 26270 535
rect 26290 515 26300 535
rect 26260 485 26300 515
rect 26260 465 26270 485
rect 26290 465 26300 485
rect 26260 450 26300 465
rect 26490 535 26530 550
rect 26490 515 26500 535
rect 26520 515 26530 535
rect 26490 485 26530 515
rect 26490 465 26500 485
rect 26520 465 26530 485
rect 26490 450 26530 465
rect 26880 535 26920 550
rect 26880 515 26890 535
rect 26910 515 26920 535
rect 26880 500 26920 515
rect 26935 535 26975 550
rect 26935 515 26945 535
rect 26965 515 26975 535
rect 26935 500 26975 515
rect 26990 535 27030 550
rect 26990 515 27000 535
rect 27020 515 27030 535
rect 26990 500 27030 515
rect 27045 535 27085 550
rect 27045 515 27055 535
rect 27075 515 27085 535
rect 27045 500 27085 515
rect 27100 535 27140 550
rect 27100 515 27110 535
rect 27130 515 27140 535
rect 27100 500 27140 515
rect 27155 535 27195 550
rect 27155 515 27165 535
rect 27185 515 27195 535
rect 27155 500 27195 515
rect 27210 535 27250 550
rect 27210 515 27220 535
rect 27240 515 27250 535
rect 27210 500 27250 515
rect 27265 535 27305 550
rect 27265 515 27275 535
rect 27295 515 27305 535
rect 27265 500 27305 515
rect 27320 535 27360 550
rect 27320 515 27330 535
rect 27350 515 27360 535
rect 27320 500 27360 515
rect 27375 535 27415 550
rect 27375 515 27385 535
rect 27405 515 27415 535
rect 27375 500 27415 515
rect 27430 535 27470 550
rect 27430 515 27440 535
rect 27460 515 27470 535
rect 27430 500 27470 515
rect 27485 535 27525 550
rect 27485 515 27495 535
rect 27515 515 27525 535
rect 27485 500 27525 515
rect 27540 535 27580 550
rect 27540 515 27550 535
rect 27570 515 27580 535
rect 27540 500 27580 515
<< pdiff >>
rect 26255 4830 26295 4858
rect 26255 4810 26265 4830
rect 26285 4810 26295 4830
rect 26255 4795 26295 4810
rect 26315 4835 26355 4858
rect 26315 4815 26325 4835
rect 26345 4815 26355 4835
rect 26315 4795 26355 4815
rect 26375 4835 26415 4858
rect 26375 4815 26385 4835
rect 26405 4815 26415 4835
rect 26375 4795 26415 4815
rect 26435 4830 26475 4858
rect 26435 4810 26445 4830
rect 26465 4810 26475 4830
rect 26435 4795 26475 4810
rect 26505 4845 26545 4875
rect 26505 4825 26515 4845
rect 26535 4825 26545 4845
rect 26505 4795 26545 4825
rect 26565 4845 26605 4875
rect 26565 4825 26575 4845
rect 26595 4825 26605 4845
rect 26565 4795 26605 4825
rect 26625 4845 26665 4875
rect 26625 4825 26635 4845
rect 26655 4825 26665 4845
rect 26625 4795 26665 4825
rect 26685 4845 26725 4875
rect 26685 4825 26695 4845
rect 26715 4825 26725 4845
rect 26685 4795 26725 4825
rect 26745 4845 26785 4875
rect 26745 4825 26755 4845
rect 26775 4825 26785 4845
rect 26745 4795 26785 4825
rect 26805 4845 26845 4875
rect 26805 4825 26815 4845
rect 26835 4825 26845 4845
rect 26805 4795 26845 4825
rect 26865 4845 26905 4875
rect 26865 4825 26875 4845
rect 26895 4825 26905 4845
rect 26865 4795 26905 4825
rect 27235 4830 27275 4850
rect 27235 4810 27245 4830
rect 27265 4810 27275 4830
rect 27235 4790 27275 4810
rect 27295 4830 27335 4850
rect 27295 4810 27305 4830
rect 27325 4810 27335 4830
rect 27295 4790 27335 4810
rect 27355 4830 27395 4850
rect 27355 4810 27365 4830
rect 27385 4810 27395 4830
rect 27355 4790 27395 4810
rect 27415 4830 27455 4850
rect 27415 4810 27425 4830
rect 27445 4810 27455 4830
rect 27415 4790 27455 4810
rect 27475 4830 27515 4850
rect 27475 4810 27485 4830
rect 27505 4810 27515 4830
rect 27475 4790 27515 4810
rect 27535 4830 27575 4850
rect 27535 4810 27545 4830
rect 27565 4810 27575 4830
rect 27535 4790 27575 4810
rect 27595 4830 27635 4850
rect 27595 4810 27605 4830
rect 27625 4810 27635 4830
rect 27595 4790 27635 4810
rect 27655 4830 27695 4850
rect 27655 4810 27665 4830
rect 27685 4810 27695 4830
rect 27655 4790 27695 4810
rect 27715 4830 27755 4850
rect 27715 4810 27725 4830
rect 27745 4810 27755 4830
rect 27715 4790 27755 4810
rect 16205 4325 16245 4353
rect 16205 4305 16215 4325
rect 16235 4305 16245 4325
rect 16205 4290 16245 4305
rect 16265 4330 16305 4353
rect 16265 4310 16275 4330
rect 16295 4310 16305 4330
rect 16265 4290 16305 4310
rect 16325 4330 16365 4353
rect 16325 4310 16335 4330
rect 16355 4310 16365 4330
rect 16325 4290 16365 4310
rect 16385 4325 16425 4353
rect 16385 4305 16395 4325
rect 16415 4305 16425 4325
rect 16385 4290 16425 4305
rect 16535 4340 16575 4370
rect 16535 4320 16545 4340
rect 16565 4320 16575 4340
rect 16535 4290 16575 4320
rect 16595 4340 16635 4370
rect 16595 4320 16605 4340
rect 16625 4320 16635 4340
rect 16595 4290 16635 4320
rect 16655 4340 16695 4370
rect 16655 4320 16665 4340
rect 16685 4320 16695 4340
rect 16655 4290 16695 4320
rect 16715 4340 16755 4370
rect 16715 4320 16725 4340
rect 16745 4320 16755 4340
rect 16715 4290 16755 4320
rect 16775 4340 16815 4370
rect 16775 4320 16785 4340
rect 16805 4320 16815 4340
rect 16775 4290 16815 4320
rect 16835 4340 16875 4370
rect 16835 4320 16845 4340
rect 16865 4320 16875 4340
rect 16835 4290 16875 4320
rect 16895 4340 16935 4370
rect 26250 4415 26290 4430
rect 26250 4395 26260 4415
rect 26280 4395 26290 4415
rect 26250 4380 26290 4395
rect 26305 4415 26345 4430
rect 26305 4395 26315 4415
rect 26335 4395 26345 4415
rect 26305 4380 26345 4395
rect 26360 4415 26400 4430
rect 26360 4395 26370 4415
rect 26390 4395 26400 4415
rect 26360 4380 26400 4395
rect 26415 4415 26455 4430
rect 26415 4395 26425 4415
rect 26445 4395 26455 4415
rect 26415 4380 26455 4395
rect 26470 4415 26510 4430
rect 26470 4395 26480 4415
rect 26500 4395 26510 4415
rect 26470 4380 26510 4395
rect 26525 4415 26565 4430
rect 26525 4395 26535 4415
rect 26555 4395 26565 4415
rect 26525 4380 26565 4395
rect 26580 4415 26620 4430
rect 26580 4395 26590 4415
rect 26610 4395 26620 4415
rect 26580 4380 26620 4395
rect 26635 4415 26675 4430
rect 26635 4395 26645 4415
rect 26665 4395 26675 4415
rect 26635 4380 26675 4395
rect 26690 4415 26730 4430
rect 26690 4395 26700 4415
rect 26720 4395 26730 4415
rect 26690 4380 26730 4395
rect 26745 4415 26785 4430
rect 26745 4395 26755 4415
rect 26775 4395 26785 4415
rect 26745 4380 26785 4395
rect 26800 4415 26840 4430
rect 26800 4395 26810 4415
rect 26830 4395 26840 4415
rect 26800 4380 26840 4395
rect 26855 4415 26895 4430
rect 26855 4395 26865 4415
rect 26885 4395 26895 4415
rect 26855 4380 26895 4395
rect 26910 4415 26950 4430
rect 26910 4395 26920 4415
rect 26940 4395 26950 4415
rect 26910 4380 26950 4395
rect 26965 4415 27005 4430
rect 26965 4395 26975 4415
rect 26995 4395 27005 4415
rect 26965 4380 27005 4395
rect 27020 4415 27060 4430
rect 27020 4395 27030 4415
rect 27050 4395 27060 4415
rect 27020 4380 27060 4395
rect 27075 4415 27115 4430
rect 27075 4395 27085 4415
rect 27105 4395 27115 4415
rect 27075 4380 27115 4395
rect 27130 4415 27170 4430
rect 27130 4395 27140 4415
rect 27160 4395 27170 4415
rect 27130 4380 27170 4395
rect 27185 4415 27225 4430
rect 27185 4395 27195 4415
rect 27215 4395 27225 4415
rect 27185 4380 27225 4395
rect 27240 4415 27280 4430
rect 27240 4395 27250 4415
rect 27270 4395 27280 4415
rect 27240 4380 27280 4395
rect 27295 4415 27335 4430
rect 27295 4395 27305 4415
rect 27325 4395 27335 4415
rect 27295 4380 27335 4395
rect 27350 4415 27390 4430
rect 27350 4395 27360 4415
rect 27380 4395 27390 4415
rect 27350 4380 27390 4395
rect 27405 4415 27445 4430
rect 27405 4395 27415 4415
rect 27435 4395 27445 4415
rect 27405 4380 27445 4395
rect 27460 4415 27500 4430
rect 27460 4395 27470 4415
rect 27490 4395 27500 4415
rect 27460 4380 27500 4395
rect 16895 4320 16905 4340
rect 16925 4320 16935 4340
rect 16895 4290 16935 4320
rect 17185 4325 17225 4345
rect 17185 4305 17195 4325
rect 17215 4305 17225 4325
rect 17185 4285 17225 4305
rect 17245 4325 17285 4345
rect 17245 4305 17255 4325
rect 17275 4305 17285 4325
rect 17245 4285 17285 4305
rect 17305 4325 17345 4345
rect 17305 4305 17315 4325
rect 17335 4305 17345 4325
rect 17305 4285 17345 4305
rect 17365 4325 17405 4345
rect 17365 4305 17375 4325
rect 17395 4305 17405 4325
rect 17365 4285 17405 4305
rect 17425 4325 17465 4345
rect 17425 4305 17435 4325
rect 17455 4305 17465 4325
rect 17425 4285 17465 4305
rect 17485 4325 17525 4345
rect 17485 4305 17495 4325
rect 17515 4305 17525 4325
rect 17485 4285 17525 4305
rect 17545 4325 17585 4345
rect 17545 4305 17555 4325
rect 17575 4305 17585 4325
rect 17545 4285 17585 4305
rect 17605 4325 17645 4345
rect 17605 4305 17615 4325
rect 17635 4305 17645 4325
rect 17605 4285 17645 4305
rect 17665 4325 17705 4345
rect 17665 4305 17675 4325
rect 17695 4305 17705 4325
rect 17665 4285 17705 4305
rect 16250 4090 16290 4105
rect 16250 4070 16260 4090
rect 16280 4070 16290 4090
rect 16250 4055 16290 4070
rect 16305 4090 16345 4105
rect 16305 4070 16315 4090
rect 16335 4070 16345 4090
rect 16305 4055 16345 4070
rect 16360 4090 16400 4105
rect 16360 4070 16370 4090
rect 16390 4070 16400 4090
rect 16360 4055 16400 4070
rect 16415 4090 16455 4105
rect 16415 4070 16425 4090
rect 16445 4070 16455 4090
rect 16415 4055 16455 4070
rect 16470 4090 16510 4105
rect 16470 4070 16480 4090
rect 16500 4070 16510 4090
rect 16470 4055 16510 4070
rect 16525 4090 16565 4105
rect 16525 4070 16535 4090
rect 16555 4070 16565 4090
rect 16525 4055 16565 4070
rect 16580 4090 16620 4105
rect 16580 4070 16590 4090
rect 16610 4070 16620 4090
rect 16580 4055 16620 4070
rect 16635 4090 16675 4105
rect 16635 4070 16645 4090
rect 16665 4070 16675 4090
rect 16635 4055 16675 4070
rect 16690 4090 16730 4105
rect 16690 4070 16700 4090
rect 16720 4070 16730 4090
rect 16690 4055 16730 4070
rect 16745 4090 16785 4105
rect 16745 4070 16755 4090
rect 16775 4070 16785 4090
rect 16745 4055 16785 4070
rect 16800 4090 16840 4105
rect 16800 4070 16810 4090
rect 16830 4070 16840 4090
rect 16800 4055 16840 4070
rect 16855 4090 16895 4105
rect 16855 4070 16865 4090
rect 16885 4070 16895 4090
rect 16855 4055 16895 4070
rect 16910 4090 16950 4105
rect 16910 4070 16920 4090
rect 16940 4070 16950 4090
rect 16910 4055 16950 4070
rect 16965 4090 17005 4105
rect 16965 4070 16975 4090
rect 16995 4070 17005 4090
rect 16965 4055 17005 4070
rect 17020 4090 17060 4105
rect 17020 4070 17030 4090
rect 17050 4070 17060 4090
rect 17020 4055 17060 4070
rect 17075 4090 17115 4105
rect 17075 4070 17085 4090
rect 17105 4070 17115 4090
rect 17075 4055 17115 4070
rect 17130 4090 17170 4105
rect 17130 4070 17140 4090
rect 17160 4070 17170 4090
rect 17130 4055 17170 4070
rect 17185 4090 17225 4105
rect 17185 4070 17195 4090
rect 17215 4070 17225 4090
rect 17185 4055 17225 4070
rect 17240 4090 17280 4105
rect 17240 4070 17250 4090
rect 17270 4070 17280 4090
rect 17240 4055 17280 4070
rect 17295 4090 17335 4105
rect 17295 4070 17305 4090
rect 17325 4070 17335 4090
rect 17295 4055 17335 4070
rect 17350 4090 17390 4105
rect 17350 4070 17360 4090
rect 17380 4070 17390 4090
rect 17350 4055 17390 4070
rect 17405 4090 17445 4105
rect 17405 4070 17415 4090
rect 17435 4070 17445 4090
rect 17405 4055 17445 4070
rect 17460 4090 17500 4105
rect 17460 4070 17470 4090
rect 17490 4070 17500 4090
rect 17460 4055 17500 4070
rect 26200 4005 26240 4020
rect 26200 3985 26210 4005
rect 26230 3985 26240 4005
rect 26200 3970 26240 3985
rect 26255 4005 26295 4020
rect 26255 3985 26265 4005
rect 26285 3985 26295 4005
rect 26255 3970 26295 3985
rect 26310 4005 26350 4020
rect 26310 3985 26320 4005
rect 26340 3985 26350 4005
rect 26310 3970 26350 3985
rect 26365 4005 26405 4020
rect 26365 3985 26375 4005
rect 26395 3985 26405 4005
rect 26365 3970 26405 3985
rect 26420 4005 26460 4020
rect 26420 3985 26430 4005
rect 26450 3985 26460 4005
rect 26420 3970 26460 3985
rect 26475 4005 26515 4020
rect 26475 3985 26485 4005
rect 26505 3985 26515 4005
rect 26475 3970 26515 3985
rect 26530 4005 26570 4020
rect 26530 3985 26540 4005
rect 26560 3985 26570 4005
rect 26530 3970 26570 3985
rect 26585 4005 26625 4020
rect 26585 3985 26595 4005
rect 26615 3985 26625 4005
rect 26585 3970 26625 3985
rect 26640 4005 26680 4020
rect 26640 3985 26650 4005
rect 26670 3985 26680 4005
rect 26640 3970 26680 3985
rect 26695 4005 26735 4020
rect 26695 3985 26705 4005
rect 26725 3985 26735 4005
rect 26695 3970 26735 3985
rect 26750 4005 26790 4020
rect 26750 3985 26760 4005
rect 26780 3985 26790 4005
rect 26750 3970 26790 3985
rect 26805 4005 26845 4020
rect 26805 3985 26815 4005
rect 26835 3985 26845 4005
rect 26805 3970 26845 3985
rect 26860 4005 26900 4020
rect 26860 3985 26870 4005
rect 26890 3985 26900 4005
rect 26860 3970 26900 3985
rect 26930 4005 26970 4020
rect 26930 3985 26940 4005
rect 26960 3985 26970 4005
rect 26930 3970 26970 3985
rect 26985 4005 27025 4020
rect 26985 3985 26995 4005
rect 27015 3985 27025 4005
rect 26985 3970 27025 3985
rect 27040 4005 27080 4020
rect 27040 3985 27050 4005
rect 27070 3985 27080 4005
rect 27040 3970 27080 3985
rect 27095 4005 27135 4020
rect 27095 3985 27105 4005
rect 27125 3985 27135 4005
rect 27095 3970 27135 3985
rect 27150 4005 27190 4020
rect 27150 3985 27160 4005
rect 27180 3985 27190 4005
rect 27150 3970 27190 3985
rect 27205 4005 27245 4020
rect 27205 3985 27215 4005
rect 27235 3985 27245 4005
rect 27205 3970 27245 3985
rect 27260 4005 27300 4020
rect 27260 3985 27270 4005
rect 27290 3985 27300 4005
rect 27260 3970 27300 3985
rect 27315 4005 27355 4020
rect 27315 3985 27325 4005
rect 27345 3985 27355 4005
rect 27315 3970 27355 3985
rect 27370 4005 27410 4020
rect 27370 3985 27380 4005
rect 27400 3985 27410 4005
rect 27370 3970 27410 3985
rect 27425 4005 27465 4020
rect 27425 3985 27435 4005
rect 27455 3985 27465 4005
rect 27425 3970 27465 3985
rect 27480 4005 27520 4020
rect 27480 3985 27490 4005
rect 27510 3985 27520 4005
rect 27480 3970 27520 3985
rect 27535 4005 27575 4020
rect 27535 3985 27545 4005
rect 27565 3985 27575 4005
rect 27535 3970 27575 3985
rect 27590 4005 27630 4020
rect 27590 3985 27600 4005
rect 27620 3985 27630 4005
rect 27590 3970 27630 3985
rect 16195 3785 16235 3800
rect 16195 3765 16205 3785
rect 16225 3765 16235 3785
rect 16195 3750 16235 3765
rect 16250 3785 16290 3800
rect 16250 3765 16260 3785
rect 16280 3765 16290 3785
rect 16250 3750 16290 3765
rect 16305 3785 16345 3800
rect 16305 3765 16315 3785
rect 16335 3765 16345 3785
rect 16305 3750 16345 3765
rect 16360 3785 16400 3800
rect 16360 3765 16370 3785
rect 16390 3765 16400 3785
rect 16360 3750 16400 3765
rect 16415 3785 16455 3800
rect 16415 3765 16425 3785
rect 16445 3765 16455 3785
rect 16415 3750 16455 3765
rect 16470 3785 16510 3800
rect 16470 3765 16480 3785
rect 16500 3765 16510 3785
rect 16470 3750 16510 3765
rect 16525 3785 16565 3800
rect 16525 3765 16535 3785
rect 16555 3765 16565 3785
rect 16525 3750 16565 3765
rect 16580 3785 16620 3800
rect 16580 3765 16590 3785
rect 16610 3765 16620 3785
rect 16580 3750 16620 3765
rect 16635 3785 16675 3800
rect 16635 3765 16645 3785
rect 16665 3765 16675 3785
rect 16635 3750 16675 3765
rect 16690 3785 16730 3800
rect 16690 3765 16700 3785
rect 16720 3765 16730 3785
rect 16690 3750 16730 3765
rect 16745 3785 16785 3800
rect 16745 3765 16755 3785
rect 16775 3765 16785 3785
rect 16745 3750 16785 3765
rect 16800 3785 16840 3800
rect 16800 3765 16810 3785
rect 16830 3765 16840 3785
rect 16800 3750 16840 3765
rect 16855 3785 16895 3800
rect 16935 3785 16975 3800
rect 16855 3765 16865 3785
rect 16885 3765 16895 3785
rect 16935 3765 16945 3785
rect 16965 3765 16975 3785
rect 16855 3750 16895 3765
rect 16935 3750 16975 3765
rect 16990 3785 17030 3800
rect 16990 3765 17000 3785
rect 17020 3765 17030 3785
rect 16990 3750 17030 3765
rect 17045 3785 17085 3800
rect 17045 3765 17055 3785
rect 17075 3765 17085 3785
rect 17045 3750 17085 3765
rect 17100 3785 17140 3800
rect 17100 3765 17110 3785
rect 17130 3765 17140 3785
rect 17100 3750 17140 3765
rect 17155 3785 17195 3800
rect 17155 3765 17165 3785
rect 17185 3765 17195 3785
rect 17155 3750 17195 3765
rect 17210 3785 17250 3800
rect 17210 3765 17220 3785
rect 17240 3765 17250 3785
rect 17210 3750 17250 3765
rect 17265 3785 17305 3800
rect 17265 3765 17275 3785
rect 17295 3765 17305 3785
rect 17265 3750 17305 3765
rect 17320 3785 17360 3800
rect 17320 3765 17330 3785
rect 17350 3765 17360 3785
rect 17320 3750 17360 3765
rect 17375 3785 17415 3800
rect 17375 3765 17385 3785
rect 17405 3765 17415 3785
rect 17375 3750 17415 3765
rect 17430 3785 17470 3800
rect 17430 3765 17440 3785
rect 17460 3765 17470 3785
rect 17430 3750 17470 3765
rect 17485 3785 17525 3800
rect 17485 3765 17495 3785
rect 17515 3765 17525 3785
rect 17485 3750 17525 3765
rect 17540 3785 17580 3800
rect 17540 3765 17550 3785
rect 17570 3765 17580 3785
rect 17540 3750 17580 3765
rect 17595 3785 17635 3800
rect 17595 3765 17605 3785
rect 17625 3765 17635 3785
rect 17595 3750 17635 3765
rect 15005 3570 15045 3585
rect 15005 3550 15015 3570
rect 15035 3550 15045 3570
rect 15005 3520 15045 3550
rect 15005 3500 15015 3520
rect 15035 3500 15045 3520
rect 15005 3470 15045 3500
rect 15005 3450 15015 3470
rect 15035 3450 15045 3470
rect 15005 3420 15045 3450
rect 15005 3400 15015 3420
rect 15035 3400 15045 3420
rect 15005 3370 15045 3400
rect 15005 3350 15015 3370
rect 15035 3350 15045 3370
rect 15005 3320 15045 3350
rect 15005 3300 15015 3320
rect 15035 3300 15045 3320
rect 15005 3270 15045 3300
rect 15005 3250 15015 3270
rect 15035 3250 15045 3270
rect 15005 3220 15045 3250
rect 15005 3200 15015 3220
rect 15035 3200 15045 3220
rect 15005 3170 15045 3200
rect 15005 3150 15015 3170
rect 15035 3150 15045 3170
rect 15005 3120 15045 3150
rect 15005 3100 15015 3120
rect 15035 3100 15045 3120
rect 15005 3070 15045 3100
rect 15005 3050 15015 3070
rect 15035 3050 15045 3070
rect 15005 3020 15045 3050
rect 15005 3000 15015 3020
rect 15035 3000 15045 3020
rect 15005 2985 15045 3000
rect 15060 3570 15100 3585
rect 15060 3550 15070 3570
rect 15090 3550 15100 3570
rect 15060 3520 15100 3550
rect 15060 3500 15070 3520
rect 15090 3500 15100 3520
rect 15060 3470 15100 3500
rect 15060 3450 15070 3470
rect 15090 3450 15100 3470
rect 15060 3420 15100 3450
rect 15060 3400 15070 3420
rect 15090 3400 15100 3420
rect 15060 3370 15100 3400
rect 15060 3350 15070 3370
rect 15090 3350 15100 3370
rect 15060 3320 15100 3350
rect 15060 3300 15070 3320
rect 15090 3300 15100 3320
rect 15060 3270 15100 3300
rect 15060 3250 15070 3270
rect 15090 3250 15100 3270
rect 15060 3220 15100 3250
rect 15060 3200 15070 3220
rect 15090 3200 15100 3220
rect 15060 3170 15100 3200
rect 15060 3150 15070 3170
rect 15090 3150 15100 3170
rect 15060 3120 15100 3150
rect 15060 3100 15070 3120
rect 15090 3100 15100 3120
rect 15060 3070 15100 3100
rect 15060 3050 15070 3070
rect 15090 3050 15100 3070
rect 15060 3020 15100 3050
rect 15060 3000 15070 3020
rect 15090 3000 15100 3020
rect 15060 2985 15100 3000
rect 15115 3570 15155 3585
rect 15115 3550 15125 3570
rect 15145 3550 15155 3570
rect 15115 3520 15155 3550
rect 15115 3500 15125 3520
rect 15145 3500 15155 3520
rect 15115 3470 15155 3500
rect 15115 3450 15125 3470
rect 15145 3450 15155 3470
rect 15115 3420 15155 3450
rect 15115 3400 15125 3420
rect 15145 3400 15155 3420
rect 15115 3370 15155 3400
rect 15115 3350 15125 3370
rect 15145 3350 15155 3370
rect 15115 3320 15155 3350
rect 15115 3300 15125 3320
rect 15145 3300 15155 3320
rect 15115 3270 15155 3300
rect 15115 3250 15125 3270
rect 15145 3250 15155 3270
rect 15115 3220 15155 3250
rect 15115 3200 15125 3220
rect 15145 3200 15155 3220
rect 15115 3170 15155 3200
rect 15115 3150 15125 3170
rect 15145 3150 15155 3170
rect 15115 3120 15155 3150
rect 15115 3100 15125 3120
rect 15145 3100 15155 3120
rect 15115 3070 15155 3100
rect 15115 3050 15125 3070
rect 15145 3050 15155 3070
rect 15115 3020 15155 3050
rect 15115 3000 15125 3020
rect 15145 3000 15155 3020
rect 15115 2985 15155 3000
rect 15170 3570 15210 3585
rect 15170 3550 15180 3570
rect 15200 3550 15210 3570
rect 15170 3520 15210 3550
rect 15170 3500 15180 3520
rect 15200 3500 15210 3520
rect 15170 3470 15210 3500
rect 15170 3450 15180 3470
rect 15200 3450 15210 3470
rect 15170 3420 15210 3450
rect 15170 3400 15180 3420
rect 15200 3400 15210 3420
rect 15170 3370 15210 3400
rect 15170 3350 15180 3370
rect 15200 3350 15210 3370
rect 15170 3320 15210 3350
rect 15170 3300 15180 3320
rect 15200 3300 15210 3320
rect 15170 3270 15210 3300
rect 15170 3250 15180 3270
rect 15200 3250 15210 3270
rect 15170 3220 15210 3250
rect 15170 3200 15180 3220
rect 15200 3200 15210 3220
rect 15170 3170 15210 3200
rect 15170 3150 15180 3170
rect 15200 3150 15210 3170
rect 15170 3120 15210 3150
rect 15170 3100 15180 3120
rect 15200 3100 15210 3120
rect 15170 3070 15210 3100
rect 15170 3050 15180 3070
rect 15200 3050 15210 3070
rect 15170 3020 15210 3050
rect 15170 3000 15180 3020
rect 15200 3000 15210 3020
rect 15170 2985 15210 3000
rect 15225 3570 15265 3585
rect 15225 3550 15235 3570
rect 15255 3550 15265 3570
rect 15225 3520 15265 3550
rect 15225 3500 15235 3520
rect 15255 3500 15265 3520
rect 15225 3470 15265 3500
rect 15225 3450 15235 3470
rect 15255 3450 15265 3470
rect 15225 3420 15265 3450
rect 15225 3400 15235 3420
rect 15255 3400 15265 3420
rect 15225 3370 15265 3400
rect 15225 3350 15235 3370
rect 15255 3350 15265 3370
rect 15225 3320 15265 3350
rect 15225 3300 15235 3320
rect 15255 3300 15265 3320
rect 15225 3270 15265 3300
rect 15225 3250 15235 3270
rect 15255 3250 15265 3270
rect 15225 3220 15265 3250
rect 15225 3200 15235 3220
rect 15255 3200 15265 3220
rect 15225 3170 15265 3200
rect 15225 3150 15235 3170
rect 15255 3150 15265 3170
rect 15225 3120 15265 3150
rect 15225 3100 15235 3120
rect 15255 3100 15265 3120
rect 15225 3070 15265 3100
rect 15225 3050 15235 3070
rect 15255 3050 15265 3070
rect 15225 3020 15265 3050
rect 15225 3000 15235 3020
rect 15255 3000 15265 3020
rect 15225 2985 15265 3000
rect 15280 3570 15320 3585
rect 15280 3550 15290 3570
rect 15310 3550 15320 3570
rect 15280 3520 15320 3550
rect 15280 3500 15290 3520
rect 15310 3500 15320 3520
rect 15280 3470 15320 3500
rect 15280 3450 15290 3470
rect 15310 3450 15320 3470
rect 15280 3420 15320 3450
rect 15280 3400 15290 3420
rect 15310 3400 15320 3420
rect 15280 3370 15320 3400
rect 15280 3350 15290 3370
rect 15310 3350 15320 3370
rect 15280 3320 15320 3350
rect 15280 3300 15290 3320
rect 15310 3300 15320 3320
rect 15280 3270 15320 3300
rect 15280 3250 15290 3270
rect 15310 3250 15320 3270
rect 15280 3220 15320 3250
rect 15280 3200 15290 3220
rect 15310 3200 15320 3220
rect 15280 3170 15320 3200
rect 15280 3150 15290 3170
rect 15310 3150 15320 3170
rect 15280 3120 15320 3150
rect 15280 3100 15290 3120
rect 15310 3100 15320 3120
rect 15280 3070 15320 3100
rect 15280 3050 15290 3070
rect 15310 3050 15320 3070
rect 15280 3020 15320 3050
rect 15280 3000 15290 3020
rect 15310 3000 15320 3020
rect 15280 2985 15320 3000
rect 15335 3570 15375 3585
rect 15335 3550 15345 3570
rect 15365 3550 15375 3570
rect 15335 3520 15375 3550
rect 15335 3500 15345 3520
rect 15365 3500 15375 3520
rect 15335 3470 15375 3500
rect 15335 3450 15345 3470
rect 15365 3450 15375 3470
rect 15335 3420 15375 3450
rect 15335 3400 15345 3420
rect 15365 3400 15375 3420
rect 15335 3370 15375 3400
rect 15335 3350 15345 3370
rect 15365 3350 15375 3370
rect 15335 3320 15375 3350
rect 15335 3300 15345 3320
rect 15365 3300 15375 3320
rect 15335 3270 15375 3300
rect 15335 3250 15345 3270
rect 15365 3250 15375 3270
rect 15335 3220 15375 3250
rect 15335 3200 15345 3220
rect 15365 3200 15375 3220
rect 15335 3170 15375 3200
rect 15335 3150 15345 3170
rect 15365 3150 15375 3170
rect 15335 3120 15375 3150
rect 15335 3100 15345 3120
rect 15365 3100 15375 3120
rect 15335 3070 15375 3100
rect 15335 3050 15345 3070
rect 15365 3050 15375 3070
rect 15335 3020 15375 3050
rect 15335 3000 15345 3020
rect 15365 3000 15375 3020
rect 15335 2985 15375 3000
rect 15390 3570 15430 3585
rect 15390 3550 15400 3570
rect 15420 3550 15430 3570
rect 15390 3520 15430 3550
rect 15390 3500 15400 3520
rect 15420 3500 15430 3520
rect 15390 3470 15430 3500
rect 15390 3450 15400 3470
rect 15420 3450 15430 3470
rect 15390 3420 15430 3450
rect 15390 3400 15400 3420
rect 15420 3400 15430 3420
rect 15390 3370 15430 3400
rect 15390 3350 15400 3370
rect 15420 3350 15430 3370
rect 15390 3320 15430 3350
rect 15390 3300 15400 3320
rect 15420 3300 15430 3320
rect 15390 3270 15430 3300
rect 15390 3250 15400 3270
rect 15420 3250 15430 3270
rect 15390 3220 15430 3250
rect 15390 3200 15400 3220
rect 15420 3200 15430 3220
rect 15390 3170 15430 3200
rect 15390 3150 15400 3170
rect 15420 3150 15430 3170
rect 15390 3120 15430 3150
rect 15390 3100 15400 3120
rect 15420 3100 15430 3120
rect 15390 3070 15430 3100
rect 15390 3050 15400 3070
rect 15420 3050 15430 3070
rect 15390 3020 15430 3050
rect 15390 3000 15400 3020
rect 15420 3000 15430 3020
rect 15390 2985 15430 3000
rect 15445 3570 15485 3585
rect 15445 3550 15455 3570
rect 15475 3550 15485 3570
rect 15445 3520 15485 3550
rect 15445 3500 15455 3520
rect 15475 3500 15485 3520
rect 15445 3470 15485 3500
rect 15445 3450 15455 3470
rect 15475 3450 15485 3470
rect 15445 3420 15485 3450
rect 15445 3400 15455 3420
rect 15475 3400 15485 3420
rect 15445 3370 15485 3400
rect 15445 3350 15455 3370
rect 15475 3350 15485 3370
rect 15445 3320 15485 3350
rect 15445 3300 15455 3320
rect 15475 3300 15485 3320
rect 15445 3270 15485 3300
rect 15445 3250 15455 3270
rect 15475 3250 15485 3270
rect 15445 3220 15485 3250
rect 15445 3200 15455 3220
rect 15475 3200 15485 3220
rect 15445 3170 15485 3200
rect 15445 3150 15455 3170
rect 15475 3150 15485 3170
rect 15445 3120 15485 3150
rect 15445 3100 15455 3120
rect 15475 3100 15485 3120
rect 15445 3070 15485 3100
rect 15445 3050 15455 3070
rect 15475 3050 15485 3070
rect 15445 3020 15485 3050
rect 15445 3000 15455 3020
rect 15475 3000 15485 3020
rect 15445 2985 15485 3000
rect 15500 3570 15540 3585
rect 15500 3550 15510 3570
rect 15530 3550 15540 3570
rect 15500 3520 15540 3550
rect 15500 3500 15510 3520
rect 15530 3500 15540 3520
rect 15500 3470 15540 3500
rect 15500 3450 15510 3470
rect 15530 3450 15540 3470
rect 15500 3420 15540 3450
rect 15500 3400 15510 3420
rect 15530 3400 15540 3420
rect 15500 3370 15540 3400
rect 15500 3350 15510 3370
rect 15530 3350 15540 3370
rect 15500 3320 15540 3350
rect 15500 3300 15510 3320
rect 15530 3300 15540 3320
rect 15500 3270 15540 3300
rect 15500 3250 15510 3270
rect 15530 3250 15540 3270
rect 15500 3220 15540 3250
rect 15500 3200 15510 3220
rect 15530 3200 15540 3220
rect 15500 3170 15540 3200
rect 15500 3150 15510 3170
rect 15530 3150 15540 3170
rect 15500 3120 15540 3150
rect 15500 3100 15510 3120
rect 15530 3100 15540 3120
rect 15500 3070 15540 3100
rect 15500 3050 15510 3070
rect 15530 3050 15540 3070
rect 15500 3020 15540 3050
rect 15500 3000 15510 3020
rect 15530 3000 15540 3020
rect 15500 2985 15540 3000
rect 15555 3570 15595 3585
rect 15555 3550 15565 3570
rect 15585 3550 15595 3570
rect 15555 3520 15595 3550
rect 15555 3500 15565 3520
rect 15585 3500 15595 3520
rect 15555 3470 15595 3500
rect 15555 3450 15565 3470
rect 15585 3450 15595 3470
rect 15555 3420 15595 3450
rect 15555 3400 15565 3420
rect 15585 3400 15595 3420
rect 15555 3370 15595 3400
rect 15555 3350 15565 3370
rect 15585 3350 15595 3370
rect 15555 3320 15595 3350
rect 15555 3300 15565 3320
rect 15585 3300 15595 3320
rect 15555 3270 15595 3300
rect 15555 3250 15565 3270
rect 15585 3250 15595 3270
rect 15555 3220 15595 3250
rect 15555 3200 15565 3220
rect 15585 3200 15595 3220
rect 15555 3170 15595 3200
rect 15555 3150 15565 3170
rect 15585 3150 15595 3170
rect 15555 3120 15595 3150
rect 15555 3100 15565 3120
rect 15585 3100 15595 3120
rect 15555 3070 15595 3100
rect 15555 3050 15565 3070
rect 15585 3050 15595 3070
rect 15555 3020 15595 3050
rect 15555 3000 15565 3020
rect 15585 3000 15595 3020
rect 15555 2985 15595 3000
rect 15610 3570 15650 3585
rect 15610 3550 15620 3570
rect 15640 3550 15650 3570
rect 15610 3520 15650 3550
rect 15610 3500 15620 3520
rect 15640 3500 15650 3520
rect 15610 3470 15650 3500
rect 15610 3450 15620 3470
rect 15640 3450 15650 3470
rect 15610 3420 15650 3450
rect 15610 3400 15620 3420
rect 15640 3400 15650 3420
rect 15610 3370 15650 3400
rect 15610 3350 15620 3370
rect 15640 3350 15650 3370
rect 15610 3320 15650 3350
rect 15610 3300 15620 3320
rect 15640 3300 15650 3320
rect 15610 3270 15650 3300
rect 15610 3250 15620 3270
rect 15640 3250 15650 3270
rect 15610 3220 15650 3250
rect 15610 3200 15620 3220
rect 15640 3200 15650 3220
rect 15610 3170 15650 3200
rect 15610 3150 15620 3170
rect 15640 3150 15650 3170
rect 15610 3120 15650 3150
rect 15610 3100 15620 3120
rect 15640 3100 15650 3120
rect 15610 3070 15650 3100
rect 15610 3050 15620 3070
rect 15640 3050 15650 3070
rect 15610 3020 15650 3050
rect 15610 3000 15620 3020
rect 15640 3000 15650 3020
rect 15610 2985 15650 3000
rect 15665 3570 15705 3585
rect 15665 3550 15675 3570
rect 15695 3550 15705 3570
rect 15665 3520 15705 3550
rect 18145 3570 18185 3585
rect 18145 3550 18155 3570
rect 18175 3550 18185 3570
rect 15665 3500 15675 3520
rect 15695 3500 15705 3520
rect 15665 3470 15705 3500
rect 15665 3450 15675 3470
rect 15695 3450 15705 3470
rect 15665 3420 15705 3450
rect 15665 3400 15675 3420
rect 15695 3400 15705 3420
rect 15665 3370 15705 3400
rect 15665 3350 15675 3370
rect 15695 3350 15705 3370
rect 15665 3320 15705 3350
rect 15665 3300 15675 3320
rect 15695 3300 15705 3320
rect 15665 3270 15705 3300
rect 15665 3250 15675 3270
rect 15695 3250 15705 3270
rect 15665 3220 15705 3250
rect 15665 3200 15675 3220
rect 15695 3200 15705 3220
rect 15665 3170 15705 3200
rect 15665 3150 15675 3170
rect 15695 3150 15705 3170
rect 15665 3120 15705 3150
rect 16220 3510 16260 3525
rect 16220 3490 16230 3510
rect 16250 3490 16260 3510
rect 16220 3460 16260 3490
rect 16220 3440 16230 3460
rect 16250 3440 16260 3460
rect 16220 3410 16260 3440
rect 16220 3390 16230 3410
rect 16250 3390 16260 3410
rect 16220 3360 16260 3390
rect 16220 3340 16230 3360
rect 16250 3340 16260 3360
rect 16220 3310 16260 3340
rect 16220 3290 16230 3310
rect 16250 3290 16260 3310
rect 16220 3260 16260 3290
rect 16220 3240 16230 3260
rect 16250 3240 16260 3260
rect 16220 3210 16260 3240
rect 16220 3190 16230 3210
rect 16250 3190 16260 3210
rect 16220 3160 16260 3190
rect 16220 3140 16230 3160
rect 16250 3140 16260 3160
rect 16220 3125 16260 3140
rect 16280 3510 16320 3525
rect 16280 3490 16290 3510
rect 16310 3490 16320 3510
rect 16280 3460 16320 3490
rect 16280 3440 16290 3460
rect 16310 3440 16320 3460
rect 16280 3410 16320 3440
rect 16280 3390 16290 3410
rect 16310 3390 16320 3410
rect 16280 3360 16320 3390
rect 16280 3340 16290 3360
rect 16310 3340 16320 3360
rect 16280 3310 16320 3340
rect 16280 3290 16290 3310
rect 16310 3290 16320 3310
rect 16280 3260 16320 3290
rect 16280 3240 16290 3260
rect 16310 3240 16320 3260
rect 16280 3210 16320 3240
rect 16280 3190 16290 3210
rect 16310 3190 16320 3210
rect 16280 3160 16320 3190
rect 16280 3140 16290 3160
rect 16310 3140 16320 3160
rect 16280 3125 16320 3140
rect 16340 3510 16380 3525
rect 16340 3490 16350 3510
rect 16370 3490 16380 3510
rect 16340 3460 16380 3490
rect 16340 3440 16350 3460
rect 16370 3440 16380 3460
rect 16340 3410 16380 3440
rect 16340 3390 16350 3410
rect 16370 3390 16380 3410
rect 16340 3360 16380 3390
rect 16340 3340 16350 3360
rect 16370 3340 16380 3360
rect 16340 3310 16380 3340
rect 16340 3290 16350 3310
rect 16370 3290 16380 3310
rect 16340 3260 16380 3290
rect 16340 3240 16350 3260
rect 16370 3240 16380 3260
rect 16340 3210 16380 3240
rect 16340 3190 16350 3210
rect 16370 3190 16380 3210
rect 16340 3160 16380 3190
rect 16340 3140 16350 3160
rect 16370 3140 16380 3160
rect 16340 3125 16380 3140
rect 16400 3510 16440 3525
rect 16400 3490 16410 3510
rect 16430 3490 16440 3510
rect 16400 3460 16440 3490
rect 16400 3440 16410 3460
rect 16430 3440 16440 3460
rect 16400 3410 16440 3440
rect 16400 3390 16410 3410
rect 16430 3390 16440 3410
rect 16400 3360 16440 3390
rect 16400 3340 16410 3360
rect 16430 3340 16440 3360
rect 16400 3310 16440 3340
rect 16400 3290 16410 3310
rect 16430 3290 16440 3310
rect 16400 3260 16440 3290
rect 16400 3240 16410 3260
rect 16430 3240 16440 3260
rect 16400 3210 16440 3240
rect 16400 3190 16410 3210
rect 16430 3190 16440 3210
rect 16400 3160 16440 3190
rect 16400 3140 16410 3160
rect 16430 3140 16440 3160
rect 16400 3125 16440 3140
rect 16460 3510 16500 3525
rect 16460 3490 16470 3510
rect 16490 3490 16500 3510
rect 16460 3460 16500 3490
rect 16460 3440 16470 3460
rect 16490 3440 16500 3460
rect 16460 3410 16500 3440
rect 16460 3390 16470 3410
rect 16490 3390 16500 3410
rect 16460 3360 16500 3390
rect 16460 3340 16470 3360
rect 16490 3340 16500 3360
rect 16460 3310 16500 3340
rect 16460 3290 16470 3310
rect 16490 3290 16500 3310
rect 16460 3260 16500 3290
rect 16460 3240 16470 3260
rect 16490 3240 16500 3260
rect 16460 3210 16500 3240
rect 16460 3190 16470 3210
rect 16490 3190 16500 3210
rect 16460 3160 16500 3190
rect 16460 3140 16470 3160
rect 16490 3140 16500 3160
rect 16460 3125 16500 3140
rect 16520 3510 16560 3525
rect 16520 3490 16530 3510
rect 16550 3490 16560 3510
rect 16520 3460 16560 3490
rect 16520 3440 16530 3460
rect 16550 3440 16560 3460
rect 16520 3410 16560 3440
rect 16520 3390 16530 3410
rect 16550 3390 16560 3410
rect 16520 3360 16560 3390
rect 16520 3340 16530 3360
rect 16550 3340 16560 3360
rect 16520 3310 16560 3340
rect 16520 3290 16530 3310
rect 16550 3290 16560 3310
rect 16520 3260 16560 3290
rect 16520 3240 16530 3260
rect 16550 3240 16560 3260
rect 16520 3210 16560 3240
rect 16520 3190 16530 3210
rect 16550 3190 16560 3210
rect 16520 3160 16560 3190
rect 16520 3140 16530 3160
rect 16550 3140 16560 3160
rect 16520 3125 16560 3140
rect 16580 3510 16620 3525
rect 16580 3490 16590 3510
rect 16610 3490 16620 3510
rect 16580 3460 16620 3490
rect 16580 3440 16590 3460
rect 16610 3440 16620 3460
rect 16580 3410 16620 3440
rect 16580 3390 16590 3410
rect 16610 3390 16620 3410
rect 16580 3360 16620 3390
rect 16580 3340 16590 3360
rect 16610 3340 16620 3360
rect 16580 3310 16620 3340
rect 16580 3290 16590 3310
rect 16610 3290 16620 3310
rect 16580 3260 16620 3290
rect 16580 3240 16590 3260
rect 16610 3240 16620 3260
rect 16580 3210 16620 3240
rect 16580 3190 16590 3210
rect 16610 3190 16620 3210
rect 16580 3160 16620 3190
rect 16580 3140 16590 3160
rect 16610 3140 16620 3160
rect 16580 3125 16620 3140
rect 16640 3510 16680 3525
rect 16640 3490 16650 3510
rect 16670 3490 16680 3510
rect 16640 3460 16680 3490
rect 16640 3440 16650 3460
rect 16670 3440 16680 3460
rect 16640 3410 16680 3440
rect 16640 3390 16650 3410
rect 16670 3390 16680 3410
rect 16640 3360 16680 3390
rect 16640 3340 16650 3360
rect 16670 3340 16680 3360
rect 16640 3310 16680 3340
rect 16640 3290 16650 3310
rect 16670 3290 16680 3310
rect 16640 3260 16680 3290
rect 16640 3240 16650 3260
rect 16670 3240 16680 3260
rect 16640 3210 16680 3240
rect 16640 3190 16650 3210
rect 16670 3190 16680 3210
rect 16640 3160 16680 3190
rect 16640 3140 16650 3160
rect 16670 3140 16680 3160
rect 16640 3125 16680 3140
rect 16700 3510 16740 3525
rect 16700 3490 16710 3510
rect 16730 3490 16740 3510
rect 16700 3460 16740 3490
rect 16700 3440 16710 3460
rect 16730 3440 16740 3460
rect 16700 3410 16740 3440
rect 16700 3390 16710 3410
rect 16730 3390 16740 3410
rect 16700 3360 16740 3390
rect 16700 3340 16710 3360
rect 16730 3340 16740 3360
rect 16700 3310 16740 3340
rect 16700 3290 16710 3310
rect 16730 3290 16740 3310
rect 16700 3260 16740 3290
rect 16700 3240 16710 3260
rect 16730 3240 16740 3260
rect 16700 3210 16740 3240
rect 16700 3190 16710 3210
rect 16730 3190 16740 3210
rect 16700 3160 16740 3190
rect 16700 3140 16710 3160
rect 16730 3140 16740 3160
rect 16700 3125 16740 3140
rect 16760 3510 16800 3525
rect 16760 3490 16770 3510
rect 16790 3490 16800 3510
rect 16760 3460 16800 3490
rect 16760 3440 16770 3460
rect 16790 3440 16800 3460
rect 16760 3410 16800 3440
rect 16760 3390 16770 3410
rect 16790 3390 16800 3410
rect 16760 3360 16800 3390
rect 16760 3340 16770 3360
rect 16790 3340 16800 3360
rect 16760 3310 16800 3340
rect 16760 3290 16770 3310
rect 16790 3290 16800 3310
rect 16760 3260 16800 3290
rect 16760 3240 16770 3260
rect 16790 3240 16800 3260
rect 16760 3210 16800 3240
rect 16760 3190 16770 3210
rect 16790 3190 16800 3210
rect 16760 3160 16800 3190
rect 16760 3140 16770 3160
rect 16790 3140 16800 3160
rect 16760 3125 16800 3140
rect 16820 3510 16860 3525
rect 16820 3490 16830 3510
rect 16850 3490 16860 3510
rect 16820 3460 16860 3490
rect 16820 3440 16830 3460
rect 16850 3440 16860 3460
rect 16820 3410 16860 3440
rect 16820 3390 16830 3410
rect 16850 3390 16860 3410
rect 16820 3360 16860 3390
rect 16820 3340 16830 3360
rect 16850 3340 16860 3360
rect 16820 3310 16860 3340
rect 16820 3290 16830 3310
rect 16850 3290 16860 3310
rect 16820 3260 16860 3290
rect 16820 3240 16830 3260
rect 16850 3240 16860 3260
rect 16820 3210 16860 3240
rect 16820 3190 16830 3210
rect 16850 3190 16860 3210
rect 16820 3160 16860 3190
rect 16820 3140 16830 3160
rect 16850 3140 16860 3160
rect 16820 3125 16860 3140
rect 16880 3510 16920 3525
rect 16880 3490 16890 3510
rect 16910 3490 16920 3510
rect 16880 3460 16920 3490
rect 16880 3440 16890 3460
rect 16910 3440 16920 3460
rect 16880 3410 16920 3440
rect 16880 3390 16890 3410
rect 16910 3390 16920 3410
rect 16880 3360 16920 3390
rect 16880 3340 16890 3360
rect 16910 3340 16920 3360
rect 16880 3310 16920 3340
rect 16880 3290 16890 3310
rect 16910 3290 16920 3310
rect 16880 3260 16920 3290
rect 16880 3240 16890 3260
rect 16910 3240 16920 3260
rect 16880 3210 16920 3240
rect 16880 3190 16890 3210
rect 16910 3190 16920 3210
rect 16880 3160 16920 3190
rect 16880 3140 16890 3160
rect 16910 3140 16920 3160
rect 16880 3125 16920 3140
rect 16940 3510 16980 3525
rect 16940 3490 16950 3510
rect 16970 3490 16980 3510
rect 16940 3460 16980 3490
rect 16940 3440 16950 3460
rect 16970 3440 16980 3460
rect 16940 3410 16980 3440
rect 16940 3390 16950 3410
rect 16970 3390 16980 3410
rect 16940 3360 16980 3390
rect 16940 3340 16950 3360
rect 16970 3340 16980 3360
rect 16940 3310 16980 3340
rect 16940 3290 16950 3310
rect 16970 3290 16980 3310
rect 16940 3260 16980 3290
rect 16940 3240 16950 3260
rect 16970 3240 16980 3260
rect 16940 3210 16980 3240
rect 16940 3190 16950 3210
rect 16970 3190 16980 3210
rect 16940 3160 16980 3190
rect 16940 3140 16950 3160
rect 16970 3140 16980 3160
rect 16940 3125 16980 3140
rect 17000 3510 17040 3525
rect 17000 3490 17010 3510
rect 17030 3490 17040 3510
rect 17000 3460 17040 3490
rect 17000 3440 17010 3460
rect 17030 3440 17040 3460
rect 17000 3410 17040 3440
rect 17000 3390 17010 3410
rect 17030 3390 17040 3410
rect 17000 3360 17040 3390
rect 17000 3340 17010 3360
rect 17030 3340 17040 3360
rect 17000 3310 17040 3340
rect 17000 3290 17010 3310
rect 17030 3290 17040 3310
rect 17000 3260 17040 3290
rect 17000 3240 17010 3260
rect 17030 3240 17040 3260
rect 17000 3210 17040 3240
rect 17000 3190 17010 3210
rect 17030 3190 17040 3210
rect 17000 3160 17040 3190
rect 17000 3140 17010 3160
rect 17030 3140 17040 3160
rect 17000 3125 17040 3140
rect 17060 3510 17100 3525
rect 17060 3490 17070 3510
rect 17090 3490 17100 3510
rect 17060 3460 17100 3490
rect 17060 3440 17070 3460
rect 17090 3440 17100 3460
rect 17060 3410 17100 3440
rect 17060 3390 17070 3410
rect 17090 3390 17100 3410
rect 17060 3360 17100 3390
rect 17060 3340 17070 3360
rect 17090 3340 17100 3360
rect 17060 3310 17100 3340
rect 17060 3290 17070 3310
rect 17090 3290 17100 3310
rect 17060 3260 17100 3290
rect 17060 3240 17070 3260
rect 17090 3240 17100 3260
rect 17060 3210 17100 3240
rect 17060 3190 17070 3210
rect 17090 3190 17100 3210
rect 17060 3160 17100 3190
rect 17060 3140 17070 3160
rect 17090 3140 17100 3160
rect 17060 3125 17100 3140
rect 17120 3510 17160 3525
rect 17120 3490 17130 3510
rect 17150 3490 17160 3510
rect 17120 3460 17160 3490
rect 17120 3440 17130 3460
rect 17150 3440 17160 3460
rect 17120 3410 17160 3440
rect 17120 3390 17130 3410
rect 17150 3390 17160 3410
rect 17120 3360 17160 3390
rect 17120 3340 17130 3360
rect 17150 3340 17160 3360
rect 17120 3310 17160 3340
rect 17120 3290 17130 3310
rect 17150 3290 17160 3310
rect 17120 3260 17160 3290
rect 17120 3240 17130 3260
rect 17150 3240 17160 3260
rect 17120 3210 17160 3240
rect 17120 3190 17130 3210
rect 17150 3190 17160 3210
rect 17120 3160 17160 3190
rect 17120 3140 17130 3160
rect 17150 3140 17160 3160
rect 17120 3125 17160 3140
rect 17180 3510 17220 3525
rect 17180 3490 17190 3510
rect 17210 3490 17220 3510
rect 17180 3460 17220 3490
rect 17180 3440 17190 3460
rect 17210 3440 17220 3460
rect 17180 3410 17220 3440
rect 17180 3390 17190 3410
rect 17210 3390 17220 3410
rect 17180 3360 17220 3390
rect 17180 3340 17190 3360
rect 17210 3340 17220 3360
rect 17180 3310 17220 3340
rect 17180 3290 17190 3310
rect 17210 3290 17220 3310
rect 17180 3260 17220 3290
rect 17180 3240 17190 3260
rect 17210 3240 17220 3260
rect 17180 3210 17220 3240
rect 17180 3190 17190 3210
rect 17210 3190 17220 3210
rect 17180 3160 17220 3190
rect 17180 3140 17190 3160
rect 17210 3140 17220 3160
rect 17180 3125 17220 3140
rect 17240 3510 17280 3525
rect 17240 3490 17250 3510
rect 17270 3490 17280 3510
rect 17240 3460 17280 3490
rect 17240 3440 17250 3460
rect 17270 3440 17280 3460
rect 17240 3410 17280 3440
rect 17240 3390 17250 3410
rect 17270 3390 17280 3410
rect 17240 3360 17280 3390
rect 17240 3340 17250 3360
rect 17270 3340 17280 3360
rect 17240 3310 17280 3340
rect 17240 3290 17250 3310
rect 17270 3290 17280 3310
rect 17240 3260 17280 3290
rect 17240 3240 17250 3260
rect 17270 3240 17280 3260
rect 17240 3210 17280 3240
rect 17240 3190 17250 3210
rect 17270 3190 17280 3210
rect 17240 3160 17280 3190
rect 17240 3140 17250 3160
rect 17270 3140 17280 3160
rect 17240 3125 17280 3140
rect 17300 3510 17340 3525
rect 17300 3490 17310 3510
rect 17330 3490 17340 3510
rect 17300 3460 17340 3490
rect 17300 3440 17310 3460
rect 17330 3440 17340 3460
rect 17300 3410 17340 3440
rect 17300 3390 17310 3410
rect 17330 3390 17340 3410
rect 17300 3360 17340 3390
rect 17300 3340 17310 3360
rect 17330 3340 17340 3360
rect 17300 3310 17340 3340
rect 17300 3290 17310 3310
rect 17330 3290 17340 3310
rect 17300 3260 17340 3290
rect 17300 3240 17310 3260
rect 17330 3240 17340 3260
rect 17300 3210 17340 3240
rect 17300 3190 17310 3210
rect 17330 3190 17340 3210
rect 17300 3160 17340 3190
rect 17300 3140 17310 3160
rect 17330 3140 17340 3160
rect 17300 3125 17340 3140
rect 17360 3510 17400 3525
rect 17360 3490 17370 3510
rect 17390 3490 17400 3510
rect 17360 3460 17400 3490
rect 17360 3440 17370 3460
rect 17390 3440 17400 3460
rect 17360 3410 17400 3440
rect 17360 3390 17370 3410
rect 17390 3390 17400 3410
rect 17360 3360 17400 3390
rect 17360 3340 17370 3360
rect 17390 3340 17400 3360
rect 17360 3310 17400 3340
rect 17360 3290 17370 3310
rect 17390 3290 17400 3310
rect 17360 3260 17400 3290
rect 17360 3240 17370 3260
rect 17390 3240 17400 3260
rect 17360 3210 17400 3240
rect 17360 3190 17370 3210
rect 17390 3190 17400 3210
rect 17360 3160 17400 3190
rect 17360 3140 17370 3160
rect 17390 3140 17400 3160
rect 17360 3125 17400 3140
rect 17420 3510 17460 3525
rect 17420 3490 17430 3510
rect 17450 3490 17460 3510
rect 17420 3460 17460 3490
rect 17420 3440 17430 3460
rect 17450 3440 17460 3460
rect 17420 3410 17460 3440
rect 17420 3390 17430 3410
rect 17450 3390 17460 3410
rect 17420 3360 17460 3390
rect 17420 3340 17430 3360
rect 17450 3340 17460 3360
rect 17420 3310 17460 3340
rect 17420 3290 17430 3310
rect 17450 3290 17460 3310
rect 17420 3260 17460 3290
rect 17420 3240 17430 3260
rect 17450 3240 17460 3260
rect 17420 3210 17460 3240
rect 17420 3190 17430 3210
rect 17450 3190 17460 3210
rect 17420 3160 17460 3190
rect 17420 3140 17430 3160
rect 17450 3140 17460 3160
rect 17420 3125 17460 3140
rect 17480 3510 17520 3525
rect 17480 3490 17490 3510
rect 17510 3490 17520 3510
rect 17480 3460 17520 3490
rect 17480 3440 17490 3460
rect 17510 3440 17520 3460
rect 17480 3410 17520 3440
rect 17480 3390 17490 3410
rect 17510 3390 17520 3410
rect 17480 3360 17520 3390
rect 17480 3340 17490 3360
rect 17510 3340 17520 3360
rect 17480 3310 17520 3340
rect 17480 3290 17490 3310
rect 17510 3290 17520 3310
rect 17480 3260 17520 3290
rect 17480 3240 17490 3260
rect 17510 3240 17520 3260
rect 17480 3210 17520 3240
rect 17480 3190 17490 3210
rect 17510 3190 17520 3210
rect 17480 3160 17520 3190
rect 17480 3140 17490 3160
rect 17510 3140 17520 3160
rect 17480 3125 17520 3140
rect 17540 3510 17580 3525
rect 17540 3490 17550 3510
rect 17570 3490 17580 3510
rect 17540 3460 17580 3490
rect 17540 3440 17550 3460
rect 17570 3440 17580 3460
rect 17540 3410 17580 3440
rect 17540 3390 17550 3410
rect 17570 3390 17580 3410
rect 17540 3360 17580 3390
rect 17540 3340 17550 3360
rect 17570 3340 17580 3360
rect 17540 3310 17580 3340
rect 17540 3290 17550 3310
rect 17570 3290 17580 3310
rect 17540 3260 17580 3290
rect 17540 3240 17550 3260
rect 17570 3240 17580 3260
rect 17540 3210 17580 3240
rect 17540 3190 17550 3210
rect 17570 3190 17580 3210
rect 17540 3160 17580 3190
rect 17540 3140 17550 3160
rect 17570 3140 17580 3160
rect 17540 3125 17580 3140
rect 18145 3520 18185 3550
rect 18145 3500 18155 3520
rect 18175 3500 18185 3520
rect 18145 3470 18185 3500
rect 18145 3450 18155 3470
rect 18175 3450 18185 3470
rect 18145 3420 18185 3450
rect 18145 3400 18155 3420
rect 18175 3400 18185 3420
rect 18145 3370 18185 3400
rect 18145 3350 18155 3370
rect 18175 3350 18185 3370
rect 18145 3320 18185 3350
rect 18145 3300 18155 3320
rect 18175 3300 18185 3320
rect 18145 3270 18185 3300
rect 18145 3250 18155 3270
rect 18175 3250 18185 3270
rect 18145 3220 18185 3250
rect 18145 3200 18155 3220
rect 18175 3200 18185 3220
rect 18145 3170 18185 3200
rect 18145 3150 18155 3170
rect 18175 3150 18185 3170
rect 15665 3100 15675 3120
rect 15695 3100 15705 3120
rect 18145 3120 18185 3150
rect 18145 3100 18155 3120
rect 18175 3100 18185 3120
rect 15665 3070 15705 3100
rect 18145 3070 18185 3100
rect 15665 3050 15675 3070
rect 15695 3050 15705 3070
rect 15665 3020 15705 3050
rect 15665 3000 15675 3020
rect 15695 3000 15705 3020
rect 15665 2985 15705 3000
rect 18145 3050 18155 3070
rect 18175 3050 18185 3070
rect 18145 3020 18185 3050
rect 18145 3000 18155 3020
rect 18175 3000 18185 3020
rect 18145 2985 18185 3000
rect 18200 3570 18240 3585
rect 18200 3550 18210 3570
rect 18230 3550 18240 3570
rect 18200 3520 18240 3550
rect 18200 3500 18210 3520
rect 18230 3500 18240 3520
rect 18200 3470 18240 3500
rect 18200 3450 18210 3470
rect 18230 3450 18240 3470
rect 18200 3420 18240 3450
rect 18200 3400 18210 3420
rect 18230 3400 18240 3420
rect 18200 3370 18240 3400
rect 18200 3350 18210 3370
rect 18230 3350 18240 3370
rect 18200 3320 18240 3350
rect 18200 3300 18210 3320
rect 18230 3300 18240 3320
rect 18200 3270 18240 3300
rect 18200 3250 18210 3270
rect 18230 3250 18240 3270
rect 18200 3220 18240 3250
rect 18200 3200 18210 3220
rect 18230 3200 18240 3220
rect 18200 3170 18240 3200
rect 18200 3150 18210 3170
rect 18230 3150 18240 3170
rect 18200 3120 18240 3150
rect 18200 3100 18210 3120
rect 18230 3100 18240 3120
rect 18200 3070 18240 3100
rect 18200 3050 18210 3070
rect 18230 3050 18240 3070
rect 18200 3020 18240 3050
rect 18200 3000 18210 3020
rect 18230 3000 18240 3020
rect 18200 2985 18240 3000
rect 18255 3570 18295 3585
rect 18255 3550 18265 3570
rect 18285 3550 18295 3570
rect 18255 3520 18295 3550
rect 18255 3500 18265 3520
rect 18285 3500 18295 3520
rect 18255 3470 18295 3500
rect 18255 3450 18265 3470
rect 18285 3450 18295 3470
rect 18255 3420 18295 3450
rect 18255 3400 18265 3420
rect 18285 3400 18295 3420
rect 18255 3370 18295 3400
rect 18255 3350 18265 3370
rect 18285 3350 18295 3370
rect 18255 3320 18295 3350
rect 18255 3300 18265 3320
rect 18285 3300 18295 3320
rect 18255 3270 18295 3300
rect 18255 3250 18265 3270
rect 18285 3250 18295 3270
rect 18255 3220 18295 3250
rect 18255 3200 18265 3220
rect 18285 3200 18295 3220
rect 18255 3170 18295 3200
rect 18255 3150 18265 3170
rect 18285 3150 18295 3170
rect 18255 3120 18295 3150
rect 18255 3100 18265 3120
rect 18285 3100 18295 3120
rect 18255 3070 18295 3100
rect 18255 3050 18265 3070
rect 18285 3050 18295 3070
rect 18255 3020 18295 3050
rect 18255 3000 18265 3020
rect 18285 3000 18295 3020
rect 18255 2985 18295 3000
rect 18310 3570 18350 3585
rect 18310 3550 18320 3570
rect 18340 3550 18350 3570
rect 18310 3520 18350 3550
rect 18310 3500 18320 3520
rect 18340 3500 18350 3520
rect 18310 3470 18350 3500
rect 18310 3450 18320 3470
rect 18340 3450 18350 3470
rect 18310 3420 18350 3450
rect 18310 3400 18320 3420
rect 18340 3400 18350 3420
rect 18310 3370 18350 3400
rect 18310 3350 18320 3370
rect 18340 3350 18350 3370
rect 18310 3320 18350 3350
rect 18310 3300 18320 3320
rect 18340 3300 18350 3320
rect 18310 3270 18350 3300
rect 18310 3250 18320 3270
rect 18340 3250 18350 3270
rect 18310 3220 18350 3250
rect 18310 3200 18320 3220
rect 18340 3200 18350 3220
rect 18310 3170 18350 3200
rect 18310 3150 18320 3170
rect 18340 3150 18350 3170
rect 18310 3120 18350 3150
rect 18310 3100 18320 3120
rect 18340 3100 18350 3120
rect 18310 3070 18350 3100
rect 18310 3050 18320 3070
rect 18340 3050 18350 3070
rect 18310 3020 18350 3050
rect 18310 3000 18320 3020
rect 18340 3000 18350 3020
rect 18310 2985 18350 3000
rect 18365 3570 18405 3585
rect 18365 3550 18375 3570
rect 18395 3550 18405 3570
rect 18365 3520 18405 3550
rect 18365 3500 18375 3520
rect 18395 3500 18405 3520
rect 18365 3470 18405 3500
rect 18365 3450 18375 3470
rect 18395 3450 18405 3470
rect 18365 3420 18405 3450
rect 18365 3400 18375 3420
rect 18395 3400 18405 3420
rect 18365 3370 18405 3400
rect 18365 3350 18375 3370
rect 18395 3350 18405 3370
rect 18365 3320 18405 3350
rect 18365 3300 18375 3320
rect 18395 3300 18405 3320
rect 18365 3270 18405 3300
rect 18365 3250 18375 3270
rect 18395 3250 18405 3270
rect 18365 3220 18405 3250
rect 18365 3200 18375 3220
rect 18395 3200 18405 3220
rect 18365 3170 18405 3200
rect 18365 3150 18375 3170
rect 18395 3150 18405 3170
rect 18365 3120 18405 3150
rect 18365 3100 18375 3120
rect 18395 3100 18405 3120
rect 18365 3070 18405 3100
rect 18365 3050 18375 3070
rect 18395 3050 18405 3070
rect 18365 3020 18405 3050
rect 18365 3000 18375 3020
rect 18395 3000 18405 3020
rect 18365 2985 18405 3000
rect 18420 3570 18460 3585
rect 18420 3550 18430 3570
rect 18450 3550 18460 3570
rect 18420 3520 18460 3550
rect 18420 3500 18430 3520
rect 18450 3500 18460 3520
rect 18420 3470 18460 3500
rect 18420 3450 18430 3470
rect 18450 3450 18460 3470
rect 18420 3420 18460 3450
rect 18420 3400 18430 3420
rect 18450 3400 18460 3420
rect 18420 3370 18460 3400
rect 18420 3350 18430 3370
rect 18450 3350 18460 3370
rect 18420 3320 18460 3350
rect 18420 3300 18430 3320
rect 18450 3300 18460 3320
rect 18420 3270 18460 3300
rect 18420 3250 18430 3270
rect 18450 3250 18460 3270
rect 18420 3220 18460 3250
rect 18420 3200 18430 3220
rect 18450 3200 18460 3220
rect 18420 3170 18460 3200
rect 18420 3150 18430 3170
rect 18450 3150 18460 3170
rect 18420 3120 18460 3150
rect 18420 3100 18430 3120
rect 18450 3100 18460 3120
rect 18420 3070 18460 3100
rect 18420 3050 18430 3070
rect 18450 3050 18460 3070
rect 18420 3020 18460 3050
rect 18420 3000 18430 3020
rect 18450 3000 18460 3020
rect 18420 2985 18460 3000
rect 18475 3570 18515 3585
rect 18475 3550 18485 3570
rect 18505 3550 18515 3570
rect 18475 3520 18515 3550
rect 18475 3500 18485 3520
rect 18505 3500 18515 3520
rect 18475 3470 18515 3500
rect 18475 3450 18485 3470
rect 18505 3450 18515 3470
rect 18475 3420 18515 3450
rect 18475 3400 18485 3420
rect 18505 3400 18515 3420
rect 18475 3370 18515 3400
rect 18475 3350 18485 3370
rect 18505 3350 18515 3370
rect 18475 3320 18515 3350
rect 18475 3300 18485 3320
rect 18505 3300 18515 3320
rect 18475 3270 18515 3300
rect 18475 3250 18485 3270
rect 18505 3250 18515 3270
rect 18475 3220 18515 3250
rect 18475 3200 18485 3220
rect 18505 3200 18515 3220
rect 18475 3170 18515 3200
rect 18475 3150 18485 3170
rect 18505 3150 18515 3170
rect 18475 3120 18515 3150
rect 18475 3100 18485 3120
rect 18505 3100 18515 3120
rect 18475 3070 18515 3100
rect 18475 3050 18485 3070
rect 18505 3050 18515 3070
rect 18475 3020 18515 3050
rect 18475 3000 18485 3020
rect 18505 3000 18515 3020
rect 18475 2985 18515 3000
rect 18530 3570 18570 3585
rect 18530 3550 18540 3570
rect 18560 3550 18570 3570
rect 18530 3520 18570 3550
rect 18530 3500 18540 3520
rect 18560 3500 18570 3520
rect 18530 3470 18570 3500
rect 18530 3450 18540 3470
rect 18560 3450 18570 3470
rect 18530 3420 18570 3450
rect 18530 3400 18540 3420
rect 18560 3400 18570 3420
rect 18530 3370 18570 3400
rect 18530 3350 18540 3370
rect 18560 3350 18570 3370
rect 18530 3320 18570 3350
rect 18530 3300 18540 3320
rect 18560 3300 18570 3320
rect 18530 3270 18570 3300
rect 18530 3250 18540 3270
rect 18560 3250 18570 3270
rect 18530 3220 18570 3250
rect 18530 3200 18540 3220
rect 18560 3200 18570 3220
rect 18530 3170 18570 3200
rect 18530 3150 18540 3170
rect 18560 3150 18570 3170
rect 18530 3120 18570 3150
rect 18530 3100 18540 3120
rect 18560 3100 18570 3120
rect 18530 3070 18570 3100
rect 18530 3050 18540 3070
rect 18560 3050 18570 3070
rect 18530 3020 18570 3050
rect 18530 3000 18540 3020
rect 18560 3000 18570 3020
rect 18530 2985 18570 3000
rect 18585 3570 18625 3585
rect 18585 3550 18595 3570
rect 18615 3550 18625 3570
rect 18585 3520 18625 3550
rect 18585 3500 18595 3520
rect 18615 3500 18625 3520
rect 18585 3470 18625 3500
rect 18585 3450 18595 3470
rect 18615 3450 18625 3470
rect 18585 3420 18625 3450
rect 18585 3400 18595 3420
rect 18615 3400 18625 3420
rect 18585 3370 18625 3400
rect 18585 3350 18595 3370
rect 18615 3350 18625 3370
rect 18585 3320 18625 3350
rect 18585 3300 18595 3320
rect 18615 3300 18625 3320
rect 18585 3270 18625 3300
rect 18585 3250 18595 3270
rect 18615 3250 18625 3270
rect 18585 3220 18625 3250
rect 18585 3200 18595 3220
rect 18615 3200 18625 3220
rect 18585 3170 18625 3200
rect 18585 3150 18595 3170
rect 18615 3150 18625 3170
rect 18585 3120 18625 3150
rect 18585 3100 18595 3120
rect 18615 3100 18625 3120
rect 18585 3070 18625 3100
rect 18585 3050 18595 3070
rect 18615 3050 18625 3070
rect 18585 3020 18625 3050
rect 18585 3000 18595 3020
rect 18615 3000 18625 3020
rect 18585 2985 18625 3000
rect 18640 3570 18680 3585
rect 18640 3550 18650 3570
rect 18670 3550 18680 3570
rect 18640 3520 18680 3550
rect 18640 3500 18650 3520
rect 18670 3500 18680 3520
rect 18640 3470 18680 3500
rect 18640 3450 18650 3470
rect 18670 3450 18680 3470
rect 18640 3420 18680 3450
rect 18640 3400 18650 3420
rect 18670 3400 18680 3420
rect 18640 3370 18680 3400
rect 18640 3350 18650 3370
rect 18670 3350 18680 3370
rect 18640 3320 18680 3350
rect 18640 3300 18650 3320
rect 18670 3300 18680 3320
rect 18640 3270 18680 3300
rect 18640 3250 18650 3270
rect 18670 3250 18680 3270
rect 18640 3220 18680 3250
rect 18640 3200 18650 3220
rect 18670 3200 18680 3220
rect 18640 3170 18680 3200
rect 18640 3150 18650 3170
rect 18670 3150 18680 3170
rect 18640 3120 18680 3150
rect 18640 3100 18650 3120
rect 18670 3100 18680 3120
rect 18640 3070 18680 3100
rect 18640 3050 18650 3070
rect 18670 3050 18680 3070
rect 18640 3020 18680 3050
rect 18640 3000 18650 3020
rect 18670 3000 18680 3020
rect 18640 2985 18680 3000
rect 18695 3570 18735 3585
rect 18695 3550 18705 3570
rect 18725 3550 18735 3570
rect 18695 3520 18735 3550
rect 18695 3500 18705 3520
rect 18725 3500 18735 3520
rect 18695 3470 18735 3500
rect 18695 3450 18705 3470
rect 18725 3450 18735 3470
rect 18695 3420 18735 3450
rect 18695 3400 18705 3420
rect 18725 3400 18735 3420
rect 18695 3370 18735 3400
rect 18695 3350 18705 3370
rect 18725 3350 18735 3370
rect 18695 3320 18735 3350
rect 18695 3300 18705 3320
rect 18725 3300 18735 3320
rect 18695 3270 18735 3300
rect 18695 3250 18705 3270
rect 18725 3250 18735 3270
rect 18695 3220 18735 3250
rect 18695 3200 18705 3220
rect 18725 3200 18735 3220
rect 18695 3170 18735 3200
rect 18695 3150 18705 3170
rect 18725 3150 18735 3170
rect 18695 3120 18735 3150
rect 18695 3100 18705 3120
rect 18725 3100 18735 3120
rect 18695 3070 18735 3100
rect 18695 3050 18705 3070
rect 18725 3050 18735 3070
rect 18695 3020 18735 3050
rect 18695 3000 18705 3020
rect 18725 3000 18735 3020
rect 18695 2985 18735 3000
rect 18750 3570 18790 3585
rect 18750 3550 18760 3570
rect 18780 3550 18790 3570
rect 18750 3520 18790 3550
rect 18750 3500 18760 3520
rect 18780 3500 18790 3520
rect 18750 3470 18790 3500
rect 18750 3450 18760 3470
rect 18780 3450 18790 3470
rect 18750 3420 18790 3450
rect 18750 3400 18760 3420
rect 18780 3400 18790 3420
rect 18750 3370 18790 3400
rect 18750 3350 18760 3370
rect 18780 3350 18790 3370
rect 18750 3320 18790 3350
rect 18750 3300 18760 3320
rect 18780 3300 18790 3320
rect 18750 3270 18790 3300
rect 18750 3250 18760 3270
rect 18780 3250 18790 3270
rect 18750 3220 18790 3250
rect 18750 3200 18760 3220
rect 18780 3200 18790 3220
rect 18750 3170 18790 3200
rect 18750 3150 18760 3170
rect 18780 3150 18790 3170
rect 18750 3120 18790 3150
rect 18750 3100 18760 3120
rect 18780 3100 18790 3120
rect 18750 3070 18790 3100
rect 18750 3050 18760 3070
rect 18780 3050 18790 3070
rect 18750 3020 18790 3050
rect 18750 3000 18760 3020
rect 18780 3000 18790 3020
rect 18750 2985 18790 3000
rect 18805 3570 18845 3585
rect 18805 3550 18815 3570
rect 18835 3550 18845 3570
rect 18805 3520 18845 3550
rect 25005 3570 25045 3585
rect 25005 3550 25015 3570
rect 25035 3550 25045 3570
rect 25005 3520 25045 3550
rect 18805 3500 18815 3520
rect 18835 3500 18845 3520
rect 18805 3470 18845 3500
rect 18805 3450 18815 3470
rect 18835 3450 18845 3470
rect 18805 3420 18845 3450
rect 18805 3400 18815 3420
rect 18835 3400 18845 3420
rect 18805 3370 18845 3400
rect 18805 3350 18815 3370
rect 18835 3350 18845 3370
rect 18805 3320 18845 3350
rect 18805 3300 18815 3320
rect 18835 3300 18845 3320
rect 18805 3270 18845 3300
rect 18805 3250 18815 3270
rect 18835 3250 18845 3270
rect 18805 3220 18845 3250
rect 18805 3200 18815 3220
rect 18835 3200 18845 3220
rect 18805 3170 18845 3200
rect 18805 3150 18815 3170
rect 18835 3150 18845 3170
rect 18805 3120 18845 3150
rect 18805 3100 18815 3120
rect 18835 3100 18845 3120
rect 18805 3070 18845 3100
rect 18805 3050 18815 3070
rect 18835 3050 18845 3070
rect 18805 3020 18845 3050
rect 18805 3000 18815 3020
rect 18835 3000 18845 3020
rect 18805 2985 18845 3000
rect 25005 3500 25015 3520
rect 25035 3500 25045 3520
rect 25005 3470 25045 3500
rect 25005 3450 25015 3470
rect 25035 3450 25045 3470
rect 25005 3420 25045 3450
rect 25005 3400 25015 3420
rect 25035 3400 25045 3420
rect 25005 3370 25045 3400
rect 25005 3350 25015 3370
rect 25035 3350 25045 3370
rect 25005 3320 25045 3350
rect 25005 3300 25015 3320
rect 25035 3300 25045 3320
rect 25005 3270 25045 3300
rect 25005 3250 25015 3270
rect 25035 3250 25045 3270
rect 25005 3220 25045 3250
rect 25005 3200 25015 3220
rect 25035 3200 25045 3220
rect 25005 3170 25045 3200
rect 25005 3150 25015 3170
rect 25035 3150 25045 3170
rect 25005 3120 25045 3150
rect 25005 3100 25015 3120
rect 25035 3100 25045 3120
rect 25005 3070 25045 3100
rect 25005 3050 25015 3070
rect 25035 3050 25045 3070
rect 25005 3020 25045 3050
rect 25005 3000 25015 3020
rect 25035 3000 25045 3020
rect 25005 2985 25045 3000
rect 25060 3570 25100 3585
rect 25060 3550 25070 3570
rect 25090 3550 25100 3570
rect 25060 3520 25100 3550
rect 25060 3500 25070 3520
rect 25090 3500 25100 3520
rect 25060 3470 25100 3500
rect 25060 3450 25070 3470
rect 25090 3450 25100 3470
rect 25060 3420 25100 3450
rect 25060 3400 25070 3420
rect 25090 3400 25100 3420
rect 25060 3370 25100 3400
rect 25060 3350 25070 3370
rect 25090 3350 25100 3370
rect 25060 3320 25100 3350
rect 25060 3300 25070 3320
rect 25090 3300 25100 3320
rect 25060 3270 25100 3300
rect 25060 3250 25070 3270
rect 25090 3250 25100 3270
rect 25060 3220 25100 3250
rect 25060 3200 25070 3220
rect 25090 3200 25100 3220
rect 25060 3170 25100 3200
rect 25060 3150 25070 3170
rect 25090 3150 25100 3170
rect 25060 3120 25100 3150
rect 25060 3100 25070 3120
rect 25090 3100 25100 3120
rect 25060 3070 25100 3100
rect 25060 3050 25070 3070
rect 25090 3050 25100 3070
rect 25060 3020 25100 3050
rect 25060 3000 25070 3020
rect 25090 3000 25100 3020
rect 25060 2985 25100 3000
rect 25115 3570 25155 3585
rect 25115 3550 25125 3570
rect 25145 3550 25155 3570
rect 25115 3520 25155 3550
rect 25115 3500 25125 3520
rect 25145 3500 25155 3520
rect 25115 3470 25155 3500
rect 25115 3450 25125 3470
rect 25145 3450 25155 3470
rect 25115 3420 25155 3450
rect 25115 3400 25125 3420
rect 25145 3400 25155 3420
rect 25115 3370 25155 3400
rect 25115 3350 25125 3370
rect 25145 3350 25155 3370
rect 25115 3320 25155 3350
rect 25115 3300 25125 3320
rect 25145 3300 25155 3320
rect 25115 3270 25155 3300
rect 25115 3250 25125 3270
rect 25145 3250 25155 3270
rect 25115 3220 25155 3250
rect 25115 3200 25125 3220
rect 25145 3200 25155 3220
rect 25115 3170 25155 3200
rect 25115 3150 25125 3170
rect 25145 3150 25155 3170
rect 25115 3120 25155 3150
rect 25115 3100 25125 3120
rect 25145 3100 25155 3120
rect 25115 3070 25155 3100
rect 25115 3050 25125 3070
rect 25145 3050 25155 3070
rect 25115 3020 25155 3050
rect 25115 3000 25125 3020
rect 25145 3000 25155 3020
rect 25115 2985 25155 3000
rect 25170 3570 25210 3585
rect 25170 3550 25180 3570
rect 25200 3550 25210 3570
rect 25170 3520 25210 3550
rect 25170 3500 25180 3520
rect 25200 3500 25210 3520
rect 25170 3470 25210 3500
rect 25170 3450 25180 3470
rect 25200 3450 25210 3470
rect 25170 3420 25210 3450
rect 25170 3400 25180 3420
rect 25200 3400 25210 3420
rect 25170 3370 25210 3400
rect 25170 3350 25180 3370
rect 25200 3350 25210 3370
rect 25170 3320 25210 3350
rect 25170 3300 25180 3320
rect 25200 3300 25210 3320
rect 25170 3270 25210 3300
rect 25170 3250 25180 3270
rect 25200 3250 25210 3270
rect 25170 3220 25210 3250
rect 25170 3200 25180 3220
rect 25200 3200 25210 3220
rect 25170 3170 25210 3200
rect 25170 3150 25180 3170
rect 25200 3150 25210 3170
rect 25170 3120 25210 3150
rect 25170 3100 25180 3120
rect 25200 3100 25210 3120
rect 25170 3070 25210 3100
rect 25170 3050 25180 3070
rect 25200 3050 25210 3070
rect 25170 3020 25210 3050
rect 25170 3000 25180 3020
rect 25200 3000 25210 3020
rect 25170 2985 25210 3000
rect 25225 3570 25265 3585
rect 25225 3550 25235 3570
rect 25255 3550 25265 3570
rect 25225 3520 25265 3550
rect 25225 3500 25235 3520
rect 25255 3500 25265 3520
rect 25225 3470 25265 3500
rect 25225 3450 25235 3470
rect 25255 3450 25265 3470
rect 25225 3420 25265 3450
rect 25225 3400 25235 3420
rect 25255 3400 25265 3420
rect 25225 3370 25265 3400
rect 25225 3350 25235 3370
rect 25255 3350 25265 3370
rect 25225 3320 25265 3350
rect 25225 3300 25235 3320
rect 25255 3300 25265 3320
rect 25225 3270 25265 3300
rect 25225 3250 25235 3270
rect 25255 3250 25265 3270
rect 25225 3220 25265 3250
rect 25225 3200 25235 3220
rect 25255 3200 25265 3220
rect 25225 3170 25265 3200
rect 25225 3150 25235 3170
rect 25255 3150 25265 3170
rect 25225 3120 25265 3150
rect 25225 3100 25235 3120
rect 25255 3100 25265 3120
rect 25225 3070 25265 3100
rect 25225 3050 25235 3070
rect 25255 3050 25265 3070
rect 25225 3020 25265 3050
rect 25225 3000 25235 3020
rect 25255 3000 25265 3020
rect 25225 2985 25265 3000
rect 25280 3570 25320 3585
rect 25280 3550 25290 3570
rect 25310 3550 25320 3570
rect 25280 3520 25320 3550
rect 25280 3500 25290 3520
rect 25310 3500 25320 3520
rect 25280 3470 25320 3500
rect 25280 3450 25290 3470
rect 25310 3450 25320 3470
rect 25280 3420 25320 3450
rect 25280 3400 25290 3420
rect 25310 3400 25320 3420
rect 25280 3370 25320 3400
rect 25280 3350 25290 3370
rect 25310 3350 25320 3370
rect 25280 3320 25320 3350
rect 25280 3300 25290 3320
rect 25310 3300 25320 3320
rect 25280 3270 25320 3300
rect 25280 3250 25290 3270
rect 25310 3250 25320 3270
rect 25280 3220 25320 3250
rect 25280 3200 25290 3220
rect 25310 3200 25320 3220
rect 25280 3170 25320 3200
rect 25280 3150 25290 3170
rect 25310 3150 25320 3170
rect 25280 3120 25320 3150
rect 25280 3100 25290 3120
rect 25310 3100 25320 3120
rect 25280 3070 25320 3100
rect 25280 3050 25290 3070
rect 25310 3050 25320 3070
rect 25280 3020 25320 3050
rect 25280 3000 25290 3020
rect 25310 3000 25320 3020
rect 25280 2985 25320 3000
rect 25335 3570 25375 3585
rect 25335 3550 25345 3570
rect 25365 3550 25375 3570
rect 25335 3520 25375 3550
rect 25335 3500 25345 3520
rect 25365 3500 25375 3520
rect 25335 3470 25375 3500
rect 25335 3450 25345 3470
rect 25365 3450 25375 3470
rect 25335 3420 25375 3450
rect 25335 3400 25345 3420
rect 25365 3400 25375 3420
rect 25335 3370 25375 3400
rect 25335 3350 25345 3370
rect 25365 3350 25375 3370
rect 25335 3320 25375 3350
rect 25335 3300 25345 3320
rect 25365 3300 25375 3320
rect 25335 3270 25375 3300
rect 25335 3250 25345 3270
rect 25365 3250 25375 3270
rect 25335 3220 25375 3250
rect 25335 3200 25345 3220
rect 25365 3200 25375 3220
rect 25335 3170 25375 3200
rect 25335 3150 25345 3170
rect 25365 3150 25375 3170
rect 25335 3120 25375 3150
rect 25335 3100 25345 3120
rect 25365 3100 25375 3120
rect 25335 3070 25375 3100
rect 25335 3050 25345 3070
rect 25365 3050 25375 3070
rect 25335 3020 25375 3050
rect 25335 3000 25345 3020
rect 25365 3000 25375 3020
rect 25335 2985 25375 3000
rect 25390 3570 25430 3585
rect 25390 3550 25400 3570
rect 25420 3550 25430 3570
rect 25390 3520 25430 3550
rect 25390 3500 25400 3520
rect 25420 3500 25430 3520
rect 25390 3470 25430 3500
rect 25390 3450 25400 3470
rect 25420 3450 25430 3470
rect 25390 3420 25430 3450
rect 25390 3400 25400 3420
rect 25420 3400 25430 3420
rect 25390 3370 25430 3400
rect 25390 3350 25400 3370
rect 25420 3350 25430 3370
rect 25390 3320 25430 3350
rect 25390 3300 25400 3320
rect 25420 3300 25430 3320
rect 25390 3270 25430 3300
rect 25390 3250 25400 3270
rect 25420 3250 25430 3270
rect 25390 3220 25430 3250
rect 25390 3200 25400 3220
rect 25420 3200 25430 3220
rect 25390 3170 25430 3200
rect 25390 3150 25400 3170
rect 25420 3150 25430 3170
rect 25390 3120 25430 3150
rect 25390 3100 25400 3120
rect 25420 3100 25430 3120
rect 25390 3070 25430 3100
rect 25390 3050 25400 3070
rect 25420 3050 25430 3070
rect 25390 3020 25430 3050
rect 25390 3000 25400 3020
rect 25420 3000 25430 3020
rect 25390 2985 25430 3000
rect 25445 3570 25485 3585
rect 25445 3550 25455 3570
rect 25475 3550 25485 3570
rect 25445 3520 25485 3550
rect 25445 3500 25455 3520
rect 25475 3500 25485 3520
rect 25445 3470 25485 3500
rect 25445 3450 25455 3470
rect 25475 3450 25485 3470
rect 25445 3420 25485 3450
rect 25445 3400 25455 3420
rect 25475 3400 25485 3420
rect 25445 3370 25485 3400
rect 25445 3350 25455 3370
rect 25475 3350 25485 3370
rect 25445 3320 25485 3350
rect 25445 3300 25455 3320
rect 25475 3300 25485 3320
rect 25445 3270 25485 3300
rect 25445 3250 25455 3270
rect 25475 3250 25485 3270
rect 25445 3220 25485 3250
rect 25445 3200 25455 3220
rect 25475 3200 25485 3220
rect 25445 3170 25485 3200
rect 25445 3150 25455 3170
rect 25475 3150 25485 3170
rect 25445 3120 25485 3150
rect 25445 3100 25455 3120
rect 25475 3100 25485 3120
rect 25445 3070 25485 3100
rect 25445 3050 25455 3070
rect 25475 3050 25485 3070
rect 25445 3020 25485 3050
rect 25445 3000 25455 3020
rect 25475 3000 25485 3020
rect 25445 2985 25485 3000
rect 25500 3570 25540 3585
rect 25500 3550 25510 3570
rect 25530 3550 25540 3570
rect 25500 3520 25540 3550
rect 25500 3500 25510 3520
rect 25530 3500 25540 3520
rect 25500 3470 25540 3500
rect 25500 3450 25510 3470
rect 25530 3450 25540 3470
rect 25500 3420 25540 3450
rect 25500 3400 25510 3420
rect 25530 3400 25540 3420
rect 25500 3370 25540 3400
rect 25500 3350 25510 3370
rect 25530 3350 25540 3370
rect 25500 3320 25540 3350
rect 25500 3300 25510 3320
rect 25530 3300 25540 3320
rect 25500 3270 25540 3300
rect 25500 3250 25510 3270
rect 25530 3250 25540 3270
rect 25500 3220 25540 3250
rect 25500 3200 25510 3220
rect 25530 3200 25540 3220
rect 25500 3170 25540 3200
rect 25500 3150 25510 3170
rect 25530 3150 25540 3170
rect 25500 3120 25540 3150
rect 25500 3100 25510 3120
rect 25530 3100 25540 3120
rect 25500 3070 25540 3100
rect 25500 3050 25510 3070
rect 25530 3050 25540 3070
rect 25500 3020 25540 3050
rect 25500 3000 25510 3020
rect 25530 3000 25540 3020
rect 25500 2985 25540 3000
rect 25555 3570 25595 3585
rect 25555 3550 25565 3570
rect 25585 3550 25595 3570
rect 25555 3520 25595 3550
rect 25555 3500 25565 3520
rect 25585 3500 25595 3520
rect 25555 3470 25595 3500
rect 25555 3450 25565 3470
rect 25585 3450 25595 3470
rect 25555 3420 25595 3450
rect 25555 3400 25565 3420
rect 25585 3400 25595 3420
rect 25555 3370 25595 3400
rect 25555 3350 25565 3370
rect 25585 3350 25595 3370
rect 25555 3320 25595 3350
rect 25555 3300 25565 3320
rect 25585 3300 25595 3320
rect 25555 3270 25595 3300
rect 25555 3250 25565 3270
rect 25585 3250 25595 3270
rect 25555 3220 25595 3250
rect 25555 3200 25565 3220
rect 25585 3200 25595 3220
rect 25555 3170 25595 3200
rect 25555 3150 25565 3170
rect 25585 3150 25595 3170
rect 25555 3120 25595 3150
rect 25555 3100 25565 3120
rect 25585 3100 25595 3120
rect 25555 3070 25595 3100
rect 25555 3050 25565 3070
rect 25585 3050 25595 3070
rect 25555 3020 25595 3050
rect 25555 3000 25565 3020
rect 25585 3000 25595 3020
rect 25555 2985 25595 3000
rect 25610 3570 25650 3585
rect 25610 3550 25620 3570
rect 25640 3550 25650 3570
rect 25610 3520 25650 3550
rect 25610 3500 25620 3520
rect 25640 3500 25650 3520
rect 25610 3470 25650 3500
rect 25610 3450 25620 3470
rect 25640 3450 25650 3470
rect 25610 3420 25650 3450
rect 25610 3400 25620 3420
rect 25640 3400 25650 3420
rect 25610 3370 25650 3400
rect 25610 3350 25620 3370
rect 25640 3350 25650 3370
rect 25610 3320 25650 3350
rect 25610 3300 25620 3320
rect 25640 3300 25650 3320
rect 25610 3270 25650 3300
rect 25610 3250 25620 3270
rect 25640 3250 25650 3270
rect 25610 3220 25650 3250
rect 25610 3200 25620 3220
rect 25640 3200 25650 3220
rect 25610 3170 25650 3200
rect 25610 3150 25620 3170
rect 25640 3150 25650 3170
rect 25610 3120 25650 3150
rect 25610 3100 25620 3120
rect 25640 3100 25650 3120
rect 25610 3070 25650 3100
rect 25610 3050 25620 3070
rect 25640 3050 25650 3070
rect 25610 3020 25650 3050
rect 25610 3000 25620 3020
rect 25640 3000 25650 3020
rect 25610 2985 25650 3000
rect 25665 3570 25705 3585
rect 25665 3550 25675 3570
rect 25695 3550 25705 3570
rect 25665 3520 25705 3550
rect 25665 3500 25675 3520
rect 25695 3500 25705 3520
rect 25665 3470 25705 3500
rect 25665 3450 25675 3470
rect 25695 3450 25705 3470
rect 25665 3420 25705 3450
rect 25665 3400 25675 3420
rect 25695 3400 25705 3420
rect 25665 3370 25705 3400
rect 25665 3350 25675 3370
rect 25695 3350 25705 3370
rect 25665 3320 25705 3350
rect 25665 3300 25675 3320
rect 25695 3300 25705 3320
rect 25665 3270 25705 3300
rect 25665 3250 25675 3270
rect 25695 3250 25705 3270
rect 25665 3220 25705 3250
rect 25665 3200 25675 3220
rect 25695 3200 25705 3220
rect 25665 3170 25705 3200
rect 25665 3150 25675 3170
rect 25695 3150 25705 3170
rect 25665 3120 25705 3150
rect 25665 3100 25675 3120
rect 25695 3100 25705 3120
rect 26220 3590 26260 3605
rect 26220 3570 26230 3590
rect 26250 3570 26260 3590
rect 26220 3540 26260 3570
rect 26220 3520 26230 3540
rect 26250 3520 26260 3540
rect 26220 3490 26260 3520
rect 26220 3470 26230 3490
rect 26250 3470 26260 3490
rect 26220 3440 26260 3470
rect 26220 3420 26230 3440
rect 26250 3420 26260 3440
rect 26220 3390 26260 3420
rect 26220 3370 26230 3390
rect 26250 3370 26260 3390
rect 26220 3340 26260 3370
rect 26220 3320 26230 3340
rect 26250 3320 26260 3340
rect 26220 3290 26260 3320
rect 26220 3270 26230 3290
rect 26250 3270 26260 3290
rect 26220 3240 26260 3270
rect 26220 3220 26230 3240
rect 26250 3220 26260 3240
rect 26220 3205 26260 3220
rect 26280 3590 26320 3605
rect 26280 3570 26290 3590
rect 26310 3570 26320 3590
rect 26280 3540 26320 3570
rect 26280 3520 26290 3540
rect 26310 3520 26320 3540
rect 26280 3490 26320 3520
rect 26280 3470 26290 3490
rect 26310 3470 26320 3490
rect 26280 3440 26320 3470
rect 26280 3420 26290 3440
rect 26310 3420 26320 3440
rect 26280 3390 26320 3420
rect 26280 3370 26290 3390
rect 26310 3370 26320 3390
rect 26280 3340 26320 3370
rect 26280 3320 26290 3340
rect 26310 3320 26320 3340
rect 26280 3290 26320 3320
rect 26280 3270 26290 3290
rect 26310 3270 26320 3290
rect 26280 3240 26320 3270
rect 26280 3220 26290 3240
rect 26310 3220 26320 3240
rect 26280 3205 26320 3220
rect 26340 3590 26380 3605
rect 26340 3570 26350 3590
rect 26370 3570 26380 3590
rect 26340 3540 26380 3570
rect 26340 3520 26350 3540
rect 26370 3520 26380 3540
rect 26340 3490 26380 3520
rect 26340 3470 26350 3490
rect 26370 3470 26380 3490
rect 26340 3440 26380 3470
rect 26340 3420 26350 3440
rect 26370 3420 26380 3440
rect 26340 3390 26380 3420
rect 26340 3370 26350 3390
rect 26370 3370 26380 3390
rect 26340 3340 26380 3370
rect 26340 3320 26350 3340
rect 26370 3320 26380 3340
rect 26340 3290 26380 3320
rect 26340 3270 26350 3290
rect 26370 3270 26380 3290
rect 26340 3240 26380 3270
rect 26340 3220 26350 3240
rect 26370 3220 26380 3240
rect 26340 3205 26380 3220
rect 26400 3590 26440 3605
rect 26400 3570 26410 3590
rect 26430 3570 26440 3590
rect 26400 3540 26440 3570
rect 26400 3520 26410 3540
rect 26430 3520 26440 3540
rect 26400 3490 26440 3520
rect 26400 3470 26410 3490
rect 26430 3470 26440 3490
rect 26400 3440 26440 3470
rect 26400 3420 26410 3440
rect 26430 3420 26440 3440
rect 26400 3390 26440 3420
rect 26400 3370 26410 3390
rect 26430 3370 26440 3390
rect 26400 3340 26440 3370
rect 26400 3320 26410 3340
rect 26430 3320 26440 3340
rect 26400 3290 26440 3320
rect 26400 3270 26410 3290
rect 26430 3270 26440 3290
rect 26400 3240 26440 3270
rect 26400 3220 26410 3240
rect 26430 3220 26440 3240
rect 26400 3205 26440 3220
rect 26460 3590 26500 3605
rect 26460 3570 26470 3590
rect 26490 3570 26500 3590
rect 26460 3540 26500 3570
rect 26460 3520 26470 3540
rect 26490 3520 26500 3540
rect 26460 3490 26500 3520
rect 26460 3470 26470 3490
rect 26490 3470 26500 3490
rect 26460 3440 26500 3470
rect 26460 3420 26470 3440
rect 26490 3420 26500 3440
rect 26460 3390 26500 3420
rect 26460 3370 26470 3390
rect 26490 3370 26500 3390
rect 26460 3340 26500 3370
rect 26460 3320 26470 3340
rect 26490 3320 26500 3340
rect 26460 3290 26500 3320
rect 26460 3270 26470 3290
rect 26490 3270 26500 3290
rect 26460 3240 26500 3270
rect 26460 3220 26470 3240
rect 26490 3220 26500 3240
rect 26460 3205 26500 3220
rect 26520 3590 26560 3605
rect 26520 3570 26530 3590
rect 26550 3570 26560 3590
rect 26520 3540 26560 3570
rect 26520 3520 26530 3540
rect 26550 3520 26560 3540
rect 26520 3490 26560 3520
rect 26520 3470 26530 3490
rect 26550 3470 26560 3490
rect 26520 3440 26560 3470
rect 26520 3420 26530 3440
rect 26550 3420 26560 3440
rect 26520 3390 26560 3420
rect 26520 3370 26530 3390
rect 26550 3370 26560 3390
rect 26520 3340 26560 3370
rect 26520 3320 26530 3340
rect 26550 3320 26560 3340
rect 26520 3290 26560 3320
rect 26520 3270 26530 3290
rect 26550 3270 26560 3290
rect 26520 3240 26560 3270
rect 26520 3220 26530 3240
rect 26550 3220 26560 3240
rect 26520 3205 26560 3220
rect 26580 3590 26620 3605
rect 26580 3570 26590 3590
rect 26610 3570 26620 3590
rect 26580 3540 26620 3570
rect 26580 3520 26590 3540
rect 26610 3520 26620 3540
rect 26580 3490 26620 3520
rect 26580 3470 26590 3490
rect 26610 3470 26620 3490
rect 26580 3440 26620 3470
rect 26580 3420 26590 3440
rect 26610 3420 26620 3440
rect 26580 3390 26620 3420
rect 26580 3370 26590 3390
rect 26610 3370 26620 3390
rect 26580 3340 26620 3370
rect 26580 3320 26590 3340
rect 26610 3320 26620 3340
rect 26580 3290 26620 3320
rect 26580 3270 26590 3290
rect 26610 3270 26620 3290
rect 26580 3240 26620 3270
rect 26580 3220 26590 3240
rect 26610 3220 26620 3240
rect 26580 3205 26620 3220
rect 26640 3590 26680 3605
rect 26640 3570 26650 3590
rect 26670 3570 26680 3590
rect 26640 3540 26680 3570
rect 26640 3520 26650 3540
rect 26670 3520 26680 3540
rect 26640 3490 26680 3520
rect 26640 3470 26650 3490
rect 26670 3470 26680 3490
rect 26640 3440 26680 3470
rect 26640 3420 26650 3440
rect 26670 3420 26680 3440
rect 26640 3390 26680 3420
rect 26640 3370 26650 3390
rect 26670 3370 26680 3390
rect 26640 3340 26680 3370
rect 26640 3320 26650 3340
rect 26670 3320 26680 3340
rect 26640 3290 26680 3320
rect 26640 3270 26650 3290
rect 26670 3270 26680 3290
rect 26640 3240 26680 3270
rect 26640 3220 26650 3240
rect 26670 3220 26680 3240
rect 26640 3205 26680 3220
rect 26700 3590 26740 3605
rect 26700 3570 26710 3590
rect 26730 3570 26740 3590
rect 26700 3540 26740 3570
rect 26700 3520 26710 3540
rect 26730 3520 26740 3540
rect 26700 3490 26740 3520
rect 26700 3470 26710 3490
rect 26730 3470 26740 3490
rect 26700 3440 26740 3470
rect 26700 3420 26710 3440
rect 26730 3420 26740 3440
rect 26700 3390 26740 3420
rect 26700 3370 26710 3390
rect 26730 3370 26740 3390
rect 26700 3340 26740 3370
rect 26700 3320 26710 3340
rect 26730 3320 26740 3340
rect 26700 3290 26740 3320
rect 26700 3270 26710 3290
rect 26730 3270 26740 3290
rect 26700 3240 26740 3270
rect 26700 3220 26710 3240
rect 26730 3220 26740 3240
rect 26700 3205 26740 3220
rect 26760 3590 26800 3605
rect 26760 3570 26770 3590
rect 26790 3570 26800 3590
rect 26760 3540 26800 3570
rect 26760 3520 26770 3540
rect 26790 3520 26800 3540
rect 26760 3490 26800 3520
rect 26760 3470 26770 3490
rect 26790 3470 26800 3490
rect 26760 3440 26800 3470
rect 26760 3420 26770 3440
rect 26790 3420 26800 3440
rect 26760 3390 26800 3420
rect 26760 3370 26770 3390
rect 26790 3370 26800 3390
rect 26760 3340 26800 3370
rect 26760 3320 26770 3340
rect 26790 3320 26800 3340
rect 26760 3290 26800 3320
rect 26760 3270 26770 3290
rect 26790 3270 26800 3290
rect 26760 3240 26800 3270
rect 26760 3220 26770 3240
rect 26790 3220 26800 3240
rect 26760 3205 26800 3220
rect 26820 3590 26860 3605
rect 26820 3570 26830 3590
rect 26850 3570 26860 3590
rect 26820 3540 26860 3570
rect 26820 3520 26830 3540
rect 26850 3520 26860 3540
rect 26820 3490 26860 3520
rect 26820 3470 26830 3490
rect 26850 3470 26860 3490
rect 26820 3440 26860 3470
rect 26820 3420 26830 3440
rect 26850 3420 26860 3440
rect 26820 3390 26860 3420
rect 26820 3370 26830 3390
rect 26850 3370 26860 3390
rect 26820 3340 26860 3370
rect 26820 3320 26830 3340
rect 26850 3320 26860 3340
rect 26820 3290 26860 3320
rect 26820 3270 26830 3290
rect 26850 3270 26860 3290
rect 26820 3240 26860 3270
rect 26820 3220 26830 3240
rect 26850 3220 26860 3240
rect 26820 3205 26860 3220
rect 26880 3590 26920 3605
rect 26880 3570 26890 3590
rect 26910 3570 26920 3590
rect 26880 3540 26920 3570
rect 26880 3520 26890 3540
rect 26910 3520 26920 3540
rect 26880 3490 26920 3520
rect 26880 3470 26890 3490
rect 26910 3470 26920 3490
rect 26880 3440 26920 3470
rect 26880 3420 26890 3440
rect 26910 3420 26920 3440
rect 26880 3390 26920 3420
rect 26880 3370 26890 3390
rect 26910 3370 26920 3390
rect 26880 3340 26920 3370
rect 26880 3320 26890 3340
rect 26910 3320 26920 3340
rect 26880 3290 26920 3320
rect 26880 3270 26890 3290
rect 26910 3270 26920 3290
rect 26880 3240 26920 3270
rect 26880 3220 26890 3240
rect 26910 3220 26920 3240
rect 26880 3205 26920 3220
rect 26940 3590 26980 3605
rect 26940 3570 26950 3590
rect 26970 3570 26980 3590
rect 26940 3540 26980 3570
rect 26940 3520 26950 3540
rect 26970 3520 26980 3540
rect 26940 3490 26980 3520
rect 26940 3470 26950 3490
rect 26970 3470 26980 3490
rect 26940 3440 26980 3470
rect 26940 3420 26950 3440
rect 26970 3420 26980 3440
rect 26940 3390 26980 3420
rect 26940 3370 26950 3390
rect 26970 3370 26980 3390
rect 26940 3340 26980 3370
rect 26940 3320 26950 3340
rect 26970 3320 26980 3340
rect 26940 3290 26980 3320
rect 26940 3270 26950 3290
rect 26970 3270 26980 3290
rect 26940 3240 26980 3270
rect 26940 3220 26950 3240
rect 26970 3220 26980 3240
rect 26940 3205 26980 3220
rect 27000 3590 27040 3605
rect 27000 3570 27010 3590
rect 27030 3570 27040 3590
rect 27000 3540 27040 3570
rect 27000 3520 27010 3540
rect 27030 3520 27040 3540
rect 27000 3490 27040 3520
rect 27000 3470 27010 3490
rect 27030 3470 27040 3490
rect 27000 3440 27040 3470
rect 27000 3420 27010 3440
rect 27030 3420 27040 3440
rect 27000 3390 27040 3420
rect 27000 3370 27010 3390
rect 27030 3370 27040 3390
rect 27000 3340 27040 3370
rect 27000 3320 27010 3340
rect 27030 3320 27040 3340
rect 27000 3290 27040 3320
rect 27000 3270 27010 3290
rect 27030 3270 27040 3290
rect 27000 3240 27040 3270
rect 27000 3220 27010 3240
rect 27030 3220 27040 3240
rect 27000 3205 27040 3220
rect 27060 3590 27100 3605
rect 27060 3570 27070 3590
rect 27090 3570 27100 3590
rect 27060 3540 27100 3570
rect 27060 3520 27070 3540
rect 27090 3520 27100 3540
rect 27060 3490 27100 3520
rect 27060 3470 27070 3490
rect 27090 3470 27100 3490
rect 27060 3440 27100 3470
rect 27060 3420 27070 3440
rect 27090 3420 27100 3440
rect 27060 3390 27100 3420
rect 27060 3370 27070 3390
rect 27090 3370 27100 3390
rect 27060 3340 27100 3370
rect 27060 3320 27070 3340
rect 27090 3320 27100 3340
rect 27060 3290 27100 3320
rect 27060 3270 27070 3290
rect 27090 3270 27100 3290
rect 27060 3240 27100 3270
rect 27060 3220 27070 3240
rect 27090 3220 27100 3240
rect 27060 3205 27100 3220
rect 27120 3590 27160 3605
rect 27120 3570 27130 3590
rect 27150 3570 27160 3590
rect 27120 3540 27160 3570
rect 27120 3520 27130 3540
rect 27150 3520 27160 3540
rect 27120 3490 27160 3520
rect 27120 3470 27130 3490
rect 27150 3470 27160 3490
rect 27120 3440 27160 3470
rect 27120 3420 27130 3440
rect 27150 3420 27160 3440
rect 27120 3390 27160 3420
rect 27120 3370 27130 3390
rect 27150 3370 27160 3390
rect 27120 3340 27160 3370
rect 27120 3320 27130 3340
rect 27150 3320 27160 3340
rect 27120 3290 27160 3320
rect 27120 3270 27130 3290
rect 27150 3270 27160 3290
rect 27120 3240 27160 3270
rect 27120 3220 27130 3240
rect 27150 3220 27160 3240
rect 27120 3205 27160 3220
rect 27180 3590 27220 3605
rect 27180 3570 27190 3590
rect 27210 3570 27220 3590
rect 27180 3540 27220 3570
rect 27180 3520 27190 3540
rect 27210 3520 27220 3540
rect 27180 3490 27220 3520
rect 27180 3470 27190 3490
rect 27210 3470 27220 3490
rect 27180 3440 27220 3470
rect 27180 3420 27190 3440
rect 27210 3420 27220 3440
rect 27180 3390 27220 3420
rect 27180 3370 27190 3390
rect 27210 3370 27220 3390
rect 27180 3340 27220 3370
rect 27180 3320 27190 3340
rect 27210 3320 27220 3340
rect 27180 3290 27220 3320
rect 27180 3270 27190 3290
rect 27210 3270 27220 3290
rect 27180 3240 27220 3270
rect 27180 3220 27190 3240
rect 27210 3220 27220 3240
rect 27180 3205 27220 3220
rect 27240 3590 27280 3605
rect 27240 3570 27250 3590
rect 27270 3570 27280 3590
rect 27240 3540 27280 3570
rect 27240 3520 27250 3540
rect 27270 3520 27280 3540
rect 27240 3490 27280 3520
rect 27240 3470 27250 3490
rect 27270 3470 27280 3490
rect 27240 3440 27280 3470
rect 27240 3420 27250 3440
rect 27270 3420 27280 3440
rect 27240 3390 27280 3420
rect 27240 3370 27250 3390
rect 27270 3370 27280 3390
rect 27240 3340 27280 3370
rect 27240 3320 27250 3340
rect 27270 3320 27280 3340
rect 27240 3290 27280 3320
rect 27240 3270 27250 3290
rect 27270 3270 27280 3290
rect 27240 3240 27280 3270
rect 27240 3220 27250 3240
rect 27270 3220 27280 3240
rect 27240 3205 27280 3220
rect 27300 3590 27340 3605
rect 27300 3570 27310 3590
rect 27330 3570 27340 3590
rect 27300 3540 27340 3570
rect 27300 3520 27310 3540
rect 27330 3520 27340 3540
rect 27300 3490 27340 3520
rect 27300 3470 27310 3490
rect 27330 3470 27340 3490
rect 27300 3440 27340 3470
rect 27300 3420 27310 3440
rect 27330 3420 27340 3440
rect 27300 3390 27340 3420
rect 27300 3370 27310 3390
rect 27330 3370 27340 3390
rect 27300 3340 27340 3370
rect 27300 3320 27310 3340
rect 27330 3320 27340 3340
rect 27300 3290 27340 3320
rect 27300 3270 27310 3290
rect 27330 3270 27340 3290
rect 27300 3240 27340 3270
rect 27300 3220 27310 3240
rect 27330 3220 27340 3240
rect 27300 3205 27340 3220
rect 27360 3590 27400 3605
rect 27360 3570 27370 3590
rect 27390 3570 27400 3590
rect 27360 3540 27400 3570
rect 27360 3520 27370 3540
rect 27390 3520 27400 3540
rect 27360 3490 27400 3520
rect 27360 3470 27370 3490
rect 27390 3470 27400 3490
rect 27360 3440 27400 3470
rect 27360 3420 27370 3440
rect 27390 3420 27400 3440
rect 27360 3390 27400 3420
rect 27360 3370 27370 3390
rect 27390 3370 27400 3390
rect 27360 3340 27400 3370
rect 27360 3320 27370 3340
rect 27390 3320 27400 3340
rect 27360 3290 27400 3320
rect 27360 3270 27370 3290
rect 27390 3270 27400 3290
rect 27360 3240 27400 3270
rect 27360 3220 27370 3240
rect 27390 3220 27400 3240
rect 27360 3205 27400 3220
rect 27420 3590 27460 3605
rect 27420 3570 27430 3590
rect 27450 3570 27460 3590
rect 27420 3540 27460 3570
rect 27420 3520 27430 3540
rect 27450 3520 27460 3540
rect 27420 3490 27460 3520
rect 27420 3470 27430 3490
rect 27450 3470 27460 3490
rect 27420 3440 27460 3470
rect 27420 3420 27430 3440
rect 27450 3420 27460 3440
rect 27420 3390 27460 3420
rect 27420 3370 27430 3390
rect 27450 3370 27460 3390
rect 27420 3340 27460 3370
rect 27420 3320 27430 3340
rect 27450 3320 27460 3340
rect 27420 3290 27460 3320
rect 27420 3270 27430 3290
rect 27450 3270 27460 3290
rect 27420 3240 27460 3270
rect 27420 3220 27430 3240
rect 27450 3220 27460 3240
rect 27420 3205 27460 3220
rect 27480 3590 27520 3605
rect 27480 3570 27490 3590
rect 27510 3570 27520 3590
rect 27480 3540 27520 3570
rect 27480 3520 27490 3540
rect 27510 3520 27520 3540
rect 27480 3490 27520 3520
rect 27480 3470 27490 3490
rect 27510 3470 27520 3490
rect 27480 3440 27520 3470
rect 27480 3420 27490 3440
rect 27510 3420 27520 3440
rect 27480 3390 27520 3420
rect 27480 3370 27490 3390
rect 27510 3370 27520 3390
rect 27480 3340 27520 3370
rect 27480 3320 27490 3340
rect 27510 3320 27520 3340
rect 27480 3290 27520 3320
rect 27480 3270 27490 3290
rect 27510 3270 27520 3290
rect 27480 3240 27520 3270
rect 27480 3220 27490 3240
rect 27510 3220 27520 3240
rect 27480 3205 27520 3220
rect 27540 3590 27580 3605
rect 27540 3570 27550 3590
rect 27570 3570 27580 3590
rect 27540 3540 27580 3570
rect 27540 3520 27550 3540
rect 27570 3520 27580 3540
rect 27540 3490 27580 3520
rect 27540 3470 27550 3490
rect 27570 3470 27580 3490
rect 27540 3440 27580 3470
rect 27540 3420 27550 3440
rect 27570 3420 27580 3440
rect 27540 3390 27580 3420
rect 27540 3370 27550 3390
rect 27570 3370 27580 3390
rect 27540 3340 27580 3370
rect 27540 3320 27550 3340
rect 27570 3320 27580 3340
rect 27540 3290 27580 3320
rect 27540 3270 27550 3290
rect 27570 3270 27580 3290
rect 27540 3240 27580 3270
rect 27540 3220 27550 3240
rect 27570 3220 27580 3240
rect 27540 3205 27580 3220
rect 25665 3070 25705 3100
rect 25665 3050 25675 3070
rect 25695 3050 25705 3070
rect 25665 3020 25705 3050
rect 25665 3000 25675 3020
rect 25695 3000 25705 3020
rect 25665 2985 25705 3000
rect 28145 3650 28185 3665
rect 28145 3630 28155 3650
rect 28175 3630 28185 3650
rect 28145 3600 28185 3630
rect 28145 3580 28155 3600
rect 28175 3580 28185 3600
rect 28145 3550 28185 3580
rect 28145 3530 28155 3550
rect 28175 3530 28185 3550
rect 28145 3500 28185 3530
rect 28145 3480 28155 3500
rect 28175 3480 28185 3500
rect 28145 3450 28185 3480
rect 28145 3430 28155 3450
rect 28175 3430 28185 3450
rect 28145 3400 28185 3430
rect 28145 3380 28155 3400
rect 28175 3380 28185 3400
rect 28145 3350 28185 3380
rect 28145 3330 28155 3350
rect 28175 3330 28185 3350
rect 28145 3300 28185 3330
rect 28145 3280 28155 3300
rect 28175 3280 28185 3300
rect 28145 3250 28185 3280
rect 28145 3230 28155 3250
rect 28175 3230 28185 3250
rect 28145 3200 28185 3230
rect 28145 3180 28155 3200
rect 28175 3180 28185 3200
rect 28145 3150 28185 3180
rect 28145 3130 28155 3150
rect 28175 3130 28185 3150
rect 28145 3100 28185 3130
rect 28145 3080 28155 3100
rect 28175 3080 28185 3100
rect 28145 3065 28185 3080
rect 28200 3650 28240 3665
rect 28200 3630 28210 3650
rect 28230 3630 28240 3650
rect 28200 3600 28240 3630
rect 28200 3580 28210 3600
rect 28230 3580 28240 3600
rect 28200 3550 28240 3580
rect 28200 3530 28210 3550
rect 28230 3530 28240 3550
rect 28200 3500 28240 3530
rect 28200 3480 28210 3500
rect 28230 3480 28240 3500
rect 28200 3450 28240 3480
rect 28200 3430 28210 3450
rect 28230 3430 28240 3450
rect 28200 3400 28240 3430
rect 28200 3380 28210 3400
rect 28230 3380 28240 3400
rect 28200 3350 28240 3380
rect 28200 3330 28210 3350
rect 28230 3330 28240 3350
rect 28200 3300 28240 3330
rect 28200 3280 28210 3300
rect 28230 3280 28240 3300
rect 28200 3250 28240 3280
rect 28200 3230 28210 3250
rect 28230 3230 28240 3250
rect 28200 3200 28240 3230
rect 28200 3180 28210 3200
rect 28230 3180 28240 3200
rect 28200 3150 28240 3180
rect 28200 3130 28210 3150
rect 28230 3130 28240 3150
rect 28200 3100 28240 3130
rect 28200 3080 28210 3100
rect 28230 3080 28240 3100
rect 28200 3065 28240 3080
rect 28255 3650 28295 3665
rect 28255 3630 28265 3650
rect 28285 3630 28295 3650
rect 28255 3600 28295 3630
rect 28255 3580 28265 3600
rect 28285 3580 28295 3600
rect 28255 3550 28295 3580
rect 28255 3530 28265 3550
rect 28285 3530 28295 3550
rect 28255 3500 28295 3530
rect 28255 3480 28265 3500
rect 28285 3480 28295 3500
rect 28255 3450 28295 3480
rect 28255 3430 28265 3450
rect 28285 3430 28295 3450
rect 28255 3400 28295 3430
rect 28255 3380 28265 3400
rect 28285 3380 28295 3400
rect 28255 3350 28295 3380
rect 28255 3330 28265 3350
rect 28285 3330 28295 3350
rect 28255 3300 28295 3330
rect 28255 3280 28265 3300
rect 28285 3280 28295 3300
rect 28255 3250 28295 3280
rect 28255 3230 28265 3250
rect 28285 3230 28295 3250
rect 28255 3200 28295 3230
rect 28255 3180 28265 3200
rect 28285 3180 28295 3200
rect 28255 3150 28295 3180
rect 28255 3130 28265 3150
rect 28285 3130 28295 3150
rect 28255 3100 28295 3130
rect 28255 3080 28265 3100
rect 28285 3080 28295 3100
rect 28255 3065 28295 3080
rect 28310 3650 28350 3665
rect 28310 3630 28320 3650
rect 28340 3630 28350 3650
rect 28310 3600 28350 3630
rect 28310 3580 28320 3600
rect 28340 3580 28350 3600
rect 28310 3550 28350 3580
rect 28310 3530 28320 3550
rect 28340 3530 28350 3550
rect 28310 3500 28350 3530
rect 28310 3480 28320 3500
rect 28340 3480 28350 3500
rect 28310 3450 28350 3480
rect 28310 3430 28320 3450
rect 28340 3430 28350 3450
rect 28310 3400 28350 3430
rect 28310 3380 28320 3400
rect 28340 3380 28350 3400
rect 28310 3350 28350 3380
rect 28310 3330 28320 3350
rect 28340 3330 28350 3350
rect 28310 3300 28350 3330
rect 28310 3280 28320 3300
rect 28340 3280 28350 3300
rect 28310 3250 28350 3280
rect 28310 3230 28320 3250
rect 28340 3230 28350 3250
rect 28310 3200 28350 3230
rect 28310 3180 28320 3200
rect 28340 3180 28350 3200
rect 28310 3150 28350 3180
rect 28310 3130 28320 3150
rect 28340 3130 28350 3150
rect 28310 3100 28350 3130
rect 28310 3080 28320 3100
rect 28340 3080 28350 3100
rect 28310 3065 28350 3080
rect 28365 3650 28405 3665
rect 28365 3630 28375 3650
rect 28395 3630 28405 3650
rect 28365 3600 28405 3630
rect 28365 3580 28375 3600
rect 28395 3580 28405 3600
rect 28365 3550 28405 3580
rect 28365 3530 28375 3550
rect 28395 3530 28405 3550
rect 28365 3500 28405 3530
rect 28365 3480 28375 3500
rect 28395 3480 28405 3500
rect 28365 3450 28405 3480
rect 28365 3430 28375 3450
rect 28395 3430 28405 3450
rect 28365 3400 28405 3430
rect 28365 3380 28375 3400
rect 28395 3380 28405 3400
rect 28365 3350 28405 3380
rect 28365 3330 28375 3350
rect 28395 3330 28405 3350
rect 28365 3300 28405 3330
rect 28365 3280 28375 3300
rect 28395 3280 28405 3300
rect 28365 3250 28405 3280
rect 28365 3230 28375 3250
rect 28395 3230 28405 3250
rect 28365 3200 28405 3230
rect 28365 3180 28375 3200
rect 28395 3180 28405 3200
rect 28365 3150 28405 3180
rect 28365 3130 28375 3150
rect 28395 3130 28405 3150
rect 28365 3100 28405 3130
rect 28365 3080 28375 3100
rect 28395 3080 28405 3100
rect 28365 3065 28405 3080
rect 28420 3650 28460 3665
rect 28420 3630 28430 3650
rect 28450 3630 28460 3650
rect 28420 3600 28460 3630
rect 28420 3580 28430 3600
rect 28450 3580 28460 3600
rect 28420 3550 28460 3580
rect 28420 3530 28430 3550
rect 28450 3530 28460 3550
rect 28420 3500 28460 3530
rect 28420 3480 28430 3500
rect 28450 3480 28460 3500
rect 28420 3450 28460 3480
rect 28420 3430 28430 3450
rect 28450 3430 28460 3450
rect 28420 3400 28460 3430
rect 28420 3380 28430 3400
rect 28450 3380 28460 3400
rect 28420 3350 28460 3380
rect 28420 3330 28430 3350
rect 28450 3330 28460 3350
rect 28420 3300 28460 3330
rect 28420 3280 28430 3300
rect 28450 3280 28460 3300
rect 28420 3250 28460 3280
rect 28420 3230 28430 3250
rect 28450 3230 28460 3250
rect 28420 3200 28460 3230
rect 28420 3180 28430 3200
rect 28450 3180 28460 3200
rect 28420 3150 28460 3180
rect 28420 3130 28430 3150
rect 28450 3130 28460 3150
rect 28420 3100 28460 3130
rect 28420 3080 28430 3100
rect 28450 3080 28460 3100
rect 28420 3065 28460 3080
rect 28475 3650 28515 3665
rect 28475 3630 28485 3650
rect 28505 3630 28515 3650
rect 28475 3600 28515 3630
rect 28475 3580 28485 3600
rect 28505 3580 28515 3600
rect 28475 3550 28515 3580
rect 28475 3530 28485 3550
rect 28505 3530 28515 3550
rect 28475 3500 28515 3530
rect 28475 3480 28485 3500
rect 28505 3480 28515 3500
rect 28475 3450 28515 3480
rect 28475 3430 28485 3450
rect 28505 3430 28515 3450
rect 28475 3400 28515 3430
rect 28475 3380 28485 3400
rect 28505 3380 28515 3400
rect 28475 3350 28515 3380
rect 28475 3330 28485 3350
rect 28505 3330 28515 3350
rect 28475 3300 28515 3330
rect 28475 3280 28485 3300
rect 28505 3280 28515 3300
rect 28475 3250 28515 3280
rect 28475 3230 28485 3250
rect 28505 3230 28515 3250
rect 28475 3200 28515 3230
rect 28475 3180 28485 3200
rect 28505 3180 28515 3200
rect 28475 3150 28515 3180
rect 28475 3130 28485 3150
rect 28505 3130 28515 3150
rect 28475 3100 28515 3130
rect 28475 3080 28485 3100
rect 28505 3080 28515 3100
rect 28475 3065 28515 3080
rect 28530 3650 28570 3665
rect 28530 3630 28540 3650
rect 28560 3630 28570 3650
rect 28530 3600 28570 3630
rect 28530 3580 28540 3600
rect 28560 3580 28570 3600
rect 28530 3550 28570 3580
rect 28530 3530 28540 3550
rect 28560 3530 28570 3550
rect 28530 3500 28570 3530
rect 28530 3480 28540 3500
rect 28560 3480 28570 3500
rect 28530 3450 28570 3480
rect 28530 3430 28540 3450
rect 28560 3430 28570 3450
rect 28530 3400 28570 3430
rect 28530 3380 28540 3400
rect 28560 3380 28570 3400
rect 28530 3350 28570 3380
rect 28530 3330 28540 3350
rect 28560 3330 28570 3350
rect 28530 3300 28570 3330
rect 28530 3280 28540 3300
rect 28560 3280 28570 3300
rect 28530 3250 28570 3280
rect 28530 3230 28540 3250
rect 28560 3230 28570 3250
rect 28530 3200 28570 3230
rect 28530 3180 28540 3200
rect 28560 3180 28570 3200
rect 28530 3150 28570 3180
rect 28530 3130 28540 3150
rect 28560 3130 28570 3150
rect 28530 3100 28570 3130
rect 28530 3080 28540 3100
rect 28560 3080 28570 3100
rect 28530 3065 28570 3080
rect 28585 3650 28625 3665
rect 28585 3630 28595 3650
rect 28615 3630 28625 3650
rect 28585 3600 28625 3630
rect 28585 3580 28595 3600
rect 28615 3580 28625 3600
rect 28585 3550 28625 3580
rect 28585 3530 28595 3550
rect 28615 3530 28625 3550
rect 28585 3500 28625 3530
rect 28585 3480 28595 3500
rect 28615 3480 28625 3500
rect 28585 3450 28625 3480
rect 28585 3430 28595 3450
rect 28615 3430 28625 3450
rect 28585 3400 28625 3430
rect 28585 3380 28595 3400
rect 28615 3380 28625 3400
rect 28585 3350 28625 3380
rect 28585 3330 28595 3350
rect 28615 3330 28625 3350
rect 28585 3300 28625 3330
rect 28585 3280 28595 3300
rect 28615 3280 28625 3300
rect 28585 3250 28625 3280
rect 28585 3230 28595 3250
rect 28615 3230 28625 3250
rect 28585 3200 28625 3230
rect 28585 3180 28595 3200
rect 28615 3180 28625 3200
rect 28585 3150 28625 3180
rect 28585 3130 28595 3150
rect 28615 3130 28625 3150
rect 28585 3100 28625 3130
rect 28585 3080 28595 3100
rect 28615 3080 28625 3100
rect 28585 3065 28625 3080
rect 28640 3650 28680 3665
rect 28640 3630 28650 3650
rect 28670 3630 28680 3650
rect 28640 3600 28680 3630
rect 28640 3580 28650 3600
rect 28670 3580 28680 3600
rect 28640 3550 28680 3580
rect 28640 3530 28650 3550
rect 28670 3530 28680 3550
rect 28640 3500 28680 3530
rect 28640 3480 28650 3500
rect 28670 3480 28680 3500
rect 28640 3450 28680 3480
rect 28640 3430 28650 3450
rect 28670 3430 28680 3450
rect 28640 3400 28680 3430
rect 28640 3380 28650 3400
rect 28670 3380 28680 3400
rect 28640 3350 28680 3380
rect 28640 3330 28650 3350
rect 28670 3330 28680 3350
rect 28640 3300 28680 3330
rect 28640 3280 28650 3300
rect 28670 3280 28680 3300
rect 28640 3250 28680 3280
rect 28640 3230 28650 3250
rect 28670 3230 28680 3250
rect 28640 3200 28680 3230
rect 28640 3180 28650 3200
rect 28670 3180 28680 3200
rect 28640 3150 28680 3180
rect 28640 3130 28650 3150
rect 28670 3130 28680 3150
rect 28640 3100 28680 3130
rect 28640 3080 28650 3100
rect 28670 3080 28680 3100
rect 28640 3065 28680 3080
rect 28695 3650 28735 3665
rect 28695 3630 28705 3650
rect 28725 3630 28735 3650
rect 28695 3600 28735 3630
rect 28695 3580 28705 3600
rect 28725 3580 28735 3600
rect 28695 3550 28735 3580
rect 28695 3530 28705 3550
rect 28725 3530 28735 3550
rect 28695 3500 28735 3530
rect 28695 3480 28705 3500
rect 28725 3480 28735 3500
rect 28695 3450 28735 3480
rect 28695 3430 28705 3450
rect 28725 3430 28735 3450
rect 28695 3400 28735 3430
rect 28695 3380 28705 3400
rect 28725 3380 28735 3400
rect 28695 3350 28735 3380
rect 28695 3330 28705 3350
rect 28725 3330 28735 3350
rect 28695 3300 28735 3330
rect 28695 3280 28705 3300
rect 28725 3280 28735 3300
rect 28695 3250 28735 3280
rect 28695 3230 28705 3250
rect 28725 3230 28735 3250
rect 28695 3200 28735 3230
rect 28695 3180 28705 3200
rect 28725 3180 28735 3200
rect 28695 3150 28735 3180
rect 28695 3130 28705 3150
rect 28725 3130 28735 3150
rect 28695 3100 28735 3130
rect 28695 3080 28705 3100
rect 28725 3080 28735 3100
rect 28695 3065 28735 3080
rect 28750 3650 28790 3665
rect 28750 3630 28760 3650
rect 28780 3630 28790 3650
rect 28750 3600 28790 3630
rect 28750 3580 28760 3600
rect 28780 3580 28790 3600
rect 28750 3550 28790 3580
rect 28750 3530 28760 3550
rect 28780 3530 28790 3550
rect 28750 3500 28790 3530
rect 28750 3480 28760 3500
rect 28780 3480 28790 3500
rect 28750 3450 28790 3480
rect 28750 3430 28760 3450
rect 28780 3430 28790 3450
rect 28750 3400 28790 3430
rect 28750 3380 28760 3400
rect 28780 3380 28790 3400
rect 28750 3350 28790 3380
rect 28750 3330 28760 3350
rect 28780 3330 28790 3350
rect 28750 3300 28790 3330
rect 28750 3280 28760 3300
rect 28780 3280 28790 3300
rect 28750 3250 28790 3280
rect 28750 3230 28760 3250
rect 28780 3230 28790 3250
rect 28750 3200 28790 3230
rect 28750 3180 28760 3200
rect 28780 3180 28790 3200
rect 28750 3150 28790 3180
rect 28750 3130 28760 3150
rect 28780 3130 28790 3150
rect 28750 3100 28790 3130
rect 28750 3080 28760 3100
rect 28780 3080 28790 3100
rect 28750 3065 28790 3080
rect 28805 3650 28845 3665
rect 28805 3630 28815 3650
rect 28835 3630 28845 3650
rect 28805 3600 28845 3630
rect 28805 3580 28815 3600
rect 28835 3580 28845 3600
rect 28805 3550 28845 3580
rect 28805 3530 28815 3550
rect 28835 3530 28845 3550
rect 28805 3500 28845 3530
rect 28805 3480 28815 3500
rect 28835 3480 28845 3500
rect 28805 3450 28845 3480
rect 28805 3430 28815 3450
rect 28835 3430 28845 3450
rect 28805 3400 28845 3430
rect 28805 3380 28815 3400
rect 28835 3380 28845 3400
rect 28805 3350 28845 3380
rect 28805 3330 28815 3350
rect 28835 3330 28845 3350
rect 28805 3300 28845 3330
rect 28805 3280 28815 3300
rect 28835 3280 28845 3300
rect 28805 3250 28845 3280
rect 28805 3230 28815 3250
rect 28835 3230 28845 3250
rect 28805 3200 28845 3230
rect 28805 3180 28815 3200
rect 28835 3180 28845 3200
rect 28805 3150 28845 3180
rect 28805 3130 28815 3150
rect 28835 3130 28845 3150
rect 28805 3100 28845 3130
rect 28805 3080 28815 3100
rect 28835 3080 28845 3100
rect 28805 3065 28845 3080
rect 2995 2915 3035 2930
rect 2995 2895 3005 2915
rect 3025 2895 3035 2915
rect 2995 2865 3035 2895
rect 2995 2845 3005 2865
rect 3025 2845 3035 2865
rect 2995 2830 3035 2845
rect 3085 2915 3125 2930
rect 3085 2895 3095 2915
rect 3115 2895 3125 2915
rect 3085 2865 3125 2895
rect 3085 2845 3095 2865
rect 3115 2845 3125 2865
rect 3085 2830 3125 2845
rect 3175 2915 3215 2930
rect 3175 2895 3185 2915
rect 3205 2895 3215 2915
rect 3175 2865 3215 2895
rect 3175 2845 3185 2865
rect 3205 2845 3215 2865
rect 3175 2830 3215 2845
rect 3265 2915 3305 2930
rect 3265 2895 3275 2915
rect 3295 2895 3305 2915
rect 3265 2865 3305 2895
rect 3265 2845 3275 2865
rect 3295 2845 3305 2865
rect 3265 2830 3305 2845
rect 3355 2915 3395 2930
rect 3355 2895 3365 2915
rect 3385 2895 3395 2915
rect 3355 2865 3395 2895
rect 3355 2845 3365 2865
rect 3385 2845 3395 2865
rect 3355 2830 3395 2845
rect 3445 2915 3485 2930
rect 3445 2895 3455 2915
rect 3475 2895 3485 2915
rect 3445 2865 3485 2895
rect 3445 2845 3455 2865
rect 3475 2845 3485 2865
rect 3445 2830 3485 2845
rect 3535 2915 3575 2930
rect 3535 2895 3545 2915
rect 3565 2895 3575 2915
rect 3535 2865 3575 2895
rect 3535 2845 3545 2865
rect 3565 2845 3575 2865
rect 3535 2830 3575 2845
rect 3625 2915 3665 2930
rect 3625 2895 3635 2915
rect 3655 2895 3665 2915
rect 3625 2865 3665 2895
rect 3625 2845 3635 2865
rect 3655 2845 3665 2865
rect 3625 2830 3665 2845
rect 3715 2915 3755 2930
rect 3715 2895 3725 2915
rect 3745 2895 3755 2915
rect 3715 2865 3755 2895
rect 3715 2845 3725 2865
rect 3745 2845 3755 2865
rect 3715 2830 3755 2845
rect 3805 2915 3845 2930
rect 3805 2895 3815 2915
rect 3835 2895 3845 2915
rect 3805 2865 3845 2895
rect 3805 2845 3815 2865
rect 3835 2845 3845 2865
rect 3805 2830 3845 2845
rect 3895 2915 3935 2930
rect 3895 2895 3905 2915
rect 3925 2895 3935 2915
rect 3895 2865 3935 2895
rect 3895 2845 3905 2865
rect 3925 2845 3935 2865
rect 3895 2830 3935 2845
rect 3985 2915 4025 2930
rect 3985 2895 3995 2915
rect 4015 2895 4025 2915
rect 3985 2865 4025 2895
rect 3985 2845 3995 2865
rect 4015 2845 4025 2865
rect 3985 2830 4025 2845
rect 4075 2915 4115 2930
rect 4075 2895 4085 2915
rect 4105 2895 4115 2915
rect 4075 2865 4115 2895
rect 4075 2845 4085 2865
rect 4105 2845 4115 2865
rect 4075 2830 4115 2845
rect 4165 2915 4205 2930
rect 4165 2895 4175 2915
rect 4195 2895 4205 2915
rect 4165 2865 4205 2895
rect 4165 2845 4175 2865
rect 4195 2845 4205 2865
rect 4165 2830 4205 2845
rect 4255 2915 4295 2930
rect 4255 2895 4265 2915
rect 4285 2895 4295 2915
rect 4255 2865 4295 2895
rect 4255 2845 4265 2865
rect 4285 2845 4295 2865
rect 4255 2830 4295 2845
rect 4345 2915 4385 2930
rect 4345 2895 4355 2915
rect 4375 2895 4385 2915
rect 4345 2865 4385 2895
rect 4345 2845 4355 2865
rect 4375 2845 4385 2865
rect 4345 2830 4385 2845
rect 4435 2915 4475 2930
rect 4435 2895 4445 2915
rect 4465 2895 4475 2915
rect 4435 2865 4475 2895
rect 4435 2845 4445 2865
rect 4465 2845 4475 2865
rect 4435 2830 4475 2845
rect 4525 2915 4565 2930
rect 4525 2895 4535 2915
rect 4555 2895 4565 2915
rect 4525 2865 4565 2895
rect 4525 2845 4535 2865
rect 4555 2845 4565 2865
rect 4525 2830 4565 2845
rect 4615 2915 4655 2930
rect 4615 2895 4625 2915
rect 4645 2895 4655 2915
rect 4615 2865 4655 2895
rect 4615 2845 4625 2865
rect 4645 2845 4655 2865
rect 4615 2830 4655 2845
rect 4705 2915 4745 2930
rect 4705 2895 4715 2915
rect 4735 2895 4745 2915
rect 4705 2865 4745 2895
rect 4705 2845 4715 2865
rect 4735 2845 4745 2865
rect 4705 2830 4745 2845
rect 4795 2915 4835 2930
rect 4795 2895 4805 2915
rect 4825 2895 4835 2915
rect 4795 2865 4835 2895
rect 4795 2845 4805 2865
rect 4825 2845 4835 2865
rect 4795 2830 4835 2845
rect 4885 2915 4925 2930
rect 4885 2895 4895 2915
rect 4915 2895 4925 2915
rect 4885 2865 4925 2895
rect 4885 2845 4895 2865
rect 4915 2845 4925 2865
rect 4885 2830 4925 2845
rect 4975 2915 5015 2930
rect 4975 2895 4985 2915
rect 5005 2895 5015 2915
rect 4975 2865 5015 2895
rect 4975 2845 4985 2865
rect 5005 2845 5015 2865
rect 4975 2830 5015 2845
rect 16015 2830 16055 2845
rect 16015 2810 16025 2830
rect 16045 2810 16055 2830
rect 16015 2780 16055 2810
rect 16015 2760 16025 2780
rect 16045 2760 16055 2780
rect 16015 2730 16055 2760
rect 16015 2710 16025 2730
rect 16045 2710 16055 2730
rect 3175 2685 3215 2700
rect 3175 2665 3185 2685
rect 3205 2665 3215 2685
rect 3175 2635 3215 2665
rect 3175 2615 3185 2635
rect 3205 2615 3215 2635
rect 3175 2585 3215 2615
rect 3175 2565 3185 2585
rect 3205 2565 3215 2585
rect 3175 2535 3215 2565
rect 3175 2515 3185 2535
rect 3205 2515 3215 2535
rect 3175 2485 3215 2515
rect 3175 2465 3185 2485
rect 3205 2465 3215 2485
rect 3175 2435 3215 2465
rect 3175 2415 3185 2435
rect 3205 2415 3215 2435
rect 3175 2400 3215 2415
rect 3265 2685 3305 2700
rect 3265 2665 3275 2685
rect 3295 2665 3305 2685
rect 3265 2635 3305 2665
rect 3265 2615 3275 2635
rect 3295 2615 3305 2635
rect 3265 2585 3305 2615
rect 3265 2565 3275 2585
rect 3295 2565 3305 2585
rect 3265 2535 3305 2565
rect 3265 2515 3275 2535
rect 3295 2515 3305 2535
rect 3265 2485 3305 2515
rect 3265 2465 3275 2485
rect 3295 2465 3305 2485
rect 3265 2435 3305 2465
rect 3265 2415 3275 2435
rect 3295 2415 3305 2435
rect 3265 2400 3305 2415
rect 3355 2685 3395 2700
rect 3355 2665 3365 2685
rect 3385 2665 3395 2685
rect 3355 2635 3395 2665
rect 3355 2615 3365 2635
rect 3385 2615 3395 2635
rect 3355 2585 3395 2615
rect 3355 2565 3365 2585
rect 3385 2565 3395 2585
rect 3355 2535 3395 2565
rect 3355 2515 3365 2535
rect 3385 2515 3395 2535
rect 3355 2485 3395 2515
rect 3355 2465 3365 2485
rect 3385 2465 3395 2485
rect 3355 2435 3395 2465
rect 3355 2415 3365 2435
rect 3385 2415 3395 2435
rect 3355 2400 3395 2415
rect 3445 2685 3485 2700
rect 3445 2665 3455 2685
rect 3475 2665 3485 2685
rect 3445 2635 3485 2665
rect 3445 2615 3455 2635
rect 3475 2615 3485 2635
rect 3445 2585 3485 2615
rect 3445 2565 3455 2585
rect 3475 2565 3485 2585
rect 3445 2535 3485 2565
rect 3445 2515 3455 2535
rect 3475 2515 3485 2535
rect 3445 2485 3485 2515
rect 3445 2465 3455 2485
rect 3475 2465 3485 2485
rect 3445 2435 3485 2465
rect 3445 2415 3455 2435
rect 3475 2415 3485 2435
rect 3445 2400 3485 2415
rect 3535 2685 3575 2700
rect 3535 2665 3545 2685
rect 3565 2665 3575 2685
rect 3535 2635 3575 2665
rect 3535 2615 3545 2635
rect 3565 2615 3575 2635
rect 3535 2585 3575 2615
rect 3535 2565 3545 2585
rect 3565 2565 3575 2585
rect 3535 2535 3575 2565
rect 3535 2515 3545 2535
rect 3565 2515 3575 2535
rect 3535 2485 3575 2515
rect 3535 2465 3545 2485
rect 3565 2465 3575 2485
rect 3535 2435 3575 2465
rect 3535 2415 3545 2435
rect 3565 2415 3575 2435
rect 3535 2400 3575 2415
rect 3625 2685 3665 2700
rect 3625 2665 3635 2685
rect 3655 2665 3665 2685
rect 3625 2635 3665 2665
rect 3625 2615 3635 2635
rect 3655 2615 3665 2635
rect 3625 2585 3665 2615
rect 3625 2565 3635 2585
rect 3655 2565 3665 2585
rect 3625 2535 3665 2565
rect 3625 2515 3635 2535
rect 3655 2515 3665 2535
rect 3625 2485 3665 2515
rect 3625 2465 3635 2485
rect 3655 2465 3665 2485
rect 3625 2435 3665 2465
rect 3625 2415 3635 2435
rect 3655 2415 3665 2435
rect 3625 2400 3665 2415
rect 3715 2685 3755 2700
rect 3715 2665 3725 2685
rect 3745 2665 3755 2685
rect 3715 2635 3755 2665
rect 3715 2615 3725 2635
rect 3745 2615 3755 2635
rect 3715 2585 3755 2615
rect 3715 2565 3725 2585
rect 3745 2565 3755 2585
rect 3715 2535 3755 2565
rect 3715 2515 3725 2535
rect 3745 2515 3755 2535
rect 3715 2485 3755 2515
rect 3715 2465 3725 2485
rect 3745 2465 3755 2485
rect 3715 2435 3755 2465
rect 3715 2415 3725 2435
rect 3745 2415 3755 2435
rect 3715 2400 3755 2415
rect 3805 2685 3845 2700
rect 3805 2665 3815 2685
rect 3835 2665 3845 2685
rect 3805 2635 3845 2665
rect 3805 2615 3815 2635
rect 3835 2615 3845 2635
rect 3805 2585 3845 2615
rect 3805 2565 3815 2585
rect 3835 2565 3845 2585
rect 3805 2535 3845 2565
rect 3805 2515 3815 2535
rect 3835 2515 3845 2535
rect 3805 2485 3845 2515
rect 3805 2465 3815 2485
rect 3835 2465 3845 2485
rect 3805 2435 3845 2465
rect 3805 2415 3815 2435
rect 3835 2415 3845 2435
rect 3805 2400 3845 2415
rect 3895 2685 3935 2700
rect 3895 2665 3905 2685
rect 3925 2665 3935 2685
rect 3895 2635 3935 2665
rect 3895 2615 3905 2635
rect 3925 2615 3935 2635
rect 3895 2585 3935 2615
rect 3895 2565 3905 2585
rect 3925 2565 3935 2585
rect 3895 2535 3935 2565
rect 3895 2515 3905 2535
rect 3925 2515 3935 2535
rect 3895 2485 3935 2515
rect 3895 2465 3905 2485
rect 3925 2465 3935 2485
rect 3895 2435 3935 2465
rect 3895 2415 3905 2435
rect 3925 2415 3935 2435
rect 3895 2400 3935 2415
rect 3985 2685 4025 2700
rect 3985 2665 3995 2685
rect 4015 2665 4025 2685
rect 3985 2635 4025 2665
rect 3985 2615 3995 2635
rect 4015 2615 4025 2635
rect 3985 2585 4025 2615
rect 3985 2565 3995 2585
rect 4015 2565 4025 2585
rect 3985 2535 4025 2565
rect 3985 2515 3995 2535
rect 4015 2515 4025 2535
rect 3985 2485 4025 2515
rect 3985 2465 3995 2485
rect 4015 2465 4025 2485
rect 3985 2435 4025 2465
rect 3985 2415 3995 2435
rect 4015 2415 4025 2435
rect 3985 2400 4025 2415
rect 4075 2685 4115 2700
rect 4075 2665 4085 2685
rect 4105 2665 4115 2685
rect 4075 2635 4115 2665
rect 4075 2615 4085 2635
rect 4105 2615 4115 2635
rect 4075 2585 4115 2615
rect 4075 2565 4085 2585
rect 4105 2565 4115 2585
rect 4075 2535 4115 2565
rect 4075 2515 4085 2535
rect 4105 2515 4115 2535
rect 4075 2485 4115 2515
rect 4075 2465 4085 2485
rect 4105 2465 4115 2485
rect 4075 2435 4115 2465
rect 4075 2415 4085 2435
rect 4105 2415 4115 2435
rect 4075 2400 4115 2415
rect 4165 2685 4205 2700
rect 4165 2665 4175 2685
rect 4195 2665 4205 2685
rect 4165 2635 4205 2665
rect 4165 2615 4175 2635
rect 4195 2615 4205 2635
rect 4165 2585 4205 2615
rect 4165 2565 4175 2585
rect 4195 2565 4205 2585
rect 4165 2535 4205 2565
rect 4165 2515 4175 2535
rect 4195 2515 4205 2535
rect 4165 2485 4205 2515
rect 4165 2465 4175 2485
rect 4195 2465 4205 2485
rect 4165 2435 4205 2465
rect 4165 2415 4175 2435
rect 4195 2415 4205 2435
rect 4165 2400 4205 2415
rect 4255 2685 4295 2700
rect 4255 2665 4265 2685
rect 4285 2665 4295 2685
rect 4255 2635 4295 2665
rect 4255 2615 4265 2635
rect 4285 2615 4295 2635
rect 4255 2585 4295 2615
rect 4255 2565 4265 2585
rect 4285 2565 4295 2585
rect 4255 2535 4295 2565
rect 4255 2515 4265 2535
rect 4285 2515 4295 2535
rect 4255 2485 4295 2515
rect 4255 2465 4265 2485
rect 4285 2465 4295 2485
rect 4255 2435 4295 2465
rect 4255 2415 4265 2435
rect 4285 2415 4295 2435
rect 4255 2400 4295 2415
rect 4345 2685 4385 2700
rect 4345 2665 4355 2685
rect 4375 2665 4385 2685
rect 4345 2635 4385 2665
rect 4345 2615 4355 2635
rect 4375 2615 4385 2635
rect 4345 2585 4385 2615
rect 4345 2565 4355 2585
rect 4375 2565 4385 2585
rect 4345 2535 4385 2565
rect 4345 2515 4355 2535
rect 4375 2515 4385 2535
rect 4345 2485 4385 2515
rect 4345 2465 4355 2485
rect 4375 2465 4385 2485
rect 4345 2435 4385 2465
rect 4345 2415 4355 2435
rect 4375 2415 4385 2435
rect 4345 2400 4385 2415
rect 4435 2685 4475 2700
rect 4435 2665 4445 2685
rect 4465 2665 4475 2685
rect 4435 2635 4475 2665
rect 4435 2615 4445 2635
rect 4465 2615 4475 2635
rect 4435 2585 4475 2615
rect 4435 2565 4445 2585
rect 4465 2565 4475 2585
rect 4435 2535 4475 2565
rect 4435 2515 4445 2535
rect 4465 2515 4475 2535
rect 4435 2485 4475 2515
rect 4435 2465 4445 2485
rect 4465 2465 4475 2485
rect 4435 2435 4475 2465
rect 4435 2415 4445 2435
rect 4465 2415 4475 2435
rect 4435 2400 4475 2415
rect 4525 2685 4565 2700
rect 4525 2665 4535 2685
rect 4555 2665 4565 2685
rect 4525 2635 4565 2665
rect 4525 2615 4535 2635
rect 4555 2615 4565 2635
rect 4525 2585 4565 2615
rect 4525 2565 4535 2585
rect 4555 2565 4565 2585
rect 4525 2535 4565 2565
rect 4525 2515 4535 2535
rect 4555 2515 4565 2535
rect 4525 2485 4565 2515
rect 4525 2465 4535 2485
rect 4555 2465 4565 2485
rect 4525 2435 4565 2465
rect 4525 2415 4535 2435
rect 4555 2415 4565 2435
rect 4525 2400 4565 2415
rect 4615 2685 4655 2700
rect 4615 2665 4625 2685
rect 4645 2665 4655 2685
rect 4615 2635 4655 2665
rect 4615 2615 4625 2635
rect 4645 2615 4655 2635
rect 4615 2585 4655 2615
rect 4615 2565 4625 2585
rect 4645 2565 4655 2585
rect 4615 2535 4655 2565
rect 4615 2515 4625 2535
rect 4645 2515 4655 2535
rect 4615 2485 4655 2515
rect 4615 2465 4625 2485
rect 4645 2465 4655 2485
rect 4615 2435 4655 2465
rect 4615 2415 4625 2435
rect 4645 2415 4655 2435
rect 4615 2400 4655 2415
rect 4705 2685 4745 2700
rect 4705 2665 4715 2685
rect 4735 2665 4745 2685
rect 4705 2635 4745 2665
rect 4705 2615 4715 2635
rect 4735 2615 4745 2635
rect 4705 2585 4745 2615
rect 4705 2565 4715 2585
rect 4735 2565 4745 2585
rect 4705 2535 4745 2565
rect 4705 2515 4715 2535
rect 4735 2515 4745 2535
rect 4705 2485 4745 2515
rect 4705 2465 4715 2485
rect 4735 2465 4745 2485
rect 4705 2435 4745 2465
rect 4705 2415 4715 2435
rect 4735 2415 4745 2435
rect 4705 2400 4745 2415
rect 4795 2685 4835 2700
rect 4795 2665 4805 2685
rect 4825 2665 4835 2685
rect 16015 2680 16055 2710
rect 4795 2635 4835 2665
rect 16015 2660 16025 2680
rect 16045 2660 16055 2680
rect 4795 2615 4805 2635
rect 4825 2615 4835 2635
rect 15005 2640 15045 2655
rect 4795 2585 4835 2615
rect 4795 2565 4805 2585
rect 4825 2565 4835 2585
rect 4795 2535 4835 2565
rect 4795 2515 4805 2535
rect 4825 2515 4835 2535
rect 4795 2485 4835 2515
rect 4795 2465 4805 2485
rect 4825 2465 4835 2485
rect 4795 2435 4835 2465
rect 4795 2415 4805 2435
rect 4825 2415 4835 2435
rect 4795 2400 4835 2415
rect 15005 2620 15015 2640
rect 15035 2620 15045 2640
rect 15005 2590 15045 2620
rect 15005 2570 15015 2590
rect 15035 2570 15045 2590
rect 15005 2540 15045 2570
rect 15005 2520 15015 2540
rect 15035 2520 15045 2540
rect 15005 2490 15045 2520
rect 15005 2470 15015 2490
rect 15035 2470 15045 2490
rect 15005 2455 15045 2470
rect 15060 2640 15100 2655
rect 15060 2620 15070 2640
rect 15090 2620 15100 2640
rect 15060 2590 15100 2620
rect 15060 2570 15070 2590
rect 15090 2570 15100 2590
rect 15060 2540 15100 2570
rect 15060 2520 15070 2540
rect 15090 2520 15100 2540
rect 15060 2490 15100 2520
rect 15060 2470 15070 2490
rect 15090 2470 15100 2490
rect 15060 2455 15100 2470
rect 15115 2640 15155 2655
rect 15115 2620 15125 2640
rect 15145 2620 15155 2640
rect 15115 2590 15155 2620
rect 15115 2570 15125 2590
rect 15145 2570 15155 2590
rect 15115 2540 15155 2570
rect 15115 2520 15125 2540
rect 15145 2520 15155 2540
rect 15115 2490 15155 2520
rect 15115 2470 15125 2490
rect 15145 2470 15155 2490
rect 15115 2455 15155 2470
rect 15170 2640 15210 2655
rect 15170 2620 15180 2640
rect 15200 2620 15210 2640
rect 15170 2590 15210 2620
rect 15170 2570 15180 2590
rect 15200 2570 15210 2590
rect 15170 2540 15210 2570
rect 15170 2520 15180 2540
rect 15200 2520 15210 2540
rect 15170 2490 15210 2520
rect 15170 2470 15180 2490
rect 15200 2470 15210 2490
rect 15170 2455 15210 2470
rect 15225 2640 15265 2655
rect 15225 2620 15235 2640
rect 15255 2620 15265 2640
rect 15225 2590 15265 2620
rect 15225 2570 15235 2590
rect 15255 2570 15265 2590
rect 15225 2540 15265 2570
rect 15225 2520 15235 2540
rect 15255 2520 15265 2540
rect 15225 2490 15265 2520
rect 15225 2470 15235 2490
rect 15255 2470 15265 2490
rect 15225 2455 15265 2470
rect 15280 2640 15320 2655
rect 15280 2620 15290 2640
rect 15310 2620 15320 2640
rect 15280 2590 15320 2620
rect 15280 2570 15290 2590
rect 15310 2570 15320 2590
rect 15280 2540 15320 2570
rect 15280 2520 15290 2540
rect 15310 2520 15320 2540
rect 15280 2490 15320 2520
rect 15280 2470 15290 2490
rect 15310 2470 15320 2490
rect 15280 2455 15320 2470
rect 15335 2640 15375 2655
rect 15335 2620 15345 2640
rect 15365 2620 15375 2640
rect 15335 2590 15375 2620
rect 15335 2570 15345 2590
rect 15365 2570 15375 2590
rect 15335 2540 15375 2570
rect 15335 2520 15345 2540
rect 15365 2520 15375 2540
rect 15335 2490 15375 2520
rect 15335 2470 15345 2490
rect 15365 2470 15375 2490
rect 15335 2455 15375 2470
rect 15390 2640 15430 2655
rect 15390 2620 15400 2640
rect 15420 2620 15430 2640
rect 15390 2590 15430 2620
rect 15390 2570 15400 2590
rect 15420 2570 15430 2590
rect 15390 2540 15430 2570
rect 15390 2520 15400 2540
rect 15420 2520 15430 2540
rect 15390 2490 15430 2520
rect 15390 2470 15400 2490
rect 15420 2470 15430 2490
rect 15390 2455 15430 2470
rect 15445 2640 15485 2655
rect 15445 2620 15455 2640
rect 15475 2620 15485 2640
rect 15445 2590 15485 2620
rect 15445 2570 15455 2590
rect 15475 2570 15485 2590
rect 15445 2540 15485 2570
rect 15445 2520 15455 2540
rect 15475 2520 15485 2540
rect 15445 2490 15485 2520
rect 15445 2470 15455 2490
rect 15475 2470 15485 2490
rect 15445 2455 15485 2470
rect 15500 2640 15540 2655
rect 15500 2620 15510 2640
rect 15530 2620 15540 2640
rect 15500 2590 15540 2620
rect 15500 2570 15510 2590
rect 15530 2570 15540 2590
rect 15500 2540 15540 2570
rect 15500 2520 15510 2540
rect 15530 2520 15540 2540
rect 15500 2490 15540 2520
rect 15500 2470 15510 2490
rect 15530 2470 15540 2490
rect 15500 2455 15540 2470
rect 15555 2640 15595 2655
rect 15555 2620 15565 2640
rect 15585 2620 15595 2640
rect 15555 2590 15595 2620
rect 15555 2570 15565 2590
rect 15585 2570 15595 2590
rect 15555 2540 15595 2570
rect 15555 2520 15565 2540
rect 15585 2520 15595 2540
rect 15555 2490 15595 2520
rect 15555 2470 15565 2490
rect 15585 2470 15595 2490
rect 15555 2455 15595 2470
rect 15610 2640 15650 2655
rect 15610 2620 15620 2640
rect 15640 2620 15650 2640
rect 15610 2590 15650 2620
rect 15610 2570 15620 2590
rect 15640 2570 15650 2590
rect 15610 2540 15650 2570
rect 15610 2520 15620 2540
rect 15640 2520 15650 2540
rect 15610 2490 15650 2520
rect 15610 2470 15620 2490
rect 15640 2470 15650 2490
rect 15610 2455 15650 2470
rect 15665 2640 15705 2655
rect 15665 2620 15675 2640
rect 15695 2620 15705 2640
rect 15665 2590 15705 2620
rect 15665 2570 15675 2590
rect 15695 2570 15705 2590
rect 15665 2540 15705 2570
rect 15665 2520 15675 2540
rect 15695 2520 15705 2540
rect 15665 2490 15705 2520
rect 16015 2630 16055 2660
rect 16015 2610 16025 2630
rect 16045 2610 16055 2630
rect 16015 2580 16055 2610
rect 16015 2560 16025 2580
rect 16045 2560 16055 2580
rect 16015 2530 16055 2560
rect 16015 2510 16025 2530
rect 16045 2510 16055 2530
rect 16015 2495 16055 2510
rect 16075 2830 16115 2845
rect 16075 2810 16085 2830
rect 16105 2810 16115 2830
rect 16075 2780 16115 2810
rect 16075 2760 16085 2780
rect 16105 2760 16115 2780
rect 16075 2730 16115 2760
rect 16075 2710 16085 2730
rect 16105 2710 16115 2730
rect 16075 2680 16115 2710
rect 16075 2660 16085 2680
rect 16105 2660 16115 2680
rect 16075 2630 16115 2660
rect 16075 2610 16085 2630
rect 16105 2610 16115 2630
rect 16075 2580 16115 2610
rect 16075 2560 16085 2580
rect 16105 2560 16115 2580
rect 16075 2530 16115 2560
rect 16075 2510 16085 2530
rect 16105 2510 16115 2530
rect 16075 2495 16115 2510
rect 16135 2830 16175 2845
rect 16135 2810 16145 2830
rect 16165 2810 16175 2830
rect 16135 2780 16175 2810
rect 16135 2760 16145 2780
rect 16165 2760 16175 2780
rect 16135 2730 16175 2760
rect 16135 2710 16145 2730
rect 16165 2710 16175 2730
rect 16135 2680 16175 2710
rect 16135 2660 16145 2680
rect 16165 2660 16175 2680
rect 16135 2630 16175 2660
rect 16135 2610 16145 2630
rect 16165 2610 16175 2630
rect 16135 2580 16175 2610
rect 16135 2560 16145 2580
rect 16165 2560 16175 2580
rect 16135 2530 16175 2560
rect 16135 2510 16145 2530
rect 16165 2510 16175 2530
rect 16135 2495 16175 2510
rect 16195 2830 16235 2845
rect 16195 2810 16205 2830
rect 16225 2810 16235 2830
rect 16195 2780 16235 2810
rect 16195 2760 16205 2780
rect 16225 2760 16235 2780
rect 16195 2730 16235 2760
rect 16195 2710 16205 2730
rect 16225 2710 16235 2730
rect 16195 2680 16235 2710
rect 16195 2660 16205 2680
rect 16225 2660 16235 2680
rect 16195 2630 16235 2660
rect 16195 2610 16205 2630
rect 16225 2610 16235 2630
rect 16195 2580 16235 2610
rect 16195 2560 16205 2580
rect 16225 2560 16235 2580
rect 16195 2530 16235 2560
rect 16195 2510 16205 2530
rect 16225 2510 16235 2530
rect 16195 2495 16235 2510
rect 16255 2830 16295 2845
rect 16255 2810 16265 2830
rect 16285 2810 16295 2830
rect 16255 2780 16295 2810
rect 16255 2760 16265 2780
rect 16285 2760 16295 2780
rect 16255 2730 16295 2760
rect 16255 2710 16265 2730
rect 16285 2710 16295 2730
rect 16255 2680 16295 2710
rect 16255 2660 16265 2680
rect 16285 2660 16295 2680
rect 16255 2630 16295 2660
rect 16255 2610 16265 2630
rect 16285 2610 16295 2630
rect 16255 2580 16295 2610
rect 16255 2560 16265 2580
rect 16285 2560 16295 2580
rect 16255 2530 16295 2560
rect 16255 2510 16265 2530
rect 16285 2510 16295 2530
rect 16255 2495 16295 2510
rect 16315 2830 16355 2845
rect 16315 2810 16325 2830
rect 16345 2810 16355 2830
rect 16315 2780 16355 2810
rect 16315 2760 16325 2780
rect 16345 2760 16355 2780
rect 16315 2730 16355 2760
rect 16315 2710 16325 2730
rect 16345 2710 16355 2730
rect 16315 2680 16355 2710
rect 16315 2660 16325 2680
rect 16345 2660 16355 2680
rect 16315 2630 16355 2660
rect 16315 2610 16325 2630
rect 16345 2610 16355 2630
rect 16315 2580 16355 2610
rect 16315 2560 16325 2580
rect 16345 2560 16355 2580
rect 16315 2530 16355 2560
rect 16315 2510 16325 2530
rect 16345 2510 16355 2530
rect 16315 2495 16355 2510
rect 16375 2830 16415 2845
rect 16375 2810 16385 2830
rect 16405 2810 16415 2830
rect 16375 2780 16415 2810
rect 16375 2760 16385 2780
rect 16405 2760 16415 2780
rect 16375 2730 16415 2760
rect 16375 2710 16385 2730
rect 16405 2710 16415 2730
rect 16375 2680 16415 2710
rect 16375 2660 16385 2680
rect 16405 2660 16415 2680
rect 16375 2630 16415 2660
rect 16375 2610 16385 2630
rect 16405 2610 16415 2630
rect 16375 2580 16415 2610
rect 16375 2560 16385 2580
rect 16405 2560 16415 2580
rect 16375 2530 16415 2560
rect 16375 2510 16385 2530
rect 16405 2510 16415 2530
rect 16375 2495 16415 2510
rect 16435 2830 16475 2845
rect 16435 2810 16445 2830
rect 16465 2810 16475 2830
rect 16435 2780 16475 2810
rect 16435 2760 16445 2780
rect 16465 2760 16475 2780
rect 16435 2730 16475 2760
rect 16435 2710 16445 2730
rect 16465 2710 16475 2730
rect 16435 2680 16475 2710
rect 16435 2660 16445 2680
rect 16465 2660 16475 2680
rect 16435 2630 16475 2660
rect 16435 2610 16445 2630
rect 16465 2610 16475 2630
rect 16435 2580 16475 2610
rect 16435 2560 16445 2580
rect 16465 2560 16475 2580
rect 16435 2530 16475 2560
rect 16435 2510 16445 2530
rect 16465 2510 16475 2530
rect 16435 2495 16475 2510
rect 16495 2830 16535 2845
rect 16495 2810 16505 2830
rect 16525 2810 16535 2830
rect 16495 2780 16535 2810
rect 16495 2760 16505 2780
rect 16525 2760 16535 2780
rect 16495 2730 16535 2760
rect 16495 2710 16505 2730
rect 16525 2710 16535 2730
rect 16495 2680 16535 2710
rect 16495 2660 16505 2680
rect 16525 2660 16535 2680
rect 16495 2630 16535 2660
rect 16495 2610 16505 2630
rect 16525 2610 16535 2630
rect 16495 2580 16535 2610
rect 16495 2560 16505 2580
rect 16525 2560 16535 2580
rect 16495 2530 16535 2560
rect 16495 2510 16505 2530
rect 16525 2510 16535 2530
rect 16495 2495 16535 2510
rect 16555 2830 16595 2845
rect 16555 2810 16565 2830
rect 16585 2810 16595 2830
rect 16555 2780 16595 2810
rect 16555 2760 16565 2780
rect 16585 2760 16595 2780
rect 16555 2730 16595 2760
rect 16555 2710 16565 2730
rect 16585 2710 16595 2730
rect 16555 2680 16595 2710
rect 16555 2660 16565 2680
rect 16585 2660 16595 2680
rect 16555 2630 16595 2660
rect 16555 2610 16565 2630
rect 16585 2610 16595 2630
rect 16555 2580 16595 2610
rect 16555 2560 16565 2580
rect 16585 2560 16595 2580
rect 16555 2530 16595 2560
rect 16555 2510 16565 2530
rect 16585 2510 16595 2530
rect 16555 2495 16595 2510
rect 16615 2830 16655 2845
rect 16615 2810 16625 2830
rect 16645 2810 16655 2830
rect 16615 2780 16655 2810
rect 16615 2760 16625 2780
rect 16645 2760 16655 2780
rect 16615 2730 16655 2760
rect 16615 2710 16625 2730
rect 16645 2710 16655 2730
rect 16615 2680 16655 2710
rect 16615 2660 16625 2680
rect 16645 2660 16655 2680
rect 16615 2630 16655 2660
rect 16615 2610 16625 2630
rect 16645 2610 16655 2630
rect 16615 2580 16655 2610
rect 16615 2560 16625 2580
rect 16645 2560 16655 2580
rect 16615 2530 16655 2560
rect 16615 2510 16625 2530
rect 16645 2510 16655 2530
rect 16615 2495 16655 2510
rect 16675 2830 16715 2845
rect 16675 2810 16685 2830
rect 16705 2810 16715 2830
rect 16675 2780 16715 2810
rect 16675 2760 16685 2780
rect 16705 2760 16715 2780
rect 16675 2730 16715 2760
rect 16675 2710 16685 2730
rect 16705 2710 16715 2730
rect 16675 2680 16715 2710
rect 16675 2660 16685 2680
rect 16705 2660 16715 2680
rect 16675 2630 16715 2660
rect 16675 2610 16685 2630
rect 16705 2610 16715 2630
rect 16675 2580 16715 2610
rect 16675 2560 16685 2580
rect 16705 2560 16715 2580
rect 16675 2530 16715 2560
rect 16675 2510 16685 2530
rect 16705 2510 16715 2530
rect 16675 2495 16715 2510
rect 16735 2830 16775 2845
rect 16735 2810 16745 2830
rect 16765 2810 16775 2830
rect 16735 2780 16775 2810
rect 16735 2760 16745 2780
rect 16765 2760 16775 2780
rect 16735 2730 16775 2760
rect 16735 2710 16745 2730
rect 16765 2710 16775 2730
rect 16735 2680 16775 2710
rect 16735 2660 16745 2680
rect 16765 2660 16775 2680
rect 16735 2630 16775 2660
rect 16735 2610 16745 2630
rect 16765 2610 16775 2630
rect 16735 2580 16775 2610
rect 16735 2560 16745 2580
rect 16765 2560 16775 2580
rect 16735 2530 16775 2560
rect 16735 2510 16745 2530
rect 16765 2510 16775 2530
rect 16735 2495 16775 2510
rect 17025 2830 17065 2845
rect 17025 2810 17035 2830
rect 17055 2810 17065 2830
rect 17025 2780 17065 2810
rect 17025 2760 17035 2780
rect 17055 2760 17065 2780
rect 17025 2730 17065 2760
rect 17025 2710 17035 2730
rect 17055 2710 17065 2730
rect 17025 2680 17065 2710
rect 17025 2660 17035 2680
rect 17055 2660 17065 2680
rect 17025 2630 17065 2660
rect 17025 2610 17035 2630
rect 17055 2610 17065 2630
rect 17025 2580 17065 2610
rect 17025 2560 17035 2580
rect 17055 2560 17065 2580
rect 17025 2530 17065 2560
rect 17025 2510 17035 2530
rect 17055 2510 17065 2530
rect 17025 2495 17065 2510
rect 17085 2830 17125 2845
rect 17085 2810 17095 2830
rect 17115 2810 17125 2830
rect 17085 2780 17125 2810
rect 17085 2760 17095 2780
rect 17115 2760 17125 2780
rect 17085 2730 17125 2760
rect 17085 2710 17095 2730
rect 17115 2710 17125 2730
rect 17085 2680 17125 2710
rect 17085 2660 17095 2680
rect 17115 2660 17125 2680
rect 17085 2630 17125 2660
rect 17085 2610 17095 2630
rect 17115 2610 17125 2630
rect 17085 2580 17125 2610
rect 17085 2560 17095 2580
rect 17115 2560 17125 2580
rect 17085 2530 17125 2560
rect 17085 2510 17095 2530
rect 17115 2510 17125 2530
rect 17085 2495 17125 2510
rect 17145 2830 17185 2845
rect 17145 2810 17155 2830
rect 17175 2810 17185 2830
rect 17145 2780 17185 2810
rect 17145 2760 17155 2780
rect 17175 2760 17185 2780
rect 17145 2730 17185 2760
rect 17145 2710 17155 2730
rect 17175 2710 17185 2730
rect 17145 2680 17185 2710
rect 17145 2660 17155 2680
rect 17175 2660 17185 2680
rect 17145 2630 17185 2660
rect 17145 2610 17155 2630
rect 17175 2610 17185 2630
rect 17145 2580 17185 2610
rect 17145 2560 17155 2580
rect 17175 2560 17185 2580
rect 17145 2530 17185 2560
rect 17145 2510 17155 2530
rect 17175 2510 17185 2530
rect 17145 2495 17185 2510
rect 17205 2830 17245 2845
rect 17205 2810 17215 2830
rect 17235 2810 17245 2830
rect 17205 2780 17245 2810
rect 17205 2760 17215 2780
rect 17235 2760 17245 2780
rect 17205 2730 17245 2760
rect 17205 2710 17215 2730
rect 17235 2710 17245 2730
rect 17205 2680 17245 2710
rect 17205 2660 17215 2680
rect 17235 2660 17245 2680
rect 17205 2630 17245 2660
rect 17205 2610 17215 2630
rect 17235 2610 17245 2630
rect 17205 2580 17245 2610
rect 17205 2560 17215 2580
rect 17235 2560 17245 2580
rect 17205 2530 17245 2560
rect 17205 2510 17215 2530
rect 17235 2510 17245 2530
rect 17205 2495 17245 2510
rect 17265 2830 17305 2845
rect 17265 2810 17275 2830
rect 17295 2810 17305 2830
rect 17265 2780 17305 2810
rect 17265 2760 17275 2780
rect 17295 2760 17305 2780
rect 17265 2730 17305 2760
rect 17265 2710 17275 2730
rect 17295 2710 17305 2730
rect 17265 2680 17305 2710
rect 17265 2660 17275 2680
rect 17295 2660 17305 2680
rect 17265 2630 17305 2660
rect 17265 2610 17275 2630
rect 17295 2610 17305 2630
rect 17265 2580 17305 2610
rect 17265 2560 17275 2580
rect 17295 2560 17305 2580
rect 17265 2530 17305 2560
rect 17265 2510 17275 2530
rect 17295 2510 17305 2530
rect 17265 2495 17305 2510
rect 17325 2830 17365 2845
rect 17325 2810 17335 2830
rect 17355 2810 17365 2830
rect 17325 2780 17365 2810
rect 17325 2760 17335 2780
rect 17355 2760 17365 2780
rect 17325 2730 17365 2760
rect 17325 2710 17335 2730
rect 17355 2710 17365 2730
rect 17325 2680 17365 2710
rect 17325 2660 17335 2680
rect 17355 2660 17365 2680
rect 17325 2630 17365 2660
rect 17325 2610 17335 2630
rect 17355 2610 17365 2630
rect 17325 2580 17365 2610
rect 17325 2560 17335 2580
rect 17355 2560 17365 2580
rect 17325 2530 17365 2560
rect 17325 2510 17335 2530
rect 17355 2510 17365 2530
rect 17325 2495 17365 2510
rect 17385 2830 17425 2845
rect 17385 2810 17395 2830
rect 17415 2810 17425 2830
rect 17385 2780 17425 2810
rect 17385 2760 17395 2780
rect 17415 2760 17425 2780
rect 17385 2730 17425 2760
rect 17385 2710 17395 2730
rect 17415 2710 17425 2730
rect 17385 2680 17425 2710
rect 17385 2660 17395 2680
rect 17415 2660 17425 2680
rect 17385 2630 17425 2660
rect 17385 2610 17395 2630
rect 17415 2610 17425 2630
rect 17385 2580 17425 2610
rect 17385 2560 17395 2580
rect 17415 2560 17425 2580
rect 17385 2530 17425 2560
rect 17385 2510 17395 2530
rect 17415 2510 17425 2530
rect 17385 2495 17425 2510
rect 17445 2830 17485 2845
rect 17445 2810 17455 2830
rect 17475 2810 17485 2830
rect 17445 2780 17485 2810
rect 17445 2760 17455 2780
rect 17475 2760 17485 2780
rect 17445 2730 17485 2760
rect 17445 2710 17455 2730
rect 17475 2710 17485 2730
rect 17445 2680 17485 2710
rect 17445 2660 17455 2680
rect 17475 2660 17485 2680
rect 17445 2630 17485 2660
rect 17445 2610 17455 2630
rect 17475 2610 17485 2630
rect 17445 2580 17485 2610
rect 17445 2560 17455 2580
rect 17475 2560 17485 2580
rect 17445 2530 17485 2560
rect 17445 2510 17455 2530
rect 17475 2510 17485 2530
rect 17445 2495 17485 2510
rect 17505 2830 17545 2845
rect 17505 2810 17515 2830
rect 17535 2810 17545 2830
rect 17505 2780 17545 2810
rect 17505 2760 17515 2780
rect 17535 2760 17545 2780
rect 17505 2730 17545 2760
rect 17505 2710 17515 2730
rect 17535 2710 17545 2730
rect 17505 2680 17545 2710
rect 17505 2660 17515 2680
rect 17535 2660 17545 2680
rect 17505 2630 17545 2660
rect 17505 2610 17515 2630
rect 17535 2610 17545 2630
rect 17505 2580 17545 2610
rect 17505 2560 17515 2580
rect 17535 2560 17545 2580
rect 17505 2530 17545 2560
rect 17505 2510 17515 2530
rect 17535 2510 17545 2530
rect 17505 2495 17545 2510
rect 17565 2830 17605 2845
rect 17565 2810 17575 2830
rect 17595 2810 17605 2830
rect 17565 2780 17605 2810
rect 17565 2760 17575 2780
rect 17595 2760 17605 2780
rect 17565 2730 17605 2760
rect 17565 2710 17575 2730
rect 17595 2710 17605 2730
rect 17565 2680 17605 2710
rect 17565 2660 17575 2680
rect 17595 2660 17605 2680
rect 17565 2630 17605 2660
rect 17565 2610 17575 2630
rect 17595 2610 17605 2630
rect 17565 2580 17605 2610
rect 17565 2560 17575 2580
rect 17595 2560 17605 2580
rect 17565 2530 17605 2560
rect 17565 2510 17575 2530
rect 17595 2510 17605 2530
rect 17565 2495 17605 2510
rect 17625 2830 17665 2845
rect 17625 2810 17635 2830
rect 17655 2810 17665 2830
rect 17625 2780 17665 2810
rect 17625 2760 17635 2780
rect 17655 2760 17665 2780
rect 17625 2730 17665 2760
rect 17625 2710 17635 2730
rect 17655 2710 17665 2730
rect 17625 2680 17665 2710
rect 17625 2660 17635 2680
rect 17655 2660 17665 2680
rect 17625 2630 17665 2660
rect 17625 2610 17635 2630
rect 17655 2610 17665 2630
rect 17625 2580 17665 2610
rect 17625 2560 17635 2580
rect 17655 2560 17665 2580
rect 17625 2530 17665 2560
rect 17625 2510 17635 2530
rect 17655 2510 17665 2530
rect 17625 2495 17665 2510
rect 17685 2830 17725 2845
rect 17685 2810 17695 2830
rect 17715 2810 17725 2830
rect 17685 2780 17725 2810
rect 17685 2760 17695 2780
rect 17715 2760 17725 2780
rect 17685 2730 17725 2760
rect 17685 2710 17695 2730
rect 17715 2710 17725 2730
rect 17685 2680 17725 2710
rect 17685 2660 17695 2680
rect 17715 2660 17725 2680
rect 17685 2630 17725 2660
rect 17685 2610 17695 2630
rect 17715 2610 17725 2630
rect 17685 2580 17725 2610
rect 17685 2560 17695 2580
rect 17715 2560 17725 2580
rect 17685 2530 17725 2560
rect 17685 2510 17695 2530
rect 17715 2510 17725 2530
rect 17685 2495 17725 2510
rect 17745 2830 17785 2845
rect 17745 2810 17755 2830
rect 17775 2810 17785 2830
rect 17745 2780 17785 2810
rect 17745 2760 17755 2780
rect 17775 2760 17785 2780
rect 17745 2730 17785 2760
rect 17745 2710 17755 2730
rect 17775 2710 17785 2730
rect 17745 2680 17785 2710
rect 17745 2660 17755 2680
rect 17775 2660 17785 2680
rect 26015 2830 26055 2845
rect 26015 2810 26025 2830
rect 26045 2810 26055 2830
rect 26015 2780 26055 2810
rect 26015 2760 26025 2780
rect 26045 2760 26055 2780
rect 26015 2730 26055 2760
rect 26015 2710 26025 2730
rect 26045 2710 26055 2730
rect 26015 2680 26055 2710
rect 17745 2630 17785 2660
rect 26015 2660 26025 2680
rect 26045 2660 26055 2680
rect 17745 2610 17755 2630
rect 17775 2610 17785 2630
rect 17745 2580 17785 2610
rect 17745 2560 17755 2580
rect 17775 2560 17785 2580
rect 17745 2530 17785 2560
rect 17745 2510 17755 2530
rect 17775 2510 17785 2530
rect 17745 2495 17785 2510
rect 18145 2640 18185 2655
rect 18145 2620 18155 2640
rect 18175 2620 18185 2640
rect 18145 2590 18185 2620
rect 18145 2570 18155 2590
rect 18175 2570 18185 2590
rect 18145 2540 18185 2570
rect 18145 2520 18155 2540
rect 18175 2520 18185 2540
rect 15665 2470 15675 2490
rect 15695 2470 15705 2490
rect 18145 2490 18185 2520
rect 18145 2470 18155 2490
rect 18175 2470 18185 2490
rect 15665 2455 15705 2470
rect 18145 2455 18185 2470
rect 18200 2640 18240 2655
rect 18200 2620 18210 2640
rect 18230 2620 18240 2640
rect 18200 2590 18240 2620
rect 18200 2570 18210 2590
rect 18230 2570 18240 2590
rect 18200 2540 18240 2570
rect 18200 2520 18210 2540
rect 18230 2520 18240 2540
rect 18200 2490 18240 2520
rect 18200 2470 18210 2490
rect 18230 2470 18240 2490
rect 18200 2455 18240 2470
rect 18255 2640 18295 2655
rect 18255 2620 18265 2640
rect 18285 2620 18295 2640
rect 18255 2590 18295 2620
rect 18255 2570 18265 2590
rect 18285 2570 18295 2590
rect 18255 2540 18295 2570
rect 18255 2520 18265 2540
rect 18285 2520 18295 2540
rect 18255 2490 18295 2520
rect 18255 2470 18265 2490
rect 18285 2470 18295 2490
rect 18255 2455 18295 2470
rect 18310 2640 18350 2655
rect 18310 2620 18320 2640
rect 18340 2620 18350 2640
rect 18310 2590 18350 2620
rect 18310 2570 18320 2590
rect 18340 2570 18350 2590
rect 18310 2540 18350 2570
rect 18310 2520 18320 2540
rect 18340 2520 18350 2540
rect 18310 2490 18350 2520
rect 18310 2470 18320 2490
rect 18340 2470 18350 2490
rect 18310 2455 18350 2470
rect 18365 2640 18405 2655
rect 18365 2620 18375 2640
rect 18395 2620 18405 2640
rect 18365 2590 18405 2620
rect 18365 2570 18375 2590
rect 18395 2570 18405 2590
rect 18365 2540 18405 2570
rect 18365 2520 18375 2540
rect 18395 2520 18405 2540
rect 18365 2490 18405 2520
rect 18365 2470 18375 2490
rect 18395 2470 18405 2490
rect 18365 2455 18405 2470
rect 18420 2640 18460 2655
rect 18420 2620 18430 2640
rect 18450 2620 18460 2640
rect 18420 2590 18460 2620
rect 18420 2570 18430 2590
rect 18450 2570 18460 2590
rect 18420 2540 18460 2570
rect 18420 2520 18430 2540
rect 18450 2520 18460 2540
rect 18420 2490 18460 2520
rect 18420 2470 18430 2490
rect 18450 2470 18460 2490
rect 18420 2455 18460 2470
rect 18475 2640 18515 2655
rect 18475 2620 18485 2640
rect 18505 2620 18515 2640
rect 18475 2590 18515 2620
rect 18475 2570 18485 2590
rect 18505 2570 18515 2590
rect 18475 2540 18515 2570
rect 18475 2520 18485 2540
rect 18505 2520 18515 2540
rect 18475 2490 18515 2520
rect 18475 2470 18485 2490
rect 18505 2470 18515 2490
rect 18475 2455 18515 2470
rect 18530 2640 18570 2655
rect 18530 2620 18540 2640
rect 18560 2620 18570 2640
rect 18530 2590 18570 2620
rect 18530 2570 18540 2590
rect 18560 2570 18570 2590
rect 18530 2540 18570 2570
rect 18530 2520 18540 2540
rect 18560 2520 18570 2540
rect 18530 2490 18570 2520
rect 18530 2470 18540 2490
rect 18560 2470 18570 2490
rect 18530 2455 18570 2470
rect 18585 2640 18625 2655
rect 18585 2620 18595 2640
rect 18615 2620 18625 2640
rect 18585 2590 18625 2620
rect 18585 2570 18595 2590
rect 18615 2570 18625 2590
rect 18585 2540 18625 2570
rect 18585 2520 18595 2540
rect 18615 2520 18625 2540
rect 18585 2490 18625 2520
rect 18585 2470 18595 2490
rect 18615 2470 18625 2490
rect 18585 2455 18625 2470
rect 18640 2640 18680 2655
rect 18640 2620 18650 2640
rect 18670 2620 18680 2640
rect 18640 2590 18680 2620
rect 18640 2570 18650 2590
rect 18670 2570 18680 2590
rect 18640 2540 18680 2570
rect 18640 2520 18650 2540
rect 18670 2520 18680 2540
rect 18640 2490 18680 2520
rect 18640 2470 18650 2490
rect 18670 2470 18680 2490
rect 18640 2455 18680 2470
rect 18695 2640 18735 2655
rect 18695 2620 18705 2640
rect 18725 2620 18735 2640
rect 18695 2590 18735 2620
rect 18695 2570 18705 2590
rect 18725 2570 18735 2590
rect 18695 2540 18735 2570
rect 18695 2520 18705 2540
rect 18725 2520 18735 2540
rect 18695 2490 18735 2520
rect 18695 2470 18705 2490
rect 18725 2470 18735 2490
rect 18695 2455 18735 2470
rect 18750 2640 18790 2655
rect 18750 2620 18760 2640
rect 18780 2620 18790 2640
rect 18750 2590 18790 2620
rect 18750 2570 18760 2590
rect 18780 2570 18790 2590
rect 18750 2540 18790 2570
rect 18750 2520 18760 2540
rect 18780 2520 18790 2540
rect 18750 2490 18790 2520
rect 18750 2470 18760 2490
rect 18780 2470 18790 2490
rect 18750 2455 18790 2470
rect 18805 2640 18845 2655
rect 18805 2620 18815 2640
rect 18835 2620 18845 2640
rect 25005 2640 25045 2655
rect 18805 2590 18845 2620
rect 18805 2570 18815 2590
rect 18835 2570 18845 2590
rect 18805 2540 18845 2570
rect 18805 2520 18815 2540
rect 18835 2520 18845 2540
rect 18805 2490 18845 2520
rect 18805 2470 18815 2490
rect 18835 2470 18845 2490
rect 18805 2455 18845 2470
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 4025 1985 4065 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 3945 1935 3985 1965
rect 4025 1935 4065 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 3945 1900 3985 1915
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 5225 1985 5265 2000
rect 5225 1965 5235 1985
rect 5255 1965 5265 1985
rect 5225 1935 5265 1965
rect 25005 2620 25015 2640
rect 25035 2620 25045 2640
rect 25005 2590 25045 2620
rect 25005 2570 25015 2590
rect 25035 2570 25045 2590
rect 25005 2540 25045 2570
rect 25005 2520 25015 2540
rect 25035 2520 25045 2540
rect 25005 2490 25045 2520
rect 25005 2470 25015 2490
rect 25035 2470 25045 2490
rect 25005 2455 25045 2470
rect 25060 2640 25100 2655
rect 25060 2620 25070 2640
rect 25090 2620 25100 2640
rect 25060 2590 25100 2620
rect 25060 2570 25070 2590
rect 25090 2570 25100 2590
rect 25060 2540 25100 2570
rect 25060 2520 25070 2540
rect 25090 2520 25100 2540
rect 25060 2490 25100 2520
rect 25060 2470 25070 2490
rect 25090 2470 25100 2490
rect 25060 2455 25100 2470
rect 25115 2640 25155 2655
rect 25115 2620 25125 2640
rect 25145 2620 25155 2640
rect 25115 2590 25155 2620
rect 25115 2570 25125 2590
rect 25145 2570 25155 2590
rect 25115 2540 25155 2570
rect 25115 2520 25125 2540
rect 25145 2520 25155 2540
rect 25115 2490 25155 2520
rect 25115 2470 25125 2490
rect 25145 2470 25155 2490
rect 25115 2455 25155 2470
rect 25170 2640 25210 2655
rect 25170 2620 25180 2640
rect 25200 2620 25210 2640
rect 25170 2590 25210 2620
rect 25170 2570 25180 2590
rect 25200 2570 25210 2590
rect 25170 2540 25210 2570
rect 25170 2520 25180 2540
rect 25200 2520 25210 2540
rect 25170 2490 25210 2520
rect 25170 2470 25180 2490
rect 25200 2470 25210 2490
rect 25170 2455 25210 2470
rect 25225 2640 25265 2655
rect 25225 2620 25235 2640
rect 25255 2620 25265 2640
rect 25225 2590 25265 2620
rect 25225 2570 25235 2590
rect 25255 2570 25265 2590
rect 25225 2540 25265 2570
rect 25225 2520 25235 2540
rect 25255 2520 25265 2540
rect 25225 2490 25265 2520
rect 25225 2470 25235 2490
rect 25255 2470 25265 2490
rect 25225 2455 25265 2470
rect 25280 2640 25320 2655
rect 25280 2620 25290 2640
rect 25310 2620 25320 2640
rect 25280 2590 25320 2620
rect 25280 2570 25290 2590
rect 25310 2570 25320 2590
rect 25280 2540 25320 2570
rect 25280 2520 25290 2540
rect 25310 2520 25320 2540
rect 25280 2490 25320 2520
rect 25280 2470 25290 2490
rect 25310 2470 25320 2490
rect 25280 2455 25320 2470
rect 25335 2640 25375 2655
rect 25335 2620 25345 2640
rect 25365 2620 25375 2640
rect 25335 2590 25375 2620
rect 25335 2570 25345 2590
rect 25365 2570 25375 2590
rect 25335 2540 25375 2570
rect 25335 2520 25345 2540
rect 25365 2520 25375 2540
rect 25335 2490 25375 2520
rect 25335 2470 25345 2490
rect 25365 2470 25375 2490
rect 25335 2455 25375 2470
rect 25390 2640 25430 2655
rect 25390 2620 25400 2640
rect 25420 2620 25430 2640
rect 25390 2590 25430 2620
rect 25390 2570 25400 2590
rect 25420 2570 25430 2590
rect 25390 2540 25430 2570
rect 25390 2520 25400 2540
rect 25420 2520 25430 2540
rect 25390 2490 25430 2520
rect 25390 2470 25400 2490
rect 25420 2470 25430 2490
rect 25390 2455 25430 2470
rect 25445 2640 25485 2655
rect 25445 2620 25455 2640
rect 25475 2620 25485 2640
rect 25445 2590 25485 2620
rect 25445 2570 25455 2590
rect 25475 2570 25485 2590
rect 25445 2540 25485 2570
rect 25445 2520 25455 2540
rect 25475 2520 25485 2540
rect 25445 2490 25485 2520
rect 25445 2470 25455 2490
rect 25475 2470 25485 2490
rect 25445 2455 25485 2470
rect 25500 2640 25540 2655
rect 25500 2620 25510 2640
rect 25530 2620 25540 2640
rect 25500 2590 25540 2620
rect 25500 2570 25510 2590
rect 25530 2570 25540 2590
rect 25500 2540 25540 2570
rect 25500 2520 25510 2540
rect 25530 2520 25540 2540
rect 25500 2490 25540 2520
rect 25500 2470 25510 2490
rect 25530 2470 25540 2490
rect 25500 2455 25540 2470
rect 25555 2640 25595 2655
rect 25555 2620 25565 2640
rect 25585 2620 25595 2640
rect 25555 2590 25595 2620
rect 25555 2570 25565 2590
rect 25585 2570 25595 2590
rect 25555 2540 25595 2570
rect 25555 2520 25565 2540
rect 25585 2520 25595 2540
rect 25555 2490 25595 2520
rect 25555 2470 25565 2490
rect 25585 2470 25595 2490
rect 25555 2455 25595 2470
rect 25610 2640 25650 2655
rect 25610 2620 25620 2640
rect 25640 2620 25650 2640
rect 25610 2590 25650 2620
rect 25610 2570 25620 2590
rect 25640 2570 25650 2590
rect 25610 2540 25650 2570
rect 25610 2520 25620 2540
rect 25640 2520 25650 2540
rect 25610 2490 25650 2520
rect 25610 2470 25620 2490
rect 25640 2470 25650 2490
rect 25610 2455 25650 2470
rect 25665 2640 25705 2655
rect 25665 2620 25675 2640
rect 25695 2620 25705 2640
rect 25665 2590 25705 2620
rect 25665 2570 25675 2590
rect 25695 2570 25705 2590
rect 25665 2540 25705 2570
rect 25665 2520 25675 2540
rect 25695 2520 25705 2540
rect 25665 2490 25705 2520
rect 26015 2630 26055 2660
rect 26015 2610 26025 2630
rect 26045 2610 26055 2630
rect 26015 2580 26055 2610
rect 26015 2560 26025 2580
rect 26045 2560 26055 2580
rect 26015 2530 26055 2560
rect 26015 2510 26025 2530
rect 26045 2510 26055 2530
rect 26015 2495 26055 2510
rect 26075 2830 26115 2845
rect 26075 2810 26085 2830
rect 26105 2810 26115 2830
rect 26075 2780 26115 2810
rect 26075 2760 26085 2780
rect 26105 2760 26115 2780
rect 26075 2730 26115 2760
rect 26075 2710 26085 2730
rect 26105 2710 26115 2730
rect 26075 2680 26115 2710
rect 26075 2660 26085 2680
rect 26105 2660 26115 2680
rect 26075 2630 26115 2660
rect 26075 2610 26085 2630
rect 26105 2610 26115 2630
rect 26075 2580 26115 2610
rect 26075 2560 26085 2580
rect 26105 2560 26115 2580
rect 26075 2530 26115 2560
rect 26075 2510 26085 2530
rect 26105 2510 26115 2530
rect 26075 2495 26115 2510
rect 26135 2830 26175 2845
rect 26135 2810 26145 2830
rect 26165 2810 26175 2830
rect 26135 2780 26175 2810
rect 26135 2760 26145 2780
rect 26165 2760 26175 2780
rect 26135 2730 26175 2760
rect 26135 2710 26145 2730
rect 26165 2710 26175 2730
rect 26135 2680 26175 2710
rect 26135 2660 26145 2680
rect 26165 2660 26175 2680
rect 26135 2630 26175 2660
rect 26135 2610 26145 2630
rect 26165 2610 26175 2630
rect 26135 2580 26175 2610
rect 26135 2560 26145 2580
rect 26165 2560 26175 2580
rect 26135 2530 26175 2560
rect 26135 2510 26145 2530
rect 26165 2510 26175 2530
rect 26135 2495 26175 2510
rect 26195 2830 26235 2845
rect 26195 2810 26205 2830
rect 26225 2810 26235 2830
rect 26195 2780 26235 2810
rect 26195 2760 26205 2780
rect 26225 2760 26235 2780
rect 26195 2730 26235 2760
rect 26195 2710 26205 2730
rect 26225 2710 26235 2730
rect 26195 2680 26235 2710
rect 26195 2660 26205 2680
rect 26225 2660 26235 2680
rect 26195 2630 26235 2660
rect 26195 2610 26205 2630
rect 26225 2610 26235 2630
rect 26195 2580 26235 2610
rect 26195 2560 26205 2580
rect 26225 2560 26235 2580
rect 26195 2530 26235 2560
rect 26195 2510 26205 2530
rect 26225 2510 26235 2530
rect 26195 2495 26235 2510
rect 26255 2830 26295 2845
rect 26255 2810 26265 2830
rect 26285 2810 26295 2830
rect 26255 2780 26295 2810
rect 26255 2760 26265 2780
rect 26285 2760 26295 2780
rect 26255 2730 26295 2760
rect 26255 2710 26265 2730
rect 26285 2710 26295 2730
rect 26255 2680 26295 2710
rect 26255 2660 26265 2680
rect 26285 2660 26295 2680
rect 26255 2630 26295 2660
rect 26255 2610 26265 2630
rect 26285 2610 26295 2630
rect 26255 2580 26295 2610
rect 26255 2560 26265 2580
rect 26285 2560 26295 2580
rect 26255 2530 26295 2560
rect 26255 2510 26265 2530
rect 26285 2510 26295 2530
rect 26255 2495 26295 2510
rect 26315 2830 26355 2845
rect 26315 2810 26325 2830
rect 26345 2810 26355 2830
rect 26315 2780 26355 2810
rect 26315 2760 26325 2780
rect 26345 2760 26355 2780
rect 26315 2730 26355 2760
rect 26315 2710 26325 2730
rect 26345 2710 26355 2730
rect 26315 2680 26355 2710
rect 26315 2660 26325 2680
rect 26345 2660 26355 2680
rect 26315 2630 26355 2660
rect 26315 2610 26325 2630
rect 26345 2610 26355 2630
rect 26315 2580 26355 2610
rect 26315 2560 26325 2580
rect 26345 2560 26355 2580
rect 26315 2530 26355 2560
rect 26315 2510 26325 2530
rect 26345 2510 26355 2530
rect 26315 2495 26355 2510
rect 26375 2830 26415 2845
rect 26375 2810 26385 2830
rect 26405 2810 26415 2830
rect 26375 2780 26415 2810
rect 26375 2760 26385 2780
rect 26405 2760 26415 2780
rect 26375 2730 26415 2760
rect 26375 2710 26385 2730
rect 26405 2710 26415 2730
rect 26375 2680 26415 2710
rect 26375 2660 26385 2680
rect 26405 2660 26415 2680
rect 26375 2630 26415 2660
rect 26375 2610 26385 2630
rect 26405 2610 26415 2630
rect 26375 2580 26415 2610
rect 26375 2560 26385 2580
rect 26405 2560 26415 2580
rect 26375 2530 26415 2560
rect 26375 2510 26385 2530
rect 26405 2510 26415 2530
rect 26375 2495 26415 2510
rect 26435 2830 26475 2845
rect 26435 2810 26445 2830
rect 26465 2810 26475 2830
rect 26435 2780 26475 2810
rect 26435 2760 26445 2780
rect 26465 2760 26475 2780
rect 26435 2730 26475 2760
rect 26435 2710 26445 2730
rect 26465 2710 26475 2730
rect 26435 2680 26475 2710
rect 26435 2660 26445 2680
rect 26465 2660 26475 2680
rect 26435 2630 26475 2660
rect 26435 2610 26445 2630
rect 26465 2610 26475 2630
rect 26435 2580 26475 2610
rect 26435 2560 26445 2580
rect 26465 2560 26475 2580
rect 26435 2530 26475 2560
rect 26435 2510 26445 2530
rect 26465 2510 26475 2530
rect 26435 2495 26475 2510
rect 26495 2830 26535 2845
rect 26495 2810 26505 2830
rect 26525 2810 26535 2830
rect 26495 2780 26535 2810
rect 26495 2760 26505 2780
rect 26525 2760 26535 2780
rect 26495 2730 26535 2760
rect 26495 2710 26505 2730
rect 26525 2710 26535 2730
rect 26495 2680 26535 2710
rect 26495 2660 26505 2680
rect 26525 2660 26535 2680
rect 26495 2630 26535 2660
rect 26495 2610 26505 2630
rect 26525 2610 26535 2630
rect 26495 2580 26535 2610
rect 26495 2560 26505 2580
rect 26525 2560 26535 2580
rect 26495 2530 26535 2560
rect 26495 2510 26505 2530
rect 26525 2510 26535 2530
rect 26495 2495 26535 2510
rect 26555 2830 26595 2845
rect 26555 2810 26565 2830
rect 26585 2810 26595 2830
rect 26555 2780 26595 2810
rect 26555 2760 26565 2780
rect 26585 2760 26595 2780
rect 26555 2730 26595 2760
rect 26555 2710 26565 2730
rect 26585 2710 26595 2730
rect 26555 2680 26595 2710
rect 26555 2660 26565 2680
rect 26585 2660 26595 2680
rect 26555 2630 26595 2660
rect 26555 2610 26565 2630
rect 26585 2610 26595 2630
rect 26555 2580 26595 2610
rect 26555 2560 26565 2580
rect 26585 2560 26595 2580
rect 26555 2530 26595 2560
rect 26555 2510 26565 2530
rect 26585 2510 26595 2530
rect 26555 2495 26595 2510
rect 26615 2830 26655 2845
rect 26615 2810 26625 2830
rect 26645 2810 26655 2830
rect 26615 2780 26655 2810
rect 26615 2760 26625 2780
rect 26645 2760 26655 2780
rect 26615 2730 26655 2760
rect 26615 2710 26625 2730
rect 26645 2710 26655 2730
rect 26615 2680 26655 2710
rect 26615 2660 26625 2680
rect 26645 2660 26655 2680
rect 26615 2630 26655 2660
rect 26615 2610 26625 2630
rect 26645 2610 26655 2630
rect 26615 2580 26655 2610
rect 26615 2560 26625 2580
rect 26645 2560 26655 2580
rect 26615 2530 26655 2560
rect 26615 2510 26625 2530
rect 26645 2510 26655 2530
rect 26615 2495 26655 2510
rect 26675 2830 26715 2845
rect 26675 2810 26685 2830
rect 26705 2810 26715 2830
rect 26675 2780 26715 2810
rect 26675 2760 26685 2780
rect 26705 2760 26715 2780
rect 26675 2730 26715 2760
rect 26675 2710 26685 2730
rect 26705 2710 26715 2730
rect 26675 2680 26715 2710
rect 26675 2660 26685 2680
rect 26705 2660 26715 2680
rect 26675 2630 26715 2660
rect 26675 2610 26685 2630
rect 26705 2610 26715 2630
rect 26675 2580 26715 2610
rect 26675 2560 26685 2580
rect 26705 2560 26715 2580
rect 26675 2530 26715 2560
rect 26675 2510 26685 2530
rect 26705 2510 26715 2530
rect 26675 2495 26715 2510
rect 26735 2830 26775 2845
rect 26735 2810 26745 2830
rect 26765 2810 26775 2830
rect 26735 2780 26775 2810
rect 26735 2760 26745 2780
rect 26765 2760 26775 2780
rect 26735 2730 26775 2760
rect 26735 2710 26745 2730
rect 26765 2710 26775 2730
rect 26735 2680 26775 2710
rect 26735 2660 26745 2680
rect 26765 2660 26775 2680
rect 26735 2630 26775 2660
rect 26735 2610 26745 2630
rect 26765 2610 26775 2630
rect 26735 2580 26775 2610
rect 26735 2560 26745 2580
rect 26765 2560 26775 2580
rect 26735 2530 26775 2560
rect 26735 2510 26745 2530
rect 26765 2510 26775 2530
rect 26735 2495 26775 2510
rect 25665 2470 25675 2490
rect 25695 2470 25705 2490
rect 25665 2455 25705 2470
rect 27035 2830 27075 2845
rect 27035 2810 27045 2830
rect 27065 2810 27075 2830
rect 27035 2780 27075 2810
rect 27035 2760 27045 2780
rect 27065 2760 27075 2780
rect 27035 2730 27075 2760
rect 27035 2710 27045 2730
rect 27065 2710 27075 2730
rect 27035 2680 27075 2710
rect 27035 2660 27045 2680
rect 27065 2660 27075 2680
rect 27035 2630 27075 2660
rect 27035 2610 27045 2630
rect 27065 2610 27075 2630
rect 27035 2580 27075 2610
rect 27035 2560 27045 2580
rect 27065 2560 27075 2580
rect 27035 2530 27075 2560
rect 27035 2510 27045 2530
rect 27065 2510 27075 2530
rect 27035 2495 27075 2510
rect 27095 2830 27135 2845
rect 27095 2810 27105 2830
rect 27125 2810 27135 2830
rect 27095 2780 27135 2810
rect 27095 2760 27105 2780
rect 27125 2760 27135 2780
rect 27095 2730 27135 2760
rect 27095 2710 27105 2730
rect 27125 2710 27135 2730
rect 27095 2680 27135 2710
rect 27095 2660 27105 2680
rect 27125 2660 27135 2680
rect 27095 2630 27135 2660
rect 27095 2610 27105 2630
rect 27125 2610 27135 2630
rect 27095 2580 27135 2610
rect 27095 2560 27105 2580
rect 27125 2560 27135 2580
rect 27095 2530 27135 2560
rect 27095 2510 27105 2530
rect 27125 2510 27135 2530
rect 27095 2495 27135 2510
rect 27155 2830 27195 2845
rect 27155 2810 27165 2830
rect 27185 2810 27195 2830
rect 27155 2780 27195 2810
rect 27155 2760 27165 2780
rect 27185 2760 27195 2780
rect 27155 2730 27195 2760
rect 27155 2710 27165 2730
rect 27185 2710 27195 2730
rect 27155 2680 27195 2710
rect 27155 2660 27165 2680
rect 27185 2660 27195 2680
rect 27155 2630 27195 2660
rect 27155 2610 27165 2630
rect 27185 2610 27195 2630
rect 27155 2580 27195 2610
rect 27155 2560 27165 2580
rect 27185 2560 27195 2580
rect 27155 2530 27195 2560
rect 27155 2510 27165 2530
rect 27185 2510 27195 2530
rect 27155 2495 27195 2510
rect 27215 2830 27255 2845
rect 27215 2810 27225 2830
rect 27245 2810 27255 2830
rect 27215 2780 27255 2810
rect 27215 2760 27225 2780
rect 27245 2760 27255 2780
rect 27215 2730 27255 2760
rect 27215 2710 27225 2730
rect 27245 2710 27255 2730
rect 27215 2680 27255 2710
rect 27215 2660 27225 2680
rect 27245 2660 27255 2680
rect 27215 2630 27255 2660
rect 27215 2610 27225 2630
rect 27245 2610 27255 2630
rect 27215 2580 27255 2610
rect 27215 2560 27225 2580
rect 27245 2560 27255 2580
rect 27215 2530 27255 2560
rect 27215 2510 27225 2530
rect 27245 2510 27255 2530
rect 27215 2495 27255 2510
rect 27275 2830 27315 2845
rect 27275 2810 27285 2830
rect 27305 2810 27315 2830
rect 27275 2780 27315 2810
rect 27275 2760 27285 2780
rect 27305 2760 27315 2780
rect 27275 2730 27315 2760
rect 27275 2710 27285 2730
rect 27305 2710 27315 2730
rect 27275 2680 27315 2710
rect 27275 2660 27285 2680
rect 27305 2660 27315 2680
rect 27275 2630 27315 2660
rect 27275 2610 27285 2630
rect 27305 2610 27315 2630
rect 27275 2580 27315 2610
rect 27275 2560 27285 2580
rect 27305 2560 27315 2580
rect 27275 2530 27315 2560
rect 27275 2510 27285 2530
rect 27305 2510 27315 2530
rect 27275 2495 27315 2510
rect 27335 2830 27375 2845
rect 27335 2810 27345 2830
rect 27365 2810 27375 2830
rect 27335 2780 27375 2810
rect 27335 2760 27345 2780
rect 27365 2760 27375 2780
rect 27335 2730 27375 2760
rect 27335 2710 27345 2730
rect 27365 2710 27375 2730
rect 27335 2680 27375 2710
rect 27335 2660 27345 2680
rect 27365 2660 27375 2680
rect 27335 2630 27375 2660
rect 27335 2610 27345 2630
rect 27365 2610 27375 2630
rect 27335 2580 27375 2610
rect 27335 2560 27345 2580
rect 27365 2560 27375 2580
rect 27335 2530 27375 2560
rect 27335 2510 27345 2530
rect 27365 2510 27375 2530
rect 27335 2495 27375 2510
rect 27395 2830 27435 2845
rect 27395 2810 27405 2830
rect 27425 2810 27435 2830
rect 27395 2780 27435 2810
rect 27395 2760 27405 2780
rect 27425 2760 27435 2780
rect 27395 2730 27435 2760
rect 27395 2710 27405 2730
rect 27425 2710 27435 2730
rect 27395 2680 27435 2710
rect 27395 2660 27405 2680
rect 27425 2660 27435 2680
rect 27395 2630 27435 2660
rect 27395 2610 27405 2630
rect 27425 2610 27435 2630
rect 27395 2580 27435 2610
rect 27395 2560 27405 2580
rect 27425 2560 27435 2580
rect 27395 2530 27435 2560
rect 27395 2510 27405 2530
rect 27425 2510 27435 2530
rect 27395 2495 27435 2510
rect 27455 2830 27495 2845
rect 27455 2810 27465 2830
rect 27485 2810 27495 2830
rect 27455 2780 27495 2810
rect 27455 2760 27465 2780
rect 27485 2760 27495 2780
rect 27455 2730 27495 2760
rect 27455 2710 27465 2730
rect 27485 2710 27495 2730
rect 27455 2680 27495 2710
rect 27455 2660 27465 2680
rect 27485 2660 27495 2680
rect 27455 2630 27495 2660
rect 27455 2610 27465 2630
rect 27485 2610 27495 2630
rect 27455 2580 27495 2610
rect 27455 2560 27465 2580
rect 27485 2560 27495 2580
rect 27455 2530 27495 2560
rect 27455 2510 27465 2530
rect 27485 2510 27495 2530
rect 27455 2495 27495 2510
rect 27515 2830 27555 2845
rect 27515 2810 27525 2830
rect 27545 2810 27555 2830
rect 27515 2780 27555 2810
rect 27515 2760 27525 2780
rect 27545 2760 27555 2780
rect 27515 2730 27555 2760
rect 27515 2710 27525 2730
rect 27545 2710 27555 2730
rect 27515 2680 27555 2710
rect 27515 2660 27525 2680
rect 27545 2660 27555 2680
rect 27515 2630 27555 2660
rect 27515 2610 27525 2630
rect 27545 2610 27555 2630
rect 27515 2580 27555 2610
rect 27515 2560 27525 2580
rect 27545 2560 27555 2580
rect 27515 2530 27555 2560
rect 27515 2510 27525 2530
rect 27545 2510 27555 2530
rect 27515 2495 27555 2510
rect 27575 2830 27615 2845
rect 27575 2810 27585 2830
rect 27605 2810 27615 2830
rect 27575 2780 27615 2810
rect 27575 2760 27585 2780
rect 27605 2760 27615 2780
rect 27575 2730 27615 2760
rect 27575 2710 27585 2730
rect 27605 2710 27615 2730
rect 27575 2680 27615 2710
rect 27575 2660 27585 2680
rect 27605 2660 27615 2680
rect 27575 2630 27615 2660
rect 27575 2610 27585 2630
rect 27605 2610 27615 2630
rect 27575 2580 27615 2610
rect 27575 2560 27585 2580
rect 27605 2560 27615 2580
rect 27575 2530 27615 2560
rect 27575 2510 27585 2530
rect 27605 2510 27615 2530
rect 27575 2495 27615 2510
rect 27635 2830 27675 2845
rect 27635 2810 27645 2830
rect 27665 2810 27675 2830
rect 27635 2780 27675 2810
rect 27635 2760 27645 2780
rect 27665 2760 27675 2780
rect 27635 2730 27675 2760
rect 27635 2710 27645 2730
rect 27665 2710 27675 2730
rect 27635 2680 27675 2710
rect 27635 2660 27645 2680
rect 27665 2660 27675 2680
rect 27635 2630 27675 2660
rect 27635 2610 27645 2630
rect 27665 2610 27675 2630
rect 27635 2580 27675 2610
rect 27635 2560 27645 2580
rect 27665 2560 27675 2580
rect 27635 2530 27675 2560
rect 27635 2510 27645 2530
rect 27665 2510 27675 2530
rect 27635 2495 27675 2510
rect 27695 2830 27735 2845
rect 27695 2810 27705 2830
rect 27725 2810 27735 2830
rect 27695 2780 27735 2810
rect 27695 2760 27705 2780
rect 27725 2760 27735 2780
rect 27695 2730 27735 2760
rect 27695 2710 27705 2730
rect 27725 2710 27735 2730
rect 27695 2680 27735 2710
rect 27695 2660 27705 2680
rect 27725 2660 27735 2680
rect 27695 2630 27735 2660
rect 27695 2610 27705 2630
rect 27725 2610 27735 2630
rect 27695 2580 27735 2610
rect 27695 2560 27705 2580
rect 27725 2560 27735 2580
rect 27695 2530 27735 2560
rect 27695 2510 27705 2530
rect 27725 2510 27735 2530
rect 27695 2495 27735 2510
rect 27755 2830 27795 2845
rect 27755 2810 27765 2830
rect 27785 2810 27795 2830
rect 27755 2780 27795 2810
rect 27755 2760 27765 2780
rect 27785 2760 27795 2780
rect 27755 2730 27795 2760
rect 27755 2710 27765 2730
rect 27785 2710 27795 2730
rect 27755 2680 27795 2710
rect 27755 2660 27765 2680
rect 27785 2660 27795 2680
rect 27755 2630 27795 2660
rect 27755 2610 27765 2630
rect 27785 2610 27795 2630
rect 27755 2580 27795 2610
rect 27755 2560 27765 2580
rect 27785 2560 27795 2580
rect 27755 2530 27795 2560
rect 27755 2510 27765 2530
rect 27785 2510 27795 2530
rect 27755 2495 27795 2510
rect 28145 2690 28185 2705
rect 28145 2670 28155 2690
rect 28175 2670 28185 2690
rect 28145 2640 28185 2670
rect 28145 2620 28155 2640
rect 28175 2620 28185 2640
rect 28145 2590 28185 2620
rect 28145 2570 28155 2590
rect 28175 2570 28185 2590
rect 28145 2540 28185 2570
rect 28145 2520 28155 2540
rect 28175 2520 28185 2540
rect 28145 2505 28185 2520
rect 28200 2690 28240 2705
rect 28200 2670 28210 2690
rect 28230 2670 28240 2690
rect 28200 2640 28240 2670
rect 28200 2620 28210 2640
rect 28230 2620 28240 2640
rect 28200 2590 28240 2620
rect 28200 2570 28210 2590
rect 28230 2570 28240 2590
rect 28200 2540 28240 2570
rect 28200 2520 28210 2540
rect 28230 2520 28240 2540
rect 28200 2505 28240 2520
rect 28255 2690 28295 2705
rect 28255 2670 28265 2690
rect 28285 2670 28295 2690
rect 28255 2640 28295 2670
rect 28255 2620 28265 2640
rect 28285 2620 28295 2640
rect 28255 2590 28295 2620
rect 28255 2570 28265 2590
rect 28285 2570 28295 2590
rect 28255 2540 28295 2570
rect 28255 2520 28265 2540
rect 28285 2520 28295 2540
rect 28255 2505 28295 2520
rect 28310 2690 28350 2705
rect 28310 2670 28320 2690
rect 28340 2670 28350 2690
rect 28310 2640 28350 2670
rect 28310 2620 28320 2640
rect 28340 2620 28350 2640
rect 28310 2590 28350 2620
rect 28310 2570 28320 2590
rect 28340 2570 28350 2590
rect 28310 2540 28350 2570
rect 28310 2520 28320 2540
rect 28340 2520 28350 2540
rect 28310 2505 28350 2520
rect 28365 2690 28405 2705
rect 28365 2670 28375 2690
rect 28395 2670 28405 2690
rect 28365 2640 28405 2670
rect 28365 2620 28375 2640
rect 28395 2620 28405 2640
rect 28365 2590 28405 2620
rect 28365 2570 28375 2590
rect 28395 2570 28405 2590
rect 28365 2540 28405 2570
rect 28365 2520 28375 2540
rect 28395 2520 28405 2540
rect 28365 2505 28405 2520
rect 28420 2690 28460 2705
rect 28420 2670 28430 2690
rect 28450 2670 28460 2690
rect 28420 2640 28460 2670
rect 28420 2620 28430 2640
rect 28450 2620 28460 2640
rect 28420 2590 28460 2620
rect 28420 2570 28430 2590
rect 28450 2570 28460 2590
rect 28420 2540 28460 2570
rect 28420 2520 28430 2540
rect 28450 2520 28460 2540
rect 28420 2505 28460 2520
rect 28475 2690 28515 2705
rect 28475 2670 28485 2690
rect 28505 2670 28515 2690
rect 28475 2640 28515 2670
rect 28475 2620 28485 2640
rect 28505 2620 28515 2640
rect 28475 2590 28515 2620
rect 28475 2570 28485 2590
rect 28505 2570 28515 2590
rect 28475 2540 28515 2570
rect 28475 2520 28485 2540
rect 28505 2520 28515 2540
rect 28475 2505 28515 2520
rect 28530 2690 28570 2705
rect 28530 2670 28540 2690
rect 28560 2670 28570 2690
rect 28530 2640 28570 2670
rect 28530 2620 28540 2640
rect 28560 2620 28570 2640
rect 28530 2590 28570 2620
rect 28530 2570 28540 2590
rect 28560 2570 28570 2590
rect 28530 2540 28570 2570
rect 28530 2520 28540 2540
rect 28560 2520 28570 2540
rect 28530 2505 28570 2520
rect 28585 2690 28625 2705
rect 28585 2670 28595 2690
rect 28615 2670 28625 2690
rect 28585 2640 28625 2670
rect 28585 2620 28595 2640
rect 28615 2620 28625 2640
rect 28585 2590 28625 2620
rect 28585 2570 28595 2590
rect 28615 2570 28625 2590
rect 28585 2540 28625 2570
rect 28585 2520 28595 2540
rect 28615 2520 28625 2540
rect 28585 2505 28625 2520
rect 28640 2690 28680 2705
rect 28640 2670 28650 2690
rect 28670 2670 28680 2690
rect 28640 2640 28680 2670
rect 28640 2620 28650 2640
rect 28670 2620 28680 2640
rect 28640 2590 28680 2620
rect 28640 2570 28650 2590
rect 28670 2570 28680 2590
rect 28640 2540 28680 2570
rect 28640 2520 28650 2540
rect 28670 2520 28680 2540
rect 28640 2505 28680 2520
rect 28695 2690 28735 2705
rect 28695 2670 28705 2690
rect 28725 2670 28735 2690
rect 28695 2640 28735 2670
rect 28695 2620 28705 2640
rect 28725 2620 28735 2640
rect 28695 2590 28735 2620
rect 28695 2570 28705 2590
rect 28725 2570 28735 2590
rect 28695 2540 28735 2570
rect 28695 2520 28705 2540
rect 28725 2520 28735 2540
rect 28695 2505 28735 2520
rect 28750 2690 28790 2705
rect 28750 2670 28760 2690
rect 28780 2670 28790 2690
rect 28750 2640 28790 2670
rect 28750 2620 28760 2640
rect 28780 2620 28790 2640
rect 28750 2590 28790 2620
rect 28750 2570 28760 2590
rect 28780 2570 28790 2590
rect 28750 2540 28790 2570
rect 28750 2520 28760 2540
rect 28780 2520 28790 2540
rect 28750 2505 28790 2520
rect 28805 2690 28845 2705
rect 28805 2670 28815 2690
rect 28835 2670 28845 2690
rect 28805 2640 28845 2670
rect 28805 2620 28815 2640
rect 28835 2620 28845 2640
rect 28805 2590 28845 2620
rect 28805 2570 28815 2590
rect 28835 2570 28845 2590
rect 28805 2540 28845 2570
rect 28805 2520 28815 2540
rect 28835 2520 28845 2540
rect 28805 2505 28845 2520
rect 5225 1915 5235 1935
rect 5255 1915 5265 1935
rect 5225 1900 5265 1915
<< ndiffc >>
rect 15015 2230 15035 2250
rect 15015 2180 15035 2200
rect 15015 2130 15035 2150
rect 15015 2080 15035 2100
rect 15015 2030 15035 2050
rect 15015 1980 15035 2000
rect 15070 2230 15090 2250
rect 15070 2180 15090 2200
rect 15070 2130 15090 2150
rect 15070 2080 15090 2100
rect 15070 2030 15090 2050
rect 15070 1980 15090 2000
rect 15125 2230 15145 2250
rect 15125 2180 15145 2200
rect 15125 2130 15145 2150
rect 15125 2080 15145 2100
rect 15125 2030 15145 2050
rect 15125 1980 15145 2000
rect 15180 2230 15200 2250
rect 15180 2180 15200 2200
rect 15180 2130 15200 2150
rect 15180 2080 15200 2100
rect 15180 2030 15200 2050
rect 15180 1980 15200 2000
rect 15235 2230 15255 2250
rect 15235 2180 15255 2200
rect 15235 2130 15255 2150
rect 15235 2080 15255 2100
rect 15235 2030 15255 2050
rect 15235 1980 15255 2000
rect 15290 2230 15310 2250
rect 15290 2180 15310 2200
rect 15290 2130 15310 2150
rect 15290 2080 15310 2100
rect 15290 2030 15310 2050
rect 15290 1980 15310 2000
rect 15345 2230 15365 2250
rect 15345 2180 15365 2200
rect 15345 2130 15365 2150
rect 15345 2080 15365 2100
rect 15345 2030 15365 2050
rect 15345 1980 15365 2000
rect 15400 2230 15420 2250
rect 15400 2180 15420 2200
rect 15400 2130 15420 2150
rect 15400 2080 15420 2100
rect 15400 2030 15420 2050
rect 15400 1980 15420 2000
rect 15455 2230 15475 2250
rect 15455 2180 15475 2200
rect 15455 2130 15475 2150
rect 15455 2080 15475 2100
rect 15455 2030 15475 2050
rect 15455 1980 15475 2000
rect 15510 2230 15530 2250
rect 15510 2180 15530 2200
rect 15510 2130 15530 2150
rect 15510 2080 15530 2100
rect 15510 2030 15530 2050
rect 15510 1980 15530 2000
rect 15565 2230 15585 2250
rect 15565 2180 15585 2200
rect 15565 2130 15585 2150
rect 15565 2080 15585 2100
rect 15565 2030 15585 2050
rect 15565 1980 15585 2000
rect 15620 2230 15640 2250
rect 15620 2180 15640 2200
rect 15620 2130 15640 2150
rect 15620 2080 15640 2100
rect 15620 2030 15640 2050
rect 15620 1980 15640 2000
rect 15675 2230 15695 2250
rect 15675 2180 15695 2200
rect 18155 2230 18175 2250
rect 18155 2180 18175 2200
rect 15675 2130 15695 2150
rect 18155 2130 18175 2150
rect 15675 2080 15695 2100
rect 15675 2030 15695 2050
rect 15675 1980 15695 2000
rect 16285 2095 16305 2115
rect 16285 2045 16305 2065
rect 16285 1995 16305 2015
rect 16340 2095 16360 2115
rect 16340 2045 16360 2065
rect 16340 1995 16360 2015
rect 16395 2095 16415 2115
rect 16395 2045 16415 2065
rect 16395 1995 16415 2015
rect 16450 2095 16470 2115
rect 16450 2045 16470 2065
rect 16450 1995 16470 2015
rect 16505 2095 16525 2115
rect 16505 2045 16525 2065
rect 16505 1995 16525 2015
rect 16560 2095 16580 2115
rect 16560 2045 16580 2065
rect 16560 1995 16580 2015
rect 16615 2095 16635 2115
rect 16615 2045 16635 2065
rect 16615 1995 16635 2015
rect 16670 2095 16690 2115
rect 16670 2045 16690 2065
rect 16670 1995 16690 2015
rect 16725 2095 16745 2115
rect 16725 2045 16745 2065
rect 16725 1995 16745 2015
rect 16780 2095 16800 2115
rect 16780 2045 16800 2065
rect 16780 1995 16800 2015
rect 16835 2095 16855 2115
rect 16835 2045 16855 2065
rect 16835 1995 16855 2015
rect 16890 2095 16910 2115
rect 16890 2045 16910 2065
rect 16890 1995 16910 2015
rect 16945 2095 16965 2115
rect 16945 2045 16965 2065
rect 16945 1995 16965 2015
rect 17000 2095 17020 2115
rect 17000 2045 17020 2065
rect 17000 1995 17020 2015
rect 17055 2095 17075 2115
rect 17055 2045 17075 2065
rect 17055 1995 17075 2015
rect 17110 2095 17130 2115
rect 17110 2045 17130 2065
rect 17110 1995 17130 2015
rect 17165 2095 17185 2115
rect 17165 2045 17185 2065
rect 17165 1995 17185 2015
rect 17220 2095 17240 2115
rect 17220 2045 17240 2065
rect 17220 1995 17240 2015
rect 17275 2095 17295 2115
rect 17275 2045 17295 2065
rect 17275 1995 17295 2015
rect 17330 2095 17350 2115
rect 17330 2045 17350 2065
rect 17330 1995 17350 2015
rect 17385 2095 17405 2115
rect 17385 2045 17405 2065
rect 17385 1995 17405 2015
rect 17440 2095 17460 2115
rect 17440 2045 17460 2065
rect 17440 1995 17460 2015
rect 17495 2095 17515 2115
rect 17495 2045 17515 2065
rect 17495 1995 17515 2015
rect 18155 2080 18175 2100
rect 18155 2030 18175 2050
rect 18155 1980 18175 2000
rect 18210 2230 18230 2250
rect 18210 2180 18230 2200
rect 18210 2130 18230 2150
rect 18210 2080 18230 2100
rect 18210 2030 18230 2050
rect 18210 1980 18230 2000
rect 18265 2230 18285 2250
rect 18265 2180 18285 2200
rect 18265 2130 18285 2150
rect 18265 2080 18285 2100
rect 18265 2030 18285 2050
rect 18265 1980 18285 2000
rect 18320 2230 18340 2250
rect 18320 2180 18340 2200
rect 18320 2130 18340 2150
rect 18320 2080 18340 2100
rect 18320 2030 18340 2050
rect 18320 1980 18340 2000
rect 18375 2230 18395 2250
rect 18375 2180 18395 2200
rect 18375 2130 18395 2150
rect 18375 2080 18395 2100
rect 18375 2030 18395 2050
rect 18375 1980 18395 2000
rect 18430 2230 18450 2250
rect 18430 2180 18450 2200
rect 18430 2130 18450 2150
rect 18430 2080 18450 2100
rect 18430 2030 18450 2050
rect 18430 1980 18450 2000
rect 18485 2230 18505 2250
rect 18485 2180 18505 2200
rect 18485 2130 18505 2150
rect 18485 2080 18505 2100
rect 18485 2030 18505 2050
rect 18485 1980 18505 2000
rect 18540 2230 18560 2250
rect 18540 2180 18560 2200
rect 18540 2130 18560 2150
rect 18540 2080 18560 2100
rect 18540 2030 18560 2050
rect 18540 1980 18560 2000
rect 18595 2230 18615 2250
rect 18595 2180 18615 2200
rect 18595 2130 18615 2150
rect 18595 2080 18615 2100
rect 18595 2030 18615 2050
rect 18595 1980 18615 2000
rect 18650 2230 18670 2250
rect 18650 2180 18670 2200
rect 18650 2130 18670 2150
rect 18650 2080 18670 2100
rect 18650 2030 18670 2050
rect 18650 1980 18670 2000
rect 18705 2230 18725 2250
rect 18705 2180 18725 2200
rect 18705 2130 18725 2150
rect 18705 2080 18725 2100
rect 18705 2030 18725 2050
rect 18705 1980 18725 2000
rect 18760 2230 18780 2250
rect 18760 2180 18780 2200
rect 18760 2130 18780 2150
rect 18760 2080 18780 2100
rect 18760 2030 18780 2050
rect 18760 1980 18780 2000
rect 18815 2230 18835 2250
rect 18815 2180 18835 2200
rect 18815 2130 18835 2150
rect 18815 2080 18835 2100
rect 18815 2030 18835 2050
rect 25015 2230 25035 2250
rect 25015 2180 25035 2200
rect 25015 2130 25035 2150
rect 25015 2080 25035 2100
rect 25015 2030 25035 2050
rect 18815 1980 18835 2000
rect 25015 1980 25035 2000
rect 25070 2230 25090 2250
rect 25070 2180 25090 2200
rect 25070 2130 25090 2150
rect 25070 2080 25090 2100
rect 25070 2030 25090 2050
rect 25070 1980 25090 2000
rect 25125 2230 25145 2250
rect 25125 2180 25145 2200
rect 25125 2130 25145 2150
rect 25125 2080 25145 2100
rect 25125 2030 25145 2050
rect 25125 1980 25145 2000
rect 25180 2230 25200 2250
rect 25180 2180 25200 2200
rect 25180 2130 25200 2150
rect 25180 2080 25200 2100
rect 25180 2030 25200 2050
rect 25180 1980 25200 2000
rect 25235 2230 25255 2250
rect 25235 2180 25255 2200
rect 25235 2130 25255 2150
rect 25235 2080 25255 2100
rect 25235 2030 25255 2050
rect 25235 1980 25255 2000
rect 25290 2230 25310 2250
rect 25290 2180 25310 2200
rect 25290 2130 25310 2150
rect 25290 2080 25310 2100
rect 25290 2030 25310 2050
rect 25290 1980 25310 2000
rect 25345 2230 25365 2250
rect 25345 2180 25365 2200
rect 25345 2130 25365 2150
rect 25345 2080 25365 2100
rect 25345 2030 25365 2050
rect 25345 1980 25365 2000
rect 25400 2230 25420 2250
rect 25400 2180 25420 2200
rect 25400 2130 25420 2150
rect 25400 2080 25420 2100
rect 25400 2030 25420 2050
rect 25400 1980 25420 2000
rect 25455 2230 25475 2250
rect 25455 2180 25475 2200
rect 25455 2130 25475 2150
rect 25455 2080 25475 2100
rect 25455 2030 25475 2050
rect 25455 1980 25475 2000
rect 25510 2230 25530 2250
rect 25510 2180 25530 2200
rect 25510 2130 25530 2150
rect 25510 2080 25530 2100
rect 25510 2030 25530 2050
rect 25510 1980 25530 2000
rect 25565 2230 25585 2250
rect 25565 2180 25585 2200
rect 25565 2130 25585 2150
rect 25565 2080 25585 2100
rect 25565 2030 25585 2050
rect 25565 1980 25585 2000
rect 25620 2230 25640 2250
rect 25620 2180 25640 2200
rect 25620 2130 25640 2150
rect 25620 2080 25640 2100
rect 25620 2030 25640 2050
rect 25620 1980 25640 2000
rect 25675 2230 25695 2250
rect 25675 2180 25695 2200
rect 25675 2130 25695 2150
rect 25675 2080 25695 2100
rect 25675 2030 25695 2050
rect 25675 1980 25695 2000
rect 26285 2095 26305 2115
rect 26285 2045 26305 2065
rect 26285 1995 26305 2015
rect 26340 2095 26360 2115
rect 26340 2045 26360 2065
rect 26340 1995 26360 2015
rect 26395 2095 26415 2115
rect 26395 2045 26415 2065
rect 26395 1995 26415 2015
rect 26450 2095 26470 2115
rect 26450 2045 26470 2065
rect 26450 1995 26470 2015
rect 26505 2095 26525 2115
rect 26505 2045 26525 2065
rect 26505 1995 26525 2015
rect 26560 2095 26580 2115
rect 26560 2045 26580 2065
rect 26560 1995 26580 2015
rect 26615 2095 26635 2115
rect 26615 2045 26635 2065
rect 26615 1995 26635 2015
rect 26670 2095 26690 2115
rect 26670 2045 26690 2065
rect 26670 1995 26690 2015
rect 26725 2095 26745 2115
rect 26725 2045 26745 2065
rect 26725 1995 26745 2015
rect 26780 2095 26800 2115
rect 26780 2045 26800 2065
rect 26780 1995 26800 2015
rect 26835 2095 26855 2115
rect 26835 2045 26855 2065
rect 26835 1995 26855 2015
rect 26890 2095 26910 2115
rect 26890 2045 26910 2065
rect 26890 1995 26910 2015
rect 26945 2095 26965 2115
rect 26945 2045 26965 2065
rect 26945 1995 26965 2015
rect 27000 2095 27020 2115
rect 27000 2045 27020 2065
rect 27000 1995 27020 2015
rect 27055 2095 27075 2115
rect 27055 2045 27075 2065
rect 27055 1995 27075 2015
rect 27110 2095 27130 2115
rect 27110 2045 27130 2065
rect 27110 1995 27130 2015
rect 27165 2095 27185 2115
rect 27165 2045 27185 2065
rect 27165 1995 27185 2015
rect 27220 2095 27240 2115
rect 27220 2045 27240 2065
rect 27220 1995 27240 2015
rect 27275 2095 27295 2115
rect 27275 2045 27295 2065
rect 27275 1995 27295 2015
rect 27330 2095 27350 2115
rect 27330 2045 27350 2065
rect 27330 1995 27350 2015
rect 27385 2095 27405 2115
rect 27385 2045 27405 2065
rect 27385 1995 27405 2015
rect 27440 2095 27460 2115
rect 27440 2045 27460 2065
rect 27440 1995 27460 2015
rect 27495 2095 27515 2115
rect 27495 2045 27515 2065
rect 27495 1995 27515 2015
rect 28155 2210 28175 2230
rect 28155 2160 28175 2180
rect 28155 2110 28175 2130
rect 28155 2060 28175 2080
rect 28155 2010 28175 2030
rect 28155 1960 28175 1980
rect 28210 2210 28230 2230
rect 28210 2160 28230 2180
rect 28210 2110 28230 2130
rect 28210 2060 28230 2080
rect 28210 2010 28230 2030
rect 28210 1960 28230 1980
rect 28265 2210 28285 2230
rect 28265 2160 28285 2180
rect 28265 2110 28285 2130
rect 28265 2060 28285 2080
rect 28265 2010 28285 2030
rect 28265 1960 28285 1980
rect 28320 2210 28340 2230
rect 28320 2160 28340 2180
rect 28320 2110 28340 2130
rect 28320 2060 28340 2080
rect 28320 2010 28340 2030
rect 28320 1960 28340 1980
rect 28375 2210 28395 2230
rect 28375 2160 28395 2180
rect 28375 2110 28395 2130
rect 28375 2060 28395 2080
rect 28375 2010 28395 2030
rect 28375 1960 28395 1980
rect 28430 2210 28450 2230
rect 28430 2160 28450 2180
rect 28430 2110 28450 2130
rect 28430 2060 28450 2080
rect 28430 2010 28450 2030
rect 28430 1960 28450 1980
rect 28485 2210 28505 2230
rect 28485 2160 28505 2180
rect 28485 2110 28505 2130
rect 28485 2060 28505 2080
rect 28485 2010 28505 2030
rect 28485 1960 28505 1980
rect 28540 2210 28560 2230
rect 28540 2160 28560 2180
rect 28540 2110 28560 2130
rect 28540 2060 28560 2080
rect 28540 2010 28560 2030
rect 28540 1960 28560 1980
rect 28595 2210 28615 2230
rect 28595 2160 28615 2180
rect 28595 2110 28615 2130
rect 28595 2060 28615 2080
rect 28595 2010 28615 2030
rect 28595 1960 28615 1980
rect 28650 2210 28670 2230
rect 28650 2160 28670 2180
rect 28650 2110 28670 2130
rect 28650 2060 28670 2080
rect 28650 2010 28670 2030
rect 28650 1960 28670 1980
rect 28705 2210 28725 2230
rect 28705 2160 28725 2180
rect 28705 2110 28725 2130
rect 28705 2060 28725 2080
rect 28705 2010 28725 2030
rect 28705 1960 28725 1980
rect 28760 2210 28780 2230
rect 28760 2160 28780 2180
rect 28760 2110 28780 2130
rect 28760 2060 28780 2080
rect 28760 2010 28780 2030
rect 28760 1960 28780 1980
rect 28815 2210 28835 2230
rect 28815 2160 28835 2180
rect 28815 2110 28835 2130
rect 28815 2060 28835 2080
rect 28815 2010 28835 2030
rect 28815 1960 28835 1980
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 4815 1630 4835 1650
rect 15015 1620 15035 1640
rect 2845 1420 2865 1440
rect 2845 1370 2865 1390
rect 2845 1320 2865 1340
rect 2845 1270 2865 1290
rect 2845 1220 2865 1240
rect 3385 1420 3405 1440
rect 3385 1370 3405 1390
rect 3385 1320 3405 1340
rect 3385 1270 3405 1290
rect 3385 1220 3405 1240
rect 3925 1420 3945 1440
rect 3925 1370 3945 1390
rect 3925 1320 3945 1340
rect 3925 1270 3945 1290
rect 3925 1220 3945 1240
rect 4065 1420 4085 1440
rect 4065 1370 4085 1390
rect 4065 1320 4085 1340
rect 4065 1270 4085 1290
rect 4065 1220 4085 1240
rect 4605 1420 4625 1440
rect 4605 1370 4625 1390
rect 4605 1320 4625 1340
rect 4605 1270 4625 1290
rect 4605 1220 4625 1240
rect 5145 1420 5165 1440
rect 5145 1370 5165 1390
rect 5145 1320 5165 1340
rect 5145 1270 5165 1290
rect 5145 1220 5165 1240
rect 2955 1040 2975 1060
rect 2955 990 2975 1010
rect 3995 1040 4015 1060
rect 3995 990 4015 1010
rect 5035 1040 5055 1060
rect 5035 990 5055 1010
rect 15015 1570 15035 1590
rect 15015 1520 15035 1540
rect 15015 1470 15035 1490
rect 15015 1420 15035 1440
rect 15015 1370 15035 1390
rect 15015 1320 15035 1340
rect 15015 1270 15035 1290
rect 15015 1220 15035 1240
rect 15015 1170 15035 1190
rect 15015 1120 15035 1140
rect 15015 1070 15035 1090
rect 15015 1020 15035 1040
rect 15015 970 15035 990
rect 15115 1620 15135 1640
rect 15115 1570 15135 1590
rect 15115 1520 15135 1540
rect 15115 1470 15135 1490
rect 15115 1420 15135 1440
rect 15115 1370 15135 1390
rect 15115 1320 15135 1340
rect 15115 1270 15135 1290
rect 15115 1220 15135 1240
rect 15115 1170 15135 1190
rect 15115 1120 15135 1140
rect 15115 1070 15135 1090
rect 15115 1020 15135 1040
rect 15115 970 15135 990
rect 15215 1620 15235 1640
rect 15215 1570 15235 1590
rect 15215 1520 15235 1540
rect 15215 1470 15235 1490
rect 15215 1420 15235 1440
rect 15215 1370 15235 1390
rect 15215 1320 15235 1340
rect 15215 1270 15235 1290
rect 15215 1220 15235 1240
rect 15215 1170 15235 1190
rect 15215 1120 15235 1140
rect 15215 1070 15235 1090
rect 15215 1020 15235 1040
rect 15215 970 15235 990
rect 15315 1620 15335 1640
rect 15315 1570 15335 1590
rect 15315 1520 15335 1540
rect 15315 1470 15335 1490
rect 15315 1420 15335 1440
rect 15315 1370 15335 1390
rect 15315 1320 15335 1340
rect 15315 1270 15335 1290
rect 15315 1220 15335 1240
rect 15315 1170 15335 1190
rect 15315 1120 15335 1140
rect 15315 1070 15335 1090
rect 15315 1020 15335 1040
rect 15315 970 15335 990
rect 15415 1620 15435 1640
rect 15415 1570 15435 1590
rect 15415 1520 15435 1540
rect 15415 1470 15435 1490
rect 15415 1420 15435 1440
rect 15415 1370 15435 1390
rect 15415 1320 15435 1340
rect 15415 1270 15435 1290
rect 15415 1220 15435 1240
rect 15415 1170 15435 1190
rect 15415 1120 15435 1140
rect 15415 1070 15435 1090
rect 15415 1020 15435 1040
rect 15415 970 15435 990
rect 15515 1620 15535 1640
rect 15515 1570 15535 1590
rect 15515 1520 15535 1540
rect 15515 1470 15535 1490
rect 15515 1420 15535 1440
rect 15515 1370 15535 1390
rect 15515 1320 15535 1340
rect 15515 1270 15535 1290
rect 15515 1220 15535 1240
rect 15515 1170 15535 1190
rect 15515 1120 15535 1140
rect 15515 1070 15535 1090
rect 15515 1020 15535 1040
rect 15515 970 15535 990
rect 15615 1620 15635 1640
rect 15615 1570 15635 1590
rect 15615 1520 15635 1540
rect 16040 1630 16060 1650
rect 16040 1580 16060 1600
rect 16040 1530 16060 1550
rect 16095 1630 16115 1650
rect 16095 1580 16115 1600
rect 16095 1530 16115 1550
rect 16150 1630 16170 1650
rect 16150 1580 16170 1600
rect 16150 1530 16170 1550
rect 16205 1630 16225 1650
rect 16205 1580 16225 1600
rect 16205 1530 16225 1550
rect 16260 1630 16280 1650
rect 16260 1580 16280 1600
rect 16260 1530 16280 1550
rect 16315 1630 16335 1650
rect 16315 1580 16335 1600
rect 16315 1530 16335 1550
rect 16370 1630 16390 1650
rect 16370 1580 16390 1600
rect 16370 1530 16390 1550
rect 16425 1630 16445 1650
rect 16425 1580 16445 1600
rect 16425 1530 16445 1550
rect 16480 1630 16500 1650
rect 16480 1580 16500 1600
rect 16480 1530 16500 1550
rect 16535 1630 16555 1650
rect 16535 1580 16555 1600
rect 16535 1530 16555 1550
rect 16590 1630 16610 1650
rect 16590 1580 16610 1600
rect 16590 1530 16610 1550
rect 16645 1630 16665 1650
rect 16645 1580 16665 1600
rect 16645 1530 16665 1550
rect 16700 1630 16720 1650
rect 16780 1630 16800 1650
rect 16700 1580 16720 1600
rect 16780 1580 16800 1600
rect 16700 1530 16720 1550
rect 16780 1530 16800 1550
rect 16835 1630 16855 1650
rect 16835 1580 16855 1600
rect 16835 1530 16855 1550
rect 16890 1630 16910 1650
rect 16890 1580 16910 1600
rect 16890 1530 16910 1550
rect 16945 1630 16965 1650
rect 16945 1580 16965 1600
rect 16945 1530 16965 1550
rect 17000 1630 17020 1650
rect 17080 1630 17100 1650
rect 17000 1580 17020 1600
rect 17080 1580 17100 1600
rect 17000 1530 17020 1550
rect 17080 1530 17100 1550
rect 17135 1630 17155 1650
rect 17135 1580 17155 1600
rect 17135 1530 17155 1550
rect 17190 1630 17210 1650
rect 17190 1580 17210 1600
rect 17190 1530 17210 1550
rect 17245 1630 17265 1650
rect 17245 1580 17265 1600
rect 17245 1530 17265 1550
rect 17300 1630 17320 1650
rect 17300 1580 17320 1600
rect 17300 1530 17320 1550
rect 17355 1630 17375 1650
rect 17355 1580 17375 1600
rect 17355 1530 17375 1550
rect 17410 1630 17430 1650
rect 17410 1580 17430 1600
rect 17410 1530 17430 1550
rect 17465 1630 17485 1650
rect 17465 1580 17485 1600
rect 17465 1530 17485 1550
rect 17520 1630 17540 1650
rect 17520 1580 17540 1600
rect 17520 1530 17540 1550
rect 17575 1630 17595 1650
rect 17575 1580 17595 1600
rect 17575 1530 17595 1550
rect 17630 1630 17650 1650
rect 17630 1580 17650 1600
rect 17630 1530 17650 1550
rect 17685 1630 17705 1650
rect 17685 1580 17705 1600
rect 17685 1530 17705 1550
rect 17740 1630 17760 1650
rect 17740 1580 17760 1600
rect 17740 1530 17760 1550
rect 18215 1620 18235 1640
rect 18215 1570 18235 1590
rect 18215 1520 18235 1540
rect 15615 1470 15635 1490
rect 18215 1470 18235 1490
rect 15615 1420 15635 1440
rect 15615 1370 15635 1390
rect 15615 1320 15635 1340
rect 15615 1270 15635 1290
rect 18215 1420 18235 1440
rect 18215 1370 18235 1390
rect 18215 1320 18235 1340
rect 18215 1270 18235 1290
rect 15615 1220 15635 1240
rect 15615 1170 15635 1190
rect 18215 1220 18235 1240
rect 15615 1120 15635 1140
rect 15615 1070 15635 1090
rect 15615 1020 15635 1040
rect 15615 970 15635 990
rect 16215 1150 16235 1170
rect 16215 1100 16235 1120
rect 16215 1050 16235 1070
rect 16215 1000 16235 1020
rect 16215 950 16235 970
rect 16270 1150 16290 1170
rect 16270 1100 16290 1120
rect 16270 1050 16290 1070
rect 16270 1000 16290 1020
rect 16270 950 16290 970
rect 16325 1150 16345 1170
rect 16325 1100 16345 1120
rect 16325 1050 16345 1070
rect 16325 1000 16345 1020
rect 16325 950 16345 970
rect 16380 1150 16400 1170
rect 16380 1100 16400 1120
rect 16380 1050 16400 1070
rect 16380 1000 16400 1020
rect 16380 950 16400 970
rect 16435 1150 16455 1170
rect 16435 1100 16455 1120
rect 16435 1050 16455 1070
rect 16435 1000 16455 1020
rect 16435 950 16455 970
rect 16490 1150 16510 1170
rect 16490 1100 16510 1120
rect 16490 1050 16510 1070
rect 16490 1000 16510 1020
rect 16490 950 16510 970
rect 16545 1150 16565 1170
rect 16545 1100 16565 1120
rect 16545 1050 16565 1070
rect 16545 1000 16565 1020
rect 16545 950 16565 970
rect 16600 1150 16620 1170
rect 16600 1100 16620 1120
rect 16600 1050 16620 1070
rect 16600 1000 16620 1020
rect 16600 950 16620 970
rect 16655 1150 16675 1170
rect 16655 1100 16675 1120
rect 16655 1050 16675 1070
rect 16655 1000 16675 1020
rect 16655 950 16675 970
rect 16710 1150 16730 1170
rect 16710 1100 16730 1120
rect 16710 1050 16730 1070
rect 16710 1000 16730 1020
rect 16710 950 16730 970
rect 16765 1150 16785 1170
rect 16765 1100 16785 1120
rect 16765 1050 16785 1070
rect 16765 1000 16785 1020
rect 16765 950 16785 970
rect 16820 1150 16840 1170
rect 16820 1100 16840 1120
rect 16820 1050 16840 1070
rect 16820 1000 16840 1020
rect 16820 950 16840 970
rect 16875 1150 16895 1170
rect 16875 1100 16895 1120
rect 16875 1050 16895 1070
rect 16875 1000 16895 1020
rect 16875 950 16895 970
rect 16930 1150 16950 1170
rect 16930 1100 16950 1120
rect 16930 1050 16950 1070
rect 16930 1000 16950 1020
rect 16930 950 16950 970
rect 16985 1150 17005 1170
rect 16985 1100 17005 1120
rect 16985 1050 17005 1070
rect 16985 1000 17005 1020
rect 16985 950 17005 970
rect 17040 1150 17060 1170
rect 17040 1100 17060 1120
rect 17040 1050 17060 1070
rect 17040 1000 17060 1020
rect 17040 950 17060 970
rect 17095 1150 17115 1170
rect 17095 1100 17115 1120
rect 17095 1050 17115 1070
rect 17095 1000 17115 1020
rect 17095 950 17115 970
rect 17150 1150 17170 1170
rect 17150 1100 17170 1120
rect 17150 1050 17170 1070
rect 17150 1000 17170 1020
rect 17150 950 17170 970
rect 17205 1150 17225 1170
rect 17205 1100 17225 1120
rect 17205 1050 17225 1070
rect 17205 1000 17225 1020
rect 17205 950 17225 970
rect 17260 1150 17280 1170
rect 17260 1100 17280 1120
rect 17260 1050 17280 1070
rect 17260 1000 17280 1020
rect 17260 950 17280 970
rect 17315 1150 17335 1170
rect 17315 1100 17335 1120
rect 17315 1050 17335 1070
rect 17315 1000 17335 1020
rect 17315 950 17335 970
rect 17370 1150 17390 1170
rect 17370 1100 17390 1120
rect 17370 1050 17390 1070
rect 17370 1000 17390 1020
rect 17370 950 17390 970
rect 17425 1150 17445 1170
rect 17425 1100 17445 1120
rect 17425 1050 17445 1070
rect 17425 1000 17445 1020
rect 17425 950 17445 970
rect 17480 1150 17500 1170
rect 17480 1100 17500 1120
rect 17480 1050 17500 1070
rect 17480 1000 17500 1020
rect 17480 950 17500 970
rect 17535 1150 17555 1170
rect 17535 1100 17555 1120
rect 17535 1050 17555 1070
rect 17535 1000 17555 1020
rect 17535 950 17555 970
rect 17590 1150 17610 1170
rect 17590 1100 17610 1120
rect 17590 1050 17610 1070
rect 17590 1000 17610 1020
rect 17590 950 17610 970
rect 18215 1170 18235 1190
rect 18215 1120 18235 1140
rect 18215 1070 18235 1090
rect 18215 1020 18235 1040
rect 18215 970 18235 990
rect 18315 1620 18335 1640
rect 18315 1570 18335 1590
rect 18315 1520 18335 1540
rect 18315 1470 18335 1490
rect 18315 1420 18335 1440
rect 18315 1370 18335 1390
rect 18315 1320 18335 1340
rect 18315 1270 18335 1290
rect 18315 1220 18335 1240
rect 18315 1170 18335 1190
rect 18315 1120 18335 1140
rect 18315 1070 18335 1090
rect 18315 1020 18335 1040
rect 18315 970 18335 990
rect 18415 1620 18435 1640
rect 18415 1570 18435 1590
rect 18415 1520 18435 1540
rect 18415 1470 18435 1490
rect 18415 1420 18435 1440
rect 18415 1370 18435 1390
rect 18415 1320 18435 1340
rect 18415 1270 18435 1290
rect 18415 1220 18435 1240
rect 18415 1170 18435 1190
rect 18415 1120 18435 1140
rect 18415 1070 18435 1090
rect 18415 1020 18435 1040
rect 18415 970 18435 990
rect 18515 1620 18535 1640
rect 18515 1570 18535 1590
rect 18515 1520 18535 1540
rect 18515 1470 18535 1490
rect 18515 1420 18535 1440
rect 18515 1370 18535 1390
rect 18515 1320 18535 1340
rect 18515 1270 18535 1290
rect 18515 1220 18535 1240
rect 18515 1170 18535 1190
rect 18515 1120 18535 1140
rect 18515 1070 18535 1090
rect 18515 1020 18535 1040
rect 18515 970 18535 990
rect 18615 1620 18635 1640
rect 18615 1570 18635 1590
rect 18615 1520 18635 1540
rect 18615 1470 18635 1490
rect 18615 1420 18635 1440
rect 18615 1370 18635 1390
rect 18615 1320 18635 1340
rect 18615 1270 18635 1290
rect 18615 1220 18635 1240
rect 18615 1170 18635 1190
rect 18615 1120 18635 1140
rect 18615 1070 18635 1090
rect 18615 1020 18635 1040
rect 18615 970 18635 990
rect 18715 1620 18735 1640
rect 18715 1570 18735 1590
rect 18715 1520 18735 1540
rect 18715 1470 18735 1490
rect 18715 1420 18735 1440
rect 18715 1370 18735 1390
rect 18715 1320 18735 1340
rect 18715 1270 18735 1290
rect 18715 1220 18735 1240
rect 18715 1170 18735 1190
rect 18715 1120 18735 1140
rect 18715 1070 18735 1090
rect 18715 1020 18735 1040
rect 18715 970 18735 990
rect 18815 1620 18835 1640
rect 25015 1620 25035 1640
rect 18815 1570 18835 1590
rect 18815 1520 18835 1540
rect 18815 1470 18835 1490
rect 18815 1420 18835 1440
rect 18815 1370 18835 1390
rect 18815 1320 18835 1340
rect 18815 1270 18835 1290
rect 18815 1220 18835 1240
rect 18815 1170 18835 1190
rect 18815 1120 18835 1140
rect 18815 1070 18835 1090
rect 18815 1020 18835 1040
rect 18815 970 18835 990
rect 25015 1570 25035 1590
rect 25015 1520 25035 1540
rect 25015 1470 25035 1490
rect 25015 1420 25035 1440
rect 25015 1370 25035 1390
rect 25015 1320 25035 1340
rect 25015 1270 25035 1290
rect 25015 1220 25035 1240
rect 25015 1170 25035 1190
rect 25015 1120 25035 1140
rect 25015 1070 25035 1090
rect 25015 1020 25035 1040
rect 25015 970 25035 990
rect 25115 1620 25135 1640
rect 25115 1570 25135 1590
rect 25115 1520 25135 1540
rect 25115 1470 25135 1490
rect 25115 1420 25135 1440
rect 25115 1370 25135 1390
rect 25115 1320 25135 1340
rect 25115 1270 25135 1290
rect 25115 1220 25135 1240
rect 25115 1170 25135 1190
rect 25115 1120 25135 1140
rect 25115 1070 25135 1090
rect 25115 1020 25135 1040
rect 25115 970 25135 990
rect 25215 1620 25235 1640
rect 25215 1570 25235 1590
rect 25215 1520 25235 1540
rect 25215 1470 25235 1490
rect 25215 1420 25235 1440
rect 25215 1370 25235 1390
rect 25215 1320 25235 1340
rect 25215 1270 25235 1290
rect 25215 1220 25235 1240
rect 25215 1170 25235 1190
rect 25215 1120 25235 1140
rect 25215 1070 25235 1090
rect 25215 1020 25235 1040
rect 25215 970 25235 990
rect 25315 1620 25335 1640
rect 25315 1570 25335 1590
rect 25315 1520 25335 1540
rect 25315 1470 25335 1490
rect 25315 1420 25335 1440
rect 25315 1370 25335 1390
rect 25315 1320 25335 1340
rect 25315 1270 25335 1290
rect 25315 1220 25335 1240
rect 25315 1170 25335 1190
rect 25315 1120 25335 1140
rect 25315 1070 25335 1090
rect 25315 1020 25335 1040
rect 25315 970 25335 990
rect 25415 1620 25435 1640
rect 25415 1570 25435 1590
rect 25415 1520 25435 1540
rect 25415 1470 25435 1490
rect 25415 1420 25435 1440
rect 25415 1370 25435 1390
rect 25415 1320 25435 1340
rect 25415 1270 25435 1290
rect 25415 1220 25435 1240
rect 25415 1170 25435 1190
rect 25415 1120 25435 1140
rect 25415 1070 25435 1090
rect 25415 1020 25435 1040
rect 25415 970 25435 990
rect 25515 1620 25535 1640
rect 25515 1570 25535 1590
rect 25515 1520 25535 1540
rect 25515 1470 25535 1490
rect 25515 1420 25535 1440
rect 25515 1370 25535 1390
rect 25515 1320 25535 1340
rect 25515 1270 25535 1290
rect 25515 1220 25535 1240
rect 25515 1170 25535 1190
rect 25515 1120 25535 1140
rect 25515 1070 25535 1090
rect 25515 1020 25535 1040
rect 25515 970 25535 990
rect 25615 1620 25635 1640
rect 25615 1570 25635 1590
rect 25615 1520 25635 1540
rect 25615 1470 25635 1490
rect 25615 1420 25635 1440
rect 25615 1370 25635 1390
rect 26040 1630 26060 1650
rect 26040 1580 26060 1600
rect 26040 1530 26060 1550
rect 26095 1630 26115 1650
rect 26095 1580 26115 1600
rect 26095 1530 26115 1550
rect 26150 1630 26170 1650
rect 26150 1580 26170 1600
rect 26150 1530 26170 1550
rect 26205 1630 26225 1650
rect 26205 1580 26225 1600
rect 26205 1530 26225 1550
rect 26260 1630 26280 1650
rect 26260 1580 26280 1600
rect 26260 1530 26280 1550
rect 26315 1630 26335 1650
rect 26315 1580 26335 1600
rect 26315 1530 26335 1550
rect 26370 1630 26390 1650
rect 26370 1580 26390 1600
rect 26370 1530 26390 1550
rect 26425 1630 26445 1650
rect 26425 1580 26445 1600
rect 26425 1530 26445 1550
rect 26480 1630 26500 1650
rect 26480 1580 26500 1600
rect 26480 1530 26500 1550
rect 26535 1630 26555 1650
rect 26535 1580 26555 1600
rect 26535 1530 26555 1550
rect 26590 1630 26610 1650
rect 26590 1580 26610 1600
rect 26590 1530 26610 1550
rect 26645 1630 26665 1650
rect 26645 1580 26665 1600
rect 26645 1530 26665 1550
rect 26700 1630 26720 1650
rect 26780 1630 26800 1650
rect 26700 1580 26720 1600
rect 26780 1580 26800 1600
rect 26700 1530 26720 1550
rect 26780 1530 26800 1550
rect 26835 1630 26855 1650
rect 26835 1580 26855 1600
rect 26835 1530 26855 1550
rect 26890 1630 26910 1650
rect 26890 1580 26910 1600
rect 26890 1530 26910 1550
rect 26945 1630 26965 1650
rect 26945 1580 26965 1600
rect 26945 1530 26965 1550
rect 27000 1630 27020 1650
rect 27080 1630 27100 1650
rect 27000 1580 27020 1600
rect 27080 1580 27100 1600
rect 27000 1530 27020 1550
rect 27080 1530 27100 1550
rect 27135 1630 27155 1650
rect 27135 1580 27155 1600
rect 27135 1530 27155 1550
rect 27190 1630 27210 1650
rect 27190 1580 27210 1600
rect 27190 1530 27210 1550
rect 27245 1630 27265 1650
rect 27245 1580 27265 1600
rect 27245 1530 27265 1550
rect 27300 1630 27320 1650
rect 27300 1580 27320 1600
rect 27300 1530 27320 1550
rect 27355 1630 27375 1650
rect 27355 1580 27375 1600
rect 27355 1530 27375 1550
rect 27410 1630 27430 1650
rect 27410 1580 27430 1600
rect 27410 1530 27430 1550
rect 27465 1630 27485 1650
rect 27465 1580 27485 1600
rect 27465 1530 27485 1550
rect 27520 1630 27540 1650
rect 27520 1580 27540 1600
rect 27520 1530 27540 1550
rect 27575 1630 27595 1650
rect 27575 1580 27595 1600
rect 27575 1530 27595 1550
rect 27630 1630 27650 1650
rect 27630 1580 27650 1600
rect 27630 1530 27650 1550
rect 27685 1630 27705 1650
rect 27685 1580 27705 1600
rect 27685 1530 27705 1550
rect 27740 1630 27760 1650
rect 27740 1580 27760 1600
rect 27740 1530 27760 1550
rect 25615 1320 25635 1340
rect 25615 1270 25635 1290
rect 25615 1220 25635 1240
rect 25615 1170 25635 1190
rect 25615 1120 25635 1140
rect 25615 1070 25635 1090
rect 25615 1020 25635 1040
rect 25615 970 25635 990
rect 3005 845 3025 865
rect 3005 795 3025 815
rect 3095 845 3115 865
rect 3095 795 3115 815
rect 3185 845 3205 865
rect 3185 795 3205 815
rect 3275 845 3295 865
rect 3275 795 3295 815
rect 3365 845 3385 865
rect 3365 795 3385 815
rect 3455 845 3475 865
rect 3455 795 3475 815
rect 3545 845 3565 865
rect 3545 795 3565 815
rect 3635 845 3655 865
rect 3635 795 3655 815
rect 3725 845 3745 865
rect 3725 795 3745 815
rect 3815 845 3835 865
rect 3815 795 3835 815
rect 3905 845 3925 865
rect 3905 795 3925 815
rect 3995 845 4015 865
rect 3995 795 4015 815
rect 4085 845 4105 865
rect 4085 795 4105 815
rect 4175 845 4195 865
rect 4175 795 4195 815
rect 4265 845 4285 865
rect 4265 795 4285 815
rect 4355 845 4375 865
rect 4355 795 4375 815
rect 4445 845 4465 865
rect 4445 795 4465 815
rect 4535 845 4555 865
rect 4535 795 4555 815
rect 4625 845 4645 865
rect 4625 795 4645 815
rect 4715 845 4735 865
rect 4715 795 4735 815
rect 4805 845 4825 865
rect 4805 795 4825 815
rect 4895 845 4915 865
rect 4895 795 4915 815
rect 4985 845 5005 865
rect 4985 795 5005 815
rect 26215 1050 26235 1070
rect 26215 1000 26235 1020
rect 26215 950 26235 970
rect 26215 900 26235 920
rect 26215 850 26235 870
rect 26270 1050 26290 1070
rect 26270 1000 26290 1020
rect 26270 950 26290 970
rect 26270 900 26290 920
rect 26270 850 26290 870
rect 26325 1050 26345 1070
rect 26325 1000 26345 1020
rect 26325 950 26345 970
rect 26325 900 26345 920
rect 26325 850 26345 870
rect 26380 1050 26400 1070
rect 26380 1000 26400 1020
rect 26380 950 26400 970
rect 26380 900 26400 920
rect 26380 850 26400 870
rect 26435 1050 26455 1070
rect 26435 1000 26455 1020
rect 26435 950 26455 970
rect 26435 900 26455 920
rect 26435 850 26455 870
rect 26490 1050 26510 1070
rect 26490 1000 26510 1020
rect 26490 950 26510 970
rect 26490 900 26510 920
rect 26490 850 26510 870
rect 26545 1050 26565 1070
rect 26545 1000 26565 1020
rect 26545 950 26565 970
rect 26545 900 26565 920
rect 26545 850 26565 870
rect 26600 1050 26620 1070
rect 26600 1000 26620 1020
rect 26600 950 26620 970
rect 26600 900 26620 920
rect 26600 850 26620 870
rect 26655 1050 26675 1070
rect 26655 1000 26675 1020
rect 26655 950 26675 970
rect 26655 900 26675 920
rect 26655 850 26675 870
rect 26710 1050 26730 1070
rect 26710 1000 26730 1020
rect 26710 950 26730 970
rect 26710 900 26730 920
rect 26710 850 26730 870
rect 26765 1050 26785 1070
rect 26765 1000 26785 1020
rect 26765 950 26785 970
rect 26765 900 26785 920
rect 26765 850 26785 870
rect 26820 1050 26840 1070
rect 26820 1000 26840 1020
rect 26820 950 26840 970
rect 26820 900 26840 920
rect 26820 850 26840 870
rect 26875 1050 26895 1070
rect 26875 1000 26895 1020
rect 26875 950 26895 970
rect 26875 900 26895 920
rect 26875 850 26895 870
rect 26930 1050 26950 1070
rect 26930 1000 26950 1020
rect 26930 950 26950 970
rect 26930 900 26950 920
rect 26930 850 26950 870
rect 26985 1050 27005 1070
rect 26985 1000 27005 1020
rect 26985 950 27005 970
rect 26985 900 27005 920
rect 26985 850 27005 870
rect 27040 1050 27060 1070
rect 27040 1000 27060 1020
rect 27040 950 27060 970
rect 27040 900 27060 920
rect 27040 850 27060 870
rect 27095 1050 27115 1070
rect 27095 1000 27115 1020
rect 27095 950 27115 970
rect 27095 900 27115 920
rect 27095 850 27115 870
rect 27150 1050 27170 1070
rect 27150 1000 27170 1020
rect 27150 950 27170 970
rect 27150 900 27170 920
rect 27150 850 27170 870
rect 27205 1050 27225 1070
rect 27205 1000 27225 1020
rect 27205 950 27225 970
rect 27205 900 27225 920
rect 27205 850 27225 870
rect 27260 1050 27280 1070
rect 27260 1000 27280 1020
rect 27260 950 27280 970
rect 27260 900 27280 920
rect 27260 850 27280 870
rect 27315 1050 27335 1070
rect 27315 1000 27335 1020
rect 27315 950 27335 970
rect 27315 900 27335 920
rect 27315 850 27335 870
rect 27370 1050 27390 1070
rect 27370 1000 27390 1020
rect 27370 950 27390 970
rect 27370 900 27390 920
rect 27370 850 27390 870
rect 27425 1050 27445 1070
rect 27425 1000 27445 1020
rect 27425 950 27445 970
rect 27425 900 27445 920
rect 27425 850 27445 870
rect 27480 1050 27500 1070
rect 27480 1000 27500 1020
rect 27480 950 27500 970
rect 27480 900 27500 920
rect 27480 850 27500 870
rect 27535 1050 27555 1070
rect 27535 1000 27555 1020
rect 27535 950 27555 970
rect 27535 900 27555 920
rect 27535 850 27555 870
rect 27590 1050 27610 1070
rect 27590 1000 27610 1020
rect 27590 950 27610 970
rect 27590 900 27610 920
rect 27590 850 27610 870
rect 28215 1620 28235 1640
rect 28215 1570 28235 1590
rect 28215 1520 28235 1540
rect 28215 1470 28235 1490
rect 28215 1420 28235 1440
rect 28215 1370 28235 1390
rect 28215 1320 28235 1340
rect 28215 1270 28235 1290
rect 28215 1220 28235 1240
rect 28215 1170 28235 1190
rect 28215 1120 28235 1140
rect 28215 1070 28235 1090
rect 28215 1020 28235 1040
rect 28215 970 28235 990
rect 28315 1620 28335 1640
rect 28315 1570 28335 1590
rect 28315 1520 28335 1540
rect 28315 1470 28335 1490
rect 28315 1420 28335 1440
rect 28315 1370 28335 1390
rect 28315 1320 28335 1340
rect 28315 1270 28335 1290
rect 28315 1220 28335 1240
rect 28315 1170 28335 1190
rect 28315 1120 28335 1140
rect 28315 1070 28335 1090
rect 28315 1020 28335 1040
rect 28315 970 28335 990
rect 28415 1620 28435 1640
rect 28415 1570 28435 1590
rect 28415 1520 28435 1540
rect 28415 1470 28435 1490
rect 28415 1420 28435 1440
rect 28415 1370 28435 1390
rect 28415 1320 28435 1340
rect 28415 1270 28435 1290
rect 28415 1220 28435 1240
rect 28415 1170 28435 1190
rect 28415 1120 28435 1140
rect 28415 1070 28435 1090
rect 28415 1020 28435 1040
rect 28415 970 28435 990
rect 28515 1620 28535 1640
rect 28515 1570 28535 1590
rect 28515 1520 28535 1540
rect 28515 1470 28535 1490
rect 28515 1420 28535 1440
rect 28515 1370 28535 1390
rect 28515 1320 28535 1340
rect 28515 1270 28535 1290
rect 28515 1220 28535 1240
rect 28515 1170 28535 1190
rect 28515 1120 28535 1140
rect 28515 1070 28535 1090
rect 28515 1020 28535 1040
rect 28515 970 28535 990
rect 28615 1620 28635 1640
rect 28615 1570 28635 1590
rect 28615 1520 28635 1540
rect 28615 1470 28635 1490
rect 28615 1420 28635 1440
rect 28615 1370 28635 1390
rect 28615 1320 28635 1340
rect 28615 1270 28635 1290
rect 28615 1220 28635 1240
rect 28615 1170 28635 1190
rect 28615 1120 28635 1140
rect 28615 1070 28635 1090
rect 28615 1020 28635 1040
rect 28615 970 28635 990
rect 28715 1620 28735 1640
rect 28715 1570 28735 1590
rect 28715 1520 28735 1540
rect 28715 1470 28735 1490
rect 28715 1420 28735 1440
rect 28715 1370 28735 1390
rect 28715 1320 28735 1340
rect 28715 1270 28735 1290
rect 28715 1220 28735 1240
rect 28715 1170 28735 1190
rect 28715 1120 28735 1140
rect 28715 1070 28735 1090
rect 28715 1020 28735 1040
rect 28715 970 28735 990
rect 28815 1620 28835 1640
rect 28815 1570 28835 1590
rect 28815 1520 28835 1540
rect 28815 1470 28835 1490
rect 28815 1420 28835 1440
rect 28815 1370 28835 1390
rect 28815 1320 28835 1340
rect 28815 1270 28835 1290
rect 28815 1220 28835 1240
rect 28815 1170 28835 1190
rect 28815 1120 28835 1140
rect 28815 1070 28835 1090
rect 28815 1020 28835 1040
rect 28815 970 28835 990
rect 16270 715 16290 735
rect 16270 665 16290 685
rect 16500 715 16520 735
rect 16890 715 16910 735
rect 16945 715 16965 735
rect 17000 715 17020 735
rect 17055 715 17075 735
rect 17110 715 17130 735
rect 17165 715 17185 735
rect 17220 715 17240 735
rect 17275 715 17295 735
rect 17330 715 17350 735
rect 17385 715 17405 735
rect 17440 715 17460 735
rect 17495 715 17515 735
rect 17550 715 17570 735
rect 16500 665 16520 685
rect 26270 515 26290 535
rect 26270 465 26290 485
rect 26500 515 26520 535
rect 26500 465 26520 485
rect 26890 515 26910 535
rect 26945 515 26965 535
rect 27000 515 27020 535
rect 27055 515 27075 535
rect 27110 515 27130 535
rect 27165 515 27185 535
rect 27220 515 27240 535
rect 27275 515 27295 535
rect 27330 515 27350 535
rect 27385 515 27405 535
rect 27440 515 27460 535
rect 27495 515 27515 535
rect 27550 515 27570 535
<< pdiffc >>
rect 26265 4810 26285 4830
rect 26325 4815 26345 4835
rect 26385 4815 26405 4835
rect 26445 4810 26465 4830
rect 26515 4825 26535 4845
rect 26575 4825 26595 4845
rect 26635 4825 26655 4845
rect 26695 4825 26715 4845
rect 26755 4825 26775 4845
rect 26815 4825 26835 4845
rect 26875 4825 26895 4845
rect 27245 4810 27265 4830
rect 27305 4810 27325 4830
rect 27365 4810 27385 4830
rect 27425 4810 27445 4830
rect 27485 4810 27505 4830
rect 27545 4810 27565 4830
rect 27605 4810 27625 4830
rect 27665 4810 27685 4830
rect 27725 4810 27745 4830
rect 16215 4305 16235 4325
rect 16275 4310 16295 4330
rect 16335 4310 16355 4330
rect 16395 4305 16415 4325
rect 16545 4320 16565 4340
rect 16605 4320 16625 4340
rect 16665 4320 16685 4340
rect 16725 4320 16745 4340
rect 16785 4320 16805 4340
rect 16845 4320 16865 4340
rect 26260 4395 26280 4415
rect 26315 4395 26335 4415
rect 26370 4395 26390 4415
rect 26425 4395 26445 4415
rect 26480 4395 26500 4415
rect 26535 4395 26555 4415
rect 26590 4395 26610 4415
rect 26645 4395 26665 4415
rect 26700 4395 26720 4415
rect 26755 4395 26775 4415
rect 26810 4395 26830 4415
rect 26865 4395 26885 4415
rect 26920 4395 26940 4415
rect 26975 4395 26995 4415
rect 27030 4395 27050 4415
rect 27085 4395 27105 4415
rect 27140 4395 27160 4415
rect 27195 4395 27215 4415
rect 27250 4395 27270 4415
rect 27305 4395 27325 4415
rect 27360 4395 27380 4415
rect 27415 4395 27435 4415
rect 27470 4395 27490 4415
rect 16905 4320 16925 4340
rect 17195 4305 17215 4325
rect 17255 4305 17275 4325
rect 17315 4305 17335 4325
rect 17375 4305 17395 4325
rect 17435 4305 17455 4325
rect 17495 4305 17515 4325
rect 17555 4305 17575 4325
rect 17615 4305 17635 4325
rect 17675 4305 17695 4325
rect 16260 4070 16280 4090
rect 16315 4070 16335 4090
rect 16370 4070 16390 4090
rect 16425 4070 16445 4090
rect 16480 4070 16500 4090
rect 16535 4070 16555 4090
rect 16590 4070 16610 4090
rect 16645 4070 16665 4090
rect 16700 4070 16720 4090
rect 16755 4070 16775 4090
rect 16810 4070 16830 4090
rect 16865 4070 16885 4090
rect 16920 4070 16940 4090
rect 16975 4070 16995 4090
rect 17030 4070 17050 4090
rect 17085 4070 17105 4090
rect 17140 4070 17160 4090
rect 17195 4070 17215 4090
rect 17250 4070 17270 4090
rect 17305 4070 17325 4090
rect 17360 4070 17380 4090
rect 17415 4070 17435 4090
rect 17470 4070 17490 4090
rect 26210 3985 26230 4005
rect 26265 3985 26285 4005
rect 26320 3985 26340 4005
rect 26375 3985 26395 4005
rect 26430 3985 26450 4005
rect 26485 3985 26505 4005
rect 26540 3985 26560 4005
rect 26595 3985 26615 4005
rect 26650 3985 26670 4005
rect 26705 3985 26725 4005
rect 26760 3985 26780 4005
rect 26815 3985 26835 4005
rect 26870 3985 26890 4005
rect 26940 3985 26960 4005
rect 26995 3985 27015 4005
rect 27050 3985 27070 4005
rect 27105 3985 27125 4005
rect 27160 3985 27180 4005
rect 27215 3985 27235 4005
rect 27270 3985 27290 4005
rect 27325 3985 27345 4005
rect 27380 3985 27400 4005
rect 27435 3985 27455 4005
rect 27490 3985 27510 4005
rect 27545 3985 27565 4005
rect 27600 3985 27620 4005
rect 16205 3765 16225 3785
rect 16260 3765 16280 3785
rect 16315 3765 16335 3785
rect 16370 3765 16390 3785
rect 16425 3765 16445 3785
rect 16480 3765 16500 3785
rect 16535 3765 16555 3785
rect 16590 3765 16610 3785
rect 16645 3765 16665 3785
rect 16700 3765 16720 3785
rect 16755 3765 16775 3785
rect 16810 3765 16830 3785
rect 16865 3765 16885 3785
rect 16945 3765 16965 3785
rect 17000 3765 17020 3785
rect 17055 3765 17075 3785
rect 17110 3765 17130 3785
rect 17165 3765 17185 3785
rect 17220 3765 17240 3785
rect 17275 3765 17295 3785
rect 17330 3765 17350 3785
rect 17385 3765 17405 3785
rect 17440 3765 17460 3785
rect 17495 3765 17515 3785
rect 17550 3765 17570 3785
rect 17605 3765 17625 3785
rect 15015 3550 15035 3570
rect 15015 3500 15035 3520
rect 15015 3450 15035 3470
rect 15015 3400 15035 3420
rect 15015 3350 15035 3370
rect 15015 3300 15035 3320
rect 15015 3250 15035 3270
rect 15015 3200 15035 3220
rect 15015 3150 15035 3170
rect 15015 3100 15035 3120
rect 15015 3050 15035 3070
rect 15015 3000 15035 3020
rect 15070 3550 15090 3570
rect 15070 3500 15090 3520
rect 15070 3450 15090 3470
rect 15070 3400 15090 3420
rect 15070 3350 15090 3370
rect 15070 3300 15090 3320
rect 15070 3250 15090 3270
rect 15070 3200 15090 3220
rect 15070 3150 15090 3170
rect 15070 3100 15090 3120
rect 15070 3050 15090 3070
rect 15070 3000 15090 3020
rect 15125 3550 15145 3570
rect 15125 3500 15145 3520
rect 15125 3450 15145 3470
rect 15125 3400 15145 3420
rect 15125 3350 15145 3370
rect 15125 3300 15145 3320
rect 15125 3250 15145 3270
rect 15125 3200 15145 3220
rect 15125 3150 15145 3170
rect 15125 3100 15145 3120
rect 15125 3050 15145 3070
rect 15125 3000 15145 3020
rect 15180 3550 15200 3570
rect 15180 3500 15200 3520
rect 15180 3450 15200 3470
rect 15180 3400 15200 3420
rect 15180 3350 15200 3370
rect 15180 3300 15200 3320
rect 15180 3250 15200 3270
rect 15180 3200 15200 3220
rect 15180 3150 15200 3170
rect 15180 3100 15200 3120
rect 15180 3050 15200 3070
rect 15180 3000 15200 3020
rect 15235 3550 15255 3570
rect 15235 3500 15255 3520
rect 15235 3450 15255 3470
rect 15235 3400 15255 3420
rect 15235 3350 15255 3370
rect 15235 3300 15255 3320
rect 15235 3250 15255 3270
rect 15235 3200 15255 3220
rect 15235 3150 15255 3170
rect 15235 3100 15255 3120
rect 15235 3050 15255 3070
rect 15235 3000 15255 3020
rect 15290 3550 15310 3570
rect 15290 3500 15310 3520
rect 15290 3450 15310 3470
rect 15290 3400 15310 3420
rect 15290 3350 15310 3370
rect 15290 3300 15310 3320
rect 15290 3250 15310 3270
rect 15290 3200 15310 3220
rect 15290 3150 15310 3170
rect 15290 3100 15310 3120
rect 15290 3050 15310 3070
rect 15290 3000 15310 3020
rect 15345 3550 15365 3570
rect 15345 3500 15365 3520
rect 15345 3450 15365 3470
rect 15345 3400 15365 3420
rect 15345 3350 15365 3370
rect 15345 3300 15365 3320
rect 15345 3250 15365 3270
rect 15345 3200 15365 3220
rect 15345 3150 15365 3170
rect 15345 3100 15365 3120
rect 15345 3050 15365 3070
rect 15345 3000 15365 3020
rect 15400 3550 15420 3570
rect 15400 3500 15420 3520
rect 15400 3450 15420 3470
rect 15400 3400 15420 3420
rect 15400 3350 15420 3370
rect 15400 3300 15420 3320
rect 15400 3250 15420 3270
rect 15400 3200 15420 3220
rect 15400 3150 15420 3170
rect 15400 3100 15420 3120
rect 15400 3050 15420 3070
rect 15400 3000 15420 3020
rect 15455 3550 15475 3570
rect 15455 3500 15475 3520
rect 15455 3450 15475 3470
rect 15455 3400 15475 3420
rect 15455 3350 15475 3370
rect 15455 3300 15475 3320
rect 15455 3250 15475 3270
rect 15455 3200 15475 3220
rect 15455 3150 15475 3170
rect 15455 3100 15475 3120
rect 15455 3050 15475 3070
rect 15455 3000 15475 3020
rect 15510 3550 15530 3570
rect 15510 3500 15530 3520
rect 15510 3450 15530 3470
rect 15510 3400 15530 3420
rect 15510 3350 15530 3370
rect 15510 3300 15530 3320
rect 15510 3250 15530 3270
rect 15510 3200 15530 3220
rect 15510 3150 15530 3170
rect 15510 3100 15530 3120
rect 15510 3050 15530 3070
rect 15510 3000 15530 3020
rect 15565 3550 15585 3570
rect 15565 3500 15585 3520
rect 15565 3450 15585 3470
rect 15565 3400 15585 3420
rect 15565 3350 15585 3370
rect 15565 3300 15585 3320
rect 15565 3250 15585 3270
rect 15565 3200 15585 3220
rect 15565 3150 15585 3170
rect 15565 3100 15585 3120
rect 15565 3050 15585 3070
rect 15565 3000 15585 3020
rect 15620 3550 15640 3570
rect 15620 3500 15640 3520
rect 15620 3450 15640 3470
rect 15620 3400 15640 3420
rect 15620 3350 15640 3370
rect 15620 3300 15640 3320
rect 15620 3250 15640 3270
rect 15620 3200 15640 3220
rect 15620 3150 15640 3170
rect 15620 3100 15640 3120
rect 15620 3050 15640 3070
rect 15620 3000 15640 3020
rect 15675 3550 15695 3570
rect 18155 3550 18175 3570
rect 15675 3500 15695 3520
rect 15675 3450 15695 3470
rect 15675 3400 15695 3420
rect 15675 3350 15695 3370
rect 15675 3300 15695 3320
rect 15675 3250 15695 3270
rect 15675 3200 15695 3220
rect 15675 3150 15695 3170
rect 16230 3490 16250 3510
rect 16230 3440 16250 3460
rect 16230 3390 16250 3410
rect 16230 3340 16250 3360
rect 16230 3290 16250 3310
rect 16230 3240 16250 3260
rect 16230 3190 16250 3210
rect 16230 3140 16250 3160
rect 16290 3490 16310 3510
rect 16290 3440 16310 3460
rect 16290 3390 16310 3410
rect 16290 3340 16310 3360
rect 16290 3290 16310 3310
rect 16290 3240 16310 3260
rect 16290 3190 16310 3210
rect 16290 3140 16310 3160
rect 16350 3490 16370 3510
rect 16350 3440 16370 3460
rect 16350 3390 16370 3410
rect 16350 3340 16370 3360
rect 16350 3290 16370 3310
rect 16350 3240 16370 3260
rect 16350 3190 16370 3210
rect 16350 3140 16370 3160
rect 16410 3490 16430 3510
rect 16410 3440 16430 3460
rect 16410 3390 16430 3410
rect 16410 3340 16430 3360
rect 16410 3290 16430 3310
rect 16410 3240 16430 3260
rect 16410 3190 16430 3210
rect 16410 3140 16430 3160
rect 16470 3490 16490 3510
rect 16470 3440 16490 3460
rect 16470 3390 16490 3410
rect 16470 3340 16490 3360
rect 16470 3290 16490 3310
rect 16470 3240 16490 3260
rect 16470 3190 16490 3210
rect 16470 3140 16490 3160
rect 16530 3490 16550 3510
rect 16530 3440 16550 3460
rect 16530 3390 16550 3410
rect 16530 3340 16550 3360
rect 16530 3290 16550 3310
rect 16530 3240 16550 3260
rect 16530 3190 16550 3210
rect 16530 3140 16550 3160
rect 16590 3490 16610 3510
rect 16590 3440 16610 3460
rect 16590 3390 16610 3410
rect 16590 3340 16610 3360
rect 16590 3290 16610 3310
rect 16590 3240 16610 3260
rect 16590 3190 16610 3210
rect 16590 3140 16610 3160
rect 16650 3490 16670 3510
rect 16650 3440 16670 3460
rect 16650 3390 16670 3410
rect 16650 3340 16670 3360
rect 16650 3290 16670 3310
rect 16650 3240 16670 3260
rect 16650 3190 16670 3210
rect 16650 3140 16670 3160
rect 16710 3490 16730 3510
rect 16710 3440 16730 3460
rect 16710 3390 16730 3410
rect 16710 3340 16730 3360
rect 16710 3290 16730 3310
rect 16710 3240 16730 3260
rect 16710 3190 16730 3210
rect 16710 3140 16730 3160
rect 16770 3490 16790 3510
rect 16770 3440 16790 3460
rect 16770 3390 16790 3410
rect 16770 3340 16790 3360
rect 16770 3290 16790 3310
rect 16770 3240 16790 3260
rect 16770 3190 16790 3210
rect 16770 3140 16790 3160
rect 16830 3490 16850 3510
rect 16830 3440 16850 3460
rect 16830 3390 16850 3410
rect 16830 3340 16850 3360
rect 16830 3290 16850 3310
rect 16830 3240 16850 3260
rect 16830 3190 16850 3210
rect 16830 3140 16850 3160
rect 16890 3490 16910 3510
rect 16890 3440 16910 3460
rect 16890 3390 16910 3410
rect 16890 3340 16910 3360
rect 16890 3290 16910 3310
rect 16890 3240 16910 3260
rect 16890 3190 16910 3210
rect 16890 3140 16910 3160
rect 16950 3490 16970 3510
rect 16950 3440 16970 3460
rect 16950 3390 16970 3410
rect 16950 3340 16970 3360
rect 16950 3290 16970 3310
rect 16950 3240 16970 3260
rect 16950 3190 16970 3210
rect 16950 3140 16970 3160
rect 17010 3490 17030 3510
rect 17010 3440 17030 3460
rect 17010 3390 17030 3410
rect 17010 3340 17030 3360
rect 17010 3290 17030 3310
rect 17010 3240 17030 3260
rect 17010 3190 17030 3210
rect 17010 3140 17030 3160
rect 17070 3490 17090 3510
rect 17070 3440 17090 3460
rect 17070 3390 17090 3410
rect 17070 3340 17090 3360
rect 17070 3290 17090 3310
rect 17070 3240 17090 3260
rect 17070 3190 17090 3210
rect 17070 3140 17090 3160
rect 17130 3490 17150 3510
rect 17130 3440 17150 3460
rect 17130 3390 17150 3410
rect 17130 3340 17150 3360
rect 17130 3290 17150 3310
rect 17130 3240 17150 3260
rect 17130 3190 17150 3210
rect 17130 3140 17150 3160
rect 17190 3490 17210 3510
rect 17190 3440 17210 3460
rect 17190 3390 17210 3410
rect 17190 3340 17210 3360
rect 17190 3290 17210 3310
rect 17190 3240 17210 3260
rect 17190 3190 17210 3210
rect 17190 3140 17210 3160
rect 17250 3490 17270 3510
rect 17250 3440 17270 3460
rect 17250 3390 17270 3410
rect 17250 3340 17270 3360
rect 17250 3290 17270 3310
rect 17250 3240 17270 3260
rect 17250 3190 17270 3210
rect 17250 3140 17270 3160
rect 17310 3490 17330 3510
rect 17310 3440 17330 3460
rect 17310 3390 17330 3410
rect 17310 3340 17330 3360
rect 17310 3290 17330 3310
rect 17310 3240 17330 3260
rect 17310 3190 17330 3210
rect 17310 3140 17330 3160
rect 17370 3490 17390 3510
rect 17370 3440 17390 3460
rect 17370 3390 17390 3410
rect 17370 3340 17390 3360
rect 17370 3290 17390 3310
rect 17370 3240 17390 3260
rect 17370 3190 17390 3210
rect 17370 3140 17390 3160
rect 17430 3490 17450 3510
rect 17430 3440 17450 3460
rect 17430 3390 17450 3410
rect 17430 3340 17450 3360
rect 17430 3290 17450 3310
rect 17430 3240 17450 3260
rect 17430 3190 17450 3210
rect 17430 3140 17450 3160
rect 17490 3490 17510 3510
rect 17490 3440 17510 3460
rect 17490 3390 17510 3410
rect 17490 3340 17510 3360
rect 17490 3290 17510 3310
rect 17490 3240 17510 3260
rect 17490 3190 17510 3210
rect 17490 3140 17510 3160
rect 17550 3490 17570 3510
rect 17550 3440 17570 3460
rect 17550 3390 17570 3410
rect 17550 3340 17570 3360
rect 17550 3290 17570 3310
rect 17550 3240 17570 3260
rect 17550 3190 17570 3210
rect 17550 3140 17570 3160
rect 18155 3500 18175 3520
rect 18155 3450 18175 3470
rect 18155 3400 18175 3420
rect 18155 3350 18175 3370
rect 18155 3300 18175 3320
rect 18155 3250 18175 3270
rect 18155 3200 18175 3220
rect 18155 3150 18175 3170
rect 15675 3100 15695 3120
rect 18155 3100 18175 3120
rect 15675 3050 15695 3070
rect 15675 3000 15695 3020
rect 18155 3050 18175 3070
rect 18155 3000 18175 3020
rect 18210 3550 18230 3570
rect 18210 3500 18230 3520
rect 18210 3450 18230 3470
rect 18210 3400 18230 3420
rect 18210 3350 18230 3370
rect 18210 3300 18230 3320
rect 18210 3250 18230 3270
rect 18210 3200 18230 3220
rect 18210 3150 18230 3170
rect 18210 3100 18230 3120
rect 18210 3050 18230 3070
rect 18210 3000 18230 3020
rect 18265 3550 18285 3570
rect 18265 3500 18285 3520
rect 18265 3450 18285 3470
rect 18265 3400 18285 3420
rect 18265 3350 18285 3370
rect 18265 3300 18285 3320
rect 18265 3250 18285 3270
rect 18265 3200 18285 3220
rect 18265 3150 18285 3170
rect 18265 3100 18285 3120
rect 18265 3050 18285 3070
rect 18265 3000 18285 3020
rect 18320 3550 18340 3570
rect 18320 3500 18340 3520
rect 18320 3450 18340 3470
rect 18320 3400 18340 3420
rect 18320 3350 18340 3370
rect 18320 3300 18340 3320
rect 18320 3250 18340 3270
rect 18320 3200 18340 3220
rect 18320 3150 18340 3170
rect 18320 3100 18340 3120
rect 18320 3050 18340 3070
rect 18320 3000 18340 3020
rect 18375 3550 18395 3570
rect 18375 3500 18395 3520
rect 18375 3450 18395 3470
rect 18375 3400 18395 3420
rect 18375 3350 18395 3370
rect 18375 3300 18395 3320
rect 18375 3250 18395 3270
rect 18375 3200 18395 3220
rect 18375 3150 18395 3170
rect 18375 3100 18395 3120
rect 18375 3050 18395 3070
rect 18375 3000 18395 3020
rect 18430 3550 18450 3570
rect 18430 3500 18450 3520
rect 18430 3450 18450 3470
rect 18430 3400 18450 3420
rect 18430 3350 18450 3370
rect 18430 3300 18450 3320
rect 18430 3250 18450 3270
rect 18430 3200 18450 3220
rect 18430 3150 18450 3170
rect 18430 3100 18450 3120
rect 18430 3050 18450 3070
rect 18430 3000 18450 3020
rect 18485 3550 18505 3570
rect 18485 3500 18505 3520
rect 18485 3450 18505 3470
rect 18485 3400 18505 3420
rect 18485 3350 18505 3370
rect 18485 3300 18505 3320
rect 18485 3250 18505 3270
rect 18485 3200 18505 3220
rect 18485 3150 18505 3170
rect 18485 3100 18505 3120
rect 18485 3050 18505 3070
rect 18485 3000 18505 3020
rect 18540 3550 18560 3570
rect 18540 3500 18560 3520
rect 18540 3450 18560 3470
rect 18540 3400 18560 3420
rect 18540 3350 18560 3370
rect 18540 3300 18560 3320
rect 18540 3250 18560 3270
rect 18540 3200 18560 3220
rect 18540 3150 18560 3170
rect 18540 3100 18560 3120
rect 18540 3050 18560 3070
rect 18540 3000 18560 3020
rect 18595 3550 18615 3570
rect 18595 3500 18615 3520
rect 18595 3450 18615 3470
rect 18595 3400 18615 3420
rect 18595 3350 18615 3370
rect 18595 3300 18615 3320
rect 18595 3250 18615 3270
rect 18595 3200 18615 3220
rect 18595 3150 18615 3170
rect 18595 3100 18615 3120
rect 18595 3050 18615 3070
rect 18595 3000 18615 3020
rect 18650 3550 18670 3570
rect 18650 3500 18670 3520
rect 18650 3450 18670 3470
rect 18650 3400 18670 3420
rect 18650 3350 18670 3370
rect 18650 3300 18670 3320
rect 18650 3250 18670 3270
rect 18650 3200 18670 3220
rect 18650 3150 18670 3170
rect 18650 3100 18670 3120
rect 18650 3050 18670 3070
rect 18650 3000 18670 3020
rect 18705 3550 18725 3570
rect 18705 3500 18725 3520
rect 18705 3450 18725 3470
rect 18705 3400 18725 3420
rect 18705 3350 18725 3370
rect 18705 3300 18725 3320
rect 18705 3250 18725 3270
rect 18705 3200 18725 3220
rect 18705 3150 18725 3170
rect 18705 3100 18725 3120
rect 18705 3050 18725 3070
rect 18705 3000 18725 3020
rect 18760 3550 18780 3570
rect 18760 3500 18780 3520
rect 18760 3450 18780 3470
rect 18760 3400 18780 3420
rect 18760 3350 18780 3370
rect 18760 3300 18780 3320
rect 18760 3250 18780 3270
rect 18760 3200 18780 3220
rect 18760 3150 18780 3170
rect 18760 3100 18780 3120
rect 18760 3050 18780 3070
rect 18760 3000 18780 3020
rect 18815 3550 18835 3570
rect 25015 3550 25035 3570
rect 18815 3500 18835 3520
rect 18815 3450 18835 3470
rect 18815 3400 18835 3420
rect 18815 3350 18835 3370
rect 18815 3300 18835 3320
rect 18815 3250 18835 3270
rect 18815 3200 18835 3220
rect 18815 3150 18835 3170
rect 18815 3100 18835 3120
rect 18815 3050 18835 3070
rect 18815 3000 18835 3020
rect 25015 3500 25035 3520
rect 25015 3450 25035 3470
rect 25015 3400 25035 3420
rect 25015 3350 25035 3370
rect 25015 3300 25035 3320
rect 25015 3250 25035 3270
rect 25015 3200 25035 3220
rect 25015 3150 25035 3170
rect 25015 3100 25035 3120
rect 25015 3050 25035 3070
rect 25015 3000 25035 3020
rect 25070 3550 25090 3570
rect 25070 3500 25090 3520
rect 25070 3450 25090 3470
rect 25070 3400 25090 3420
rect 25070 3350 25090 3370
rect 25070 3300 25090 3320
rect 25070 3250 25090 3270
rect 25070 3200 25090 3220
rect 25070 3150 25090 3170
rect 25070 3100 25090 3120
rect 25070 3050 25090 3070
rect 25070 3000 25090 3020
rect 25125 3550 25145 3570
rect 25125 3500 25145 3520
rect 25125 3450 25145 3470
rect 25125 3400 25145 3420
rect 25125 3350 25145 3370
rect 25125 3300 25145 3320
rect 25125 3250 25145 3270
rect 25125 3200 25145 3220
rect 25125 3150 25145 3170
rect 25125 3100 25145 3120
rect 25125 3050 25145 3070
rect 25125 3000 25145 3020
rect 25180 3550 25200 3570
rect 25180 3500 25200 3520
rect 25180 3450 25200 3470
rect 25180 3400 25200 3420
rect 25180 3350 25200 3370
rect 25180 3300 25200 3320
rect 25180 3250 25200 3270
rect 25180 3200 25200 3220
rect 25180 3150 25200 3170
rect 25180 3100 25200 3120
rect 25180 3050 25200 3070
rect 25180 3000 25200 3020
rect 25235 3550 25255 3570
rect 25235 3500 25255 3520
rect 25235 3450 25255 3470
rect 25235 3400 25255 3420
rect 25235 3350 25255 3370
rect 25235 3300 25255 3320
rect 25235 3250 25255 3270
rect 25235 3200 25255 3220
rect 25235 3150 25255 3170
rect 25235 3100 25255 3120
rect 25235 3050 25255 3070
rect 25235 3000 25255 3020
rect 25290 3550 25310 3570
rect 25290 3500 25310 3520
rect 25290 3450 25310 3470
rect 25290 3400 25310 3420
rect 25290 3350 25310 3370
rect 25290 3300 25310 3320
rect 25290 3250 25310 3270
rect 25290 3200 25310 3220
rect 25290 3150 25310 3170
rect 25290 3100 25310 3120
rect 25290 3050 25310 3070
rect 25290 3000 25310 3020
rect 25345 3550 25365 3570
rect 25345 3500 25365 3520
rect 25345 3450 25365 3470
rect 25345 3400 25365 3420
rect 25345 3350 25365 3370
rect 25345 3300 25365 3320
rect 25345 3250 25365 3270
rect 25345 3200 25365 3220
rect 25345 3150 25365 3170
rect 25345 3100 25365 3120
rect 25345 3050 25365 3070
rect 25345 3000 25365 3020
rect 25400 3550 25420 3570
rect 25400 3500 25420 3520
rect 25400 3450 25420 3470
rect 25400 3400 25420 3420
rect 25400 3350 25420 3370
rect 25400 3300 25420 3320
rect 25400 3250 25420 3270
rect 25400 3200 25420 3220
rect 25400 3150 25420 3170
rect 25400 3100 25420 3120
rect 25400 3050 25420 3070
rect 25400 3000 25420 3020
rect 25455 3550 25475 3570
rect 25455 3500 25475 3520
rect 25455 3450 25475 3470
rect 25455 3400 25475 3420
rect 25455 3350 25475 3370
rect 25455 3300 25475 3320
rect 25455 3250 25475 3270
rect 25455 3200 25475 3220
rect 25455 3150 25475 3170
rect 25455 3100 25475 3120
rect 25455 3050 25475 3070
rect 25455 3000 25475 3020
rect 25510 3550 25530 3570
rect 25510 3500 25530 3520
rect 25510 3450 25530 3470
rect 25510 3400 25530 3420
rect 25510 3350 25530 3370
rect 25510 3300 25530 3320
rect 25510 3250 25530 3270
rect 25510 3200 25530 3220
rect 25510 3150 25530 3170
rect 25510 3100 25530 3120
rect 25510 3050 25530 3070
rect 25510 3000 25530 3020
rect 25565 3550 25585 3570
rect 25565 3500 25585 3520
rect 25565 3450 25585 3470
rect 25565 3400 25585 3420
rect 25565 3350 25585 3370
rect 25565 3300 25585 3320
rect 25565 3250 25585 3270
rect 25565 3200 25585 3220
rect 25565 3150 25585 3170
rect 25565 3100 25585 3120
rect 25565 3050 25585 3070
rect 25565 3000 25585 3020
rect 25620 3550 25640 3570
rect 25620 3500 25640 3520
rect 25620 3450 25640 3470
rect 25620 3400 25640 3420
rect 25620 3350 25640 3370
rect 25620 3300 25640 3320
rect 25620 3250 25640 3270
rect 25620 3200 25640 3220
rect 25620 3150 25640 3170
rect 25620 3100 25640 3120
rect 25620 3050 25640 3070
rect 25620 3000 25640 3020
rect 25675 3550 25695 3570
rect 25675 3500 25695 3520
rect 25675 3450 25695 3470
rect 25675 3400 25695 3420
rect 25675 3350 25695 3370
rect 25675 3300 25695 3320
rect 25675 3250 25695 3270
rect 25675 3200 25695 3220
rect 25675 3150 25695 3170
rect 25675 3100 25695 3120
rect 26230 3570 26250 3590
rect 26230 3520 26250 3540
rect 26230 3470 26250 3490
rect 26230 3420 26250 3440
rect 26230 3370 26250 3390
rect 26230 3320 26250 3340
rect 26230 3270 26250 3290
rect 26230 3220 26250 3240
rect 26290 3570 26310 3590
rect 26290 3520 26310 3540
rect 26290 3470 26310 3490
rect 26290 3420 26310 3440
rect 26290 3370 26310 3390
rect 26290 3320 26310 3340
rect 26290 3270 26310 3290
rect 26290 3220 26310 3240
rect 26350 3570 26370 3590
rect 26350 3520 26370 3540
rect 26350 3470 26370 3490
rect 26350 3420 26370 3440
rect 26350 3370 26370 3390
rect 26350 3320 26370 3340
rect 26350 3270 26370 3290
rect 26350 3220 26370 3240
rect 26410 3570 26430 3590
rect 26410 3520 26430 3540
rect 26410 3470 26430 3490
rect 26410 3420 26430 3440
rect 26410 3370 26430 3390
rect 26410 3320 26430 3340
rect 26410 3270 26430 3290
rect 26410 3220 26430 3240
rect 26470 3570 26490 3590
rect 26470 3520 26490 3540
rect 26470 3470 26490 3490
rect 26470 3420 26490 3440
rect 26470 3370 26490 3390
rect 26470 3320 26490 3340
rect 26470 3270 26490 3290
rect 26470 3220 26490 3240
rect 26530 3570 26550 3590
rect 26530 3520 26550 3540
rect 26530 3470 26550 3490
rect 26530 3420 26550 3440
rect 26530 3370 26550 3390
rect 26530 3320 26550 3340
rect 26530 3270 26550 3290
rect 26530 3220 26550 3240
rect 26590 3570 26610 3590
rect 26590 3520 26610 3540
rect 26590 3470 26610 3490
rect 26590 3420 26610 3440
rect 26590 3370 26610 3390
rect 26590 3320 26610 3340
rect 26590 3270 26610 3290
rect 26590 3220 26610 3240
rect 26650 3570 26670 3590
rect 26650 3520 26670 3540
rect 26650 3470 26670 3490
rect 26650 3420 26670 3440
rect 26650 3370 26670 3390
rect 26650 3320 26670 3340
rect 26650 3270 26670 3290
rect 26650 3220 26670 3240
rect 26710 3570 26730 3590
rect 26710 3520 26730 3540
rect 26710 3470 26730 3490
rect 26710 3420 26730 3440
rect 26710 3370 26730 3390
rect 26710 3320 26730 3340
rect 26710 3270 26730 3290
rect 26710 3220 26730 3240
rect 26770 3570 26790 3590
rect 26770 3520 26790 3540
rect 26770 3470 26790 3490
rect 26770 3420 26790 3440
rect 26770 3370 26790 3390
rect 26770 3320 26790 3340
rect 26770 3270 26790 3290
rect 26770 3220 26790 3240
rect 26830 3570 26850 3590
rect 26830 3520 26850 3540
rect 26830 3470 26850 3490
rect 26830 3420 26850 3440
rect 26830 3370 26850 3390
rect 26830 3320 26850 3340
rect 26830 3270 26850 3290
rect 26830 3220 26850 3240
rect 26890 3570 26910 3590
rect 26890 3520 26910 3540
rect 26890 3470 26910 3490
rect 26890 3420 26910 3440
rect 26890 3370 26910 3390
rect 26890 3320 26910 3340
rect 26890 3270 26910 3290
rect 26890 3220 26910 3240
rect 26950 3570 26970 3590
rect 26950 3520 26970 3540
rect 26950 3470 26970 3490
rect 26950 3420 26970 3440
rect 26950 3370 26970 3390
rect 26950 3320 26970 3340
rect 26950 3270 26970 3290
rect 26950 3220 26970 3240
rect 27010 3570 27030 3590
rect 27010 3520 27030 3540
rect 27010 3470 27030 3490
rect 27010 3420 27030 3440
rect 27010 3370 27030 3390
rect 27010 3320 27030 3340
rect 27010 3270 27030 3290
rect 27010 3220 27030 3240
rect 27070 3570 27090 3590
rect 27070 3520 27090 3540
rect 27070 3470 27090 3490
rect 27070 3420 27090 3440
rect 27070 3370 27090 3390
rect 27070 3320 27090 3340
rect 27070 3270 27090 3290
rect 27070 3220 27090 3240
rect 27130 3570 27150 3590
rect 27130 3520 27150 3540
rect 27130 3470 27150 3490
rect 27130 3420 27150 3440
rect 27130 3370 27150 3390
rect 27130 3320 27150 3340
rect 27130 3270 27150 3290
rect 27130 3220 27150 3240
rect 27190 3570 27210 3590
rect 27190 3520 27210 3540
rect 27190 3470 27210 3490
rect 27190 3420 27210 3440
rect 27190 3370 27210 3390
rect 27190 3320 27210 3340
rect 27190 3270 27210 3290
rect 27190 3220 27210 3240
rect 27250 3570 27270 3590
rect 27250 3520 27270 3540
rect 27250 3470 27270 3490
rect 27250 3420 27270 3440
rect 27250 3370 27270 3390
rect 27250 3320 27270 3340
rect 27250 3270 27270 3290
rect 27250 3220 27270 3240
rect 27310 3570 27330 3590
rect 27310 3520 27330 3540
rect 27310 3470 27330 3490
rect 27310 3420 27330 3440
rect 27310 3370 27330 3390
rect 27310 3320 27330 3340
rect 27310 3270 27330 3290
rect 27310 3220 27330 3240
rect 27370 3570 27390 3590
rect 27370 3520 27390 3540
rect 27370 3470 27390 3490
rect 27370 3420 27390 3440
rect 27370 3370 27390 3390
rect 27370 3320 27390 3340
rect 27370 3270 27390 3290
rect 27370 3220 27390 3240
rect 27430 3570 27450 3590
rect 27430 3520 27450 3540
rect 27430 3470 27450 3490
rect 27430 3420 27450 3440
rect 27430 3370 27450 3390
rect 27430 3320 27450 3340
rect 27430 3270 27450 3290
rect 27430 3220 27450 3240
rect 27490 3570 27510 3590
rect 27490 3520 27510 3540
rect 27490 3470 27510 3490
rect 27490 3420 27510 3440
rect 27490 3370 27510 3390
rect 27490 3320 27510 3340
rect 27490 3270 27510 3290
rect 27490 3220 27510 3240
rect 27550 3570 27570 3590
rect 27550 3520 27570 3540
rect 27550 3470 27570 3490
rect 27550 3420 27570 3440
rect 27550 3370 27570 3390
rect 27550 3320 27570 3340
rect 27550 3270 27570 3290
rect 27550 3220 27570 3240
rect 25675 3050 25695 3070
rect 25675 3000 25695 3020
rect 28155 3630 28175 3650
rect 28155 3580 28175 3600
rect 28155 3530 28175 3550
rect 28155 3480 28175 3500
rect 28155 3430 28175 3450
rect 28155 3380 28175 3400
rect 28155 3330 28175 3350
rect 28155 3280 28175 3300
rect 28155 3230 28175 3250
rect 28155 3180 28175 3200
rect 28155 3130 28175 3150
rect 28155 3080 28175 3100
rect 28210 3630 28230 3650
rect 28210 3580 28230 3600
rect 28210 3530 28230 3550
rect 28210 3480 28230 3500
rect 28210 3430 28230 3450
rect 28210 3380 28230 3400
rect 28210 3330 28230 3350
rect 28210 3280 28230 3300
rect 28210 3230 28230 3250
rect 28210 3180 28230 3200
rect 28210 3130 28230 3150
rect 28210 3080 28230 3100
rect 28265 3630 28285 3650
rect 28265 3580 28285 3600
rect 28265 3530 28285 3550
rect 28265 3480 28285 3500
rect 28265 3430 28285 3450
rect 28265 3380 28285 3400
rect 28265 3330 28285 3350
rect 28265 3280 28285 3300
rect 28265 3230 28285 3250
rect 28265 3180 28285 3200
rect 28265 3130 28285 3150
rect 28265 3080 28285 3100
rect 28320 3630 28340 3650
rect 28320 3580 28340 3600
rect 28320 3530 28340 3550
rect 28320 3480 28340 3500
rect 28320 3430 28340 3450
rect 28320 3380 28340 3400
rect 28320 3330 28340 3350
rect 28320 3280 28340 3300
rect 28320 3230 28340 3250
rect 28320 3180 28340 3200
rect 28320 3130 28340 3150
rect 28320 3080 28340 3100
rect 28375 3630 28395 3650
rect 28375 3580 28395 3600
rect 28375 3530 28395 3550
rect 28375 3480 28395 3500
rect 28375 3430 28395 3450
rect 28375 3380 28395 3400
rect 28375 3330 28395 3350
rect 28375 3280 28395 3300
rect 28375 3230 28395 3250
rect 28375 3180 28395 3200
rect 28375 3130 28395 3150
rect 28375 3080 28395 3100
rect 28430 3630 28450 3650
rect 28430 3580 28450 3600
rect 28430 3530 28450 3550
rect 28430 3480 28450 3500
rect 28430 3430 28450 3450
rect 28430 3380 28450 3400
rect 28430 3330 28450 3350
rect 28430 3280 28450 3300
rect 28430 3230 28450 3250
rect 28430 3180 28450 3200
rect 28430 3130 28450 3150
rect 28430 3080 28450 3100
rect 28485 3630 28505 3650
rect 28485 3580 28505 3600
rect 28485 3530 28505 3550
rect 28485 3480 28505 3500
rect 28485 3430 28505 3450
rect 28485 3380 28505 3400
rect 28485 3330 28505 3350
rect 28485 3280 28505 3300
rect 28485 3230 28505 3250
rect 28485 3180 28505 3200
rect 28485 3130 28505 3150
rect 28485 3080 28505 3100
rect 28540 3630 28560 3650
rect 28540 3580 28560 3600
rect 28540 3530 28560 3550
rect 28540 3480 28560 3500
rect 28540 3430 28560 3450
rect 28540 3380 28560 3400
rect 28540 3330 28560 3350
rect 28540 3280 28560 3300
rect 28540 3230 28560 3250
rect 28540 3180 28560 3200
rect 28540 3130 28560 3150
rect 28540 3080 28560 3100
rect 28595 3630 28615 3650
rect 28595 3580 28615 3600
rect 28595 3530 28615 3550
rect 28595 3480 28615 3500
rect 28595 3430 28615 3450
rect 28595 3380 28615 3400
rect 28595 3330 28615 3350
rect 28595 3280 28615 3300
rect 28595 3230 28615 3250
rect 28595 3180 28615 3200
rect 28595 3130 28615 3150
rect 28595 3080 28615 3100
rect 28650 3630 28670 3650
rect 28650 3580 28670 3600
rect 28650 3530 28670 3550
rect 28650 3480 28670 3500
rect 28650 3430 28670 3450
rect 28650 3380 28670 3400
rect 28650 3330 28670 3350
rect 28650 3280 28670 3300
rect 28650 3230 28670 3250
rect 28650 3180 28670 3200
rect 28650 3130 28670 3150
rect 28650 3080 28670 3100
rect 28705 3630 28725 3650
rect 28705 3580 28725 3600
rect 28705 3530 28725 3550
rect 28705 3480 28725 3500
rect 28705 3430 28725 3450
rect 28705 3380 28725 3400
rect 28705 3330 28725 3350
rect 28705 3280 28725 3300
rect 28705 3230 28725 3250
rect 28705 3180 28725 3200
rect 28705 3130 28725 3150
rect 28705 3080 28725 3100
rect 28760 3630 28780 3650
rect 28760 3580 28780 3600
rect 28760 3530 28780 3550
rect 28760 3480 28780 3500
rect 28760 3430 28780 3450
rect 28760 3380 28780 3400
rect 28760 3330 28780 3350
rect 28760 3280 28780 3300
rect 28760 3230 28780 3250
rect 28760 3180 28780 3200
rect 28760 3130 28780 3150
rect 28760 3080 28780 3100
rect 28815 3630 28835 3650
rect 28815 3580 28835 3600
rect 28815 3530 28835 3550
rect 28815 3480 28835 3500
rect 28815 3430 28835 3450
rect 28815 3380 28835 3400
rect 28815 3330 28835 3350
rect 28815 3280 28835 3300
rect 28815 3230 28835 3250
rect 28815 3180 28835 3200
rect 28815 3130 28835 3150
rect 28815 3080 28835 3100
rect 3005 2895 3025 2915
rect 3005 2845 3025 2865
rect 3095 2895 3115 2915
rect 3095 2845 3115 2865
rect 3185 2895 3205 2915
rect 3185 2845 3205 2865
rect 3275 2895 3295 2915
rect 3275 2845 3295 2865
rect 3365 2895 3385 2915
rect 3365 2845 3385 2865
rect 3455 2895 3475 2915
rect 3455 2845 3475 2865
rect 3545 2895 3565 2915
rect 3545 2845 3565 2865
rect 3635 2895 3655 2915
rect 3635 2845 3655 2865
rect 3725 2895 3745 2915
rect 3725 2845 3745 2865
rect 3815 2895 3835 2915
rect 3815 2845 3835 2865
rect 3905 2895 3925 2915
rect 3905 2845 3925 2865
rect 3995 2895 4015 2915
rect 3995 2845 4015 2865
rect 4085 2895 4105 2915
rect 4085 2845 4105 2865
rect 4175 2895 4195 2915
rect 4175 2845 4195 2865
rect 4265 2895 4285 2915
rect 4265 2845 4285 2865
rect 4355 2895 4375 2915
rect 4355 2845 4375 2865
rect 4445 2895 4465 2915
rect 4445 2845 4465 2865
rect 4535 2895 4555 2915
rect 4535 2845 4555 2865
rect 4625 2895 4645 2915
rect 4625 2845 4645 2865
rect 4715 2895 4735 2915
rect 4715 2845 4735 2865
rect 4805 2895 4825 2915
rect 4805 2845 4825 2865
rect 4895 2895 4915 2915
rect 4895 2845 4915 2865
rect 4985 2895 5005 2915
rect 4985 2845 5005 2865
rect 16025 2810 16045 2830
rect 16025 2760 16045 2780
rect 16025 2710 16045 2730
rect 3185 2665 3205 2685
rect 3185 2615 3205 2635
rect 3185 2565 3205 2585
rect 3185 2515 3205 2535
rect 3185 2465 3205 2485
rect 3185 2415 3205 2435
rect 3275 2665 3295 2685
rect 3275 2615 3295 2635
rect 3275 2565 3295 2585
rect 3275 2515 3295 2535
rect 3275 2465 3295 2485
rect 3275 2415 3295 2435
rect 3365 2665 3385 2685
rect 3365 2615 3385 2635
rect 3365 2565 3385 2585
rect 3365 2515 3385 2535
rect 3365 2465 3385 2485
rect 3365 2415 3385 2435
rect 3455 2665 3475 2685
rect 3455 2615 3475 2635
rect 3455 2565 3475 2585
rect 3455 2515 3475 2535
rect 3455 2465 3475 2485
rect 3455 2415 3475 2435
rect 3545 2665 3565 2685
rect 3545 2615 3565 2635
rect 3545 2565 3565 2585
rect 3545 2515 3565 2535
rect 3545 2465 3565 2485
rect 3545 2415 3565 2435
rect 3635 2665 3655 2685
rect 3635 2615 3655 2635
rect 3635 2565 3655 2585
rect 3635 2515 3655 2535
rect 3635 2465 3655 2485
rect 3635 2415 3655 2435
rect 3725 2665 3745 2685
rect 3725 2615 3745 2635
rect 3725 2565 3745 2585
rect 3725 2515 3745 2535
rect 3725 2465 3745 2485
rect 3725 2415 3745 2435
rect 3815 2665 3835 2685
rect 3815 2615 3835 2635
rect 3815 2565 3835 2585
rect 3815 2515 3835 2535
rect 3815 2465 3835 2485
rect 3815 2415 3835 2435
rect 3905 2665 3925 2685
rect 3905 2615 3925 2635
rect 3905 2565 3925 2585
rect 3905 2515 3925 2535
rect 3905 2465 3925 2485
rect 3905 2415 3925 2435
rect 3995 2665 4015 2685
rect 3995 2615 4015 2635
rect 3995 2565 4015 2585
rect 3995 2515 4015 2535
rect 3995 2465 4015 2485
rect 3995 2415 4015 2435
rect 4085 2665 4105 2685
rect 4085 2615 4105 2635
rect 4085 2565 4105 2585
rect 4085 2515 4105 2535
rect 4085 2465 4105 2485
rect 4085 2415 4105 2435
rect 4175 2665 4195 2685
rect 4175 2615 4195 2635
rect 4175 2565 4195 2585
rect 4175 2515 4195 2535
rect 4175 2465 4195 2485
rect 4175 2415 4195 2435
rect 4265 2665 4285 2685
rect 4265 2615 4285 2635
rect 4265 2565 4285 2585
rect 4265 2515 4285 2535
rect 4265 2465 4285 2485
rect 4265 2415 4285 2435
rect 4355 2665 4375 2685
rect 4355 2615 4375 2635
rect 4355 2565 4375 2585
rect 4355 2515 4375 2535
rect 4355 2465 4375 2485
rect 4355 2415 4375 2435
rect 4445 2665 4465 2685
rect 4445 2615 4465 2635
rect 4445 2565 4465 2585
rect 4445 2515 4465 2535
rect 4445 2465 4465 2485
rect 4445 2415 4465 2435
rect 4535 2665 4555 2685
rect 4535 2615 4555 2635
rect 4535 2565 4555 2585
rect 4535 2515 4555 2535
rect 4535 2465 4555 2485
rect 4535 2415 4555 2435
rect 4625 2665 4645 2685
rect 4625 2615 4645 2635
rect 4625 2565 4645 2585
rect 4625 2515 4645 2535
rect 4625 2465 4645 2485
rect 4625 2415 4645 2435
rect 4715 2665 4735 2685
rect 4715 2615 4735 2635
rect 4715 2565 4735 2585
rect 4715 2515 4735 2535
rect 4715 2465 4735 2485
rect 4715 2415 4735 2435
rect 4805 2665 4825 2685
rect 16025 2660 16045 2680
rect 4805 2615 4825 2635
rect 4805 2565 4825 2585
rect 4805 2515 4825 2535
rect 4805 2465 4825 2485
rect 4805 2415 4825 2435
rect 15015 2620 15035 2640
rect 15015 2570 15035 2590
rect 15015 2520 15035 2540
rect 15015 2470 15035 2490
rect 15070 2620 15090 2640
rect 15070 2570 15090 2590
rect 15070 2520 15090 2540
rect 15070 2470 15090 2490
rect 15125 2620 15145 2640
rect 15125 2570 15145 2590
rect 15125 2520 15145 2540
rect 15125 2470 15145 2490
rect 15180 2620 15200 2640
rect 15180 2570 15200 2590
rect 15180 2520 15200 2540
rect 15180 2470 15200 2490
rect 15235 2620 15255 2640
rect 15235 2570 15255 2590
rect 15235 2520 15255 2540
rect 15235 2470 15255 2490
rect 15290 2620 15310 2640
rect 15290 2570 15310 2590
rect 15290 2520 15310 2540
rect 15290 2470 15310 2490
rect 15345 2620 15365 2640
rect 15345 2570 15365 2590
rect 15345 2520 15365 2540
rect 15345 2470 15365 2490
rect 15400 2620 15420 2640
rect 15400 2570 15420 2590
rect 15400 2520 15420 2540
rect 15400 2470 15420 2490
rect 15455 2620 15475 2640
rect 15455 2570 15475 2590
rect 15455 2520 15475 2540
rect 15455 2470 15475 2490
rect 15510 2620 15530 2640
rect 15510 2570 15530 2590
rect 15510 2520 15530 2540
rect 15510 2470 15530 2490
rect 15565 2620 15585 2640
rect 15565 2570 15585 2590
rect 15565 2520 15585 2540
rect 15565 2470 15585 2490
rect 15620 2620 15640 2640
rect 15620 2570 15640 2590
rect 15620 2520 15640 2540
rect 15620 2470 15640 2490
rect 15675 2620 15695 2640
rect 15675 2570 15695 2590
rect 15675 2520 15695 2540
rect 16025 2610 16045 2630
rect 16025 2560 16045 2580
rect 16025 2510 16045 2530
rect 16085 2810 16105 2830
rect 16085 2760 16105 2780
rect 16085 2710 16105 2730
rect 16085 2660 16105 2680
rect 16085 2610 16105 2630
rect 16085 2560 16105 2580
rect 16085 2510 16105 2530
rect 16145 2810 16165 2830
rect 16145 2760 16165 2780
rect 16145 2710 16165 2730
rect 16145 2660 16165 2680
rect 16145 2610 16165 2630
rect 16145 2560 16165 2580
rect 16145 2510 16165 2530
rect 16205 2810 16225 2830
rect 16205 2760 16225 2780
rect 16205 2710 16225 2730
rect 16205 2660 16225 2680
rect 16205 2610 16225 2630
rect 16205 2560 16225 2580
rect 16205 2510 16225 2530
rect 16265 2810 16285 2830
rect 16265 2760 16285 2780
rect 16265 2710 16285 2730
rect 16265 2660 16285 2680
rect 16265 2610 16285 2630
rect 16265 2560 16285 2580
rect 16265 2510 16285 2530
rect 16325 2810 16345 2830
rect 16325 2760 16345 2780
rect 16325 2710 16345 2730
rect 16325 2660 16345 2680
rect 16325 2610 16345 2630
rect 16325 2560 16345 2580
rect 16325 2510 16345 2530
rect 16385 2810 16405 2830
rect 16385 2760 16405 2780
rect 16385 2710 16405 2730
rect 16385 2660 16405 2680
rect 16385 2610 16405 2630
rect 16385 2560 16405 2580
rect 16385 2510 16405 2530
rect 16445 2810 16465 2830
rect 16445 2760 16465 2780
rect 16445 2710 16465 2730
rect 16445 2660 16465 2680
rect 16445 2610 16465 2630
rect 16445 2560 16465 2580
rect 16445 2510 16465 2530
rect 16505 2810 16525 2830
rect 16505 2760 16525 2780
rect 16505 2710 16525 2730
rect 16505 2660 16525 2680
rect 16505 2610 16525 2630
rect 16505 2560 16525 2580
rect 16505 2510 16525 2530
rect 16565 2810 16585 2830
rect 16565 2760 16585 2780
rect 16565 2710 16585 2730
rect 16565 2660 16585 2680
rect 16565 2610 16585 2630
rect 16565 2560 16585 2580
rect 16565 2510 16585 2530
rect 16625 2810 16645 2830
rect 16625 2760 16645 2780
rect 16625 2710 16645 2730
rect 16625 2660 16645 2680
rect 16625 2610 16645 2630
rect 16625 2560 16645 2580
rect 16625 2510 16645 2530
rect 16685 2810 16705 2830
rect 16685 2760 16705 2780
rect 16685 2710 16705 2730
rect 16685 2660 16705 2680
rect 16685 2610 16705 2630
rect 16685 2560 16705 2580
rect 16685 2510 16705 2530
rect 16745 2810 16765 2830
rect 16745 2760 16765 2780
rect 16745 2710 16765 2730
rect 16745 2660 16765 2680
rect 16745 2610 16765 2630
rect 16745 2560 16765 2580
rect 16745 2510 16765 2530
rect 17035 2810 17055 2830
rect 17035 2760 17055 2780
rect 17035 2710 17055 2730
rect 17035 2660 17055 2680
rect 17035 2610 17055 2630
rect 17035 2560 17055 2580
rect 17035 2510 17055 2530
rect 17095 2810 17115 2830
rect 17095 2760 17115 2780
rect 17095 2710 17115 2730
rect 17095 2660 17115 2680
rect 17095 2610 17115 2630
rect 17095 2560 17115 2580
rect 17095 2510 17115 2530
rect 17155 2810 17175 2830
rect 17155 2760 17175 2780
rect 17155 2710 17175 2730
rect 17155 2660 17175 2680
rect 17155 2610 17175 2630
rect 17155 2560 17175 2580
rect 17155 2510 17175 2530
rect 17215 2810 17235 2830
rect 17215 2760 17235 2780
rect 17215 2710 17235 2730
rect 17215 2660 17235 2680
rect 17215 2610 17235 2630
rect 17215 2560 17235 2580
rect 17215 2510 17235 2530
rect 17275 2810 17295 2830
rect 17275 2760 17295 2780
rect 17275 2710 17295 2730
rect 17275 2660 17295 2680
rect 17275 2610 17295 2630
rect 17275 2560 17295 2580
rect 17275 2510 17295 2530
rect 17335 2810 17355 2830
rect 17335 2760 17355 2780
rect 17335 2710 17355 2730
rect 17335 2660 17355 2680
rect 17335 2610 17355 2630
rect 17335 2560 17355 2580
rect 17335 2510 17355 2530
rect 17395 2810 17415 2830
rect 17395 2760 17415 2780
rect 17395 2710 17415 2730
rect 17395 2660 17415 2680
rect 17395 2610 17415 2630
rect 17395 2560 17415 2580
rect 17395 2510 17415 2530
rect 17455 2810 17475 2830
rect 17455 2760 17475 2780
rect 17455 2710 17475 2730
rect 17455 2660 17475 2680
rect 17455 2610 17475 2630
rect 17455 2560 17475 2580
rect 17455 2510 17475 2530
rect 17515 2810 17535 2830
rect 17515 2760 17535 2780
rect 17515 2710 17535 2730
rect 17515 2660 17535 2680
rect 17515 2610 17535 2630
rect 17515 2560 17535 2580
rect 17515 2510 17535 2530
rect 17575 2810 17595 2830
rect 17575 2760 17595 2780
rect 17575 2710 17595 2730
rect 17575 2660 17595 2680
rect 17575 2610 17595 2630
rect 17575 2560 17595 2580
rect 17575 2510 17595 2530
rect 17635 2810 17655 2830
rect 17635 2760 17655 2780
rect 17635 2710 17655 2730
rect 17635 2660 17655 2680
rect 17635 2610 17655 2630
rect 17635 2560 17655 2580
rect 17635 2510 17655 2530
rect 17695 2810 17715 2830
rect 17695 2760 17715 2780
rect 17695 2710 17715 2730
rect 17695 2660 17715 2680
rect 17695 2610 17715 2630
rect 17695 2560 17715 2580
rect 17695 2510 17715 2530
rect 17755 2810 17775 2830
rect 17755 2760 17775 2780
rect 17755 2710 17775 2730
rect 17755 2660 17775 2680
rect 26025 2810 26045 2830
rect 26025 2760 26045 2780
rect 26025 2710 26045 2730
rect 26025 2660 26045 2680
rect 17755 2610 17775 2630
rect 17755 2560 17775 2580
rect 17755 2510 17775 2530
rect 18155 2620 18175 2640
rect 18155 2570 18175 2590
rect 18155 2520 18175 2540
rect 15675 2470 15695 2490
rect 18155 2470 18175 2490
rect 18210 2620 18230 2640
rect 18210 2570 18230 2590
rect 18210 2520 18230 2540
rect 18210 2470 18230 2490
rect 18265 2620 18285 2640
rect 18265 2570 18285 2590
rect 18265 2520 18285 2540
rect 18265 2470 18285 2490
rect 18320 2620 18340 2640
rect 18320 2570 18340 2590
rect 18320 2520 18340 2540
rect 18320 2470 18340 2490
rect 18375 2620 18395 2640
rect 18375 2570 18395 2590
rect 18375 2520 18395 2540
rect 18375 2470 18395 2490
rect 18430 2620 18450 2640
rect 18430 2570 18450 2590
rect 18430 2520 18450 2540
rect 18430 2470 18450 2490
rect 18485 2620 18505 2640
rect 18485 2570 18505 2590
rect 18485 2520 18505 2540
rect 18485 2470 18505 2490
rect 18540 2620 18560 2640
rect 18540 2570 18560 2590
rect 18540 2520 18560 2540
rect 18540 2470 18560 2490
rect 18595 2620 18615 2640
rect 18595 2570 18615 2590
rect 18595 2520 18615 2540
rect 18595 2470 18615 2490
rect 18650 2620 18670 2640
rect 18650 2570 18670 2590
rect 18650 2520 18670 2540
rect 18650 2470 18670 2490
rect 18705 2620 18725 2640
rect 18705 2570 18725 2590
rect 18705 2520 18725 2540
rect 18705 2470 18725 2490
rect 18760 2620 18780 2640
rect 18760 2570 18780 2590
rect 18760 2520 18780 2540
rect 18760 2470 18780 2490
rect 18815 2620 18835 2640
rect 18815 2570 18835 2590
rect 18815 2520 18835 2540
rect 18815 2470 18835 2490
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 4035 1965 4055 1985
rect 3955 1915 3975 1935
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 5235 1965 5255 1985
rect 25015 2620 25035 2640
rect 25015 2570 25035 2590
rect 25015 2520 25035 2540
rect 25015 2470 25035 2490
rect 25070 2620 25090 2640
rect 25070 2570 25090 2590
rect 25070 2520 25090 2540
rect 25070 2470 25090 2490
rect 25125 2620 25145 2640
rect 25125 2570 25145 2590
rect 25125 2520 25145 2540
rect 25125 2470 25145 2490
rect 25180 2620 25200 2640
rect 25180 2570 25200 2590
rect 25180 2520 25200 2540
rect 25180 2470 25200 2490
rect 25235 2620 25255 2640
rect 25235 2570 25255 2590
rect 25235 2520 25255 2540
rect 25235 2470 25255 2490
rect 25290 2620 25310 2640
rect 25290 2570 25310 2590
rect 25290 2520 25310 2540
rect 25290 2470 25310 2490
rect 25345 2620 25365 2640
rect 25345 2570 25365 2590
rect 25345 2520 25365 2540
rect 25345 2470 25365 2490
rect 25400 2620 25420 2640
rect 25400 2570 25420 2590
rect 25400 2520 25420 2540
rect 25400 2470 25420 2490
rect 25455 2620 25475 2640
rect 25455 2570 25475 2590
rect 25455 2520 25475 2540
rect 25455 2470 25475 2490
rect 25510 2620 25530 2640
rect 25510 2570 25530 2590
rect 25510 2520 25530 2540
rect 25510 2470 25530 2490
rect 25565 2620 25585 2640
rect 25565 2570 25585 2590
rect 25565 2520 25585 2540
rect 25565 2470 25585 2490
rect 25620 2620 25640 2640
rect 25620 2570 25640 2590
rect 25620 2520 25640 2540
rect 25620 2470 25640 2490
rect 25675 2620 25695 2640
rect 25675 2570 25695 2590
rect 25675 2520 25695 2540
rect 26025 2610 26045 2630
rect 26025 2560 26045 2580
rect 26025 2510 26045 2530
rect 26085 2810 26105 2830
rect 26085 2760 26105 2780
rect 26085 2710 26105 2730
rect 26085 2660 26105 2680
rect 26085 2610 26105 2630
rect 26085 2560 26105 2580
rect 26085 2510 26105 2530
rect 26145 2810 26165 2830
rect 26145 2760 26165 2780
rect 26145 2710 26165 2730
rect 26145 2660 26165 2680
rect 26145 2610 26165 2630
rect 26145 2560 26165 2580
rect 26145 2510 26165 2530
rect 26205 2810 26225 2830
rect 26205 2760 26225 2780
rect 26205 2710 26225 2730
rect 26205 2660 26225 2680
rect 26205 2610 26225 2630
rect 26205 2560 26225 2580
rect 26205 2510 26225 2530
rect 26265 2810 26285 2830
rect 26265 2760 26285 2780
rect 26265 2710 26285 2730
rect 26265 2660 26285 2680
rect 26265 2610 26285 2630
rect 26265 2560 26285 2580
rect 26265 2510 26285 2530
rect 26325 2810 26345 2830
rect 26325 2760 26345 2780
rect 26325 2710 26345 2730
rect 26325 2660 26345 2680
rect 26325 2610 26345 2630
rect 26325 2560 26345 2580
rect 26325 2510 26345 2530
rect 26385 2810 26405 2830
rect 26385 2760 26405 2780
rect 26385 2710 26405 2730
rect 26385 2660 26405 2680
rect 26385 2610 26405 2630
rect 26385 2560 26405 2580
rect 26385 2510 26405 2530
rect 26445 2810 26465 2830
rect 26445 2760 26465 2780
rect 26445 2710 26465 2730
rect 26445 2660 26465 2680
rect 26445 2610 26465 2630
rect 26445 2560 26465 2580
rect 26445 2510 26465 2530
rect 26505 2810 26525 2830
rect 26505 2760 26525 2780
rect 26505 2710 26525 2730
rect 26505 2660 26525 2680
rect 26505 2610 26525 2630
rect 26505 2560 26525 2580
rect 26505 2510 26525 2530
rect 26565 2810 26585 2830
rect 26565 2760 26585 2780
rect 26565 2710 26585 2730
rect 26565 2660 26585 2680
rect 26565 2610 26585 2630
rect 26565 2560 26585 2580
rect 26565 2510 26585 2530
rect 26625 2810 26645 2830
rect 26625 2760 26645 2780
rect 26625 2710 26645 2730
rect 26625 2660 26645 2680
rect 26625 2610 26645 2630
rect 26625 2560 26645 2580
rect 26625 2510 26645 2530
rect 26685 2810 26705 2830
rect 26685 2760 26705 2780
rect 26685 2710 26705 2730
rect 26685 2660 26705 2680
rect 26685 2610 26705 2630
rect 26685 2560 26705 2580
rect 26685 2510 26705 2530
rect 26745 2810 26765 2830
rect 26745 2760 26765 2780
rect 26745 2710 26765 2730
rect 26745 2660 26765 2680
rect 26745 2610 26765 2630
rect 26745 2560 26765 2580
rect 26745 2510 26765 2530
rect 25675 2470 25695 2490
rect 27045 2810 27065 2830
rect 27045 2760 27065 2780
rect 27045 2710 27065 2730
rect 27045 2660 27065 2680
rect 27045 2610 27065 2630
rect 27045 2560 27065 2580
rect 27045 2510 27065 2530
rect 27105 2810 27125 2830
rect 27105 2760 27125 2780
rect 27105 2710 27125 2730
rect 27105 2660 27125 2680
rect 27105 2610 27125 2630
rect 27105 2560 27125 2580
rect 27105 2510 27125 2530
rect 27165 2810 27185 2830
rect 27165 2760 27185 2780
rect 27165 2710 27185 2730
rect 27165 2660 27185 2680
rect 27165 2610 27185 2630
rect 27165 2560 27185 2580
rect 27165 2510 27185 2530
rect 27225 2810 27245 2830
rect 27225 2760 27245 2780
rect 27225 2710 27245 2730
rect 27225 2660 27245 2680
rect 27225 2610 27245 2630
rect 27225 2560 27245 2580
rect 27225 2510 27245 2530
rect 27285 2810 27305 2830
rect 27285 2760 27305 2780
rect 27285 2710 27305 2730
rect 27285 2660 27305 2680
rect 27285 2610 27305 2630
rect 27285 2560 27305 2580
rect 27285 2510 27305 2530
rect 27345 2810 27365 2830
rect 27345 2760 27365 2780
rect 27345 2710 27365 2730
rect 27345 2660 27365 2680
rect 27345 2610 27365 2630
rect 27345 2560 27365 2580
rect 27345 2510 27365 2530
rect 27405 2810 27425 2830
rect 27405 2760 27425 2780
rect 27405 2710 27425 2730
rect 27405 2660 27425 2680
rect 27405 2610 27425 2630
rect 27405 2560 27425 2580
rect 27405 2510 27425 2530
rect 27465 2810 27485 2830
rect 27465 2760 27485 2780
rect 27465 2710 27485 2730
rect 27465 2660 27485 2680
rect 27465 2610 27485 2630
rect 27465 2560 27485 2580
rect 27465 2510 27485 2530
rect 27525 2810 27545 2830
rect 27525 2760 27545 2780
rect 27525 2710 27545 2730
rect 27525 2660 27545 2680
rect 27525 2610 27545 2630
rect 27525 2560 27545 2580
rect 27525 2510 27545 2530
rect 27585 2810 27605 2830
rect 27585 2760 27605 2780
rect 27585 2710 27605 2730
rect 27585 2660 27605 2680
rect 27585 2610 27605 2630
rect 27585 2560 27605 2580
rect 27585 2510 27605 2530
rect 27645 2810 27665 2830
rect 27645 2760 27665 2780
rect 27645 2710 27665 2730
rect 27645 2660 27665 2680
rect 27645 2610 27665 2630
rect 27645 2560 27665 2580
rect 27645 2510 27665 2530
rect 27705 2810 27725 2830
rect 27705 2760 27725 2780
rect 27705 2710 27725 2730
rect 27705 2660 27725 2680
rect 27705 2610 27725 2630
rect 27705 2560 27725 2580
rect 27705 2510 27725 2530
rect 27765 2810 27785 2830
rect 27765 2760 27785 2780
rect 27765 2710 27785 2730
rect 27765 2660 27785 2680
rect 27765 2610 27785 2630
rect 27765 2560 27785 2580
rect 27765 2510 27785 2530
rect 28155 2670 28175 2690
rect 28155 2620 28175 2640
rect 28155 2570 28175 2590
rect 28155 2520 28175 2540
rect 28210 2670 28230 2690
rect 28210 2620 28230 2640
rect 28210 2570 28230 2590
rect 28210 2520 28230 2540
rect 28265 2670 28285 2690
rect 28265 2620 28285 2640
rect 28265 2570 28285 2590
rect 28265 2520 28285 2540
rect 28320 2670 28340 2690
rect 28320 2620 28340 2640
rect 28320 2570 28340 2590
rect 28320 2520 28340 2540
rect 28375 2670 28395 2690
rect 28375 2620 28395 2640
rect 28375 2570 28395 2590
rect 28375 2520 28395 2540
rect 28430 2670 28450 2690
rect 28430 2620 28450 2640
rect 28430 2570 28450 2590
rect 28430 2520 28450 2540
rect 28485 2670 28505 2690
rect 28485 2620 28505 2640
rect 28485 2570 28505 2590
rect 28485 2520 28505 2540
rect 28540 2670 28560 2690
rect 28540 2620 28560 2640
rect 28540 2570 28560 2590
rect 28540 2520 28560 2540
rect 28595 2670 28615 2690
rect 28595 2620 28615 2640
rect 28595 2570 28615 2590
rect 28595 2520 28615 2540
rect 28650 2670 28670 2690
rect 28650 2620 28670 2640
rect 28650 2570 28670 2590
rect 28650 2520 28670 2540
rect 28705 2670 28725 2690
rect 28705 2620 28725 2640
rect 28705 2570 28725 2590
rect 28705 2520 28725 2540
rect 28760 2670 28780 2690
rect 28760 2620 28780 2640
rect 28760 2570 28780 2590
rect 28760 2520 28780 2540
rect 28815 2670 28835 2690
rect 28815 2620 28835 2640
rect 28815 2570 28835 2590
rect 28815 2520 28835 2540
rect 5235 1915 5255 1935
<< psubdiff >>
rect 29035 3680 29315 3700
rect 29035 3375 29055 3680
rect 29035 2980 29055 3280
rect 29295 3375 29315 3680
rect 29295 2980 29315 3280
rect 29035 2960 29135 2980
rect 29215 2960 29315 2980
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 14965 2250 15005 2265
rect 14965 2230 14975 2250
rect 14995 2230 15005 2250
rect 14965 2200 15005 2230
rect 14965 2180 14975 2200
rect 14995 2180 15005 2200
rect 14965 2150 15005 2180
rect 14965 2130 14975 2150
rect 14995 2130 15005 2150
rect 14965 2100 15005 2130
rect 14965 2080 14975 2100
rect 14995 2080 15005 2100
rect 14965 2050 15005 2080
rect 14965 2030 14975 2050
rect 14995 2030 15005 2050
rect 14965 2000 15005 2030
rect 14965 1980 14975 2000
rect 14995 1980 15005 2000
rect 14965 1965 15005 1980
rect 15705 2250 15745 2265
rect 15705 2230 15715 2250
rect 15735 2230 15745 2250
rect 15705 2200 15745 2230
rect 15705 2180 15715 2200
rect 15735 2180 15745 2200
rect 18105 2250 18145 2265
rect 18105 2230 18115 2250
rect 18135 2230 18145 2250
rect 18105 2200 18145 2230
rect 15705 2150 15745 2180
rect 18105 2180 18115 2200
rect 18135 2180 18145 2200
rect 15705 2130 15715 2150
rect 15735 2130 15745 2150
rect 18105 2150 18145 2180
rect 18105 2130 18115 2150
rect 18135 2130 18145 2150
rect 15705 2100 15745 2130
rect 15705 2080 15715 2100
rect 15735 2080 15745 2100
rect 15705 2050 15745 2080
rect 15705 2030 15715 2050
rect 15735 2030 15745 2050
rect 15705 2000 15745 2030
rect 15705 1980 15715 2000
rect 15735 1980 15745 2000
rect 16235 2115 16275 2130
rect 16235 2095 16245 2115
rect 16265 2095 16275 2115
rect 16235 2065 16275 2095
rect 16235 2045 16245 2065
rect 16265 2045 16275 2065
rect 16235 2015 16275 2045
rect 16235 1995 16245 2015
rect 16265 1995 16275 2015
rect 16235 1980 16275 1995
rect 17525 2115 17565 2130
rect 17525 2095 17535 2115
rect 17555 2095 17565 2115
rect 17525 2065 17565 2095
rect 17525 2045 17535 2065
rect 17555 2045 17565 2065
rect 17525 2015 17565 2045
rect 17525 1995 17535 2015
rect 17555 1995 17565 2015
rect 17525 1980 17565 1995
rect 18105 2100 18145 2130
rect 18105 2080 18115 2100
rect 18135 2080 18145 2100
rect 18105 2050 18145 2080
rect 18105 2030 18115 2050
rect 18135 2030 18145 2050
rect 18105 2000 18145 2030
rect 18105 1980 18115 2000
rect 18135 1980 18145 2000
rect 15705 1965 15745 1980
rect 18105 1965 18145 1980
rect 18845 2250 18885 2265
rect 18845 2230 18855 2250
rect 18875 2230 18885 2250
rect 18845 2200 18885 2230
rect 18845 2180 18855 2200
rect 18875 2180 18885 2200
rect 18845 2150 18885 2180
rect 18845 2130 18855 2150
rect 18875 2130 18885 2150
rect 18845 2100 18885 2130
rect 18845 2080 18855 2100
rect 18875 2080 18885 2100
rect 18845 2050 18885 2080
rect 18845 2030 18855 2050
rect 18875 2030 18885 2050
rect 18845 2000 18885 2030
rect 28995 2665 29135 2685
rect 29215 2665 29350 2685
rect 28095 2320 28455 2340
rect 28535 2320 28895 2340
rect 24965 2250 25005 2265
rect 24965 2230 24975 2250
rect 24995 2230 25005 2250
rect 24965 2200 25005 2230
rect 24965 2180 24975 2200
rect 24995 2180 25005 2200
rect 24965 2150 25005 2180
rect 24965 2130 24975 2150
rect 24995 2130 25005 2150
rect 24965 2100 25005 2130
rect 24965 2080 24975 2100
rect 24995 2080 25005 2100
rect 24965 2050 25005 2080
rect 24965 2030 24975 2050
rect 24995 2030 25005 2050
rect 18845 1980 18855 2000
rect 18875 1980 18885 2000
rect 18845 1965 18885 1980
rect 24965 2000 25005 2030
rect 24965 1980 24975 2000
rect 24995 1980 25005 2000
rect 24965 1965 25005 1980
rect 25705 2250 25745 2265
rect 25705 2230 25715 2250
rect 25735 2230 25745 2250
rect 25705 2200 25745 2230
rect 25705 2180 25715 2200
rect 25735 2180 25745 2200
rect 25705 2150 25745 2180
rect 25705 2130 25715 2150
rect 25735 2130 25745 2150
rect 25705 2100 25745 2130
rect 25705 2080 25715 2100
rect 25735 2080 25745 2100
rect 25705 2050 25745 2080
rect 25705 2030 25715 2050
rect 25735 2030 25745 2050
rect 25705 2000 25745 2030
rect 25705 1980 25715 2000
rect 25735 1980 25745 2000
rect 25705 1965 25745 1980
rect 26225 2205 26860 2225
rect 26940 2205 27575 2225
rect 26225 2090 26245 2205
rect 26225 1905 26245 2010
rect 27555 2090 27575 2205
rect 27555 1905 27575 2010
rect 26225 1885 26860 1905
rect 26940 1885 27575 1905
rect 28095 2135 28115 2320
rect 28095 1870 28115 2055
rect 28875 2135 28895 2320
rect 28875 1870 28895 2055
rect 28995 2335 29015 2665
rect 28995 1925 29015 2255
rect 29330 2335 29350 2665
rect 29330 1925 29350 2255
rect 28995 1905 29135 1925
rect 29215 1905 29350 1925
rect 28095 1850 28455 1870
rect 28535 1850 28895 1870
rect 25940 1800 26860 1820
rect 26940 1800 27860 1820
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
rect 3980 1650 4030 1665
rect 3980 1630 3995 1650
rect 4015 1630 4030 1650
rect 3980 1615 4030 1630
rect 14965 1640 15005 1655
rect 14965 1620 14975 1640
rect 14995 1620 15005 1640
rect 5065 1060 5105 1075
rect 5065 1040 5075 1060
rect 5095 1040 5105 1060
rect 5065 1010 5105 1040
rect 5065 990 5075 1010
rect 5095 990 5105 1010
rect 5065 975 5105 990
rect 14965 1590 15005 1620
rect 14965 1570 14975 1590
rect 14995 1570 15005 1590
rect 14965 1540 15005 1570
rect 14965 1520 14975 1540
rect 14995 1520 15005 1540
rect 14965 1490 15005 1520
rect 14965 1470 14975 1490
rect 14995 1470 15005 1490
rect 14965 1440 15005 1470
rect 14965 1420 14975 1440
rect 14995 1420 15005 1440
rect 14965 1390 15005 1420
rect 14965 1370 14975 1390
rect 14995 1370 15005 1390
rect 14965 1340 15005 1370
rect 14965 1320 14975 1340
rect 14995 1320 15005 1340
rect 14965 1290 15005 1320
rect 14965 1270 14975 1290
rect 14995 1270 15005 1290
rect 14965 1240 15005 1270
rect 14965 1220 14975 1240
rect 14995 1220 15005 1240
rect 14965 1190 15005 1220
rect 14965 1170 14975 1190
rect 14995 1170 15005 1190
rect 14965 1140 15005 1170
rect 14965 1120 14975 1140
rect 14995 1120 15005 1140
rect 14965 1090 15005 1120
rect 14965 1070 14975 1090
rect 14995 1070 15005 1090
rect 14965 1040 15005 1070
rect 14965 1020 14975 1040
rect 14995 1020 15005 1040
rect 14965 990 15005 1020
rect 14965 970 14975 990
rect 14995 970 15005 990
rect 14965 955 15005 970
rect 15645 1640 15685 1655
rect 15645 1620 15655 1640
rect 15675 1620 15685 1640
rect 15645 1590 15685 1620
rect 15645 1570 15655 1590
rect 15675 1570 15685 1590
rect 15645 1540 15685 1570
rect 15645 1520 15655 1540
rect 15675 1520 15685 1540
rect 15645 1490 15685 1520
rect 15990 1650 16030 1665
rect 15990 1630 16000 1650
rect 16020 1630 16030 1650
rect 15990 1600 16030 1630
rect 15990 1580 16000 1600
rect 16020 1580 16030 1600
rect 15990 1550 16030 1580
rect 15990 1530 16000 1550
rect 16020 1530 16030 1550
rect 15990 1515 16030 1530
rect 16730 1650 16770 1665
rect 16730 1630 16740 1650
rect 16760 1630 16770 1650
rect 16730 1600 16770 1630
rect 16730 1580 16740 1600
rect 16760 1580 16770 1600
rect 16730 1550 16770 1580
rect 16730 1530 16740 1550
rect 16760 1530 16770 1550
rect 16730 1515 16770 1530
rect 17030 1650 17070 1665
rect 17030 1630 17040 1650
rect 17060 1630 17070 1650
rect 17030 1600 17070 1630
rect 17030 1580 17040 1600
rect 17060 1580 17070 1600
rect 17030 1550 17070 1580
rect 17030 1530 17040 1550
rect 17060 1530 17070 1550
rect 17030 1515 17070 1530
rect 17770 1650 17810 1665
rect 17770 1630 17780 1650
rect 17800 1630 17810 1650
rect 17770 1600 17810 1630
rect 17770 1580 17780 1600
rect 17800 1580 17810 1600
rect 17770 1550 17810 1580
rect 17770 1530 17780 1550
rect 17800 1530 17810 1550
rect 17770 1515 17810 1530
rect 18165 1640 18205 1655
rect 18165 1620 18175 1640
rect 18195 1620 18205 1640
rect 18165 1590 18205 1620
rect 18165 1570 18175 1590
rect 18195 1570 18205 1590
rect 18165 1540 18205 1570
rect 18165 1520 18175 1540
rect 18195 1520 18205 1540
rect 15645 1470 15655 1490
rect 15675 1470 15685 1490
rect 15645 1440 15685 1470
rect 18165 1490 18205 1520
rect 18165 1470 18175 1490
rect 18195 1470 18205 1490
rect 15645 1420 15655 1440
rect 15675 1420 15685 1440
rect 15645 1390 15685 1420
rect 15645 1370 15655 1390
rect 15675 1370 15685 1390
rect 15645 1340 15685 1370
rect 15645 1320 15655 1340
rect 15675 1320 15685 1340
rect 15645 1290 15685 1320
rect 15645 1270 15655 1290
rect 15675 1270 15685 1290
rect 15645 1240 15685 1270
rect 18165 1440 18205 1470
rect 18165 1420 18175 1440
rect 18195 1420 18205 1440
rect 18165 1390 18205 1420
rect 18165 1370 18175 1390
rect 18195 1370 18205 1390
rect 18165 1340 18205 1370
rect 18165 1320 18175 1340
rect 18195 1320 18205 1340
rect 18165 1290 18205 1320
rect 18165 1270 18175 1290
rect 18195 1270 18205 1290
rect 15645 1220 15655 1240
rect 15675 1220 15685 1240
rect 15645 1190 15685 1220
rect 15645 1170 15655 1190
rect 15675 1170 15685 1190
rect 18165 1240 18205 1270
rect 18165 1220 18175 1240
rect 18195 1220 18205 1240
rect 18165 1190 18205 1220
rect 15645 1140 15685 1170
rect 15645 1120 15655 1140
rect 15675 1120 15685 1140
rect 15645 1090 15685 1120
rect 15645 1070 15655 1090
rect 15675 1070 15685 1090
rect 15645 1040 15685 1070
rect 15645 1020 15655 1040
rect 15675 1020 15685 1040
rect 15645 990 15685 1020
rect 15645 970 15655 990
rect 15675 970 15685 990
rect 15645 955 15685 970
rect 16165 1170 16205 1185
rect 16165 1150 16175 1170
rect 16195 1150 16205 1170
rect 16165 1120 16205 1150
rect 16165 1100 16175 1120
rect 16195 1100 16205 1120
rect 16165 1070 16205 1100
rect 16165 1050 16175 1070
rect 16195 1050 16205 1070
rect 16165 1020 16205 1050
rect 16165 1000 16175 1020
rect 16195 1000 16205 1020
rect 16165 970 16205 1000
rect 16165 950 16175 970
rect 16195 950 16205 970
rect 16165 935 16205 950
rect 17620 1170 17660 1185
rect 17620 1150 17630 1170
rect 17650 1150 17660 1170
rect 17620 1120 17660 1150
rect 17620 1100 17630 1120
rect 17650 1100 17660 1120
rect 17620 1070 17660 1100
rect 17620 1050 17630 1070
rect 17650 1050 17660 1070
rect 17620 1020 17660 1050
rect 17620 1000 17630 1020
rect 17650 1000 17660 1020
rect 17620 970 17660 1000
rect 17620 950 17630 970
rect 17650 950 17660 970
rect 18165 1170 18175 1190
rect 18195 1170 18205 1190
rect 18165 1140 18205 1170
rect 18165 1120 18175 1140
rect 18195 1120 18205 1140
rect 18165 1090 18205 1120
rect 18165 1070 18175 1090
rect 18195 1070 18205 1090
rect 18165 1040 18205 1070
rect 18165 1020 18175 1040
rect 18195 1020 18205 1040
rect 18165 990 18205 1020
rect 18165 970 18175 990
rect 18195 970 18205 990
rect 18165 955 18205 970
rect 18845 1640 18885 1655
rect 18845 1620 18855 1640
rect 18875 1620 18885 1640
rect 18845 1590 18885 1620
rect 24965 1640 25005 1655
rect 24965 1620 24975 1640
rect 24995 1620 25005 1640
rect 18845 1570 18855 1590
rect 18875 1570 18885 1590
rect 18845 1540 18885 1570
rect 18845 1520 18855 1540
rect 18875 1520 18885 1540
rect 18845 1490 18885 1520
rect 18845 1470 18855 1490
rect 18875 1470 18885 1490
rect 18845 1440 18885 1470
rect 18845 1420 18855 1440
rect 18875 1420 18885 1440
rect 18845 1390 18885 1420
rect 18845 1370 18855 1390
rect 18875 1370 18885 1390
rect 18845 1340 18885 1370
rect 18845 1320 18855 1340
rect 18875 1320 18885 1340
rect 18845 1290 18885 1320
rect 18845 1270 18855 1290
rect 18875 1270 18885 1290
rect 18845 1240 18885 1270
rect 18845 1220 18855 1240
rect 18875 1220 18885 1240
rect 18845 1190 18885 1220
rect 18845 1170 18855 1190
rect 18875 1170 18885 1190
rect 18845 1140 18885 1170
rect 18845 1120 18855 1140
rect 18875 1120 18885 1140
rect 18845 1090 18885 1120
rect 18845 1070 18855 1090
rect 18875 1070 18885 1090
rect 18845 1040 18885 1070
rect 18845 1020 18855 1040
rect 18875 1020 18885 1040
rect 18845 990 18885 1020
rect 18845 970 18855 990
rect 18875 970 18885 990
rect 18845 955 18885 970
rect 17620 935 17660 950
rect 24965 1590 25005 1620
rect 24965 1570 24975 1590
rect 24995 1570 25005 1590
rect 24965 1540 25005 1570
rect 24965 1520 24975 1540
rect 24995 1520 25005 1540
rect 24965 1490 25005 1520
rect 24965 1470 24975 1490
rect 24995 1470 25005 1490
rect 24965 1440 25005 1470
rect 24965 1420 24975 1440
rect 24995 1420 25005 1440
rect 24965 1390 25005 1420
rect 24965 1370 24975 1390
rect 24995 1370 25005 1390
rect 24965 1340 25005 1370
rect 24965 1320 24975 1340
rect 24995 1320 25005 1340
rect 24965 1290 25005 1320
rect 24965 1270 24975 1290
rect 24995 1270 25005 1290
rect 24965 1240 25005 1270
rect 24965 1220 24975 1240
rect 24995 1220 25005 1240
rect 24965 1190 25005 1220
rect 24965 1170 24975 1190
rect 24995 1170 25005 1190
rect 24965 1140 25005 1170
rect 24965 1120 24975 1140
rect 24995 1120 25005 1140
rect 24965 1090 25005 1120
rect 24965 1070 24975 1090
rect 24995 1070 25005 1090
rect 24965 1040 25005 1070
rect 24965 1020 24975 1040
rect 24995 1020 25005 1040
rect 24965 990 25005 1020
rect 24965 970 24975 990
rect 24995 970 25005 990
rect 24965 955 25005 970
rect 25645 1640 25685 1655
rect 25645 1620 25655 1640
rect 25675 1620 25685 1640
rect 25645 1590 25685 1620
rect 25645 1570 25655 1590
rect 25675 1570 25685 1590
rect 25645 1540 25685 1570
rect 25645 1520 25655 1540
rect 25675 1520 25685 1540
rect 25645 1490 25685 1520
rect 25645 1470 25655 1490
rect 25675 1470 25685 1490
rect 25645 1440 25685 1470
rect 25645 1420 25655 1440
rect 25675 1420 25685 1440
rect 25645 1390 25685 1420
rect 25645 1370 25655 1390
rect 25675 1370 25685 1390
rect 25645 1340 25685 1370
rect 25940 1630 25960 1800
rect 25940 1380 25960 1550
rect 26730 1650 26770 1665
rect 26730 1630 26740 1650
rect 26760 1630 26770 1650
rect 26730 1600 26770 1630
rect 26730 1580 26740 1600
rect 26760 1580 26770 1600
rect 26730 1550 26770 1580
rect 26730 1530 26740 1550
rect 26760 1530 26770 1550
rect 26730 1515 26770 1530
rect 27030 1650 27070 1665
rect 27030 1630 27040 1650
rect 27060 1630 27070 1650
rect 27030 1600 27070 1630
rect 27030 1580 27040 1600
rect 27060 1580 27070 1600
rect 27030 1550 27070 1580
rect 27030 1530 27040 1550
rect 27060 1530 27070 1550
rect 27030 1515 27070 1530
rect 27840 1630 27860 1800
rect 27840 1380 27860 1550
rect 25940 1360 26860 1380
rect 26940 1360 27860 1380
rect 28155 1730 28485 1750
rect 28565 1730 28895 1750
rect 25645 1320 25655 1340
rect 25675 1320 25685 1340
rect 25645 1290 25685 1320
rect 25645 1270 25655 1290
rect 25675 1270 25685 1290
rect 25645 1240 25685 1270
rect 25645 1220 25655 1240
rect 25675 1220 25685 1240
rect 25645 1190 25685 1220
rect 28155 1345 28175 1730
rect 25645 1170 25655 1190
rect 25675 1170 25685 1190
rect 25645 1140 25685 1170
rect 25645 1120 25655 1140
rect 25675 1120 25685 1140
rect 25645 1090 25685 1120
rect 25645 1070 25655 1090
rect 25675 1070 25685 1090
rect 25645 1040 25685 1070
rect 25645 1020 25655 1040
rect 25675 1020 25685 1040
rect 25645 990 25685 1020
rect 25645 970 25655 990
rect 25675 970 25685 990
rect 25645 955 25685 970
rect 26155 1175 26845 1195
rect 26925 1175 27675 1195
rect 26155 980 26175 1175
rect 2955 865 2995 880
rect 2955 845 2965 865
rect 2985 845 2995 865
rect 2955 815 2995 845
rect 2955 795 2965 815
rect 2985 795 2995 815
rect 2955 780 2995 795
rect 5015 865 5055 880
rect 5015 845 5025 865
rect 5045 845 5055 865
rect 5015 815 5055 845
rect 5015 795 5025 815
rect 5045 795 5055 815
rect 5015 780 5055 795
rect 26155 755 26175 900
rect 27655 980 27675 1175
rect 27655 755 27675 900
rect 28155 880 28175 1265
rect 28875 1345 28895 1730
rect 28875 880 28895 1265
rect 28155 860 28485 880
rect 28565 860 28895 880
rect 28985 1675 29065 1695
rect 29145 1675 29220 1695
rect 28985 1300 29005 1675
rect 28985 860 29005 1220
rect 29200 1300 29220 1675
rect 29200 860 29220 1220
rect 28985 840 29065 860
rect 29145 840 29220 860
rect 16840 735 16880 750
rect 16840 715 16850 735
rect 16870 715 16880 735
rect 16840 700 16880 715
rect 17580 735 17620 750
rect 26155 735 26845 755
rect 26925 735 27675 755
rect 17580 715 17590 735
rect 17610 715 17620 735
rect 17580 700 17620 715
rect 26210 625 26355 645
rect 26435 625 26585 645
rect 26210 555 26230 625
rect 26565 555 26585 625
rect 26210 415 26230 475
rect 26565 415 26585 475
rect 26210 395 26355 415
rect 26435 395 26585 415
rect 26830 625 27190 645
rect 27270 625 27630 645
rect 26830 555 26850 625
rect 27610 555 27630 625
rect 26830 425 26850 475
rect 27610 425 27630 475
rect 26830 405 27190 425
rect 27270 405 27630 425
<< nsubdiff >>
rect 26205 4950 26520 4970
rect 26600 4950 26955 4970
rect 26205 4865 26225 4950
rect 26935 4865 26955 4950
rect 26205 4715 26225 4785
rect 26935 4715 26955 4785
rect 26205 4695 26520 4715
rect 26600 4695 26955 4715
rect 27185 4925 27460 4945
rect 27540 4925 27805 4945
rect 27185 4860 27205 4925
rect 27785 4865 27805 4925
rect 27185 4715 27205 4780
rect 27785 4715 27805 4780
rect 27185 4695 27460 4715
rect 27540 4695 27805 4715
rect 26200 4505 26835 4525
rect 26915 4505 27550 4525
rect 26200 4445 26220 4505
rect 27530 4445 27550 4505
rect 16165 4325 16205 4353
rect 16165 4305 16175 4325
rect 16195 4305 16205 4325
rect 16165 4290 16205 4305
rect 16425 4325 16465 4353
rect 16425 4305 16435 4325
rect 16455 4305 16465 4325
rect 16425 4290 16465 4305
rect 16495 4340 16535 4370
rect 16495 4320 16505 4340
rect 16525 4320 16535 4340
rect 16495 4290 16535 4320
rect 16935 4340 16975 4370
rect 16935 4320 16945 4340
rect 16965 4320 16975 4340
rect 16935 4290 16975 4320
rect 17145 4325 17185 4345
rect 17145 4305 17155 4325
rect 17175 4305 17185 4325
rect 17145 4285 17185 4305
rect 17705 4325 17745 4345
rect 17705 4305 17715 4325
rect 17735 4305 17745 4325
rect 17705 4285 17745 4305
rect 26200 4305 26220 4365
rect 27530 4305 27550 4365
rect 26200 4285 26835 4305
rect 26915 4285 27550 4305
rect 16210 4090 16250 4105
rect 16210 4070 16220 4090
rect 16240 4070 16250 4090
rect 16210 4055 16250 4070
rect 17500 4090 17540 4105
rect 17500 4070 17510 4090
rect 17530 4070 17540 4090
rect 17500 4055 17540 4070
rect 26150 4095 26875 4115
rect 26955 4095 27680 4115
rect 26150 4035 26170 4095
rect 27660 4035 27680 4095
rect 26150 3895 26170 3955
rect 27660 3895 27680 3955
rect 26150 3875 26875 3895
rect 26955 3875 27680 3895
rect 16155 3785 16195 3800
rect 16155 3765 16165 3785
rect 16185 3765 16195 3785
rect 16155 3750 16195 3765
rect 16895 3785 16935 3800
rect 16895 3765 16905 3785
rect 16925 3765 16935 3785
rect 16895 3750 16935 3765
rect 17635 3785 17675 3800
rect 17635 3765 17645 3785
rect 17665 3765 17675 3785
rect 17635 3750 17675 3765
rect 28095 3740 28455 3760
rect 28535 3740 28895 3760
rect 26170 3680 26860 3700
rect 26940 3680 27630 3700
rect 14965 3570 15005 3585
rect 14965 3550 14975 3570
rect 14995 3550 15005 3570
rect 14965 3520 15005 3550
rect 14965 3500 14975 3520
rect 14995 3500 15005 3520
rect 14965 3470 15005 3500
rect 14965 3450 14975 3470
rect 14995 3450 15005 3470
rect 14965 3420 15005 3450
rect 14965 3400 14975 3420
rect 14995 3400 15005 3420
rect 14965 3370 15005 3400
rect 14965 3350 14975 3370
rect 14995 3350 15005 3370
rect 14965 3320 15005 3350
rect 14965 3300 14975 3320
rect 14995 3300 15005 3320
rect 14965 3270 15005 3300
rect 14965 3250 14975 3270
rect 14995 3250 15005 3270
rect 14965 3220 15005 3250
rect 14965 3200 14975 3220
rect 14995 3200 15005 3220
rect 14965 3170 15005 3200
rect 14965 3150 14975 3170
rect 14995 3150 15005 3170
rect 14965 3120 15005 3150
rect 14965 3100 14975 3120
rect 14995 3100 15005 3120
rect 14965 3070 15005 3100
rect 14965 3050 14975 3070
rect 14995 3050 15005 3070
rect 14965 3020 15005 3050
rect 14965 3000 14975 3020
rect 14995 3000 15005 3020
rect 14965 2985 15005 3000
rect 15705 3570 15745 3585
rect 15705 3550 15715 3570
rect 15735 3550 15745 3570
rect 15705 3520 15745 3550
rect 18105 3570 18145 3585
rect 18105 3550 18115 3570
rect 18135 3550 18145 3570
rect 15705 3500 15715 3520
rect 15735 3500 15745 3520
rect 15705 3470 15745 3500
rect 15705 3450 15715 3470
rect 15735 3450 15745 3470
rect 15705 3420 15745 3450
rect 15705 3400 15715 3420
rect 15735 3400 15745 3420
rect 15705 3370 15745 3400
rect 15705 3350 15715 3370
rect 15735 3350 15745 3370
rect 15705 3320 15745 3350
rect 15705 3300 15715 3320
rect 15735 3300 15745 3320
rect 15705 3270 15745 3300
rect 15705 3250 15715 3270
rect 15735 3250 15745 3270
rect 15705 3220 15745 3250
rect 15705 3200 15715 3220
rect 15735 3200 15745 3220
rect 15705 3170 15745 3200
rect 15705 3150 15715 3170
rect 15735 3150 15745 3170
rect 15705 3120 15745 3150
rect 16180 3510 16220 3525
rect 16180 3490 16190 3510
rect 16210 3490 16220 3510
rect 16180 3460 16220 3490
rect 16180 3440 16190 3460
rect 16210 3440 16220 3460
rect 16180 3410 16220 3440
rect 16180 3390 16190 3410
rect 16210 3390 16220 3410
rect 16180 3360 16220 3390
rect 16180 3340 16190 3360
rect 16210 3340 16220 3360
rect 16180 3310 16220 3340
rect 16180 3290 16190 3310
rect 16210 3290 16220 3310
rect 16180 3260 16220 3290
rect 16180 3240 16190 3260
rect 16210 3240 16220 3260
rect 16180 3210 16220 3240
rect 16180 3190 16190 3210
rect 16210 3190 16220 3210
rect 16180 3160 16220 3190
rect 16180 3140 16190 3160
rect 16210 3140 16220 3160
rect 16180 3125 16220 3140
rect 17580 3510 17620 3525
rect 17580 3490 17590 3510
rect 17610 3490 17620 3510
rect 17580 3460 17620 3490
rect 17580 3440 17590 3460
rect 17610 3440 17620 3460
rect 17580 3410 17620 3440
rect 17580 3390 17590 3410
rect 17610 3390 17620 3410
rect 17580 3360 17620 3390
rect 17580 3340 17590 3360
rect 17610 3340 17620 3360
rect 17580 3310 17620 3340
rect 17580 3290 17590 3310
rect 17610 3290 17620 3310
rect 17580 3260 17620 3290
rect 17580 3240 17590 3260
rect 17610 3240 17620 3260
rect 17580 3210 17620 3240
rect 17580 3190 17590 3210
rect 17610 3190 17620 3210
rect 17580 3160 17620 3190
rect 17580 3140 17590 3160
rect 17610 3140 17620 3160
rect 17580 3125 17620 3140
rect 18105 3520 18145 3550
rect 18105 3500 18115 3520
rect 18135 3500 18145 3520
rect 18105 3470 18145 3500
rect 18105 3450 18115 3470
rect 18135 3450 18145 3470
rect 18105 3420 18145 3450
rect 18105 3400 18115 3420
rect 18135 3400 18145 3420
rect 18105 3370 18145 3400
rect 18105 3350 18115 3370
rect 18135 3350 18145 3370
rect 18105 3320 18145 3350
rect 18105 3300 18115 3320
rect 18135 3300 18145 3320
rect 18105 3270 18145 3300
rect 18105 3250 18115 3270
rect 18135 3250 18145 3270
rect 18105 3220 18145 3250
rect 18105 3200 18115 3220
rect 18135 3200 18145 3220
rect 18105 3170 18145 3200
rect 18105 3150 18115 3170
rect 18135 3150 18145 3170
rect 15705 3100 15715 3120
rect 15735 3100 15745 3120
rect 18105 3120 18145 3150
rect 18105 3100 18115 3120
rect 18135 3100 18145 3120
rect 15705 3070 15745 3100
rect 18105 3070 18145 3100
rect 15705 3050 15715 3070
rect 15735 3050 15745 3070
rect 15705 3020 15745 3050
rect 15705 3000 15715 3020
rect 15735 3000 15745 3020
rect 15705 2985 15745 3000
rect 18105 3050 18115 3070
rect 18135 3050 18145 3070
rect 18105 3020 18145 3050
rect 18105 3000 18115 3020
rect 18135 3000 18145 3020
rect 18105 2985 18145 3000
rect 18845 3570 18885 3585
rect 18845 3550 18855 3570
rect 18875 3550 18885 3570
rect 18845 3520 18885 3550
rect 24965 3570 25005 3585
rect 24965 3550 24975 3570
rect 24995 3550 25005 3570
rect 24965 3520 25005 3550
rect 18845 3500 18855 3520
rect 18875 3500 18885 3520
rect 18845 3470 18885 3500
rect 18845 3450 18855 3470
rect 18875 3450 18885 3470
rect 18845 3420 18885 3450
rect 18845 3400 18855 3420
rect 18875 3400 18885 3420
rect 18845 3370 18885 3400
rect 18845 3350 18855 3370
rect 18875 3350 18885 3370
rect 18845 3320 18885 3350
rect 18845 3300 18855 3320
rect 18875 3300 18885 3320
rect 18845 3270 18885 3300
rect 18845 3250 18855 3270
rect 18875 3250 18885 3270
rect 18845 3220 18885 3250
rect 18845 3200 18855 3220
rect 18875 3200 18885 3220
rect 18845 3170 18885 3200
rect 18845 3150 18855 3170
rect 18875 3150 18885 3170
rect 18845 3120 18885 3150
rect 18845 3100 18855 3120
rect 18875 3100 18885 3120
rect 18845 3070 18885 3100
rect 18845 3050 18855 3070
rect 18875 3050 18885 3070
rect 18845 3020 18885 3050
rect 18845 3000 18855 3020
rect 18875 3000 18885 3020
rect 18845 2985 18885 3000
rect 24965 3500 24975 3520
rect 24995 3500 25005 3520
rect 24965 3470 25005 3500
rect 24965 3450 24975 3470
rect 24995 3450 25005 3470
rect 24965 3420 25005 3450
rect 24965 3400 24975 3420
rect 24995 3400 25005 3420
rect 24965 3370 25005 3400
rect 24965 3350 24975 3370
rect 24995 3350 25005 3370
rect 24965 3320 25005 3350
rect 24965 3300 24975 3320
rect 24995 3300 25005 3320
rect 24965 3270 25005 3300
rect 24965 3250 24975 3270
rect 24995 3250 25005 3270
rect 24965 3220 25005 3250
rect 24965 3200 24975 3220
rect 24995 3200 25005 3220
rect 24965 3170 25005 3200
rect 24965 3150 24975 3170
rect 24995 3150 25005 3170
rect 24965 3120 25005 3150
rect 24965 3100 24975 3120
rect 24995 3100 25005 3120
rect 24965 3070 25005 3100
rect 24965 3050 24975 3070
rect 24995 3050 25005 3070
rect 24965 3020 25005 3050
rect 24965 3000 24975 3020
rect 24995 3000 25005 3020
rect 24965 2985 25005 3000
rect 25705 3570 25745 3585
rect 25705 3550 25715 3570
rect 25735 3550 25745 3570
rect 25705 3520 25745 3550
rect 25705 3500 25715 3520
rect 25735 3500 25745 3520
rect 25705 3470 25745 3500
rect 25705 3450 25715 3470
rect 25735 3450 25745 3470
rect 25705 3420 25745 3450
rect 25705 3400 25715 3420
rect 25735 3400 25745 3420
rect 25705 3370 25745 3400
rect 25705 3350 25715 3370
rect 25735 3350 25745 3370
rect 25705 3320 25745 3350
rect 25705 3300 25715 3320
rect 25735 3300 25745 3320
rect 25705 3270 25745 3300
rect 25705 3250 25715 3270
rect 25735 3250 25745 3270
rect 25705 3220 25745 3250
rect 25705 3200 25715 3220
rect 25735 3200 25745 3220
rect 25705 3170 25745 3200
rect 25705 3150 25715 3170
rect 25735 3150 25745 3170
rect 25705 3120 25745 3150
rect 25705 3100 25715 3120
rect 25735 3100 25745 3120
rect 26170 3445 26190 3680
rect 26170 3130 26190 3365
rect 27610 3445 27630 3680
rect 27610 3130 27630 3365
rect 26170 3110 26860 3130
rect 26940 3110 27630 3130
rect 28095 3410 28115 3740
rect 25705 3070 25745 3100
rect 25705 3050 25715 3070
rect 25735 3050 25745 3070
rect 25705 3020 25745 3050
rect 25705 3000 25715 3020
rect 25735 3000 25745 3020
rect 25705 2985 25745 3000
rect 28095 2990 28115 3315
rect 28875 3410 28895 3740
rect 28875 2990 28895 3315
rect 28095 2970 28455 2990
rect 28535 2970 28895 2990
rect 2955 2915 2995 2930
rect 2955 2895 2965 2915
rect 2985 2895 2995 2915
rect 2955 2865 2995 2895
rect 2955 2845 2965 2865
rect 2985 2845 2995 2865
rect 2955 2830 2995 2845
rect 5015 2915 5055 2930
rect 5015 2895 5025 2915
rect 5045 2895 5055 2915
rect 26985 2920 27375 2940
rect 27455 2920 27845 2940
rect 5015 2865 5055 2895
rect 5015 2845 5025 2865
rect 5045 2845 5055 2865
rect 5015 2830 5055 2845
rect 15975 2830 16015 2845
rect 15975 2810 15985 2830
rect 16005 2810 16015 2830
rect 15975 2780 16015 2810
rect 15975 2760 15985 2780
rect 16005 2760 16015 2780
rect 15975 2730 16015 2760
rect 15975 2710 15985 2730
rect 16005 2710 16015 2730
rect 3135 2685 3175 2700
rect 3135 2665 3145 2685
rect 3165 2665 3175 2685
rect 3135 2635 3175 2665
rect 3135 2615 3145 2635
rect 3165 2615 3175 2635
rect 3135 2585 3175 2615
rect 3135 2565 3145 2585
rect 3165 2565 3175 2585
rect 3135 2535 3175 2565
rect 3135 2515 3145 2535
rect 3165 2515 3175 2535
rect 3135 2485 3175 2515
rect 3135 2465 3145 2485
rect 3165 2465 3175 2485
rect 3135 2435 3175 2465
rect 3135 2415 3145 2435
rect 3165 2415 3175 2435
rect 3135 2400 3175 2415
rect 4835 2685 4875 2700
rect 4835 2665 4845 2685
rect 4865 2665 4875 2685
rect 15975 2680 16015 2710
rect 4835 2635 4875 2665
rect 15975 2660 15985 2680
rect 16005 2660 16015 2680
rect 4835 2615 4845 2635
rect 4865 2615 4875 2635
rect 14965 2640 15005 2655
rect 4835 2585 4875 2615
rect 4835 2565 4845 2585
rect 4865 2565 4875 2585
rect 4835 2535 4875 2565
rect 4835 2515 4845 2535
rect 4865 2515 4875 2535
rect 4835 2485 4875 2515
rect 4835 2465 4845 2485
rect 4865 2465 4875 2485
rect 4835 2435 4875 2465
rect 4835 2415 4845 2435
rect 4865 2415 4875 2435
rect 4835 2400 4875 2415
rect 14965 2620 14975 2640
rect 14995 2620 15005 2640
rect 14965 2590 15005 2620
rect 14965 2570 14975 2590
rect 14995 2570 15005 2590
rect 14965 2540 15005 2570
rect 14965 2520 14975 2540
rect 14995 2520 15005 2540
rect 14965 2490 15005 2520
rect 14965 2470 14975 2490
rect 14995 2470 15005 2490
rect 14965 2455 15005 2470
rect 15705 2640 15745 2655
rect 15705 2620 15715 2640
rect 15735 2620 15745 2640
rect 15705 2590 15745 2620
rect 15705 2570 15715 2590
rect 15735 2570 15745 2590
rect 15705 2540 15745 2570
rect 15705 2520 15715 2540
rect 15735 2520 15745 2540
rect 15705 2490 15745 2520
rect 15975 2630 16015 2660
rect 15975 2610 15985 2630
rect 16005 2610 16015 2630
rect 15975 2580 16015 2610
rect 15975 2560 15985 2580
rect 16005 2560 16015 2580
rect 15975 2530 16015 2560
rect 15975 2510 15985 2530
rect 16005 2510 16015 2530
rect 15975 2495 16015 2510
rect 16775 2830 16815 2845
rect 16775 2810 16785 2830
rect 16805 2810 16815 2830
rect 16775 2780 16815 2810
rect 16775 2760 16785 2780
rect 16805 2760 16815 2780
rect 16775 2730 16815 2760
rect 16775 2710 16785 2730
rect 16805 2710 16815 2730
rect 16775 2680 16815 2710
rect 16775 2660 16785 2680
rect 16805 2660 16815 2680
rect 16775 2630 16815 2660
rect 16775 2610 16785 2630
rect 16805 2610 16815 2630
rect 16775 2580 16815 2610
rect 16775 2560 16785 2580
rect 16805 2560 16815 2580
rect 16775 2530 16815 2560
rect 16775 2510 16785 2530
rect 16805 2510 16815 2530
rect 16775 2495 16815 2510
rect 16985 2830 17025 2845
rect 16985 2810 16995 2830
rect 17015 2810 17025 2830
rect 16985 2780 17025 2810
rect 16985 2760 16995 2780
rect 17015 2760 17025 2780
rect 16985 2730 17025 2760
rect 16985 2710 16995 2730
rect 17015 2710 17025 2730
rect 16985 2680 17025 2710
rect 16985 2660 16995 2680
rect 17015 2660 17025 2680
rect 16985 2630 17025 2660
rect 16985 2610 16995 2630
rect 17015 2610 17025 2630
rect 16985 2580 17025 2610
rect 16985 2560 16995 2580
rect 17015 2560 17025 2580
rect 16985 2530 17025 2560
rect 16985 2510 16995 2530
rect 17015 2510 17025 2530
rect 16985 2495 17025 2510
rect 17785 2830 17825 2845
rect 17785 2810 17795 2830
rect 17815 2810 17825 2830
rect 17785 2780 17825 2810
rect 17785 2760 17795 2780
rect 17815 2760 17825 2780
rect 17785 2730 17825 2760
rect 17785 2710 17795 2730
rect 17815 2710 17825 2730
rect 17785 2680 17825 2710
rect 17785 2660 17795 2680
rect 17815 2660 17825 2680
rect 25975 2830 26015 2845
rect 25975 2810 25985 2830
rect 26005 2810 26015 2830
rect 25975 2780 26015 2810
rect 25975 2760 25985 2780
rect 26005 2760 26015 2780
rect 25975 2730 26015 2760
rect 25975 2710 25985 2730
rect 26005 2710 26015 2730
rect 25975 2680 26015 2710
rect 17785 2630 17825 2660
rect 25975 2660 25985 2680
rect 26005 2660 26015 2680
rect 17785 2610 17795 2630
rect 17815 2610 17825 2630
rect 17785 2580 17825 2610
rect 17785 2560 17795 2580
rect 17815 2560 17825 2580
rect 17785 2530 17825 2560
rect 17785 2510 17795 2530
rect 17815 2510 17825 2530
rect 17785 2495 17825 2510
rect 18105 2640 18145 2655
rect 18105 2620 18115 2640
rect 18135 2620 18145 2640
rect 18105 2590 18145 2620
rect 18105 2570 18115 2590
rect 18135 2570 18145 2590
rect 18105 2540 18145 2570
rect 18105 2520 18115 2540
rect 18135 2520 18145 2540
rect 15705 2470 15715 2490
rect 15735 2470 15745 2490
rect 18105 2490 18145 2520
rect 18105 2470 18115 2490
rect 18135 2470 18145 2490
rect 15705 2455 15745 2470
rect 18105 2455 18145 2470
rect 18845 2640 18885 2655
rect 18845 2620 18855 2640
rect 18875 2620 18885 2640
rect 24965 2640 25005 2655
rect 18845 2590 18885 2620
rect 18845 2570 18855 2590
rect 18875 2570 18885 2590
rect 18845 2540 18885 2570
rect 18845 2520 18855 2540
rect 18875 2520 18885 2540
rect 18845 2490 18885 2520
rect 18845 2470 18855 2490
rect 18875 2470 18885 2490
rect 18845 2455 18885 2470
rect 3985 1985 4025 2000
rect 3985 1965 3995 1985
rect 4015 1965 4025 1985
rect 3985 1935 4025 1965
rect 3985 1915 3995 1935
rect 4015 1915 4025 1935
rect 3985 1900 4025 1915
rect 24965 2620 24975 2640
rect 24995 2620 25005 2640
rect 24965 2590 25005 2620
rect 24965 2570 24975 2590
rect 24995 2570 25005 2590
rect 24965 2540 25005 2570
rect 24965 2520 24975 2540
rect 24995 2520 25005 2540
rect 24965 2490 25005 2520
rect 24965 2470 24975 2490
rect 24995 2470 25005 2490
rect 24965 2455 25005 2470
rect 25705 2640 25745 2655
rect 25705 2620 25715 2640
rect 25735 2620 25745 2640
rect 25705 2590 25745 2620
rect 25705 2570 25715 2590
rect 25735 2570 25745 2590
rect 25705 2540 25745 2570
rect 25705 2520 25715 2540
rect 25735 2520 25745 2540
rect 25705 2490 25745 2520
rect 25975 2630 26015 2660
rect 25975 2610 25985 2630
rect 26005 2610 26015 2630
rect 25975 2580 26015 2610
rect 25975 2560 25985 2580
rect 26005 2560 26015 2580
rect 25975 2530 26015 2560
rect 25975 2510 25985 2530
rect 26005 2510 26015 2530
rect 25975 2495 26015 2510
rect 26775 2830 26815 2845
rect 26775 2810 26785 2830
rect 26805 2810 26815 2830
rect 26775 2780 26815 2810
rect 26775 2760 26785 2780
rect 26805 2760 26815 2780
rect 26775 2730 26815 2760
rect 26775 2710 26785 2730
rect 26805 2710 26815 2730
rect 26775 2680 26815 2710
rect 26775 2660 26785 2680
rect 26805 2660 26815 2680
rect 26775 2630 26815 2660
rect 26775 2610 26785 2630
rect 26805 2610 26815 2630
rect 26775 2580 26815 2610
rect 26775 2560 26785 2580
rect 26805 2560 26815 2580
rect 26775 2530 26815 2560
rect 26775 2510 26785 2530
rect 26805 2510 26815 2530
rect 26775 2495 26815 2510
rect 26985 2710 27005 2920
rect 25705 2470 25715 2490
rect 25735 2470 25745 2490
rect 25705 2455 25745 2470
rect 26985 2420 27005 2630
rect 27825 2710 27845 2920
rect 27825 2420 27845 2630
rect 26985 2400 27375 2420
rect 27455 2400 27845 2420
rect 28095 2780 28455 2800
rect 28535 2780 28895 2800
rect 28095 2645 28115 2780
rect 28095 2430 28115 2565
rect 28875 2645 28895 2780
rect 28875 2430 28895 2565
rect 28095 2410 28455 2430
rect 28535 2410 28895 2430
<< psubdiffcont >>
rect 29035 3280 29055 3375
rect 29295 3280 29315 3375
rect 29135 2960 29215 2980
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 14975 2230 14995 2250
rect 14975 2180 14995 2200
rect 14975 2130 14995 2150
rect 14975 2080 14995 2100
rect 14975 2030 14995 2050
rect 14975 1980 14995 2000
rect 15715 2230 15735 2250
rect 15715 2180 15735 2200
rect 18115 2230 18135 2250
rect 18115 2180 18135 2200
rect 15715 2130 15735 2150
rect 18115 2130 18135 2150
rect 15715 2080 15735 2100
rect 15715 2030 15735 2050
rect 15715 1980 15735 2000
rect 16245 2095 16265 2115
rect 16245 2045 16265 2065
rect 16245 1995 16265 2015
rect 17535 2095 17555 2115
rect 17535 2045 17555 2065
rect 17535 1995 17555 2015
rect 18115 2080 18135 2100
rect 18115 2030 18135 2050
rect 18115 1980 18135 2000
rect 18855 2230 18875 2250
rect 18855 2180 18875 2200
rect 18855 2130 18875 2150
rect 18855 2080 18875 2100
rect 18855 2030 18875 2050
rect 29135 2665 29215 2685
rect 28455 2320 28535 2340
rect 24975 2230 24995 2250
rect 24975 2180 24995 2200
rect 24975 2130 24995 2150
rect 24975 2080 24995 2100
rect 24975 2030 24995 2050
rect 18855 1980 18875 2000
rect 24975 1980 24995 2000
rect 25715 2230 25735 2250
rect 25715 2180 25735 2200
rect 25715 2130 25735 2150
rect 25715 2080 25735 2100
rect 25715 2030 25735 2050
rect 25715 1980 25735 2000
rect 26860 2205 26940 2225
rect 26225 2010 26245 2090
rect 27555 2010 27575 2090
rect 26860 1885 26940 1905
rect 28095 2055 28115 2135
rect 28875 2055 28895 2135
rect 28995 2255 29015 2335
rect 29330 2255 29350 2335
rect 29135 1905 29215 1925
rect 28455 1850 28535 1870
rect 26860 1800 26940 1820
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 3995 1630 4015 1650
rect 14975 1620 14995 1640
rect 5075 1040 5095 1060
rect 5075 990 5095 1010
rect 14975 1570 14995 1590
rect 14975 1520 14995 1540
rect 14975 1470 14995 1490
rect 14975 1420 14995 1440
rect 14975 1370 14995 1390
rect 14975 1320 14995 1340
rect 14975 1270 14995 1290
rect 14975 1220 14995 1240
rect 14975 1170 14995 1190
rect 14975 1120 14995 1140
rect 14975 1070 14995 1090
rect 14975 1020 14995 1040
rect 14975 970 14995 990
rect 15655 1620 15675 1640
rect 15655 1570 15675 1590
rect 15655 1520 15675 1540
rect 16000 1630 16020 1650
rect 16000 1580 16020 1600
rect 16000 1530 16020 1550
rect 16740 1630 16760 1650
rect 16740 1580 16760 1600
rect 16740 1530 16760 1550
rect 17040 1630 17060 1650
rect 17040 1580 17060 1600
rect 17040 1530 17060 1550
rect 17780 1630 17800 1650
rect 17780 1580 17800 1600
rect 17780 1530 17800 1550
rect 18175 1620 18195 1640
rect 18175 1570 18195 1590
rect 18175 1520 18195 1540
rect 15655 1470 15675 1490
rect 18175 1470 18195 1490
rect 15655 1420 15675 1440
rect 15655 1370 15675 1390
rect 15655 1320 15675 1340
rect 15655 1270 15675 1290
rect 18175 1420 18195 1440
rect 18175 1370 18195 1390
rect 18175 1320 18195 1340
rect 18175 1270 18195 1290
rect 15655 1220 15675 1240
rect 15655 1170 15675 1190
rect 18175 1220 18195 1240
rect 15655 1120 15675 1140
rect 15655 1070 15675 1090
rect 15655 1020 15675 1040
rect 15655 970 15675 990
rect 16175 1150 16195 1170
rect 16175 1100 16195 1120
rect 16175 1050 16195 1070
rect 16175 1000 16195 1020
rect 16175 950 16195 970
rect 17630 1150 17650 1170
rect 17630 1100 17650 1120
rect 17630 1050 17650 1070
rect 17630 1000 17650 1020
rect 17630 950 17650 970
rect 18175 1170 18195 1190
rect 18175 1120 18195 1140
rect 18175 1070 18195 1090
rect 18175 1020 18195 1040
rect 18175 970 18195 990
rect 18855 1620 18875 1640
rect 24975 1620 24995 1640
rect 18855 1570 18875 1590
rect 18855 1520 18875 1540
rect 18855 1470 18875 1490
rect 18855 1420 18875 1440
rect 18855 1370 18875 1390
rect 18855 1320 18875 1340
rect 18855 1270 18875 1290
rect 18855 1220 18875 1240
rect 18855 1170 18875 1190
rect 18855 1120 18875 1140
rect 18855 1070 18875 1090
rect 18855 1020 18875 1040
rect 18855 970 18875 990
rect 24975 1570 24995 1590
rect 24975 1520 24995 1540
rect 24975 1470 24995 1490
rect 24975 1420 24995 1440
rect 24975 1370 24995 1390
rect 24975 1320 24995 1340
rect 24975 1270 24995 1290
rect 24975 1220 24995 1240
rect 24975 1170 24995 1190
rect 24975 1120 24995 1140
rect 24975 1070 24995 1090
rect 24975 1020 24995 1040
rect 24975 970 24995 990
rect 25655 1620 25675 1640
rect 25655 1570 25675 1590
rect 25655 1520 25675 1540
rect 25655 1470 25675 1490
rect 25655 1420 25675 1440
rect 25655 1370 25675 1390
rect 25940 1550 25960 1630
rect 26740 1630 26760 1650
rect 26740 1580 26760 1600
rect 26740 1530 26760 1550
rect 27040 1630 27060 1650
rect 27040 1580 27060 1600
rect 27040 1530 27060 1550
rect 27840 1550 27860 1630
rect 26860 1360 26940 1380
rect 28485 1730 28565 1750
rect 25655 1320 25675 1340
rect 25655 1270 25675 1290
rect 25655 1220 25675 1240
rect 28155 1265 28175 1345
rect 25655 1170 25675 1190
rect 25655 1120 25675 1140
rect 25655 1070 25675 1090
rect 25655 1020 25675 1040
rect 25655 970 25675 990
rect 26845 1175 26925 1195
rect 26155 900 26175 980
rect 2965 845 2985 865
rect 2965 795 2985 815
rect 5025 845 5045 865
rect 5025 795 5045 815
rect 27655 900 27675 980
rect 28875 1265 28895 1345
rect 28485 860 28565 880
rect 29065 1675 29145 1695
rect 28985 1220 29005 1300
rect 29200 1220 29220 1300
rect 29065 840 29145 860
rect 16850 715 16870 735
rect 26845 735 26925 755
rect 17590 715 17610 735
rect 26355 625 26435 645
rect 26210 475 26230 555
rect 26565 475 26585 555
rect 26355 395 26435 415
rect 27190 625 27270 645
rect 26830 475 26850 555
rect 27610 475 27630 555
rect 27190 405 27270 425
<< nsubdiffcont >>
rect 26520 4950 26600 4970
rect 26205 4785 26225 4865
rect 26935 4785 26955 4865
rect 26520 4695 26600 4715
rect 27460 4925 27540 4945
rect 27185 4780 27205 4860
rect 27785 4780 27805 4865
rect 27460 4695 27540 4715
rect 26835 4505 26915 4525
rect 16175 4305 16195 4325
rect 16435 4305 16455 4325
rect 16505 4320 16525 4340
rect 26200 4365 26220 4445
rect 16945 4320 16965 4340
rect 17155 4305 17175 4325
rect 17715 4305 17735 4325
rect 27530 4365 27550 4445
rect 26835 4285 26915 4305
rect 16220 4070 16240 4090
rect 17510 4070 17530 4090
rect 26875 4095 26955 4115
rect 26150 3955 26170 4035
rect 27660 3955 27680 4035
rect 26875 3875 26955 3895
rect 16165 3765 16185 3785
rect 16905 3765 16925 3785
rect 17645 3765 17665 3785
rect 28455 3740 28535 3760
rect 26860 3680 26940 3700
rect 14975 3550 14995 3570
rect 14975 3500 14995 3520
rect 14975 3450 14995 3470
rect 14975 3400 14995 3420
rect 14975 3350 14995 3370
rect 14975 3300 14995 3320
rect 14975 3250 14995 3270
rect 14975 3200 14995 3220
rect 14975 3150 14995 3170
rect 14975 3100 14995 3120
rect 14975 3050 14995 3070
rect 14975 3000 14995 3020
rect 15715 3550 15735 3570
rect 18115 3550 18135 3570
rect 15715 3500 15735 3520
rect 15715 3450 15735 3470
rect 15715 3400 15735 3420
rect 15715 3350 15735 3370
rect 15715 3300 15735 3320
rect 15715 3250 15735 3270
rect 15715 3200 15735 3220
rect 15715 3150 15735 3170
rect 16190 3490 16210 3510
rect 16190 3440 16210 3460
rect 16190 3390 16210 3410
rect 16190 3340 16210 3360
rect 16190 3290 16210 3310
rect 16190 3240 16210 3260
rect 16190 3190 16210 3210
rect 16190 3140 16210 3160
rect 17590 3490 17610 3510
rect 17590 3440 17610 3460
rect 17590 3390 17610 3410
rect 17590 3340 17610 3360
rect 17590 3290 17610 3310
rect 17590 3240 17610 3260
rect 17590 3190 17610 3210
rect 17590 3140 17610 3160
rect 18115 3500 18135 3520
rect 18115 3450 18135 3470
rect 18115 3400 18135 3420
rect 18115 3350 18135 3370
rect 18115 3300 18135 3320
rect 18115 3250 18135 3270
rect 18115 3200 18135 3220
rect 18115 3150 18135 3170
rect 15715 3100 15735 3120
rect 18115 3100 18135 3120
rect 15715 3050 15735 3070
rect 15715 3000 15735 3020
rect 18115 3050 18135 3070
rect 18115 3000 18135 3020
rect 18855 3550 18875 3570
rect 24975 3550 24995 3570
rect 18855 3500 18875 3520
rect 18855 3450 18875 3470
rect 18855 3400 18875 3420
rect 18855 3350 18875 3370
rect 18855 3300 18875 3320
rect 18855 3250 18875 3270
rect 18855 3200 18875 3220
rect 18855 3150 18875 3170
rect 18855 3100 18875 3120
rect 18855 3050 18875 3070
rect 18855 3000 18875 3020
rect 24975 3500 24995 3520
rect 24975 3450 24995 3470
rect 24975 3400 24995 3420
rect 24975 3350 24995 3370
rect 24975 3300 24995 3320
rect 24975 3250 24995 3270
rect 24975 3200 24995 3220
rect 24975 3150 24995 3170
rect 24975 3100 24995 3120
rect 24975 3050 24995 3070
rect 24975 3000 24995 3020
rect 25715 3550 25735 3570
rect 25715 3500 25735 3520
rect 25715 3450 25735 3470
rect 25715 3400 25735 3420
rect 25715 3350 25735 3370
rect 25715 3300 25735 3320
rect 25715 3250 25735 3270
rect 25715 3200 25735 3220
rect 25715 3150 25735 3170
rect 25715 3100 25735 3120
rect 26170 3365 26190 3445
rect 27610 3365 27630 3445
rect 26860 3110 26940 3130
rect 28095 3315 28115 3410
rect 25715 3050 25735 3070
rect 25715 3000 25735 3020
rect 28875 3315 28895 3410
rect 28455 2970 28535 2990
rect 2965 2895 2985 2915
rect 2965 2845 2985 2865
rect 5025 2895 5045 2915
rect 27375 2920 27455 2940
rect 5025 2845 5045 2865
rect 15985 2810 16005 2830
rect 15985 2760 16005 2780
rect 15985 2710 16005 2730
rect 3145 2665 3165 2685
rect 3145 2615 3165 2635
rect 3145 2565 3165 2585
rect 3145 2515 3165 2535
rect 3145 2465 3165 2485
rect 3145 2415 3165 2435
rect 4845 2665 4865 2685
rect 15985 2660 16005 2680
rect 4845 2615 4865 2635
rect 4845 2565 4865 2585
rect 4845 2515 4865 2535
rect 4845 2465 4865 2485
rect 4845 2415 4865 2435
rect 14975 2620 14995 2640
rect 14975 2570 14995 2590
rect 14975 2520 14995 2540
rect 14975 2470 14995 2490
rect 15715 2620 15735 2640
rect 15715 2570 15735 2590
rect 15715 2520 15735 2540
rect 15985 2610 16005 2630
rect 15985 2560 16005 2580
rect 15985 2510 16005 2530
rect 16785 2810 16805 2830
rect 16785 2760 16805 2780
rect 16785 2710 16805 2730
rect 16785 2660 16805 2680
rect 16785 2610 16805 2630
rect 16785 2560 16805 2580
rect 16785 2510 16805 2530
rect 16995 2810 17015 2830
rect 16995 2760 17015 2780
rect 16995 2710 17015 2730
rect 16995 2660 17015 2680
rect 16995 2610 17015 2630
rect 16995 2560 17015 2580
rect 16995 2510 17015 2530
rect 17795 2810 17815 2830
rect 17795 2760 17815 2780
rect 17795 2710 17815 2730
rect 17795 2660 17815 2680
rect 25985 2810 26005 2830
rect 25985 2760 26005 2780
rect 25985 2710 26005 2730
rect 25985 2660 26005 2680
rect 17795 2610 17815 2630
rect 17795 2560 17815 2580
rect 17795 2510 17815 2530
rect 18115 2620 18135 2640
rect 18115 2570 18135 2590
rect 18115 2520 18135 2540
rect 15715 2470 15735 2490
rect 18115 2470 18135 2490
rect 18855 2620 18875 2640
rect 18855 2570 18875 2590
rect 18855 2520 18875 2540
rect 18855 2470 18875 2490
rect 3995 1965 4015 1985
rect 3995 1915 4015 1935
rect 24975 2620 24995 2640
rect 24975 2570 24995 2590
rect 24975 2520 24995 2540
rect 24975 2470 24995 2490
rect 25715 2620 25735 2640
rect 25715 2570 25735 2590
rect 25715 2520 25735 2540
rect 25985 2610 26005 2630
rect 25985 2560 26005 2580
rect 25985 2510 26005 2530
rect 26785 2810 26805 2830
rect 26785 2760 26805 2780
rect 26785 2710 26805 2730
rect 26785 2660 26805 2680
rect 26785 2610 26805 2630
rect 26785 2560 26805 2580
rect 26785 2510 26805 2530
rect 26985 2630 27005 2710
rect 25715 2470 25735 2490
rect 27825 2630 27845 2710
rect 27375 2400 27455 2420
rect 28455 2780 28535 2800
rect 28095 2565 28115 2645
rect 28875 2565 28895 2645
rect 28455 2410 28535 2430
<< poly >>
rect 26865 4920 26905 4930
rect 26865 4905 26875 4920
rect 26845 4900 26875 4905
rect 26895 4900 26905 4920
rect 26845 4890 26905 4900
rect 26545 4875 26565 4890
rect 26605 4875 26625 4890
rect 26665 4875 26685 4890
rect 26725 4875 26745 4890
rect 26785 4875 26805 4890
rect 26845 4875 26865 4890
rect 26295 4858 26315 4875
rect 26355 4858 26375 4873
rect 26415 4858 26435 4873
rect 26295 4780 26315 4795
rect 26355 4780 26375 4795
rect 26415 4780 26435 4795
rect 26545 4780 26565 4795
rect 26605 4785 26625 4795
rect 26665 4785 26685 4795
rect 26725 4785 26745 4795
rect 26785 4785 26805 4795
rect 26345 4770 26385 4780
rect 26605 4770 26805 4785
rect 26845 4780 26865 4795
rect 26345 4750 26355 4770
rect 26375 4750 26385 4770
rect 26345 4740 26385 4750
rect 26685 4765 26725 4770
rect 26685 4745 26695 4765
rect 26715 4745 26725 4765
rect 26685 4735 26725 4745
rect 27275 4850 27295 4865
rect 27335 4850 27355 4865
rect 27395 4850 27415 4865
rect 27455 4850 27475 4865
rect 27515 4850 27535 4865
rect 27575 4850 27595 4865
rect 27635 4850 27655 4865
rect 27695 4850 27715 4865
rect 27275 4780 27295 4790
rect 27335 4780 27355 4790
rect 27395 4780 27415 4790
rect 27455 4780 27475 4790
rect 27515 4780 27535 4790
rect 27575 4780 27595 4790
rect 27635 4780 27655 4790
rect 27695 4780 27715 4790
rect 27275 4765 27715 4780
rect 27358 4745 27366 4765
rect 27384 4745 27392 4765
rect 27358 4735 27392 4745
rect 16597 4460 16633 4470
rect 16597 4440 16605 4460
rect 16625 4440 16633 4460
rect 16597 4430 16633 4440
rect 16717 4460 16753 4470
rect 16717 4440 16725 4460
rect 16745 4440 16753 4460
rect 16717 4430 16753 4440
rect 16837 4460 16873 4470
rect 16837 4440 16845 4460
rect 16865 4440 16873 4460
rect 16837 4430 16873 4440
rect 16535 4415 16575 4425
rect 16165 4400 16205 4410
rect 16165 4380 16175 4400
rect 16195 4380 16205 4400
rect 16425 4400 16465 4410
rect 16425 4380 16435 4400
rect 16455 4380 16465 4400
rect 16535 4395 16545 4415
rect 16565 4400 16575 4415
rect 16895 4415 16935 4425
rect 16895 4400 16905 4415
rect 16565 4395 16595 4400
rect 16535 4385 16595 4395
rect 16875 4395 16905 4400
rect 16925 4395 16935 4415
rect 16875 4385 16935 4395
rect 16165 4365 16265 4380
rect 16245 4353 16265 4365
rect 16305 4353 16325 4368
rect 16365 4365 16465 4380
rect 16575 4370 16595 4385
rect 16635 4370 16655 4385
rect 16695 4370 16715 4385
rect 16755 4370 16775 4385
rect 16815 4370 16835 4385
rect 16875 4370 16895 4385
rect 16365 4353 16385 4365
rect 26290 4430 26305 4445
rect 26345 4430 26360 4445
rect 26400 4430 26415 4445
rect 26455 4430 26470 4445
rect 26510 4430 26525 4445
rect 26565 4430 26580 4445
rect 26620 4430 26635 4445
rect 26675 4430 26690 4445
rect 26730 4430 26745 4445
rect 26785 4430 26800 4445
rect 26840 4430 26855 4445
rect 26895 4430 26910 4445
rect 26950 4430 26965 4445
rect 27005 4430 27020 4445
rect 27060 4430 27075 4445
rect 27115 4430 27130 4445
rect 27170 4430 27185 4445
rect 27225 4430 27240 4445
rect 27280 4430 27295 4445
rect 27335 4430 27350 4445
rect 27390 4430 27405 4445
rect 27445 4430 27460 4445
rect 26290 4365 26305 4380
rect 26345 4370 26360 4380
rect 26400 4370 26415 4380
rect 26455 4370 26470 4380
rect 26510 4370 26525 4380
rect 26565 4370 26580 4380
rect 26620 4370 26635 4380
rect 26675 4370 26690 4380
rect 26730 4370 26745 4380
rect 26785 4370 26800 4380
rect 26840 4370 26855 4380
rect 26895 4370 26910 4380
rect 26950 4370 26965 4380
rect 27005 4370 27020 4380
rect 27060 4370 27075 4380
rect 27115 4370 27130 4380
rect 27170 4370 27185 4380
rect 27225 4370 27240 4380
rect 27280 4370 27295 4380
rect 27335 4370 27350 4380
rect 27390 4370 27405 4380
rect 17225 4345 17245 4360
rect 17285 4345 17305 4360
rect 17345 4345 17365 4360
rect 17405 4345 17425 4360
rect 17465 4345 17485 4360
rect 17525 4345 17545 4360
rect 17585 4345 17605 4360
rect 17645 4345 17665 4360
rect 16245 4275 16265 4290
rect 16305 4275 16325 4290
rect 16365 4275 16385 4290
rect 16575 4275 16595 4290
rect 16635 4280 16655 4290
rect 16695 4280 16715 4290
rect 16755 4280 16775 4290
rect 16815 4280 16835 4290
rect 16295 4265 16335 4275
rect 16635 4265 16835 4280
rect 16875 4275 16895 4290
rect 26345 4355 27405 4370
rect 27445 4365 27460 4380
rect 26362 4335 26370 4355
rect 26390 4335 26398 4355
rect 26362 4325 26398 4335
rect 17225 4275 17245 4285
rect 17285 4275 17305 4285
rect 17345 4275 17365 4285
rect 17405 4275 17425 4285
rect 17465 4275 17485 4285
rect 17525 4275 17545 4285
rect 17585 4275 17605 4285
rect 17645 4275 17665 4285
rect 16295 4245 16305 4265
rect 16325 4245 16335 4265
rect 16295 4235 16335 4245
rect 16715 4260 16755 4265
rect 17225 4260 17665 4275
rect 16715 4240 16725 4260
rect 16745 4240 16755 4260
rect 16715 4230 16755 4240
rect 17308 4240 17316 4260
rect 17334 4240 17342 4260
rect 17308 4230 17342 4240
rect 16210 4150 16250 4160
rect 16210 4130 16220 4150
rect 16240 4130 16250 4150
rect 17500 4150 17540 4160
rect 17500 4130 17510 4150
rect 17530 4130 17540 4150
rect 16210 4115 16305 4130
rect 16290 4105 16305 4115
rect 16345 4105 16360 4120
rect 16400 4105 16415 4120
rect 16455 4105 16470 4120
rect 16510 4105 16525 4120
rect 16565 4105 16580 4120
rect 16620 4105 16635 4120
rect 16675 4105 16690 4120
rect 16730 4105 16745 4120
rect 16785 4105 16800 4120
rect 16840 4105 16855 4120
rect 16895 4105 16910 4120
rect 16950 4105 16965 4120
rect 17005 4105 17020 4120
rect 17060 4105 17075 4120
rect 17115 4105 17130 4120
rect 17170 4105 17185 4120
rect 17225 4105 17240 4120
rect 17280 4105 17295 4120
rect 17335 4105 17350 4120
rect 17390 4105 17405 4120
rect 17445 4115 17540 4130
rect 17445 4105 17460 4115
rect 16290 4040 16305 4055
rect 16345 4045 16360 4055
rect 16400 4045 16415 4055
rect 16455 4045 16470 4055
rect 16510 4045 16525 4055
rect 16565 4045 16580 4055
rect 16620 4045 16635 4055
rect 16675 4045 16690 4055
rect 16730 4045 16745 4055
rect 16785 4045 16800 4055
rect 16840 4045 16855 4055
rect 16895 4045 16910 4055
rect 16950 4045 16965 4055
rect 17005 4045 17020 4055
rect 17060 4045 17075 4055
rect 17115 4045 17130 4055
rect 17170 4045 17185 4055
rect 17225 4045 17240 4055
rect 17280 4045 17295 4055
rect 17335 4045 17350 4055
rect 17390 4045 17405 4055
rect 16345 4030 17405 4045
rect 17445 4040 17460 4055
rect 26280 4065 26310 4075
rect 26280 4045 26285 4065
rect 26305 4045 26310 4065
rect 26480 4065 26510 4075
rect 26480 4045 26485 4065
rect 26505 4045 26510 4065
rect 27008 4065 27038 4075
rect 27008 4045 27013 4065
rect 27033 4045 27038 4065
rect 27205 4065 27245 4075
rect 27205 4045 27215 4065
rect 27235 4045 27245 4065
rect 27425 4065 27465 4075
rect 27425 4045 27435 4065
rect 27455 4045 27465 4065
rect 26280 4035 26310 4045
rect 16362 4010 16370 4030
rect 16390 4010 16398 4030
rect 16362 4000 16398 4010
rect 26240 4020 26255 4035
rect 26295 4020 26310 4035
rect 26350 4020 26365 4035
rect 26405 4020 26420 4035
rect 26460 4030 26530 4045
rect 26460 4020 26475 4030
rect 26515 4020 26530 4030
rect 26570 4020 26585 4035
rect 26625 4020 26640 4035
rect 26680 4030 26750 4045
rect 27008 4035 27040 4045
rect 26680 4020 26695 4030
rect 26735 4020 26750 4030
rect 26790 4020 26805 4035
rect 26845 4020 26860 4035
rect 26970 4020 26985 4035
rect 27025 4020 27040 4035
rect 27080 4020 27095 4035
rect 27135 4020 27150 4035
rect 27190 4030 27260 4045
rect 27190 4020 27205 4030
rect 27245 4020 27260 4030
rect 27300 4020 27315 4035
rect 27355 4020 27370 4035
rect 27410 4030 27480 4045
rect 27410 4020 27425 4030
rect 27465 4020 27480 4030
rect 27520 4020 27535 4035
rect 27575 4020 27590 4035
rect 26240 3955 26255 3970
rect 26295 3955 26310 3970
rect 26350 3960 26365 3970
rect 26405 3960 26420 3970
rect 26350 3955 26420 3960
rect 26460 3955 26475 3970
rect 26515 3955 26530 3970
rect 26570 3960 26585 3970
rect 26625 3960 26640 3970
rect 26570 3955 26640 3960
rect 26680 3955 26695 3970
rect 26735 3955 26750 3970
rect 26790 3955 26805 3970
rect 26845 3955 26860 3970
rect 26970 3955 26985 3970
rect 27025 3955 27040 3970
rect 27080 3960 27095 3970
rect 27135 3960 27150 3970
rect 27080 3955 27150 3960
rect 27190 3955 27205 3970
rect 27245 3955 27260 3970
rect 27300 3960 27315 3970
rect 27355 3960 27370 3970
rect 27300 3955 27370 3960
rect 27410 3955 27425 3970
rect 27465 3955 27480 3970
rect 27520 3955 27535 3970
rect 27575 3955 27590 3970
rect 26350 3945 26439 3955
rect 26570 3945 26659 3955
rect 26407 3925 26413 3945
rect 26430 3925 26439 3945
rect 26407 3915 26439 3925
rect 26627 3925 26633 3945
rect 26650 3925 26659 3945
rect 26627 3915 26659 3925
rect 26771 3945 26805 3955
rect 27080 3945 27169 3955
rect 27300 3945 27389 3955
rect 26771 3925 26780 3945
rect 26797 3925 26805 3945
rect 26771 3915 26805 3925
rect 27137 3925 27143 3945
rect 27160 3925 27169 3945
rect 27137 3915 27169 3925
rect 27357 3925 27363 3945
rect 27380 3925 27389 3945
rect 27357 3915 27389 3925
rect 27501 3945 27535 3955
rect 27501 3925 27510 3945
rect 27527 3925 27535 3945
rect 27501 3915 27535 3925
rect 16155 3845 16195 3855
rect 16155 3825 16165 3845
rect 16185 3825 16195 3845
rect 16271 3845 16303 3855
rect 16271 3825 16277 3845
rect 16294 3825 16303 3845
rect 16470 3845 16510 3855
rect 16470 3825 16480 3845
rect 16500 3825 16510 3845
rect 16690 3845 16730 3855
rect 16690 3825 16700 3845
rect 16720 3825 16730 3845
rect 16895 3845 16935 3855
rect 16895 3825 16905 3845
rect 16925 3825 16935 3845
rect 17011 3845 17043 3855
rect 17011 3825 17017 3845
rect 17034 3825 17043 3845
rect 17210 3845 17250 3855
rect 17210 3825 17220 3845
rect 17240 3825 17250 3845
rect 17430 3845 17470 3855
rect 17430 3825 17440 3845
rect 17460 3825 17470 3845
rect 17635 3845 17675 3855
rect 17635 3825 17645 3845
rect 17665 3825 17675 3845
rect 16155 3810 16250 3825
rect 16271 3815 16305 3825
rect 16235 3800 16250 3810
rect 16290 3800 16305 3815
rect 16345 3800 16360 3815
rect 16400 3800 16415 3815
rect 16455 3810 16525 3825
rect 16455 3800 16470 3810
rect 16510 3800 16525 3810
rect 16565 3800 16580 3815
rect 16620 3800 16635 3815
rect 16675 3810 16745 3825
rect 16675 3800 16690 3810
rect 16730 3800 16745 3810
rect 16785 3800 16800 3815
rect 16840 3810 16990 3825
rect 17011 3815 17045 3825
rect 16840 3800 16855 3810
rect 16975 3800 16990 3810
rect 17030 3800 17045 3815
rect 17085 3800 17100 3815
rect 17140 3800 17155 3815
rect 17195 3810 17265 3825
rect 17195 3800 17210 3810
rect 17250 3800 17265 3810
rect 17305 3800 17320 3815
rect 17360 3800 17375 3815
rect 17415 3810 17485 3825
rect 17415 3800 17430 3810
rect 17470 3800 17485 3810
rect 17525 3800 17540 3815
rect 17580 3810 17675 3825
rect 17580 3800 17595 3810
rect 16235 3735 16250 3750
rect 16290 3735 16305 3750
rect 16345 3740 16360 3750
rect 16400 3740 16415 3750
rect 16345 3735 16415 3740
rect 16455 3735 16470 3750
rect 16510 3735 16525 3750
rect 16565 3740 16580 3750
rect 16620 3740 16635 3750
rect 16565 3735 16635 3740
rect 16675 3735 16690 3750
rect 16730 3735 16745 3750
rect 16785 3735 16800 3750
rect 16840 3735 16855 3750
rect 16975 3735 16990 3750
rect 17030 3735 17045 3750
rect 17085 3740 17100 3750
rect 17140 3740 17155 3750
rect 17085 3735 17155 3740
rect 17195 3735 17210 3750
rect 17250 3735 17265 3750
rect 17305 3740 17320 3750
rect 17360 3740 17375 3750
rect 17305 3735 17375 3740
rect 17415 3735 17430 3750
rect 17470 3735 17485 3750
rect 17525 3735 17540 3750
rect 17580 3735 17595 3750
rect 16345 3725 16434 3735
rect 16565 3725 16654 3735
rect 16402 3705 16408 3725
rect 16425 3705 16434 3725
rect 16402 3695 16434 3705
rect 16622 3705 16628 3725
rect 16645 3705 16654 3725
rect 16622 3695 16654 3705
rect 16766 3725 16800 3735
rect 17085 3725 17174 3735
rect 17305 3725 17394 3735
rect 16766 3705 16775 3725
rect 16792 3705 16800 3725
rect 16766 3695 16800 3705
rect 17142 3705 17148 3725
rect 17165 3705 17174 3725
rect 17142 3695 17174 3705
rect 17362 3705 17368 3725
rect 17385 3705 17394 3725
rect 17362 3695 17394 3705
rect 17506 3725 17540 3735
rect 17506 3705 17515 3725
rect 17532 3705 17540 3725
rect 17506 3695 17540 3705
rect 15045 3585 15060 3600
rect 15100 3585 15115 3600
rect 15155 3585 15170 3600
rect 15210 3585 15225 3600
rect 15265 3585 15280 3600
rect 15320 3585 15335 3600
rect 15375 3585 15390 3600
rect 15430 3585 15445 3600
rect 15485 3585 15500 3600
rect 15540 3585 15555 3600
rect 15595 3585 15610 3600
rect 15650 3585 15665 3600
rect 18185 3585 18200 3600
rect 18240 3585 18255 3600
rect 18295 3585 18310 3600
rect 18350 3585 18365 3600
rect 18405 3585 18420 3600
rect 18460 3585 18475 3600
rect 18515 3585 18530 3600
rect 18570 3585 18585 3600
rect 18625 3585 18640 3600
rect 18680 3585 18695 3600
rect 18735 3585 18750 3600
rect 18790 3585 18805 3600
rect 25045 3585 25060 3600
rect 25100 3585 25115 3600
rect 25155 3585 25170 3600
rect 25210 3585 25225 3600
rect 25265 3585 25280 3600
rect 25320 3585 25335 3600
rect 25375 3585 25390 3600
rect 25430 3585 25445 3600
rect 25485 3585 25500 3600
rect 25540 3585 25555 3600
rect 25595 3585 25610 3600
rect 25650 3585 25665 3600
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 3035 2930 3085 2945
rect 3125 2930 3175 2945
rect 3215 2930 3265 2945
rect 3305 2930 3355 2945
rect 3395 2930 3445 2945
rect 3485 2930 3535 2945
rect 3575 2930 3625 2945
rect 3665 2930 3715 2945
rect 3755 2930 3805 2945
rect 3845 2930 3895 2945
rect 3935 2930 3985 2945
rect 4025 2930 4075 2945
rect 4115 2930 4165 2945
rect 4205 2930 4255 2945
rect 4295 2930 4345 2945
rect 4385 2930 4435 2945
rect 4475 2930 4525 2945
rect 4565 2930 4615 2945
rect 4655 2930 4705 2945
rect 4745 2930 4795 2945
rect 4835 2930 4885 2945
rect 4925 2930 4975 2945
rect 16180 3570 16220 3580
rect 16180 3550 16190 3570
rect 16210 3550 16220 3570
rect 17580 3570 17620 3580
rect 17580 3550 17590 3570
rect 17610 3550 17620 3570
rect 16180 3535 16280 3550
rect 16260 3525 16280 3535
rect 16320 3525 16340 3540
rect 16380 3525 16400 3540
rect 16440 3525 16460 3540
rect 16500 3525 16520 3540
rect 16560 3525 16580 3540
rect 16620 3525 16640 3540
rect 16680 3525 16700 3540
rect 16740 3525 16760 3540
rect 16800 3525 16820 3540
rect 16860 3525 16880 3540
rect 16920 3525 16940 3540
rect 16980 3525 17000 3540
rect 17040 3525 17060 3540
rect 17100 3525 17120 3540
rect 17160 3525 17180 3540
rect 17220 3525 17240 3540
rect 17280 3525 17300 3540
rect 17340 3525 17360 3540
rect 17400 3525 17420 3540
rect 17460 3525 17480 3540
rect 17520 3535 17620 3550
rect 17520 3525 17540 3535
rect 16260 3110 16280 3125
rect 16320 3115 16340 3125
rect 16380 3115 16400 3125
rect 16440 3115 16460 3125
rect 16500 3115 16520 3125
rect 16560 3115 16580 3125
rect 16620 3115 16640 3125
rect 16680 3115 16700 3125
rect 16740 3115 16760 3125
rect 16800 3115 16820 3125
rect 16860 3115 16880 3125
rect 16920 3115 16940 3125
rect 16980 3115 17000 3125
rect 17040 3115 17060 3125
rect 17100 3115 17120 3125
rect 17160 3115 17180 3125
rect 17220 3115 17240 3125
rect 17280 3115 17300 3125
rect 17340 3115 17360 3125
rect 17400 3115 17420 3125
rect 17460 3115 17480 3125
rect 16320 3100 17480 3115
rect 17520 3110 17540 3125
rect 16823 3080 16831 3100
rect 16849 3080 16857 3100
rect 16823 3070 16857 3080
rect 15045 2975 15060 2985
rect 14965 2960 15060 2975
rect 15100 2975 15115 2985
rect 15155 2975 15170 2985
rect 15210 2975 15225 2985
rect 15265 2975 15280 2985
rect 15320 2975 15335 2985
rect 15375 2975 15390 2985
rect 15430 2975 15445 2985
rect 15485 2975 15500 2985
rect 15540 2975 15555 2985
rect 15595 2975 15610 2985
rect 15100 2960 15610 2975
rect 15650 2975 15665 2985
rect 18185 2975 18200 2985
rect 15650 2960 15745 2975
rect 14965 2940 14975 2960
rect 14995 2940 15005 2960
rect 14965 2930 15005 2940
rect 15503 2940 15511 2960
rect 15529 2940 15537 2960
rect 15503 2930 15537 2940
rect 15705 2940 15715 2960
rect 15735 2940 15745 2960
rect 15705 2930 15745 2940
rect 18105 2960 18200 2975
rect 18240 2975 18255 2985
rect 18295 2975 18310 2985
rect 18350 2975 18365 2985
rect 18405 2975 18420 2985
rect 18460 2975 18475 2985
rect 18515 2975 18530 2985
rect 18570 2975 18585 2985
rect 18625 2975 18640 2985
rect 18680 2975 18695 2985
rect 18735 2975 18750 2985
rect 18240 2960 18750 2975
rect 18790 2975 18805 2985
rect 18790 2960 18885 2975
rect 18105 2940 18115 2960
rect 18135 2940 18145 2960
rect 18105 2930 18145 2940
rect 18313 2940 18321 2960
rect 18339 2940 18347 2960
rect 18313 2930 18347 2940
rect 18845 2940 18855 2960
rect 18875 2940 18885 2960
rect 26260 3605 26280 3620
rect 26320 3605 26340 3620
rect 26380 3605 26400 3620
rect 26440 3605 26460 3620
rect 26500 3605 26520 3620
rect 26560 3605 26580 3620
rect 26620 3605 26640 3620
rect 26680 3605 26700 3620
rect 26740 3605 26760 3620
rect 26800 3605 26820 3620
rect 26860 3605 26880 3620
rect 26920 3605 26940 3620
rect 26980 3605 27000 3620
rect 27040 3605 27060 3620
rect 27100 3605 27120 3620
rect 27160 3605 27180 3620
rect 27220 3605 27240 3620
rect 27280 3605 27300 3620
rect 27340 3605 27360 3620
rect 27400 3605 27420 3620
rect 27460 3605 27480 3620
rect 27520 3605 27540 3620
rect 26260 3190 26280 3205
rect 26320 3195 26340 3205
rect 26380 3195 26400 3205
rect 26440 3195 26460 3205
rect 26500 3195 26520 3205
rect 26560 3195 26580 3205
rect 26620 3195 26640 3205
rect 26680 3195 26700 3205
rect 26740 3195 26760 3205
rect 26800 3195 26820 3205
rect 26860 3195 26880 3205
rect 26920 3195 26940 3205
rect 26980 3195 27000 3205
rect 27040 3195 27060 3205
rect 27100 3195 27120 3205
rect 27160 3195 27180 3205
rect 27220 3195 27240 3205
rect 27280 3195 27300 3205
rect 27340 3195 27360 3205
rect 27400 3195 27420 3205
rect 27460 3195 27480 3205
rect 26320 3180 27480 3195
rect 27520 3190 27540 3205
rect 26823 3160 26831 3180
rect 26849 3160 26857 3180
rect 26823 3150 26857 3160
rect 28185 3665 28200 3680
rect 28240 3665 28255 3680
rect 28295 3665 28310 3680
rect 28350 3665 28365 3680
rect 28405 3665 28420 3680
rect 28460 3665 28475 3680
rect 28515 3665 28530 3680
rect 28570 3665 28585 3680
rect 28625 3665 28640 3680
rect 28680 3665 28695 3680
rect 28735 3665 28750 3680
rect 28790 3665 28805 3680
rect 28185 3050 28200 3065
rect 28240 3055 28255 3065
rect 28295 3055 28310 3065
rect 28350 3055 28365 3065
rect 28405 3055 28420 3065
rect 28460 3055 28475 3065
rect 28515 3055 28530 3065
rect 28570 3055 28585 3065
rect 28625 3055 28640 3065
rect 28680 3055 28695 3065
rect 28735 3055 28750 3065
rect 28240 3040 28750 3055
rect 28790 3050 28805 3065
rect 28313 3020 28321 3040
rect 28339 3020 28347 3040
rect 28313 3010 28347 3020
rect 25045 2975 25060 2985
rect 24965 2960 25060 2975
rect 25100 2975 25115 2985
rect 25155 2975 25170 2985
rect 25210 2975 25225 2985
rect 25265 2975 25280 2985
rect 25320 2975 25335 2985
rect 25375 2975 25390 2985
rect 25430 2975 25445 2985
rect 25485 2975 25500 2985
rect 25540 2975 25555 2985
rect 25595 2975 25610 2985
rect 25100 2960 25610 2975
rect 25650 2975 25665 2985
rect 25650 2960 25745 2975
rect 24965 2940 24975 2960
rect 24995 2940 25005 2960
rect 18845 2930 18885 2940
rect 24965 2930 25005 2940
rect 25503 2940 25511 2960
rect 25529 2940 25537 2960
rect 25503 2930 25537 2940
rect 25705 2940 25715 2960
rect 25735 2940 25745 2960
rect 25705 2930 25745 2940
rect 15975 2890 16015 2900
rect 15975 2870 15985 2890
rect 16005 2870 16015 2890
rect 16775 2890 16815 2900
rect 16775 2870 16785 2890
rect 16805 2870 16815 2890
rect 15975 2855 16075 2870
rect 16055 2845 16075 2855
rect 16115 2845 16135 2860
rect 16175 2845 16195 2860
rect 16235 2845 16255 2860
rect 16295 2845 16315 2860
rect 16355 2845 16375 2860
rect 16415 2845 16435 2860
rect 16475 2845 16495 2860
rect 16535 2845 16555 2860
rect 16595 2845 16615 2860
rect 16655 2845 16675 2860
rect 16715 2855 16815 2870
rect 16985 2890 17025 2900
rect 16985 2870 16995 2890
rect 17015 2870 17025 2890
rect 17785 2890 17825 2900
rect 17785 2870 17795 2890
rect 17815 2870 17825 2890
rect 16985 2855 17085 2870
rect 16715 2845 16735 2855
rect 17065 2845 17085 2855
rect 17125 2845 17145 2860
rect 17185 2845 17205 2860
rect 17245 2845 17265 2860
rect 17305 2845 17325 2860
rect 17365 2845 17385 2860
rect 17425 2845 17445 2860
rect 17485 2845 17505 2860
rect 17545 2845 17565 2860
rect 17605 2845 17625 2860
rect 17665 2845 17685 2860
rect 17725 2855 17825 2870
rect 25975 2890 26015 2900
rect 25975 2870 25985 2890
rect 26005 2870 26015 2890
rect 26775 2890 26815 2900
rect 26775 2870 26785 2890
rect 26805 2870 26815 2890
rect 25975 2855 26075 2870
rect 17725 2845 17745 2855
rect 26055 2845 26075 2855
rect 26115 2845 26135 2860
rect 26175 2845 26195 2860
rect 26235 2845 26255 2860
rect 26295 2845 26315 2860
rect 26355 2845 26375 2860
rect 26415 2845 26435 2860
rect 26475 2845 26495 2860
rect 26535 2845 26555 2860
rect 26595 2845 26615 2860
rect 26655 2845 26675 2860
rect 26715 2855 26815 2870
rect 26715 2845 26735 2855
rect 3035 2815 3085 2830
rect 2995 2805 3085 2815
rect 3125 2820 3175 2830
rect 3215 2820 3265 2830
rect 3305 2820 3355 2830
rect 3395 2820 3445 2830
rect 3485 2820 3535 2830
rect 3575 2820 3625 2830
rect 3665 2820 3715 2830
rect 3755 2820 3805 2830
rect 3845 2820 3895 2830
rect 3935 2820 3985 2830
rect 4025 2820 4075 2830
rect 4115 2820 4165 2830
rect 4205 2820 4255 2830
rect 4295 2820 4345 2830
rect 4385 2820 4435 2830
rect 4475 2820 4525 2830
rect 4565 2820 4615 2830
rect 4655 2820 4705 2830
rect 4745 2820 4795 2830
rect 4835 2820 4885 2830
rect 3125 2805 4885 2820
rect 4925 2815 4975 2830
rect 4925 2805 5015 2815
rect 2995 2785 3005 2805
rect 3025 2800 3085 2805
rect 4925 2800 4985 2805
rect 3025 2785 3035 2800
rect 2995 2775 3035 2785
rect 4975 2785 4985 2800
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2730 3215 2745
rect 4795 2745 4835 2755
rect 4795 2730 4805 2745
rect 3205 2725 3265 2730
rect 3175 2715 3265 2725
rect 4745 2725 4805 2730
rect 4825 2725 4835 2745
rect 4745 2715 4835 2725
rect 3215 2700 3265 2715
rect 3305 2700 3355 2715
rect 3395 2700 3445 2715
rect 3485 2700 3535 2715
rect 3575 2700 3625 2715
rect 3665 2700 3715 2715
rect 3755 2700 3805 2715
rect 3845 2700 3895 2715
rect 3935 2700 3985 2715
rect 4025 2700 4075 2715
rect 4115 2700 4165 2715
rect 4205 2700 4255 2715
rect 4295 2700 4345 2715
rect 4385 2700 4435 2715
rect 4475 2700 4525 2715
rect 4565 2700 4615 2715
rect 4655 2700 4705 2715
rect 4745 2700 4795 2715
rect 15045 2655 15060 2670
rect 15100 2655 15115 2670
rect 15155 2655 15170 2670
rect 15210 2655 15225 2670
rect 15265 2655 15280 2670
rect 15320 2655 15335 2670
rect 15375 2655 15390 2670
rect 15430 2655 15445 2670
rect 15485 2655 15500 2670
rect 15540 2655 15555 2670
rect 15595 2655 15610 2670
rect 15650 2655 15665 2670
rect 3215 2385 3265 2400
rect 3305 2390 3355 2400
rect 3395 2390 3445 2400
rect 3485 2390 3535 2400
rect 3575 2390 3625 2400
rect 3665 2390 3715 2400
rect 3755 2390 3805 2400
rect 3845 2390 3895 2400
rect 3935 2390 3985 2400
rect 4025 2390 4075 2400
rect 4115 2390 4165 2400
rect 4205 2390 4255 2400
rect 4295 2390 4345 2400
rect 4385 2390 4435 2400
rect 4475 2390 4525 2400
rect 4565 2390 4615 2400
rect 4655 2390 4705 2400
rect 3305 2375 4705 2390
rect 4745 2385 4795 2400
rect 3355 2370 3395 2375
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 3355 2340 3395 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 5205 2000 5225 2015
rect 18185 2655 18200 2670
rect 18240 2655 18255 2670
rect 18295 2655 18310 2670
rect 18350 2655 18365 2670
rect 18405 2655 18420 2670
rect 18460 2655 18475 2670
rect 18515 2655 18530 2670
rect 18570 2655 18585 2670
rect 18625 2655 18640 2670
rect 18680 2655 18695 2670
rect 18735 2655 18750 2670
rect 18790 2655 18805 2670
rect 25045 2655 25060 2670
rect 25100 2655 25115 2670
rect 25155 2655 25170 2670
rect 25210 2655 25225 2670
rect 25265 2655 25280 2670
rect 25320 2655 25335 2670
rect 25375 2655 25390 2670
rect 25430 2655 25445 2670
rect 25485 2655 25500 2670
rect 25540 2655 25555 2670
rect 25595 2655 25610 2670
rect 25650 2655 25665 2670
rect 16055 2480 16075 2495
rect 16115 2485 16135 2495
rect 16175 2485 16195 2495
rect 16235 2485 16255 2495
rect 16295 2485 16315 2495
rect 16355 2485 16375 2495
rect 16415 2485 16435 2495
rect 16475 2485 16495 2495
rect 16535 2485 16555 2495
rect 16595 2485 16615 2495
rect 16655 2485 16675 2495
rect 16115 2470 16675 2485
rect 16715 2480 16735 2495
rect 17065 2480 17085 2495
rect 17125 2485 17145 2495
rect 17185 2485 17205 2495
rect 17245 2485 17265 2495
rect 17305 2485 17325 2495
rect 17365 2485 17385 2495
rect 17425 2485 17445 2495
rect 17485 2485 17505 2495
rect 17545 2485 17565 2495
rect 17605 2485 17625 2495
rect 17665 2485 17685 2495
rect 17125 2470 17685 2485
rect 17725 2480 17745 2495
rect 15045 2445 15060 2455
rect 14965 2430 15060 2445
rect 15100 2445 15115 2455
rect 15155 2445 15170 2455
rect 15210 2445 15225 2455
rect 15265 2445 15280 2455
rect 15320 2445 15335 2455
rect 15375 2445 15390 2455
rect 15430 2445 15445 2455
rect 15485 2445 15500 2455
rect 15540 2445 15555 2455
rect 15595 2445 15610 2455
rect 15100 2430 15610 2445
rect 15650 2445 15665 2455
rect 16378 2450 16386 2470
rect 16404 2450 16412 2470
rect 15650 2430 15745 2445
rect 16378 2440 16412 2450
rect 17388 2450 17396 2470
rect 17414 2450 17422 2470
rect 17388 2440 17422 2450
rect 18185 2445 18200 2455
rect 14965 2410 14975 2430
rect 14995 2410 15005 2430
rect 14965 2400 15005 2410
rect 15595 2380 15610 2430
rect 15705 2410 15715 2430
rect 15735 2410 15745 2430
rect 15705 2400 15745 2410
rect 18105 2430 18200 2445
rect 18240 2445 18255 2455
rect 18295 2445 18310 2455
rect 18350 2445 18365 2455
rect 18405 2445 18420 2455
rect 18460 2445 18475 2455
rect 18515 2445 18530 2455
rect 18570 2445 18585 2455
rect 18625 2445 18640 2455
rect 18680 2445 18695 2455
rect 18735 2445 18750 2455
rect 18240 2430 18750 2445
rect 18790 2445 18805 2455
rect 18790 2430 18885 2445
rect 18105 2410 18115 2430
rect 18135 2410 18145 2430
rect 18105 2400 18145 2410
rect 18240 2380 18255 2430
rect 18845 2410 18855 2430
rect 18875 2410 18885 2430
rect 18845 2400 18885 2410
rect 15585 2370 15625 2380
rect 15585 2350 15595 2370
rect 15615 2350 15625 2370
rect 15585 2340 15625 2350
rect 18225 2370 18265 2380
rect 18225 2350 18235 2370
rect 18255 2350 18265 2370
rect 18225 2340 18265 2350
rect 14965 2310 15005 2320
rect 14965 2290 14975 2310
rect 14995 2290 15005 2310
rect 15595 2290 15610 2340
rect 15705 2310 15745 2320
rect 15705 2290 15715 2310
rect 15735 2290 15745 2310
rect 14965 2275 15060 2290
rect 15045 2265 15060 2275
rect 15100 2275 15610 2290
rect 15100 2265 15115 2275
rect 15155 2265 15170 2275
rect 15210 2265 15225 2275
rect 15265 2265 15280 2275
rect 15320 2265 15335 2275
rect 15375 2265 15390 2275
rect 15430 2265 15445 2275
rect 15485 2265 15500 2275
rect 15540 2265 15555 2275
rect 15595 2265 15610 2275
rect 15650 2275 15745 2290
rect 18105 2310 18145 2320
rect 18105 2290 18115 2310
rect 18135 2290 18145 2310
rect 18240 2290 18255 2340
rect 18845 2310 18885 2320
rect 18845 2290 18855 2310
rect 18875 2290 18885 2310
rect 18105 2275 18200 2290
rect 15650 2265 15665 2275
rect 18185 2265 18200 2275
rect 18240 2275 18750 2290
rect 18240 2265 18255 2275
rect 18295 2265 18310 2275
rect 18350 2265 18365 2275
rect 18405 2265 18420 2275
rect 18460 2265 18475 2275
rect 18515 2265 18530 2275
rect 18570 2265 18585 2275
rect 18625 2265 18640 2275
rect 18680 2265 18695 2275
rect 18735 2265 18750 2275
rect 18790 2275 18885 2290
rect 18790 2265 18805 2275
rect 16828 2175 16862 2185
rect 16828 2155 16836 2175
rect 16854 2155 16862 2175
rect 16315 2130 16330 2145
rect 16370 2140 17430 2155
rect 16370 2130 16385 2140
rect 16425 2130 16440 2140
rect 16480 2130 16495 2140
rect 16535 2130 16550 2140
rect 16590 2130 16605 2140
rect 16645 2130 16660 2140
rect 16700 2130 16715 2140
rect 16755 2130 16770 2140
rect 16810 2130 16825 2140
rect 16865 2130 16880 2140
rect 16920 2130 16935 2140
rect 16975 2130 16990 2140
rect 17030 2130 17045 2140
rect 17085 2130 17100 2140
rect 17140 2130 17155 2140
rect 17195 2130 17210 2140
rect 17250 2130 17265 2140
rect 17305 2130 17320 2140
rect 17360 2130 17375 2140
rect 17415 2130 17430 2140
rect 17470 2130 17485 2145
rect 16315 1970 16330 1980
rect 15045 1950 15060 1965
rect 15100 1950 15115 1965
rect 15155 1950 15170 1965
rect 15210 1950 15225 1965
rect 15265 1950 15280 1965
rect 15320 1950 15335 1965
rect 15375 1950 15390 1965
rect 15430 1950 15445 1965
rect 15485 1950 15500 1965
rect 15540 1950 15555 1965
rect 15595 1950 15610 1965
rect 15650 1950 15665 1965
rect 16235 1955 16330 1970
rect 16370 1965 16385 1980
rect 16425 1965 16440 1980
rect 16480 1965 16495 1980
rect 16535 1965 16550 1980
rect 16590 1965 16605 1980
rect 16645 1965 16660 1980
rect 16700 1965 16715 1980
rect 16755 1965 16770 1980
rect 16810 1965 16825 1980
rect 16865 1965 16880 1980
rect 16920 1965 16935 1980
rect 16975 1965 16990 1980
rect 17030 1965 17045 1980
rect 17085 1965 17100 1980
rect 17140 1965 17155 1980
rect 17195 1965 17210 1980
rect 17250 1965 17265 1980
rect 17305 1965 17320 1980
rect 17360 1965 17375 1980
rect 17415 1965 17430 1980
rect 17470 1970 17485 1980
rect 17470 1955 17565 1970
rect 27075 2845 27095 2860
rect 27135 2845 27155 2860
rect 27195 2845 27215 2860
rect 27255 2845 27275 2860
rect 27315 2845 27335 2860
rect 27375 2845 27395 2860
rect 27435 2845 27455 2860
rect 27495 2845 27515 2860
rect 27555 2845 27575 2860
rect 27615 2845 27635 2860
rect 27675 2845 27695 2860
rect 27735 2845 27755 2860
rect 26055 2480 26075 2495
rect 26115 2485 26135 2495
rect 26175 2485 26195 2495
rect 26235 2485 26255 2495
rect 26295 2485 26315 2495
rect 26355 2485 26375 2495
rect 26415 2485 26435 2495
rect 26475 2485 26495 2495
rect 26535 2485 26555 2495
rect 26595 2485 26615 2495
rect 26655 2485 26675 2495
rect 26115 2470 26675 2485
rect 26715 2480 26735 2495
rect 25045 2445 25060 2455
rect 24965 2430 25060 2445
rect 25100 2445 25115 2455
rect 25155 2445 25170 2455
rect 25210 2445 25225 2455
rect 25265 2445 25280 2455
rect 25320 2445 25335 2455
rect 25375 2445 25390 2455
rect 25430 2445 25445 2455
rect 25485 2445 25500 2455
rect 25540 2445 25555 2455
rect 25595 2445 25610 2455
rect 25100 2430 25610 2445
rect 25650 2445 25665 2455
rect 26378 2450 26386 2470
rect 26404 2450 26412 2470
rect 25650 2430 25745 2445
rect 26378 2440 26412 2450
rect 24965 2410 24975 2430
rect 24995 2410 25005 2430
rect 24965 2400 25005 2410
rect 25595 2380 25610 2430
rect 25705 2410 25715 2430
rect 25735 2410 25745 2430
rect 25705 2400 25745 2410
rect 27075 2480 27095 2495
rect 27135 2485 27155 2495
rect 27195 2485 27215 2495
rect 27255 2485 27275 2495
rect 27315 2485 27335 2495
rect 27375 2485 27395 2495
rect 27435 2485 27455 2495
rect 27495 2485 27515 2495
rect 27555 2485 27575 2495
rect 27615 2485 27635 2495
rect 27675 2485 27695 2495
rect 27135 2470 27695 2485
rect 27735 2480 27755 2495
rect 27398 2450 27406 2470
rect 27424 2450 27432 2470
rect 27398 2440 27432 2450
rect 28185 2705 28200 2720
rect 28240 2705 28255 2720
rect 28295 2705 28310 2720
rect 28350 2705 28365 2720
rect 28405 2705 28420 2720
rect 28460 2705 28475 2720
rect 28515 2705 28530 2720
rect 28570 2705 28585 2720
rect 28625 2705 28640 2720
rect 28680 2705 28695 2720
rect 28735 2705 28750 2720
rect 28790 2705 28805 2720
rect 28185 2490 28200 2505
rect 28240 2495 28255 2505
rect 28295 2495 28310 2505
rect 28350 2495 28365 2505
rect 28405 2495 28420 2505
rect 28460 2495 28475 2505
rect 28515 2495 28530 2505
rect 28570 2495 28585 2505
rect 28625 2495 28640 2505
rect 28680 2495 28695 2505
rect 28735 2495 28750 2505
rect 28240 2480 28750 2495
rect 28790 2490 28805 2505
rect 28313 2460 28321 2480
rect 28339 2460 28347 2480
rect 28313 2450 28347 2460
rect 25585 2370 25625 2380
rect 25585 2350 25595 2370
rect 25615 2350 25625 2370
rect 25585 2340 25625 2350
rect 24965 2310 25005 2320
rect 24965 2290 24975 2310
rect 24995 2290 25005 2310
rect 25595 2290 25610 2340
rect 25705 2310 25745 2320
rect 25705 2290 25715 2310
rect 25735 2290 25745 2310
rect 24965 2275 25060 2290
rect 25045 2265 25060 2275
rect 25100 2275 25610 2290
rect 25100 2265 25115 2275
rect 25155 2265 25170 2275
rect 25210 2265 25225 2275
rect 25265 2265 25280 2275
rect 25320 2265 25335 2275
rect 25375 2265 25390 2275
rect 25430 2265 25445 2275
rect 25485 2265 25500 2275
rect 25540 2265 25555 2275
rect 25595 2265 25610 2275
rect 25650 2275 25745 2290
rect 25650 2265 25665 2275
rect 26828 2175 26862 2185
rect 26828 2155 26836 2175
rect 26854 2155 26862 2175
rect 26315 2130 26330 2145
rect 26370 2140 27430 2155
rect 26370 2130 26385 2140
rect 26425 2130 26440 2140
rect 26480 2130 26495 2140
rect 26535 2130 26550 2140
rect 26590 2130 26605 2140
rect 26645 2130 26660 2140
rect 26700 2130 26715 2140
rect 26755 2130 26770 2140
rect 26810 2130 26825 2140
rect 26865 2130 26880 2140
rect 26920 2130 26935 2140
rect 26975 2130 26990 2140
rect 27030 2130 27045 2140
rect 27085 2130 27100 2140
rect 27140 2130 27155 2140
rect 27195 2130 27210 2140
rect 27250 2130 27265 2140
rect 27305 2130 27320 2140
rect 27360 2130 27375 2140
rect 27415 2130 27430 2140
rect 27470 2130 27485 2145
rect 16235 1935 16245 1955
rect 16265 1935 16275 1955
rect 16235 1925 16275 1935
rect 17525 1935 17535 1955
rect 17555 1935 17565 1955
rect 18185 1950 18200 1965
rect 18240 1950 18255 1965
rect 18295 1950 18310 1965
rect 18350 1950 18365 1965
rect 18405 1950 18420 1965
rect 18460 1950 18475 1965
rect 18515 1950 18530 1965
rect 18570 1950 18585 1965
rect 18625 1950 18640 1965
rect 18680 1950 18695 1965
rect 18735 1950 18750 1965
rect 18790 1950 18805 1965
rect 25045 1950 25060 1965
rect 25100 1950 25115 1965
rect 25155 1950 25170 1965
rect 25210 1950 25225 1965
rect 25265 1950 25280 1965
rect 25320 1950 25335 1965
rect 25375 1950 25390 1965
rect 25430 1950 25445 1965
rect 25485 1950 25500 1965
rect 25540 1950 25555 1965
rect 25595 1950 25610 1965
rect 25650 1950 25665 1965
rect 17525 1925 17565 1935
rect 26315 1965 26330 1980
rect 26370 1965 26385 1980
rect 26425 1965 26440 1980
rect 26480 1965 26495 1980
rect 26535 1965 26550 1980
rect 26590 1965 26605 1980
rect 26645 1965 26660 1980
rect 26700 1965 26715 1980
rect 26755 1965 26770 1980
rect 26810 1965 26825 1980
rect 26865 1965 26880 1980
rect 26920 1965 26935 1980
rect 26975 1965 26990 1980
rect 27030 1965 27045 1980
rect 27085 1965 27100 1980
rect 27140 1965 27155 1980
rect 27195 1965 27210 1980
rect 27250 1965 27265 1980
rect 27305 1965 27320 1980
rect 27360 1965 27375 1980
rect 27415 1965 27430 1980
rect 27470 1965 27485 1980
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2765 1875 2805 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2765 1855 2775 1875
rect 2795 1855 2805 1875
rect 2765 1845 2805 1855
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1890 3945 1900
rect 4065 1890 4085 1900
rect 3855 1875 3895 1885
rect 3925 1875 4085 1890
rect 4125 1885 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 4365 1890 4385 1900
rect 4115 1875 4155 1885
rect 4185 1875 4385 1890
rect 4425 1890 4445 1900
rect 4485 1890 4505 1900
rect 4425 1875 4505 1890
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4725 1890 4745 1900
rect 4545 1875 4745 1890
rect 4785 1890 4805 1900
rect 4845 1890 4865 1900
rect 4785 1875 4865 1890
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 5085 1890 5105 1900
rect 4905 1875 5105 1890
rect 5145 1885 5165 1900
rect 5205 1885 5225 1900
rect 28313 2290 28347 2300
rect 28313 2270 28321 2290
rect 28339 2270 28347 2290
rect 28185 2245 28200 2260
rect 28240 2255 28750 2270
rect 28240 2245 28255 2255
rect 28295 2245 28310 2255
rect 28350 2245 28365 2255
rect 28405 2245 28420 2255
rect 28460 2245 28475 2255
rect 28515 2245 28530 2255
rect 28570 2245 28585 2255
rect 28625 2245 28640 2255
rect 28680 2245 28695 2255
rect 28735 2245 28750 2255
rect 28790 2245 28805 2260
rect 5135 1875 5175 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1875
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5245 1885
rect 5205 1855 5215 1875
rect 5235 1855 5245 1875
rect 5205 1845 5245 1855
rect 28185 1930 28200 1945
rect 28240 1930 28255 1945
rect 28295 1930 28310 1945
rect 28350 1930 28365 1945
rect 28405 1930 28420 1945
rect 28460 1930 28475 1945
rect 28515 1930 28530 1945
rect 28570 1930 28585 1945
rect 28625 1930 28640 1945
rect 28680 1930 28695 1945
rect 28735 1930 28750 1945
rect 28790 1930 28805 1945
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1720 4785 1735
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4245 1705 4785 1720
rect 16237 1710 16269 1720
rect 4245 1665 4265 1705
rect 4305 1665 4325 1680
rect 4365 1665 4385 1680
rect 4425 1665 4445 1705
rect 4485 1665 4505 1705
rect 4545 1665 4565 1680
rect 4605 1665 4625 1680
rect 4665 1665 4685 1705
rect 4725 1665 4745 1705
rect 15408 1700 15442 1710
rect 15408 1680 15416 1700
rect 15434 1680 15442 1700
rect 16237 1690 16243 1710
rect 16260 1690 16269 1710
rect 16457 1710 16489 1720
rect 16457 1690 16463 1710
rect 16480 1690 16489 1710
rect 16180 1680 16269 1690
rect 16400 1680 16489 1690
rect 16601 1710 16635 1720
rect 16601 1690 16610 1710
rect 16627 1690 16635 1710
rect 16867 1710 16899 1720
rect 16867 1695 16876 1710
rect 16601 1680 16635 1690
rect 16865 1690 16876 1695
rect 16893 1690 16899 1710
rect 17277 1710 17309 1720
rect 17277 1690 17283 1710
rect 17300 1690 17309 1710
rect 17497 1710 17529 1720
rect 17497 1690 17503 1710
rect 17520 1690 17529 1710
rect 16865 1680 16899 1690
rect 17220 1680 17309 1690
rect 17440 1680 17529 1690
rect 17641 1710 17675 1720
rect 17641 1690 17650 1710
rect 17667 1690 17675 1710
rect 17641 1680 17675 1690
rect 18408 1700 18442 1710
rect 18408 1680 18416 1700
rect 18434 1680 18442 1700
rect 25408 1700 25442 1710
rect 25408 1680 25416 1700
rect 25434 1680 25442 1700
rect 4785 1665 4805 1680
rect 15045 1655 15105 1670
rect 15145 1665 15505 1680
rect 15145 1655 15205 1665
rect 15245 1655 15305 1665
rect 15345 1655 15405 1665
rect 15445 1655 15505 1665
rect 15545 1655 15605 1670
rect 16070 1665 16085 1680
rect 16125 1665 16140 1680
rect 16180 1675 16250 1680
rect 16180 1665 16195 1675
rect 16235 1665 16250 1675
rect 16290 1665 16305 1680
rect 16345 1665 16360 1680
rect 16400 1675 16470 1680
rect 16400 1665 16415 1675
rect 16455 1665 16470 1675
rect 16510 1665 16525 1680
rect 16565 1665 16580 1680
rect 16620 1665 16635 1680
rect 16675 1665 16690 1680
rect 16810 1665 16825 1680
rect 16865 1665 16880 1680
rect 16920 1665 16935 1680
rect 16975 1665 16990 1680
rect 17110 1665 17125 1680
rect 17165 1665 17180 1680
rect 17220 1675 17290 1680
rect 17220 1665 17235 1675
rect 17275 1665 17290 1675
rect 17330 1665 17345 1680
rect 17385 1665 17400 1680
rect 17440 1675 17510 1680
rect 17440 1665 17455 1675
rect 17495 1665 17510 1675
rect 17550 1665 17565 1680
rect 17605 1665 17620 1680
rect 17660 1665 17675 1680
rect 17715 1665 17730 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4245 1600 4265 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4305 1575 4325 1615
rect 4365 1575 4385 1615
rect 4425 1600 4445 1615
rect 4485 1600 4505 1615
rect 4545 1575 4565 1615
rect 4605 1575 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4785 1600 4805 1615
rect 4785 1590 4845 1600
rect 4785 1575 4815 1590
rect 4305 1570 4815 1575
rect 4835 1570 4845 1590
rect 4305 1560 4845 1570
rect 2925 1495 2965 1505
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1470 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1470 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1470 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1470 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1470 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1470 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 3765 1470 3805 1475
rect 4205 1495 4245 1505
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1470 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1470 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1470 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1470 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1470 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1470 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1470 5085 1475
rect 2875 1455 3375 1470
rect 3415 1455 3915 1470
rect 4095 1455 4595 1470
rect 4635 1455 5135 1470
rect 2875 1190 3375 1205
rect 3415 1190 3915 1205
rect 4095 1190 4595 1205
rect 4635 1190 5135 1205
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2985 1075 3985 1090
rect 4025 1075 5025 1090
rect 2985 960 3985 975
rect 4025 960 5025 975
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 18245 1655 18305 1670
rect 18345 1665 18705 1680
rect 18345 1655 18405 1665
rect 18445 1655 18505 1665
rect 18545 1655 18605 1665
rect 18645 1655 18705 1665
rect 18745 1655 18805 1670
rect 25045 1655 25105 1670
rect 25145 1665 25505 1680
rect 25145 1655 25205 1665
rect 25245 1655 25305 1665
rect 25345 1655 25405 1665
rect 25445 1655 25505 1665
rect 25545 1655 25605 1670
rect 16070 1505 16085 1515
rect 15990 1490 16085 1505
rect 16125 1500 16140 1515
rect 16180 1500 16195 1515
rect 16235 1500 16250 1515
rect 16290 1505 16305 1515
rect 16345 1505 16360 1515
rect 16106 1490 16140 1500
rect 16290 1490 16360 1505
rect 16400 1500 16415 1515
rect 16455 1500 16470 1515
rect 16510 1505 16525 1515
rect 16565 1505 16580 1515
rect 16510 1490 16580 1505
rect 16620 1500 16635 1515
rect 16675 1505 16690 1515
rect 16810 1505 16825 1515
rect 16675 1490 16825 1505
rect 16865 1500 16880 1515
rect 16920 1500 16935 1515
rect 16975 1505 16990 1515
rect 17110 1505 17125 1515
rect 16920 1490 16954 1500
rect 16975 1490 17125 1505
rect 17165 1500 17180 1515
rect 17220 1500 17235 1515
rect 17275 1500 17290 1515
rect 17330 1505 17345 1515
rect 17385 1505 17400 1515
rect 17146 1490 17180 1500
rect 17330 1490 17400 1505
rect 17440 1500 17455 1515
rect 17495 1500 17510 1515
rect 17550 1505 17565 1515
rect 17605 1505 17620 1515
rect 17550 1490 17620 1505
rect 17660 1500 17675 1515
rect 17715 1505 17730 1515
rect 17715 1490 17810 1505
rect 15990 1470 16000 1490
rect 16020 1470 16030 1490
rect 15990 1460 16030 1470
rect 16106 1470 16112 1490
rect 16129 1470 16138 1490
rect 16106 1460 16138 1470
rect 16305 1470 16315 1490
rect 16335 1470 16345 1490
rect 16305 1460 16345 1470
rect 16525 1470 16535 1490
rect 16555 1470 16565 1490
rect 16525 1460 16565 1470
rect 16730 1470 16740 1490
rect 16760 1470 16770 1490
rect 16730 1460 16770 1470
rect 16922 1470 16928 1490
rect 16945 1470 16954 1490
rect 16922 1460 16954 1470
rect 17030 1470 17040 1490
rect 17060 1470 17070 1490
rect 17030 1460 17070 1470
rect 17146 1470 17152 1490
rect 17169 1470 17178 1490
rect 17146 1460 17178 1470
rect 17345 1470 17355 1490
rect 17375 1470 17385 1490
rect 17345 1460 17385 1470
rect 17565 1470 17575 1490
rect 17595 1470 17605 1490
rect 17565 1460 17605 1470
rect 17770 1470 17780 1490
rect 17800 1470 17810 1490
rect 17770 1460 17810 1470
rect 17595 1245 17635 1255
rect 17595 1240 17605 1245
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 17510 1225 17605 1240
rect 17625 1225 17635 1245
rect 16245 1185 16260 1200
rect 16300 1195 17360 1210
rect 16300 1185 16315 1195
rect 16355 1185 16370 1195
rect 16410 1185 16425 1195
rect 16465 1185 16480 1195
rect 16520 1185 16535 1195
rect 16575 1185 16590 1195
rect 16630 1185 16645 1195
rect 16685 1185 16700 1195
rect 16740 1185 16755 1195
rect 16795 1185 16810 1195
rect 16850 1185 16865 1195
rect 16905 1185 16920 1195
rect 16960 1185 16975 1195
rect 17015 1185 17030 1195
rect 17070 1185 17085 1195
rect 17125 1185 17140 1195
rect 17180 1185 17195 1195
rect 17235 1185 17250 1195
rect 17290 1185 17305 1195
rect 17345 1185 17360 1195
rect 17400 1195 17470 1210
rect 17400 1185 17415 1195
rect 17455 1185 17470 1195
rect 17510 1185 17525 1225
rect 17595 1215 17635 1225
rect 17565 1185 17580 1200
rect 15045 945 15105 955
rect 14965 930 15105 945
rect 15145 940 15205 955
rect 15245 940 15305 955
rect 15345 940 15405 955
rect 15445 940 15505 955
rect 15545 945 15605 955
rect 15545 930 15685 945
rect 18245 945 18305 955
rect 14965 910 14975 930
rect 14995 910 15005 930
rect 2995 890 3085 905
rect 3035 880 3085 890
rect 3125 890 4885 905
rect 3125 880 3175 890
rect 3215 880 3265 890
rect 3305 880 3355 890
rect 3395 880 3445 890
rect 3485 880 3535 890
rect 3575 880 3625 890
rect 3665 880 3715 890
rect 3755 880 3805 890
rect 3845 880 3895 890
rect 3935 880 3985 890
rect 4025 880 4075 890
rect 4115 880 4165 890
rect 4205 880 4255 890
rect 4295 880 4345 890
rect 4385 880 4435 890
rect 4475 880 4525 890
rect 4565 880 4615 890
rect 4655 880 4705 890
rect 4745 880 4795 890
rect 4835 880 4885 890
rect 4925 890 5015 905
rect 14965 900 15005 910
rect 15645 910 15655 930
rect 15675 910 15685 930
rect 16245 920 16260 935
rect 16300 920 16315 935
rect 16355 920 16370 935
rect 16410 920 16425 935
rect 16465 920 16480 935
rect 16520 920 16535 935
rect 16575 920 16590 935
rect 16630 920 16645 935
rect 16685 920 16700 935
rect 16740 920 16755 935
rect 16795 920 16810 935
rect 16850 920 16865 935
rect 16905 920 16920 935
rect 16960 920 16975 935
rect 17015 920 17030 935
rect 17070 920 17085 935
rect 17125 920 17140 935
rect 17180 920 17195 935
rect 17235 920 17250 935
rect 17290 920 17305 935
rect 17345 920 17360 935
rect 17400 920 17415 935
rect 17455 920 17470 935
rect 17510 920 17525 935
rect 17565 920 17580 935
rect 18165 930 18305 945
rect 18345 940 18405 955
rect 18445 940 18505 955
rect 18545 940 18605 955
rect 18645 940 18705 955
rect 18745 945 18805 955
rect 18745 930 18885 945
rect 15645 900 15685 910
rect 16165 910 16260 920
rect 16165 890 16175 910
rect 16195 905 16260 910
rect 17565 910 17660 920
rect 17565 905 17630 910
rect 16195 890 16205 905
rect 4925 880 4975 890
rect 16165 880 16205 890
rect 17620 890 17630 905
rect 17650 890 17660 910
rect 18165 910 18175 930
rect 18195 910 18205 930
rect 18165 900 18205 910
rect 18845 910 18855 930
rect 18875 910 18885 930
rect 26237 1710 26269 1720
rect 26237 1690 26243 1710
rect 26260 1690 26269 1710
rect 26457 1710 26489 1720
rect 26457 1690 26463 1710
rect 26480 1690 26489 1710
rect 26180 1680 26269 1690
rect 26400 1680 26489 1690
rect 26601 1710 26635 1720
rect 26601 1690 26610 1710
rect 26627 1690 26635 1710
rect 26867 1710 26899 1720
rect 26867 1695 26876 1710
rect 26601 1680 26635 1690
rect 26865 1690 26876 1695
rect 26893 1690 26899 1710
rect 27277 1710 27309 1720
rect 27277 1690 27283 1710
rect 27300 1690 27309 1710
rect 27497 1710 27529 1720
rect 27497 1690 27503 1710
rect 27520 1690 27529 1710
rect 26865 1680 26899 1690
rect 27220 1680 27309 1690
rect 27440 1680 27529 1690
rect 27641 1710 27675 1720
rect 27641 1690 27650 1710
rect 27667 1690 27675 1710
rect 27641 1680 27675 1690
rect 26070 1665 26085 1680
rect 26125 1665 26140 1680
rect 26180 1675 26250 1680
rect 26180 1665 26195 1675
rect 26235 1665 26250 1675
rect 26290 1665 26305 1680
rect 26345 1665 26360 1680
rect 26400 1675 26470 1680
rect 26400 1665 26415 1675
rect 26455 1665 26470 1675
rect 26510 1665 26525 1680
rect 26565 1665 26580 1680
rect 26620 1665 26635 1680
rect 26675 1665 26690 1680
rect 26810 1665 26825 1680
rect 26865 1665 26880 1680
rect 26920 1665 26935 1680
rect 26975 1665 26990 1680
rect 27110 1665 27125 1680
rect 27165 1665 27180 1680
rect 27220 1675 27290 1680
rect 27220 1665 27235 1675
rect 27275 1665 27290 1675
rect 27330 1665 27345 1680
rect 27385 1665 27400 1680
rect 27440 1675 27510 1680
rect 27440 1665 27455 1675
rect 27495 1665 27510 1675
rect 27550 1665 27565 1680
rect 27605 1665 27620 1680
rect 27660 1665 27675 1680
rect 27715 1665 27730 1680
rect 26070 1500 26085 1515
rect 26125 1500 26140 1515
rect 26180 1500 26195 1515
rect 26235 1500 26250 1515
rect 26290 1505 26305 1515
rect 26345 1505 26360 1515
rect 26106 1490 26140 1500
rect 26290 1490 26360 1505
rect 26400 1500 26415 1515
rect 26455 1500 26470 1515
rect 26510 1505 26525 1515
rect 26565 1505 26580 1515
rect 26510 1490 26580 1505
rect 26620 1500 26635 1515
rect 26675 1505 26690 1515
rect 26810 1505 26825 1515
rect 26675 1490 26825 1505
rect 26865 1500 26880 1515
rect 26920 1500 26935 1515
rect 26975 1505 26990 1515
rect 27110 1505 27125 1515
rect 26920 1490 26954 1500
rect 26975 1490 27125 1505
rect 27165 1500 27180 1515
rect 27220 1500 27235 1515
rect 27275 1500 27290 1515
rect 27330 1505 27345 1515
rect 27385 1505 27400 1515
rect 27146 1490 27180 1500
rect 27330 1490 27400 1505
rect 27440 1500 27455 1515
rect 27495 1500 27510 1515
rect 27550 1505 27565 1515
rect 27605 1505 27620 1515
rect 27550 1490 27620 1505
rect 27660 1500 27675 1515
rect 27715 1500 27730 1515
rect 26106 1470 26112 1490
rect 26129 1470 26138 1490
rect 26106 1460 26138 1470
rect 26305 1470 26315 1490
rect 26335 1470 26345 1490
rect 26305 1460 26345 1470
rect 26525 1470 26535 1490
rect 26555 1470 26565 1490
rect 26525 1460 26565 1470
rect 26730 1470 26740 1490
rect 26760 1470 26770 1490
rect 26730 1460 26770 1470
rect 26922 1470 26928 1490
rect 26945 1470 26954 1490
rect 26922 1460 26954 1470
rect 27030 1470 27040 1490
rect 27060 1470 27070 1490
rect 27030 1460 27070 1470
rect 27146 1470 27152 1490
rect 27169 1470 27178 1490
rect 27146 1460 27178 1470
rect 27345 1470 27355 1490
rect 27375 1470 27385 1490
rect 27345 1460 27385 1470
rect 27565 1470 27575 1490
rect 27595 1470 27605 1490
rect 27565 1460 27605 1470
rect 28408 1700 28442 1710
rect 28408 1680 28416 1700
rect 28434 1680 28442 1700
rect 28245 1655 28305 1670
rect 28345 1665 28705 1680
rect 28345 1655 28405 1665
rect 28445 1655 28505 1665
rect 28545 1655 28605 1665
rect 28645 1655 28705 1665
rect 28745 1655 28805 1670
rect 27595 1145 27635 1155
rect 27595 1140 27605 1145
rect 26815 1130 26845 1140
rect 26815 1110 26820 1130
rect 26840 1110 26845 1130
rect 27510 1125 27605 1140
rect 27625 1125 27635 1145
rect 26245 1085 26260 1100
rect 26300 1095 27360 1110
rect 26300 1085 26315 1095
rect 26355 1085 26370 1095
rect 26410 1085 26425 1095
rect 26465 1085 26480 1095
rect 26520 1085 26535 1095
rect 26575 1085 26590 1095
rect 26630 1085 26645 1095
rect 26685 1085 26700 1095
rect 26740 1085 26755 1095
rect 26795 1085 26810 1095
rect 26850 1085 26865 1095
rect 26905 1085 26920 1095
rect 26960 1085 26975 1095
rect 27015 1085 27030 1095
rect 27070 1085 27085 1095
rect 27125 1085 27140 1095
rect 27180 1085 27195 1095
rect 27235 1085 27250 1095
rect 27290 1085 27305 1095
rect 27345 1085 27360 1095
rect 27400 1095 27470 1110
rect 27400 1085 27415 1095
rect 27455 1085 27470 1095
rect 27510 1085 27525 1125
rect 27595 1115 27635 1125
rect 27565 1085 27580 1100
rect 25045 945 25105 955
rect 24965 930 25105 945
rect 25145 940 25205 955
rect 25245 940 25305 955
rect 25345 940 25405 955
rect 25445 940 25505 955
rect 25545 945 25605 955
rect 25545 930 25685 945
rect 24965 910 24975 930
rect 24995 910 25005 930
rect 18845 900 18885 910
rect 24965 900 25005 910
rect 25645 910 25655 930
rect 25675 910 25685 930
rect 25645 900 25685 910
rect 17620 880 17660 890
rect 16305 795 16345 805
rect 3035 765 3085 780
rect 3125 755 3175 780
rect 3215 765 3265 780
rect 3305 765 3355 780
rect 3395 765 3445 780
rect 3485 765 3535 780
rect 3575 765 3625 780
rect 3665 765 3715 780
rect 3755 765 3805 780
rect 3845 765 3895 780
rect 3935 765 3985 780
rect 4025 765 4075 780
rect 4115 765 4165 780
rect 4205 765 4255 780
rect 4295 765 4345 780
rect 4385 765 4435 780
rect 4475 765 4525 780
rect 4565 765 4615 780
rect 4655 765 4705 780
rect 4745 765 4795 780
rect 4835 765 4885 780
rect 4925 765 4975 780
rect 16305 775 16315 795
rect 16335 775 16345 795
rect 16305 765 16345 775
rect 16375 795 16415 805
rect 16375 775 16385 795
rect 16405 775 16415 795
rect 16375 765 16415 775
rect 16445 795 16485 805
rect 16445 775 16455 795
rect 16475 775 16485 795
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 16445 765 16485 775
rect 3125 750 3140 755
rect 3130 735 3140 750
rect 3160 750 3175 755
rect 16300 750 16490 765
rect 16920 760 17485 775
rect 16920 750 16935 760
rect 16975 750 16990 760
rect 17030 750 17045 760
rect 17085 750 17100 760
rect 17140 750 17155 760
rect 17195 750 17210 760
rect 17250 750 17265 760
rect 17305 750 17320 760
rect 17360 750 17375 760
rect 17415 750 17430 760
rect 17470 750 17485 760
rect 17525 750 17540 765
rect 26245 820 26260 835
rect 26300 820 26315 835
rect 26355 820 26370 835
rect 26410 820 26425 835
rect 26465 820 26480 835
rect 26520 820 26535 835
rect 26575 820 26590 835
rect 26630 820 26645 835
rect 26685 820 26700 835
rect 26740 820 26755 835
rect 26795 820 26810 835
rect 26850 820 26865 835
rect 26905 820 26920 835
rect 26960 820 26975 835
rect 27015 820 27030 835
rect 27070 820 27085 835
rect 27125 820 27140 835
rect 27180 820 27195 835
rect 27235 820 27250 835
rect 27290 820 27305 835
rect 27345 820 27360 835
rect 27400 820 27415 835
rect 27455 820 27470 835
rect 27510 820 27525 835
rect 27565 820 27580 835
rect 26195 810 26260 820
rect 26195 790 26205 810
rect 26225 805 26260 810
rect 27565 810 27625 820
rect 27565 805 27595 810
rect 26225 790 26235 805
rect 26195 780 26235 790
rect 27585 790 27595 805
rect 27615 790 27625 810
rect 27585 780 27625 790
rect 28245 940 28305 955
rect 28345 940 28405 955
rect 28445 940 28505 955
rect 28545 940 28605 955
rect 28645 940 28705 955
rect 28745 940 28805 955
rect 3160 735 3170 750
rect 3130 725 3170 735
rect 16920 690 16935 700
rect 16840 675 16935 690
rect 16975 685 16990 700
rect 17030 685 17045 700
rect 17085 685 17100 700
rect 17140 685 17155 700
rect 17195 685 17210 700
rect 17250 685 17265 700
rect 17305 685 17320 700
rect 17360 685 17375 700
rect 17415 685 17430 700
rect 17470 685 17485 700
rect 17525 690 17540 700
rect 17525 675 17620 690
rect 16840 655 16850 675
rect 16870 655 16880 675
rect 16300 635 16490 650
rect 16840 645 16880 655
rect 17580 655 17590 675
rect 17610 655 17620 675
rect 17580 645 17620 655
rect 26305 595 26345 605
rect 26305 575 26315 595
rect 26335 575 26345 595
rect 26305 565 26345 575
rect 26375 595 26415 605
rect 26375 575 26385 595
rect 26405 575 26415 595
rect 26375 565 26415 575
rect 26445 595 26485 605
rect 26445 575 26455 595
rect 26475 575 26485 595
rect 26445 565 26485 575
rect 26300 550 26490 565
rect 26300 435 26490 450
rect 26935 595 26975 605
rect 26935 575 26945 595
rect 26965 575 26975 595
rect 27155 595 27195 605
rect 27155 575 27165 595
rect 27185 575 27195 595
rect 27375 595 27415 605
rect 27375 575 27385 595
rect 27405 575 27415 595
rect 26920 560 27485 575
rect 26920 550 26935 560
rect 26975 550 26990 560
rect 27030 550 27045 560
rect 27085 550 27100 560
rect 27140 550 27155 560
rect 27195 550 27210 560
rect 27250 550 27265 560
rect 27305 550 27320 560
rect 27360 550 27375 560
rect 27415 550 27430 560
rect 27470 550 27485 560
rect 27525 550 27540 565
rect 26920 485 26935 500
rect 26975 485 26990 500
rect 27030 485 27045 500
rect 27085 485 27100 500
rect 27140 485 27155 500
rect 27195 485 27210 500
rect 27250 485 27265 500
rect 27305 485 27320 500
rect 27360 485 27375 500
rect 27415 485 27430 500
rect 27470 485 27485 500
rect 27525 485 27540 500
<< polycont >>
rect 26875 4900 26895 4920
rect 26355 4750 26375 4770
rect 26695 4745 26715 4765
rect 27366 4745 27384 4765
rect 16605 4440 16625 4460
rect 16725 4440 16745 4460
rect 16845 4440 16865 4460
rect 16175 4380 16195 4400
rect 16435 4380 16455 4400
rect 16545 4395 16565 4415
rect 16905 4395 16925 4415
rect 26370 4335 26390 4355
rect 16305 4245 16325 4265
rect 16725 4240 16745 4260
rect 17316 4240 17334 4260
rect 16220 4130 16240 4150
rect 17510 4130 17530 4150
rect 26285 4045 26305 4065
rect 26485 4045 26505 4065
rect 27013 4045 27033 4065
rect 27215 4045 27235 4065
rect 27435 4045 27455 4065
rect 16370 4010 16390 4030
rect 26413 3925 26430 3945
rect 26633 3925 26650 3945
rect 26780 3925 26797 3945
rect 27143 3925 27160 3945
rect 27363 3925 27380 3945
rect 27510 3925 27527 3945
rect 16165 3825 16185 3845
rect 16277 3825 16294 3845
rect 16480 3825 16500 3845
rect 16700 3825 16720 3845
rect 16905 3825 16925 3845
rect 17017 3825 17034 3845
rect 17220 3825 17240 3845
rect 17440 3825 17460 3845
rect 17645 3825 17665 3845
rect 16408 3705 16425 3725
rect 16628 3705 16645 3725
rect 16775 3705 16792 3725
rect 17148 3705 17165 3725
rect 17368 3705 17385 3725
rect 17515 3705 17532 3725
rect 3145 2955 3165 2975
rect 4845 2955 4865 2975
rect 16190 3550 16210 3570
rect 17590 3550 17610 3570
rect 16831 3080 16849 3100
rect 14975 2940 14995 2960
rect 15511 2940 15529 2960
rect 15715 2940 15735 2960
rect 18115 2940 18135 2960
rect 18321 2940 18339 2960
rect 18855 2940 18875 2960
rect 26831 3160 26849 3180
rect 28321 3020 28339 3040
rect 24975 2940 24995 2960
rect 25511 2940 25529 2960
rect 25715 2940 25735 2960
rect 15985 2870 16005 2890
rect 16785 2870 16805 2890
rect 16995 2870 17015 2890
rect 17795 2870 17815 2890
rect 25985 2870 26005 2890
rect 26785 2870 26805 2890
rect 3005 2785 3025 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 4805 2725 4825 2745
rect 3365 2350 3385 2370
rect 3895 2355 3915 2375
rect 16386 2450 16404 2470
rect 17396 2450 17414 2470
rect 14975 2410 14995 2430
rect 15715 2410 15735 2430
rect 18115 2410 18135 2430
rect 18855 2410 18875 2430
rect 15595 2350 15615 2370
rect 18235 2350 18255 2370
rect 14975 2290 14995 2310
rect 15715 2290 15735 2310
rect 18115 2290 18135 2310
rect 18855 2290 18875 2310
rect 16836 2155 16854 2175
rect 26386 2450 26404 2470
rect 24975 2410 24995 2430
rect 25715 2410 25735 2430
rect 27406 2450 27424 2470
rect 28321 2460 28339 2480
rect 25595 2350 25615 2370
rect 24975 2290 24995 2310
rect 25715 2290 25735 2310
rect 26836 2155 26854 2175
rect 16245 1935 16265 1955
rect 17535 1935 17555 1955
rect 2630 1855 2650 1875
rect 2775 1855 2795 1875
rect 28321 2270 28339 2290
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 3995 1850 4015 1870
rect 4125 1855 4145 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 5215 1855 5235 1875
rect 3235 1735 3255 1755
rect 4755 1735 4775 1755
rect 15416 1680 15434 1700
rect 16243 1690 16260 1710
rect 16463 1690 16480 1710
rect 16610 1690 16627 1710
rect 16876 1690 16893 1710
rect 17283 1690 17300 1710
rect 17503 1690 17520 1710
rect 17650 1690 17667 1710
rect 18416 1680 18434 1700
rect 25416 1680 25434 1700
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 3005 905 3025 925
rect 4985 905 5005 925
rect 16000 1470 16020 1490
rect 16112 1470 16129 1490
rect 16315 1470 16335 1490
rect 16535 1470 16555 1490
rect 16740 1470 16760 1490
rect 16928 1470 16945 1490
rect 17040 1470 17060 1490
rect 17152 1470 17169 1490
rect 17355 1470 17375 1490
rect 17575 1470 17595 1490
rect 17780 1470 17800 1490
rect 16820 1210 16840 1230
rect 17605 1225 17625 1245
rect 14975 910 14995 930
rect 15655 910 15675 930
rect 16175 890 16195 910
rect 17630 890 17650 910
rect 18175 910 18195 930
rect 18855 910 18875 930
rect 26243 1690 26260 1710
rect 26463 1690 26480 1710
rect 26610 1690 26627 1710
rect 26876 1690 26893 1710
rect 27283 1690 27300 1710
rect 27503 1690 27520 1710
rect 27650 1690 27667 1710
rect 26112 1470 26129 1490
rect 26315 1470 26335 1490
rect 26535 1470 26555 1490
rect 26740 1470 26760 1490
rect 26928 1470 26945 1490
rect 27040 1470 27060 1490
rect 27152 1470 27169 1490
rect 27355 1470 27375 1490
rect 27575 1470 27595 1490
rect 28416 1680 28434 1700
rect 26820 1110 26840 1130
rect 27605 1125 27625 1145
rect 24975 910 24995 930
rect 25655 910 25675 930
rect 16315 775 16335 795
rect 16385 775 16405 795
rect 16455 775 16475 795
rect 16945 775 16965 795
rect 17165 775 17185 795
rect 17385 775 17405 795
rect 3140 735 3160 755
rect 26205 790 26225 810
rect 27595 790 27615 810
rect 16850 655 16870 675
rect 17590 655 17610 675
rect 26315 575 26335 595
rect 26385 575 26405 595
rect 26455 575 26475 595
rect 26945 575 26965 595
rect 27165 575 27185 595
rect 27385 575 27405 595
<< xpolycontact >>
rect 14554 3300 14695 3520
rect 91 3170 311 3205
rect 925 3170 1145 3205
rect 1306 3165 1526 3200
rect 2110 3165 2330 3200
rect 91 3110 311 3145
rect 925 3110 1145 3145
rect 1306 3105 1526 3140
rect 2110 3105 2330 3140
rect 91 3030 311 3065
rect 895 3030 1115 3065
rect 1306 3045 1526 3080
rect 2110 3045 2330 3080
rect 91 2970 311 3005
rect 895 2970 1115 3005
rect 1306 2985 1526 3020
rect 2110 2985 2330 3020
rect 1306 2925 1526 2960
rect 2110 2925 2330 2960
rect 14554 2940 14695 3160
rect 19105 3300 19246 3520
rect 19105 2940 19246 3160
rect 24554 3300 24695 3520
rect 24554 2940 24695 3160
rect 29105 3400 29246 3620
rect 29105 3040 29246 3260
rect 1306 2865 1526 2900
rect 2110 2865 2330 2900
rect 96 2820 315 2855
rect 504 2820 724 2855
rect 1306 2805 1526 2840
rect 1740 2805 1960 2840
rect 96 2760 315 2795
rect 504 2760 724 2795
rect 14640 2405 14675 2625
rect 14640 2010 14675 2230
rect 14700 2405 14735 2625
rect 14700 2010 14735 2230
rect 14760 2405 14795 2625
rect 14760 2010 14795 2230
rect 14820 2405 14855 2625
rect 18995 2405 19030 2625
rect 14820 2010 14855 2230
rect 18995 2010 19030 2230
rect 19055 2405 19090 2625
rect 19055 2010 19090 2230
rect 19115 2405 19150 2625
rect 19115 2010 19150 2230
rect 19175 2405 19210 2625
rect 19175 2010 19210 2230
rect 24640 2405 24675 2625
rect 24640 2010 24675 2230
rect 24700 2405 24735 2625
rect 24700 2010 24735 2230
rect 24760 2405 24795 2625
rect 24760 2010 24795 2230
rect 24820 2405 24855 2625
rect 24820 2010 24855 2230
rect 29065 2385 29100 2605
rect 29065 1990 29100 2210
rect 29125 2385 29160 2605
rect 29125 1990 29160 2210
rect 29185 2385 29220 2605
rect 29185 1990 29220 2210
rect 29245 2385 29280 2605
rect 29245 1990 29280 2210
rect 14820 1385 14855 1605
rect 14820 910 14855 1130
rect 14880 1385 14915 1605
rect 14880 910 14915 1130
rect 18935 1385 18970 1605
rect 18935 910 18970 1130
rect 18995 1385 19030 1605
rect 18995 910 19030 1130
rect 24820 1385 24855 1605
rect 24820 910 24855 1130
rect 24880 1385 24915 1605
rect 24880 910 24915 1130
rect 29055 1385 29090 1605
rect 29055 910 29090 1130
rect 29115 1385 29150 1605
rect 29115 910 29150 1130
<< ppolyres >>
rect 14554 3160 14695 3300
rect 19105 3160 19246 3300
rect 24554 3160 24695 3300
rect 29105 3260 29246 3400
rect 315 2820 504 2855
rect 315 2760 504 2795
<< xpolyres >>
rect 311 3170 925 3205
rect 1526 3165 2110 3200
rect 311 3110 925 3145
rect 1526 3105 2110 3140
rect 311 3030 895 3065
rect 1526 3045 2110 3080
rect 311 2970 895 3005
rect 1526 2985 2110 3020
rect 1526 2925 2110 2960
rect 1526 2865 2110 2900
rect 1526 2805 1740 2840
rect 14640 2230 14675 2405
rect 14700 2230 14735 2405
rect 14760 2230 14795 2405
rect 14820 2230 14855 2405
rect 18995 2230 19030 2405
rect 19055 2230 19090 2405
rect 19115 2230 19150 2405
rect 19175 2230 19210 2405
rect 24640 2230 24675 2405
rect 24700 2230 24735 2405
rect 24760 2230 24795 2405
rect 24820 2230 24855 2405
rect 29065 2210 29100 2385
rect 29125 2210 29160 2385
rect 29185 2210 29220 2385
rect 29245 2210 29280 2385
rect 14820 1130 14855 1385
rect 14880 1130 14915 1385
rect 18935 1130 18970 1385
rect 18995 1130 19030 1385
rect 24820 1130 24855 1385
rect 24880 1130 24915 1385
rect 29055 1130 29090 1385
rect 29115 1130 29150 1385
<< locali >>
rect 26565 4970 26605 4990
rect 26685 4970 26725 4990
rect 26805 4970 26845 4990
rect 26205 4950 26520 4970
rect 26600 4950 26955 4970
rect 26205 4865 26225 4950
rect 26505 4920 26545 4930
rect 26505 4900 26515 4920
rect 26535 4900 26545 4920
rect 26505 4890 26545 4900
rect 26572 4920 26598 4930
rect 26572 4900 26575 4920
rect 26595 4900 26598 4920
rect 26572 4890 26598 4900
rect 26625 4920 26665 4930
rect 26625 4900 26635 4920
rect 26655 4900 26665 4920
rect 26625 4890 26665 4900
rect 26692 4920 26718 4930
rect 26692 4900 26695 4920
rect 26715 4900 26718 4920
rect 26692 4890 26718 4900
rect 26745 4920 26785 4930
rect 26745 4900 26755 4920
rect 26775 4900 26785 4920
rect 26745 4890 26785 4900
rect 26812 4920 26838 4930
rect 26812 4900 26815 4920
rect 26835 4900 26838 4920
rect 26812 4890 26838 4900
rect 26865 4920 26905 4930
rect 26865 4900 26875 4920
rect 26895 4900 26905 4920
rect 26865 4890 26905 4900
rect 26325 4853 26345 4875
rect 26515 4870 26535 4890
rect 26575 4870 26595 4890
rect 26635 4870 26655 4890
rect 26695 4870 26715 4890
rect 26755 4870 26775 4890
rect 26815 4870 26835 4890
rect 26875 4870 26895 4890
rect 26260 4830 26290 4853
rect 26260 4810 26265 4830
rect 26285 4810 26290 4830
rect 26260 4800 26290 4810
rect 26320 4835 26350 4853
rect 26320 4815 26325 4835
rect 26345 4815 26350 4835
rect 26320 4800 26350 4815
rect 26380 4835 26410 4853
rect 26380 4815 26385 4835
rect 26405 4815 26410 4835
rect 26380 4800 26410 4815
rect 26440 4830 26470 4853
rect 26440 4810 26445 4830
rect 26465 4810 26470 4830
rect 26440 4800 26470 4810
rect 26510 4845 26540 4870
rect 26510 4825 26515 4845
rect 26535 4825 26540 4845
rect 26510 4800 26540 4825
rect 26570 4845 26600 4870
rect 26570 4825 26575 4845
rect 26595 4825 26600 4845
rect 26570 4800 26600 4825
rect 26630 4845 26660 4870
rect 26630 4825 26635 4845
rect 26655 4825 26660 4845
rect 26630 4800 26660 4825
rect 26690 4845 26720 4870
rect 26690 4825 26695 4845
rect 26715 4825 26720 4845
rect 26690 4800 26720 4825
rect 26750 4845 26780 4870
rect 26750 4825 26755 4845
rect 26775 4825 26780 4845
rect 26750 4800 26780 4825
rect 26810 4845 26840 4870
rect 26810 4825 26815 4845
rect 26835 4825 26840 4845
rect 26810 4800 26840 4825
rect 26870 4845 26900 4870
rect 26870 4825 26875 4845
rect 26895 4825 26900 4845
rect 26870 4800 26900 4825
rect 26935 4865 26955 4950
rect 26205 4715 26225 4785
rect 26385 4780 26405 4800
rect 26345 4770 26405 4780
rect 26345 4750 26355 4770
rect 26375 4760 26405 4770
rect 26685 4765 26725 4775
rect 26375 4750 26385 4760
rect 26345 4740 26385 4750
rect 26685 4745 26695 4765
rect 26715 4745 26725 4765
rect 26685 4735 26725 4745
rect 26935 4715 26955 4785
rect 26205 4695 26520 4715
rect 26600 4695 26955 4715
rect 27185 4925 27460 4945
rect 27540 4925 27805 4945
rect 27185 4860 27205 4925
rect 27235 4895 27275 4905
rect 27235 4875 27245 4895
rect 27265 4875 27275 4895
rect 27235 4865 27275 4875
rect 27355 4895 27395 4905
rect 27355 4875 27365 4895
rect 27385 4875 27395 4895
rect 27355 4865 27395 4875
rect 27475 4895 27515 4905
rect 27475 4875 27485 4895
rect 27505 4875 27515 4895
rect 27475 4865 27515 4875
rect 27595 4895 27635 4905
rect 27595 4875 27605 4895
rect 27625 4875 27635 4895
rect 27595 4865 27635 4875
rect 27715 4895 27755 4905
rect 27715 4875 27725 4895
rect 27745 4875 27755 4895
rect 27715 4865 27755 4875
rect 27785 4865 27805 4925
rect 27245 4845 27265 4865
rect 27365 4845 27385 4865
rect 27485 4845 27505 4865
rect 27605 4845 27625 4865
rect 27725 4845 27745 4865
rect 27240 4830 27270 4845
rect 27240 4810 27245 4830
rect 27265 4810 27270 4830
rect 27240 4795 27270 4810
rect 27300 4830 27330 4845
rect 27300 4810 27305 4830
rect 27325 4810 27330 4830
rect 27300 4795 27330 4810
rect 27360 4830 27390 4845
rect 27360 4810 27365 4830
rect 27385 4810 27390 4830
rect 27360 4795 27390 4810
rect 27420 4830 27450 4845
rect 27420 4810 27425 4830
rect 27445 4810 27450 4830
rect 27420 4795 27450 4810
rect 27480 4830 27510 4845
rect 27480 4810 27485 4830
rect 27505 4810 27510 4830
rect 27480 4795 27510 4810
rect 27540 4830 27570 4845
rect 27540 4810 27545 4830
rect 27565 4810 27570 4830
rect 27540 4795 27570 4810
rect 27600 4830 27630 4845
rect 27600 4810 27605 4830
rect 27625 4810 27630 4830
rect 27600 4795 27630 4810
rect 27660 4830 27690 4845
rect 27660 4810 27665 4830
rect 27685 4810 27690 4830
rect 27660 4795 27690 4810
rect 27720 4830 27750 4845
rect 27720 4810 27725 4830
rect 27745 4810 27750 4830
rect 27720 4795 27750 4810
rect 27185 4715 27205 4780
rect 27305 4775 27325 4795
rect 27425 4775 27445 4795
rect 27545 4775 27565 4795
rect 27665 4775 27685 4795
rect 27295 4765 27335 4775
rect 27295 4745 27305 4765
rect 27325 4745 27335 4765
rect 27295 4735 27335 4745
rect 27358 4765 27392 4775
rect 27358 4745 27366 4765
rect 27384 4745 27392 4765
rect 27358 4735 27392 4745
rect 27415 4765 27455 4775
rect 27415 4745 27425 4765
rect 27445 4745 27455 4765
rect 27415 4735 27455 4745
rect 27535 4765 27575 4775
rect 27535 4745 27545 4765
rect 27565 4745 27575 4765
rect 27535 4735 27575 4745
rect 27655 4765 27695 4775
rect 27655 4745 27665 4765
rect 27685 4745 27695 4765
rect 27655 4735 27695 4745
rect 27785 4715 27805 4780
rect 27185 4695 27460 4715
rect 27540 4695 27805 4715
rect 26200 4505 26835 4525
rect 26915 4505 27550 4525
rect 16597 4460 16633 4470
rect 16597 4440 16605 4460
rect 16625 4440 16633 4460
rect 16597 4430 16633 4440
rect 16717 4460 16753 4470
rect 16717 4440 16725 4460
rect 16745 4440 16753 4460
rect 16717 4430 16753 4440
rect 16837 4460 16873 4470
rect 16837 4440 16845 4460
rect 16865 4440 16873 4460
rect 16837 4430 16873 4440
rect 26200 4445 26220 4505
rect 26360 4475 26400 4485
rect 26360 4455 26370 4475
rect 26390 4455 26400 4475
rect 26360 4445 26400 4455
rect 26470 4475 26510 4485
rect 26470 4455 26480 4475
rect 26500 4455 26510 4475
rect 26470 4445 26510 4455
rect 26580 4475 26620 4485
rect 26580 4455 26590 4475
rect 26610 4455 26620 4475
rect 26580 4445 26620 4455
rect 26690 4475 26730 4485
rect 26690 4455 26700 4475
rect 26720 4455 26730 4475
rect 26690 4445 26730 4455
rect 26800 4475 26840 4485
rect 26800 4455 26810 4475
rect 26830 4455 26840 4475
rect 26800 4445 26840 4455
rect 26910 4475 26950 4485
rect 26910 4455 26920 4475
rect 26940 4455 26950 4475
rect 26910 4445 26950 4455
rect 27020 4475 27060 4485
rect 27020 4455 27030 4475
rect 27050 4455 27060 4475
rect 27020 4445 27060 4455
rect 27130 4475 27170 4485
rect 27130 4455 27140 4475
rect 27160 4455 27170 4475
rect 27130 4445 27170 4455
rect 27240 4475 27280 4485
rect 27240 4455 27250 4475
rect 27270 4455 27280 4475
rect 27240 4445 27280 4455
rect 27350 4475 27390 4485
rect 27350 4455 27360 4475
rect 27380 4455 27390 4475
rect 27350 4445 27390 4455
rect 27530 4445 27550 4505
rect 16535 4415 16575 4425
rect 16165 4400 16205 4410
rect 16165 4380 16175 4400
rect 16195 4380 16205 4400
rect 16165 4370 16205 4380
rect 16425 4400 16465 4410
rect 16425 4380 16435 4400
rect 16455 4380 16465 4400
rect 16535 4395 16545 4415
rect 16565 4395 16575 4415
rect 16535 4385 16575 4395
rect 16425 4370 16465 4380
rect 16175 4348 16195 4370
rect 16435 4348 16455 4370
rect 16545 4365 16565 4385
rect 16605 4365 16625 4430
rect 16655 4415 16695 4425
rect 16655 4395 16665 4415
rect 16685 4395 16695 4415
rect 16655 4385 16695 4395
rect 16665 4365 16685 4385
rect 16725 4365 16745 4430
rect 16775 4415 16815 4425
rect 16775 4395 16785 4415
rect 16805 4395 16815 4415
rect 16775 4385 16815 4395
rect 16785 4365 16805 4385
rect 16845 4365 16865 4430
rect 16895 4415 16935 4425
rect 16895 4395 16905 4415
rect 16925 4395 16935 4415
rect 16895 4385 16935 4395
rect 17185 4390 17225 4400
rect 16905 4365 16925 4385
rect 17185 4370 17195 4390
rect 17215 4370 17225 4390
rect 16170 4325 16240 4348
rect 16170 4305 16175 4325
rect 16195 4305 16215 4325
rect 16235 4305 16240 4325
rect 16170 4295 16240 4305
rect 16270 4330 16300 4348
rect 16270 4310 16275 4330
rect 16295 4310 16300 4330
rect 16270 4295 16300 4310
rect 16330 4330 16360 4348
rect 16330 4310 16335 4330
rect 16355 4310 16360 4330
rect 16330 4295 16360 4310
rect 16390 4325 16460 4348
rect 16390 4305 16395 4325
rect 16415 4305 16435 4325
rect 16455 4305 16460 4325
rect 16390 4295 16460 4305
rect 16500 4340 16570 4365
rect 16500 4320 16505 4340
rect 16525 4320 16545 4340
rect 16565 4320 16570 4340
rect 16500 4295 16570 4320
rect 16600 4340 16630 4365
rect 16600 4320 16605 4340
rect 16625 4320 16630 4340
rect 16600 4295 16630 4320
rect 16660 4340 16690 4365
rect 16660 4320 16665 4340
rect 16685 4320 16690 4340
rect 16660 4295 16690 4320
rect 16720 4340 16750 4365
rect 16720 4320 16725 4340
rect 16745 4320 16750 4340
rect 16720 4295 16750 4320
rect 16780 4340 16810 4365
rect 16780 4320 16785 4340
rect 16805 4320 16810 4340
rect 16780 4295 16810 4320
rect 16840 4340 16870 4365
rect 16840 4320 16845 4340
rect 16865 4320 16870 4340
rect 16840 4295 16870 4320
rect 16900 4340 16970 4365
rect 17185 4360 17225 4370
rect 17305 4390 17345 4400
rect 17305 4370 17315 4390
rect 17335 4370 17345 4390
rect 17305 4360 17345 4370
rect 17425 4390 17465 4400
rect 17425 4370 17435 4390
rect 17455 4370 17465 4390
rect 17425 4360 17465 4370
rect 17545 4390 17585 4400
rect 17545 4370 17555 4390
rect 17575 4370 17585 4390
rect 17545 4360 17585 4370
rect 17665 4390 17705 4400
rect 17665 4370 17675 4390
rect 17695 4370 17705 4390
rect 17665 4360 17705 4370
rect 26370 4425 26390 4445
rect 26480 4425 26500 4445
rect 26590 4425 26610 4445
rect 26700 4425 26720 4445
rect 26810 4425 26830 4445
rect 26920 4425 26940 4445
rect 27030 4425 27050 4445
rect 27140 4425 27160 4445
rect 27250 4425 27270 4445
rect 27360 4425 27380 4445
rect 26255 4415 26285 4425
rect 26255 4395 26260 4415
rect 26280 4395 26285 4415
rect 26255 4385 26285 4395
rect 26310 4415 26340 4425
rect 26310 4395 26315 4415
rect 26335 4395 26340 4415
rect 26310 4385 26340 4395
rect 26365 4415 26395 4425
rect 26365 4395 26370 4415
rect 26390 4395 26395 4415
rect 26365 4385 26395 4395
rect 26420 4415 26450 4425
rect 26420 4395 26425 4415
rect 26445 4395 26450 4415
rect 26420 4385 26450 4395
rect 26475 4415 26505 4425
rect 26475 4395 26480 4415
rect 26500 4395 26505 4415
rect 26475 4385 26505 4395
rect 26530 4415 26560 4425
rect 26530 4395 26535 4415
rect 26555 4395 26560 4415
rect 26530 4385 26560 4395
rect 26585 4415 26615 4425
rect 26585 4395 26590 4415
rect 26610 4395 26615 4415
rect 26585 4385 26615 4395
rect 26640 4415 26670 4425
rect 26640 4395 26645 4415
rect 26665 4395 26670 4415
rect 26640 4385 26670 4395
rect 26695 4415 26725 4425
rect 26695 4395 26700 4415
rect 26720 4395 26725 4415
rect 26695 4385 26725 4395
rect 26750 4415 26780 4425
rect 26750 4395 26755 4415
rect 26775 4395 26780 4415
rect 26750 4385 26780 4395
rect 26805 4415 26835 4425
rect 26805 4395 26810 4415
rect 26830 4395 26835 4415
rect 26805 4385 26835 4395
rect 26860 4415 26890 4425
rect 26860 4395 26865 4415
rect 26885 4395 26890 4415
rect 26860 4385 26890 4395
rect 26915 4415 26945 4425
rect 26915 4395 26920 4415
rect 26940 4395 26945 4415
rect 26915 4385 26945 4395
rect 26970 4415 27000 4425
rect 26970 4395 26975 4415
rect 26995 4395 27000 4415
rect 26970 4385 27000 4395
rect 27025 4415 27055 4425
rect 27025 4395 27030 4415
rect 27050 4395 27055 4415
rect 27025 4385 27055 4395
rect 27080 4415 27110 4425
rect 27080 4395 27085 4415
rect 27105 4395 27110 4415
rect 27080 4385 27110 4395
rect 27135 4415 27165 4425
rect 27135 4395 27140 4415
rect 27160 4395 27165 4415
rect 27135 4385 27165 4395
rect 27190 4415 27220 4425
rect 27190 4395 27195 4415
rect 27215 4395 27220 4415
rect 27190 4385 27220 4395
rect 27245 4415 27275 4425
rect 27245 4395 27250 4415
rect 27270 4395 27275 4415
rect 27245 4385 27275 4395
rect 27300 4415 27330 4425
rect 27300 4395 27305 4415
rect 27325 4395 27330 4415
rect 27300 4385 27330 4395
rect 27355 4415 27385 4425
rect 27355 4395 27360 4415
rect 27380 4395 27385 4415
rect 27355 4385 27385 4395
rect 27410 4415 27440 4425
rect 27410 4395 27415 4415
rect 27435 4395 27440 4415
rect 27410 4385 27440 4395
rect 27465 4415 27495 4425
rect 27465 4395 27470 4415
rect 27490 4395 27495 4415
rect 27465 4385 27495 4395
rect 26315 4365 26335 4385
rect 26425 4365 26445 4385
rect 26535 4365 26555 4385
rect 26645 4365 26665 4385
rect 26755 4365 26775 4385
rect 26865 4365 26885 4385
rect 26975 4365 26995 4385
rect 27085 4365 27105 4385
rect 27195 4365 27215 4385
rect 27305 4365 27325 4385
rect 27415 4365 27435 4385
rect 17195 4340 17215 4360
rect 17315 4340 17335 4360
rect 17435 4340 17455 4360
rect 17555 4340 17575 4360
rect 17675 4340 17695 4360
rect 16900 4320 16905 4340
rect 16925 4320 16945 4340
rect 16965 4320 16970 4340
rect 16900 4295 16970 4320
rect 17150 4325 17220 4340
rect 17150 4305 17155 4325
rect 17175 4305 17195 4325
rect 17215 4305 17220 4325
rect 16335 4275 16355 4295
rect 17150 4290 17220 4305
rect 17250 4325 17280 4340
rect 17250 4305 17255 4325
rect 17275 4305 17280 4325
rect 17250 4290 17280 4305
rect 17310 4325 17340 4340
rect 17310 4305 17315 4325
rect 17335 4305 17340 4325
rect 17310 4290 17340 4305
rect 17370 4325 17400 4340
rect 17370 4305 17375 4325
rect 17395 4305 17400 4325
rect 17370 4290 17400 4305
rect 17430 4325 17460 4340
rect 17430 4305 17435 4325
rect 17455 4305 17460 4325
rect 17430 4290 17460 4305
rect 17490 4325 17520 4340
rect 17490 4305 17495 4325
rect 17515 4305 17520 4325
rect 17490 4290 17520 4305
rect 17550 4325 17580 4340
rect 17550 4305 17555 4325
rect 17575 4305 17580 4325
rect 17550 4290 17580 4305
rect 17610 4325 17640 4340
rect 17610 4305 17615 4325
rect 17635 4305 17640 4325
rect 17610 4290 17640 4305
rect 17670 4325 17740 4340
rect 17670 4305 17675 4325
rect 17695 4305 17715 4325
rect 17735 4305 17740 4325
rect 17670 4290 17740 4305
rect 26200 4305 26220 4365
rect 26305 4355 26345 4365
rect 26305 4335 26315 4355
rect 26335 4335 26345 4355
rect 26305 4325 26345 4335
rect 26362 4355 26398 4365
rect 26362 4335 26370 4355
rect 26390 4335 26398 4355
rect 26362 4325 26398 4335
rect 26415 4355 26455 4365
rect 26415 4335 26425 4355
rect 26445 4335 26455 4355
rect 26415 4325 26455 4335
rect 26525 4355 26565 4365
rect 26525 4335 26535 4355
rect 26555 4335 26565 4355
rect 26525 4325 26565 4335
rect 26635 4355 26675 4365
rect 26635 4335 26645 4355
rect 26665 4335 26675 4355
rect 26635 4325 26675 4335
rect 26745 4355 26785 4365
rect 26745 4335 26755 4355
rect 26775 4335 26785 4355
rect 26745 4325 26785 4335
rect 26855 4355 26895 4365
rect 26855 4335 26865 4355
rect 26885 4335 26895 4355
rect 26855 4325 26895 4335
rect 26965 4355 27005 4365
rect 26965 4335 26975 4355
rect 26995 4335 27005 4355
rect 26965 4325 27005 4335
rect 27075 4355 27115 4365
rect 27075 4335 27085 4355
rect 27105 4335 27115 4355
rect 27075 4325 27115 4335
rect 27185 4355 27225 4365
rect 27185 4335 27195 4355
rect 27215 4335 27225 4355
rect 27185 4325 27225 4335
rect 27295 4355 27335 4365
rect 27295 4335 27305 4355
rect 27325 4335 27335 4355
rect 27295 4325 27335 4335
rect 27405 4355 27445 4365
rect 27405 4335 27415 4355
rect 27435 4335 27445 4355
rect 27405 4325 27445 4335
rect 27530 4305 27550 4365
rect 16295 4265 16355 4275
rect 17255 4270 17275 4290
rect 17375 4270 17395 4290
rect 17495 4270 17515 4290
rect 17615 4270 17635 4290
rect 26200 4285 26835 4305
rect 26915 4285 27550 4305
rect 16295 4245 16305 4265
rect 16325 4255 16355 4265
rect 16715 4260 16755 4270
rect 16325 4245 16335 4255
rect 16295 4235 16335 4245
rect 16715 4240 16725 4260
rect 16745 4240 16755 4260
rect 16715 4230 16755 4240
rect 17245 4260 17285 4270
rect 17245 4240 17255 4260
rect 17275 4240 17285 4260
rect 17245 4230 17285 4240
rect 17308 4260 17342 4270
rect 17308 4240 17316 4260
rect 17334 4240 17342 4260
rect 17308 4230 17342 4240
rect 17365 4260 17405 4270
rect 17365 4240 17375 4260
rect 17395 4240 17405 4260
rect 17365 4230 17405 4240
rect 17485 4260 17525 4270
rect 17485 4240 17495 4260
rect 17515 4240 17525 4260
rect 17485 4230 17525 4240
rect 17605 4260 17645 4270
rect 17605 4240 17615 4260
rect 17635 4240 17645 4260
rect 17605 4230 17645 4240
rect 26420 4210 26460 4250
rect 26635 4210 26675 4250
rect 26855 4210 26895 4250
rect 27075 4210 27115 4250
rect 27295 4210 27335 4250
rect 16210 4150 16250 4160
rect 16210 4130 16220 4150
rect 16240 4130 16250 4150
rect 16210 4120 16250 4130
rect 16360 4150 16400 4160
rect 16360 4130 16370 4150
rect 16390 4130 16400 4150
rect 16360 4120 16400 4130
rect 16470 4150 16510 4160
rect 16470 4130 16480 4150
rect 16500 4130 16510 4150
rect 16470 4120 16510 4130
rect 16580 4150 16620 4160
rect 16580 4130 16590 4150
rect 16610 4130 16620 4150
rect 16580 4120 16620 4130
rect 16690 4150 16730 4160
rect 16690 4130 16700 4150
rect 16720 4130 16730 4150
rect 16690 4120 16730 4130
rect 16800 4150 16840 4160
rect 16800 4130 16810 4150
rect 16830 4130 16840 4150
rect 16800 4120 16840 4130
rect 16910 4150 16950 4160
rect 16910 4130 16920 4150
rect 16940 4130 16950 4150
rect 16910 4120 16950 4130
rect 17020 4150 17060 4160
rect 17020 4130 17030 4150
rect 17050 4130 17060 4150
rect 17020 4120 17060 4130
rect 17130 4150 17170 4160
rect 17130 4130 17140 4150
rect 17160 4130 17170 4150
rect 17130 4120 17170 4130
rect 17240 4150 17280 4160
rect 17240 4130 17250 4150
rect 17270 4130 17280 4150
rect 17240 4120 17280 4130
rect 17350 4150 17390 4160
rect 17350 4130 17360 4150
rect 17380 4130 17390 4150
rect 17350 4120 17390 4130
rect 17500 4150 17540 4160
rect 17500 4130 17510 4150
rect 17530 4130 17540 4150
rect 17500 4120 17540 4130
rect 16220 4100 16240 4120
rect 16370 4100 16390 4120
rect 16480 4100 16500 4120
rect 16590 4100 16610 4120
rect 16700 4100 16720 4120
rect 16810 4100 16830 4120
rect 16920 4100 16940 4120
rect 17030 4100 17050 4120
rect 17140 4100 17160 4120
rect 17250 4100 17270 4120
rect 17360 4100 17380 4120
rect 17510 4100 17530 4120
rect 26325 4115 26355 4130
rect 26425 4115 26455 4130
rect 26535 4115 26565 4130
rect 26645 4115 26675 4130
rect 26755 4115 26785 4130
rect 27055 4115 27085 4130
rect 27155 4115 27185 4130
rect 27265 4115 27295 4130
rect 27375 4115 27405 4130
rect 27485 4115 27515 4130
rect 16215 4090 16285 4100
rect 16215 4070 16220 4090
rect 16240 4070 16260 4090
rect 16280 4070 16285 4090
rect 16215 4060 16285 4070
rect 16310 4090 16340 4100
rect 16310 4070 16315 4090
rect 16335 4070 16340 4090
rect 16310 4060 16340 4070
rect 16365 4090 16395 4100
rect 16365 4070 16370 4090
rect 16390 4070 16395 4090
rect 16365 4060 16395 4070
rect 16420 4090 16450 4100
rect 16420 4070 16425 4090
rect 16445 4070 16450 4090
rect 16420 4060 16450 4070
rect 16475 4090 16505 4100
rect 16475 4070 16480 4090
rect 16500 4070 16505 4090
rect 16475 4060 16505 4070
rect 16530 4090 16560 4100
rect 16530 4070 16535 4090
rect 16555 4070 16560 4090
rect 16530 4060 16560 4070
rect 16585 4090 16615 4100
rect 16585 4070 16590 4090
rect 16610 4070 16615 4090
rect 16585 4060 16615 4070
rect 16640 4090 16670 4100
rect 16640 4070 16645 4090
rect 16665 4070 16670 4090
rect 16640 4060 16670 4070
rect 16695 4090 16725 4100
rect 16695 4070 16700 4090
rect 16720 4070 16725 4090
rect 16695 4060 16725 4070
rect 16750 4090 16780 4100
rect 16750 4070 16755 4090
rect 16775 4070 16780 4090
rect 16750 4060 16780 4070
rect 16805 4090 16835 4100
rect 16805 4070 16810 4090
rect 16830 4070 16835 4090
rect 16805 4060 16835 4070
rect 16860 4090 16890 4100
rect 16860 4070 16865 4090
rect 16885 4070 16890 4090
rect 16860 4060 16890 4070
rect 16915 4090 16945 4100
rect 16915 4070 16920 4090
rect 16940 4070 16945 4090
rect 16915 4060 16945 4070
rect 16970 4090 17000 4100
rect 16970 4070 16975 4090
rect 16995 4070 17000 4090
rect 16970 4060 17000 4070
rect 17025 4090 17055 4100
rect 17025 4070 17030 4090
rect 17050 4070 17055 4090
rect 17025 4060 17055 4070
rect 17080 4090 17110 4100
rect 17080 4070 17085 4090
rect 17105 4070 17110 4090
rect 17080 4060 17110 4070
rect 17135 4090 17165 4100
rect 17135 4070 17140 4090
rect 17160 4070 17165 4090
rect 17135 4060 17165 4070
rect 17190 4090 17220 4100
rect 17190 4070 17195 4090
rect 17215 4070 17220 4090
rect 17190 4060 17220 4070
rect 17245 4090 17275 4100
rect 17245 4070 17250 4090
rect 17270 4070 17275 4090
rect 17245 4060 17275 4070
rect 17300 4090 17330 4100
rect 17300 4070 17305 4090
rect 17325 4070 17330 4090
rect 17300 4060 17330 4070
rect 17355 4090 17385 4100
rect 17355 4070 17360 4090
rect 17380 4070 17385 4090
rect 17355 4060 17385 4070
rect 17410 4090 17440 4100
rect 17410 4070 17415 4090
rect 17435 4070 17440 4090
rect 17410 4060 17440 4070
rect 17465 4090 17535 4100
rect 17465 4070 17470 4090
rect 17490 4070 17510 4090
rect 17530 4070 17535 4090
rect 17465 4060 17535 4070
rect 26150 4095 26875 4115
rect 26955 4095 27680 4115
rect 16315 4040 16335 4060
rect 16425 4040 16445 4060
rect 16535 4040 16555 4060
rect 16645 4040 16665 4060
rect 16755 4040 16775 4060
rect 16865 4040 16885 4060
rect 16975 4040 16995 4060
rect 17085 4040 17105 4060
rect 17195 4040 17215 4060
rect 17305 4040 17325 4060
rect 17415 4040 17435 4060
rect 16305 4030 16345 4040
rect 16305 4010 16315 4030
rect 16335 4010 16345 4030
rect 16305 4000 16345 4010
rect 16362 4030 16398 4040
rect 16362 4010 16370 4030
rect 16390 4010 16398 4030
rect 16362 4000 16398 4010
rect 16415 4030 16455 4040
rect 16415 4010 16425 4030
rect 16445 4010 16455 4030
rect 16415 4000 16455 4010
rect 16525 4030 16565 4040
rect 16525 4010 16535 4030
rect 16555 4010 16565 4030
rect 16525 4000 16565 4010
rect 16635 4030 16675 4040
rect 16635 4010 16645 4030
rect 16665 4010 16675 4030
rect 16635 4000 16675 4010
rect 16745 4030 16785 4040
rect 16745 4010 16755 4030
rect 16775 4010 16785 4030
rect 16745 4000 16785 4010
rect 16855 4030 16895 4040
rect 16855 4010 16865 4030
rect 16885 4010 16895 4030
rect 16855 4000 16895 4010
rect 16965 4030 17005 4040
rect 16965 4010 16975 4030
rect 16995 4010 17005 4030
rect 16965 4000 17005 4010
rect 17075 4030 17115 4040
rect 17075 4010 17085 4030
rect 17105 4010 17115 4030
rect 17075 4000 17115 4010
rect 17185 4030 17225 4040
rect 17185 4010 17195 4030
rect 17215 4010 17225 4030
rect 17185 4000 17225 4010
rect 17295 4030 17335 4040
rect 17295 4010 17305 4030
rect 17325 4010 17335 4030
rect 17295 4000 17335 4010
rect 17405 4030 17445 4040
rect 17405 4010 17415 4030
rect 17435 4010 17445 4030
rect 17405 4000 17445 4010
rect 26150 4035 26170 4095
rect 26280 4065 26310 4075
rect 26280 4045 26285 4065
rect 26305 4045 26310 4065
rect 26280 4035 26310 4045
rect 26327 4065 26353 4075
rect 26327 4045 26330 4065
rect 26350 4045 26353 4065
rect 26327 4035 26353 4045
rect 26370 4065 26400 4075
rect 26370 4045 26375 4065
rect 26395 4045 26400 4065
rect 26370 4035 26400 4045
rect 26427 4065 26453 4075
rect 26427 4045 26430 4065
rect 26450 4045 26453 4065
rect 26427 4035 26453 4045
rect 26480 4065 26510 4075
rect 26480 4045 26485 4065
rect 26505 4045 26510 4065
rect 26480 4035 26510 4045
rect 26537 4065 26563 4075
rect 26537 4045 26540 4065
rect 26560 4045 26563 4065
rect 26537 4035 26563 4045
rect 26647 4065 26673 4075
rect 26647 4045 26650 4065
rect 26670 4045 26673 4065
rect 26647 4035 26673 4045
rect 26757 4065 26783 4075
rect 26757 4045 26760 4065
rect 26780 4045 26783 4065
rect 26757 4035 26783 4045
rect 27008 4065 27038 4075
rect 27008 4045 27013 4065
rect 27033 4045 27038 4065
rect 27008 4035 27038 4045
rect 27057 4065 27083 4075
rect 27057 4045 27060 4065
rect 27080 4045 27083 4065
rect 27057 4035 27083 4045
rect 27157 4065 27183 4075
rect 27157 4045 27160 4065
rect 27180 4045 27183 4065
rect 27157 4035 27183 4045
rect 27205 4065 27245 4075
rect 27205 4045 27215 4065
rect 27235 4045 27245 4065
rect 27205 4035 27245 4045
rect 27267 4065 27293 4075
rect 27267 4045 27270 4065
rect 27290 4045 27293 4065
rect 27267 4035 27293 4045
rect 27377 4065 27403 4075
rect 27377 4045 27380 4065
rect 27400 4045 27403 4065
rect 27377 4035 27403 4045
rect 27425 4065 27465 4075
rect 27425 4045 27435 4065
rect 27455 4045 27465 4065
rect 27425 4035 27465 4045
rect 27487 4065 27513 4075
rect 27487 4045 27490 4065
rect 27510 4045 27513 4065
rect 27487 4035 27513 4045
rect 27660 4035 27680 4095
rect 27875 4040 27905 4070
rect 16415 3940 16455 3980
rect 16635 3940 16675 3980
rect 16855 3940 16895 3980
rect 17075 3940 17115 3980
rect 17295 3940 17335 3980
rect 26327 4015 26345 4035
rect 26375 4015 26395 4035
rect 26430 4015 26450 4035
rect 26540 4015 26560 4035
rect 26650 4015 26670 4035
rect 26760 4015 26780 4035
rect 27057 4015 27075 4035
rect 27160 4015 27180 4035
rect 27270 4015 27290 4035
rect 27380 4015 27400 4035
rect 27490 4015 27510 4035
rect 26205 4005 26235 4015
rect 26205 3985 26210 4005
rect 26230 3985 26235 4005
rect 26205 3975 26235 3985
rect 26260 4005 26290 4015
rect 26260 3985 26265 4005
rect 26285 3985 26290 4005
rect 26260 3975 26290 3985
rect 26315 4005 26345 4015
rect 26315 3985 26320 4005
rect 26340 3985 26345 4005
rect 26315 3975 26345 3985
rect 26370 4005 26400 4015
rect 26370 3985 26375 4005
rect 26395 3985 26400 4005
rect 26370 3975 26400 3985
rect 26425 4005 26455 4015
rect 26425 3985 26430 4005
rect 26450 3985 26455 4005
rect 26425 3975 26455 3985
rect 26480 4005 26510 4015
rect 26480 3985 26485 4005
rect 26505 3985 26510 4005
rect 26480 3975 26510 3985
rect 26535 4005 26565 4015
rect 26535 3985 26540 4005
rect 26560 3985 26565 4005
rect 26535 3975 26565 3985
rect 26590 4005 26620 4015
rect 26590 3985 26595 4005
rect 26615 3985 26620 4005
rect 26590 3975 26620 3985
rect 26645 4005 26675 4015
rect 26645 3985 26650 4005
rect 26670 3985 26675 4005
rect 26645 3975 26675 3985
rect 26700 4005 26730 4015
rect 26700 3985 26705 4005
rect 26725 3985 26730 4005
rect 26700 3975 26730 3985
rect 26755 4005 26785 4015
rect 26755 3985 26760 4005
rect 26780 3985 26785 4005
rect 26755 3975 26785 3985
rect 26810 4005 26840 4015
rect 26810 3985 26815 4005
rect 26835 3985 26840 4005
rect 26810 3975 26840 3985
rect 26865 4005 26895 4015
rect 26865 3985 26870 4005
rect 26890 3985 26895 4005
rect 26865 3975 26895 3985
rect 26935 4005 26965 4015
rect 26935 3985 26940 4005
rect 26960 3985 26965 4005
rect 26935 3975 26965 3985
rect 26990 4005 27020 4015
rect 26990 3985 26995 4005
rect 27015 3985 27020 4005
rect 26990 3975 27020 3985
rect 27045 4005 27075 4015
rect 27045 3985 27050 4005
rect 27070 3985 27075 4005
rect 27045 3975 27075 3985
rect 27100 4005 27130 4015
rect 27100 3985 27105 4005
rect 27125 3985 27130 4005
rect 27100 3975 27130 3985
rect 27155 4005 27185 4015
rect 27155 3985 27160 4005
rect 27180 3985 27185 4005
rect 27155 3975 27185 3985
rect 27210 4005 27240 4015
rect 27210 3985 27215 4005
rect 27235 3985 27240 4005
rect 27210 3975 27240 3985
rect 27265 4005 27295 4015
rect 27265 3985 27270 4005
rect 27290 3985 27295 4005
rect 27265 3975 27295 3985
rect 27320 4005 27350 4015
rect 27320 3985 27325 4005
rect 27345 3985 27350 4005
rect 27320 3975 27350 3985
rect 27375 4005 27405 4015
rect 27375 3985 27380 4005
rect 27400 3985 27405 4005
rect 27375 3975 27405 3985
rect 27430 4005 27460 4015
rect 27430 3985 27435 4005
rect 27455 3985 27460 4005
rect 27430 3975 27460 3985
rect 27485 4005 27515 4015
rect 27485 3985 27490 4005
rect 27510 3985 27515 4005
rect 27485 3975 27515 3985
rect 27540 4005 27570 4015
rect 27540 3985 27545 4005
rect 27565 3985 27570 4005
rect 27540 3975 27570 3985
rect 27595 4005 27625 4015
rect 27595 3985 27600 4005
rect 27620 3985 27625 4005
rect 27595 3975 27625 3985
rect 26265 3955 26285 3975
rect 26370 3955 26390 3975
rect 26485 3955 26505 3975
rect 26590 3955 26610 3975
rect 26705 3955 26725 3975
rect 26820 3955 26840 3975
rect 26995 3955 27015 3975
rect 27100 3955 27120 3975
rect 27215 3955 27235 3975
rect 27320 3955 27340 3975
rect 27435 3955 27455 3975
rect 27550 3955 27570 3975
rect 16310 3905 16350 3915
rect 16310 3885 16320 3905
rect 16340 3885 16350 3905
rect 16310 3875 16350 3885
rect 16415 3905 16455 3915
rect 16415 3885 16425 3905
rect 16445 3885 16455 3905
rect 16415 3875 16455 3885
rect 16525 3905 16565 3915
rect 16525 3885 16535 3905
rect 16555 3885 16565 3905
rect 16525 3875 16565 3885
rect 16635 3905 16675 3915
rect 16635 3885 16645 3905
rect 16665 3885 16675 3905
rect 16635 3875 16675 3885
rect 16745 3905 16785 3915
rect 16745 3885 16755 3905
rect 16775 3885 16785 3905
rect 16745 3875 16785 3885
rect 17050 3905 17090 3915
rect 17050 3885 17060 3905
rect 17080 3885 17090 3905
rect 17050 3875 17090 3885
rect 17155 3905 17195 3915
rect 17155 3885 17165 3905
rect 17185 3885 17195 3905
rect 17155 3875 17195 3885
rect 17265 3905 17305 3915
rect 17265 3885 17275 3905
rect 17295 3885 17305 3905
rect 17265 3875 17305 3885
rect 17375 3905 17415 3915
rect 17375 3885 17385 3905
rect 17405 3885 17415 3905
rect 17375 3875 17415 3885
rect 17485 3905 17525 3915
rect 17485 3885 17495 3905
rect 17515 3885 17525 3905
rect 17485 3875 17525 3885
rect 26150 3895 26170 3955
rect 26255 3945 26295 3955
rect 26255 3925 26265 3945
rect 26285 3925 26295 3945
rect 26255 3915 26295 3925
rect 26350 3945 26390 3955
rect 26350 3925 26360 3945
rect 26380 3925 26390 3945
rect 26350 3915 26390 3925
rect 26407 3945 26439 3955
rect 26407 3925 26413 3945
rect 26430 3925 26439 3945
rect 26407 3915 26439 3925
rect 26475 3945 26515 3955
rect 26475 3925 26485 3945
rect 26505 3925 26515 3945
rect 26475 3915 26515 3925
rect 26570 3945 26610 3955
rect 26570 3925 26580 3945
rect 26600 3925 26610 3945
rect 26570 3915 26610 3925
rect 26627 3945 26659 3955
rect 26627 3925 26633 3945
rect 26650 3925 26659 3945
rect 26627 3915 26659 3925
rect 26695 3945 26735 3955
rect 26695 3925 26705 3945
rect 26725 3925 26735 3945
rect 26695 3915 26735 3925
rect 26771 3945 26803 3955
rect 26771 3925 26780 3945
rect 26797 3925 26803 3945
rect 26771 3915 26803 3925
rect 26820 3945 26860 3955
rect 26820 3925 26830 3945
rect 26850 3925 26860 3945
rect 26820 3915 26860 3925
rect 26985 3945 27025 3955
rect 26985 3925 26995 3945
rect 27015 3925 27025 3945
rect 26985 3915 27025 3925
rect 27080 3945 27120 3955
rect 27080 3925 27090 3945
rect 27110 3925 27120 3945
rect 27080 3915 27120 3925
rect 27137 3945 27169 3955
rect 27137 3925 27143 3945
rect 27160 3925 27169 3945
rect 27137 3915 27169 3925
rect 27205 3945 27245 3955
rect 27205 3925 27215 3945
rect 27235 3925 27245 3945
rect 27205 3915 27245 3925
rect 27300 3945 27340 3955
rect 27300 3925 27310 3945
rect 27330 3925 27340 3945
rect 27300 3915 27340 3925
rect 27357 3945 27389 3955
rect 27357 3925 27363 3945
rect 27380 3925 27389 3945
rect 27357 3915 27389 3925
rect 27425 3945 27465 3955
rect 27425 3925 27435 3945
rect 27455 3925 27465 3945
rect 27425 3915 27465 3925
rect 27501 3945 27533 3955
rect 27501 3925 27510 3945
rect 27527 3925 27533 3945
rect 27501 3915 27533 3925
rect 27550 3945 27590 3955
rect 27550 3925 27560 3945
rect 27580 3925 27590 3945
rect 27550 3915 27590 3925
rect 27660 3895 27680 3955
rect 26150 3875 26875 3895
rect 26955 3875 27680 3895
rect 16155 3845 16195 3855
rect 16155 3825 16165 3845
rect 16185 3825 16195 3845
rect 16155 3815 16195 3825
rect 16271 3845 16303 3855
rect 16271 3825 16277 3845
rect 16294 3825 16303 3845
rect 16271 3815 16303 3825
rect 16165 3795 16185 3815
rect 16320 3795 16340 3875
rect 16360 3845 16400 3855
rect 16360 3825 16370 3845
rect 16390 3825 16400 3845
rect 16360 3815 16400 3825
rect 16370 3795 16390 3815
rect 16425 3795 16445 3875
rect 16470 3845 16510 3855
rect 16470 3825 16480 3845
rect 16500 3825 16510 3845
rect 16470 3815 16510 3825
rect 16535 3795 16555 3875
rect 16645 3795 16665 3875
rect 16690 3845 16730 3855
rect 16690 3825 16700 3845
rect 16720 3825 16730 3845
rect 16690 3815 16730 3825
rect 16755 3795 16775 3875
rect 16800 3845 16840 3855
rect 16800 3825 16810 3845
rect 16830 3825 16840 3845
rect 16800 3815 16840 3825
rect 16895 3845 16935 3855
rect 16895 3825 16905 3845
rect 16925 3825 16935 3845
rect 16895 3815 16935 3825
rect 17011 3845 17043 3855
rect 17011 3825 17017 3845
rect 17034 3825 17043 3845
rect 17011 3815 17043 3825
rect 16810 3795 16830 3815
rect 16905 3795 16925 3815
rect 17060 3795 17080 3875
rect 17165 3795 17185 3875
rect 17210 3845 17250 3855
rect 17210 3825 17220 3845
rect 17240 3825 17250 3845
rect 17210 3815 17250 3825
rect 17275 3795 17295 3875
rect 17385 3795 17405 3875
rect 17430 3845 17470 3855
rect 17430 3825 17440 3845
rect 17460 3825 17470 3845
rect 17430 3815 17470 3825
rect 17495 3795 17515 3875
rect 26260 3860 26290 3875
rect 26365 3860 26395 3875
rect 26480 3860 26510 3875
rect 26585 3860 26615 3875
rect 26700 3860 26730 3875
rect 26815 3860 26845 3875
rect 26990 3860 27020 3875
rect 27210 3860 27240 3875
rect 27430 3860 27460 3875
rect 17635 3845 17675 3855
rect 17635 3825 17645 3845
rect 17665 3825 17675 3845
rect 17635 3815 17675 3825
rect 17865 3820 17895 3850
rect 17645 3795 17665 3815
rect 27975 3795 28005 3825
rect 16155 3785 16230 3795
rect 16155 3765 16165 3785
rect 16185 3765 16205 3785
rect 16225 3765 16230 3785
rect 16155 3755 16230 3765
rect 16255 3785 16285 3795
rect 16255 3765 16260 3785
rect 16280 3765 16285 3785
rect 16255 3755 16285 3765
rect 16310 3785 16340 3795
rect 16310 3765 16315 3785
rect 16335 3765 16340 3785
rect 16310 3755 16340 3765
rect 16365 3785 16395 3795
rect 16365 3765 16370 3785
rect 16390 3765 16395 3785
rect 16365 3755 16395 3765
rect 16420 3785 16450 3795
rect 16420 3765 16425 3785
rect 16445 3765 16450 3785
rect 16420 3755 16450 3765
rect 16475 3785 16505 3795
rect 16475 3765 16480 3785
rect 16500 3765 16505 3785
rect 16475 3755 16505 3765
rect 16530 3785 16560 3795
rect 16530 3765 16535 3785
rect 16555 3765 16560 3785
rect 16530 3755 16560 3765
rect 16585 3785 16615 3795
rect 16585 3765 16590 3785
rect 16610 3765 16615 3785
rect 16585 3755 16615 3765
rect 16640 3785 16670 3795
rect 16640 3765 16645 3785
rect 16665 3765 16670 3785
rect 16640 3755 16670 3765
rect 16695 3785 16725 3795
rect 16695 3765 16700 3785
rect 16720 3765 16725 3785
rect 16695 3755 16725 3765
rect 16750 3785 16780 3795
rect 16750 3765 16755 3785
rect 16775 3765 16780 3785
rect 16750 3755 16780 3765
rect 16805 3785 16835 3795
rect 16805 3765 16810 3785
rect 16830 3765 16835 3785
rect 16805 3755 16835 3765
rect 16860 3785 16970 3795
rect 16860 3765 16865 3785
rect 16885 3765 16905 3785
rect 16925 3765 16945 3785
rect 16965 3765 16970 3785
rect 16860 3755 16970 3765
rect 16995 3785 17025 3795
rect 16995 3765 17000 3785
rect 17020 3765 17025 3785
rect 16995 3755 17025 3765
rect 17050 3785 17080 3795
rect 17050 3765 17055 3785
rect 17075 3765 17080 3785
rect 17050 3755 17080 3765
rect 17105 3785 17135 3795
rect 17105 3765 17110 3785
rect 17130 3765 17135 3785
rect 17105 3755 17135 3765
rect 17160 3785 17190 3795
rect 17160 3765 17165 3785
rect 17185 3765 17190 3785
rect 17160 3755 17190 3765
rect 17215 3785 17245 3795
rect 17215 3765 17220 3785
rect 17240 3765 17245 3785
rect 17215 3755 17245 3765
rect 17270 3785 17300 3795
rect 17270 3765 17275 3785
rect 17295 3765 17300 3785
rect 17270 3755 17300 3765
rect 17325 3785 17355 3795
rect 17325 3765 17330 3785
rect 17350 3765 17355 3785
rect 17325 3755 17355 3765
rect 17380 3785 17410 3795
rect 17380 3765 17385 3785
rect 17405 3765 17410 3785
rect 17380 3755 17410 3765
rect 17435 3785 17465 3795
rect 17435 3765 17440 3785
rect 17460 3765 17465 3785
rect 17435 3755 17465 3765
rect 17490 3785 17520 3795
rect 17490 3765 17495 3785
rect 17515 3765 17520 3785
rect 17490 3755 17520 3765
rect 17545 3785 17575 3795
rect 17545 3765 17550 3785
rect 17570 3765 17575 3785
rect 17545 3755 17575 3765
rect 17600 3785 17675 3795
rect 17600 3765 17605 3785
rect 17625 3765 17645 3785
rect 17665 3765 17675 3785
rect 17600 3755 17675 3765
rect 16260 3675 16280 3755
rect 16365 3675 16385 3755
rect 16402 3725 16434 3735
rect 16402 3705 16408 3725
rect 16425 3705 16434 3725
rect 16402 3695 16434 3705
rect 16480 3675 16500 3755
rect 16585 3675 16605 3755
rect 16622 3725 16654 3735
rect 16622 3705 16628 3725
rect 16645 3705 16654 3725
rect 16622 3695 16654 3705
rect 16700 3675 16720 3755
rect 16766 3725 16798 3735
rect 16766 3705 16775 3725
rect 16792 3705 16798 3725
rect 16766 3695 16798 3705
rect 16815 3675 16835 3755
rect 17000 3685 17020 3755
rect 16990 3675 17030 3685
rect 16250 3665 16290 3675
rect 16250 3645 16260 3665
rect 16280 3645 16290 3665
rect 14610 3605 14640 3635
rect 15060 3630 15100 3640
rect 15060 3610 15070 3630
rect 15090 3610 15100 3630
rect 15060 3600 15100 3610
rect 15170 3630 15210 3640
rect 15170 3610 15180 3630
rect 15200 3610 15210 3630
rect 15170 3600 15210 3610
rect 15280 3630 15320 3640
rect 15280 3610 15290 3630
rect 15310 3610 15320 3630
rect 15280 3600 15320 3610
rect 15390 3630 15430 3640
rect 15390 3610 15400 3630
rect 15420 3610 15430 3630
rect 15390 3600 15430 3610
rect 15500 3630 15540 3640
rect 15500 3610 15510 3630
rect 15530 3610 15540 3630
rect 15500 3600 15540 3610
rect 15610 3630 15650 3640
rect 16250 3635 16290 3645
rect 16355 3665 16395 3675
rect 16355 3645 16365 3665
rect 16385 3645 16395 3665
rect 16355 3635 16395 3645
rect 16470 3665 16510 3675
rect 16470 3645 16480 3665
rect 16500 3645 16510 3665
rect 16470 3635 16510 3645
rect 16575 3665 16615 3675
rect 16575 3645 16585 3665
rect 16605 3645 16615 3665
rect 16575 3635 16615 3645
rect 16690 3665 16730 3675
rect 16690 3645 16700 3665
rect 16720 3645 16730 3665
rect 16690 3635 16730 3645
rect 16805 3665 16845 3675
rect 16805 3645 16815 3665
rect 16835 3645 16845 3665
rect 16990 3655 17000 3675
rect 17020 3655 17030 3675
rect 16990 3645 17030 3655
rect 16805 3635 16845 3645
rect 17105 3640 17125 3755
rect 17142 3725 17174 3735
rect 17142 3705 17148 3725
rect 17165 3705 17174 3725
rect 17142 3695 17174 3705
rect 17220 3685 17240 3755
rect 17210 3675 17250 3685
rect 17210 3655 17220 3675
rect 17240 3655 17250 3675
rect 17210 3645 17250 3655
rect 17325 3640 17345 3755
rect 17362 3725 17394 3735
rect 17362 3705 17368 3725
rect 17385 3705 17394 3725
rect 17362 3695 17394 3705
rect 17440 3685 17460 3755
rect 17506 3725 17538 3735
rect 17506 3705 17515 3725
rect 17532 3705 17538 3725
rect 17506 3695 17538 3705
rect 17430 3675 17470 3685
rect 17430 3655 17440 3675
rect 17460 3655 17470 3675
rect 17430 3645 17470 3655
rect 17555 3640 17575 3755
rect 27095 3750 27125 3780
rect 27315 3750 27345 3780
rect 27545 3750 27575 3780
rect 27920 3750 27950 3780
rect 28095 3740 28455 3760
rect 28535 3740 28895 3760
rect 26170 3680 26860 3700
rect 26940 3680 27630 3700
rect 17965 3650 17995 3680
rect 15610 3610 15620 3630
rect 15640 3610 15650 3630
rect 15610 3600 15650 3610
rect 17095 3600 17135 3640
rect 17315 3600 17355 3640
rect 17545 3600 17585 3640
rect 17910 3605 17940 3635
rect 18200 3630 18240 3640
rect 18200 3610 18210 3630
rect 18230 3610 18240 3630
rect 18200 3600 18240 3610
rect 18310 3630 18350 3640
rect 18310 3610 18320 3630
rect 18340 3610 18350 3630
rect 18310 3600 18350 3610
rect 18420 3630 18460 3640
rect 18420 3610 18430 3630
rect 18450 3610 18460 3630
rect 18420 3600 18460 3610
rect 18530 3630 18570 3640
rect 18530 3610 18540 3630
rect 18560 3610 18570 3630
rect 18530 3600 18570 3610
rect 18640 3630 18680 3640
rect 18640 3610 18650 3630
rect 18670 3610 18680 3630
rect 18640 3600 18680 3610
rect 18750 3630 18790 3640
rect 18750 3610 18760 3630
rect 18780 3610 18790 3630
rect 18750 3600 18790 3610
rect 19160 3605 19190 3635
rect 24610 3605 24640 3635
rect 25060 3630 25100 3640
rect 25060 3610 25070 3630
rect 25090 3610 25100 3630
rect 25060 3600 25100 3610
rect 25170 3630 25210 3640
rect 25170 3610 25180 3630
rect 25200 3610 25210 3630
rect 25170 3600 25210 3610
rect 25280 3630 25320 3640
rect 25280 3610 25290 3630
rect 25310 3610 25320 3630
rect 25280 3600 25320 3610
rect 25390 3630 25430 3640
rect 25390 3610 25400 3630
rect 25420 3610 25430 3630
rect 25390 3600 25430 3610
rect 25500 3630 25540 3640
rect 25500 3610 25510 3630
rect 25530 3610 25540 3630
rect 25500 3600 25540 3610
rect 25610 3630 25650 3640
rect 25610 3610 25620 3630
rect 25640 3610 25650 3630
rect 25610 3600 25650 3610
rect 15070 3580 15090 3600
rect 15180 3580 15200 3600
rect 15290 3580 15310 3600
rect 15400 3580 15420 3600
rect 15510 3580 15530 3600
rect 15620 3580 15640 3600
rect 18210 3580 18230 3600
rect 18320 3580 18340 3600
rect 18430 3580 18450 3600
rect 18540 3580 18560 3600
rect 18650 3580 18670 3600
rect 18760 3580 18780 3600
rect 25070 3580 25090 3600
rect 25180 3580 25200 3600
rect 25290 3580 25310 3600
rect 25400 3580 25420 3600
rect 25510 3580 25530 3600
rect 25620 3580 25640 3600
rect 14970 3570 15040 3580
rect 1266 3495 1296 3525
rect 14554 3520 14695 3560
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1210 3310 1240 3340
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 5365 3305 5395 3335
rect 14970 3550 14975 3570
rect 14995 3550 15015 3570
rect 15035 3550 15040 3570
rect 14970 3520 15040 3550
rect 14970 3500 14975 3520
rect 14995 3500 15015 3520
rect 15035 3500 15040 3520
rect 14970 3470 15040 3500
rect 14970 3450 14975 3470
rect 14995 3450 15015 3470
rect 15035 3450 15040 3470
rect 14970 3420 15040 3450
rect 14970 3400 14975 3420
rect 14995 3400 15015 3420
rect 15035 3400 15040 3420
rect 14970 3370 15040 3400
rect 14970 3350 14975 3370
rect 14995 3350 15015 3370
rect 15035 3350 15040 3370
rect 14970 3320 15040 3350
rect 14970 3300 14975 3320
rect 14995 3300 15015 3320
rect 15035 3300 15040 3320
rect 1165 3255 1195 3285
rect 4890 3255 4920 3285
rect 5415 3255 5445 3285
rect 14970 3270 15040 3300
rect 14970 3250 14975 3270
rect 14995 3250 15015 3270
rect 15035 3250 15040 3270
rect 2740 3210 2770 3240
rect 14970 3220 15040 3250
rect 46 3200 91 3205
rect 46 3175 56 3200
rect 81 3175 91 3200
rect 46 3170 91 3175
rect 14970 3200 14975 3220
rect 14995 3200 15015 3220
rect 15035 3200 15040 3220
rect 1110 3145 1145 3170
rect 1261 3195 1306 3200
rect 1261 3170 1271 3195
rect 1296 3170 1306 3195
rect 1261 3165 1306 3170
rect 2330 3165 2370 3200
rect 46 3140 91 3145
rect 46 3115 56 3140
rect 81 3115 91 3140
rect 46 3110 91 3115
rect 1261 3135 1306 3140
rect 1261 3110 1271 3135
rect 1296 3110 1306 3135
rect 1261 3105 1306 3110
rect 1165 3070 1195 3100
rect 2295 3080 2330 3105
rect 46 3060 91 3065
rect 46 3035 56 3060
rect 81 3035 91 3060
rect 46 3030 91 3035
rect 1080 3005 1115 3030
rect 46 3000 91 3005
rect 46 2975 56 3000
rect 81 2975 91 3000
rect 46 2970 91 2975
rect 1266 3045 1306 3080
rect 910 2910 1120 2915
rect 910 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1120 2910
rect 910 2875 1120 2880
rect 1266 2900 1286 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 14970 3170 15040 3200
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 5320 3110 5350 3140
rect 3990 3050 4020 3080
rect 2330 2985 2370 3020
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 1306 2960 1341 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3080 2975 3120 2985
rect 3080 2955 3090 2975
rect 3110 2955 3120 2975
rect 3080 2945 3120 2955
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2975 3305 2985
rect 3265 2955 3275 2975
rect 3295 2955 3305 2975
rect 3265 2945 3305 2955
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2975 3665 2985
rect 3625 2955 3635 2975
rect 3655 2955 3665 2975
rect 3625 2945 3665 2955
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2975 4205 2985
rect 4165 2955 4175 2975
rect 4195 2955 4205 2975
rect 4165 2945 4205 2955
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2975 4565 2985
rect 4525 2955 4535 2975
rect 4555 2955 4565 2975
rect 4525 2945 4565 2955
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 3095 2925 3115 2945
rect 3275 2925 3295 2945
rect 3455 2925 3475 2945
rect 3635 2925 3655 2945
rect 3815 2925 3835 2945
rect 3995 2925 4015 2945
rect 4175 2925 4195 2945
rect 4355 2925 4375 2945
rect 4535 2925 4555 2945
rect 4715 2925 4735 2945
rect 4895 2925 4915 2945
rect 14970 3150 14975 3170
rect 14995 3150 15015 3170
rect 15035 3150 15040 3170
rect 14970 3120 15040 3150
rect 14970 3100 14975 3120
rect 14995 3100 15015 3120
rect 15035 3100 15040 3120
rect 14970 3070 15040 3100
rect 14970 3050 14975 3070
rect 14995 3050 15015 3070
rect 15035 3050 15040 3070
rect 14970 3020 15040 3050
rect 14970 3000 14975 3020
rect 14995 3000 15015 3020
rect 15035 3000 15040 3020
rect 14970 2990 15040 3000
rect 15065 3570 15095 3580
rect 15065 3550 15070 3570
rect 15090 3550 15095 3570
rect 15065 3520 15095 3550
rect 15065 3500 15070 3520
rect 15090 3500 15095 3520
rect 15065 3470 15095 3500
rect 15065 3450 15070 3470
rect 15090 3450 15095 3470
rect 15065 3420 15095 3450
rect 15065 3400 15070 3420
rect 15090 3400 15095 3420
rect 15065 3370 15095 3400
rect 15065 3350 15070 3370
rect 15090 3350 15095 3370
rect 15065 3320 15095 3350
rect 15065 3300 15070 3320
rect 15090 3300 15095 3320
rect 15065 3270 15095 3300
rect 15065 3250 15070 3270
rect 15090 3250 15095 3270
rect 15065 3220 15095 3250
rect 15065 3200 15070 3220
rect 15090 3200 15095 3220
rect 15065 3170 15095 3200
rect 15065 3150 15070 3170
rect 15090 3150 15095 3170
rect 15065 3120 15095 3150
rect 15065 3100 15070 3120
rect 15090 3100 15095 3120
rect 15065 3070 15095 3100
rect 15065 3050 15070 3070
rect 15090 3050 15095 3070
rect 15065 3020 15095 3050
rect 15065 3000 15070 3020
rect 15090 3000 15095 3020
rect 15065 2990 15095 3000
rect 15120 3570 15150 3580
rect 15120 3550 15125 3570
rect 15145 3550 15150 3570
rect 15120 3520 15150 3550
rect 15120 3500 15125 3520
rect 15145 3500 15150 3520
rect 15120 3470 15150 3500
rect 15120 3450 15125 3470
rect 15145 3450 15150 3470
rect 15120 3420 15150 3450
rect 15120 3400 15125 3420
rect 15145 3400 15150 3420
rect 15120 3370 15150 3400
rect 15120 3350 15125 3370
rect 15145 3350 15150 3370
rect 15120 3320 15150 3350
rect 15120 3300 15125 3320
rect 15145 3300 15150 3320
rect 15120 3270 15150 3300
rect 15120 3250 15125 3270
rect 15145 3250 15150 3270
rect 15120 3220 15150 3250
rect 15120 3200 15125 3220
rect 15145 3200 15150 3220
rect 15120 3170 15150 3200
rect 15120 3150 15125 3170
rect 15145 3150 15150 3170
rect 15120 3120 15150 3150
rect 15120 3100 15125 3120
rect 15145 3100 15150 3120
rect 15120 3070 15150 3100
rect 15120 3050 15125 3070
rect 15145 3050 15150 3070
rect 15120 3020 15150 3050
rect 15120 3000 15125 3020
rect 15145 3000 15150 3020
rect 15120 2990 15150 3000
rect 15175 3570 15205 3580
rect 15175 3550 15180 3570
rect 15200 3550 15205 3570
rect 15175 3520 15205 3550
rect 15175 3500 15180 3520
rect 15200 3500 15205 3520
rect 15175 3470 15205 3500
rect 15175 3450 15180 3470
rect 15200 3450 15205 3470
rect 15175 3420 15205 3450
rect 15175 3400 15180 3420
rect 15200 3400 15205 3420
rect 15175 3370 15205 3400
rect 15175 3350 15180 3370
rect 15200 3350 15205 3370
rect 15175 3320 15205 3350
rect 15175 3300 15180 3320
rect 15200 3300 15205 3320
rect 15175 3270 15205 3300
rect 15175 3250 15180 3270
rect 15200 3250 15205 3270
rect 15175 3220 15205 3250
rect 15175 3200 15180 3220
rect 15200 3200 15205 3220
rect 15175 3170 15205 3200
rect 15175 3150 15180 3170
rect 15200 3150 15205 3170
rect 15175 3120 15205 3150
rect 15175 3100 15180 3120
rect 15200 3100 15205 3120
rect 15175 3070 15205 3100
rect 15175 3050 15180 3070
rect 15200 3050 15205 3070
rect 15175 3020 15205 3050
rect 15175 3000 15180 3020
rect 15200 3000 15205 3020
rect 15175 2990 15205 3000
rect 15230 3570 15260 3580
rect 15230 3550 15235 3570
rect 15255 3550 15260 3570
rect 15230 3520 15260 3550
rect 15230 3500 15235 3520
rect 15255 3500 15260 3520
rect 15230 3470 15260 3500
rect 15230 3450 15235 3470
rect 15255 3450 15260 3470
rect 15230 3420 15260 3450
rect 15230 3400 15235 3420
rect 15255 3400 15260 3420
rect 15230 3370 15260 3400
rect 15230 3350 15235 3370
rect 15255 3350 15260 3370
rect 15230 3320 15260 3350
rect 15230 3300 15235 3320
rect 15255 3300 15260 3320
rect 15230 3270 15260 3300
rect 15230 3250 15235 3270
rect 15255 3250 15260 3270
rect 15230 3220 15260 3250
rect 15230 3200 15235 3220
rect 15255 3200 15260 3220
rect 15230 3170 15260 3200
rect 15230 3150 15235 3170
rect 15255 3150 15260 3170
rect 15230 3120 15260 3150
rect 15230 3100 15235 3120
rect 15255 3100 15260 3120
rect 15230 3070 15260 3100
rect 15230 3050 15235 3070
rect 15255 3050 15260 3070
rect 15230 3020 15260 3050
rect 15230 3000 15235 3020
rect 15255 3000 15260 3020
rect 15230 2990 15260 3000
rect 15285 3570 15315 3580
rect 15285 3550 15290 3570
rect 15310 3550 15315 3570
rect 15285 3520 15315 3550
rect 15285 3500 15290 3520
rect 15310 3500 15315 3520
rect 15285 3470 15315 3500
rect 15285 3450 15290 3470
rect 15310 3450 15315 3470
rect 15285 3420 15315 3450
rect 15285 3400 15290 3420
rect 15310 3400 15315 3420
rect 15285 3370 15315 3400
rect 15285 3350 15290 3370
rect 15310 3350 15315 3370
rect 15285 3320 15315 3350
rect 15285 3300 15290 3320
rect 15310 3300 15315 3320
rect 15285 3270 15315 3300
rect 15285 3250 15290 3270
rect 15310 3250 15315 3270
rect 15285 3220 15315 3250
rect 15285 3200 15290 3220
rect 15310 3200 15315 3220
rect 15285 3170 15315 3200
rect 15285 3150 15290 3170
rect 15310 3150 15315 3170
rect 15285 3120 15315 3150
rect 15285 3100 15290 3120
rect 15310 3100 15315 3120
rect 15285 3070 15315 3100
rect 15285 3050 15290 3070
rect 15310 3050 15315 3070
rect 15285 3020 15315 3050
rect 15285 3000 15290 3020
rect 15310 3000 15315 3020
rect 15285 2990 15315 3000
rect 15340 3570 15370 3580
rect 15340 3550 15345 3570
rect 15365 3550 15370 3570
rect 15340 3520 15370 3550
rect 15340 3500 15345 3520
rect 15365 3500 15370 3520
rect 15340 3470 15370 3500
rect 15340 3450 15345 3470
rect 15365 3450 15370 3470
rect 15340 3420 15370 3450
rect 15340 3400 15345 3420
rect 15365 3400 15370 3420
rect 15340 3370 15370 3400
rect 15340 3350 15345 3370
rect 15365 3350 15370 3370
rect 15340 3320 15370 3350
rect 15340 3300 15345 3320
rect 15365 3300 15370 3320
rect 15340 3270 15370 3300
rect 15340 3250 15345 3270
rect 15365 3250 15370 3270
rect 15340 3220 15370 3250
rect 15340 3200 15345 3220
rect 15365 3200 15370 3220
rect 15340 3170 15370 3200
rect 15340 3150 15345 3170
rect 15365 3150 15370 3170
rect 15340 3120 15370 3150
rect 15340 3100 15345 3120
rect 15365 3100 15370 3120
rect 15340 3070 15370 3100
rect 15340 3050 15345 3070
rect 15365 3050 15370 3070
rect 15340 3020 15370 3050
rect 15340 3000 15345 3020
rect 15365 3000 15370 3020
rect 15340 2990 15370 3000
rect 15395 3570 15425 3580
rect 15395 3550 15400 3570
rect 15420 3550 15425 3570
rect 15395 3520 15425 3550
rect 15395 3500 15400 3520
rect 15420 3500 15425 3520
rect 15395 3470 15425 3500
rect 15395 3450 15400 3470
rect 15420 3450 15425 3470
rect 15395 3420 15425 3450
rect 15395 3400 15400 3420
rect 15420 3400 15425 3420
rect 15395 3370 15425 3400
rect 15395 3350 15400 3370
rect 15420 3350 15425 3370
rect 15395 3320 15425 3350
rect 15395 3300 15400 3320
rect 15420 3300 15425 3320
rect 15395 3270 15425 3300
rect 15395 3250 15400 3270
rect 15420 3250 15425 3270
rect 15395 3220 15425 3250
rect 15395 3200 15400 3220
rect 15420 3200 15425 3220
rect 15395 3170 15425 3200
rect 15395 3150 15400 3170
rect 15420 3150 15425 3170
rect 15395 3120 15425 3150
rect 15395 3100 15400 3120
rect 15420 3100 15425 3120
rect 15395 3070 15425 3100
rect 15395 3050 15400 3070
rect 15420 3050 15425 3070
rect 15395 3020 15425 3050
rect 15395 3000 15400 3020
rect 15420 3000 15425 3020
rect 15395 2990 15425 3000
rect 15450 3570 15480 3580
rect 15450 3550 15455 3570
rect 15475 3550 15480 3570
rect 15450 3520 15480 3550
rect 15450 3500 15455 3520
rect 15475 3500 15480 3520
rect 15450 3470 15480 3500
rect 15450 3450 15455 3470
rect 15475 3450 15480 3470
rect 15450 3420 15480 3450
rect 15450 3400 15455 3420
rect 15475 3400 15480 3420
rect 15450 3370 15480 3400
rect 15450 3350 15455 3370
rect 15475 3350 15480 3370
rect 15450 3320 15480 3350
rect 15450 3300 15455 3320
rect 15475 3300 15480 3320
rect 15450 3270 15480 3300
rect 15450 3250 15455 3270
rect 15475 3250 15480 3270
rect 15450 3220 15480 3250
rect 15450 3200 15455 3220
rect 15475 3200 15480 3220
rect 15450 3170 15480 3200
rect 15450 3150 15455 3170
rect 15475 3150 15480 3170
rect 15450 3120 15480 3150
rect 15450 3100 15455 3120
rect 15475 3100 15480 3120
rect 15450 3070 15480 3100
rect 15450 3050 15455 3070
rect 15475 3050 15480 3070
rect 15450 3020 15480 3050
rect 15450 3000 15455 3020
rect 15475 3000 15480 3020
rect 15450 2990 15480 3000
rect 15505 3570 15535 3580
rect 15505 3550 15510 3570
rect 15530 3550 15535 3570
rect 15505 3520 15535 3550
rect 15505 3500 15510 3520
rect 15530 3500 15535 3520
rect 15505 3470 15535 3500
rect 15505 3450 15510 3470
rect 15530 3450 15535 3470
rect 15505 3420 15535 3450
rect 15505 3400 15510 3420
rect 15530 3400 15535 3420
rect 15505 3370 15535 3400
rect 15505 3350 15510 3370
rect 15530 3350 15535 3370
rect 15505 3320 15535 3350
rect 15505 3300 15510 3320
rect 15530 3300 15535 3320
rect 15505 3270 15535 3300
rect 15505 3250 15510 3270
rect 15530 3250 15535 3270
rect 15505 3220 15535 3250
rect 15505 3200 15510 3220
rect 15530 3200 15535 3220
rect 15505 3170 15535 3200
rect 15505 3150 15510 3170
rect 15530 3150 15535 3170
rect 15505 3120 15535 3150
rect 15505 3100 15510 3120
rect 15530 3100 15535 3120
rect 15505 3070 15535 3100
rect 15505 3050 15510 3070
rect 15530 3050 15535 3070
rect 15505 3020 15535 3050
rect 15505 3000 15510 3020
rect 15530 3000 15535 3020
rect 15505 2990 15535 3000
rect 15560 3570 15590 3580
rect 15560 3550 15565 3570
rect 15585 3550 15590 3570
rect 15560 3520 15590 3550
rect 15560 3500 15565 3520
rect 15585 3500 15590 3520
rect 15560 3470 15590 3500
rect 15560 3450 15565 3470
rect 15585 3450 15590 3470
rect 15560 3420 15590 3450
rect 15560 3400 15565 3420
rect 15585 3400 15590 3420
rect 15560 3370 15590 3400
rect 15560 3350 15565 3370
rect 15585 3350 15590 3370
rect 15560 3320 15590 3350
rect 15560 3300 15565 3320
rect 15585 3300 15590 3320
rect 15560 3270 15590 3300
rect 15560 3250 15565 3270
rect 15585 3250 15590 3270
rect 15560 3220 15590 3250
rect 15560 3200 15565 3220
rect 15585 3200 15590 3220
rect 15560 3170 15590 3200
rect 15560 3150 15565 3170
rect 15585 3150 15590 3170
rect 15560 3120 15590 3150
rect 15560 3100 15565 3120
rect 15585 3100 15590 3120
rect 15560 3070 15590 3100
rect 15560 3050 15565 3070
rect 15585 3050 15590 3070
rect 15560 3020 15590 3050
rect 15560 3000 15565 3020
rect 15585 3000 15590 3020
rect 15560 2990 15590 3000
rect 15615 3570 15645 3580
rect 15615 3550 15620 3570
rect 15640 3550 15645 3570
rect 15615 3520 15645 3550
rect 15615 3500 15620 3520
rect 15640 3500 15645 3520
rect 15615 3470 15645 3500
rect 15615 3450 15620 3470
rect 15640 3450 15645 3470
rect 15615 3420 15645 3450
rect 15615 3400 15620 3420
rect 15640 3400 15645 3420
rect 15615 3370 15645 3400
rect 15615 3350 15620 3370
rect 15640 3350 15645 3370
rect 15615 3320 15645 3350
rect 15615 3300 15620 3320
rect 15640 3300 15645 3320
rect 15615 3270 15645 3300
rect 15615 3250 15620 3270
rect 15640 3250 15645 3270
rect 15615 3220 15645 3250
rect 15615 3200 15620 3220
rect 15640 3200 15645 3220
rect 15615 3170 15645 3200
rect 15615 3150 15620 3170
rect 15640 3150 15645 3170
rect 15615 3120 15645 3150
rect 15615 3100 15620 3120
rect 15640 3100 15645 3120
rect 15615 3070 15645 3100
rect 15615 3050 15620 3070
rect 15640 3050 15645 3070
rect 15615 3020 15645 3050
rect 15615 3000 15620 3020
rect 15640 3000 15645 3020
rect 15615 2990 15645 3000
rect 15670 3570 15740 3580
rect 15670 3550 15675 3570
rect 15695 3550 15715 3570
rect 15735 3550 15740 3570
rect 15670 3520 15740 3550
rect 16180 3570 16220 3580
rect 16180 3550 16190 3570
rect 16210 3550 16220 3570
rect 16180 3540 16220 3550
rect 16340 3570 16380 3580
rect 16340 3550 16350 3570
rect 16370 3550 16380 3570
rect 16340 3540 16380 3550
rect 16460 3570 16500 3580
rect 16460 3550 16470 3570
rect 16490 3550 16500 3570
rect 16460 3540 16500 3550
rect 16580 3570 16620 3580
rect 16580 3550 16590 3570
rect 16610 3550 16620 3570
rect 16580 3540 16620 3550
rect 16700 3570 16740 3580
rect 16700 3550 16710 3570
rect 16730 3550 16740 3570
rect 16700 3540 16740 3550
rect 16820 3570 16860 3580
rect 16820 3550 16830 3570
rect 16850 3550 16860 3570
rect 16820 3540 16860 3550
rect 16940 3570 16980 3580
rect 16940 3550 16950 3570
rect 16970 3550 16980 3570
rect 16940 3540 16980 3550
rect 17060 3570 17100 3580
rect 17060 3550 17070 3570
rect 17090 3550 17100 3570
rect 17060 3540 17100 3550
rect 17180 3570 17220 3580
rect 17180 3550 17190 3570
rect 17210 3550 17220 3570
rect 17180 3540 17220 3550
rect 17300 3570 17340 3580
rect 17300 3550 17310 3570
rect 17330 3550 17340 3570
rect 17300 3540 17340 3550
rect 17420 3570 17460 3580
rect 17420 3550 17430 3570
rect 17450 3550 17460 3570
rect 17420 3540 17460 3550
rect 17580 3570 17620 3580
rect 17580 3550 17590 3570
rect 17610 3550 17620 3570
rect 17580 3540 17620 3550
rect 18110 3570 18180 3580
rect 18110 3550 18115 3570
rect 18135 3550 18155 3570
rect 18175 3550 18180 3570
rect 16190 3520 16210 3540
rect 16350 3520 16370 3540
rect 16470 3520 16490 3540
rect 16590 3520 16610 3540
rect 16710 3520 16730 3540
rect 16830 3520 16850 3540
rect 16950 3520 16970 3540
rect 17070 3520 17090 3540
rect 17190 3520 17210 3540
rect 17310 3520 17330 3540
rect 17430 3520 17450 3540
rect 17590 3520 17610 3540
rect 18110 3520 18180 3550
rect 15670 3500 15675 3520
rect 15695 3500 15715 3520
rect 15735 3500 15740 3520
rect 15670 3470 15740 3500
rect 15670 3450 15675 3470
rect 15695 3450 15715 3470
rect 15735 3450 15740 3470
rect 15670 3420 15740 3450
rect 15670 3400 15675 3420
rect 15695 3400 15715 3420
rect 15735 3400 15740 3420
rect 15670 3370 15740 3400
rect 15670 3350 15675 3370
rect 15695 3350 15715 3370
rect 15735 3350 15740 3370
rect 15670 3320 15740 3350
rect 15670 3300 15675 3320
rect 15695 3300 15715 3320
rect 15735 3300 15740 3320
rect 15670 3270 15740 3300
rect 15670 3250 15675 3270
rect 15695 3250 15715 3270
rect 15735 3250 15740 3270
rect 15670 3220 15740 3250
rect 15670 3200 15675 3220
rect 15695 3200 15715 3220
rect 15735 3200 15740 3220
rect 15670 3170 15740 3200
rect 15670 3150 15675 3170
rect 15695 3150 15715 3170
rect 15735 3150 15740 3170
rect 15670 3120 15740 3150
rect 16185 3510 16255 3520
rect 16185 3490 16190 3510
rect 16210 3490 16230 3510
rect 16250 3490 16255 3510
rect 16185 3460 16255 3490
rect 16185 3440 16190 3460
rect 16210 3440 16230 3460
rect 16250 3440 16255 3460
rect 16185 3410 16255 3440
rect 16185 3390 16190 3410
rect 16210 3390 16230 3410
rect 16250 3390 16255 3410
rect 16185 3360 16255 3390
rect 16185 3340 16190 3360
rect 16210 3340 16230 3360
rect 16250 3340 16255 3360
rect 16185 3310 16255 3340
rect 16185 3290 16190 3310
rect 16210 3290 16230 3310
rect 16250 3290 16255 3310
rect 16185 3260 16255 3290
rect 16185 3240 16190 3260
rect 16210 3240 16230 3260
rect 16250 3240 16255 3260
rect 16185 3210 16255 3240
rect 16185 3190 16190 3210
rect 16210 3190 16230 3210
rect 16250 3190 16255 3210
rect 16185 3160 16255 3190
rect 16185 3140 16190 3160
rect 16210 3140 16230 3160
rect 16250 3140 16255 3160
rect 16185 3130 16255 3140
rect 16285 3510 16315 3520
rect 16285 3490 16290 3510
rect 16310 3490 16315 3510
rect 16285 3460 16315 3490
rect 16285 3440 16290 3460
rect 16310 3440 16315 3460
rect 16285 3410 16315 3440
rect 16285 3390 16290 3410
rect 16310 3390 16315 3410
rect 16285 3360 16315 3390
rect 16285 3340 16290 3360
rect 16310 3340 16315 3360
rect 16285 3310 16315 3340
rect 16285 3290 16290 3310
rect 16310 3290 16315 3310
rect 16285 3260 16315 3290
rect 16285 3240 16290 3260
rect 16310 3240 16315 3260
rect 16285 3210 16315 3240
rect 16285 3190 16290 3210
rect 16310 3190 16315 3210
rect 16285 3160 16315 3190
rect 16285 3140 16290 3160
rect 16310 3140 16315 3160
rect 16285 3130 16315 3140
rect 16345 3510 16375 3520
rect 16345 3490 16350 3510
rect 16370 3490 16375 3510
rect 16345 3460 16375 3490
rect 16345 3440 16350 3460
rect 16370 3440 16375 3460
rect 16345 3410 16375 3440
rect 16345 3390 16350 3410
rect 16370 3390 16375 3410
rect 16345 3360 16375 3390
rect 16345 3340 16350 3360
rect 16370 3340 16375 3360
rect 16345 3310 16375 3340
rect 16345 3290 16350 3310
rect 16370 3290 16375 3310
rect 16345 3260 16375 3290
rect 16345 3240 16350 3260
rect 16370 3240 16375 3260
rect 16345 3210 16375 3240
rect 16345 3190 16350 3210
rect 16370 3190 16375 3210
rect 16345 3160 16375 3190
rect 16345 3140 16350 3160
rect 16370 3140 16375 3160
rect 16345 3130 16375 3140
rect 16405 3510 16435 3520
rect 16405 3490 16410 3510
rect 16430 3490 16435 3510
rect 16405 3460 16435 3490
rect 16405 3440 16410 3460
rect 16430 3440 16435 3460
rect 16405 3410 16435 3440
rect 16405 3390 16410 3410
rect 16430 3390 16435 3410
rect 16405 3360 16435 3390
rect 16405 3340 16410 3360
rect 16430 3340 16435 3360
rect 16405 3310 16435 3340
rect 16405 3290 16410 3310
rect 16430 3290 16435 3310
rect 16405 3260 16435 3290
rect 16405 3240 16410 3260
rect 16430 3240 16435 3260
rect 16405 3210 16435 3240
rect 16405 3190 16410 3210
rect 16430 3190 16435 3210
rect 16405 3160 16435 3190
rect 16405 3140 16410 3160
rect 16430 3140 16435 3160
rect 16405 3130 16435 3140
rect 16465 3510 16495 3520
rect 16465 3490 16470 3510
rect 16490 3490 16495 3510
rect 16465 3460 16495 3490
rect 16465 3440 16470 3460
rect 16490 3440 16495 3460
rect 16465 3410 16495 3440
rect 16465 3390 16470 3410
rect 16490 3390 16495 3410
rect 16465 3360 16495 3390
rect 16465 3340 16470 3360
rect 16490 3340 16495 3360
rect 16465 3310 16495 3340
rect 16465 3290 16470 3310
rect 16490 3290 16495 3310
rect 16465 3260 16495 3290
rect 16465 3240 16470 3260
rect 16490 3240 16495 3260
rect 16465 3210 16495 3240
rect 16465 3190 16470 3210
rect 16490 3190 16495 3210
rect 16465 3160 16495 3190
rect 16465 3140 16470 3160
rect 16490 3140 16495 3160
rect 16465 3130 16495 3140
rect 16525 3510 16555 3520
rect 16525 3490 16530 3510
rect 16550 3490 16555 3510
rect 16525 3460 16555 3490
rect 16525 3440 16530 3460
rect 16550 3440 16555 3460
rect 16525 3410 16555 3440
rect 16525 3390 16530 3410
rect 16550 3390 16555 3410
rect 16525 3360 16555 3390
rect 16525 3340 16530 3360
rect 16550 3340 16555 3360
rect 16525 3310 16555 3340
rect 16525 3290 16530 3310
rect 16550 3290 16555 3310
rect 16525 3260 16555 3290
rect 16525 3240 16530 3260
rect 16550 3240 16555 3260
rect 16525 3210 16555 3240
rect 16525 3190 16530 3210
rect 16550 3190 16555 3210
rect 16525 3160 16555 3190
rect 16525 3140 16530 3160
rect 16550 3140 16555 3160
rect 16525 3130 16555 3140
rect 16585 3510 16615 3520
rect 16585 3490 16590 3510
rect 16610 3490 16615 3510
rect 16585 3460 16615 3490
rect 16585 3440 16590 3460
rect 16610 3440 16615 3460
rect 16585 3410 16615 3440
rect 16585 3390 16590 3410
rect 16610 3390 16615 3410
rect 16585 3360 16615 3390
rect 16585 3340 16590 3360
rect 16610 3340 16615 3360
rect 16585 3310 16615 3340
rect 16585 3290 16590 3310
rect 16610 3290 16615 3310
rect 16585 3260 16615 3290
rect 16585 3240 16590 3260
rect 16610 3240 16615 3260
rect 16585 3210 16615 3240
rect 16585 3190 16590 3210
rect 16610 3190 16615 3210
rect 16585 3160 16615 3190
rect 16585 3140 16590 3160
rect 16610 3140 16615 3160
rect 16585 3130 16615 3140
rect 16645 3510 16675 3520
rect 16645 3490 16650 3510
rect 16670 3490 16675 3510
rect 16645 3460 16675 3490
rect 16645 3440 16650 3460
rect 16670 3440 16675 3460
rect 16645 3410 16675 3440
rect 16645 3390 16650 3410
rect 16670 3390 16675 3410
rect 16645 3360 16675 3390
rect 16645 3340 16650 3360
rect 16670 3340 16675 3360
rect 16645 3310 16675 3340
rect 16645 3290 16650 3310
rect 16670 3290 16675 3310
rect 16645 3260 16675 3290
rect 16645 3240 16650 3260
rect 16670 3240 16675 3260
rect 16645 3210 16675 3240
rect 16645 3190 16650 3210
rect 16670 3190 16675 3210
rect 16645 3160 16675 3190
rect 16645 3140 16650 3160
rect 16670 3140 16675 3160
rect 16645 3130 16675 3140
rect 16705 3510 16735 3520
rect 16705 3490 16710 3510
rect 16730 3490 16735 3510
rect 16705 3460 16735 3490
rect 16705 3440 16710 3460
rect 16730 3440 16735 3460
rect 16705 3410 16735 3440
rect 16705 3390 16710 3410
rect 16730 3390 16735 3410
rect 16705 3360 16735 3390
rect 16705 3340 16710 3360
rect 16730 3340 16735 3360
rect 16705 3310 16735 3340
rect 16705 3290 16710 3310
rect 16730 3290 16735 3310
rect 16705 3260 16735 3290
rect 16705 3240 16710 3260
rect 16730 3240 16735 3260
rect 16705 3210 16735 3240
rect 16705 3190 16710 3210
rect 16730 3190 16735 3210
rect 16705 3160 16735 3190
rect 16705 3140 16710 3160
rect 16730 3140 16735 3160
rect 16705 3130 16735 3140
rect 16765 3510 16795 3520
rect 16765 3490 16770 3510
rect 16790 3490 16795 3510
rect 16765 3460 16795 3490
rect 16765 3440 16770 3460
rect 16790 3440 16795 3460
rect 16765 3410 16795 3440
rect 16765 3390 16770 3410
rect 16790 3390 16795 3410
rect 16765 3360 16795 3390
rect 16765 3340 16770 3360
rect 16790 3340 16795 3360
rect 16765 3310 16795 3340
rect 16765 3290 16770 3310
rect 16790 3290 16795 3310
rect 16765 3260 16795 3290
rect 16765 3240 16770 3260
rect 16790 3240 16795 3260
rect 16765 3210 16795 3240
rect 16765 3190 16770 3210
rect 16790 3190 16795 3210
rect 16765 3160 16795 3190
rect 16765 3140 16770 3160
rect 16790 3140 16795 3160
rect 16765 3130 16795 3140
rect 16825 3510 16855 3520
rect 16825 3490 16830 3510
rect 16850 3490 16855 3510
rect 16825 3460 16855 3490
rect 16825 3440 16830 3460
rect 16850 3440 16855 3460
rect 16825 3410 16855 3440
rect 16825 3390 16830 3410
rect 16850 3390 16855 3410
rect 16825 3360 16855 3390
rect 16825 3340 16830 3360
rect 16850 3340 16855 3360
rect 16825 3310 16855 3340
rect 16825 3290 16830 3310
rect 16850 3290 16855 3310
rect 16825 3260 16855 3290
rect 16825 3240 16830 3260
rect 16850 3240 16855 3260
rect 16825 3210 16855 3240
rect 16825 3190 16830 3210
rect 16850 3190 16855 3210
rect 16825 3160 16855 3190
rect 16825 3140 16830 3160
rect 16850 3140 16855 3160
rect 16825 3130 16855 3140
rect 16885 3510 16915 3520
rect 16885 3490 16890 3510
rect 16910 3490 16915 3510
rect 16885 3460 16915 3490
rect 16885 3440 16890 3460
rect 16910 3440 16915 3460
rect 16885 3410 16915 3440
rect 16885 3390 16890 3410
rect 16910 3390 16915 3410
rect 16885 3360 16915 3390
rect 16885 3340 16890 3360
rect 16910 3340 16915 3360
rect 16885 3310 16915 3340
rect 16885 3290 16890 3310
rect 16910 3290 16915 3310
rect 16885 3260 16915 3290
rect 16885 3240 16890 3260
rect 16910 3240 16915 3260
rect 16885 3210 16915 3240
rect 16885 3190 16890 3210
rect 16910 3190 16915 3210
rect 16885 3160 16915 3190
rect 16885 3140 16890 3160
rect 16910 3140 16915 3160
rect 16885 3130 16915 3140
rect 16945 3510 16975 3520
rect 16945 3490 16950 3510
rect 16970 3490 16975 3510
rect 16945 3460 16975 3490
rect 16945 3440 16950 3460
rect 16970 3440 16975 3460
rect 16945 3410 16975 3440
rect 16945 3390 16950 3410
rect 16970 3390 16975 3410
rect 16945 3360 16975 3390
rect 16945 3340 16950 3360
rect 16970 3340 16975 3360
rect 16945 3310 16975 3340
rect 16945 3290 16950 3310
rect 16970 3290 16975 3310
rect 16945 3260 16975 3290
rect 16945 3240 16950 3260
rect 16970 3240 16975 3260
rect 16945 3210 16975 3240
rect 16945 3190 16950 3210
rect 16970 3190 16975 3210
rect 16945 3160 16975 3190
rect 16945 3140 16950 3160
rect 16970 3140 16975 3160
rect 16945 3130 16975 3140
rect 17005 3510 17035 3520
rect 17005 3490 17010 3510
rect 17030 3490 17035 3510
rect 17005 3460 17035 3490
rect 17005 3440 17010 3460
rect 17030 3440 17035 3460
rect 17005 3410 17035 3440
rect 17005 3390 17010 3410
rect 17030 3390 17035 3410
rect 17005 3360 17035 3390
rect 17005 3340 17010 3360
rect 17030 3340 17035 3360
rect 17005 3310 17035 3340
rect 17005 3290 17010 3310
rect 17030 3290 17035 3310
rect 17005 3260 17035 3290
rect 17005 3240 17010 3260
rect 17030 3240 17035 3260
rect 17005 3210 17035 3240
rect 17005 3190 17010 3210
rect 17030 3190 17035 3210
rect 17005 3160 17035 3190
rect 17005 3140 17010 3160
rect 17030 3140 17035 3160
rect 17005 3130 17035 3140
rect 17065 3510 17095 3520
rect 17065 3490 17070 3510
rect 17090 3490 17095 3510
rect 17065 3460 17095 3490
rect 17065 3440 17070 3460
rect 17090 3440 17095 3460
rect 17065 3410 17095 3440
rect 17065 3390 17070 3410
rect 17090 3390 17095 3410
rect 17065 3360 17095 3390
rect 17065 3340 17070 3360
rect 17090 3340 17095 3360
rect 17065 3310 17095 3340
rect 17065 3290 17070 3310
rect 17090 3290 17095 3310
rect 17065 3260 17095 3290
rect 17065 3240 17070 3260
rect 17090 3240 17095 3260
rect 17065 3210 17095 3240
rect 17065 3190 17070 3210
rect 17090 3190 17095 3210
rect 17065 3160 17095 3190
rect 17065 3140 17070 3160
rect 17090 3140 17095 3160
rect 17065 3130 17095 3140
rect 17125 3510 17155 3520
rect 17125 3490 17130 3510
rect 17150 3490 17155 3510
rect 17125 3460 17155 3490
rect 17125 3440 17130 3460
rect 17150 3440 17155 3460
rect 17125 3410 17155 3440
rect 17125 3390 17130 3410
rect 17150 3390 17155 3410
rect 17125 3360 17155 3390
rect 17125 3340 17130 3360
rect 17150 3340 17155 3360
rect 17125 3310 17155 3340
rect 17125 3290 17130 3310
rect 17150 3290 17155 3310
rect 17125 3260 17155 3290
rect 17125 3240 17130 3260
rect 17150 3240 17155 3260
rect 17125 3210 17155 3240
rect 17125 3190 17130 3210
rect 17150 3190 17155 3210
rect 17125 3160 17155 3190
rect 17125 3140 17130 3160
rect 17150 3140 17155 3160
rect 17125 3130 17155 3140
rect 17185 3510 17215 3520
rect 17185 3490 17190 3510
rect 17210 3490 17215 3510
rect 17185 3460 17215 3490
rect 17185 3440 17190 3460
rect 17210 3440 17215 3460
rect 17185 3410 17215 3440
rect 17185 3390 17190 3410
rect 17210 3390 17215 3410
rect 17185 3360 17215 3390
rect 17185 3340 17190 3360
rect 17210 3340 17215 3360
rect 17185 3310 17215 3340
rect 17185 3290 17190 3310
rect 17210 3290 17215 3310
rect 17185 3260 17215 3290
rect 17185 3240 17190 3260
rect 17210 3240 17215 3260
rect 17185 3210 17215 3240
rect 17185 3190 17190 3210
rect 17210 3190 17215 3210
rect 17185 3160 17215 3190
rect 17185 3140 17190 3160
rect 17210 3140 17215 3160
rect 17185 3130 17215 3140
rect 17245 3510 17275 3520
rect 17245 3490 17250 3510
rect 17270 3490 17275 3510
rect 17245 3460 17275 3490
rect 17245 3440 17250 3460
rect 17270 3440 17275 3460
rect 17245 3410 17275 3440
rect 17245 3390 17250 3410
rect 17270 3390 17275 3410
rect 17245 3360 17275 3390
rect 17245 3340 17250 3360
rect 17270 3340 17275 3360
rect 17245 3310 17275 3340
rect 17245 3290 17250 3310
rect 17270 3290 17275 3310
rect 17245 3260 17275 3290
rect 17245 3240 17250 3260
rect 17270 3240 17275 3260
rect 17245 3210 17275 3240
rect 17245 3190 17250 3210
rect 17270 3190 17275 3210
rect 17245 3160 17275 3190
rect 17245 3140 17250 3160
rect 17270 3140 17275 3160
rect 17245 3130 17275 3140
rect 17305 3510 17335 3520
rect 17305 3490 17310 3510
rect 17330 3490 17335 3510
rect 17305 3460 17335 3490
rect 17305 3440 17310 3460
rect 17330 3440 17335 3460
rect 17305 3410 17335 3440
rect 17305 3390 17310 3410
rect 17330 3390 17335 3410
rect 17305 3360 17335 3390
rect 17305 3340 17310 3360
rect 17330 3340 17335 3360
rect 17305 3310 17335 3340
rect 17305 3290 17310 3310
rect 17330 3290 17335 3310
rect 17305 3260 17335 3290
rect 17305 3240 17310 3260
rect 17330 3240 17335 3260
rect 17305 3210 17335 3240
rect 17305 3190 17310 3210
rect 17330 3190 17335 3210
rect 17305 3160 17335 3190
rect 17305 3140 17310 3160
rect 17330 3140 17335 3160
rect 17305 3130 17335 3140
rect 17365 3510 17395 3520
rect 17365 3490 17370 3510
rect 17390 3490 17395 3510
rect 17365 3460 17395 3490
rect 17365 3440 17370 3460
rect 17390 3440 17395 3460
rect 17365 3410 17395 3440
rect 17365 3390 17370 3410
rect 17390 3390 17395 3410
rect 17365 3360 17395 3390
rect 17365 3340 17370 3360
rect 17390 3340 17395 3360
rect 17365 3310 17395 3340
rect 17365 3290 17370 3310
rect 17390 3290 17395 3310
rect 17365 3260 17395 3290
rect 17365 3240 17370 3260
rect 17390 3240 17395 3260
rect 17365 3210 17395 3240
rect 17365 3190 17370 3210
rect 17390 3190 17395 3210
rect 17365 3160 17395 3190
rect 17365 3140 17370 3160
rect 17390 3140 17395 3160
rect 17365 3130 17395 3140
rect 17425 3510 17455 3520
rect 17425 3490 17430 3510
rect 17450 3490 17455 3510
rect 17425 3460 17455 3490
rect 17425 3440 17430 3460
rect 17450 3440 17455 3460
rect 17425 3410 17455 3440
rect 17425 3390 17430 3410
rect 17450 3390 17455 3410
rect 17425 3360 17455 3390
rect 17425 3340 17430 3360
rect 17450 3340 17455 3360
rect 17425 3310 17455 3340
rect 17425 3290 17430 3310
rect 17450 3290 17455 3310
rect 17425 3260 17455 3290
rect 17425 3240 17430 3260
rect 17450 3240 17455 3260
rect 17425 3210 17455 3240
rect 17425 3190 17430 3210
rect 17450 3190 17455 3210
rect 17425 3160 17455 3190
rect 17425 3140 17430 3160
rect 17450 3140 17455 3160
rect 17425 3130 17455 3140
rect 17485 3510 17515 3520
rect 17485 3490 17490 3510
rect 17510 3490 17515 3510
rect 17485 3460 17515 3490
rect 17485 3440 17490 3460
rect 17510 3440 17515 3460
rect 17485 3410 17515 3440
rect 17485 3390 17490 3410
rect 17510 3390 17515 3410
rect 17485 3360 17515 3390
rect 17485 3340 17490 3360
rect 17510 3340 17515 3360
rect 17485 3310 17515 3340
rect 17485 3290 17490 3310
rect 17510 3290 17515 3310
rect 17485 3260 17515 3290
rect 17485 3240 17490 3260
rect 17510 3240 17515 3260
rect 17485 3210 17515 3240
rect 17485 3190 17490 3210
rect 17510 3190 17515 3210
rect 17485 3160 17515 3190
rect 17485 3140 17490 3160
rect 17510 3140 17515 3160
rect 17485 3130 17515 3140
rect 17545 3510 17615 3520
rect 17545 3490 17550 3510
rect 17570 3490 17590 3510
rect 17610 3490 17615 3510
rect 17545 3460 17615 3490
rect 17545 3440 17550 3460
rect 17570 3440 17590 3460
rect 17610 3440 17615 3460
rect 17545 3410 17615 3440
rect 17545 3390 17550 3410
rect 17570 3390 17590 3410
rect 17610 3390 17615 3410
rect 17545 3360 17615 3390
rect 17545 3340 17550 3360
rect 17570 3340 17590 3360
rect 17610 3340 17615 3360
rect 17545 3310 17615 3340
rect 17545 3290 17550 3310
rect 17570 3290 17590 3310
rect 17610 3290 17615 3310
rect 17545 3260 17615 3290
rect 17545 3240 17550 3260
rect 17570 3240 17590 3260
rect 17610 3240 17615 3260
rect 17545 3210 17615 3240
rect 17545 3190 17550 3210
rect 17570 3190 17590 3210
rect 17610 3190 17615 3210
rect 17545 3160 17615 3190
rect 17545 3140 17550 3160
rect 17570 3140 17590 3160
rect 17610 3140 17615 3160
rect 17545 3130 17615 3140
rect 18110 3500 18115 3520
rect 18135 3500 18155 3520
rect 18175 3500 18180 3520
rect 18110 3470 18180 3500
rect 18110 3450 18115 3470
rect 18135 3450 18155 3470
rect 18175 3450 18180 3470
rect 18110 3420 18180 3450
rect 18110 3400 18115 3420
rect 18135 3400 18155 3420
rect 18175 3400 18180 3420
rect 18110 3370 18180 3400
rect 18110 3350 18115 3370
rect 18135 3350 18155 3370
rect 18175 3350 18180 3370
rect 18110 3320 18180 3350
rect 18110 3300 18115 3320
rect 18135 3300 18155 3320
rect 18175 3300 18180 3320
rect 18110 3270 18180 3300
rect 18110 3250 18115 3270
rect 18135 3250 18155 3270
rect 18175 3250 18180 3270
rect 18110 3220 18180 3250
rect 18110 3200 18115 3220
rect 18135 3200 18155 3220
rect 18175 3200 18180 3220
rect 18110 3170 18180 3200
rect 18110 3150 18115 3170
rect 18135 3150 18155 3170
rect 18175 3150 18180 3170
rect 15670 3100 15675 3120
rect 15695 3100 15715 3120
rect 15735 3100 15740 3120
rect 16290 3110 16310 3130
rect 16410 3110 16430 3130
rect 16530 3110 16550 3130
rect 16650 3110 16670 3130
rect 16770 3110 16790 3130
rect 16890 3110 16910 3130
rect 17010 3110 17030 3130
rect 17130 3110 17150 3130
rect 17250 3110 17270 3130
rect 17370 3110 17390 3130
rect 17490 3110 17510 3130
rect 18110 3120 18180 3150
rect 15670 3070 15740 3100
rect 16280 3100 16320 3110
rect 16280 3080 16290 3100
rect 16310 3080 16320 3100
rect 16280 3070 16320 3080
rect 16400 3100 16440 3110
rect 16400 3080 16410 3100
rect 16430 3080 16440 3100
rect 16400 3070 16440 3080
rect 16520 3100 16560 3110
rect 16520 3080 16530 3100
rect 16550 3080 16560 3100
rect 16520 3070 16560 3080
rect 16640 3100 16680 3110
rect 16640 3080 16650 3100
rect 16670 3080 16680 3100
rect 16640 3070 16680 3080
rect 16760 3100 16800 3110
rect 16760 3080 16770 3100
rect 16790 3080 16800 3100
rect 16760 3070 16800 3080
rect 16823 3100 16857 3110
rect 16823 3080 16831 3100
rect 16849 3080 16857 3100
rect 16823 3070 16857 3080
rect 16880 3100 16920 3110
rect 16880 3080 16890 3100
rect 16910 3080 16920 3100
rect 16880 3070 16920 3080
rect 17000 3100 17040 3110
rect 17000 3080 17010 3100
rect 17030 3080 17040 3100
rect 17000 3070 17040 3080
rect 17120 3100 17160 3110
rect 17120 3080 17130 3100
rect 17150 3080 17160 3100
rect 17120 3070 17160 3080
rect 17240 3100 17280 3110
rect 17240 3080 17250 3100
rect 17270 3080 17280 3100
rect 17240 3070 17280 3080
rect 17360 3100 17400 3110
rect 17360 3080 17370 3100
rect 17390 3080 17400 3100
rect 17360 3070 17400 3080
rect 17480 3100 17520 3110
rect 17480 3080 17490 3100
rect 17510 3080 17520 3100
rect 17480 3070 17520 3080
rect 18110 3100 18115 3120
rect 18135 3100 18155 3120
rect 18175 3100 18180 3120
rect 18110 3070 18180 3100
rect 15670 3050 15675 3070
rect 15695 3050 15715 3070
rect 15735 3050 15740 3070
rect 15670 3020 15740 3050
rect 15670 3000 15675 3020
rect 15695 3000 15715 3020
rect 15735 3000 15740 3020
rect 15670 2990 15740 3000
rect 18110 3050 18115 3070
rect 18135 3050 18155 3070
rect 18175 3050 18180 3070
rect 18110 3020 18180 3050
rect 18110 3000 18115 3020
rect 18135 3000 18155 3020
rect 18175 3000 18180 3020
rect 18110 2990 18180 3000
rect 18205 3570 18235 3580
rect 18205 3550 18210 3570
rect 18230 3550 18235 3570
rect 18205 3520 18235 3550
rect 18205 3500 18210 3520
rect 18230 3500 18235 3520
rect 18205 3470 18235 3500
rect 18205 3450 18210 3470
rect 18230 3450 18235 3470
rect 18205 3420 18235 3450
rect 18205 3400 18210 3420
rect 18230 3400 18235 3420
rect 18205 3370 18235 3400
rect 18205 3350 18210 3370
rect 18230 3350 18235 3370
rect 18205 3320 18235 3350
rect 18205 3300 18210 3320
rect 18230 3300 18235 3320
rect 18205 3270 18235 3300
rect 18205 3250 18210 3270
rect 18230 3250 18235 3270
rect 18205 3220 18235 3250
rect 18205 3200 18210 3220
rect 18230 3200 18235 3220
rect 18205 3170 18235 3200
rect 18205 3150 18210 3170
rect 18230 3150 18235 3170
rect 18205 3120 18235 3150
rect 18205 3100 18210 3120
rect 18230 3100 18235 3120
rect 18205 3070 18235 3100
rect 18205 3050 18210 3070
rect 18230 3050 18235 3070
rect 18205 3020 18235 3050
rect 18205 3000 18210 3020
rect 18230 3000 18235 3020
rect 18205 2990 18235 3000
rect 18260 3570 18290 3580
rect 18260 3550 18265 3570
rect 18285 3550 18290 3570
rect 18260 3520 18290 3550
rect 18260 3500 18265 3520
rect 18285 3500 18290 3520
rect 18260 3470 18290 3500
rect 18260 3450 18265 3470
rect 18285 3450 18290 3470
rect 18260 3420 18290 3450
rect 18260 3400 18265 3420
rect 18285 3400 18290 3420
rect 18260 3370 18290 3400
rect 18260 3350 18265 3370
rect 18285 3350 18290 3370
rect 18260 3320 18290 3350
rect 18260 3300 18265 3320
rect 18285 3300 18290 3320
rect 18260 3270 18290 3300
rect 18260 3250 18265 3270
rect 18285 3250 18290 3270
rect 18260 3220 18290 3250
rect 18260 3200 18265 3220
rect 18285 3200 18290 3220
rect 18260 3170 18290 3200
rect 18260 3150 18265 3170
rect 18285 3150 18290 3170
rect 18260 3120 18290 3150
rect 18260 3100 18265 3120
rect 18285 3100 18290 3120
rect 18260 3070 18290 3100
rect 18260 3050 18265 3070
rect 18285 3050 18290 3070
rect 18260 3020 18290 3050
rect 18260 3000 18265 3020
rect 18285 3000 18290 3020
rect 18260 2990 18290 3000
rect 18315 3570 18345 3580
rect 18315 3550 18320 3570
rect 18340 3550 18345 3570
rect 18315 3520 18345 3550
rect 18315 3500 18320 3520
rect 18340 3500 18345 3520
rect 18315 3470 18345 3500
rect 18315 3450 18320 3470
rect 18340 3450 18345 3470
rect 18315 3420 18345 3450
rect 18315 3400 18320 3420
rect 18340 3400 18345 3420
rect 18315 3370 18345 3400
rect 18315 3350 18320 3370
rect 18340 3350 18345 3370
rect 18315 3320 18345 3350
rect 18315 3300 18320 3320
rect 18340 3300 18345 3320
rect 18315 3270 18345 3300
rect 18315 3250 18320 3270
rect 18340 3250 18345 3270
rect 18315 3220 18345 3250
rect 18315 3200 18320 3220
rect 18340 3200 18345 3220
rect 18315 3170 18345 3200
rect 18315 3150 18320 3170
rect 18340 3150 18345 3170
rect 18315 3120 18345 3150
rect 18315 3100 18320 3120
rect 18340 3100 18345 3120
rect 18315 3070 18345 3100
rect 18315 3050 18320 3070
rect 18340 3050 18345 3070
rect 18315 3020 18345 3050
rect 18315 3000 18320 3020
rect 18340 3000 18345 3020
rect 18315 2990 18345 3000
rect 18370 3570 18400 3580
rect 18370 3550 18375 3570
rect 18395 3550 18400 3570
rect 18370 3520 18400 3550
rect 18370 3500 18375 3520
rect 18395 3500 18400 3520
rect 18370 3470 18400 3500
rect 18370 3450 18375 3470
rect 18395 3450 18400 3470
rect 18370 3420 18400 3450
rect 18370 3400 18375 3420
rect 18395 3400 18400 3420
rect 18370 3370 18400 3400
rect 18370 3350 18375 3370
rect 18395 3350 18400 3370
rect 18370 3320 18400 3350
rect 18370 3300 18375 3320
rect 18395 3300 18400 3320
rect 18370 3270 18400 3300
rect 18370 3250 18375 3270
rect 18395 3250 18400 3270
rect 18370 3220 18400 3250
rect 18370 3200 18375 3220
rect 18395 3200 18400 3220
rect 18370 3170 18400 3200
rect 18370 3150 18375 3170
rect 18395 3150 18400 3170
rect 18370 3120 18400 3150
rect 18370 3100 18375 3120
rect 18395 3100 18400 3120
rect 18370 3070 18400 3100
rect 18370 3050 18375 3070
rect 18395 3050 18400 3070
rect 18370 3020 18400 3050
rect 18370 3000 18375 3020
rect 18395 3000 18400 3020
rect 18370 2990 18400 3000
rect 18425 3570 18455 3580
rect 18425 3550 18430 3570
rect 18450 3550 18455 3570
rect 18425 3520 18455 3550
rect 18425 3500 18430 3520
rect 18450 3500 18455 3520
rect 18425 3470 18455 3500
rect 18425 3450 18430 3470
rect 18450 3450 18455 3470
rect 18425 3420 18455 3450
rect 18425 3400 18430 3420
rect 18450 3400 18455 3420
rect 18425 3370 18455 3400
rect 18425 3350 18430 3370
rect 18450 3350 18455 3370
rect 18425 3320 18455 3350
rect 18425 3300 18430 3320
rect 18450 3300 18455 3320
rect 18425 3270 18455 3300
rect 18425 3250 18430 3270
rect 18450 3250 18455 3270
rect 18425 3220 18455 3250
rect 18425 3200 18430 3220
rect 18450 3200 18455 3220
rect 18425 3170 18455 3200
rect 18425 3150 18430 3170
rect 18450 3150 18455 3170
rect 18425 3120 18455 3150
rect 18425 3100 18430 3120
rect 18450 3100 18455 3120
rect 18425 3070 18455 3100
rect 18425 3050 18430 3070
rect 18450 3050 18455 3070
rect 18425 3020 18455 3050
rect 18425 3000 18430 3020
rect 18450 3000 18455 3020
rect 18425 2990 18455 3000
rect 18480 3570 18510 3580
rect 18480 3550 18485 3570
rect 18505 3550 18510 3570
rect 18480 3520 18510 3550
rect 18480 3500 18485 3520
rect 18505 3500 18510 3520
rect 18480 3470 18510 3500
rect 18480 3450 18485 3470
rect 18505 3450 18510 3470
rect 18480 3420 18510 3450
rect 18480 3400 18485 3420
rect 18505 3400 18510 3420
rect 18480 3370 18510 3400
rect 18480 3350 18485 3370
rect 18505 3350 18510 3370
rect 18480 3320 18510 3350
rect 18480 3300 18485 3320
rect 18505 3300 18510 3320
rect 18480 3270 18510 3300
rect 18480 3250 18485 3270
rect 18505 3250 18510 3270
rect 18480 3220 18510 3250
rect 18480 3200 18485 3220
rect 18505 3200 18510 3220
rect 18480 3170 18510 3200
rect 18480 3150 18485 3170
rect 18505 3150 18510 3170
rect 18480 3120 18510 3150
rect 18480 3100 18485 3120
rect 18505 3100 18510 3120
rect 18480 3070 18510 3100
rect 18480 3050 18485 3070
rect 18505 3050 18510 3070
rect 18480 3020 18510 3050
rect 18480 3000 18485 3020
rect 18505 3000 18510 3020
rect 18480 2990 18510 3000
rect 18535 3570 18565 3580
rect 18535 3550 18540 3570
rect 18560 3550 18565 3570
rect 18535 3520 18565 3550
rect 18535 3500 18540 3520
rect 18560 3500 18565 3520
rect 18535 3470 18565 3500
rect 18535 3450 18540 3470
rect 18560 3450 18565 3470
rect 18535 3420 18565 3450
rect 18535 3400 18540 3420
rect 18560 3400 18565 3420
rect 18535 3370 18565 3400
rect 18535 3350 18540 3370
rect 18560 3350 18565 3370
rect 18535 3320 18565 3350
rect 18535 3300 18540 3320
rect 18560 3300 18565 3320
rect 18535 3270 18565 3300
rect 18535 3250 18540 3270
rect 18560 3250 18565 3270
rect 18535 3220 18565 3250
rect 18535 3200 18540 3220
rect 18560 3200 18565 3220
rect 18535 3170 18565 3200
rect 18535 3150 18540 3170
rect 18560 3150 18565 3170
rect 18535 3120 18565 3150
rect 18535 3100 18540 3120
rect 18560 3100 18565 3120
rect 18535 3070 18565 3100
rect 18535 3050 18540 3070
rect 18560 3050 18565 3070
rect 18535 3020 18565 3050
rect 18535 3000 18540 3020
rect 18560 3000 18565 3020
rect 18535 2990 18565 3000
rect 18590 3570 18620 3580
rect 18590 3550 18595 3570
rect 18615 3550 18620 3570
rect 18590 3520 18620 3550
rect 18590 3500 18595 3520
rect 18615 3500 18620 3520
rect 18590 3470 18620 3500
rect 18590 3450 18595 3470
rect 18615 3450 18620 3470
rect 18590 3420 18620 3450
rect 18590 3400 18595 3420
rect 18615 3400 18620 3420
rect 18590 3370 18620 3400
rect 18590 3350 18595 3370
rect 18615 3350 18620 3370
rect 18590 3320 18620 3350
rect 18590 3300 18595 3320
rect 18615 3300 18620 3320
rect 18590 3270 18620 3300
rect 18590 3250 18595 3270
rect 18615 3250 18620 3270
rect 18590 3220 18620 3250
rect 18590 3200 18595 3220
rect 18615 3200 18620 3220
rect 18590 3170 18620 3200
rect 18590 3150 18595 3170
rect 18615 3150 18620 3170
rect 18590 3120 18620 3150
rect 18590 3100 18595 3120
rect 18615 3100 18620 3120
rect 18590 3070 18620 3100
rect 18590 3050 18595 3070
rect 18615 3050 18620 3070
rect 18590 3020 18620 3050
rect 18590 3000 18595 3020
rect 18615 3000 18620 3020
rect 18590 2990 18620 3000
rect 18645 3570 18675 3580
rect 18645 3550 18650 3570
rect 18670 3550 18675 3570
rect 18645 3520 18675 3550
rect 18645 3500 18650 3520
rect 18670 3500 18675 3520
rect 18645 3470 18675 3500
rect 18645 3450 18650 3470
rect 18670 3450 18675 3470
rect 18645 3420 18675 3450
rect 18645 3400 18650 3420
rect 18670 3400 18675 3420
rect 18645 3370 18675 3400
rect 18645 3350 18650 3370
rect 18670 3350 18675 3370
rect 18645 3320 18675 3350
rect 18645 3300 18650 3320
rect 18670 3300 18675 3320
rect 18645 3270 18675 3300
rect 18645 3250 18650 3270
rect 18670 3250 18675 3270
rect 18645 3220 18675 3250
rect 18645 3200 18650 3220
rect 18670 3200 18675 3220
rect 18645 3170 18675 3200
rect 18645 3150 18650 3170
rect 18670 3150 18675 3170
rect 18645 3120 18675 3150
rect 18645 3100 18650 3120
rect 18670 3100 18675 3120
rect 18645 3070 18675 3100
rect 18645 3050 18650 3070
rect 18670 3050 18675 3070
rect 18645 3020 18675 3050
rect 18645 3000 18650 3020
rect 18670 3000 18675 3020
rect 18645 2990 18675 3000
rect 18700 3570 18730 3580
rect 18700 3550 18705 3570
rect 18725 3550 18730 3570
rect 18700 3520 18730 3550
rect 18700 3500 18705 3520
rect 18725 3500 18730 3520
rect 18700 3470 18730 3500
rect 18700 3450 18705 3470
rect 18725 3450 18730 3470
rect 18700 3420 18730 3450
rect 18700 3400 18705 3420
rect 18725 3400 18730 3420
rect 18700 3370 18730 3400
rect 18700 3350 18705 3370
rect 18725 3350 18730 3370
rect 18700 3320 18730 3350
rect 18700 3300 18705 3320
rect 18725 3300 18730 3320
rect 18700 3270 18730 3300
rect 18700 3250 18705 3270
rect 18725 3250 18730 3270
rect 18700 3220 18730 3250
rect 18700 3200 18705 3220
rect 18725 3200 18730 3220
rect 18700 3170 18730 3200
rect 18700 3150 18705 3170
rect 18725 3150 18730 3170
rect 18700 3120 18730 3150
rect 18700 3100 18705 3120
rect 18725 3100 18730 3120
rect 18700 3070 18730 3100
rect 18700 3050 18705 3070
rect 18725 3050 18730 3070
rect 18700 3020 18730 3050
rect 18700 3000 18705 3020
rect 18725 3000 18730 3020
rect 18700 2990 18730 3000
rect 18755 3570 18785 3580
rect 18755 3550 18760 3570
rect 18780 3550 18785 3570
rect 18755 3520 18785 3550
rect 18755 3500 18760 3520
rect 18780 3500 18785 3520
rect 18755 3470 18785 3500
rect 18755 3450 18760 3470
rect 18780 3450 18785 3470
rect 18755 3420 18785 3450
rect 18755 3400 18760 3420
rect 18780 3400 18785 3420
rect 18755 3370 18785 3400
rect 18755 3350 18760 3370
rect 18780 3350 18785 3370
rect 18755 3320 18785 3350
rect 18755 3300 18760 3320
rect 18780 3300 18785 3320
rect 18755 3270 18785 3300
rect 18755 3250 18760 3270
rect 18780 3250 18785 3270
rect 18755 3220 18785 3250
rect 18755 3200 18760 3220
rect 18780 3200 18785 3220
rect 18755 3170 18785 3200
rect 18755 3150 18760 3170
rect 18780 3150 18785 3170
rect 18755 3120 18785 3150
rect 18755 3100 18760 3120
rect 18780 3100 18785 3120
rect 18755 3070 18785 3100
rect 18755 3050 18760 3070
rect 18780 3050 18785 3070
rect 18755 3020 18785 3050
rect 18755 3000 18760 3020
rect 18780 3000 18785 3020
rect 18755 2990 18785 3000
rect 18810 3570 18880 3580
rect 18810 3550 18815 3570
rect 18835 3550 18855 3570
rect 18875 3550 18880 3570
rect 24970 3570 25040 3580
rect 18810 3520 18880 3550
rect 18810 3500 18815 3520
rect 18835 3500 18855 3520
rect 18875 3500 18880 3520
rect 18810 3470 18880 3500
rect 18810 3450 18815 3470
rect 18835 3450 18855 3470
rect 18875 3450 18880 3470
rect 18810 3420 18880 3450
rect 18810 3400 18815 3420
rect 18835 3400 18855 3420
rect 18875 3400 18880 3420
rect 18810 3370 18880 3400
rect 18810 3350 18815 3370
rect 18835 3350 18855 3370
rect 18875 3350 18880 3370
rect 18810 3320 18880 3350
rect 18810 3300 18815 3320
rect 18835 3300 18855 3320
rect 18875 3300 18880 3320
rect 19105 3520 19246 3560
rect 24554 3520 24695 3560
rect 24970 3550 24975 3570
rect 24995 3550 25015 3570
rect 25035 3550 25040 3570
rect 24970 3520 25040 3550
rect 24970 3500 24975 3520
rect 24995 3500 25015 3520
rect 25035 3500 25040 3520
rect 24970 3470 25040 3500
rect 24970 3450 24975 3470
rect 24995 3450 25015 3470
rect 25035 3450 25040 3470
rect 24970 3420 25040 3450
rect 24970 3400 24975 3420
rect 24995 3400 25015 3420
rect 25035 3400 25040 3420
rect 24970 3370 25040 3400
rect 24970 3350 24975 3370
rect 24995 3350 25015 3370
rect 25035 3350 25040 3370
rect 24970 3320 25040 3350
rect 24970 3300 24975 3320
rect 24995 3300 25015 3320
rect 25035 3300 25040 3320
rect 18810 3270 18880 3300
rect 18810 3250 18815 3270
rect 18835 3250 18855 3270
rect 18875 3250 18880 3270
rect 18810 3220 18880 3250
rect 18810 3200 18815 3220
rect 18835 3200 18855 3220
rect 18875 3200 18880 3220
rect 18810 3170 18880 3200
rect 18810 3150 18815 3170
rect 18835 3150 18855 3170
rect 18875 3150 18880 3170
rect 24970 3270 25040 3300
rect 24970 3250 24975 3270
rect 24995 3250 25015 3270
rect 25035 3250 25040 3270
rect 24970 3220 25040 3250
rect 24970 3200 24975 3220
rect 24995 3200 25015 3220
rect 25035 3200 25040 3220
rect 24970 3170 25040 3200
rect 18810 3120 18880 3150
rect 18810 3100 18815 3120
rect 18835 3100 18855 3120
rect 18875 3100 18880 3120
rect 18810 3070 18880 3100
rect 18810 3050 18815 3070
rect 18835 3050 18855 3070
rect 18875 3050 18880 3070
rect 18810 3020 18880 3050
rect 18810 3000 18815 3020
rect 18835 3000 18855 3020
rect 18875 3000 18880 3020
rect 18810 2990 18880 3000
rect 14975 2970 14995 2990
rect 15125 2970 15145 2990
rect 15235 2970 15255 2990
rect 15345 2970 15365 2990
rect 15455 2970 15475 2990
rect 15565 2970 15585 2990
rect 15715 2970 15735 2990
rect 18115 2970 18135 2990
rect 18265 2970 18285 2990
rect 18375 2970 18395 2990
rect 18485 2970 18505 2990
rect 18595 2970 18615 2990
rect 18705 2970 18725 2990
rect 18855 2970 18875 2990
rect 2960 2915 3030 2925
rect 1266 2865 1306 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2960 2895 2965 2915
rect 2985 2895 3005 2915
rect 3025 2895 3030 2915
rect 2960 2865 3030 2895
rect -55 2825 -25 2855
rect 51 2850 96 2855
rect 51 2825 61 2850
rect 86 2825 96 2850
rect 51 2820 96 2825
rect 724 2850 769 2855
rect 724 2825 734 2850
rect 759 2825 769 2850
rect 724 2820 769 2825
rect 1210 2820 1240 2850
rect 2960 2845 2965 2865
rect 2985 2845 3005 2865
rect 3025 2845 3030 2865
rect 1261 2835 1306 2840
rect 1261 2810 1271 2835
rect 1296 2810 1306 2835
rect 1261 2805 1306 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2960 2835 3030 2845
rect 3090 2915 3120 2925
rect 3090 2895 3095 2915
rect 3115 2895 3120 2915
rect 3090 2865 3120 2895
rect 3090 2845 3095 2865
rect 3115 2845 3120 2865
rect 3090 2835 3120 2845
rect 3180 2915 3210 2925
rect 3180 2895 3185 2915
rect 3205 2895 3210 2915
rect 3180 2865 3210 2895
rect 3180 2845 3185 2865
rect 3205 2845 3210 2865
rect 3180 2835 3210 2845
rect 3270 2915 3300 2925
rect 3270 2895 3275 2915
rect 3295 2895 3300 2915
rect 3270 2865 3300 2895
rect 3270 2845 3275 2865
rect 3295 2845 3300 2865
rect 3270 2835 3300 2845
rect 3360 2915 3390 2925
rect 3360 2895 3365 2915
rect 3385 2895 3390 2915
rect 3360 2865 3390 2895
rect 3360 2845 3365 2865
rect 3385 2845 3390 2865
rect 3360 2835 3390 2845
rect 3450 2915 3480 2925
rect 3450 2895 3455 2915
rect 3475 2895 3480 2915
rect 3450 2865 3480 2895
rect 3450 2845 3455 2865
rect 3475 2845 3480 2865
rect 3450 2835 3480 2845
rect 3540 2915 3570 2925
rect 3540 2895 3545 2915
rect 3565 2895 3570 2915
rect 3540 2865 3570 2895
rect 3540 2845 3545 2865
rect 3565 2845 3570 2865
rect 3540 2835 3570 2845
rect 3630 2915 3660 2925
rect 3630 2895 3635 2915
rect 3655 2895 3660 2915
rect 3630 2865 3660 2895
rect 3630 2845 3635 2865
rect 3655 2845 3660 2865
rect 3630 2835 3660 2845
rect 3720 2915 3750 2925
rect 3720 2895 3725 2915
rect 3745 2895 3750 2915
rect 3720 2865 3750 2895
rect 3720 2845 3725 2865
rect 3745 2845 3750 2865
rect 3720 2835 3750 2845
rect 3810 2915 3840 2925
rect 3810 2895 3815 2915
rect 3835 2895 3840 2915
rect 3810 2865 3840 2895
rect 3810 2845 3815 2865
rect 3835 2845 3840 2865
rect 3810 2835 3840 2845
rect 3900 2915 3930 2925
rect 3900 2895 3905 2915
rect 3925 2895 3930 2915
rect 3900 2865 3930 2895
rect 3900 2845 3905 2865
rect 3925 2845 3930 2865
rect 3900 2835 3930 2845
rect 3990 2915 4020 2925
rect 3990 2895 3995 2915
rect 4015 2895 4020 2915
rect 3990 2865 4020 2895
rect 3990 2845 3995 2865
rect 4015 2845 4020 2865
rect 3990 2835 4020 2845
rect 4080 2915 4110 2925
rect 4080 2895 4085 2915
rect 4105 2895 4110 2915
rect 4080 2865 4110 2895
rect 4080 2845 4085 2865
rect 4105 2845 4110 2865
rect 4080 2835 4110 2845
rect 4170 2915 4200 2925
rect 4170 2895 4175 2915
rect 4195 2895 4200 2915
rect 4170 2865 4200 2895
rect 4170 2845 4175 2865
rect 4195 2845 4200 2865
rect 4170 2835 4200 2845
rect 4260 2915 4290 2925
rect 4260 2895 4265 2915
rect 4285 2895 4290 2915
rect 4260 2865 4290 2895
rect 4260 2845 4265 2865
rect 4285 2845 4290 2865
rect 4260 2835 4290 2845
rect 4350 2915 4380 2925
rect 4350 2895 4355 2915
rect 4375 2895 4380 2915
rect 4350 2865 4380 2895
rect 4350 2845 4355 2865
rect 4375 2845 4380 2865
rect 4350 2835 4380 2845
rect 4440 2915 4470 2925
rect 4440 2895 4445 2915
rect 4465 2895 4470 2915
rect 4440 2865 4470 2895
rect 4440 2845 4445 2865
rect 4465 2845 4470 2865
rect 4440 2835 4470 2845
rect 4530 2915 4560 2925
rect 4530 2895 4535 2915
rect 4555 2895 4560 2915
rect 4530 2865 4560 2895
rect 4530 2845 4535 2865
rect 4555 2845 4560 2865
rect 4530 2835 4560 2845
rect 4620 2915 4650 2925
rect 4620 2895 4625 2915
rect 4645 2895 4650 2915
rect 4620 2865 4650 2895
rect 4620 2845 4625 2865
rect 4645 2845 4650 2865
rect 4620 2835 4650 2845
rect 4710 2915 4740 2925
rect 4710 2895 4715 2915
rect 4735 2895 4740 2915
rect 4710 2865 4740 2895
rect 4710 2845 4715 2865
rect 4735 2845 4740 2865
rect 4710 2835 4740 2845
rect 4800 2915 4830 2925
rect 4800 2895 4805 2915
rect 4825 2895 4830 2915
rect 4800 2865 4830 2895
rect 4800 2845 4805 2865
rect 4825 2845 4830 2865
rect 4800 2835 4830 2845
rect 4890 2915 4920 2925
rect 4890 2895 4895 2915
rect 4915 2895 4920 2915
rect 4890 2865 4920 2895
rect 4890 2845 4895 2865
rect 4915 2845 4920 2865
rect 4890 2835 4920 2845
rect 4980 2915 5050 2925
rect 4980 2895 4985 2915
rect 5005 2895 5025 2915
rect 5045 2895 5050 2915
rect 14554 2900 14695 2940
rect 14965 2960 15005 2970
rect 14965 2940 14975 2960
rect 14995 2940 15005 2960
rect 14965 2930 15005 2940
rect 15115 2960 15155 2970
rect 15115 2940 15125 2960
rect 15145 2940 15155 2960
rect 15115 2930 15155 2940
rect 15225 2960 15265 2970
rect 15225 2940 15235 2960
rect 15255 2940 15265 2960
rect 15225 2930 15265 2940
rect 15335 2960 15375 2970
rect 15335 2940 15345 2960
rect 15365 2940 15375 2960
rect 15335 2930 15375 2940
rect 15445 2960 15485 2970
rect 15445 2940 15455 2960
rect 15475 2940 15485 2960
rect 15445 2930 15485 2940
rect 15503 2960 15537 2970
rect 15503 2940 15511 2960
rect 15529 2940 15537 2960
rect 15503 2930 15537 2940
rect 15555 2960 15595 2970
rect 15555 2940 15565 2960
rect 15585 2940 15595 2960
rect 15555 2930 15595 2940
rect 15705 2960 15745 2970
rect 15705 2940 15715 2960
rect 15735 2940 15745 2960
rect 15705 2930 15745 2940
rect 18105 2960 18145 2970
rect 18105 2940 18115 2960
rect 18135 2940 18145 2960
rect 18105 2930 18145 2940
rect 18255 2960 18295 2970
rect 18255 2940 18265 2960
rect 18285 2940 18295 2960
rect 18255 2930 18295 2940
rect 18313 2960 18347 2970
rect 18313 2940 18321 2960
rect 18339 2940 18347 2960
rect 18313 2930 18347 2940
rect 18365 2960 18405 2970
rect 18365 2940 18375 2960
rect 18395 2940 18405 2960
rect 18365 2930 18405 2940
rect 18475 2960 18515 2970
rect 18475 2940 18485 2960
rect 18505 2940 18515 2960
rect 18475 2930 18515 2940
rect 18585 2960 18625 2970
rect 18585 2940 18595 2960
rect 18615 2940 18625 2960
rect 18585 2930 18625 2940
rect 18695 2960 18735 2970
rect 18695 2940 18705 2960
rect 18725 2940 18735 2960
rect 18695 2930 18735 2940
rect 18845 2960 18885 2970
rect 18845 2940 18855 2960
rect 18875 2940 18885 2960
rect 18845 2930 18885 2940
rect 19105 2900 19246 2940
rect 24970 3150 24975 3170
rect 24995 3150 25015 3170
rect 25035 3150 25040 3170
rect 24970 3120 25040 3150
rect 24970 3100 24975 3120
rect 24995 3100 25015 3120
rect 25035 3100 25040 3120
rect 24970 3070 25040 3100
rect 24970 3050 24975 3070
rect 24995 3050 25015 3070
rect 25035 3050 25040 3070
rect 24970 3020 25040 3050
rect 24970 3000 24975 3020
rect 24995 3000 25015 3020
rect 25035 3000 25040 3020
rect 24970 2990 25040 3000
rect 25065 3570 25095 3580
rect 25065 3550 25070 3570
rect 25090 3550 25095 3570
rect 25065 3520 25095 3550
rect 25065 3500 25070 3520
rect 25090 3500 25095 3520
rect 25065 3470 25095 3500
rect 25065 3450 25070 3470
rect 25090 3450 25095 3470
rect 25065 3420 25095 3450
rect 25065 3400 25070 3420
rect 25090 3400 25095 3420
rect 25065 3370 25095 3400
rect 25065 3350 25070 3370
rect 25090 3350 25095 3370
rect 25065 3320 25095 3350
rect 25065 3300 25070 3320
rect 25090 3300 25095 3320
rect 25065 3270 25095 3300
rect 25065 3250 25070 3270
rect 25090 3250 25095 3270
rect 25065 3220 25095 3250
rect 25065 3200 25070 3220
rect 25090 3200 25095 3220
rect 25065 3170 25095 3200
rect 25065 3150 25070 3170
rect 25090 3150 25095 3170
rect 25065 3120 25095 3150
rect 25065 3100 25070 3120
rect 25090 3100 25095 3120
rect 25065 3070 25095 3100
rect 25065 3050 25070 3070
rect 25090 3050 25095 3070
rect 25065 3020 25095 3050
rect 25065 3000 25070 3020
rect 25090 3000 25095 3020
rect 25065 2990 25095 3000
rect 25120 3570 25150 3580
rect 25120 3550 25125 3570
rect 25145 3550 25150 3570
rect 25120 3520 25150 3550
rect 25120 3500 25125 3520
rect 25145 3500 25150 3520
rect 25120 3470 25150 3500
rect 25120 3450 25125 3470
rect 25145 3450 25150 3470
rect 25120 3420 25150 3450
rect 25120 3400 25125 3420
rect 25145 3400 25150 3420
rect 25120 3370 25150 3400
rect 25120 3350 25125 3370
rect 25145 3350 25150 3370
rect 25120 3320 25150 3350
rect 25120 3300 25125 3320
rect 25145 3300 25150 3320
rect 25120 3270 25150 3300
rect 25120 3250 25125 3270
rect 25145 3250 25150 3270
rect 25120 3220 25150 3250
rect 25120 3200 25125 3220
rect 25145 3200 25150 3220
rect 25120 3170 25150 3200
rect 25120 3150 25125 3170
rect 25145 3150 25150 3170
rect 25120 3120 25150 3150
rect 25120 3100 25125 3120
rect 25145 3100 25150 3120
rect 25120 3070 25150 3100
rect 25120 3050 25125 3070
rect 25145 3050 25150 3070
rect 25120 3020 25150 3050
rect 25120 3000 25125 3020
rect 25145 3000 25150 3020
rect 25120 2990 25150 3000
rect 25175 3570 25205 3580
rect 25175 3550 25180 3570
rect 25200 3550 25205 3570
rect 25175 3520 25205 3550
rect 25175 3500 25180 3520
rect 25200 3500 25205 3520
rect 25175 3470 25205 3500
rect 25175 3450 25180 3470
rect 25200 3450 25205 3470
rect 25175 3420 25205 3450
rect 25175 3400 25180 3420
rect 25200 3400 25205 3420
rect 25175 3370 25205 3400
rect 25175 3350 25180 3370
rect 25200 3350 25205 3370
rect 25175 3320 25205 3350
rect 25175 3300 25180 3320
rect 25200 3300 25205 3320
rect 25175 3270 25205 3300
rect 25175 3250 25180 3270
rect 25200 3250 25205 3270
rect 25175 3220 25205 3250
rect 25175 3200 25180 3220
rect 25200 3200 25205 3220
rect 25175 3170 25205 3200
rect 25175 3150 25180 3170
rect 25200 3150 25205 3170
rect 25175 3120 25205 3150
rect 25175 3100 25180 3120
rect 25200 3100 25205 3120
rect 25175 3070 25205 3100
rect 25175 3050 25180 3070
rect 25200 3050 25205 3070
rect 25175 3020 25205 3050
rect 25175 3000 25180 3020
rect 25200 3000 25205 3020
rect 25175 2990 25205 3000
rect 25230 3570 25260 3580
rect 25230 3550 25235 3570
rect 25255 3550 25260 3570
rect 25230 3520 25260 3550
rect 25230 3500 25235 3520
rect 25255 3500 25260 3520
rect 25230 3470 25260 3500
rect 25230 3450 25235 3470
rect 25255 3450 25260 3470
rect 25230 3420 25260 3450
rect 25230 3400 25235 3420
rect 25255 3400 25260 3420
rect 25230 3370 25260 3400
rect 25230 3350 25235 3370
rect 25255 3350 25260 3370
rect 25230 3320 25260 3350
rect 25230 3300 25235 3320
rect 25255 3300 25260 3320
rect 25230 3270 25260 3300
rect 25230 3250 25235 3270
rect 25255 3250 25260 3270
rect 25230 3220 25260 3250
rect 25230 3200 25235 3220
rect 25255 3200 25260 3220
rect 25230 3170 25260 3200
rect 25230 3150 25235 3170
rect 25255 3150 25260 3170
rect 25230 3120 25260 3150
rect 25230 3100 25235 3120
rect 25255 3100 25260 3120
rect 25230 3070 25260 3100
rect 25230 3050 25235 3070
rect 25255 3050 25260 3070
rect 25230 3020 25260 3050
rect 25230 3000 25235 3020
rect 25255 3000 25260 3020
rect 25230 2990 25260 3000
rect 25285 3570 25315 3580
rect 25285 3550 25290 3570
rect 25310 3550 25315 3570
rect 25285 3520 25315 3550
rect 25285 3500 25290 3520
rect 25310 3500 25315 3520
rect 25285 3470 25315 3500
rect 25285 3450 25290 3470
rect 25310 3450 25315 3470
rect 25285 3420 25315 3450
rect 25285 3400 25290 3420
rect 25310 3400 25315 3420
rect 25285 3370 25315 3400
rect 25285 3350 25290 3370
rect 25310 3350 25315 3370
rect 25285 3320 25315 3350
rect 25285 3300 25290 3320
rect 25310 3300 25315 3320
rect 25285 3270 25315 3300
rect 25285 3250 25290 3270
rect 25310 3250 25315 3270
rect 25285 3220 25315 3250
rect 25285 3200 25290 3220
rect 25310 3200 25315 3220
rect 25285 3170 25315 3200
rect 25285 3150 25290 3170
rect 25310 3150 25315 3170
rect 25285 3120 25315 3150
rect 25285 3100 25290 3120
rect 25310 3100 25315 3120
rect 25285 3070 25315 3100
rect 25285 3050 25290 3070
rect 25310 3050 25315 3070
rect 25285 3020 25315 3050
rect 25285 3000 25290 3020
rect 25310 3000 25315 3020
rect 25285 2990 25315 3000
rect 25340 3570 25370 3580
rect 25340 3550 25345 3570
rect 25365 3550 25370 3570
rect 25340 3520 25370 3550
rect 25340 3500 25345 3520
rect 25365 3500 25370 3520
rect 25340 3470 25370 3500
rect 25340 3450 25345 3470
rect 25365 3450 25370 3470
rect 25340 3420 25370 3450
rect 25340 3400 25345 3420
rect 25365 3400 25370 3420
rect 25340 3370 25370 3400
rect 25340 3350 25345 3370
rect 25365 3350 25370 3370
rect 25340 3320 25370 3350
rect 25340 3300 25345 3320
rect 25365 3300 25370 3320
rect 25340 3270 25370 3300
rect 25340 3250 25345 3270
rect 25365 3250 25370 3270
rect 25340 3220 25370 3250
rect 25340 3200 25345 3220
rect 25365 3200 25370 3220
rect 25340 3170 25370 3200
rect 25340 3150 25345 3170
rect 25365 3150 25370 3170
rect 25340 3120 25370 3150
rect 25340 3100 25345 3120
rect 25365 3100 25370 3120
rect 25340 3070 25370 3100
rect 25340 3050 25345 3070
rect 25365 3050 25370 3070
rect 25340 3020 25370 3050
rect 25340 3000 25345 3020
rect 25365 3000 25370 3020
rect 25340 2990 25370 3000
rect 25395 3570 25425 3580
rect 25395 3550 25400 3570
rect 25420 3550 25425 3570
rect 25395 3520 25425 3550
rect 25395 3500 25400 3520
rect 25420 3500 25425 3520
rect 25395 3470 25425 3500
rect 25395 3450 25400 3470
rect 25420 3450 25425 3470
rect 25395 3420 25425 3450
rect 25395 3400 25400 3420
rect 25420 3400 25425 3420
rect 25395 3370 25425 3400
rect 25395 3350 25400 3370
rect 25420 3350 25425 3370
rect 25395 3320 25425 3350
rect 25395 3300 25400 3320
rect 25420 3300 25425 3320
rect 25395 3270 25425 3300
rect 25395 3250 25400 3270
rect 25420 3250 25425 3270
rect 25395 3220 25425 3250
rect 25395 3200 25400 3220
rect 25420 3200 25425 3220
rect 25395 3170 25425 3200
rect 25395 3150 25400 3170
rect 25420 3150 25425 3170
rect 25395 3120 25425 3150
rect 25395 3100 25400 3120
rect 25420 3100 25425 3120
rect 25395 3070 25425 3100
rect 25395 3050 25400 3070
rect 25420 3050 25425 3070
rect 25395 3020 25425 3050
rect 25395 3000 25400 3020
rect 25420 3000 25425 3020
rect 25395 2990 25425 3000
rect 25450 3570 25480 3580
rect 25450 3550 25455 3570
rect 25475 3550 25480 3570
rect 25450 3520 25480 3550
rect 25450 3500 25455 3520
rect 25475 3500 25480 3520
rect 25450 3470 25480 3500
rect 25450 3450 25455 3470
rect 25475 3450 25480 3470
rect 25450 3420 25480 3450
rect 25450 3400 25455 3420
rect 25475 3400 25480 3420
rect 25450 3370 25480 3400
rect 25450 3350 25455 3370
rect 25475 3350 25480 3370
rect 25450 3320 25480 3350
rect 25450 3300 25455 3320
rect 25475 3300 25480 3320
rect 25450 3270 25480 3300
rect 25450 3250 25455 3270
rect 25475 3250 25480 3270
rect 25450 3220 25480 3250
rect 25450 3200 25455 3220
rect 25475 3200 25480 3220
rect 25450 3170 25480 3200
rect 25450 3150 25455 3170
rect 25475 3150 25480 3170
rect 25450 3120 25480 3150
rect 25450 3100 25455 3120
rect 25475 3100 25480 3120
rect 25450 3070 25480 3100
rect 25450 3050 25455 3070
rect 25475 3050 25480 3070
rect 25450 3020 25480 3050
rect 25450 3000 25455 3020
rect 25475 3000 25480 3020
rect 25450 2990 25480 3000
rect 25505 3570 25535 3580
rect 25505 3550 25510 3570
rect 25530 3550 25535 3570
rect 25505 3520 25535 3550
rect 25505 3500 25510 3520
rect 25530 3500 25535 3520
rect 25505 3470 25535 3500
rect 25505 3450 25510 3470
rect 25530 3450 25535 3470
rect 25505 3420 25535 3450
rect 25505 3400 25510 3420
rect 25530 3400 25535 3420
rect 25505 3370 25535 3400
rect 25505 3350 25510 3370
rect 25530 3350 25535 3370
rect 25505 3320 25535 3350
rect 25505 3300 25510 3320
rect 25530 3300 25535 3320
rect 25505 3270 25535 3300
rect 25505 3250 25510 3270
rect 25530 3250 25535 3270
rect 25505 3220 25535 3250
rect 25505 3200 25510 3220
rect 25530 3200 25535 3220
rect 25505 3170 25535 3200
rect 25505 3150 25510 3170
rect 25530 3150 25535 3170
rect 25505 3120 25535 3150
rect 25505 3100 25510 3120
rect 25530 3100 25535 3120
rect 25505 3070 25535 3100
rect 25505 3050 25510 3070
rect 25530 3050 25535 3070
rect 25505 3020 25535 3050
rect 25505 3000 25510 3020
rect 25530 3000 25535 3020
rect 25505 2990 25535 3000
rect 25560 3570 25590 3580
rect 25560 3550 25565 3570
rect 25585 3550 25590 3570
rect 25560 3520 25590 3550
rect 25560 3500 25565 3520
rect 25585 3500 25590 3520
rect 25560 3470 25590 3500
rect 25560 3450 25565 3470
rect 25585 3450 25590 3470
rect 25560 3420 25590 3450
rect 25560 3400 25565 3420
rect 25585 3400 25590 3420
rect 25560 3370 25590 3400
rect 25560 3350 25565 3370
rect 25585 3350 25590 3370
rect 25560 3320 25590 3350
rect 25560 3300 25565 3320
rect 25585 3300 25590 3320
rect 25560 3270 25590 3300
rect 25560 3250 25565 3270
rect 25585 3250 25590 3270
rect 25560 3220 25590 3250
rect 25560 3200 25565 3220
rect 25585 3200 25590 3220
rect 25560 3170 25590 3200
rect 25560 3150 25565 3170
rect 25585 3150 25590 3170
rect 25560 3120 25590 3150
rect 25560 3100 25565 3120
rect 25585 3100 25590 3120
rect 25560 3070 25590 3100
rect 25560 3050 25565 3070
rect 25585 3050 25590 3070
rect 25560 3020 25590 3050
rect 25560 3000 25565 3020
rect 25585 3000 25590 3020
rect 25560 2990 25590 3000
rect 25615 3570 25645 3580
rect 25615 3550 25620 3570
rect 25640 3550 25645 3570
rect 25615 3520 25645 3550
rect 25615 3500 25620 3520
rect 25640 3500 25645 3520
rect 25615 3470 25645 3500
rect 25615 3450 25620 3470
rect 25640 3450 25645 3470
rect 25615 3420 25645 3450
rect 25615 3400 25620 3420
rect 25640 3400 25645 3420
rect 25615 3370 25645 3400
rect 25615 3350 25620 3370
rect 25640 3350 25645 3370
rect 25615 3320 25645 3350
rect 25615 3300 25620 3320
rect 25640 3300 25645 3320
rect 25615 3270 25645 3300
rect 25615 3250 25620 3270
rect 25640 3250 25645 3270
rect 25615 3220 25645 3250
rect 25615 3200 25620 3220
rect 25640 3200 25645 3220
rect 25615 3170 25645 3200
rect 25615 3150 25620 3170
rect 25640 3150 25645 3170
rect 25615 3120 25645 3150
rect 25615 3100 25620 3120
rect 25640 3100 25645 3120
rect 25615 3070 25645 3100
rect 25615 3050 25620 3070
rect 25640 3050 25645 3070
rect 25615 3020 25645 3050
rect 25615 3000 25620 3020
rect 25640 3000 25645 3020
rect 25615 2990 25645 3000
rect 25670 3570 25740 3580
rect 25670 3550 25675 3570
rect 25695 3550 25715 3570
rect 25735 3550 25740 3570
rect 25670 3520 25740 3550
rect 25670 3500 25675 3520
rect 25695 3500 25715 3520
rect 25735 3500 25740 3520
rect 25670 3470 25740 3500
rect 25670 3450 25675 3470
rect 25695 3450 25715 3470
rect 25735 3450 25740 3470
rect 25670 3420 25740 3450
rect 25670 3400 25675 3420
rect 25695 3400 25715 3420
rect 25735 3400 25740 3420
rect 25670 3370 25740 3400
rect 25670 3350 25675 3370
rect 25695 3350 25715 3370
rect 25735 3350 25740 3370
rect 25670 3320 25740 3350
rect 25670 3300 25675 3320
rect 25695 3300 25715 3320
rect 25735 3300 25740 3320
rect 25670 3270 25740 3300
rect 25670 3250 25675 3270
rect 25695 3250 25715 3270
rect 25735 3250 25740 3270
rect 25670 3220 25740 3250
rect 25670 3200 25675 3220
rect 25695 3200 25715 3220
rect 25735 3200 25740 3220
rect 25670 3170 25740 3200
rect 25670 3150 25675 3170
rect 25695 3150 25715 3170
rect 25735 3150 25740 3170
rect 25670 3120 25740 3150
rect 25670 3100 25675 3120
rect 25695 3100 25715 3120
rect 25735 3100 25740 3120
rect 26170 3445 26190 3680
rect 26340 3650 26380 3660
rect 26340 3630 26350 3650
rect 26370 3630 26380 3650
rect 26340 3620 26380 3630
rect 26460 3650 26500 3660
rect 26460 3630 26470 3650
rect 26490 3630 26500 3650
rect 26460 3620 26500 3630
rect 26580 3650 26620 3660
rect 26580 3630 26590 3650
rect 26610 3630 26620 3650
rect 26580 3620 26620 3630
rect 26700 3650 26740 3660
rect 26700 3630 26710 3650
rect 26730 3630 26740 3650
rect 26700 3620 26740 3630
rect 26820 3650 26860 3660
rect 26820 3630 26830 3650
rect 26850 3630 26860 3650
rect 26820 3620 26860 3630
rect 26940 3650 26980 3660
rect 26940 3630 26950 3650
rect 26970 3630 26980 3650
rect 26940 3620 26980 3630
rect 27060 3650 27100 3660
rect 27060 3630 27070 3650
rect 27090 3630 27100 3650
rect 27060 3620 27100 3630
rect 27180 3650 27220 3660
rect 27180 3630 27190 3650
rect 27210 3630 27220 3650
rect 27180 3620 27220 3630
rect 27300 3650 27340 3660
rect 27300 3630 27310 3650
rect 27330 3630 27340 3650
rect 27300 3620 27340 3630
rect 27420 3650 27460 3660
rect 27420 3630 27430 3650
rect 27450 3630 27460 3650
rect 27420 3620 27460 3630
rect 26350 3600 26370 3620
rect 26470 3600 26490 3620
rect 26590 3600 26610 3620
rect 26710 3600 26730 3620
rect 26830 3600 26850 3620
rect 26950 3600 26970 3620
rect 27070 3600 27090 3620
rect 27190 3600 27210 3620
rect 27310 3600 27330 3620
rect 27430 3600 27450 3620
rect 26170 3130 26190 3365
rect 26225 3590 26255 3600
rect 26225 3570 26230 3590
rect 26250 3570 26255 3590
rect 26225 3540 26255 3570
rect 26225 3520 26230 3540
rect 26250 3520 26255 3540
rect 26225 3490 26255 3520
rect 26225 3470 26230 3490
rect 26250 3470 26255 3490
rect 26225 3440 26255 3470
rect 26225 3420 26230 3440
rect 26250 3420 26255 3440
rect 26225 3390 26255 3420
rect 26225 3370 26230 3390
rect 26250 3370 26255 3390
rect 26225 3340 26255 3370
rect 26225 3320 26230 3340
rect 26250 3320 26255 3340
rect 26225 3290 26255 3320
rect 26225 3270 26230 3290
rect 26250 3270 26255 3290
rect 26225 3240 26255 3270
rect 26225 3220 26230 3240
rect 26250 3220 26255 3240
rect 26225 3210 26255 3220
rect 26285 3590 26315 3600
rect 26285 3570 26290 3590
rect 26310 3570 26315 3590
rect 26285 3540 26315 3570
rect 26285 3520 26290 3540
rect 26310 3520 26315 3540
rect 26285 3490 26315 3520
rect 26285 3470 26290 3490
rect 26310 3470 26315 3490
rect 26285 3440 26315 3470
rect 26285 3420 26290 3440
rect 26310 3420 26315 3440
rect 26285 3390 26315 3420
rect 26285 3370 26290 3390
rect 26310 3370 26315 3390
rect 26285 3340 26315 3370
rect 26285 3320 26290 3340
rect 26310 3320 26315 3340
rect 26285 3290 26315 3320
rect 26285 3270 26290 3290
rect 26310 3270 26315 3290
rect 26285 3240 26315 3270
rect 26285 3220 26290 3240
rect 26310 3220 26315 3240
rect 26285 3210 26315 3220
rect 26345 3590 26375 3600
rect 26345 3570 26350 3590
rect 26370 3570 26375 3590
rect 26345 3540 26375 3570
rect 26345 3520 26350 3540
rect 26370 3520 26375 3540
rect 26345 3490 26375 3520
rect 26345 3470 26350 3490
rect 26370 3470 26375 3490
rect 26345 3440 26375 3470
rect 26345 3420 26350 3440
rect 26370 3420 26375 3440
rect 26345 3390 26375 3420
rect 26345 3370 26350 3390
rect 26370 3370 26375 3390
rect 26345 3340 26375 3370
rect 26345 3320 26350 3340
rect 26370 3320 26375 3340
rect 26345 3290 26375 3320
rect 26345 3270 26350 3290
rect 26370 3270 26375 3290
rect 26345 3240 26375 3270
rect 26345 3220 26350 3240
rect 26370 3220 26375 3240
rect 26345 3210 26375 3220
rect 26405 3590 26435 3600
rect 26405 3570 26410 3590
rect 26430 3570 26435 3590
rect 26405 3540 26435 3570
rect 26405 3520 26410 3540
rect 26430 3520 26435 3540
rect 26405 3490 26435 3520
rect 26405 3470 26410 3490
rect 26430 3470 26435 3490
rect 26405 3440 26435 3470
rect 26405 3420 26410 3440
rect 26430 3420 26435 3440
rect 26405 3390 26435 3420
rect 26405 3370 26410 3390
rect 26430 3370 26435 3390
rect 26405 3340 26435 3370
rect 26405 3320 26410 3340
rect 26430 3320 26435 3340
rect 26405 3290 26435 3320
rect 26405 3270 26410 3290
rect 26430 3270 26435 3290
rect 26405 3240 26435 3270
rect 26405 3220 26410 3240
rect 26430 3220 26435 3240
rect 26405 3210 26435 3220
rect 26465 3590 26495 3600
rect 26465 3570 26470 3590
rect 26490 3570 26495 3590
rect 26465 3540 26495 3570
rect 26465 3520 26470 3540
rect 26490 3520 26495 3540
rect 26465 3490 26495 3520
rect 26465 3470 26470 3490
rect 26490 3470 26495 3490
rect 26465 3440 26495 3470
rect 26465 3420 26470 3440
rect 26490 3420 26495 3440
rect 26465 3390 26495 3420
rect 26465 3370 26470 3390
rect 26490 3370 26495 3390
rect 26465 3340 26495 3370
rect 26465 3320 26470 3340
rect 26490 3320 26495 3340
rect 26465 3290 26495 3320
rect 26465 3270 26470 3290
rect 26490 3270 26495 3290
rect 26465 3240 26495 3270
rect 26465 3220 26470 3240
rect 26490 3220 26495 3240
rect 26465 3210 26495 3220
rect 26525 3590 26555 3600
rect 26525 3570 26530 3590
rect 26550 3570 26555 3590
rect 26525 3540 26555 3570
rect 26525 3520 26530 3540
rect 26550 3520 26555 3540
rect 26525 3490 26555 3520
rect 26525 3470 26530 3490
rect 26550 3470 26555 3490
rect 26525 3440 26555 3470
rect 26525 3420 26530 3440
rect 26550 3420 26555 3440
rect 26525 3390 26555 3420
rect 26525 3370 26530 3390
rect 26550 3370 26555 3390
rect 26525 3340 26555 3370
rect 26525 3320 26530 3340
rect 26550 3320 26555 3340
rect 26525 3290 26555 3320
rect 26525 3270 26530 3290
rect 26550 3270 26555 3290
rect 26525 3240 26555 3270
rect 26525 3220 26530 3240
rect 26550 3220 26555 3240
rect 26525 3210 26555 3220
rect 26585 3590 26615 3600
rect 26585 3570 26590 3590
rect 26610 3570 26615 3590
rect 26585 3540 26615 3570
rect 26585 3520 26590 3540
rect 26610 3520 26615 3540
rect 26585 3490 26615 3520
rect 26585 3470 26590 3490
rect 26610 3470 26615 3490
rect 26585 3440 26615 3470
rect 26585 3420 26590 3440
rect 26610 3420 26615 3440
rect 26585 3390 26615 3420
rect 26585 3370 26590 3390
rect 26610 3370 26615 3390
rect 26585 3340 26615 3370
rect 26585 3320 26590 3340
rect 26610 3320 26615 3340
rect 26585 3290 26615 3320
rect 26585 3270 26590 3290
rect 26610 3270 26615 3290
rect 26585 3240 26615 3270
rect 26585 3220 26590 3240
rect 26610 3220 26615 3240
rect 26585 3210 26615 3220
rect 26645 3590 26675 3600
rect 26645 3570 26650 3590
rect 26670 3570 26675 3590
rect 26645 3540 26675 3570
rect 26645 3520 26650 3540
rect 26670 3520 26675 3540
rect 26645 3490 26675 3520
rect 26645 3470 26650 3490
rect 26670 3470 26675 3490
rect 26645 3440 26675 3470
rect 26645 3420 26650 3440
rect 26670 3420 26675 3440
rect 26645 3390 26675 3420
rect 26645 3370 26650 3390
rect 26670 3370 26675 3390
rect 26645 3340 26675 3370
rect 26645 3320 26650 3340
rect 26670 3320 26675 3340
rect 26645 3290 26675 3320
rect 26645 3270 26650 3290
rect 26670 3270 26675 3290
rect 26645 3240 26675 3270
rect 26645 3220 26650 3240
rect 26670 3220 26675 3240
rect 26645 3210 26675 3220
rect 26705 3590 26735 3600
rect 26705 3570 26710 3590
rect 26730 3570 26735 3590
rect 26705 3540 26735 3570
rect 26705 3520 26710 3540
rect 26730 3520 26735 3540
rect 26705 3490 26735 3520
rect 26705 3470 26710 3490
rect 26730 3470 26735 3490
rect 26705 3440 26735 3470
rect 26705 3420 26710 3440
rect 26730 3420 26735 3440
rect 26705 3390 26735 3420
rect 26705 3370 26710 3390
rect 26730 3370 26735 3390
rect 26705 3340 26735 3370
rect 26705 3320 26710 3340
rect 26730 3320 26735 3340
rect 26705 3290 26735 3320
rect 26705 3270 26710 3290
rect 26730 3270 26735 3290
rect 26705 3240 26735 3270
rect 26705 3220 26710 3240
rect 26730 3220 26735 3240
rect 26705 3210 26735 3220
rect 26765 3590 26795 3600
rect 26765 3570 26770 3590
rect 26790 3570 26795 3590
rect 26765 3540 26795 3570
rect 26765 3520 26770 3540
rect 26790 3520 26795 3540
rect 26765 3490 26795 3520
rect 26765 3470 26770 3490
rect 26790 3470 26795 3490
rect 26765 3440 26795 3470
rect 26765 3420 26770 3440
rect 26790 3420 26795 3440
rect 26765 3390 26795 3420
rect 26765 3370 26770 3390
rect 26790 3370 26795 3390
rect 26765 3340 26795 3370
rect 26765 3320 26770 3340
rect 26790 3320 26795 3340
rect 26765 3290 26795 3320
rect 26765 3270 26770 3290
rect 26790 3270 26795 3290
rect 26765 3240 26795 3270
rect 26765 3220 26770 3240
rect 26790 3220 26795 3240
rect 26765 3210 26795 3220
rect 26825 3590 26855 3600
rect 26825 3570 26830 3590
rect 26850 3570 26855 3590
rect 26825 3540 26855 3570
rect 26825 3520 26830 3540
rect 26850 3520 26855 3540
rect 26825 3490 26855 3520
rect 26825 3470 26830 3490
rect 26850 3470 26855 3490
rect 26825 3440 26855 3470
rect 26825 3420 26830 3440
rect 26850 3420 26855 3440
rect 26825 3390 26855 3420
rect 26825 3370 26830 3390
rect 26850 3370 26855 3390
rect 26825 3340 26855 3370
rect 26825 3320 26830 3340
rect 26850 3320 26855 3340
rect 26825 3290 26855 3320
rect 26825 3270 26830 3290
rect 26850 3270 26855 3290
rect 26825 3240 26855 3270
rect 26825 3220 26830 3240
rect 26850 3220 26855 3240
rect 26825 3210 26855 3220
rect 26885 3590 26915 3600
rect 26885 3570 26890 3590
rect 26910 3570 26915 3590
rect 26885 3540 26915 3570
rect 26885 3520 26890 3540
rect 26910 3520 26915 3540
rect 26885 3490 26915 3520
rect 26885 3470 26890 3490
rect 26910 3470 26915 3490
rect 26885 3440 26915 3470
rect 26885 3420 26890 3440
rect 26910 3420 26915 3440
rect 26885 3390 26915 3420
rect 26885 3370 26890 3390
rect 26910 3370 26915 3390
rect 26885 3340 26915 3370
rect 26885 3320 26890 3340
rect 26910 3320 26915 3340
rect 26885 3290 26915 3320
rect 26885 3270 26890 3290
rect 26910 3270 26915 3290
rect 26885 3240 26915 3270
rect 26885 3220 26890 3240
rect 26910 3220 26915 3240
rect 26885 3210 26915 3220
rect 26945 3590 26975 3600
rect 26945 3570 26950 3590
rect 26970 3570 26975 3590
rect 26945 3540 26975 3570
rect 26945 3520 26950 3540
rect 26970 3520 26975 3540
rect 26945 3490 26975 3520
rect 26945 3470 26950 3490
rect 26970 3470 26975 3490
rect 26945 3440 26975 3470
rect 26945 3420 26950 3440
rect 26970 3420 26975 3440
rect 26945 3390 26975 3420
rect 26945 3370 26950 3390
rect 26970 3370 26975 3390
rect 26945 3340 26975 3370
rect 26945 3320 26950 3340
rect 26970 3320 26975 3340
rect 26945 3290 26975 3320
rect 26945 3270 26950 3290
rect 26970 3270 26975 3290
rect 26945 3240 26975 3270
rect 26945 3220 26950 3240
rect 26970 3220 26975 3240
rect 26945 3210 26975 3220
rect 27005 3590 27035 3600
rect 27005 3570 27010 3590
rect 27030 3570 27035 3590
rect 27005 3540 27035 3570
rect 27005 3520 27010 3540
rect 27030 3520 27035 3540
rect 27005 3490 27035 3520
rect 27005 3470 27010 3490
rect 27030 3470 27035 3490
rect 27005 3440 27035 3470
rect 27005 3420 27010 3440
rect 27030 3420 27035 3440
rect 27005 3390 27035 3420
rect 27005 3370 27010 3390
rect 27030 3370 27035 3390
rect 27005 3340 27035 3370
rect 27005 3320 27010 3340
rect 27030 3320 27035 3340
rect 27005 3290 27035 3320
rect 27005 3270 27010 3290
rect 27030 3270 27035 3290
rect 27005 3240 27035 3270
rect 27005 3220 27010 3240
rect 27030 3220 27035 3240
rect 27005 3210 27035 3220
rect 27065 3590 27095 3600
rect 27065 3570 27070 3590
rect 27090 3570 27095 3590
rect 27065 3540 27095 3570
rect 27065 3520 27070 3540
rect 27090 3520 27095 3540
rect 27065 3490 27095 3520
rect 27065 3470 27070 3490
rect 27090 3470 27095 3490
rect 27065 3440 27095 3470
rect 27065 3420 27070 3440
rect 27090 3420 27095 3440
rect 27065 3390 27095 3420
rect 27065 3370 27070 3390
rect 27090 3370 27095 3390
rect 27065 3340 27095 3370
rect 27065 3320 27070 3340
rect 27090 3320 27095 3340
rect 27065 3290 27095 3320
rect 27065 3270 27070 3290
rect 27090 3270 27095 3290
rect 27065 3240 27095 3270
rect 27065 3220 27070 3240
rect 27090 3220 27095 3240
rect 27065 3210 27095 3220
rect 27125 3590 27155 3600
rect 27125 3570 27130 3590
rect 27150 3570 27155 3590
rect 27125 3540 27155 3570
rect 27125 3520 27130 3540
rect 27150 3520 27155 3540
rect 27125 3490 27155 3520
rect 27125 3470 27130 3490
rect 27150 3470 27155 3490
rect 27125 3440 27155 3470
rect 27125 3420 27130 3440
rect 27150 3420 27155 3440
rect 27125 3390 27155 3420
rect 27125 3370 27130 3390
rect 27150 3370 27155 3390
rect 27125 3340 27155 3370
rect 27125 3320 27130 3340
rect 27150 3320 27155 3340
rect 27125 3290 27155 3320
rect 27125 3270 27130 3290
rect 27150 3270 27155 3290
rect 27125 3240 27155 3270
rect 27125 3220 27130 3240
rect 27150 3220 27155 3240
rect 27125 3210 27155 3220
rect 27185 3590 27215 3600
rect 27185 3570 27190 3590
rect 27210 3570 27215 3590
rect 27185 3540 27215 3570
rect 27185 3520 27190 3540
rect 27210 3520 27215 3540
rect 27185 3490 27215 3520
rect 27185 3470 27190 3490
rect 27210 3470 27215 3490
rect 27185 3440 27215 3470
rect 27185 3420 27190 3440
rect 27210 3420 27215 3440
rect 27185 3390 27215 3420
rect 27185 3370 27190 3390
rect 27210 3370 27215 3390
rect 27185 3340 27215 3370
rect 27185 3320 27190 3340
rect 27210 3320 27215 3340
rect 27185 3290 27215 3320
rect 27185 3270 27190 3290
rect 27210 3270 27215 3290
rect 27185 3240 27215 3270
rect 27185 3220 27190 3240
rect 27210 3220 27215 3240
rect 27185 3210 27215 3220
rect 27245 3590 27275 3600
rect 27245 3570 27250 3590
rect 27270 3570 27275 3590
rect 27245 3540 27275 3570
rect 27245 3520 27250 3540
rect 27270 3520 27275 3540
rect 27245 3490 27275 3520
rect 27245 3470 27250 3490
rect 27270 3470 27275 3490
rect 27245 3440 27275 3470
rect 27245 3420 27250 3440
rect 27270 3420 27275 3440
rect 27245 3390 27275 3420
rect 27245 3370 27250 3390
rect 27270 3370 27275 3390
rect 27245 3340 27275 3370
rect 27245 3320 27250 3340
rect 27270 3320 27275 3340
rect 27245 3290 27275 3320
rect 27245 3270 27250 3290
rect 27270 3270 27275 3290
rect 27245 3240 27275 3270
rect 27245 3220 27250 3240
rect 27270 3220 27275 3240
rect 27245 3210 27275 3220
rect 27305 3590 27335 3600
rect 27305 3570 27310 3590
rect 27330 3570 27335 3590
rect 27305 3540 27335 3570
rect 27305 3520 27310 3540
rect 27330 3520 27335 3540
rect 27305 3490 27335 3520
rect 27305 3470 27310 3490
rect 27330 3470 27335 3490
rect 27305 3440 27335 3470
rect 27305 3420 27310 3440
rect 27330 3420 27335 3440
rect 27305 3390 27335 3420
rect 27305 3370 27310 3390
rect 27330 3370 27335 3390
rect 27305 3340 27335 3370
rect 27305 3320 27310 3340
rect 27330 3320 27335 3340
rect 27305 3290 27335 3320
rect 27305 3270 27310 3290
rect 27330 3270 27335 3290
rect 27305 3240 27335 3270
rect 27305 3220 27310 3240
rect 27330 3220 27335 3240
rect 27305 3210 27335 3220
rect 27365 3590 27395 3600
rect 27365 3570 27370 3590
rect 27390 3570 27395 3590
rect 27365 3540 27395 3570
rect 27365 3520 27370 3540
rect 27390 3520 27395 3540
rect 27365 3490 27395 3520
rect 27365 3470 27370 3490
rect 27390 3470 27395 3490
rect 27365 3440 27395 3470
rect 27365 3420 27370 3440
rect 27390 3420 27395 3440
rect 27365 3390 27395 3420
rect 27365 3370 27370 3390
rect 27390 3370 27395 3390
rect 27365 3340 27395 3370
rect 27365 3320 27370 3340
rect 27390 3320 27395 3340
rect 27365 3290 27395 3320
rect 27365 3270 27370 3290
rect 27390 3270 27395 3290
rect 27365 3240 27395 3270
rect 27365 3220 27370 3240
rect 27390 3220 27395 3240
rect 27365 3210 27395 3220
rect 27425 3590 27455 3600
rect 27425 3570 27430 3590
rect 27450 3570 27455 3590
rect 27425 3540 27455 3570
rect 27425 3520 27430 3540
rect 27450 3520 27455 3540
rect 27425 3490 27455 3520
rect 27425 3470 27430 3490
rect 27450 3470 27455 3490
rect 27425 3440 27455 3470
rect 27425 3420 27430 3440
rect 27450 3420 27455 3440
rect 27425 3390 27455 3420
rect 27425 3370 27430 3390
rect 27450 3370 27455 3390
rect 27425 3340 27455 3370
rect 27425 3320 27430 3340
rect 27450 3320 27455 3340
rect 27425 3290 27455 3320
rect 27425 3270 27430 3290
rect 27450 3270 27455 3290
rect 27425 3240 27455 3270
rect 27425 3220 27430 3240
rect 27450 3220 27455 3240
rect 27425 3210 27455 3220
rect 27485 3590 27515 3600
rect 27485 3570 27490 3590
rect 27510 3570 27515 3590
rect 27485 3540 27515 3570
rect 27485 3520 27490 3540
rect 27510 3520 27515 3540
rect 27485 3490 27515 3520
rect 27485 3470 27490 3490
rect 27510 3470 27515 3490
rect 27485 3440 27515 3470
rect 27485 3420 27490 3440
rect 27510 3420 27515 3440
rect 27485 3390 27515 3420
rect 27485 3370 27490 3390
rect 27510 3370 27515 3390
rect 27485 3340 27515 3370
rect 27485 3320 27490 3340
rect 27510 3320 27515 3340
rect 27485 3290 27515 3320
rect 27485 3270 27490 3290
rect 27510 3270 27515 3290
rect 27485 3240 27515 3270
rect 27485 3220 27490 3240
rect 27510 3220 27515 3240
rect 27485 3210 27515 3220
rect 27545 3590 27575 3600
rect 27545 3570 27550 3590
rect 27570 3570 27575 3590
rect 27545 3540 27575 3570
rect 27545 3520 27550 3540
rect 27570 3520 27575 3540
rect 27545 3490 27575 3520
rect 27545 3470 27550 3490
rect 27570 3470 27575 3490
rect 27545 3440 27575 3470
rect 27545 3420 27550 3440
rect 27570 3420 27575 3440
rect 27545 3390 27575 3420
rect 27545 3370 27550 3390
rect 27570 3370 27575 3390
rect 27545 3340 27575 3370
rect 27545 3320 27550 3340
rect 27570 3320 27575 3340
rect 27545 3290 27575 3320
rect 27545 3270 27550 3290
rect 27570 3270 27575 3290
rect 27545 3240 27575 3270
rect 27545 3220 27550 3240
rect 27570 3220 27575 3240
rect 27545 3210 27575 3220
rect 27610 3445 27630 3680
rect 26290 3190 26310 3210
rect 26410 3190 26430 3210
rect 26530 3190 26550 3210
rect 26650 3190 26670 3210
rect 26770 3190 26790 3210
rect 26890 3190 26910 3210
rect 27010 3190 27030 3210
rect 27130 3190 27150 3210
rect 27250 3190 27270 3210
rect 27370 3190 27390 3210
rect 27490 3190 27510 3210
rect 26280 3180 26320 3190
rect 26280 3160 26290 3180
rect 26310 3160 26320 3180
rect 26280 3150 26320 3160
rect 26400 3180 26440 3190
rect 26400 3160 26410 3180
rect 26430 3160 26440 3180
rect 26400 3150 26440 3160
rect 26520 3180 26560 3190
rect 26520 3160 26530 3180
rect 26550 3160 26560 3180
rect 26520 3150 26560 3160
rect 26640 3180 26680 3190
rect 26640 3160 26650 3180
rect 26670 3160 26680 3180
rect 26640 3150 26680 3160
rect 26760 3180 26800 3190
rect 26760 3160 26770 3180
rect 26790 3160 26800 3180
rect 26760 3150 26800 3160
rect 26823 3180 26857 3190
rect 26823 3160 26831 3180
rect 26849 3160 26857 3180
rect 26823 3150 26857 3160
rect 26880 3180 26920 3190
rect 26880 3160 26890 3180
rect 26910 3160 26920 3180
rect 26880 3150 26920 3160
rect 27000 3180 27040 3190
rect 27000 3160 27010 3180
rect 27030 3160 27040 3180
rect 27000 3150 27040 3160
rect 27120 3180 27160 3190
rect 27120 3160 27130 3180
rect 27150 3160 27160 3180
rect 27120 3150 27160 3160
rect 27240 3180 27280 3190
rect 27240 3160 27250 3180
rect 27270 3160 27280 3180
rect 27240 3150 27280 3160
rect 27360 3180 27400 3190
rect 27360 3160 27370 3180
rect 27390 3160 27400 3180
rect 27360 3150 27400 3160
rect 27480 3180 27520 3190
rect 27480 3160 27490 3180
rect 27510 3160 27520 3180
rect 27480 3150 27520 3160
rect 27610 3130 27630 3365
rect 26170 3110 26860 3130
rect 26940 3110 27630 3130
rect 28095 3410 28115 3740
rect 28200 3710 28240 3720
rect 28200 3690 28210 3710
rect 28230 3690 28240 3710
rect 28200 3680 28240 3690
rect 28310 3710 28350 3720
rect 28310 3690 28320 3710
rect 28340 3690 28350 3710
rect 28310 3680 28350 3690
rect 28420 3710 28460 3720
rect 28420 3690 28430 3710
rect 28450 3690 28460 3710
rect 28420 3680 28460 3690
rect 28530 3710 28570 3720
rect 28530 3690 28540 3710
rect 28560 3690 28570 3710
rect 28530 3680 28570 3690
rect 28640 3710 28680 3720
rect 28640 3690 28650 3710
rect 28670 3690 28680 3710
rect 28640 3680 28680 3690
rect 28750 3710 28790 3720
rect 28750 3690 28760 3710
rect 28780 3690 28790 3710
rect 28750 3680 28790 3690
rect 28210 3660 28230 3680
rect 28320 3660 28340 3680
rect 28430 3660 28450 3680
rect 28540 3660 28560 3680
rect 28650 3660 28670 3680
rect 28760 3660 28780 3680
rect 25670 3070 25740 3100
rect 25670 3050 25675 3070
rect 25695 3050 25715 3070
rect 25735 3050 25740 3070
rect 25670 3020 25740 3050
rect 25670 3000 25675 3020
rect 25695 3000 25715 3020
rect 25735 3000 25740 3020
rect 25670 2990 25740 3000
rect 28095 2990 28115 3315
rect 28150 3650 28180 3660
rect 28150 3630 28155 3650
rect 28175 3630 28180 3650
rect 28150 3600 28180 3630
rect 28150 3580 28155 3600
rect 28175 3580 28180 3600
rect 28150 3550 28180 3580
rect 28150 3530 28155 3550
rect 28175 3530 28180 3550
rect 28150 3500 28180 3530
rect 28150 3480 28155 3500
rect 28175 3480 28180 3500
rect 28150 3450 28180 3480
rect 28150 3430 28155 3450
rect 28175 3430 28180 3450
rect 28150 3400 28180 3430
rect 28150 3380 28155 3400
rect 28175 3380 28180 3400
rect 28150 3350 28180 3380
rect 28150 3330 28155 3350
rect 28175 3330 28180 3350
rect 28150 3300 28180 3330
rect 28150 3280 28155 3300
rect 28175 3280 28180 3300
rect 28150 3250 28180 3280
rect 28150 3230 28155 3250
rect 28175 3230 28180 3250
rect 28150 3200 28180 3230
rect 28150 3180 28155 3200
rect 28175 3180 28180 3200
rect 28150 3150 28180 3180
rect 28150 3130 28155 3150
rect 28175 3130 28180 3150
rect 28150 3100 28180 3130
rect 28150 3080 28155 3100
rect 28175 3080 28180 3100
rect 28150 3070 28180 3080
rect 28205 3650 28235 3660
rect 28205 3630 28210 3650
rect 28230 3630 28235 3650
rect 28205 3600 28235 3630
rect 28205 3580 28210 3600
rect 28230 3580 28235 3600
rect 28205 3550 28235 3580
rect 28205 3530 28210 3550
rect 28230 3530 28235 3550
rect 28205 3500 28235 3530
rect 28205 3480 28210 3500
rect 28230 3480 28235 3500
rect 28205 3450 28235 3480
rect 28205 3430 28210 3450
rect 28230 3430 28235 3450
rect 28205 3400 28235 3430
rect 28205 3380 28210 3400
rect 28230 3380 28235 3400
rect 28205 3350 28235 3380
rect 28205 3330 28210 3350
rect 28230 3330 28235 3350
rect 28205 3300 28235 3330
rect 28205 3280 28210 3300
rect 28230 3280 28235 3300
rect 28205 3250 28235 3280
rect 28205 3230 28210 3250
rect 28230 3230 28235 3250
rect 28205 3200 28235 3230
rect 28205 3180 28210 3200
rect 28230 3180 28235 3200
rect 28205 3150 28235 3180
rect 28205 3130 28210 3150
rect 28230 3130 28235 3150
rect 28205 3100 28235 3130
rect 28205 3080 28210 3100
rect 28230 3080 28235 3100
rect 28205 3070 28235 3080
rect 28260 3650 28290 3660
rect 28260 3630 28265 3650
rect 28285 3630 28290 3650
rect 28260 3600 28290 3630
rect 28260 3580 28265 3600
rect 28285 3580 28290 3600
rect 28260 3550 28290 3580
rect 28260 3530 28265 3550
rect 28285 3530 28290 3550
rect 28260 3500 28290 3530
rect 28260 3480 28265 3500
rect 28285 3480 28290 3500
rect 28260 3450 28290 3480
rect 28260 3430 28265 3450
rect 28285 3430 28290 3450
rect 28260 3400 28290 3430
rect 28260 3380 28265 3400
rect 28285 3380 28290 3400
rect 28260 3350 28290 3380
rect 28260 3330 28265 3350
rect 28285 3330 28290 3350
rect 28260 3300 28290 3330
rect 28260 3280 28265 3300
rect 28285 3280 28290 3300
rect 28260 3250 28290 3280
rect 28260 3230 28265 3250
rect 28285 3230 28290 3250
rect 28260 3200 28290 3230
rect 28260 3180 28265 3200
rect 28285 3180 28290 3200
rect 28260 3150 28290 3180
rect 28260 3130 28265 3150
rect 28285 3130 28290 3150
rect 28260 3100 28290 3130
rect 28260 3080 28265 3100
rect 28285 3080 28290 3100
rect 28260 3070 28290 3080
rect 28315 3650 28345 3660
rect 28315 3630 28320 3650
rect 28340 3630 28345 3650
rect 28315 3600 28345 3630
rect 28315 3580 28320 3600
rect 28340 3580 28345 3600
rect 28315 3550 28345 3580
rect 28315 3530 28320 3550
rect 28340 3530 28345 3550
rect 28315 3500 28345 3530
rect 28315 3480 28320 3500
rect 28340 3480 28345 3500
rect 28315 3450 28345 3480
rect 28315 3430 28320 3450
rect 28340 3430 28345 3450
rect 28315 3400 28345 3430
rect 28315 3380 28320 3400
rect 28340 3380 28345 3400
rect 28315 3350 28345 3380
rect 28315 3330 28320 3350
rect 28340 3330 28345 3350
rect 28315 3300 28345 3330
rect 28315 3280 28320 3300
rect 28340 3280 28345 3300
rect 28315 3250 28345 3280
rect 28315 3230 28320 3250
rect 28340 3230 28345 3250
rect 28315 3200 28345 3230
rect 28315 3180 28320 3200
rect 28340 3180 28345 3200
rect 28315 3150 28345 3180
rect 28315 3130 28320 3150
rect 28340 3130 28345 3150
rect 28315 3100 28345 3130
rect 28315 3080 28320 3100
rect 28340 3080 28345 3100
rect 28315 3070 28345 3080
rect 28370 3650 28400 3660
rect 28370 3630 28375 3650
rect 28395 3630 28400 3650
rect 28370 3600 28400 3630
rect 28370 3580 28375 3600
rect 28395 3580 28400 3600
rect 28370 3550 28400 3580
rect 28370 3530 28375 3550
rect 28395 3530 28400 3550
rect 28370 3500 28400 3530
rect 28370 3480 28375 3500
rect 28395 3480 28400 3500
rect 28370 3450 28400 3480
rect 28370 3430 28375 3450
rect 28395 3430 28400 3450
rect 28370 3400 28400 3430
rect 28370 3380 28375 3400
rect 28395 3380 28400 3400
rect 28370 3350 28400 3380
rect 28370 3330 28375 3350
rect 28395 3330 28400 3350
rect 28370 3300 28400 3330
rect 28370 3280 28375 3300
rect 28395 3280 28400 3300
rect 28370 3250 28400 3280
rect 28370 3230 28375 3250
rect 28395 3230 28400 3250
rect 28370 3200 28400 3230
rect 28370 3180 28375 3200
rect 28395 3180 28400 3200
rect 28370 3150 28400 3180
rect 28370 3130 28375 3150
rect 28395 3130 28400 3150
rect 28370 3100 28400 3130
rect 28370 3080 28375 3100
rect 28395 3080 28400 3100
rect 28370 3070 28400 3080
rect 28425 3650 28455 3660
rect 28425 3630 28430 3650
rect 28450 3630 28455 3650
rect 28425 3600 28455 3630
rect 28425 3580 28430 3600
rect 28450 3580 28455 3600
rect 28425 3550 28455 3580
rect 28425 3530 28430 3550
rect 28450 3530 28455 3550
rect 28425 3500 28455 3530
rect 28425 3480 28430 3500
rect 28450 3480 28455 3500
rect 28425 3450 28455 3480
rect 28425 3430 28430 3450
rect 28450 3430 28455 3450
rect 28425 3400 28455 3430
rect 28425 3380 28430 3400
rect 28450 3380 28455 3400
rect 28425 3350 28455 3380
rect 28425 3330 28430 3350
rect 28450 3330 28455 3350
rect 28425 3300 28455 3330
rect 28425 3280 28430 3300
rect 28450 3280 28455 3300
rect 28425 3250 28455 3280
rect 28425 3230 28430 3250
rect 28450 3230 28455 3250
rect 28425 3200 28455 3230
rect 28425 3180 28430 3200
rect 28450 3180 28455 3200
rect 28425 3150 28455 3180
rect 28425 3130 28430 3150
rect 28450 3130 28455 3150
rect 28425 3100 28455 3130
rect 28425 3080 28430 3100
rect 28450 3080 28455 3100
rect 28425 3070 28455 3080
rect 28480 3650 28510 3660
rect 28480 3630 28485 3650
rect 28505 3630 28510 3650
rect 28480 3600 28510 3630
rect 28480 3580 28485 3600
rect 28505 3580 28510 3600
rect 28480 3550 28510 3580
rect 28480 3530 28485 3550
rect 28505 3530 28510 3550
rect 28480 3500 28510 3530
rect 28480 3480 28485 3500
rect 28505 3480 28510 3500
rect 28480 3450 28510 3480
rect 28480 3430 28485 3450
rect 28505 3430 28510 3450
rect 28480 3400 28510 3430
rect 28480 3380 28485 3400
rect 28505 3380 28510 3400
rect 28480 3350 28510 3380
rect 28480 3330 28485 3350
rect 28505 3330 28510 3350
rect 28480 3300 28510 3330
rect 28480 3280 28485 3300
rect 28505 3280 28510 3300
rect 28480 3250 28510 3280
rect 28480 3230 28485 3250
rect 28505 3230 28510 3250
rect 28480 3200 28510 3230
rect 28480 3180 28485 3200
rect 28505 3180 28510 3200
rect 28480 3150 28510 3180
rect 28480 3130 28485 3150
rect 28505 3130 28510 3150
rect 28480 3100 28510 3130
rect 28480 3080 28485 3100
rect 28505 3080 28510 3100
rect 28480 3070 28510 3080
rect 28535 3650 28565 3660
rect 28535 3630 28540 3650
rect 28560 3630 28565 3650
rect 28535 3600 28565 3630
rect 28535 3580 28540 3600
rect 28560 3580 28565 3600
rect 28535 3550 28565 3580
rect 28535 3530 28540 3550
rect 28560 3530 28565 3550
rect 28535 3500 28565 3530
rect 28535 3480 28540 3500
rect 28560 3480 28565 3500
rect 28535 3450 28565 3480
rect 28535 3430 28540 3450
rect 28560 3430 28565 3450
rect 28535 3400 28565 3430
rect 28535 3380 28540 3400
rect 28560 3380 28565 3400
rect 28535 3350 28565 3380
rect 28535 3330 28540 3350
rect 28560 3330 28565 3350
rect 28535 3300 28565 3330
rect 28535 3280 28540 3300
rect 28560 3280 28565 3300
rect 28535 3250 28565 3280
rect 28535 3230 28540 3250
rect 28560 3230 28565 3250
rect 28535 3200 28565 3230
rect 28535 3180 28540 3200
rect 28560 3180 28565 3200
rect 28535 3150 28565 3180
rect 28535 3130 28540 3150
rect 28560 3130 28565 3150
rect 28535 3100 28565 3130
rect 28535 3080 28540 3100
rect 28560 3080 28565 3100
rect 28535 3070 28565 3080
rect 28590 3650 28620 3660
rect 28590 3630 28595 3650
rect 28615 3630 28620 3650
rect 28590 3600 28620 3630
rect 28590 3580 28595 3600
rect 28615 3580 28620 3600
rect 28590 3550 28620 3580
rect 28590 3530 28595 3550
rect 28615 3530 28620 3550
rect 28590 3500 28620 3530
rect 28590 3480 28595 3500
rect 28615 3480 28620 3500
rect 28590 3450 28620 3480
rect 28590 3430 28595 3450
rect 28615 3430 28620 3450
rect 28590 3400 28620 3430
rect 28590 3380 28595 3400
rect 28615 3380 28620 3400
rect 28590 3350 28620 3380
rect 28590 3330 28595 3350
rect 28615 3330 28620 3350
rect 28590 3300 28620 3330
rect 28590 3280 28595 3300
rect 28615 3280 28620 3300
rect 28590 3250 28620 3280
rect 28590 3230 28595 3250
rect 28615 3230 28620 3250
rect 28590 3200 28620 3230
rect 28590 3180 28595 3200
rect 28615 3180 28620 3200
rect 28590 3150 28620 3180
rect 28590 3130 28595 3150
rect 28615 3130 28620 3150
rect 28590 3100 28620 3130
rect 28590 3080 28595 3100
rect 28615 3080 28620 3100
rect 28590 3070 28620 3080
rect 28645 3650 28675 3660
rect 28645 3630 28650 3650
rect 28670 3630 28675 3650
rect 28645 3600 28675 3630
rect 28645 3580 28650 3600
rect 28670 3580 28675 3600
rect 28645 3550 28675 3580
rect 28645 3530 28650 3550
rect 28670 3530 28675 3550
rect 28645 3500 28675 3530
rect 28645 3480 28650 3500
rect 28670 3480 28675 3500
rect 28645 3450 28675 3480
rect 28645 3430 28650 3450
rect 28670 3430 28675 3450
rect 28645 3400 28675 3430
rect 28645 3380 28650 3400
rect 28670 3380 28675 3400
rect 28645 3350 28675 3380
rect 28645 3330 28650 3350
rect 28670 3330 28675 3350
rect 28645 3300 28675 3330
rect 28645 3280 28650 3300
rect 28670 3280 28675 3300
rect 28645 3250 28675 3280
rect 28645 3230 28650 3250
rect 28670 3230 28675 3250
rect 28645 3200 28675 3230
rect 28645 3180 28650 3200
rect 28670 3180 28675 3200
rect 28645 3150 28675 3180
rect 28645 3130 28650 3150
rect 28670 3130 28675 3150
rect 28645 3100 28675 3130
rect 28645 3080 28650 3100
rect 28670 3080 28675 3100
rect 28645 3070 28675 3080
rect 28700 3650 28730 3660
rect 28700 3630 28705 3650
rect 28725 3630 28730 3650
rect 28700 3600 28730 3630
rect 28700 3580 28705 3600
rect 28725 3580 28730 3600
rect 28700 3550 28730 3580
rect 28700 3530 28705 3550
rect 28725 3530 28730 3550
rect 28700 3500 28730 3530
rect 28700 3480 28705 3500
rect 28725 3480 28730 3500
rect 28700 3450 28730 3480
rect 28700 3430 28705 3450
rect 28725 3430 28730 3450
rect 28700 3400 28730 3430
rect 28700 3380 28705 3400
rect 28725 3380 28730 3400
rect 28700 3350 28730 3380
rect 28700 3330 28705 3350
rect 28725 3330 28730 3350
rect 28700 3300 28730 3330
rect 28700 3280 28705 3300
rect 28725 3280 28730 3300
rect 28700 3250 28730 3280
rect 28700 3230 28705 3250
rect 28725 3230 28730 3250
rect 28700 3200 28730 3230
rect 28700 3180 28705 3200
rect 28725 3180 28730 3200
rect 28700 3150 28730 3180
rect 28700 3130 28705 3150
rect 28725 3130 28730 3150
rect 28700 3100 28730 3130
rect 28700 3080 28705 3100
rect 28725 3080 28730 3100
rect 28700 3070 28730 3080
rect 28755 3650 28785 3660
rect 28755 3630 28760 3650
rect 28780 3630 28785 3650
rect 28755 3600 28785 3630
rect 28755 3580 28760 3600
rect 28780 3580 28785 3600
rect 28755 3550 28785 3580
rect 28755 3530 28760 3550
rect 28780 3530 28785 3550
rect 28755 3500 28785 3530
rect 28755 3480 28760 3500
rect 28780 3480 28785 3500
rect 28755 3450 28785 3480
rect 28755 3430 28760 3450
rect 28780 3430 28785 3450
rect 28755 3400 28785 3430
rect 28755 3380 28760 3400
rect 28780 3380 28785 3400
rect 28755 3350 28785 3380
rect 28755 3330 28760 3350
rect 28780 3330 28785 3350
rect 28755 3300 28785 3330
rect 28755 3280 28760 3300
rect 28780 3280 28785 3300
rect 28755 3250 28785 3280
rect 28755 3230 28760 3250
rect 28780 3230 28785 3250
rect 28755 3200 28785 3230
rect 28755 3180 28760 3200
rect 28780 3180 28785 3200
rect 28755 3150 28785 3180
rect 28755 3130 28760 3150
rect 28780 3130 28785 3150
rect 28755 3100 28785 3130
rect 28755 3080 28760 3100
rect 28780 3080 28785 3100
rect 28755 3070 28785 3080
rect 28810 3650 28840 3660
rect 28810 3630 28815 3650
rect 28835 3630 28840 3650
rect 28810 3600 28840 3630
rect 28810 3580 28815 3600
rect 28835 3580 28840 3600
rect 28810 3550 28840 3580
rect 28810 3530 28815 3550
rect 28835 3530 28840 3550
rect 28810 3500 28840 3530
rect 28810 3480 28815 3500
rect 28835 3480 28840 3500
rect 28810 3450 28840 3480
rect 28810 3430 28815 3450
rect 28835 3430 28840 3450
rect 28810 3400 28840 3430
rect 28810 3380 28815 3400
rect 28835 3380 28840 3400
rect 28810 3350 28840 3380
rect 28810 3330 28815 3350
rect 28835 3330 28840 3350
rect 28810 3300 28840 3330
rect 28810 3280 28815 3300
rect 28835 3280 28840 3300
rect 28810 3250 28840 3280
rect 28810 3230 28815 3250
rect 28835 3230 28840 3250
rect 28810 3200 28840 3230
rect 28810 3180 28815 3200
rect 28835 3180 28840 3200
rect 28810 3150 28840 3180
rect 28810 3130 28815 3150
rect 28835 3130 28840 3150
rect 28810 3100 28840 3130
rect 28810 3080 28815 3100
rect 28835 3080 28840 3100
rect 28810 3070 28840 3080
rect 28875 3410 28895 3740
rect 28265 3050 28285 3070
rect 28375 3050 28395 3070
rect 28485 3050 28505 3070
rect 28595 3050 28615 3070
rect 28705 3050 28725 3070
rect 28255 3040 28295 3050
rect 28255 3020 28265 3040
rect 28285 3020 28295 3040
rect 28255 3010 28295 3020
rect 28313 3040 28347 3050
rect 28313 3020 28321 3040
rect 28339 3020 28347 3040
rect 28313 3010 28347 3020
rect 28365 3040 28405 3050
rect 28365 3020 28375 3040
rect 28395 3020 28405 3040
rect 28365 3010 28405 3020
rect 28475 3040 28515 3050
rect 28475 3020 28485 3040
rect 28505 3020 28515 3040
rect 28475 3010 28515 3020
rect 28585 3040 28625 3050
rect 28585 3020 28595 3040
rect 28615 3020 28625 3040
rect 28585 3010 28625 3020
rect 28695 3040 28735 3050
rect 28695 3020 28705 3040
rect 28725 3020 28735 3040
rect 28695 3010 28735 3020
rect 28875 2990 28895 3315
rect 24975 2970 24995 2990
rect 25125 2970 25145 2990
rect 25235 2970 25255 2990
rect 25345 2970 25365 2990
rect 25455 2970 25475 2990
rect 25565 2970 25585 2990
rect 25715 2970 25735 2990
rect 28095 2970 28455 2990
rect 28535 2970 28895 2990
rect 29035 3680 29315 3700
rect 29035 3375 29055 3680
rect 29105 3620 29246 3660
rect 29035 2980 29055 3280
rect 29295 3375 29315 3680
rect 29105 3000 29246 3040
rect 29295 2980 29315 3280
rect 24554 2900 24695 2940
rect 24965 2960 25005 2970
rect 24965 2940 24975 2960
rect 24995 2940 25005 2960
rect 24965 2930 25005 2940
rect 25115 2960 25155 2970
rect 25115 2940 25125 2960
rect 25145 2940 25155 2960
rect 25115 2930 25155 2940
rect 25225 2960 25265 2970
rect 25225 2940 25235 2960
rect 25255 2940 25265 2960
rect 25225 2930 25265 2940
rect 25335 2960 25375 2970
rect 25335 2940 25345 2960
rect 25365 2940 25375 2960
rect 25335 2930 25375 2940
rect 25445 2960 25485 2970
rect 25445 2940 25455 2960
rect 25475 2940 25485 2960
rect 25445 2930 25485 2940
rect 25503 2960 25537 2970
rect 25503 2940 25511 2960
rect 25529 2940 25537 2960
rect 25503 2930 25537 2940
rect 25555 2960 25595 2970
rect 25555 2940 25565 2960
rect 25585 2940 25595 2960
rect 25555 2930 25595 2940
rect 25705 2960 25745 2970
rect 29035 2960 29135 2980
rect 29215 2960 29315 2980
rect 25705 2940 25715 2960
rect 25735 2940 25745 2960
rect 25705 2930 25745 2940
rect 26985 2920 27375 2940
rect 27455 2920 27845 2940
rect 4980 2865 5050 2895
rect 4980 2845 4985 2865
rect 5005 2845 5025 2865
rect 5045 2845 5050 2865
rect 15975 2890 16015 2900
rect 15975 2870 15985 2890
rect 16005 2870 16015 2890
rect 15975 2860 16015 2870
rect 16135 2890 16175 2900
rect 16135 2870 16145 2890
rect 16165 2870 16175 2890
rect 16135 2860 16175 2870
rect 16255 2890 16295 2900
rect 16255 2870 16265 2890
rect 16285 2870 16295 2890
rect 16255 2860 16295 2870
rect 16375 2890 16415 2900
rect 16375 2870 16385 2890
rect 16405 2870 16415 2890
rect 16375 2860 16415 2870
rect 16495 2890 16535 2900
rect 16495 2870 16505 2890
rect 16525 2870 16535 2890
rect 16495 2860 16535 2870
rect 16615 2890 16655 2900
rect 16615 2870 16625 2890
rect 16645 2870 16655 2890
rect 16615 2860 16655 2870
rect 16775 2890 16815 2900
rect 16775 2870 16785 2890
rect 16805 2870 16815 2890
rect 16775 2860 16815 2870
rect 16985 2890 17025 2900
rect 16985 2870 16995 2890
rect 17015 2870 17025 2890
rect 16985 2860 17025 2870
rect 17145 2890 17185 2900
rect 17145 2870 17155 2890
rect 17175 2870 17185 2890
rect 17145 2860 17185 2870
rect 17265 2890 17305 2900
rect 17265 2870 17275 2890
rect 17295 2870 17305 2890
rect 17265 2860 17305 2870
rect 17385 2890 17425 2900
rect 17385 2870 17395 2890
rect 17415 2870 17425 2890
rect 17385 2860 17425 2870
rect 17505 2890 17545 2900
rect 17505 2870 17515 2890
rect 17535 2870 17545 2890
rect 17505 2860 17545 2870
rect 17625 2890 17665 2900
rect 17625 2870 17635 2890
rect 17655 2870 17665 2890
rect 17625 2860 17665 2870
rect 17785 2890 17825 2900
rect 17785 2870 17795 2890
rect 17815 2870 17825 2890
rect 17785 2860 17825 2870
rect 25975 2890 26015 2900
rect 25975 2870 25985 2890
rect 26005 2870 26015 2890
rect 25975 2860 26015 2870
rect 26135 2890 26175 2900
rect 26135 2870 26145 2890
rect 26165 2870 26175 2890
rect 26135 2860 26175 2870
rect 26255 2890 26295 2900
rect 26255 2870 26265 2890
rect 26285 2870 26295 2890
rect 26255 2860 26295 2870
rect 26375 2890 26415 2900
rect 26375 2870 26385 2890
rect 26405 2870 26415 2890
rect 26375 2860 26415 2870
rect 26495 2890 26535 2900
rect 26495 2870 26505 2890
rect 26525 2870 26535 2890
rect 26495 2860 26535 2870
rect 26615 2890 26655 2900
rect 26615 2870 26625 2890
rect 26645 2870 26655 2890
rect 26615 2860 26655 2870
rect 26775 2890 26815 2900
rect 26775 2870 26785 2890
rect 26805 2870 26815 2890
rect 26775 2860 26815 2870
rect 4980 2835 5050 2845
rect 15985 2840 16005 2860
rect 16145 2840 16165 2860
rect 16265 2840 16285 2860
rect 16385 2840 16405 2860
rect 16505 2840 16525 2860
rect 16625 2840 16645 2860
rect 16785 2840 16805 2860
rect 16995 2840 17015 2860
rect 17155 2840 17175 2860
rect 17275 2840 17295 2860
rect 17395 2840 17415 2860
rect 17515 2840 17535 2860
rect 17635 2840 17655 2860
rect 17795 2840 17815 2860
rect 25985 2840 26005 2860
rect 26145 2840 26165 2860
rect 26265 2840 26285 2860
rect 26385 2840 26405 2860
rect 26505 2840 26525 2860
rect 26625 2840 26645 2860
rect 26785 2840 26805 2860
rect 3005 2815 3025 2835
rect 3185 2815 3205 2835
rect 3365 2815 3385 2835
rect 3545 2815 3565 2835
rect 3725 2815 3745 2835
rect 3905 2815 3925 2835
rect 4085 2815 4105 2835
rect 4265 2815 4285 2835
rect 4445 2815 4465 2835
rect 4625 2815 4645 2835
rect 4805 2815 4825 2835
rect 4985 2815 5005 2835
rect 15980 2830 16050 2840
rect 2995 2805 3035 2815
rect -10 2765 20 2795
rect 51 2790 96 2795
rect 51 2765 61 2790
rect 86 2765 96 2790
rect 51 2760 96 2765
rect 724 2790 769 2795
rect 724 2765 734 2790
rect 759 2765 769 2790
rect 724 2760 769 2765
rect 2620 2755 2660 2795
rect 2995 2785 3005 2805
rect 3025 2785 3035 2805
rect 2995 2775 3035 2785
rect 3175 2805 3215 2815
rect 3175 2785 3185 2805
rect 3205 2785 3215 2805
rect 3175 2775 3215 2785
rect 3355 2805 3395 2815
rect 3355 2785 3365 2805
rect 3385 2785 3395 2805
rect 3355 2775 3395 2785
rect 3535 2805 3575 2815
rect 3535 2785 3545 2805
rect 3565 2785 3575 2805
rect 3535 2775 3575 2785
rect 3715 2805 3755 2815
rect 3715 2785 3725 2805
rect 3745 2785 3755 2805
rect 3715 2775 3755 2785
rect 3895 2805 3935 2815
rect 3895 2785 3905 2805
rect 3925 2785 3935 2805
rect 3895 2775 3935 2785
rect 4075 2805 4115 2815
rect 4075 2785 4085 2805
rect 4105 2785 4115 2805
rect 4075 2775 4115 2785
rect 4255 2805 4295 2815
rect 4255 2785 4265 2805
rect 4285 2785 4295 2805
rect 4255 2775 4295 2785
rect 4435 2805 4475 2815
rect 4435 2785 4445 2805
rect 4465 2785 4475 2805
rect 4435 2775 4475 2785
rect 4615 2805 4655 2815
rect 4615 2785 4625 2805
rect 4645 2785 4655 2805
rect 4615 2775 4655 2785
rect 4795 2805 4835 2815
rect 4795 2785 4805 2805
rect 4825 2785 4835 2805
rect 4795 2775 4835 2785
rect 4975 2805 5015 2815
rect 4975 2785 4985 2805
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 15980 2810 15985 2830
rect 16005 2810 16025 2830
rect 16045 2810 16050 2830
rect 15980 2780 16050 2810
rect 15980 2760 15985 2780
rect 16005 2760 16025 2780
rect 16045 2760 16050 2780
rect 1266 2715 1296 2745
rect 2150 2710 2190 2750
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2725 3215 2745
rect 3175 2715 3215 2725
rect 3355 2745 3395 2755
rect 3355 2725 3365 2745
rect 3385 2725 3395 2745
rect 3355 2715 3395 2725
rect 3535 2745 3575 2755
rect 3535 2725 3545 2745
rect 3565 2725 3575 2745
rect 3535 2715 3575 2725
rect 3715 2745 3755 2755
rect 3715 2725 3725 2745
rect 3745 2725 3755 2745
rect 3715 2715 3755 2725
rect 3895 2745 3935 2755
rect 3895 2725 3905 2745
rect 3925 2725 3935 2745
rect 3895 2715 3935 2725
rect 4075 2745 4115 2755
rect 4075 2725 4085 2745
rect 4105 2725 4115 2745
rect 4075 2715 4115 2725
rect 4255 2745 4295 2755
rect 4255 2725 4265 2745
rect 4285 2725 4295 2745
rect 4255 2715 4295 2725
rect 4435 2745 4475 2755
rect 4435 2725 4445 2745
rect 4465 2725 4475 2745
rect 4435 2715 4475 2725
rect 4615 2745 4655 2755
rect 4615 2725 4625 2745
rect 4645 2725 4655 2745
rect 4615 2715 4655 2725
rect 4795 2745 4835 2755
rect 4795 2725 4805 2745
rect 4825 2725 4835 2745
rect 4795 2715 4835 2725
rect 15980 2730 16050 2760
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3185 2695 3205 2715
rect 3365 2695 3385 2715
rect 3545 2695 3565 2715
rect 3725 2695 3745 2715
rect 3905 2695 3925 2715
rect 4085 2695 4105 2715
rect 4265 2695 4285 2715
rect 4445 2695 4465 2715
rect 4625 2695 4645 2715
rect 4805 2695 4825 2715
rect 15980 2710 15985 2730
rect 16005 2710 16025 2730
rect 16045 2710 16050 2730
rect 15060 2700 15100 2710
rect 3140 2685 3210 2695
rect 3140 2665 3145 2685
rect 3165 2665 3185 2685
rect 3205 2665 3210 2685
rect 3140 2635 3210 2665
rect 3140 2615 3145 2635
rect 3165 2615 3185 2635
rect 3205 2615 3210 2635
rect 3140 2585 3210 2615
rect 3140 2565 3145 2585
rect 3165 2565 3185 2585
rect 3205 2565 3210 2585
rect 3140 2535 3210 2565
rect 3140 2515 3145 2535
rect 3165 2515 3185 2535
rect 3205 2515 3210 2535
rect 3140 2485 3210 2515
rect 3140 2465 3145 2485
rect 3165 2465 3185 2485
rect 3205 2465 3210 2485
rect 3140 2435 3210 2465
rect 3140 2415 3145 2435
rect 3165 2415 3185 2435
rect 3205 2415 3210 2435
rect 3140 2405 3210 2415
rect 3270 2685 3300 2695
rect 3270 2665 3275 2685
rect 3295 2665 3300 2685
rect 3270 2635 3300 2665
rect 3270 2615 3275 2635
rect 3295 2615 3300 2635
rect 3270 2585 3300 2615
rect 3270 2565 3275 2585
rect 3295 2565 3300 2585
rect 3270 2535 3300 2565
rect 3270 2515 3275 2535
rect 3295 2515 3300 2535
rect 3270 2485 3300 2515
rect 3270 2465 3275 2485
rect 3295 2465 3300 2485
rect 3270 2435 3300 2465
rect 3270 2415 3275 2435
rect 3295 2415 3300 2435
rect 3270 2405 3300 2415
rect 3360 2685 3390 2695
rect 3360 2665 3365 2685
rect 3385 2665 3390 2685
rect 3360 2635 3390 2665
rect 3360 2615 3365 2635
rect 3385 2615 3390 2635
rect 3360 2585 3390 2615
rect 3360 2565 3365 2585
rect 3385 2565 3390 2585
rect 3360 2535 3390 2565
rect 3360 2515 3365 2535
rect 3385 2515 3390 2535
rect 3360 2485 3390 2515
rect 3360 2465 3365 2485
rect 3385 2465 3390 2485
rect 3360 2435 3390 2465
rect 3360 2415 3365 2435
rect 3385 2415 3390 2435
rect 3360 2405 3390 2415
rect 3450 2685 3480 2695
rect 3450 2665 3455 2685
rect 3475 2665 3480 2685
rect 3450 2635 3480 2665
rect 3450 2615 3455 2635
rect 3475 2615 3480 2635
rect 3450 2585 3480 2615
rect 3450 2565 3455 2585
rect 3475 2565 3480 2585
rect 3450 2535 3480 2565
rect 3450 2515 3455 2535
rect 3475 2515 3480 2535
rect 3450 2485 3480 2515
rect 3450 2465 3455 2485
rect 3475 2465 3480 2485
rect 3450 2435 3480 2465
rect 3450 2415 3455 2435
rect 3475 2415 3480 2435
rect 3450 2405 3480 2415
rect 3540 2685 3570 2695
rect 3540 2665 3545 2685
rect 3565 2665 3570 2685
rect 3540 2635 3570 2665
rect 3540 2615 3545 2635
rect 3565 2615 3570 2635
rect 3540 2585 3570 2615
rect 3540 2565 3545 2585
rect 3565 2565 3570 2585
rect 3540 2535 3570 2565
rect 3540 2515 3545 2535
rect 3565 2515 3570 2535
rect 3540 2485 3570 2515
rect 3540 2465 3545 2485
rect 3565 2465 3570 2485
rect 3540 2435 3570 2465
rect 3540 2415 3545 2435
rect 3565 2415 3570 2435
rect 3540 2405 3570 2415
rect 3630 2685 3660 2695
rect 3630 2665 3635 2685
rect 3655 2665 3660 2685
rect 3630 2635 3660 2665
rect 3630 2615 3635 2635
rect 3655 2615 3660 2635
rect 3630 2585 3660 2615
rect 3630 2565 3635 2585
rect 3655 2565 3660 2585
rect 3630 2535 3660 2565
rect 3630 2515 3635 2535
rect 3655 2515 3660 2535
rect 3630 2485 3660 2515
rect 3630 2465 3635 2485
rect 3655 2465 3660 2485
rect 3630 2435 3660 2465
rect 3630 2415 3635 2435
rect 3655 2415 3660 2435
rect 3630 2405 3660 2415
rect 3720 2685 3750 2695
rect 3720 2665 3725 2685
rect 3745 2665 3750 2685
rect 3720 2635 3750 2665
rect 3720 2615 3725 2635
rect 3745 2615 3750 2635
rect 3720 2585 3750 2615
rect 3720 2565 3725 2585
rect 3745 2565 3750 2585
rect 3720 2535 3750 2565
rect 3720 2515 3725 2535
rect 3745 2515 3750 2535
rect 3720 2485 3750 2515
rect 3720 2465 3725 2485
rect 3745 2465 3750 2485
rect 3720 2435 3750 2465
rect 3720 2415 3725 2435
rect 3745 2415 3750 2435
rect 3720 2405 3750 2415
rect 3810 2685 3840 2695
rect 3810 2665 3815 2685
rect 3835 2665 3840 2685
rect 3810 2635 3840 2665
rect 3810 2615 3815 2635
rect 3835 2615 3840 2635
rect 3810 2585 3840 2615
rect 3810 2565 3815 2585
rect 3835 2565 3840 2585
rect 3810 2535 3840 2565
rect 3810 2515 3815 2535
rect 3835 2515 3840 2535
rect 3810 2485 3840 2515
rect 3810 2465 3815 2485
rect 3835 2465 3840 2485
rect 3810 2435 3840 2465
rect 3810 2415 3815 2435
rect 3835 2415 3840 2435
rect 3810 2405 3840 2415
rect 3900 2685 3930 2695
rect 3900 2665 3905 2685
rect 3925 2665 3930 2685
rect 3900 2635 3930 2665
rect 3900 2615 3905 2635
rect 3925 2615 3930 2635
rect 3900 2585 3930 2615
rect 3900 2565 3905 2585
rect 3925 2565 3930 2585
rect 3900 2535 3930 2565
rect 3900 2515 3905 2535
rect 3925 2515 3930 2535
rect 3900 2485 3930 2515
rect 3900 2465 3905 2485
rect 3925 2465 3930 2485
rect 3900 2435 3930 2465
rect 3900 2415 3905 2435
rect 3925 2415 3930 2435
rect 3900 2405 3930 2415
rect 3990 2685 4020 2695
rect 3990 2665 3995 2685
rect 4015 2665 4020 2685
rect 3990 2635 4020 2665
rect 3990 2615 3995 2635
rect 4015 2615 4020 2635
rect 3990 2585 4020 2615
rect 3990 2565 3995 2585
rect 4015 2565 4020 2585
rect 3990 2535 4020 2565
rect 3990 2515 3995 2535
rect 4015 2515 4020 2535
rect 3990 2485 4020 2515
rect 3990 2465 3995 2485
rect 4015 2465 4020 2485
rect 3990 2435 4020 2465
rect 3990 2415 3995 2435
rect 4015 2415 4020 2435
rect 3990 2405 4020 2415
rect 4080 2685 4110 2695
rect 4080 2665 4085 2685
rect 4105 2665 4110 2685
rect 4080 2635 4110 2665
rect 4080 2615 4085 2635
rect 4105 2615 4110 2635
rect 4080 2585 4110 2615
rect 4080 2565 4085 2585
rect 4105 2565 4110 2585
rect 4080 2535 4110 2565
rect 4080 2515 4085 2535
rect 4105 2515 4110 2535
rect 4080 2485 4110 2515
rect 4080 2465 4085 2485
rect 4105 2465 4110 2485
rect 4080 2435 4110 2465
rect 4080 2415 4085 2435
rect 4105 2415 4110 2435
rect 4080 2405 4110 2415
rect 4170 2685 4200 2695
rect 4170 2665 4175 2685
rect 4195 2665 4200 2685
rect 4170 2635 4200 2665
rect 4170 2615 4175 2635
rect 4195 2615 4200 2635
rect 4170 2585 4200 2615
rect 4170 2565 4175 2585
rect 4195 2565 4200 2585
rect 4170 2535 4200 2565
rect 4170 2515 4175 2535
rect 4195 2515 4200 2535
rect 4170 2485 4200 2515
rect 4170 2465 4175 2485
rect 4195 2465 4200 2485
rect 4170 2435 4200 2465
rect 4170 2415 4175 2435
rect 4195 2415 4200 2435
rect 4170 2405 4200 2415
rect 4260 2685 4290 2695
rect 4260 2665 4265 2685
rect 4285 2665 4290 2685
rect 4260 2635 4290 2665
rect 4260 2615 4265 2635
rect 4285 2615 4290 2635
rect 4260 2585 4290 2615
rect 4260 2565 4265 2585
rect 4285 2565 4290 2585
rect 4260 2535 4290 2565
rect 4260 2515 4265 2535
rect 4285 2515 4290 2535
rect 4260 2485 4290 2515
rect 4260 2465 4265 2485
rect 4285 2465 4290 2485
rect 4260 2435 4290 2465
rect 4260 2415 4265 2435
rect 4285 2415 4290 2435
rect 4260 2405 4290 2415
rect 4350 2685 4380 2695
rect 4350 2665 4355 2685
rect 4375 2665 4380 2685
rect 4350 2635 4380 2665
rect 4350 2615 4355 2635
rect 4375 2615 4380 2635
rect 4350 2585 4380 2615
rect 4350 2565 4355 2585
rect 4375 2565 4380 2585
rect 4350 2535 4380 2565
rect 4350 2515 4355 2535
rect 4375 2515 4380 2535
rect 4350 2485 4380 2515
rect 4350 2465 4355 2485
rect 4375 2465 4380 2485
rect 4350 2435 4380 2465
rect 4350 2415 4355 2435
rect 4375 2415 4380 2435
rect 4350 2405 4380 2415
rect 4440 2685 4470 2695
rect 4440 2665 4445 2685
rect 4465 2665 4470 2685
rect 4440 2635 4470 2665
rect 4440 2615 4445 2635
rect 4465 2615 4470 2635
rect 4440 2585 4470 2615
rect 4440 2565 4445 2585
rect 4465 2565 4470 2585
rect 4440 2535 4470 2565
rect 4440 2515 4445 2535
rect 4465 2515 4470 2535
rect 4440 2485 4470 2515
rect 4440 2465 4445 2485
rect 4465 2465 4470 2485
rect 4440 2435 4470 2465
rect 4440 2415 4445 2435
rect 4465 2415 4470 2435
rect 4440 2405 4470 2415
rect 4530 2685 4560 2695
rect 4530 2665 4535 2685
rect 4555 2665 4560 2685
rect 4530 2635 4560 2665
rect 4530 2615 4535 2635
rect 4555 2615 4560 2635
rect 4530 2585 4560 2615
rect 4530 2565 4535 2585
rect 4555 2565 4560 2585
rect 4530 2535 4560 2565
rect 4530 2515 4535 2535
rect 4555 2515 4560 2535
rect 4530 2485 4560 2515
rect 4530 2465 4535 2485
rect 4555 2465 4560 2485
rect 4530 2435 4560 2465
rect 4530 2415 4535 2435
rect 4555 2415 4560 2435
rect 4530 2405 4560 2415
rect 4620 2685 4650 2695
rect 4620 2665 4625 2685
rect 4645 2665 4650 2685
rect 4620 2635 4650 2665
rect 4620 2615 4625 2635
rect 4645 2615 4650 2635
rect 4620 2585 4650 2615
rect 4620 2565 4625 2585
rect 4645 2565 4650 2585
rect 4620 2535 4650 2565
rect 4620 2515 4625 2535
rect 4645 2515 4650 2535
rect 4620 2485 4650 2515
rect 4620 2465 4625 2485
rect 4645 2465 4650 2485
rect 4620 2435 4650 2465
rect 4620 2415 4625 2435
rect 4645 2415 4650 2435
rect 4620 2405 4650 2415
rect 4710 2685 4740 2695
rect 4710 2665 4715 2685
rect 4735 2665 4740 2685
rect 4710 2635 4740 2665
rect 4710 2615 4715 2635
rect 4735 2615 4740 2635
rect 4710 2585 4740 2615
rect 4710 2565 4715 2585
rect 4735 2565 4740 2585
rect 4710 2535 4740 2565
rect 4710 2515 4715 2535
rect 4735 2515 4740 2535
rect 4710 2485 4740 2515
rect 4710 2465 4715 2485
rect 4735 2465 4740 2485
rect 4710 2435 4740 2465
rect 4710 2415 4715 2435
rect 4735 2415 4740 2435
rect 4710 2405 4740 2415
rect 4800 2685 4870 2695
rect 4800 2665 4805 2685
rect 4825 2665 4845 2685
rect 4865 2665 4870 2685
rect 15060 2680 15070 2700
rect 15090 2680 15100 2700
rect 15060 2670 15100 2680
rect 15170 2700 15210 2710
rect 15170 2680 15180 2700
rect 15200 2680 15210 2700
rect 15170 2670 15210 2680
rect 15280 2700 15320 2710
rect 15280 2680 15290 2700
rect 15310 2680 15320 2700
rect 15280 2670 15320 2680
rect 15390 2700 15430 2710
rect 15390 2680 15400 2700
rect 15420 2680 15430 2700
rect 15390 2670 15430 2680
rect 15500 2700 15540 2710
rect 15500 2680 15510 2700
rect 15530 2680 15540 2700
rect 15500 2670 15540 2680
rect 15610 2700 15650 2710
rect 15610 2680 15620 2700
rect 15640 2680 15650 2700
rect 15610 2670 15650 2680
rect 15980 2680 16050 2710
rect 4800 2635 4870 2665
rect 4800 2615 4805 2635
rect 4825 2615 4845 2635
rect 4865 2615 4870 2635
rect 4800 2585 4870 2615
rect 4800 2565 4805 2585
rect 4825 2565 4845 2585
rect 4865 2565 4870 2585
rect 4800 2535 4870 2565
rect 4800 2515 4805 2535
rect 4825 2515 4845 2535
rect 4865 2515 4870 2535
rect 4800 2485 4870 2515
rect 4800 2465 4805 2485
rect 4825 2465 4845 2485
rect 4865 2465 4870 2485
rect 4800 2435 4870 2465
rect 4800 2415 4805 2435
rect 4825 2415 4845 2435
rect 4865 2415 4870 2435
rect 4800 2405 4870 2415
rect 14640 2645 14855 2665
rect 15070 2650 15090 2670
rect 15180 2650 15200 2670
rect 15290 2650 15310 2670
rect 15400 2650 15420 2670
rect 15510 2650 15530 2670
rect 15620 2650 15640 2670
rect 15980 2660 15985 2680
rect 16005 2660 16025 2680
rect 16045 2660 16050 2680
rect 14640 2625 14675 2645
rect 14820 2625 14855 2645
rect 14735 2575 14760 2625
rect 14970 2640 15040 2650
rect 14970 2620 14975 2640
rect 14995 2620 15015 2640
rect 15035 2620 15040 2640
rect 14970 2590 15040 2620
rect 14970 2570 14975 2590
rect 14995 2570 15015 2590
rect 15035 2570 15040 2590
rect 14970 2540 15040 2570
rect 14970 2520 14975 2540
rect 14995 2520 15015 2540
rect 15035 2520 15040 2540
rect 14970 2490 15040 2520
rect 14970 2470 14975 2490
rect 14995 2470 15015 2490
rect 15035 2470 15040 2490
rect 14970 2460 15040 2470
rect 15065 2640 15095 2650
rect 15065 2620 15070 2640
rect 15090 2620 15095 2640
rect 15065 2590 15095 2620
rect 15065 2570 15070 2590
rect 15090 2570 15095 2590
rect 15065 2540 15095 2570
rect 15065 2520 15070 2540
rect 15090 2520 15095 2540
rect 15065 2490 15095 2520
rect 15065 2470 15070 2490
rect 15090 2470 15095 2490
rect 15065 2460 15095 2470
rect 15120 2640 15150 2650
rect 15120 2620 15125 2640
rect 15145 2620 15150 2640
rect 15120 2590 15150 2620
rect 15120 2570 15125 2590
rect 15145 2570 15150 2590
rect 15120 2540 15150 2570
rect 15120 2520 15125 2540
rect 15145 2520 15150 2540
rect 15120 2490 15150 2520
rect 15120 2470 15125 2490
rect 15145 2470 15150 2490
rect 15120 2460 15150 2470
rect 15175 2640 15205 2650
rect 15175 2620 15180 2640
rect 15200 2620 15205 2640
rect 15175 2590 15205 2620
rect 15175 2570 15180 2590
rect 15200 2570 15205 2590
rect 15175 2540 15205 2570
rect 15175 2520 15180 2540
rect 15200 2520 15205 2540
rect 15175 2490 15205 2520
rect 15175 2470 15180 2490
rect 15200 2470 15205 2490
rect 15175 2460 15205 2470
rect 15230 2640 15260 2650
rect 15230 2620 15235 2640
rect 15255 2620 15260 2640
rect 15230 2590 15260 2620
rect 15230 2570 15235 2590
rect 15255 2570 15260 2590
rect 15230 2540 15260 2570
rect 15230 2520 15235 2540
rect 15255 2520 15260 2540
rect 15230 2490 15260 2520
rect 15230 2470 15235 2490
rect 15255 2470 15260 2490
rect 15230 2460 15260 2470
rect 15285 2640 15315 2650
rect 15285 2620 15290 2640
rect 15310 2620 15315 2640
rect 15285 2590 15315 2620
rect 15285 2570 15290 2590
rect 15310 2570 15315 2590
rect 15285 2540 15315 2570
rect 15285 2520 15290 2540
rect 15310 2520 15315 2540
rect 15285 2490 15315 2520
rect 15285 2470 15290 2490
rect 15310 2470 15315 2490
rect 15285 2460 15315 2470
rect 15340 2640 15370 2650
rect 15340 2620 15345 2640
rect 15365 2620 15370 2640
rect 15340 2590 15370 2620
rect 15340 2570 15345 2590
rect 15365 2570 15370 2590
rect 15340 2540 15370 2570
rect 15340 2520 15345 2540
rect 15365 2520 15370 2540
rect 15340 2490 15370 2520
rect 15340 2470 15345 2490
rect 15365 2470 15370 2490
rect 15340 2460 15370 2470
rect 15395 2640 15425 2650
rect 15395 2620 15400 2640
rect 15420 2620 15425 2640
rect 15395 2590 15425 2620
rect 15395 2570 15400 2590
rect 15420 2570 15425 2590
rect 15395 2540 15425 2570
rect 15395 2520 15400 2540
rect 15420 2520 15425 2540
rect 15395 2490 15425 2520
rect 15395 2470 15400 2490
rect 15420 2470 15425 2490
rect 15395 2460 15425 2470
rect 15450 2640 15480 2650
rect 15450 2620 15455 2640
rect 15475 2620 15480 2640
rect 15450 2590 15480 2620
rect 15450 2570 15455 2590
rect 15475 2570 15480 2590
rect 15450 2540 15480 2570
rect 15450 2520 15455 2540
rect 15475 2520 15480 2540
rect 15450 2490 15480 2520
rect 15450 2470 15455 2490
rect 15475 2470 15480 2490
rect 15450 2460 15480 2470
rect 15505 2640 15535 2650
rect 15505 2620 15510 2640
rect 15530 2620 15535 2640
rect 15505 2590 15535 2620
rect 15505 2570 15510 2590
rect 15530 2570 15535 2590
rect 15505 2540 15535 2570
rect 15505 2520 15510 2540
rect 15530 2520 15535 2540
rect 15505 2490 15535 2520
rect 15505 2470 15510 2490
rect 15530 2470 15535 2490
rect 15505 2460 15535 2470
rect 15560 2640 15590 2650
rect 15560 2620 15565 2640
rect 15585 2620 15590 2640
rect 15560 2590 15590 2620
rect 15560 2570 15565 2590
rect 15585 2570 15590 2590
rect 15560 2540 15590 2570
rect 15560 2520 15565 2540
rect 15585 2520 15590 2540
rect 15560 2490 15590 2520
rect 15560 2470 15565 2490
rect 15585 2470 15590 2490
rect 15560 2460 15590 2470
rect 15615 2640 15645 2650
rect 15615 2620 15620 2640
rect 15640 2620 15645 2640
rect 15615 2590 15645 2620
rect 15615 2570 15620 2590
rect 15640 2570 15645 2590
rect 15615 2540 15645 2570
rect 15615 2520 15620 2540
rect 15640 2520 15645 2540
rect 15615 2490 15645 2520
rect 15615 2470 15620 2490
rect 15640 2470 15645 2490
rect 15615 2460 15645 2470
rect 15670 2640 15740 2650
rect 15670 2620 15675 2640
rect 15695 2620 15715 2640
rect 15735 2620 15740 2640
rect 15670 2590 15740 2620
rect 15670 2570 15675 2590
rect 15695 2570 15715 2590
rect 15735 2570 15740 2590
rect 15670 2540 15740 2570
rect 15670 2520 15675 2540
rect 15695 2520 15715 2540
rect 15735 2520 15740 2540
rect 15670 2490 15740 2520
rect 15980 2630 16050 2660
rect 15980 2610 15985 2630
rect 16005 2610 16025 2630
rect 16045 2610 16050 2630
rect 15980 2580 16050 2610
rect 15980 2560 15985 2580
rect 16005 2560 16025 2580
rect 16045 2560 16050 2580
rect 15980 2530 16050 2560
rect 15980 2510 15985 2530
rect 16005 2510 16025 2530
rect 16045 2510 16050 2530
rect 15980 2500 16050 2510
rect 16080 2830 16110 2840
rect 16080 2810 16085 2830
rect 16105 2810 16110 2830
rect 16080 2780 16110 2810
rect 16080 2760 16085 2780
rect 16105 2760 16110 2780
rect 16080 2730 16110 2760
rect 16080 2710 16085 2730
rect 16105 2710 16110 2730
rect 16080 2680 16110 2710
rect 16080 2660 16085 2680
rect 16105 2660 16110 2680
rect 16080 2630 16110 2660
rect 16080 2610 16085 2630
rect 16105 2610 16110 2630
rect 16080 2580 16110 2610
rect 16080 2560 16085 2580
rect 16105 2560 16110 2580
rect 16080 2530 16110 2560
rect 16080 2510 16085 2530
rect 16105 2510 16110 2530
rect 16080 2500 16110 2510
rect 16140 2830 16170 2840
rect 16140 2810 16145 2830
rect 16165 2810 16170 2830
rect 16140 2780 16170 2810
rect 16140 2760 16145 2780
rect 16165 2760 16170 2780
rect 16140 2730 16170 2760
rect 16140 2710 16145 2730
rect 16165 2710 16170 2730
rect 16140 2680 16170 2710
rect 16140 2660 16145 2680
rect 16165 2660 16170 2680
rect 16140 2630 16170 2660
rect 16140 2610 16145 2630
rect 16165 2610 16170 2630
rect 16140 2580 16170 2610
rect 16140 2560 16145 2580
rect 16165 2560 16170 2580
rect 16140 2530 16170 2560
rect 16140 2510 16145 2530
rect 16165 2510 16170 2530
rect 16140 2500 16170 2510
rect 16200 2830 16230 2840
rect 16200 2810 16205 2830
rect 16225 2810 16230 2830
rect 16200 2780 16230 2810
rect 16200 2760 16205 2780
rect 16225 2760 16230 2780
rect 16200 2730 16230 2760
rect 16200 2710 16205 2730
rect 16225 2710 16230 2730
rect 16200 2680 16230 2710
rect 16200 2660 16205 2680
rect 16225 2660 16230 2680
rect 16200 2630 16230 2660
rect 16200 2610 16205 2630
rect 16225 2610 16230 2630
rect 16200 2580 16230 2610
rect 16200 2560 16205 2580
rect 16225 2560 16230 2580
rect 16200 2530 16230 2560
rect 16200 2510 16205 2530
rect 16225 2510 16230 2530
rect 16200 2500 16230 2510
rect 16260 2830 16290 2840
rect 16260 2810 16265 2830
rect 16285 2810 16290 2830
rect 16260 2780 16290 2810
rect 16260 2760 16265 2780
rect 16285 2760 16290 2780
rect 16260 2730 16290 2760
rect 16260 2710 16265 2730
rect 16285 2710 16290 2730
rect 16260 2680 16290 2710
rect 16260 2660 16265 2680
rect 16285 2660 16290 2680
rect 16260 2630 16290 2660
rect 16260 2610 16265 2630
rect 16285 2610 16290 2630
rect 16260 2580 16290 2610
rect 16260 2560 16265 2580
rect 16285 2560 16290 2580
rect 16260 2530 16290 2560
rect 16260 2510 16265 2530
rect 16285 2510 16290 2530
rect 16260 2500 16290 2510
rect 16320 2830 16350 2840
rect 16320 2810 16325 2830
rect 16345 2810 16350 2830
rect 16320 2780 16350 2810
rect 16320 2760 16325 2780
rect 16345 2760 16350 2780
rect 16320 2730 16350 2760
rect 16320 2710 16325 2730
rect 16345 2710 16350 2730
rect 16320 2680 16350 2710
rect 16320 2660 16325 2680
rect 16345 2660 16350 2680
rect 16320 2630 16350 2660
rect 16320 2610 16325 2630
rect 16345 2610 16350 2630
rect 16320 2580 16350 2610
rect 16320 2560 16325 2580
rect 16345 2560 16350 2580
rect 16320 2530 16350 2560
rect 16320 2510 16325 2530
rect 16345 2510 16350 2530
rect 16320 2500 16350 2510
rect 16380 2830 16410 2840
rect 16380 2810 16385 2830
rect 16405 2810 16410 2830
rect 16380 2780 16410 2810
rect 16380 2760 16385 2780
rect 16405 2760 16410 2780
rect 16380 2730 16410 2760
rect 16380 2710 16385 2730
rect 16405 2710 16410 2730
rect 16380 2680 16410 2710
rect 16380 2660 16385 2680
rect 16405 2660 16410 2680
rect 16380 2630 16410 2660
rect 16380 2610 16385 2630
rect 16405 2610 16410 2630
rect 16380 2580 16410 2610
rect 16380 2560 16385 2580
rect 16405 2560 16410 2580
rect 16380 2530 16410 2560
rect 16380 2510 16385 2530
rect 16405 2510 16410 2530
rect 16380 2500 16410 2510
rect 16440 2830 16470 2840
rect 16440 2810 16445 2830
rect 16465 2810 16470 2830
rect 16440 2780 16470 2810
rect 16440 2760 16445 2780
rect 16465 2760 16470 2780
rect 16440 2730 16470 2760
rect 16440 2710 16445 2730
rect 16465 2710 16470 2730
rect 16440 2680 16470 2710
rect 16440 2660 16445 2680
rect 16465 2660 16470 2680
rect 16440 2630 16470 2660
rect 16440 2610 16445 2630
rect 16465 2610 16470 2630
rect 16440 2580 16470 2610
rect 16440 2560 16445 2580
rect 16465 2560 16470 2580
rect 16440 2530 16470 2560
rect 16440 2510 16445 2530
rect 16465 2510 16470 2530
rect 16440 2500 16470 2510
rect 16500 2830 16530 2840
rect 16500 2810 16505 2830
rect 16525 2810 16530 2830
rect 16500 2780 16530 2810
rect 16500 2760 16505 2780
rect 16525 2760 16530 2780
rect 16500 2730 16530 2760
rect 16500 2710 16505 2730
rect 16525 2710 16530 2730
rect 16500 2680 16530 2710
rect 16500 2660 16505 2680
rect 16525 2660 16530 2680
rect 16500 2630 16530 2660
rect 16500 2610 16505 2630
rect 16525 2610 16530 2630
rect 16500 2580 16530 2610
rect 16500 2560 16505 2580
rect 16525 2560 16530 2580
rect 16500 2530 16530 2560
rect 16500 2510 16505 2530
rect 16525 2510 16530 2530
rect 16500 2500 16530 2510
rect 16560 2830 16590 2840
rect 16560 2810 16565 2830
rect 16585 2810 16590 2830
rect 16560 2780 16590 2810
rect 16560 2760 16565 2780
rect 16585 2760 16590 2780
rect 16560 2730 16590 2760
rect 16560 2710 16565 2730
rect 16585 2710 16590 2730
rect 16560 2680 16590 2710
rect 16560 2660 16565 2680
rect 16585 2660 16590 2680
rect 16560 2630 16590 2660
rect 16560 2610 16565 2630
rect 16585 2610 16590 2630
rect 16560 2580 16590 2610
rect 16560 2560 16565 2580
rect 16585 2560 16590 2580
rect 16560 2530 16590 2560
rect 16560 2510 16565 2530
rect 16585 2510 16590 2530
rect 16560 2500 16590 2510
rect 16620 2830 16650 2840
rect 16620 2810 16625 2830
rect 16645 2810 16650 2830
rect 16620 2780 16650 2810
rect 16620 2760 16625 2780
rect 16645 2760 16650 2780
rect 16620 2730 16650 2760
rect 16620 2710 16625 2730
rect 16645 2710 16650 2730
rect 16620 2680 16650 2710
rect 16620 2660 16625 2680
rect 16645 2660 16650 2680
rect 16620 2630 16650 2660
rect 16620 2610 16625 2630
rect 16645 2610 16650 2630
rect 16620 2580 16650 2610
rect 16620 2560 16625 2580
rect 16645 2560 16650 2580
rect 16620 2530 16650 2560
rect 16620 2510 16625 2530
rect 16645 2510 16650 2530
rect 16620 2500 16650 2510
rect 16680 2830 16710 2840
rect 16680 2810 16685 2830
rect 16705 2810 16710 2830
rect 16680 2780 16710 2810
rect 16680 2760 16685 2780
rect 16705 2760 16710 2780
rect 16680 2730 16710 2760
rect 16680 2710 16685 2730
rect 16705 2710 16710 2730
rect 16680 2680 16710 2710
rect 16680 2660 16685 2680
rect 16705 2660 16710 2680
rect 16680 2630 16710 2660
rect 16680 2610 16685 2630
rect 16705 2610 16710 2630
rect 16680 2580 16710 2610
rect 16680 2560 16685 2580
rect 16705 2560 16710 2580
rect 16680 2530 16710 2560
rect 16680 2510 16685 2530
rect 16705 2510 16710 2530
rect 16680 2500 16710 2510
rect 16740 2830 16810 2840
rect 16740 2810 16745 2830
rect 16765 2810 16785 2830
rect 16805 2810 16810 2830
rect 16740 2780 16810 2810
rect 16740 2760 16745 2780
rect 16765 2760 16785 2780
rect 16805 2760 16810 2780
rect 16740 2730 16810 2760
rect 16740 2710 16745 2730
rect 16765 2710 16785 2730
rect 16805 2710 16810 2730
rect 16740 2680 16810 2710
rect 16740 2660 16745 2680
rect 16765 2660 16785 2680
rect 16805 2660 16810 2680
rect 16740 2630 16810 2660
rect 16740 2610 16745 2630
rect 16765 2610 16785 2630
rect 16805 2610 16810 2630
rect 16740 2580 16810 2610
rect 16740 2560 16745 2580
rect 16765 2560 16785 2580
rect 16805 2560 16810 2580
rect 16740 2530 16810 2560
rect 16740 2510 16745 2530
rect 16765 2510 16785 2530
rect 16805 2510 16810 2530
rect 16740 2500 16810 2510
rect 16990 2830 17060 2840
rect 16990 2810 16995 2830
rect 17015 2810 17035 2830
rect 17055 2810 17060 2830
rect 16990 2780 17060 2810
rect 16990 2760 16995 2780
rect 17015 2760 17035 2780
rect 17055 2760 17060 2780
rect 16990 2730 17060 2760
rect 16990 2710 16995 2730
rect 17015 2710 17035 2730
rect 17055 2710 17060 2730
rect 16990 2680 17060 2710
rect 16990 2660 16995 2680
rect 17015 2660 17035 2680
rect 17055 2660 17060 2680
rect 16990 2630 17060 2660
rect 16990 2610 16995 2630
rect 17015 2610 17035 2630
rect 17055 2610 17060 2630
rect 16990 2580 17060 2610
rect 16990 2560 16995 2580
rect 17015 2560 17035 2580
rect 17055 2560 17060 2580
rect 16990 2530 17060 2560
rect 16990 2510 16995 2530
rect 17015 2510 17035 2530
rect 17055 2510 17060 2530
rect 16990 2500 17060 2510
rect 17090 2830 17120 2840
rect 17090 2810 17095 2830
rect 17115 2810 17120 2830
rect 17090 2780 17120 2810
rect 17090 2760 17095 2780
rect 17115 2760 17120 2780
rect 17090 2730 17120 2760
rect 17090 2710 17095 2730
rect 17115 2710 17120 2730
rect 17090 2680 17120 2710
rect 17090 2660 17095 2680
rect 17115 2660 17120 2680
rect 17090 2630 17120 2660
rect 17090 2610 17095 2630
rect 17115 2610 17120 2630
rect 17090 2580 17120 2610
rect 17090 2560 17095 2580
rect 17115 2560 17120 2580
rect 17090 2530 17120 2560
rect 17090 2510 17095 2530
rect 17115 2510 17120 2530
rect 17090 2500 17120 2510
rect 17150 2830 17180 2840
rect 17150 2810 17155 2830
rect 17175 2810 17180 2830
rect 17150 2780 17180 2810
rect 17150 2760 17155 2780
rect 17175 2760 17180 2780
rect 17150 2730 17180 2760
rect 17150 2710 17155 2730
rect 17175 2710 17180 2730
rect 17150 2680 17180 2710
rect 17150 2660 17155 2680
rect 17175 2660 17180 2680
rect 17150 2630 17180 2660
rect 17150 2610 17155 2630
rect 17175 2610 17180 2630
rect 17150 2580 17180 2610
rect 17150 2560 17155 2580
rect 17175 2560 17180 2580
rect 17150 2530 17180 2560
rect 17150 2510 17155 2530
rect 17175 2510 17180 2530
rect 17150 2500 17180 2510
rect 17210 2830 17240 2840
rect 17210 2810 17215 2830
rect 17235 2810 17240 2830
rect 17210 2780 17240 2810
rect 17210 2760 17215 2780
rect 17235 2760 17240 2780
rect 17210 2730 17240 2760
rect 17210 2710 17215 2730
rect 17235 2710 17240 2730
rect 17210 2680 17240 2710
rect 17210 2660 17215 2680
rect 17235 2660 17240 2680
rect 17210 2630 17240 2660
rect 17210 2610 17215 2630
rect 17235 2610 17240 2630
rect 17210 2580 17240 2610
rect 17210 2560 17215 2580
rect 17235 2560 17240 2580
rect 17210 2530 17240 2560
rect 17210 2510 17215 2530
rect 17235 2510 17240 2530
rect 17210 2500 17240 2510
rect 17270 2830 17300 2840
rect 17270 2810 17275 2830
rect 17295 2810 17300 2830
rect 17270 2780 17300 2810
rect 17270 2760 17275 2780
rect 17295 2760 17300 2780
rect 17270 2730 17300 2760
rect 17270 2710 17275 2730
rect 17295 2710 17300 2730
rect 17270 2680 17300 2710
rect 17270 2660 17275 2680
rect 17295 2660 17300 2680
rect 17270 2630 17300 2660
rect 17270 2610 17275 2630
rect 17295 2610 17300 2630
rect 17270 2580 17300 2610
rect 17270 2560 17275 2580
rect 17295 2560 17300 2580
rect 17270 2530 17300 2560
rect 17270 2510 17275 2530
rect 17295 2510 17300 2530
rect 17270 2500 17300 2510
rect 17330 2830 17360 2840
rect 17330 2810 17335 2830
rect 17355 2810 17360 2830
rect 17330 2780 17360 2810
rect 17330 2760 17335 2780
rect 17355 2760 17360 2780
rect 17330 2730 17360 2760
rect 17330 2710 17335 2730
rect 17355 2710 17360 2730
rect 17330 2680 17360 2710
rect 17330 2660 17335 2680
rect 17355 2660 17360 2680
rect 17330 2630 17360 2660
rect 17330 2610 17335 2630
rect 17355 2610 17360 2630
rect 17330 2580 17360 2610
rect 17330 2560 17335 2580
rect 17355 2560 17360 2580
rect 17330 2530 17360 2560
rect 17330 2510 17335 2530
rect 17355 2510 17360 2530
rect 17330 2500 17360 2510
rect 17390 2830 17420 2840
rect 17390 2810 17395 2830
rect 17415 2810 17420 2830
rect 17390 2780 17420 2810
rect 17390 2760 17395 2780
rect 17415 2760 17420 2780
rect 17390 2730 17420 2760
rect 17390 2710 17395 2730
rect 17415 2710 17420 2730
rect 17390 2680 17420 2710
rect 17390 2660 17395 2680
rect 17415 2660 17420 2680
rect 17390 2630 17420 2660
rect 17390 2610 17395 2630
rect 17415 2610 17420 2630
rect 17390 2580 17420 2610
rect 17390 2560 17395 2580
rect 17415 2560 17420 2580
rect 17390 2530 17420 2560
rect 17390 2510 17395 2530
rect 17415 2510 17420 2530
rect 17390 2500 17420 2510
rect 17450 2830 17480 2840
rect 17450 2810 17455 2830
rect 17475 2810 17480 2830
rect 17450 2780 17480 2810
rect 17450 2760 17455 2780
rect 17475 2760 17480 2780
rect 17450 2730 17480 2760
rect 17450 2710 17455 2730
rect 17475 2710 17480 2730
rect 17450 2680 17480 2710
rect 17450 2660 17455 2680
rect 17475 2660 17480 2680
rect 17450 2630 17480 2660
rect 17450 2610 17455 2630
rect 17475 2610 17480 2630
rect 17450 2580 17480 2610
rect 17450 2560 17455 2580
rect 17475 2560 17480 2580
rect 17450 2530 17480 2560
rect 17450 2510 17455 2530
rect 17475 2510 17480 2530
rect 17450 2500 17480 2510
rect 17510 2830 17540 2840
rect 17510 2810 17515 2830
rect 17535 2810 17540 2830
rect 17510 2780 17540 2810
rect 17510 2760 17515 2780
rect 17535 2760 17540 2780
rect 17510 2730 17540 2760
rect 17510 2710 17515 2730
rect 17535 2710 17540 2730
rect 17510 2680 17540 2710
rect 17510 2660 17515 2680
rect 17535 2660 17540 2680
rect 17510 2630 17540 2660
rect 17510 2610 17515 2630
rect 17535 2610 17540 2630
rect 17510 2580 17540 2610
rect 17510 2560 17515 2580
rect 17535 2560 17540 2580
rect 17510 2530 17540 2560
rect 17510 2510 17515 2530
rect 17535 2510 17540 2530
rect 17510 2500 17540 2510
rect 17570 2830 17600 2840
rect 17570 2810 17575 2830
rect 17595 2810 17600 2830
rect 17570 2780 17600 2810
rect 17570 2760 17575 2780
rect 17595 2760 17600 2780
rect 17570 2730 17600 2760
rect 17570 2710 17575 2730
rect 17595 2710 17600 2730
rect 17570 2680 17600 2710
rect 17570 2660 17575 2680
rect 17595 2660 17600 2680
rect 17570 2630 17600 2660
rect 17570 2610 17575 2630
rect 17595 2610 17600 2630
rect 17570 2580 17600 2610
rect 17570 2560 17575 2580
rect 17595 2560 17600 2580
rect 17570 2530 17600 2560
rect 17570 2510 17575 2530
rect 17595 2510 17600 2530
rect 17570 2500 17600 2510
rect 17630 2830 17660 2840
rect 17630 2810 17635 2830
rect 17655 2810 17660 2830
rect 17630 2780 17660 2810
rect 17630 2760 17635 2780
rect 17655 2760 17660 2780
rect 17630 2730 17660 2760
rect 17630 2710 17635 2730
rect 17655 2710 17660 2730
rect 17630 2680 17660 2710
rect 17630 2660 17635 2680
rect 17655 2660 17660 2680
rect 17630 2630 17660 2660
rect 17630 2610 17635 2630
rect 17655 2610 17660 2630
rect 17630 2580 17660 2610
rect 17630 2560 17635 2580
rect 17655 2560 17660 2580
rect 17630 2530 17660 2560
rect 17630 2510 17635 2530
rect 17655 2510 17660 2530
rect 17630 2500 17660 2510
rect 17690 2830 17720 2840
rect 17690 2810 17695 2830
rect 17715 2810 17720 2830
rect 17690 2780 17720 2810
rect 17690 2760 17695 2780
rect 17715 2760 17720 2780
rect 17690 2730 17720 2760
rect 17690 2710 17695 2730
rect 17715 2710 17720 2730
rect 17690 2680 17720 2710
rect 17690 2660 17695 2680
rect 17715 2660 17720 2680
rect 17690 2630 17720 2660
rect 17690 2610 17695 2630
rect 17715 2610 17720 2630
rect 17690 2580 17720 2610
rect 17690 2560 17695 2580
rect 17715 2560 17720 2580
rect 17690 2530 17720 2560
rect 17690 2510 17695 2530
rect 17715 2510 17720 2530
rect 17690 2500 17720 2510
rect 17750 2830 17820 2840
rect 17750 2810 17755 2830
rect 17775 2810 17795 2830
rect 17815 2810 17820 2830
rect 17750 2780 17820 2810
rect 17750 2760 17755 2780
rect 17775 2760 17795 2780
rect 17815 2760 17820 2780
rect 17750 2730 17820 2760
rect 17750 2710 17755 2730
rect 17775 2710 17795 2730
rect 17815 2710 17820 2730
rect 25980 2830 26050 2840
rect 25980 2810 25985 2830
rect 26005 2810 26025 2830
rect 26045 2810 26050 2830
rect 25980 2780 26050 2810
rect 25980 2760 25985 2780
rect 26005 2760 26025 2780
rect 26045 2760 26050 2780
rect 25980 2730 26050 2760
rect 25980 2710 25985 2730
rect 26005 2710 26025 2730
rect 26045 2710 26050 2730
rect 17750 2680 17820 2710
rect 17750 2660 17755 2680
rect 17775 2660 17795 2680
rect 17815 2660 17820 2680
rect 18200 2700 18240 2710
rect 18200 2680 18210 2700
rect 18230 2680 18240 2700
rect 18200 2670 18240 2680
rect 18310 2700 18350 2710
rect 18310 2680 18320 2700
rect 18340 2680 18350 2700
rect 18310 2670 18350 2680
rect 18420 2700 18460 2710
rect 18420 2680 18430 2700
rect 18450 2680 18460 2700
rect 18420 2670 18460 2680
rect 18530 2700 18570 2710
rect 18530 2680 18540 2700
rect 18560 2680 18570 2700
rect 18530 2670 18570 2680
rect 18640 2700 18680 2710
rect 18640 2680 18650 2700
rect 18670 2680 18680 2700
rect 18640 2670 18680 2680
rect 18750 2700 18790 2710
rect 18750 2680 18760 2700
rect 18780 2680 18790 2700
rect 18750 2670 18790 2680
rect 25060 2700 25100 2710
rect 25060 2680 25070 2700
rect 25090 2680 25100 2700
rect 25060 2670 25100 2680
rect 25170 2700 25210 2710
rect 25170 2680 25180 2700
rect 25200 2680 25210 2700
rect 25170 2670 25210 2680
rect 25280 2700 25320 2710
rect 25280 2680 25290 2700
rect 25310 2680 25320 2700
rect 25280 2670 25320 2680
rect 25390 2700 25430 2710
rect 25390 2680 25400 2700
rect 25420 2680 25430 2700
rect 25390 2670 25430 2680
rect 25500 2700 25540 2710
rect 25500 2680 25510 2700
rect 25530 2680 25540 2700
rect 25500 2670 25540 2680
rect 25610 2700 25650 2710
rect 25610 2680 25620 2700
rect 25640 2680 25650 2700
rect 25610 2670 25650 2680
rect 25980 2680 26050 2710
rect 17750 2630 17820 2660
rect 18210 2650 18230 2670
rect 18320 2650 18340 2670
rect 18430 2650 18450 2670
rect 18540 2650 18560 2670
rect 18650 2650 18670 2670
rect 18760 2650 18780 2670
rect 17750 2610 17755 2630
rect 17775 2610 17795 2630
rect 17815 2610 17820 2630
rect 17750 2580 17820 2610
rect 17750 2560 17755 2580
rect 17775 2560 17795 2580
rect 17815 2560 17820 2580
rect 17750 2530 17820 2560
rect 17750 2510 17755 2530
rect 17775 2510 17795 2530
rect 17815 2510 17820 2530
rect 17750 2500 17820 2510
rect 18110 2640 18180 2650
rect 18110 2620 18115 2640
rect 18135 2620 18155 2640
rect 18175 2620 18180 2640
rect 18110 2590 18180 2620
rect 18110 2570 18115 2590
rect 18135 2570 18155 2590
rect 18175 2570 18180 2590
rect 18110 2540 18180 2570
rect 18110 2520 18115 2540
rect 18135 2520 18155 2540
rect 18175 2520 18180 2540
rect 15670 2470 15675 2490
rect 15695 2470 15715 2490
rect 15735 2470 15740 2490
rect 16085 2480 16105 2500
rect 16205 2480 16225 2500
rect 16325 2480 16345 2500
rect 16445 2480 16465 2500
rect 16565 2480 16585 2500
rect 16685 2480 16705 2500
rect 17095 2480 17115 2500
rect 17215 2480 17235 2500
rect 17335 2480 17355 2500
rect 17455 2480 17475 2500
rect 17575 2480 17595 2500
rect 17695 2480 17715 2500
rect 18110 2490 18180 2520
rect 15670 2460 15740 2470
rect 16075 2470 16115 2480
rect 14975 2440 14995 2460
rect 15125 2440 15145 2460
rect 15235 2440 15255 2460
rect 15345 2440 15365 2460
rect 15455 2440 15475 2460
rect 15565 2440 15585 2460
rect 15715 2440 15735 2460
rect 16075 2450 16085 2470
rect 16105 2450 16115 2470
rect 16075 2440 16115 2450
rect 16195 2470 16235 2480
rect 16195 2450 16205 2470
rect 16225 2450 16235 2470
rect 16195 2440 16235 2450
rect 16315 2470 16355 2480
rect 16315 2450 16325 2470
rect 16345 2450 16355 2470
rect 16315 2440 16355 2450
rect 16378 2470 16412 2480
rect 16378 2450 16386 2470
rect 16404 2450 16412 2470
rect 16378 2440 16412 2450
rect 16435 2470 16475 2480
rect 16435 2450 16445 2470
rect 16465 2450 16475 2470
rect 16435 2440 16475 2450
rect 16555 2470 16595 2480
rect 16555 2450 16565 2470
rect 16585 2450 16595 2470
rect 16555 2440 16595 2450
rect 16675 2470 16715 2480
rect 16675 2450 16685 2470
rect 16705 2450 16715 2470
rect 16675 2440 16715 2450
rect 17085 2470 17125 2480
rect 17085 2450 17095 2470
rect 17115 2450 17125 2470
rect 17085 2440 17125 2450
rect 17205 2470 17245 2480
rect 17205 2450 17215 2470
rect 17235 2450 17245 2470
rect 17205 2440 17245 2450
rect 17325 2470 17365 2480
rect 17325 2450 17335 2470
rect 17355 2450 17365 2470
rect 17325 2440 17365 2450
rect 17388 2470 17422 2480
rect 17388 2450 17396 2470
rect 17414 2450 17422 2470
rect 17388 2440 17422 2450
rect 17445 2470 17485 2480
rect 17445 2450 17455 2470
rect 17475 2450 17485 2470
rect 17445 2440 17485 2450
rect 17565 2470 17605 2480
rect 17565 2450 17575 2470
rect 17595 2450 17605 2470
rect 17565 2440 17605 2450
rect 17685 2470 17725 2480
rect 17685 2450 17695 2470
rect 17715 2450 17725 2470
rect 18110 2470 18115 2490
rect 18135 2470 18155 2490
rect 18175 2470 18180 2490
rect 18110 2460 18180 2470
rect 18205 2640 18235 2650
rect 18205 2620 18210 2640
rect 18230 2620 18235 2640
rect 18205 2590 18235 2620
rect 18205 2570 18210 2590
rect 18230 2570 18235 2590
rect 18205 2540 18235 2570
rect 18205 2520 18210 2540
rect 18230 2520 18235 2540
rect 18205 2490 18235 2520
rect 18205 2470 18210 2490
rect 18230 2470 18235 2490
rect 18205 2460 18235 2470
rect 18260 2640 18290 2650
rect 18260 2620 18265 2640
rect 18285 2620 18290 2640
rect 18260 2590 18290 2620
rect 18260 2570 18265 2590
rect 18285 2570 18290 2590
rect 18260 2540 18290 2570
rect 18260 2520 18265 2540
rect 18285 2520 18290 2540
rect 18260 2490 18290 2520
rect 18260 2470 18265 2490
rect 18285 2470 18290 2490
rect 18260 2460 18290 2470
rect 18315 2640 18345 2650
rect 18315 2620 18320 2640
rect 18340 2620 18345 2640
rect 18315 2590 18345 2620
rect 18315 2570 18320 2590
rect 18340 2570 18345 2590
rect 18315 2540 18345 2570
rect 18315 2520 18320 2540
rect 18340 2520 18345 2540
rect 18315 2490 18345 2520
rect 18315 2470 18320 2490
rect 18340 2470 18345 2490
rect 18315 2460 18345 2470
rect 18370 2640 18400 2650
rect 18370 2620 18375 2640
rect 18395 2620 18400 2640
rect 18370 2590 18400 2620
rect 18370 2570 18375 2590
rect 18395 2570 18400 2590
rect 18370 2540 18400 2570
rect 18370 2520 18375 2540
rect 18395 2520 18400 2540
rect 18370 2490 18400 2520
rect 18370 2470 18375 2490
rect 18395 2470 18400 2490
rect 18370 2460 18400 2470
rect 18425 2640 18455 2650
rect 18425 2620 18430 2640
rect 18450 2620 18455 2640
rect 18425 2590 18455 2620
rect 18425 2570 18430 2590
rect 18450 2570 18455 2590
rect 18425 2540 18455 2570
rect 18425 2520 18430 2540
rect 18450 2520 18455 2540
rect 18425 2490 18455 2520
rect 18425 2470 18430 2490
rect 18450 2470 18455 2490
rect 18425 2460 18455 2470
rect 18480 2640 18510 2650
rect 18480 2620 18485 2640
rect 18505 2620 18510 2640
rect 18480 2590 18510 2620
rect 18480 2570 18485 2590
rect 18505 2570 18510 2590
rect 18480 2540 18510 2570
rect 18480 2520 18485 2540
rect 18505 2520 18510 2540
rect 18480 2490 18510 2520
rect 18480 2470 18485 2490
rect 18505 2470 18510 2490
rect 18480 2460 18510 2470
rect 18535 2640 18565 2650
rect 18535 2620 18540 2640
rect 18560 2620 18565 2640
rect 18535 2590 18565 2620
rect 18535 2570 18540 2590
rect 18560 2570 18565 2590
rect 18535 2540 18565 2570
rect 18535 2520 18540 2540
rect 18560 2520 18565 2540
rect 18535 2490 18565 2520
rect 18535 2470 18540 2490
rect 18560 2470 18565 2490
rect 18535 2460 18565 2470
rect 18590 2640 18620 2650
rect 18590 2620 18595 2640
rect 18615 2620 18620 2640
rect 18590 2590 18620 2620
rect 18590 2570 18595 2590
rect 18615 2570 18620 2590
rect 18590 2540 18620 2570
rect 18590 2520 18595 2540
rect 18615 2520 18620 2540
rect 18590 2490 18620 2520
rect 18590 2470 18595 2490
rect 18615 2470 18620 2490
rect 18590 2460 18620 2470
rect 18645 2640 18675 2650
rect 18645 2620 18650 2640
rect 18670 2620 18675 2640
rect 18645 2590 18675 2620
rect 18645 2570 18650 2590
rect 18670 2570 18675 2590
rect 18645 2540 18675 2570
rect 18645 2520 18650 2540
rect 18670 2520 18675 2540
rect 18645 2490 18675 2520
rect 18645 2470 18650 2490
rect 18670 2470 18675 2490
rect 18645 2460 18675 2470
rect 18700 2640 18730 2650
rect 18700 2620 18705 2640
rect 18725 2620 18730 2640
rect 18700 2590 18730 2620
rect 18700 2570 18705 2590
rect 18725 2570 18730 2590
rect 18700 2540 18730 2570
rect 18700 2520 18705 2540
rect 18725 2520 18730 2540
rect 18700 2490 18730 2520
rect 18700 2470 18705 2490
rect 18725 2470 18730 2490
rect 18700 2460 18730 2470
rect 18755 2640 18785 2650
rect 18755 2620 18760 2640
rect 18780 2620 18785 2640
rect 18755 2590 18785 2620
rect 18755 2570 18760 2590
rect 18780 2570 18785 2590
rect 18755 2540 18785 2570
rect 18755 2520 18760 2540
rect 18780 2520 18785 2540
rect 18755 2490 18785 2520
rect 18755 2470 18760 2490
rect 18780 2470 18785 2490
rect 18755 2460 18785 2470
rect 18810 2640 18880 2650
rect 18810 2620 18815 2640
rect 18835 2620 18855 2640
rect 18875 2620 18880 2640
rect 18810 2590 18880 2620
rect 18810 2570 18815 2590
rect 18835 2570 18855 2590
rect 18875 2570 18880 2590
rect 18810 2540 18880 2570
rect 18810 2520 18815 2540
rect 18835 2520 18855 2540
rect 18875 2520 18880 2540
rect 18810 2490 18880 2520
rect 18810 2470 18815 2490
rect 18835 2470 18855 2490
rect 18875 2470 18880 2490
rect 18810 2460 18880 2470
rect 18995 2645 19210 2665
rect 18995 2625 19030 2645
rect 19175 2625 19210 2645
rect 17685 2440 17725 2450
rect 18115 2440 18135 2460
rect 18265 2440 18285 2460
rect 18375 2440 18395 2460
rect 18485 2440 18505 2460
rect 18595 2440 18615 2460
rect 18705 2440 18725 2460
rect 18855 2440 18875 2460
rect 14965 2430 15005 2440
rect 14965 2410 14975 2430
rect 14995 2410 15005 2430
rect 3275 2385 3295 2405
rect 3455 2385 3475 2405
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2370 3395 2380
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 2625 2315 2655 2345
rect 3355 2340 3395 2350
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3635 2340 3655 2405
rect 3815 2385 3835 2405
rect 3995 2385 4015 2405
rect 4175 2385 4195 2405
rect 3805 2375 3845 2385
rect 3805 2355 3815 2375
rect 3835 2355 3845 2375
rect 3805 2345 3845 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2375 4205 2385
rect 4165 2355 4175 2375
rect 4195 2355 4205 2375
rect 4165 2345 4205 2355
rect 4355 2340 4375 2405
rect 4535 2385 4555 2405
rect 4715 2385 4735 2405
rect 14965 2400 15005 2410
rect 15115 2430 15155 2440
rect 15115 2410 15125 2430
rect 15145 2410 15155 2430
rect 15115 2400 15155 2410
rect 15225 2430 15265 2440
rect 15225 2410 15235 2430
rect 15255 2410 15265 2430
rect 15225 2400 15265 2410
rect 15335 2430 15375 2440
rect 15335 2410 15345 2430
rect 15365 2410 15375 2430
rect 15335 2400 15375 2410
rect 15445 2430 15485 2440
rect 15445 2410 15455 2430
rect 15475 2410 15485 2430
rect 15445 2400 15485 2410
rect 15555 2430 15595 2440
rect 15555 2410 15565 2430
rect 15585 2410 15595 2430
rect 15555 2400 15595 2410
rect 15705 2430 15745 2440
rect 15705 2410 15715 2430
rect 15735 2410 15745 2430
rect 15705 2400 15745 2410
rect 18105 2430 18145 2440
rect 18105 2410 18115 2430
rect 18135 2410 18145 2430
rect 18105 2400 18145 2410
rect 18255 2430 18295 2440
rect 18255 2410 18265 2430
rect 18285 2410 18295 2430
rect 18255 2400 18295 2410
rect 18365 2430 18405 2440
rect 18365 2410 18375 2430
rect 18395 2410 18405 2430
rect 18365 2400 18405 2410
rect 18475 2430 18515 2440
rect 18475 2410 18485 2430
rect 18505 2410 18515 2430
rect 18475 2400 18515 2410
rect 18585 2430 18625 2440
rect 18585 2410 18595 2430
rect 18615 2410 18625 2430
rect 18585 2400 18625 2410
rect 18695 2430 18735 2440
rect 18695 2410 18705 2430
rect 18725 2410 18735 2430
rect 18695 2400 18735 2410
rect 18845 2430 18885 2440
rect 18845 2410 18855 2430
rect 18875 2410 18885 2430
rect 18845 2400 18885 2410
rect 19090 2575 19115 2625
rect 24640 2645 24855 2665
rect 25070 2650 25090 2670
rect 25180 2650 25200 2670
rect 25290 2650 25310 2670
rect 25400 2650 25420 2670
rect 25510 2650 25530 2670
rect 25620 2650 25640 2670
rect 25980 2660 25985 2680
rect 26005 2660 26025 2680
rect 26045 2660 26050 2680
rect 24640 2625 24675 2645
rect 24820 2625 24855 2645
rect 24735 2575 24760 2625
rect 24970 2640 25040 2650
rect 24970 2620 24975 2640
rect 24995 2620 25015 2640
rect 25035 2620 25040 2640
rect 24970 2590 25040 2620
rect 24970 2570 24975 2590
rect 24995 2570 25015 2590
rect 25035 2570 25040 2590
rect 24970 2540 25040 2570
rect 24970 2520 24975 2540
rect 24995 2520 25015 2540
rect 25035 2520 25040 2540
rect 24970 2490 25040 2520
rect 24970 2470 24975 2490
rect 24995 2470 25015 2490
rect 25035 2470 25040 2490
rect 24970 2460 25040 2470
rect 25065 2640 25095 2650
rect 25065 2620 25070 2640
rect 25090 2620 25095 2640
rect 25065 2590 25095 2620
rect 25065 2570 25070 2590
rect 25090 2570 25095 2590
rect 25065 2540 25095 2570
rect 25065 2520 25070 2540
rect 25090 2520 25095 2540
rect 25065 2490 25095 2520
rect 25065 2470 25070 2490
rect 25090 2470 25095 2490
rect 25065 2460 25095 2470
rect 25120 2640 25150 2650
rect 25120 2620 25125 2640
rect 25145 2620 25150 2640
rect 25120 2590 25150 2620
rect 25120 2570 25125 2590
rect 25145 2570 25150 2590
rect 25120 2540 25150 2570
rect 25120 2520 25125 2540
rect 25145 2520 25150 2540
rect 25120 2490 25150 2520
rect 25120 2470 25125 2490
rect 25145 2470 25150 2490
rect 25120 2460 25150 2470
rect 25175 2640 25205 2650
rect 25175 2620 25180 2640
rect 25200 2620 25205 2640
rect 25175 2590 25205 2620
rect 25175 2570 25180 2590
rect 25200 2570 25205 2590
rect 25175 2540 25205 2570
rect 25175 2520 25180 2540
rect 25200 2520 25205 2540
rect 25175 2490 25205 2520
rect 25175 2470 25180 2490
rect 25200 2470 25205 2490
rect 25175 2460 25205 2470
rect 25230 2640 25260 2650
rect 25230 2620 25235 2640
rect 25255 2620 25260 2640
rect 25230 2590 25260 2620
rect 25230 2570 25235 2590
rect 25255 2570 25260 2590
rect 25230 2540 25260 2570
rect 25230 2520 25235 2540
rect 25255 2520 25260 2540
rect 25230 2490 25260 2520
rect 25230 2470 25235 2490
rect 25255 2470 25260 2490
rect 25230 2460 25260 2470
rect 25285 2640 25315 2650
rect 25285 2620 25290 2640
rect 25310 2620 25315 2640
rect 25285 2590 25315 2620
rect 25285 2570 25290 2590
rect 25310 2570 25315 2590
rect 25285 2540 25315 2570
rect 25285 2520 25290 2540
rect 25310 2520 25315 2540
rect 25285 2490 25315 2520
rect 25285 2470 25290 2490
rect 25310 2470 25315 2490
rect 25285 2460 25315 2470
rect 25340 2640 25370 2650
rect 25340 2620 25345 2640
rect 25365 2620 25370 2640
rect 25340 2590 25370 2620
rect 25340 2570 25345 2590
rect 25365 2570 25370 2590
rect 25340 2540 25370 2570
rect 25340 2520 25345 2540
rect 25365 2520 25370 2540
rect 25340 2490 25370 2520
rect 25340 2470 25345 2490
rect 25365 2470 25370 2490
rect 25340 2460 25370 2470
rect 25395 2640 25425 2650
rect 25395 2620 25400 2640
rect 25420 2620 25425 2640
rect 25395 2590 25425 2620
rect 25395 2570 25400 2590
rect 25420 2570 25425 2590
rect 25395 2540 25425 2570
rect 25395 2520 25400 2540
rect 25420 2520 25425 2540
rect 25395 2490 25425 2520
rect 25395 2470 25400 2490
rect 25420 2470 25425 2490
rect 25395 2460 25425 2470
rect 25450 2640 25480 2650
rect 25450 2620 25455 2640
rect 25475 2620 25480 2640
rect 25450 2590 25480 2620
rect 25450 2570 25455 2590
rect 25475 2570 25480 2590
rect 25450 2540 25480 2570
rect 25450 2520 25455 2540
rect 25475 2520 25480 2540
rect 25450 2490 25480 2520
rect 25450 2470 25455 2490
rect 25475 2470 25480 2490
rect 25450 2460 25480 2470
rect 25505 2640 25535 2650
rect 25505 2620 25510 2640
rect 25530 2620 25535 2640
rect 25505 2590 25535 2620
rect 25505 2570 25510 2590
rect 25530 2570 25535 2590
rect 25505 2540 25535 2570
rect 25505 2520 25510 2540
rect 25530 2520 25535 2540
rect 25505 2490 25535 2520
rect 25505 2470 25510 2490
rect 25530 2470 25535 2490
rect 25505 2460 25535 2470
rect 25560 2640 25590 2650
rect 25560 2620 25565 2640
rect 25585 2620 25590 2640
rect 25560 2590 25590 2620
rect 25560 2570 25565 2590
rect 25585 2570 25590 2590
rect 25560 2540 25590 2570
rect 25560 2520 25565 2540
rect 25585 2520 25590 2540
rect 25560 2490 25590 2520
rect 25560 2470 25565 2490
rect 25585 2470 25590 2490
rect 25560 2460 25590 2470
rect 25615 2640 25645 2650
rect 25615 2620 25620 2640
rect 25640 2620 25645 2640
rect 25615 2590 25645 2620
rect 25615 2570 25620 2590
rect 25640 2570 25645 2590
rect 25615 2540 25645 2570
rect 25615 2520 25620 2540
rect 25640 2520 25645 2540
rect 25615 2490 25645 2520
rect 25615 2470 25620 2490
rect 25640 2470 25645 2490
rect 25615 2460 25645 2470
rect 25670 2640 25740 2650
rect 25670 2620 25675 2640
rect 25695 2620 25715 2640
rect 25735 2620 25740 2640
rect 25670 2590 25740 2620
rect 25670 2570 25675 2590
rect 25695 2570 25715 2590
rect 25735 2570 25740 2590
rect 25670 2540 25740 2570
rect 25670 2520 25675 2540
rect 25695 2520 25715 2540
rect 25735 2520 25740 2540
rect 25670 2490 25740 2520
rect 25980 2630 26050 2660
rect 25980 2610 25985 2630
rect 26005 2610 26025 2630
rect 26045 2610 26050 2630
rect 25980 2580 26050 2610
rect 25980 2560 25985 2580
rect 26005 2560 26025 2580
rect 26045 2560 26050 2580
rect 25980 2530 26050 2560
rect 25980 2510 25985 2530
rect 26005 2510 26025 2530
rect 26045 2510 26050 2530
rect 25980 2500 26050 2510
rect 26080 2830 26110 2840
rect 26080 2810 26085 2830
rect 26105 2810 26110 2830
rect 26080 2780 26110 2810
rect 26080 2760 26085 2780
rect 26105 2760 26110 2780
rect 26080 2730 26110 2760
rect 26080 2710 26085 2730
rect 26105 2710 26110 2730
rect 26080 2680 26110 2710
rect 26080 2660 26085 2680
rect 26105 2660 26110 2680
rect 26080 2630 26110 2660
rect 26080 2610 26085 2630
rect 26105 2610 26110 2630
rect 26080 2580 26110 2610
rect 26080 2560 26085 2580
rect 26105 2560 26110 2580
rect 26080 2530 26110 2560
rect 26080 2510 26085 2530
rect 26105 2510 26110 2530
rect 26080 2500 26110 2510
rect 26140 2830 26170 2840
rect 26140 2810 26145 2830
rect 26165 2810 26170 2830
rect 26140 2780 26170 2810
rect 26140 2760 26145 2780
rect 26165 2760 26170 2780
rect 26140 2730 26170 2760
rect 26140 2710 26145 2730
rect 26165 2710 26170 2730
rect 26140 2680 26170 2710
rect 26140 2660 26145 2680
rect 26165 2660 26170 2680
rect 26140 2630 26170 2660
rect 26140 2610 26145 2630
rect 26165 2610 26170 2630
rect 26140 2580 26170 2610
rect 26140 2560 26145 2580
rect 26165 2560 26170 2580
rect 26140 2530 26170 2560
rect 26140 2510 26145 2530
rect 26165 2510 26170 2530
rect 26140 2500 26170 2510
rect 26200 2830 26230 2840
rect 26200 2810 26205 2830
rect 26225 2810 26230 2830
rect 26200 2780 26230 2810
rect 26200 2760 26205 2780
rect 26225 2760 26230 2780
rect 26200 2730 26230 2760
rect 26200 2710 26205 2730
rect 26225 2710 26230 2730
rect 26200 2680 26230 2710
rect 26200 2660 26205 2680
rect 26225 2660 26230 2680
rect 26200 2630 26230 2660
rect 26200 2610 26205 2630
rect 26225 2610 26230 2630
rect 26200 2580 26230 2610
rect 26200 2560 26205 2580
rect 26225 2560 26230 2580
rect 26200 2530 26230 2560
rect 26200 2510 26205 2530
rect 26225 2510 26230 2530
rect 26200 2500 26230 2510
rect 26260 2830 26290 2840
rect 26260 2810 26265 2830
rect 26285 2810 26290 2830
rect 26260 2780 26290 2810
rect 26260 2760 26265 2780
rect 26285 2760 26290 2780
rect 26260 2730 26290 2760
rect 26260 2710 26265 2730
rect 26285 2710 26290 2730
rect 26260 2680 26290 2710
rect 26260 2660 26265 2680
rect 26285 2660 26290 2680
rect 26260 2630 26290 2660
rect 26260 2610 26265 2630
rect 26285 2610 26290 2630
rect 26260 2580 26290 2610
rect 26260 2560 26265 2580
rect 26285 2560 26290 2580
rect 26260 2530 26290 2560
rect 26260 2510 26265 2530
rect 26285 2510 26290 2530
rect 26260 2500 26290 2510
rect 26320 2830 26350 2840
rect 26320 2810 26325 2830
rect 26345 2810 26350 2830
rect 26320 2780 26350 2810
rect 26320 2760 26325 2780
rect 26345 2760 26350 2780
rect 26320 2730 26350 2760
rect 26320 2710 26325 2730
rect 26345 2710 26350 2730
rect 26320 2680 26350 2710
rect 26320 2660 26325 2680
rect 26345 2660 26350 2680
rect 26320 2630 26350 2660
rect 26320 2610 26325 2630
rect 26345 2610 26350 2630
rect 26320 2580 26350 2610
rect 26320 2560 26325 2580
rect 26345 2560 26350 2580
rect 26320 2530 26350 2560
rect 26320 2510 26325 2530
rect 26345 2510 26350 2530
rect 26320 2500 26350 2510
rect 26380 2830 26410 2840
rect 26380 2810 26385 2830
rect 26405 2810 26410 2830
rect 26380 2780 26410 2810
rect 26380 2760 26385 2780
rect 26405 2760 26410 2780
rect 26380 2730 26410 2760
rect 26380 2710 26385 2730
rect 26405 2710 26410 2730
rect 26380 2680 26410 2710
rect 26380 2660 26385 2680
rect 26405 2660 26410 2680
rect 26380 2630 26410 2660
rect 26380 2610 26385 2630
rect 26405 2610 26410 2630
rect 26380 2580 26410 2610
rect 26380 2560 26385 2580
rect 26405 2560 26410 2580
rect 26380 2530 26410 2560
rect 26380 2510 26385 2530
rect 26405 2510 26410 2530
rect 26380 2500 26410 2510
rect 26440 2830 26470 2840
rect 26440 2810 26445 2830
rect 26465 2810 26470 2830
rect 26440 2780 26470 2810
rect 26440 2760 26445 2780
rect 26465 2760 26470 2780
rect 26440 2730 26470 2760
rect 26440 2710 26445 2730
rect 26465 2710 26470 2730
rect 26440 2680 26470 2710
rect 26440 2660 26445 2680
rect 26465 2660 26470 2680
rect 26440 2630 26470 2660
rect 26440 2610 26445 2630
rect 26465 2610 26470 2630
rect 26440 2580 26470 2610
rect 26440 2560 26445 2580
rect 26465 2560 26470 2580
rect 26440 2530 26470 2560
rect 26440 2510 26445 2530
rect 26465 2510 26470 2530
rect 26440 2500 26470 2510
rect 26500 2830 26530 2840
rect 26500 2810 26505 2830
rect 26525 2810 26530 2830
rect 26500 2780 26530 2810
rect 26500 2760 26505 2780
rect 26525 2760 26530 2780
rect 26500 2730 26530 2760
rect 26500 2710 26505 2730
rect 26525 2710 26530 2730
rect 26500 2680 26530 2710
rect 26500 2660 26505 2680
rect 26525 2660 26530 2680
rect 26500 2630 26530 2660
rect 26500 2610 26505 2630
rect 26525 2610 26530 2630
rect 26500 2580 26530 2610
rect 26500 2560 26505 2580
rect 26525 2560 26530 2580
rect 26500 2530 26530 2560
rect 26500 2510 26505 2530
rect 26525 2510 26530 2530
rect 26500 2500 26530 2510
rect 26560 2830 26590 2840
rect 26560 2810 26565 2830
rect 26585 2810 26590 2830
rect 26560 2780 26590 2810
rect 26560 2760 26565 2780
rect 26585 2760 26590 2780
rect 26560 2730 26590 2760
rect 26560 2710 26565 2730
rect 26585 2710 26590 2730
rect 26560 2680 26590 2710
rect 26560 2660 26565 2680
rect 26585 2660 26590 2680
rect 26560 2630 26590 2660
rect 26560 2610 26565 2630
rect 26585 2610 26590 2630
rect 26560 2580 26590 2610
rect 26560 2560 26565 2580
rect 26585 2560 26590 2580
rect 26560 2530 26590 2560
rect 26560 2510 26565 2530
rect 26585 2510 26590 2530
rect 26560 2500 26590 2510
rect 26620 2830 26650 2840
rect 26620 2810 26625 2830
rect 26645 2810 26650 2830
rect 26620 2780 26650 2810
rect 26620 2760 26625 2780
rect 26645 2760 26650 2780
rect 26620 2730 26650 2760
rect 26620 2710 26625 2730
rect 26645 2710 26650 2730
rect 26620 2680 26650 2710
rect 26620 2660 26625 2680
rect 26645 2660 26650 2680
rect 26620 2630 26650 2660
rect 26620 2610 26625 2630
rect 26645 2610 26650 2630
rect 26620 2580 26650 2610
rect 26620 2560 26625 2580
rect 26645 2560 26650 2580
rect 26620 2530 26650 2560
rect 26620 2510 26625 2530
rect 26645 2510 26650 2530
rect 26620 2500 26650 2510
rect 26680 2830 26710 2840
rect 26680 2810 26685 2830
rect 26705 2810 26710 2830
rect 26680 2780 26710 2810
rect 26680 2760 26685 2780
rect 26705 2760 26710 2780
rect 26680 2730 26710 2760
rect 26680 2710 26685 2730
rect 26705 2710 26710 2730
rect 26680 2680 26710 2710
rect 26680 2660 26685 2680
rect 26705 2660 26710 2680
rect 26680 2630 26710 2660
rect 26680 2610 26685 2630
rect 26705 2610 26710 2630
rect 26680 2580 26710 2610
rect 26680 2560 26685 2580
rect 26705 2560 26710 2580
rect 26680 2530 26710 2560
rect 26680 2510 26685 2530
rect 26705 2510 26710 2530
rect 26680 2500 26710 2510
rect 26740 2830 26810 2840
rect 26740 2810 26745 2830
rect 26765 2810 26785 2830
rect 26805 2810 26810 2830
rect 26740 2780 26810 2810
rect 26740 2760 26745 2780
rect 26765 2760 26785 2780
rect 26805 2760 26810 2780
rect 26740 2730 26810 2760
rect 26740 2710 26745 2730
rect 26765 2710 26785 2730
rect 26805 2710 26810 2730
rect 26740 2680 26810 2710
rect 26740 2660 26745 2680
rect 26765 2660 26785 2680
rect 26805 2660 26810 2680
rect 26740 2630 26810 2660
rect 26740 2610 26745 2630
rect 26765 2610 26785 2630
rect 26805 2610 26810 2630
rect 26740 2580 26810 2610
rect 26740 2560 26745 2580
rect 26765 2560 26785 2580
rect 26805 2560 26810 2580
rect 26740 2530 26810 2560
rect 26740 2510 26745 2530
rect 26765 2510 26785 2530
rect 26805 2510 26810 2530
rect 26740 2500 26810 2510
rect 26985 2710 27005 2920
rect 27155 2890 27195 2900
rect 27155 2870 27165 2890
rect 27185 2870 27195 2890
rect 27155 2860 27195 2870
rect 27275 2890 27315 2900
rect 27275 2870 27285 2890
rect 27305 2870 27315 2890
rect 27275 2860 27315 2870
rect 27395 2890 27435 2900
rect 27395 2870 27405 2890
rect 27425 2870 27435 2890
rect 27395 2860 27435 2870
rect 27515 2890 27555 2900
rect 27515 2870 27525 2890
rect 27545 2870 27555 2890
rect 27515 2860 27555 2870
rect 27635 2890 27675 2900
rect 27635 2870 27645 2890
rect 27665 2870 27675 2890
rect 27635 2860 27675 2870
rect 27165 2840 27185 2860
rect 27285 2840 27305 2860
rect 27405 2840 27425 2860
rect 27525 2840 27545 2860
rect 27645 2840 27665 2860
rect 25670 2470 25675 2490
rect 25695 2470 25715 2490
rect 25735 2470 25740 2490
rect 26085 2480 26105 2500
rect 26205 2480 26225 2500
rect 26325 2480 26345 2500
rect 26445 2480 26465 2500
rect 26565 2480 26585 2500
rect 26685 2480 26705 2500
rect 25670 2460 25740 2470
rect 26075 2470 26115 2480
rect 24975 2440 24995 2460
rect 25125 2440 25145 2460
rect 25235 2440 25255 2460
rect 25345 2440 25365 2460
rect 25455 2440 25475 2460
rect 25565 2440 25585 2460
rect 25715 2440 25735 2460
rect 26075 2450 26085 2470
rect 26105 2450 26115 2470
rect 26075 2440 26115 2450
rect 26195 2470 26235 2480
rect 26195 2450 26205 2470
rect 26225 2450 26235 2470
rect 26195 2440 26235 2450
rect 26315 2470 26355 2480
rect 26315 2450 26325 2470
rect 26345 2450 26355 2470
rect 26315 2440 26355 2450
rect 26378 2470 26412 2480
rect 26378 2450 26386 2470
rect 26404 2450 26412 2470
rect 26378 2440 26412 2450
rect 26435 2470 26475 2480
rect 26435 2450 26445 2470
rect 26465 2450 26475 2470
rect 26435 2440 26475 2450
rect 26555 2470 26595 2480
rect 26555 2450 26565 2470
rect 26585 2450 26595 2470
rect 26555 2440 26595 2450
rect 26675 2470 26715 2480
rect 26675 2450 26685 2470
rect 26705 2450 26715 2470
rect 26675 2440 26715 2450
rect 24965 2430 25005 2440
rect 24965 2410 24975 2430
rect 24995 2410 25005 2430
rect 24965 2400 25005 2410
rect 25115 2430 25155 2440
rect 25115 2410 25125 2430
rect 25145 2410 25155 2430
rect 25115 2400 25155 2410
rect 25225 2430 25265 2440
rect 25225 2410 25235 2430
rect 25255 2410 25265 2430
rect 25225 2400 25265 2410
rect 25335 2430 25375 2440
rect 25335 2410 25345 2430
rect 25365 2410 25375 2430
rect 25335 2400 25375 2410
rect 25445 2430 25485 2440
rect 25445 2410 25455 2430
rect 25475 2410 25485 2430
rect 25445 2400 25485 2410
rect 25555 2430 25595 2440
rect 25555 2410 25565 2430
rect 25585 2410 25595 2430
rect 25555 2400 25595 2410
rect 25705 2430 25745 2440
rect 25705 2410 25715 2430
rect 25735 2410 25745 2430
rect 25705 2400 25745 2410
rect 26985 2420 27005 2630
rect 27040 2830 27070 2840
rect 27040 2810 27045 2830
rect 27065 2810 27070 2830
rect 27040 2780 27070 2810
rect 27040 2760 27045 2780
rect 27065 2760 27070 2780
rect 27040 2730 27070 2760
rect 27040 2710 27045 2730
rect 27065 2710 27070 2730
rect 27040 2680 27070 2710
rect 27040 2660 27045 2680
rect 27065 2660 27070 2680
rect 27040 2630 27070 2660
rect 27040 2610 27045 2630
rect 27065 2610 27070 2630
rect 27040 2580 27070 2610
rect 27040 2560 27045 2580
rect 27065 2560 27070 2580
rect 27040 2530 27070 2560
rect 27040 2510 27045 2530
rect 27065 2510 27070 2530
rect 27040 2500 27070 2510
rect 27100 2830 27130 2840
rect 27100 2810 27105 2830
rect 27125 2810 27130 2830
rect 27100 2780 27130 2810
rect 27100 2760 27105 2780
rect 27125 2760 27130 2780
rect 27100 2730 27130 2760
rect 27100 2710 27105 2730
rect 27125 2710 27130 2730
rect 27100 2680 27130 2710
rect 27100 2660 27105 2680
rect 27125 2660 27130 2680
rect 27100 2630 27130 2660
rect 27100 2610 27105 2630
rect 27125 2610 27130 2630
rect 27100 2580 27130 2610
rect 27100 2560 27105 2580
rect 27125 2560 27130 2580
rect 27100 2530 27130 2560
rect 27100 2510 27105 2530
rect 27125 2510 27130 2530
rect 27100 2500 27130 2510
rect 27160 2830 27190 2840
rect 27160 2810 27165 2830
rect 27185 2810 27190 2830
rect 27160 2780 27190 2810
rect 27160 2760 27165 2780
rect 27185 2760 27190 2780
rect 27160 2730 27190 2760
rect 27160 2710 27165 2730
rect 27185 2710 27190 2730
rect 27160 2680 27190 2710
rect 27160 2660 27165 2680
rect 27185 2660 27190 2680
rect 27160 2630 27190 2660
rect 27160 2610 27165 2630
rect 27185 2610 27190 2630
rect 27160 2580 27190 2610
rect 27160 2560 27165 2580
rect 27185 2560 27190 2580
rect 27160 2530 27190 2560
rect 27160 2510 27165 2530
rect 27185 2510 27190 2530
rect 27160 2500 27190 2510
rect 27220 2830 27250 2840
rect 27220 2810 27225 2830
rect 27245 2810 27250 2830
rect 27220 2780 27250 2810
rect 27220 2760 27225 2780
rect 27245 2760 27250 2780
rect 27220 2730 27250 2760
rect 27220 2710 27225 2730
rect 27245 2710 27250 2730
rect 27220 2680 27250 2710
rect 27220 2660 27225 2680
rect 27245 2660 27250 2680
rect 27220 2630 27250 2660
rect 27220 2610 27225 2630
rect 27245 2610 27250 2630
rect 27220 2580 27250 2610
rect 27220 2560 27225 2580
rect 27245 2560 27250 2580
rect 27220 2530 27250 2560
rect 27220 2510 27225 2530
rect 27245 2510 27250 2530
rect 27220 2500 27250 2510
rect 27280 2830 27310 2840
rect 27280 2810 27285 2830
rect 27305 2810 27310 2830
rect 27280 2780 27310 2810
rect 27280 2760 27285 2780
rect 27305 2760 27310 2780
rect 27280 2730 27310 2760
rect 27280 2710 27285 2730
rect 27305 2710 27310 2730
rect 27280 2680 27310 2710
rect 27280 2660 27285 2680
rect 27305 2660 27310 2680
rect 27280 2630 27310 2660
rect 27280 2610 27285 2630
rect 27305 2610 27310 2630
rect 27280 2580 27310 2610
rect 27280 2560 27285 2580
rect 27305 2560 27310 2580
rect 27280 2530 27310 2560
rect 27280 2510 27285 2530
rect 27305 2510 27310 2530
rect 27280 2500 27310 2510
rect 27340 2830 27370 2840
rect 27340 2810 27345 2830
rect 27365 2810 27370 2830
rect 27340 2780 27370 2810
rect 27340 2760 27345 2780
rect 27365 2760 27370 2780
rect 27340 2730 27370 2760
rect 27340 2710 27345 2730
rect 27365 2710 27370 2730
rect 27340 2680 27370 2710
rect 27340 2660 27345 2680
rect 27365 2660 27370 2680
rect 27340 2630 27370 2660
rect 27340 2610 27345 2630
rect 27365 2610 27370 2630
rect 27340 2580 27370 2610
rect 27340 2560 27345 2580
rect 27365 2560 27370 2580
rect 27340 2530 27370 2560
rect 27340 2510 27345 2530
rect 27365 2510 27370 2530
rect 27340 2500 27370 2510
rect 27400 2830 27430 2840
rect 27400 2810 27405 2830
rect 27425 2810 27430 2830
rect 27400 2780 27430 2810
rect 27400 2760 27405 2780
rect 27425 2760 27430 2780
rect 27400 2730 27430 2760
rect 27400 2710 27405 2730
rect 27425 2710 27430 2730
rect 27400 2680 27430 2710
rect 27400 2660 27405 2680
rect 27425 2660 27430 2680
rect 27400 2630 27430 2660
rect 27400 2610 27405 2630
rect 27425 2610 27430 2630
rect 27400 2580 27430 2610
rect 27400 2560 27405 2580
rect 27425 2560 27430 2580
rect 27400 2530 27430 2560
rect 27400 2510 27405 2530
rect 27425 2510 27430 2530
rect 27400 2500 27430 2510
rect 27460 2830 27490 2840
rect 27460 2810 27465 2830
rect 27485 2810 27490 2830
rect 27460 2780 27490 2810
rect 27460 2760 27465 2780
rect 27485 2760 27490 2780
rect 27460 2730 27490 2760
rect 27460 2710 27465 2730
rect 27485 2710 27490 2730
rect 27460 2680 27490 2710
rect 27460 2660 27465 2680
rect 27485 2660 27490 2680
rect 27460 2630 27490 2660
rect 27460 2610 27465 2630
rect 27485 2610 27490 2630
rect 27460 2580 27490 2610
rect 27460 2560 27465 2580
rect 27485 2560 27490 2580
rect 27460 2530 27490 2560
rect 27460 2510 27465 2530
rect 27485 2510 27490 2530
rect 27460 2500 27490 2510
rect 27520 2830 27550 2840
rect 27520 2810 27525 2830
rect 27545 2810 27550 2830
rect 27520 2780 27550 2810
rect 27520 2760 27525 2780
rect 27545 2760 27550 2780
rect 27520 2730 27550 2760
rect 27520 2710 27525 2730
rect 27545 2710 27550 2730
rect 27520 2680 27550 2710
rect 27520 2660 27525 2680
rect 27545 2660 27550 2680
rect 27520 2630 27550 2660
rect 27520 2610 27525 2630
rect 27545 2610 27550 2630
rect 27520 2580 27550 2610
rect 27520 2560 27525 2580
rect 27545 2560 27550 2580
rect 27520 2530 27550 2560
rect 27520 2510 27525 2530
rect 27545 2510 27550 2530
rect 27520 2500 27550 2510
rect 27580 2830 27610 2840
rect 27580 2810 27585 2830
rect 27605 2810 27610 2830
rect 27580 2780 27610 2810
rect 27580 2760 27585 2780
rect 27605 2760 27610 2780
rect 27580 2730 27610 2760
rect 27580 2710 27585 2730
rect 27605 2710 27610 2730
rect 27580 2680 27610 2710
rect 27580 2660 27585 2680
rect 27605 2660 27610 2680
rect 27580 2630 27610 2660
rect 27580 2610 27585 2630
rect 27605 2610 27610 2630
rect 27580 2580 27610 2610
rect 27580 2560 27585 2580
rect 27605 2560 27610 2580
rect 27580 2530 27610 2560
rect 27580 2510 27585 2530
rect 27605 2510 27610 2530
rect 27580 2500 27610 2510
rect 27640 2830 27670 2840
rect 27640 2810 27645 2830
rect 27665 2810 27670 2830
rect 27640 2780 27670 2810
rect 27640 2760 27645 2780
rect 27665 2760 27670 2780
rect 27640 2730 27670 2760
rect 27640 2710 27645 2730
rect 27665 2710 27670 2730
rect 27640 2680 27670 2710
rect 27640 2660 27645 2680
rect 27665 2660 27670 2680
rect 27640 2630 27670 2660
rect 27640 2610 27645 2630
rect 27665 2610 27670 2630
rect 27640 2580 27670 2610
rect 27640 2560 27645 2580
rect 27665 2560 27670 2580
rect 27640 2530 27670 2560
rect 27640 2510 27645 2530
rect 27665 2510 27670 2530
rect 27640 2500 27670 2510
rect 27700 2830 27730 2840
rect 27700 2810 27705 2830
rect 27725 2810 27730 2830
rect 27700 2780 27730 2810
rect 27700 2760 27705 2780
rect 27725 2760 27730 2780
rect 27700 2730 27730 2760
rect 27700 2710 27705 2730
rect 27725 2710 27730 2730
rect 27700 2680 27730 2710
rect 27700 2660 27705 2680
rect 27725 2660 27730 2680
rect 27700 2630 27730 2660
rect 27700 2610 27705 2630
rect 27725 2610 27730 2630
rect 27700 2580 27730 2610
rect 27700 2560 27705 2580
rect 27725 2560 27730 2580
rect 27700 2530 27730 2560
rect 27700 2510 27705 2530
rect 27725 2510 27730 2530
rect 27700 2500 27730 2510
rect 27760 2830 27790 2840
rect 27760 2810 27765 2830
rect 27785 2810 27790 2830
rect 27760 2780 27790 2810
rect 27760 2760 27765 2780
rect 27785 2760 27790 2780
rect 27760 2730 27790 2760
rect 27760 2710 27765 2730
rect 27785 2710 27790 2730
rect 27760 2680 27790 2710
rect 27760 2660 27765 2680
rect 27785 2660 27790 2680
rect 27760 2630 27790 2660
rect 27760 2610 27765 2630
rect 27785 2610 27790 2630
rect 27760 2580 27790 2610
rect 27760 2560 27765 2580
rect 27785 2560 27790 2580
rect 27760 2530 27790 2560
rect 27760 2510 27765 2530
rect 27785 2510 27790 2530
rect 27760 2500 27790 2510
rect 27825 2710 27845 2920
rect 27105 2480 27125 2500
rect 27225 2480 27245 2500
rect 27345 2480 27365 2500
rect 27465 2480 27485 2500
rect 27585 2480 27605 2500
rect 27705 2480 27725 2500
rect 27095 2470 27135 2480
rect 27095 2450 27105 2470
rect 27125 2450 27135 2470
rect 27095 2440 27135 2450
rect 27215 2470 27255 2480
rect 27215 2450 27225 2470
rect 27245 2450 27255 2470
rect 27215 2440 27255 2450
rect 27335 2470 27375 2480
rect 27335 2450 27345 2470
rect 27365 2450 27375 2470
rect 27335 2440 27375 2450
rect 27398 2470 27432 2480
rect 27398 2450 27406 2470
rect 27424 2450 27432 2470
rect 27398 2440 27432 2450
rect 27455 2470 27495 2480
rect 27455 2450 27465 2470
rect 27485 2450 27495 2470
rect 27455 2440 27495 2450
rect 27575 2470 27615 2480
rect 27575 2450 27585 2470
rect 27605 2450 27615 2470
rect 27575 2440 27615 2450
rect 27695 2470 27735 2480
rect 27695 2450 27705 2470
rect 27725 2450 27735 2470
rect 27695 2440 27735 2450
rect 27825 2420 27845 2630
rect 26985 2400 27375 2420
rect 27455 2400 27845 2420
rect 28095 2780 28455 2800
rect 28535 2780 28895 2800
rect 28095 2645 28115 2780
rect 28200 2750 28240 2760
rect 28200 2730 28210 2750
rect 28230 2730 28240 2750
rect 28200 2720 28240 2730
rect 28310 2750 28350 2760
rect 28310 2730 28320 2750
rect 28340 2730 28350 2750
rect 28310 2720 28350 2730
rect 28420 2750 28460 2760
rect 28420 2730 28430 2750
rect 28450 2730 28460 2750
rect 28420 2720 28460 2730
rect 28530 2750 28570 2760
rect 28530 2730 28540 2750
rect 28560 2730 28570 2750
rect 28530 2720 28570 2730
rect 28640 2750 28680 2760
rect 28640 2730 28650 2750
rect 28670 2730 28680 2750
rect 28640 2720 28680 2730
rect 28750 2750 28790 2760
rect 28750 2730 28760 2750
rect 28780 2730 28790 2750
rect 28750 2720 28790 2730
rect 28210 2700 28230 2720
rect 28320 2700 28340 2720
rect 28430 2700 28450 2720
rect 28540 2700 28560 2720
rect 28650 2700 28670 2720
rect 28760 2700 28780 2720
rect 28095 2430 28115 2565
rect 28150 2690 28180 2700
rect 28150 2670 28155 2690
rect 28175 2670 28180 2690
rect 28150 2640 28180 2670
rect 28150 2620 28155 2640
rect 28175 2620 28180 2640
rect 28150 2590 28180 2620
rect 28150 2570 28155 2590
rect 28175 2570 28180 2590
rect 28150 2540 28180 2570
rect 28150 2520 28155 2540
rect 28175 2520 28180 2540
rect 28150 2510 28180 2520
rect 28205 2690 28235 2700
rect 28205 2670 28210 2690
rect 28230 2670 28235 2690
rect 28205 2640 28235 2670
rect 28205 2620 28210 2640
rect 28230 2620 28235 2640
rect 28205 2590 28235 2620
rect 28205 2570 28210 2590
rect 28230 2570 28235 2590
rect 28205 2540 28235 2570
rect 28205 2520 28210 2540
rect 28230 2520 28235 2540
rect 28205 2510 28235 2520
rect 28260 2690 28290 2700
rect 28260 2670 28265 2690
rect 28285 2670 28290 2690
rect 28260 2640 28290 2670
rect 28260 2620 28265 2640
rect 28285 2620 28290 2640
rect 28260 2590 28290 2620
rect 28260 2570 28265 2590
rect 28285 2570 28290 2590
rect 28260 2540 28290 2570
rect 28260 2520 28265 2540
rect 28285 2520 28290 2540
rect 28260 2510 28290 2520
rect 28315 2690 28345 2700
rect 28315 2670 28320 2690
rect 28340 2670 28345 2690
rect 28315 2640 28345 2670
rect 28315 2620 28320 2640
rect 28340 2620 28345 2640
rect 28315 2590 28345 2620
rect 28315 2570 28320 2590
rect 28340 2570 28345 2590
rect 28315 2540 28345 2570
rect 28315 2520 28320 2540
rect 28340 2520 28345 2540
rect 28315 2510 28345 2520
rect 28370 2690 28400 2700
rect 28370 2670 28375 2690
rect 28395 2670 28400 2690
rect 28370 2640 28400 2670
rect 28370 2620 28375 2640
rect 28395 2620 28400 2640
rect 28370 2590 28400 2620
rect 28370 2570 28375 2590
rect 28395 2570 28400 2590
rect 28370 2540 28400 2570
rect 28370 2520 28375 2540
rect 28395 2520 28400 2540
rect 28370 2510 28400 2520
rect 28425 2690 28455 2700
rect 28425 2670 28430 2690
rect 28450 2670 28455 2690
rect 28425 2640 28455 2670
rect 28425 2620 28430 2640
rect 28450 2620 28455 2640
rect 28425 2590 28455 2620
rect 28425 2570 28430 2590
rect 28450 2570 28455 2590
rect 28425 2540 28455 2570
rect 28425 2520 28430 2540
rect 28450 2520 28455 2540
rect 28425 2510 28455 2520
rect 28480 2690 28510 2700
rect 28480 2670 28485 2690
rect 28505 2670 28510 2690
rect 28480 2640 28510 2670
rect 28480 2620 28485 2640
rect 28505 2620 28510 2640
rect 28480 2590 28510 2620
rect 28480 2570 28485 2590
rect 28505 2570 28510 2590
rect 28480 2540 28510 2570
rect 28480 2520 28485 2540
rect 28505 2520 28510 2540
rect 28480 2510 28510 2520
rect 28535 2690 28565 2700
rect 28535 2670 28540 2690
rect 28560 2670 28565 2690
rect 28535 2640 28565 2670
rect 28535 2620 28540 2640
rect 28560 2620 28565 2640
rect 28535 2590 28565 2620
rect 28535 2570 28540 2590
rect 28560 2570 28565 2590
rect 28535 2540 28565 2570
rect 28535 2520 28540 2540
rect 28560 2520 28565 2540
rect 28535 2510 28565 2520
rect 28590 2690 28620 2700
rect 28590 2670 28595 2690
rect 28615 2670 28620 2690
rect 28590 2640 28620 2670
rect 28590 2620 28595 2640
rect 28615 2620 28620 2640
rect 28590 2590 28620 2620
rect 28590 2570 28595 2590
rect 28615 2570 28620 2590
rect 28590 2540 28620 2570
rect 28590 2520 28595 2540
rect 28615 2520 28620 2540
rect 28590 2510 28620 2520
rect 28645 2690 28675 2700
rect 28645 2670 28650 2690
rect 28670 2670 28675 2690
rect 28645 2640 28675 2670
rect 28645 2620 28650 2640
rect 28670 2620 28675 2640
rect 28645 2590 28675 2620
rect 28645 2570 28650 2590
rect 28670 2570 28675 2590
rect 28645 2540 28675 2570
rect 28645 2520 28650 2540
rect 28670 2520 28675 2540
rect 28645 2510 28675 2520
rect 28700 2690 28730 2700
rect 28700 2670 28705 2690
rect 28725 2670 28730 2690
rect 28700 2640 28730 2670
rect 28700 2620 28705 2640
rect 28725 2620 28730 2640
rect 28700 2590 28730 2620
rect 28700 2570 28705 2590
rect 28725 2570 28730 2590
rect 28700 2540 28730 2570
rect 28700 2520 28705 2540
rect 28725 2520 28730 2540
rect 28700 2510 28730 2520
rect 28755 2690 28785 2700
rect 28755 2670 28760 2690
rect 28780 2670 28785 2690
rect 28755 2640 28785 2670
rect 28755 2620 28760 2640
rect 28780 2620 28785 2640
rect 28755 2590 28785 2620
rect 28755 2570 28760 2590
rect 28780 2570 28785 2590
rect 28755 2540 28785 2570
rect 28755 2520 28760 2540
rect 28780 2520 28785 2540
rect 28755 2510 28785 2520
rect 28810 2690 28840 2700
rect 28810 2670 28815 2690
rect 28835 2670 28840 2690
rect 28810 2640 28840 2670
rect 28810 2620 28815 2640
rect 28835 2620 28840 2640
rect 28810 2590 28840 2620
rect 28810 2570 28815 2590
rect 28835 2570 28840 2590
rect 28810 2540 28840 2570
rect 28810 2520 28815 2540
rect 28835 2520 28840 2540
rect 28810 2510 28840 2520
rect 28875 2645 28895 2780
rect 28265 2490 28285 2510
rect 28375 2490 28395 2510
rect 28485 2490 28505 2510
rect 28595 2490 28615 2510
rect 28705 2490 28725 2510
rect 28255 2480 28295 2490
rect 28255 2460 28265 2480
rect 28285 2460 28295 2480
rect 28255 2450 28295 2460
rect 28313 2480 28347 2490
rect 28313 2460 28321 2480
rect 28339 2460 28347 2480
rect 28313 2450 28347 2460
rect 28365 2480 28405 2490
rect 28365 2460 28375 2480
rect 28395 2460 28405 2480
rect 28365 2450 28405 2460
rect 28475 2480 28515 2490
rect 28475 2460 28485 2480
rect 28505 2460 28515 2480
rect 28475 2450 28515 2460
rect 28585 2480 28625 2490
rect 28585 2460 28595 2480
rect 28615 2460 28625 2480
rect 28585 2450 28625 2460
rect 28695 2480 28735 2490
rect 28695 2460 28705 2480
rect 28725 2460 28735 2480
rect 28695 2450 28735 2460
rect 28875 2430 28895 2565
rect 28095 2410 28455 2430
rect 28535 2410 28895 2430
rect 28995 2665 29135 2685
rect 29215 2665 29350 2685
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 15585 2370 15625 2380
rect 15585 2350 15595 2370
rect 15615 2350 15625 2370
rect 15585 2340 15625 2350
rect 18225 2370 18265 2380
rect 18225 2350 18235 2370
rect 18255 2350 18265 2370
rect 18225 2340 18265 2350
rect 25585 2370 25625 2380
rect 25585 2350 25595 2370
rect 25615 2350 25625 2370
rect 25585 2340 25625 2350
rect 3625 2330 3665 2340
rect 3625 2310 3635 2330
rect 3655 2310 3665 2330
rect 3625 2300 3665 2310
rect 4345 2330 4385 2340
rect 4345 2310 4355 2330
rect 4375 2310 4385 2330
rect 28095 2320 28455 2340
rect 28535 2320 28895 2340
rect 4345 2300 4385 2310
rect 14965 2310 15005 2320
rect 2740 2260 2770 2290
rect 3445 2285 3485 2295
rect 3445 2265 3455 2285
rect 3475 2265 3485 2285
rect 3445 2255 3485 2265
rect 4525 2285 4565 2295
rect 14965 2290 14975 2310
rect 14995 2290 15005 2310
rect 4525 2265 4535 2285
rect 4555 2265 4565 2285
rect 4525 2255 4565 2265
rect 5275 2260 5305 2290
rect 14965 2280 15005 2290
rect 15115 2310 15155 2320
rect 15115 2290 15125 2310
rect 15145 2290 15155 2310
rect 15115 2280 15155 2290
rect 15225 2310 15265 2320
rect 15225 2290 15235 2310
rect 15255 2290 15265 2310
rect 15225 2280 15265 2290
rect 15335 2310 15375 2320
rect 15335 2290 15345 2310
rect 15365 2290 15375 2310
rect 15335 2280 15375 2290
rect 15445 2310 15485 2320
rect 15445 2290 15455 2310
rect 15475 2290 15485 2310
rect 15445 2280 15485 2290
rect 15555 2310 15595 2320
rect 15555 2290 15565 2310
rect 15585 2290 15595 2310
rect 15555 2280 15595 2290
rect 15705 2310 15745 2320
rect 15705 2290 15715 2310
rect 15735 2290 15745 2310
rect 15705 2280 15745 2290
rect 18105 2310 18145 2320
rect 18105 2290 18115 2310
rect 18135 2290 18145 2310
rect 18105 2280 18145 2290
rect 18255 2310 18295 2320
rect 18255 2290 18265 2310
rect 18285 2290 18295 2310
rect 18255 2280 18295 2290
rect 18365 2310 18405 2320
rect 18365 2290 18375 2310
rect 18395 2290 18405 2310
rect 18365 2280 18405 2290
rect 18475 2310 18515 2320
rect 18475 2290 18485 2310
rect 18505 2290 18515 2310
rect 18475 2280 18515 2290
rect 18585 2310 18625 2320
rect 18585 2290 18595 2310
rect 18615 2290 18625 2310
rect 18585 2280 18625 2290
rect 18695 2310 18735 2320
rect 18695 2290 18705 2310
rect 18725 2290 18735 2310
rect 18695 2280 18735 2290
rect 18845 2310 18885 2320
rect 18845 2290 18855 2310
rect 18875 2290 18885 2310
rect 18845 2280 18885 2290
rect 24965 2310 25005 2320
rect 24965 2290 24975 2310
rect 24995 2290 25005 2310
rect 24965 2280 25005 2290
rect 25115 2310 25155 2320
rect 25115 2290 25125 2310
rect 25145 2290 25155 2310
rect 25115 2280 25155 2290
rect 25225 2310 25265 2320
rect 25225 2290 25235 2310
rect 25255 2290 25265 2310
rect 25225 2280 25265 2290
rect 25335 2310 25375 2320
rect 25335 2290 25345 2310
rect 25365 2290 25375 2310
rect 25335 2280 25375 2290
rect 25445 2310 25485 2320
rect 25445 2290 25455 2310
rect 25475 2290 25485 2310
rect 25445 2280 25485 2290
rect 25555 2310 25595 2320
rect 25555 2290 25565 2310
rect 25585 2290 25595 2310
rect 25555 2280 25595 2290
rect 25705 2310 25745 2320
rect 25705 2290 25715 2310
rect 25735 2290 25745 2310
rect 25705 2280 25745 2290
rect 14975 2260 14995 2280
rect 15125 2260 15145 2280
rect 15235 2260 15255 2280
rect 15345 2260 15365 2280
rect 15455 2260 15475 2280
rect 15565 2260 15585 2280
rect 15715 2260 15735 2280
rect 18115 2260 18135 2280
rect 18265 2260 18285 2280
rect 18375 2260 18395 2280
rect 18485 2260 18505 2280
rect 18595 2260 18615 2280
rect 18705 2260 18725 2280
rect 18855 2260 18875 2280
rect 24975 2260 24995 2280
rect 25125 2260 25145 2280
rect 25235 2260 25255 2280
rect 25345 2260 25365 2280
rect 25455 2260 25475 2280
rect 25565 2260 25585 2280
rect 25715 2260 25735 2280
rect 14970 2250 15040 2260
rect 2430 2215 2460 2245
rect 3810 2215 3840 2245
rect 14970 2230 14975 2250
rect 14995 2230 15015 2250
rect 15035 2230 15040 2250
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3630 2120 3660 2150
rect 4090 2115 4120 2145
rect 5320 2115 5350 2145
rect 2745 2090 2785 2100
rect 2745 2070 2755 2090
rect 2775 2070 2785 2090
rect 2745 2060 2785 2070
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 3985 2090 4025 2100
rect 3985 2070 3995 2090
rect 4015 2070 4025 2090
rect 3985 2060 4025 2070
rect 4145 2090 4185 2100
rect 4145 2070 4155 2090
rect 4175 2070 4185 2090
rect 4145 2060 4185 2070
rect 4265 2090 4305 2100
rect 4265 2070 4275 2090
rect 4295 2070 4305 2090
rect 4265 2060 4305 2070
rect 4385 2090 4425 2100
rect 4385 2070 4395 2090
rect 4415 2070 4425 2090
rect 4385 2060 4425 2070
rect 4505 2090 4545 2100
rect 4505 2070 4515 2090
rect 4535 2070 4545 2090
rect 4505 2060 4545 2070
rect 4625 2090 4665 2100
rect 4625 2070 4635 2090
rect 4655 2070 4665 2090
rect 4625 2060 4665 2070
rect 4745 2090 4785 2100
rect 4745 2070 4755 2090
rect 4775 2070 4785 2090
rect 4745 2060 4785 2070
rect 4865 2090 4905 2100
rect 4865 2070 4875 2090
rect 4895 2070 4905 2090
rect 4865 2060 4905 2070
rect 4985 2090 5025 2100
rect 4985 2070 4995 2090
rect 5015 2070 5025 2090
rect 4985 2060 5025 2070
rect 5105 2090 5145 2100
rect 5105 2070 5115 2090
rect 5135 2070 5145 2090
rect 5105 2060 5145 2070
rect 5225 2090 5265 2100
rect 5225 2070 5235 2090
rect 5255 2070 5265 2090
rect 5225 2060 5265 2070
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2060
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3895 1995 3915 2015
rect 3995 1995 4015 2060
rect 4085 2045 4125 2055
rect 4085 2025 4095 2045
rect 4115 2025 4125 2045
rect 4085 2015 4125 2025
rect 4095 1995 4115 2015
rect 4155 1995 4175 2060
rect 4275 1995 4295 2060
rect 4395 1995 4415 2060
rect 4445 2045 4485 2055
rect 4445 2025 4455 2045
rect 4475 2025 4485 2045
rect 4445 2015 4485 2025
rect 4455 1995 4475 2015
rect 4515 1995 4535 2060
rect 4635 1995 4655 2060
rect 4755 1995 4775 2060
rect 4805 2045 4845 2055
rect 4805 2025 4815 2045
rect 4835 2025 4845 2045
rect 4805 2015 4845 2025
rect 4815 1995 4835 2015
rect 4875 1995 4895 2060
rect 4995 1995 5015 2060
rect 5115 1995 5135 2060
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5175 1995 5195 2015
rect 5235 1995 5255 2060
rect 14640 2000 14675 2010
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 4060 1995
rect 3950 1965 3955 1985
rect 3975 1965 3995 1985
rect 4015 1965 4035 1985
rect 4055 1965 4060 1985
rect 3950 1935 4060 1965
rect 3950 1915 3955 1935
rect 3975 1915 3995 1935
rect 4015 1915 4035 1935
rect 4055 1915 4060 1935
rect 3950 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 5230 1985 5260 1995
rect 5230 1965 5235 1985
rect 5255 1965 5260 1985
rect 14640 1975 14645 2000
rect 14670 1975 14675 2000
rect 14640 1965 14675 1975
rect 14700 2000 14735 2010
rect 14700 1975 14705 2000
rect 14730 1975 14735 2000
rect 14700 1965 14735 1975
rect 14760 2000 14795 2010
rect 14760 1975 14765 2000
rect 14790 1975 14795 2000
rect 14760 1965 14795 1975
rect 14820 2000 14855 2010
rect 14820 1975 14825 2000
rect 14850 1975 14855 2000
rect 14820 1965 14855 1975
rect 14970 2200 15040 2230
rect 14970 2180 14975 2200
rect 14995 2180 15015 2200
rect 15035 2180 15040 2200
rect 14970 2150 15040 2180
rect 14970 2130 14975 2150
rect 14995 2130 15015 2150
rect 15035 2130 15040 2150
rect 14970 2100 15040 2130
rect 14970 2080 14975 2100
rect 14995 2080 15015 2100
rect 15035 2080 15040 2100
rect 14970 2050 15040 2080
rect 14970 2030 14975 2050
rect 14995 2030 15015 2050
rect 15035 2030 15040 2050
rect 14970 2000 15040 2030
rect 14970 1980 14975 2000
rect 14995 1980 15015 2000
rect 15035 1980 15040 2000
rect 14970 1970 15040 1980
rect 15065 2250 15095 2260
rect 15065 2230 15070 2250
rect 15090 2230 15095 2250
rect 15065 2200 15095 2230
rect 15065 2180 15070 2200
rect 15090 2180 15095 2200
rect 15065 2150 15095 2180
rect 15065 2130 15070 2150
rect 15090 2130 15095 2150
rect 15065 2100 15095 2130
rect 15065 2080 15070 2100
rect 15090 2080 15095 2100
rect 15065 2050 15095 2080
rect 15065 2030 15070 2050
rect 15090 2030 15095 2050
rect 15065 2000 15095 2030
rect 15065 1980 15070 2000
rect 15090 1980 15095 2000
rect 15065 1970 15095 1980
rect 15120 2250 15150 2260
rect 15120 2230 15125 2250
rect 15145 2230 15150 2250
rect 15120 2200 15150 2230
rect 15120 2180 15125 2200
rect 15145 2180 15150 2200
rect 15120 2150 15150 2180
rect 15120 2130 15125 2150
rect 15145 2130 15150 2150
rect 15120 2100 15150 2130
rect 15120 2080 15125 2100
rect 15145 2080 15150 2100
rect 15120 2050 15150 2080
rect 15120 2030 15125 2050
rect 15145 2030 15150 2050
rect 15120 2000 15150 2030
rect 15120 1980 15125 2000
rect 15145 1980 15150 2000
rect 15120 1970 15150 1980
rect 15175 2250 15205 2260
rect 15175 2230 15180 2250
rect 15200 2230 15205 2250
rect 15175 2200 15205 2230
rect 15175 2180 15180 2200
rect 15200 2180 15205 2200
rect 15175 2150 15205 2180
rect 15175 2130 15180 2150
rect 15200 2130 15205 2150
rect 15175 2100 15205 2130
rect 15175 2080 15180 2100
rect 15200 2080 15205 2100
rect 15175 2050 15205 2080
rect 15175 2030 15180 2050
rect 15200 2030 15205 2050
rect 15175 2000 15205 2030
rect 15175 1980 15180 2000
rect 15200 1980 15205 2000
rect 15175 1970 15205 1980
rect 15230 2250 15260 2260
rect 15230 2230 15235 2250
rect 15255 2230 15260 2250
rect 15230 2200 15260 2230
rect 15230 2180 15235 2200
rect 15255 2180 15260 2200
rect 15230 2150 15260 2180
rect 15230 2130 15235 2150
rect 15255 2130 15260 2150
rect 15230 2100 15260 2130
rect 15230 2080 15235 2100
rect 15255 2080 15260 2100
rect 15230 2050 15260 2080
rect 15230 2030 15235 2050
rect 15255 2030 15260 2050
rect 15230 2000 15260 2030
rect 15230 1980 15235 2000
rect 15255 1980 15260 2000
rect 15230 1970 15260 1980
rect 15285 2250 15315 2260
rect 15285 2230 15290 2250
rect 15310 2230 15315 2250
rect 15285 2200 15315 2230
rect 15285 2180 15290 2200
rect 15310 2180 15315 2200
rect 15285 2150 15315 2180
rect 15285 2130 15290 2150
rect 15310 2130 15315 2150
rect 15285 2100 15315 2130
rect 15285 2080 15290 2100
rect 15310 2080 15315 2100
rect 15285 2050 15315 2080
rect 15285 2030 15290 2050
rect 15310 2030 15315 2050
rect 15285 2000 15315 2030
rect 15285 1980 15290 2000
rect 15310 1980 15315 2000
rect 15285 1970 15315 1980
rect 15340 2250 15370 2260
rect 15340 2230 15345 2250
rect 15365 2230 15370 2250
rect 15340 2200 15370 2230
rect 15340 2180 15345 2200
rect 15365 2180 15370 2200
rect 15340 2150 15370 2180
rect 15340 2130 15345 2150
rect 15365 2130 15370 2150
rect 15340 2100 15370 2130
rect 15340 2080 15345 2100
rect 15365 2080 15370 2100
rect 15340 2050 15370 2080
rect 15340 2030 15345 2050
rect 15365 2030 15370 2050
rect 15340 2000 15370 2030
rect 15340 1980 15345 2000
rect 15365 1980 15370 2000
rect 15340 1970 15370 1980
rect 15395 2250 15425 2260
rect 15395 2230 15400 2250
rect 15420 2230 15425 2250
rect 15395 2200 15425 2230
rect 15395 2180 15400 2200
rect 15420 2180 15425 2200
rect 15395 2150 15425 2180
rect 15395 2130 15400 2150
rect 15420 2130 15425 2150
rect 15395 2100 15425 2130
rect 15395 2080 15400 2100
rect 15420 2080 15425 2100
rect 15395 2050 15425 2080
rect 15395 2030 15400 2050
rect 15420 2030 15425 2050
rect 15395 2000 15425 2030
rect 15395 1980 15400 2000
rect 15420 1980 15425 2000
rect 15395 1970 15425 1980
rect 15450 2250 15480 2260
rect 15450 2230 15455 2250
rect 15475 2230 15480 2250
rect 15450 2200 15480 2230
rect 15450 2180 15455 2200
rect 15475 2180 15480 2200
rect 15450 2150 15480 2180
rect 15450 2130 15455 2150
rect 15475 2130 15480 2150
rect 15450 2100 15480 2130
rect 15450 2080 15455 2100
rect 15475 2080 15480 2100
rect 15450 2050 15480 2080
rect 15450 2030 15455 2050
rect 15475 2030 15480 2050
rect 15450 2000 15480 2030
rect 15450 1980 15455 2000
rect 15475 1980 15480 2000
rect 15450 1970 15480 1980
rect 15505 2250 15535 2260
rect 15505 2230 15510 2250
rect 15530 2230 15535 2250
rect 15505 2200 15535 2230
rect 15505 2180 15510 2200
rect 15530 2180 15535 2200
rect 15505 2150 15535 2180
rect 15505 2130 15510 2150
rect 15530 2130 15535 2150
rect 15505 2100 15535 2130
rect 15505 2080 15510 2100
rect 15530 2080 15535 2100
rect 15505 2050 15535 2080
rect 15505 2030 15510 2050
rect 15530 2030 15535 2050
rect 15505 2000 15535 2030
rect 15505 1980 15510 2000
rect 15530 1980 15535 2000
rect 15505 1970 15535 1980
rect 15560 2250 15590 2260
rect 15560 2230 15565 2250
rect 15585 2230 15590 2250
rect 15560 2200 15590 2230
rect 15560 2180 15565 2200
rect 15585 2180 15590 2200
rect 15560 2150 15590 2180
rect 15560 2130 15565 2150
rect 15585 2130 15590 2150
rect 15560 2100 15590 2130
rect 15560 2080 15565 2100
rect 15585 2080 15590 2100
rect 15560 2050 15590 2080
rect 15560 2030 15565 2050
rect 15585 2030 15590 2050
rect 15560 2000 15590 2030
rect 15560 1980 15565 2000
rect 15585 1980 15590 2000
rect 15560 1970 15590 1980
rect 15615 2250 15645 2260
rect 15615 2230 15620 2250
rect 15640 2230 15645 2250
rect 15615 2200 15645 2230
rect 15615 2180 15620 2200
rect 15640 2180 15645 2200
rect 15615 2150 15645 2180
rect 15615 2130 15620 2150
rect 15640 2130 15645 2150
rect 15615 2100 15645 2130
rect 15615 2080 15620 2100
rect 15640 2080 15645 2100
rect 15615 2050 15645 2080
rect 15615 2030 15620 2050
rect 15640 2030 15645 2050
rect 15615 2000 15645 2030
rect 15615 1980 15620 2000
rect 15640 1980 15645 2000
rect 15615 1970 15645 1980
rect 15670 2250 15740 2260
rect 15670 2230 15675 2250
rect 15695 2230 15715 2250
rect 15735 2230 15740 2250
rect 15670 2200 15740 2230
rect 15670 2180 15675 2200
rect 15695 2180 15715 2200
rect 15735 2180 15740 2200
rect 18110 2250 18180 2260
rect 18110 2230 18115 2250
rect 18135 2230 18155 2250
rect 18175 2230 18180 2250
rect 18110 2200 18180 2230
rect 15670 2150 15740 2180
rect 15670 2130 15675 2150
rect 15695 2130 15715 2150
rect 15735 2130 15740 2150
rect 16330 2175 16370 2185
rect 16330 2155 16340 2175
rect 16360 2155 16370 2175
rect 16330 2145 16370 2155
rect 16440 2175 16480 2185
rect 16440 2155 16450 2175
rect 16470 2155 16480 2175
rect 16440 2145 16480 2155
rect 16550 2175 16590 2185
rect 16550 2155 16560 2175
rect 16580 2155 16590 2175
rect 16550 2145 16590 2155
rect 16660 2175 16700 2185
rect 16660 2155 16670 2175
rect 16690 2155 16700 2175
rect 16660 2145 16700 2155
rect 16770 2175 16810 2185
rect 16770 2155 16780 2175
rect 16800 2155 16810 2175
rect 16770 2145 16810 2155
rect 16828 2175 16862 2185
rect 16828 2155 16836 2175
rect 16854 2155 16862 2175
rect 16828 2145 16862 2155
rect 16880 2175 16920 2185
rect 16880 2155 16890 2175
rect 16910 2155 16920 2175
rect 16880 2145 16920 2155
rect 16990 2175 17030 2185
rect 16990 2155 17000 2175
rect 17020 2155 17030 2175
rect 16990 2145 17030 2155
rect 17100 2175 17140 2185
rect 17100 2155 17110 2175
rect 17130 2155 17140 2175
rect 17100 2145 17140 2155
rect 17210 2175 17250 2185
rect 17210 2155 17220 2175
rect 17240 2155 17250 2175
rect 17210 2145 17250 2155
rect 17320 2175 17360 2185
rect 17320 2155 17330 2175
rect 17350 2155 17360 2175
rect 17320 2145 17360 2155
rect 17430 2175 17470 2185
rect 17430 2155 17440 2175
rect 17460 2155 17470 2175
rect 17430 2145 17470 2155
rect 18110 2180 18115 2200
rect 18135 2180 18155 2200
rect 18175 2180 18180 2200
rect 18110 2150 18180 2180
rect 15670 2100 15740 2130
rect 16340 2125 16360 2145
rect 16450 2125 16470 2145
rect 16560 2125 16580 2145
rect 16670 2125 16690 2145
rect 16780 2125 16800 2145
rect 16890 2125 16910 2145
rect 17000 2125 17020 2145
rect 17110 2125 17130 2145
rect 17220 2125 17240 2145
rect 17330 2125 17350 2145
rect 17440 2125 17460 2145
rect 18110 2130 18115 2150
rect 18135 2130 18155 2150
rect 18175 2130 18180 2150
rect 15670 2080 15675 2100
rect 15695 2080 15715 2100
rect 15735 2080 15740 2100
rect 15670 2050 15740 2080
rect 15670 2030 15675 2050
rect 15695 2030 15715 2050
rect 15735 2030 15740 2050
rect 15670 2000 15740 2030
rect 15670 1980 15675 2000
rect 15695 1980 15715 2000
rect 15735 1980 15740 2000
rect 16240 2115 16310 2125
rect 16240 2095 16245 2115
rect 16265 2095 16285 2115
rect 16305 2095 16310 2115
rect 16240 2065 16310 2095
rect 16240 2045 16245 2065
rect 16265 2045 16285 2065
rect 16305 2045 16310 2065
rect 16240 2015 16310 2045
rect 16240 1995 16245 2015
rect 16265 1995 16285 2015
rect 16305 1995 16310 2015
rect 16240 1985 16310 1995
rect 16335 2115 16365 2125
rect 16335 2095 16340 2115
rect 16360 2095 16365 2115
rect 16335 2065 16365 2095
rect 16335 2045 16340 2065
rect 16360 2045 16365 2065
rect 16335 2015 16365 2045
rect 16335 1995 16340 2015
rect 16360 1995 16365 2015
rect 16335 1985 16365 1995
rect 16390 2115 16420 2125
rect 16390 2095 16395 2115
rect 16415 2095 16420 2115
rect 16390 2065 16420 2095
rect 16390 2045 16395 2065
rect 16415 2045 16420 2065
rect 16390 2015 16420 2045
rect 16390 1995 16395 2015
rect 16415 1995 16420 2015
rect 16390 1985 16420 1995
rect 16445 2115 16475 2125
rect 16445 2095 16450 2115
rect 16470 2095 16475 2115
rect 16445 2065 16475 2095
rect 16445 2045 16450 2065
rect 16470 2045 16475 2065
rect 16445 2015 16475 2045
rect 16445 1995 16450 2015
rect 16470 1995 16475 2015
rect 16445 1985 16475 1995
rect 16500 2115 16530 2125
rect 16500 2095 16505 2115
rect 16525 2095 16530 2115
rect 16500 2065 16530 2095
rect 16500 2045 16505 2065
rect 16525 2045 16530 2065
rect 16500 2015 16530 2045
rect 16500 1995 16505 2015
rect 16525 1995 16530 2015
rect 16500 1985 16530 1995
rect 16555 2115 16585 2125
rect 16555 2095 16560 2115
rect 16580 2095 16585 2115
rect 16555 2065 16585 2095
rect 16555 2045 16560 2065
rect 16580 2045 16585 2065
rect 16555 2015 16585 2045
rect 16555 1995 16560 2015
rect 16580 1995 16585 2015
rect 16555 1985 16585 1995
rect 16610 2115 16640 2125
rect 16610 2095 16615 2115
rect 16635 2095 16640 2115
rect 16610 2065 16640 2095
rect 16610 2045 16615 2065
rect 16635 2045 16640 2065
rect 16610 2015 16640 2045
rect 16610 1995 16615 2015
rect 16635 1995 16640 2015
rect 16610 1985 16640 1995
rect 16665 2115 16695 2125
rect 16665 2095 16670 2115
rect 16690 2095 16695 2115
rect 16665 2065 16695 2095
rect 16665 2045 16670 2065
rect 16690 2045 16695 2065
rect 16665 2015 16695 2045
rect 16665 1995 16670 2015
rect 16690 1995 16695 2015
rect 16665 1985 16695 1995
rect 16720 2115 16750 2125
rect 16720 2095 16725 2115
rect 16745 2095 16750 2115
rect 16720 2065 16750 2095
rect 16720 2045 16725 2065
rect 16745 2045 16750 2065
rect 16720 2015 16750 2045
rect 16720 1995 16725 2015
rect 16745 1995 16750 2015
rect 16720 1985 16750 1995
rect 16775 2115 16805 2125
rect 16775 2095 16780 2115
rect 16800 2095 16805 2115
rect 16775 2065 16805 2095
rect 16775 2045 16780 2065
rect 16800 2045 16805 2065
rect 16775 2015 16805 2045
rect 16775 1995 16780 2015
rect 16800 1995 16805 2015
rect 16775 1985 16805 1995
rect 16830 2115 16860 2125
rect 16830 2095 16835 2115
rect 16855 2095 16860 2115
rect 16830 2065 16860 2095
rect 16830 2045 16835 2065
rect 16855 2045 16860 2065
rect 16830 2015 16860 2045
rect 16830 1995 16835 2015
rect 16855 1995 16860 2015
rect 16830 1985 16860 1995
rect 16885 2115 16915 2125
rect 16885 2095 16890 2115
rect 16910 2095 16915 2115
rect 16885 2065 16915 2095
rect 16885 2045 16890 2065
rect 16910 2045 16915 2065
rect 16885 2015 16915 2045
rect 16885 1995 16890 2015
rect 16910 1995 16915 2015
rect 16885 1985 16915 1995
rect 16940 2115 16970 2125
rect 16940 2095 16945 2115
rect 16965 2095 16970 2115
rect 16940 2065 16970 2095
rect 16940 2045 16945 2065
rect 16965 2045 16970 2065
rect 16940 2015 16970 2045
rect 16940 1995 16945 2015
rect 16965 1995 16970 2015
rect 16940 1985 16970 1995
rect 16995 2115 17025 2125
rect 16995 2095 17000 2115
rect 17020 2095 17025 2115
rect 16995 2065 17025 2095
rect 16995 2045 17000 2065
rect 17020 2045 17025 2065
rect 16995 2015 17025 2045
rect 16995 1995 17000 2015
rect 17020 1995 17025 2015
rect 16995 1985 17025 1995
rect 17050 2115 17080 2125
rect 17050 2095 17055 2115
rect 17075 2095 17080 2115
rect 17050 2065 17080 2095
rect 17050 2045 17055 2065
rect 17075 2045 17080 2065
rect 17050 2015 17080 2045
rect 17050 1995 17055 2015
rect 17075 1995 17080 2015
rect 17050 1985 17080 1995
rect 17105 2115 17135 2125
rect 17105 2095 17110 2115
rect 17130 2095 17135 2115
rect 17105 2065 17135 2095
rect 17105 2045 17110 2065
rect 17130 2045 17135 2065
rect 17105 2015 17135 2045
rect 17105 1995 17110 2015
rect 17130 1995 17135 2015
rect 17105 1985 17135 1995
rect 17160 2115 17190 2125
rect 17160 2095 17165 2115
rect 17185 2095 17190 2115
rect 17160 2065 17190 2095
rect 17160 2045 17165 2065
rect 17185 2045 17190 2065
rect 17160 2015 17190 2045
rect 17160 1995 17165 2015
rect 17185 1995 17190 2015
rect 17160 1985 17190 1995
rect 17215 2115 17245 2125
rect 17215 2095 17220 2115
rect 17240 2095 17245 2115
rect 17215 2065 17245 2095
rect 17215 2045 17220 2065
rect 17240 2045 17245 2065
rect 17215 2015 17245 2045
rect 17215 1995 17220 2015
rect 17240 1995 17245 2015
rect 17215 1985 17245 1995
rect 17270 2115 17300 2125
rect 17270 2095 17275 2115
rect 17295 2095 17300 2115
rect 17270 2065 17300 2095
rect 17270 2045 17275 2065
rect 17295 2045 17300 2065
rect 17270 2015 17300 2045
rect 17270 1995 17275 2015
rect 17295 1995 17300 2015
rect 17270 1985 17300 1995
rect 17325 2115 17355 2125
rect 17325 2095 17330 2115
rect 17350 2095 17355 2115
rect 17325 2065 17355 2095
rect 17325 2045 17330 2065
rect 17350 2045 17355 2065
rect 17325 2015 17355 2045
rect 17325 1995 17330 2015
rect 17350 1995 17355 2015
rect 17325 1985 17355 1995
rect 17380 2115 17410 2125
rect 17380 2095 17385 2115
rect 17405 2095 17410 2115
rect 17380 2065 17410 2095
rect 17380 2045 17385 2065
rect 17405 2045 17410 2065
rect 17380 2015 17410 2045
rect 17380 1995 17385 2015
rect 17405 1995 17410 2015
rect 17380 1985 17410 1995
rect 17435 2115 17465 2125
rect 17435 2095 17440 2115
rect 17460 2095 17465 2115
rect 17435 2065 17465 2095
rect 17435 2045 17440 2065
rect 17460 2045 17465 2065
rect 17435 2015 17465 2045
rect 17435 1995 17440 2015
rect 17460 1995 17465 2015
rect 17435 1985 17465 1995
rect 17490 2115 17560 2125
rect 17490 2095 17495 2115
rect 17515 2095 17535 2115
rect 17555 2095 17560 2115
rect 17490 2065 17560 2095
rect 17490 2045 17495 2065
rect 17515 2045 17535 2065
rect 17555 2045 17560 2065
rect 17490 2015 17560 2045
rect 17490 1995 17495 2015
rect 17515 1995 17535 2015
rect 17555 1995 17560 2015
rect 17490 1985 17560 1995
rect 18110 2100 18180 2130
rect 18110 2080 18115 2100
rect 18135 2080 18155 2100
rect 18175 2080 18180 2100
rect 18110 2050 18180 2080
rect 18110 2030 18115 2050
rect 18135 2030 18155 2050
rect 18175 2030 18180 2050
rect 18110 2000 18180 2030
rect 15670 1970 15740 1980
rect 5230 1935 5260 1965
rect 15070 1950 15090 1970
rect 15180 1950 15200 1970
rect 15290 1950 15310 1970
rect 15400 1950 15420 1970
rect 15510 1950 15530 1970
rect 15620 1950 15640 1970
rect 16245 1965 16265 1985
rect 16395 1965 16415 1985
rect 16505 1965 16525 1985
rect 16615 1965 16635 1985
rect 16725 1965 16745 1985
rect 16835 1965 16855 1985
rect 16945 1965 16965 1985
rect 17055 1965 17075 1985
rect 17165 1965 17185 1985
rect 17275 1965 17295 1985
rect 17385 1965 17405 1985
rect 17535 1965 17555 1985
rect 18110 1980 18115 2000
rect 18135 1980 18155 2000
rect 18175 1980 18180 2000
rect 18110 1970 18180 1980
rect 18205 2250 18235 2260
rect 18205 2230 18210 2250
rect 18230 2230 18235 2250
rect 18205 2200 18235 2230
rect 18205 2180 18210 2200
rect 18230 2180 18235 2200
rect 18205 2150 18235 2180
rect 18205 2130 18210 2150
rect 18230 2130 18235 2150
rect 18205 2100 18235 2130
rect 18205 2080 18210 2100
rect 18230 2080 18235 2100
rect 18205 2050 18235 2080
rect 18205 2030 18210 2050
rect 18230 2030 18235 2050
rect 18205 2000 18235 2030
rect 18205 1980 18210 2000
rect 18230 1980 18235 2000
rect 18205 1970 18235 1980
rect 18260 2250 18290 2260
rect 18260 2230 18265 2250
rect 18285 2230 18290 2250
rect 18260 2200 18290 2230
rect 18260 2180 18265 2200
rect 18285 2180 18290 2200
rect 18260 2150 18290 2180
rect 18260 2130 18265 2150
rect 18285 2130 18290 2150
rect 18260 2100 18290 2130
rect 18260 2080 18265 2100
rect 18285 2080 18290 2100
rect 18260 2050 18290 2080
rect 18260 2030 18265 2050
rect 18285 2030 18290 2050
rect 18260 2000 18290 2030
rect 18260 1980 18265 2000
rect 18285 1980 18290 2000
rect 18260 1970 18290 1980
rect 18315 2250 18345 2260
rect 18315 2230 18320 2250
rect 18340 2230 18345 2250
rect 18315 2200 18345 2230
rect 18315 2180 18320 2200
rect 18340 2180 18345 2200
rect 18315 2150 18345 2180
rect 18315 2130 18320 2150
rect 18340 2130 18345 2150
rect 18315 2100 18345 2130
rect 18315 2080 18320 2100
rect 18340 2080 18345 2100
rect 18315 2050 18345 2080
rect 18315 2030 18320 2050
rect 18340 2030 18345 2050
rect 18315 2000 18345 2030
rect 18315 1980 18320 2000
rect 18340 1980 18345 2000
rect 18315 1970 18345 1980
rect 18370 2250 18400 2260
rect 18370 2230 18375 2250
rect 18395 2230 18400 2250
rect 18370 2200 18400 2230
rect 18370 2180 18375 2200
rect 18395 2180 18400 2200
rect 18370 2150 18400 2180
rect 18370 2130 18375 2150
rect 18395 2130 18400 2150
rect 18370 2100 18400 2130
rect 18370 2080 18375 2100
rect 18395 2080 18400 2100
rect 18370 2050 18400 2080
rect 18370 2030 18375 2050
rect 18395 2030 18400 2050
rect 18370 2000 18400 2030
rect 18370 1980 18375 2000
rect 18395 1980 18400 2000
rect 18370 1970 18400 1980
rect 18425 2250 18455 2260
rect 18425 2230 18430 2250
rect 18450 2230 18455 2250
rect 18425 2200 18455 2230
rect 18425 2180 18430 2200
rect 18450 2180 18455 2200
rect 18425 2150 18455 2180
rect 18425 2130 18430 2150
rect 18450 2130 18455 2150
rect 18425 2100 18455 2130
rect 18425 2080 18430 2100
rect 18450 2080 18455 2100
rect 18425 2050 18455 2080
rect 18425 2030 18430 2050
rect 18450 2030 18455 2050
rect 18425 2000 18455 2030
rect 18425 1980 18430 2000
rect 18450 1980 18455 2000
rect 18425 1970 18455 1980
rect 18480 2250 18510 2260
rect 18480 2230 18485 2250
rect 18505 2230 18510 2250
rect 18480 2200 18510 2230
rect 18480 2180 18485 2200
rect 18505 2180 18510 2200
rect 18480 2150 18510 2180
rect 18480 2130 18485 2150
rect 18505 2130 18510 2150
rect 18480 2100 18510 2130
rect 18480 2080 18485 2100
rect 18505 2080 18510 2100
rect 18480 2050 18510 2080
rect 18480 2030 18485 2050
rect 18505 2030 18510 2050
rect 18480 2000 18510 2030
rect 18480 1980 18485 2000
rect 18505 1980 18510 2000
rect 18480 1970 18510 1980
rect 18535 2250 18565 2260
rect 18535 2230 18540 2250
rect 18560 2230 18565 2250
rect 18535 2200 18565 2230
rect 18535 2180 18540 2200
rect 18560 2180 18565 2200
rect 18535 2150 18565 2180
rect 18535 2130 18540 2150
rect 18560 2130 18565 2150
rect 18535 2100 18565 2130
rect 18535 2080 18540 2100
rect 18560 2080 18565 2100
rect 18535 2050 18565 2080
rect 18535 2030 18540 2050
rect 18560 2030 18565 2050
rect 18535 2000 18565 2030
rect 18535 1980 18540 2000
rect 18560 1980 18565 2000
rect 18535 1970 18565 1980
rect 18590 2250 18620 2260
rect 18590 2230 18595 2250
rect 18615 2230 18620 2250
rect 18590 2200 18620 2230
rect 18590 2180 18595 2200
rect 18615 2180 18620 2200
rect 18590 2150 18620 2180
rect 18590 2130 18595 2150
rect 18615 2130 18620 2150
rect 18590 2100 18620 2130
rect 18590 2080 18595 2100
rect 18615 2080 18620 2100
rect 18590 2050 18620 2080
rect 18590 2030 18595 2050
rect 18615 2030 18620 2050
rect 18590 2000 18620 2030
rect 18590 1980 18595 2000
rect 18615 1980 18620 2000
rect 18590 1970 18620 1980
rect 18645 2250 18675 2260
rect 18645 2230 18650 2250
rect 18670 2230 18675 2250
rect 18645 2200 18675 2230
rect 18645 2180 18650 2200
rect 18670 2180 18675 2200
rect 18645 2150 18675 2180
rect 18645 2130 18650 2150
rect 18670 2130 18675 2150
rect 18645 2100 18675 2130
rect 18645 2080 18650 2100
rect 18670 2080 18675 2100
rect 18645 2050 18675 2080
rect 18645 2030 18650 2050
rect 18670 2030 18675 2050
rect 18645 2000 18675 2030
rect 18645 1980 18650 2000
rect 18670 1980 18675 2000
rect 18645 1970 18675 1980
rect 18700 2250 18730 2260
rect 18700 2230 18705 2250
rect 18725 2230 18730 2250
rect 18700 2200 18730 2230
rect 18700 2180 18705 2200
rect 18725 2180 18730 2200
rect 18700 2150 18730 2180
rect 18700 2130 18705 2150
rect 18725 2130 18730 2150
rect 18700 2100 18730 2130
rect 18700 2080 18705 2100
rect 18725 2080 18730 2100
rect 18700 2050 18730 2080
rect 18700 2030 18705 2050
rect 18725 2030 18730 2050
rect 18700 2000 18730 2030
rect 18700 1980 18705 2000
rect 18725 1980 18730 2000
rect 18700 1970 18730 1980
rect 18755 2250 18785 2260
rect 18755 2230 18760 2250
rect 18780 2230 18785 2250
rect 18755 2200 18785 2230
rect 18755 2180 18760 2200
rect 18780 2180 18785 2200
rect 18755 2150 18785 2180
rect 18755 2130 18760 2150
rect 18780 2130 18785 2150
rect 18755 2100 18785 2130
rect 18755 2080 18760 2100
rect 18780 2080 18785 2100
rect 18755 2050 18785 2080
rect 18755 2030 18760 2050
rect 18780 2030 18785 2050
rect 18755 2000 18785 2030
rect 18755 1980 18760 2000
rect 18780 1980 18785 2000
rect 18755 1970 18785 1980
rect 18810 2250 18880 2260
rect 18810 2230 18815 2250
rect 18835 2230 18855 2250
rect 18875 2230 18880 2250
rect 24970 2250 25040 2260
rect 24970 2230 24975 2250
rect 24995 2230 25015 2250
rect 25035 2230 25040 2250
rect 18810 2200 18880 2230
rect 18810 2180 18815 2200
rect 18835 2180 18855 2200
rect 18875 2180 18880 2200
rect 18810 2150 18880 2180
rect 18810 2130 18815 2150
rect 18835 2130 18855 2150
rect 18875 2130 18880 2150
rect 18810 2100 18880 2130
rect 18810 2080 18815 2100
rect 18835 2080 18855 2100
rect 18875 2080 18880 2100
rect 18810 2050 18880 2080
rect 18810 2030 18815 2050
rect 18835 2030 18855 2050
rect 18875 2030 18880 2050
rect 18810 2000 18880 2030
rect 18810 1980 18815 2000
rect 18835 1980 18855 2000
rect 18875 1980 18880 2000
rect 18810 1970 18880 1980
rect 18995 2000 19030 2010
rect 18995 1975 19000 2000
rect 19025 1975 19030 2000
rect 16235 1955 16275 1965
rect 5230 1915 5235 1935
rect 5255 1915 5260 1935
rect 5230 1905 5260 1915
rect 15060 1940 15100 1950
rect 15060 1920 15070 1940
rect 15088 1920 15100 1940
rect 15060 1910 15100 1920
rect 15170 1940 15210 1950
rect 15170 1920 15180 1940
rect 15198 1920 15210 1940
rect 15170 1910 15210 1920
rect 15280 1940 15320 1950
rect 15280 1920 15290 1940
rect 15308 1920 15320 1940
rect 15280 1910 15320 1920
rect 15390 1940 15430 1950
rect 15390 1920 15400 1940
rect 15418 1920 15430 1940
rect 15390 1910 15430 1920
rect 15500 1940 15540 1950
rect 15500 1920 15510 1940
rect 15528 1920 15540 1940
rect 15500 1910 15540 1920
rect 15610 1940 15650 1950
rect 15610 1920 15620 1940
rect 15638 1920 15650 1940
rect 16235 1935 16245 1955
rect 16265 1935 16275 1955
rect 16235 1925 16275 1935
rect 16385 1955 16425 1965
rect 16385 1935 16395 1955
rect 16415 1935 16425 1955
rect 16385 1925 16425 1935
rect 16495 1955 16535 1965
rect 16495 1935 16505 1955
rect 16525 1935 16535 1955
rect 16495 1925 16535 1935
rect 16605 1955 16645 1965
rect 16605 1935 16615 1955
rect 16635 1935 16645 1955
rect 16605 1925 16645 1935
rect 16715 1955 16755 1965
rect 16715 1935 16725 1955
rect 16745 1935 16755 1955
rect 16715 1925 16755 1935
rect 16825 1955 16865 1965
rect 16825 1935 16835 1955
rect 16855 1935 16865 1955
rect 16825 1925 16865 1935
rect 16935 1955 16975 1965
rect 16935 1935 16945 1955
rect 16965 1935 16975 1955
rect 16935 1925 16975 1935
rect 17045 1955 17085 1965
rect 17045 1935 17055 1955
rect 17075 1935 17085 1955
rect 17045 1925 17085 1935
rect 17155 1955 17195 1965
rect 17155 1935 17165 1955
rect 17185 1935 17195 1955
rect 17155 1925 17195 1935
rect 17265 1955 17305 1965
rect 17265 1935 17275 1955
rect 17295 1935 17305 1955
rect 17265 1925 17305 1935
rect 17375 1955 17415 1965
rect 17375 1935 17385 1955
rect 17405 1935 17415 1955
rect 17375 1925 17415 1935
rect 17525 1955 17565 1965
rect 17525 1935 17535 1955
rect 17555 1935 17565 1955
rect 18210 1950 18230 1970
rect 18320 1950 18340 1970
rect 18430 1950 18450 1970
rect 18540 1950 18560 1970
rect 18650 1950 18670 1970
rect 18760 1950 18780 1970
rect 18995 1965 19030 1975
rect 19055 2000 19090 2010
rect 19055 1975 19060 2000
rect 19085 1975 19090 2000
rect 19055 1965 19090 1975
rect 19115 2000 19150 2010
rect 19115 1975 19120 2000
rect 19145 1975 19150 2000
rect 19115 1965 19150 1975
rect 19175 2000 19210 2010
rect 19175 1975 19180 2000
rect 19205 1975 19210 2000
rect 19175 1965 19210 1975
rect 24640 2000 24675 2010
rect 24640 1975 24645 2000
rect 24670 1975 24675 2000
rect 24640 1965 24675 1975
rect 24700 2000 24735 2010
rect 24700 1975 24705 2000
rect 24730 1975 24735 2000
rect 24700 1965 24735 1975
rect 24760 2000 24795 2010
rect 24760 1975 24765 2000
rect 24790 1975 24795 2000
rect 24760 1965 24795 1975
rect 24820 2000 24855 2010
rect 24820 1975 24825 2000
rect 24850 1975 24855 2000
rect 24820 1965 24855 1975
rect 24970 2200 25040 2230
rect 24970 2180 24975 2200
rect 24995 2180 25015 2200
rect 25035 2180 25040 2200
rect 24970 2150 25040 2180
rect 24970 2130 24975 2150
rect 24995 2130 25015 2150
rect 25035 2130 25040 2150
rect 24970 2100 25040 2130
rect 24970 2080 24975 2100
rect 24995 2080 25015 2100
rect 25035 2080 25040 2100
rect 24970 2050 25040 2080
rect 24970 2030 24975 2050
rect 24995 2030 25015 2050
rect 25035 2030 25040 2050
rect 24970 2000 25040 2030
rect 24970 1980 24975 2000
rect 24995 1980 25015 2000
rect 25035 1980 25040 2000
rect 24970 1970 25040 1980
rect 25065 2250 25095 2260
rect 25065 2230 25070 2250
rect 25090 2230 25095 2250
rect 25065 2200 25095 2230
rect 25065 2180 25070 2200
rect 25090 2180 25095 2200
rect 25065 2150 25095 2180
rect 25065 2130 25070 2150
rect 25090 2130 25095 2150
rect 25065 2100 25095 2130
rect 25065 2080 25070 2100
rect 25090 2080 25095 2100
rect 25065 2050 25095 2080
rect 25065 2030 25070 2050
rect 25090 2030 25095 2050
rect 25065 2000 25095 2030
rect 25065 1980 25070 2000
rect 25090 1980 25095 2000
rect 25065 1970 25095 1980
rect 25120 2250 25150 2260
rect 25120 2230 25125 2250
rect 25145 2230 25150 2250
rect 25120 2200 25150 2230
rect 25120 2180 25125 2200
rect 25145 2180 25150 2200
rect 25120 2150 25150 2180
rect 25120 2130 25125 2150
rect 25145 2130 25150 2150
rect 25120 2100 25150 2130
rect 25120 2080 25125 2100
rect 25145 2080 25150 2100
rect 25120 2050 25150 2080
rect 25120 2030 25125 2050
rect 25145 2030 25150 2050
rect 25120 2000 25150 2030
rect 25120 1980 25125 2000
rect 25145 1980 25150 2000
rect 25120 1970 25150 1980
rect 25175 2250 25205 2260
rect 25175 2230 25180 2250
rect 25200 2230 25205 2250
rect 25175 2200 25205 2230
rect 25175 2180 25180 2200
rect 25200 2180 25205 2200
rect 25175 2150 25205 2180
rect 25175 2130 25180 2150
rect 25200 2130 25205 2150
rect 25175 2100 25205 2130
rect 25175 2080 25180 2100
rect 25200 2080 25205 2100
rect 25175 2050 25205 2080
rect 25175 2030 25180 2050
rect 25200 2030 25205 2050
rect 25175 2000 25205 2030
rect 25175 1980 25180 2000
rect 25200 1980 25205 2000
rect 25175 1970 25205 1980
rect 25230 2250 25260 2260
rect 25230 2230 25235 2250
rect 25255 2230 25260 2250
rect 25230 2200 25260 2230
rect 25230 2180 25235 2200
rect 25255 2180 25260 2200
rect 25230 2150 25260 2180
rect 25230 2130 25235 2150
rect 25255 2130 25260 2150
rect 25230 2100 25260 2130
rect 25230 2080 25235 2100
rect 25255 2080 25260 2100
rect 25230 2050 25260 2080
rect 25230 2030 25235 2050
rect 25255 2030 25260 2050
rect 25230 2000 25260 2030
rect 25230 1980 25235 2000
rect 25255 1980 25260 2000
rect 25230 1970 25260 1980
rect 25285 2250 25315 2260
rect 25285 2230 25290 2250
rect 25310 2230 25315 2250
rect 25285 2200 25315 2230
rect 25285 2180 25290 2200
rect 25310 2180 25315 2200
rect 25285 2150 25315 2180
rect 25285 2130 25290 2150
rect 25310 2130 25315 2150
rect 25285 2100 25315 2130
rect 25285 2080 25290 2100
rect 25310 2080 25315 2100
rect 25285 2050 25315 2080
rect 25285 2030 25290 2050
rect 25310 2030 25315 2050
rect 25285 2000 25315 2030
rect 25285 1980 25290 2000
rect 25310 1980 25315 2000
rect 25285 1970 25315 1980
rect 25340 2250 25370 2260
rect 25340 2230 25345 2250
rect 25365 2230 25370 2250
rect 25340 2200 25370 2230
rect 25340 2180 25345 2200
rect 25365 2180 25370 2200
rect 25340 2150 25370 2180
rect 25340 2130 25345 2150
rect 25365 2130 25370 2150
rect 25340 2100 25370 2130
rect 25340 2080 25345 2100
rect 25365 2080 25370 2100
rect 25340 2050 25370 2080
rect 25340 2030 25345 2050
rect 25365 2030 25370 2050
rect 25340 2000 25370 2030
rect 25340 1980 25345 2000
rect 25365 1980 25370 2000
rect 25340 1970 25370 1980
rect 25395 2250 25425 2260
rect 25395 2230 25400 2250
rect 25420 2230 25425 2250
rect 25395 2200 25425 2230
rect 25395 2180 25400 2200
rect 25420 2180 25425 2200
rect 25395 2150 25425 2180
rect 25395 2130 25400 2150
rect 25420 2130 25425 2150
rect 25395 2100 25425 2130
rect 25395 2080 25400 2100
rect 25420 2080 25425 2100
rect 25395 2050 25425 2080
rect 25395 2030 25400 2050
rect 25420 2030 25425 2050
rect 25395 2000 25425 2030
rect 25395 1980 25400 2000
rect 25420 1980 25425 2000
rect 25395 1970 25425 1980
rect 25450 2250 25480 2260
rect 25450 2230 25455 2250
rect 25475 2230 25480 2250
rect 25450 2200 25480 2230
rect 25450 2180 25455 2200
rect 25475 2180 25480 2200
rect 25450 2150 25480 2180
rect 25450 2130 25455 2150
rect 25475 2130 25480 2150
rect 25450 2100 25480 2130
rect 25450 2080 25455 2100
rect 25475 2080 25480 2100
rect 25450 2050 25480 2080
rect 25450 2030 25455 2050
rect 25475 2030 25480 2050
rect 25450 2000 25480 2030
rect 25450 1980 25455 2000
rect 25475 1980 25480 2000
rect 25450 1970 25480 1980
rect 25505 2250 25535 2260
rect 25505 2230 25510 2250
rect 25530 2230 25535 2250
rect 25505 2200 25535 2230
rect 25505 2180 25510 2200
rect 25530 2180 25535 2200
rect 25505 2150 25535 2180
rect 25505 2130 25510 2150
rect 25530 2130 25535 2150
rect 25505 2100 25535 2130
rect 25505 2080 25510 2100
rect 25530 2080 25535 2100
rect 25505 2050 25535 2080
rect 25505 2030 25510 2050
rect 25530 2030 25535 2050
rect 25505 2000 25535 2030
rect 25505 1980 25510 2000
rect 25530 1980 25535 2000
rect 25505 1970 25535 1980
rect 25560 2250 25590 2260
rect 25560 2230 25565 2250
rect 25585 2230 25590 2250
rect 25560 2200 25590 2230
rect 25560 2180 25565 2200
rect 25585 2180 25590 2200
rect 25560 2150 25590 2180
rect 25560 2130 25565 2150
rect 25585 2130 25590 2150
rect 25560 2100 25590 2130
rect 25560 2080 25565 2100
rect 25585 2080 25590 2100
rect 25560 2050 25590 2080
rect 25560 2030 25565 2050
rect 25585 2030 25590 2050
rect 25560 2000 25590 2030
rect 25560 1980 25565 2000
rect 25585 1980 25590 2000
rect 25560 1970 25590 1980
rect 25615 2250 25645 2260
rect 25615 2230 25620 2250
rect 25640 2230 25645 2250
rect 25615 2200 25645 2230
rect 25615 2180 25620 2200
rect 25640 2180 25645 2200
rect 25615 2150 25645 2180
rect 25615 2130 25620 2150
rect 25640 2130 25645 2150
rect 25615 2100 25645 2130
rect 25615 2080 25620 2100
rect 25640 2080 25645 2100
rect 25615 2050 25645 2080
rect 25615 2030 25620 2050
rect 25640 2030 25645 2050
rect 25615 2000 25645 2030
rect 25615 1980 25620 2000
rect 25640 1980 25645 2000
rect 25615 1970 25645 1980
rect 25670 2250 25740 2260
rect 25670 2230 25675 2250
rect 25695 2230 25715 2250
rect 25735 2230 25740 2250
rect 25670 2200 25740 2230
rect 25670 2180 25675 2200
rect 25695 2180 25715 2200
rect 25735 2180 25740 2200
rect 25670 2150 25740 2180
rect 25670 2130 25675 2150
rect 25695 2130 25715 2150
rect 25735 2130 25740 2150
rect 25670 2100 25740 2130
rect 25670 2080 25675 2100
rect 25695 2080 25715 2100
rect 25735 2080 25740 2100
rect 25670 2050 25740 2080
rect 25670 2030 25675 2050
rect 25695 2030 25715 2050
rect 25735 2030 25740 2050
rect 25670 2000 25740 2030
rect 25670 1980 25675 2000
rect 25695 1980 25715 2000
rect 25735 1980 25740 2000
rect 25670 1970 25740 1980
rect 26225 2205 26860 2225
rect 26940 2205 27575 2225
rect 26225 2090 26245 2205
rect 26330 2175 26370 2185
rect 26330 2155 26340 2175
rect 26360 2155 26370 2175
rect 26330 2145 26370 2155
rect 26440 2175 26480 2185
rect 26440 2155 26450 2175
rect 26470 2155 26480 2175
rect 26440 2145 26480 2155
rect 26550 2175 26590 2185
rect 26550 2155 26560 2175
rect 26580 2155 26590 2175
rect 26550 2145 26590 2155
rect 26660 2175 26700 2185
rect 26660 2155 26670 2175
rect 26690 2155 26700 2175
rect 26660 2145 26700 2155
rect 26770 2175 26810 2185
rect 26770 2155 26780 2175
rect 26800 2155 26810 2175
rect 26770 2145 26810 2155
rect 26828 2175 26862 2185
rect 26828 2155 26836 2175
rect 26854 2155 26862 2175
rect 26828 2145 26862 2155
rect 26880 2175 26920 2185
rect 26880 2155 26890 2175
rect 26910 2155 26920 2175
rect 26880 2145 26920 2155
rect 26990 2175 27030 2185
rect 26990 2155 27000 2175
rect 27020 2155 27030 2175
rect 26990 2145 27030 2155
rect 27100 2175 27140 2185
rect 27100 2155 27110 2175
rect 27130 2155 27140 2175
rect 27100 2145 27140 2155
rect 27210 2175 27250 2185
rect 27210 2155 27220 2175
rect 27240 2155 27250 2175
rect 27210 2145 27250 2155
rect 27320 2175 27360 2185
rect 27320 2155 27330 2175
rect 27350 2155 27360 2175
rect 27320 2145 27360 2155
rect 27430 2175 27470 2185
rect 27430 2155 27440 2175
rect 27460 2155 27470 2175
rect 27430 2145 27470 2155
rect 26340 2125 26360 2145
rect 26450 2125 26470 2145
rect 26560 2125 26580 2145
rect 26670 2125 26690 2145
rect 26780 2125 26800 2145
rect 26890 2125 26910 2145
rect 27000 2125 27020 2145
rect 27110 2125 27130 2145
rect 27220 2125 27240 2145
rect 27330 2125 27350 2145
rect 27440 2125 27460 2145
rect 25070 1950 25090 1970
rect 25180 1950 25200 1970
rect 25290 1950 25310 1970
rect 25400 1950 25420 1970
rect 25510 1950 25530 1970
rect 25620 1950 25640 1970
rect 17525 1925 17565 1935
rect 18200 1940 18240 1950
rect 15610 1910 15650 1920
rect 18200 1920 18212 1940
rect 18230 1920 18240 1940
rect 18200 1910 18240 1920
rect 18310 1940 18350 1950
rect 18310 1920 18322 1940
rect 18340 1920 18350 1940
rect 18310 1910 18350 1920
rect 18420 1940 18460 1950
rect 18420 1920 18432 1940
rect 18450 1920 18460 1940
rect 18420 1910 18460 1920
rect 18530 1940 18570 1950
rect 18530 1920 18542 1940
rect 18560 1920 18570 1940
rect 18530 1910 18570 1920
rect 18640 1940 18680 1950
rect 18640 1920 18652 1940
rect 18670 1920 18680 1940
rect 18640 1910 18680 1920
rect 18750 1940 18790 1950
rect 18750 1920 18762 1940
rect 18780 1920 18790 1940
rect 18750 1910 18790 1920
rect 25060 1940 25100 1950
rect 25060 1920 25070 1940
rect 25088 1920 25100 1940
rect 25060 1910 25100 1920
rect 25170 1940 25210 1950
rect 25170 1920 25180 1940
rect 25198 1920 25210 1940
rect 25170 1910 25210 1920
rect 25280 1940 25320 1950
rect 25280 1920 25290 1940
rect 25308 1920 25320 1940
rect 25280 1910 25320 1920
rect 25390 1940 25430 1950
rect 25390 1920 25400 1940
rect 25418 1920 25430 1940
rect 25390 1910 25430 1920
rect 25500 1940 25540 1950
rect 25500 1920 25510 1940
rect 25528 1920 25540 1940
rect 25500 1910 25540 1920
rect 25610 1940 25650 1950
rect 25610 1920 25620 1940
rect 25638 1920 25650 1940
rect 25610 1910 25650 1920
rect 26225 1905 26245 2010
rect 26280 2115 26310 2125
rect 26280 2095 26285 2115
rect 26305 2095 26310 2115
rect 26280 2065 26310 2095
rect 26280 2045 26285 2065
rect 26305 2045 26310 2065
rect 26280 2015 26310 2045
rect 26280 1995 26285 2015
rect 26305 1995 26310 2015
rect 26280 1985 26310 1995
rect 26335 2115 26365 2125
rect 26335 2095 26340 2115
rect 26360 2095 26365 2115
rect 26335 2065 26365 2095
rect 26335 2045 26340 2065
rect 26360 2045 26365 2065
rect 26335 2015 26365 2045
rect 26335 1995 26340 2015
rect 26360 1995 26365 2015
rect 26335 1985 26365 1995
rect 26390 2115 26420 2125
rect 26390 2095 26395 2115
rect 26415 2095 26420 2115
rect 26390 2065 26420 2095
rect 26390 2045 26395 2065
rect 26415 2045 26420 2065
rect 26390 2015 26420 2045
rect 26390 1995 26395 2015
rect 26415 1995 26420 2015
rect 26390 1985 26420 1995
rect 26445 2115 26475 2125
rect 26445 2095 26450 2115
rect 26470 2095 26475 2115
rect 26445 2065 26475 2095
rect 26445 2045 26450 2065
rect 26470 2045 26475 2065
rect 26445 2015 26475 2045
rect 26445 1995 26450 2015
rect 26470 1995 26475 2015
rect 26445 1985 26475 1995
rect 26500 2115 26530 2125
rect 26500 2095 26505 2115
rect 26525 2095 26530 2115
rect 26500 2065 26530 2095
rect 26500 2045 26505 2065
rect 26525 2045 26530 2065
rect 26500 2015 26530 2045
rect 26500 1995 26505 2015
rect 26525 1995 26530 2015
rect 26500 1985 26530 1995
rect 26555 2115 26585 2125
rect 26555 2095 26560 2115
rect 26580 2095 26585 2115
rect 26555 2065 26585 2095
rect 26555 2045 26560 2065
rect 26580 2045 26585 2065
rect 26555 2015 26585 2045
rect 26555 1995 26560 2015
rect 26580 1995 26585 2015
rect 26555 1985 26585 1995
rect 26610 2115 26640 2125
rect 26610 2095 26615 2115
rect 26635 2095 26640 2115
rect 26610 2065 26640 2095
rect 26610 2045 26615 2065
rect 26635 2045 26640 2065
rect 26610 2015 26640 2045
rect 26610 1995 26615 2015
rect 26635 1995 26640 2015
rect 26610 1985 26640 1995
rect 26665 2115 26695 2125
rect 26665 2095 26670 2115
rect 26690 2095 26695 2115
rect 26665 2065 26695 2095
rect 26665 2045 26670 2065
rect 26690 2045 26695 2065
rect 26665 2015 26695 2045
rect 26665 1995 26670 2015
rect 26690 1995 26695 2015
rect 26665 1985 26695 1995
rect 26720 2115 26750 2125
rect 26720 2095 26725 2115
rect 26745 2095 26750 2115
rect 26720 2065 26750 2095
rect 26720 2045 26725 2065
rect 26745 2045 26750 2065
rect 26720 2015 26750 2045
rect 26720 1995 26725 2015
rect 26745 1995 26750 2015
rect 26720 1985 26750 1995
rect 26775 2115 26805 2125
rect 26775 2095 26780 2115
rect 26800 2095 26805 2115
rect 26775 2065 26805 2095
rect 26775 2045 26780 2065
rect 26800 2045 26805 2065
rect 26775 2015 26805 2045
rect 26775 1995 26780 2015
rect 26800 1995 26805 2015
rect 26775 1985 26805 1995
rect 26830 2115 26860 2125
rect 26830 2095 26835 2115
rect 26855 2095 26860 2115
rect 26830 2065 26860 2095
rect 26830 2045 26835 2065
rect 26855 2045 26860 2065
rect 26830 2015 26860 2045
rect 26830 1995 26835 2015
rect 26855 1995 26860 2015
rect 26830 1985 26860 1995
rect 26885 2115 26915 2125
rect 26885 2095 26890 2115
rect 26910 2095 26915 2115
rect 26885 2065 26915 2095
rect 26885 2045 26890 2065
rect 26910 2045 26915 2065
rect 26885 2015 26915 2045
rect 26885 1995 26890 2015
rect 26910 1995 26915 2015
rect 26885 1985 26915 1995
rect 26940 2115 26970 2125
rect 26940 2095 26945 2115
rect 26965 2095 26970 2115
rect 26940 2065 26970 2095
rect 26940 2045 26945 2065
rect 26965 2045 26970 2065
rect 26940 2015 26970 2045
rect 26940 1995 26945 2015
rect 26965 1995 26970 2015
rect 26940 1985 26970 1995
rect 26995 2115 27025 2125
rect 26995 2095 27000 2115
rect 27020 2095 27025 2115
rect 26995 2065 27025 2095
rect 26995 2045 27000 2065
rect 27020 2045 27025 2065
rect 26995 2015 27025 2045
rect 26995 1995 27000 2015
rect 27020 1995 27025 2015
rect 26995 1985 27025 1995
rect 27050 2115 27080 2125
rect 27050 2095 27055 2115
rect 27075 2095 27080 2115
rect 27050 2065 27080 2095
rect 27050 2045 27055 2065
rect 27075 2045 27080 2065
rect 27050 2015 27080 2045
rect 27050 1995 27055 2015
rect 27075 1995 27080 2015
rect 27050 1985 27080 1995
rect 27105 2115 27135 2125
rect 27105 2095 27110 2115
rect 27130 2095 27135 2115
rect 27105 2065 27135 2095
rect 27105 2045 27110 2065
rect 27130 2045 27135 2065
rect 27105 2015 27135 2045
rect 27105 1995 27110 2015
rect 27130 1995 27135 2015
rect 27105 1985 27135 1995
rect 27160 2115 27190 2125
rect 27160 2095 27165 2115
rect 27185 2095 27190 2115
rect 27160 2065 27190 2095
rect 27160 2045 27165 2065
rect 27185 2045 27190 2065
rect 27160 2015 27190 2045
rect 27160 1995 27165 2015
rect 27185 1995 27190 2015
rect 27160 1985 27190 1995
rect 27215 2115 27245 2125
rect 27215 2095 27220 2115
rect 27240 2095 27245 2115
rect 27215 2065 27245 2095
rect 27215 2045 27220 2065
rect 27240 2045 27245 2065
rect 27215 2015 27245 2045
rect 27215 1995 27220 2015
rect 27240 1995 27245 2015
rect 27215 1985 27245 1995
rect 27270 2115 27300 2125
rect 27270 2095 27275 2115
rect 27295 2095 27300 2115
rect 27270 2065 27300 2095
rect 27270 2045 27275 2065
rect 27295 2045 27300 2065
rect 27270 2015 27300 2045
rect 27270 1995 27275 2015
rect 27295 1995 27300 2015
rect 27270 1985 27300 1995
rect 27325 2115 27355 2125
rect 27325 2095 27330 2115
rect 27350 2095 27355 2115
rect 27325 2065 27355 2095
rect 27325 2045 27330 2065
rect 27350 2045 27355 2065
rect 27325 2015 27355 2045
rect 27325 1995 27330 2015
rect 27350 1995 27355 2015
rect 27325 1985 27355 1995
rect 27380 2115 27410 2125
rect 27380 2095 27385 2115
rect 27405 2095 27410 2115
rect 27380 2065 27410 2095
rect 27380 2045 27385 2065
rect 27405 2045 27410 2065
rect 27380 2015 27410 2045
rect 27380 1995 27385 2015
rect 27405 1995 27410 2015
rect 27380 1985 27410 1995
rect 27435 2115 27465 2125
rect 27435 2095 27440 2115
rect 27460 2095 27465 2115
rect 27435 2065 27465 2095
rect 27435 2045 27440 2065
rect 27460 2045 27465 2065
rect 27435 2015 27465 2045
rect 27435 1995 27440 2015
rect 27460 1995 27465 2015
rect 27435 1985 27465 1995
rect 27490 2115 27520 2125
rect 27490 2095 27495 2115
rect 27515 2095 27520 2115
rect 27490 2065 27520 2095
rect 27490 2045 27495 2065
rect 27515 2045 27520 2065
rect 27490 2015 27520 2045
rect 27490 1995 27495 2015
rect 27515 1995 27520 2015
rect 27490 1985 27520 1995
rect 27555 2090 27575 2205
rect 26395 1965 26415 1985
rect 26505 1965 26525 1985
rect 26615 1965 26635 1985
rect 26725 1965 26745 1985
rect 26835 1965 26855 1985
rect 26945 1965 26965 1985
rect 27055 1965 27075 1985
rect 27165 1965 27185 1985
rect 27275 1965 27295 1985
rect 27385 1965 27405 1985
rect 26385 1955 26425 1965
rect 26385 1935 26395 1955
rect 26415 1935 26425 1955
rect 26385 1925 26425 1935
rect 26495 1955 26535 1965
rect 26495 1935 26505 1955
rect 26525 1935 26535 1955
rect 26495 1925 26535 1935
rect 26605 1955 26645 1965
rect 26605 1935 26615 1955
rect 26635 1935 26645 1955
rect 26605 1925 26645 1935
rect 26715 1955 26755 1965
rect 26715 1935 26725 1955
rect 26745 1935 26755 1955
rect 26715 1925 26755 1935
rect 26825 1955 26865 1965
rect 26825 1935 26835 1955
rect 26855 1935 26865 1955
rect 26825 1925 26865 1935
rect 26935 1955 26975 1965
rect 26935 1935 26945 1955
rect 26965 1935 26975 1955
rect 26935 1925 26975 1935
rect 27045 1955 27085 1965
rect 27045 1935 27055 1955
rect 27075 1935 27085 1955
rect 27045 1925 27085 1935
rect 27155 1955 27195 1965
rect 27155 1935 27165 1955
rect 27185 1935 27195 1955
rect 27155 1925 27195 1935
rect 27265 1955 27305 1965
rect 27265 1935 27275 1955
rect 27295 1935 27305 1955
rect 27265 1925 27305 1935
rect 27375 1955 27415 1965
rect 27375 1935 27385 1955
rect 27405 1935 27415 1955
rect 27375 1925 27415 1935
rect 27555 1905 27575 2010
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2755 1885 2775 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2755 1875 2805 1885
rect 2755 1855 2775 1875
rect 2795 1855 2805 1875
rect 2755 1845 2805 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3995 1880 4015 1905
rect 4215 1885 4235 1905
rect 4335 1885 4355 1905
rect 4575 1885 4595 1905
rect 4695 1885 4715 1905
rect 4935 1885 4955 1905
rect 5055 1885 5075 1905
rect 5235 1885 5255 1905
rect 26225 1885 26860 1905
rect 26940 1885 27575 1905
rect 28095 2135 28115 2320
rect 28255 2290 28295 2300
rect 28255 2270 28265 2290
rect 28285 2270 28295 2290
rect 28255 2260 28295 2270
rect 28313 2290 28347 2300
rect 28313 2270 28321 2290
rect 28339 2270 28347 2290
rect 28313 2260 28347 2270
rect 28365 2290 28405 2300
rect 28365 2270 28375 2290
rect 28395 2270 28405 2290
rect 28365 2260 28405 2270
rect 28475 2290 28515 2300
rect 28475 2270 28485 2290
rect 28505 2270 28515 2290
rect 28475 2260 28515 2270
rect 28585 2290 28625 2300
rect 28585 2270 28595 2290
rect 28615 2270 28625 2290
rect 28585 2260 28625 2270
rect 28695 2290 28735 2300
rect 28695 2270 28705 2290
rect 28725 2270 28735 2290
rect 28695 2260 28735 2270
rect 28265 2240 28285 2260
rect 28375 2240 28395 2260
rect 28485 2240 28505 2260
rect 28595 2240 28615 2260
rect 28705 2240 28725 2260
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1880
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1875 4365 1885
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1875 4725 1885
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1875 5085 1885
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5255 1885
rect 5205 1855 5215 1875
rect 5235 1855 5255 1875
rect 5205 1845 5255 1855
rect 28095 1870 28115 2055
rect 28150 2230 28180 2240
rect 28150 2210 28155 2230
rect 28175 2210 28180 2230
rect 28150 2180 28180 2210
rect 28150 2160 28155 2180
rect 28175 2160 28180 2180
rect 28150 2130 28180 2160
rect 28150 2110 28155 2130
rect 28175 2110 28180 2130
rect 28150 2080 28180 2110
rect 28150 2060 28155 2080
rect 28175 2060 28180 2080
rect 28150 2030 28180 2060
rect 28150 2010 28155 2030
rect 28175 2010 28180 2030
rect 28150 1980 28180 2010
rect 28150 1960 28155 1980
rect 28175 1960 28180 1980
rect 28150 1950 28180 1960
rect 28205 2230 28235 2240
rect 28205 2210 28210 2230
rect 28230 2210 28235 2230
rect 28205 2180 28235 2210
rect 28205 2160 28210 2180
rect 28230 2160 28235 2180
rect 28205 2130 28235 2160
rect 28205 2110 28210 2130
rect 28230 2110 28235 2130
rect 28205 2080 28235 2110
rect 28205 2060 28210 2080
rect 28230 2060 28235 2080
rect 28205 2030 28235 2060
rect 28205 2010 28210 2030
rect 28230 2010 28235 2030
rect 28205 1980 28235 2010
rect 28205 1960 28210 1980
rect 28230 1960 28235 1980
rect 28205 1950 28235 1960
rect 28260 2230 28290 2240
rect 28260 2210 28265 2230
rect 28285 2210 28290 2230
rect 28260 2180 28290 2210
rect 28260 2160 28265 2180
rect 28285 2160 28290 2180
rect 28260 2130 28290 2160
rect 28260 2110 28265 2130
rect 28285 2110 28290 2130
rect 28260 2080 28290 2110
rect 28260 2060 28265 2080
rect 28285 2060 28290 2080
rect 28260 2030 28290 2060
rect 28260 2010 28265 2030
rect 28285 2010 28290 2030
rect 28260 1980 28290 2010
rect 28260 1960 28265 1980
rect 28285 1960 28290 1980
rect 28260 1950 28290 1960
rect 28315 2230 28345 2240
rect 28315 2210 28320 2230
rect 28340 2210 28345 2230
rect 28315 2180 28345 2210
rect 28315 2160 28320 2180
rect 28340 2160 28345 2180
rect 28315 2130 28345 2160
rect 28315 2110 28320 2130
rect 28340 2110 28345 2130
rect 28315 2080 28345 2110
rect 28315 2060 28320 2080
rect 28340 2060 28345 2080
rect 28315 2030 28345 2060
rect 28315 2010 28320 2030
rect 28340 2010 28345 2030
rect 28315 1980 28345 2010
rect 28315 1960 28320 1980
rect 28340 1960 28345 1980
rect 28315 1950 28345 1960
rect 28370 2230 28400 2240
rect 28370 2210 28375 2230
rect 28395 2210 28400 2230
rect 28370 2180 28400 2210
rect 28370 2160 28375 2180
rect 28395 2160 28400 2180
rect 28370 2130 28400 2160
rect 28370 2110 28375 2130
rect 28395 2110 28400 2130
rect 28370 2080 28400 2110
rect 28370 2060 28375 2080
rect 28395 2060 28400 2080
rect 28370 2030 28400 2060
rect 28370 2010 28375 2030
rect 28395 2010 28400 2030
rect 28370 1980 28400 2010
rect 28370 1960 28375 1980
rect 28395 1960 28400 1980
rect 28370 1950 28400 1960
rect 28425 2230 28455 2240
rect 28425 2210 28430 2230
rect 28450 2210 28455 2230
rect 28425 2180 28455 2210
rect 28425 2160 28430 2180
rect 28450 2160 28455 2180
rect 28425 2130 28455 2160
rect 28425 2110 28430 2130
rect 28450 2110 28455 2130
rect 28425 2080 28455 2110
rect 28425 2060 28430 2080
rect 28450 2060 28455 2080
rect 28425 2030 28455 2060
rect 28425 2010 28430 2030
rect 28450 2010 28455 2030
rect 28425 1980 28455 2010
rect 28425 1960 28430 1980
rect 28450 1960 28455 1980
rect 28425 1950 28455 1960
rect 28480 2230 28510 2240
rect 28480 2210 28485 2230
rect 28505 2210 28510 2230
rect 28480 2180 28510 2210
rect 28480 2160 28485 2180
rect 28505 2160 28510 2180
rect 28480 2130 28510 2160
rect 28480 2110 28485 2130
rect 28505 2110 28510 2130
rect 28480 2080 28510 2110
rect 28480 2060 28485 2080
rect 28505 2060 28510 2080
rect 28480 2030 28510 2060
rect 28480 2010 28485 2030
rect 28505 2010 28510 2030
rect 28480 1980 28510 2010
rect 28480 1960 28485 1980
rect 28505 1960 28510 1980
rect 28480 1950 28510 1960
rect 28535 2230 28565 2240
rect 28535 2210 28540 2230
rect 28560 2210 28565 2230
rect 28535 2180 28565 2210
rect 28535 2160 28540 2180
rect 28560 2160 28565 2180
rect 28535 2130 28565 2160
rect 28535 2110 28540 2130
rect 28560 2110 28565 2130
rect 28535 2080 28565 2110
rect 28535 2060 28540 2080
rect 28560 2060 28565 2080
rect 28535 2030 28565 2060
rect 28535 2010 28540 2030
rect 28560 2010 28565 2030
rect 28535 1980 28565 2010
rect 28535 1960 28540 1980
rect 28560 1960 28565 1980
rect 28535 1950 28565 1960
rect 28590 2230 28620 2240
rect 28590 2210 28595 2230
rect 28615 2210 28620 2230
rect 28590 2180 28620 2210
rect 28590 2160 28595 2180
rect 28615 2160 28620 2180
rect 28590 2130 28620 2160
rect 28590 2110 28595 2130
rect 28615 2110 28620 2130
rect 28590 2080 28620 2110
rect 28590 2060 28595 2080
rect 28615 2060 28620 2080
rect 28590 2030 28620 2060
rect 28590 2010 28595 2030
rect 28615 2010 28620 2030
rect 28590 1980 28620 2010
rect 28590 1960 28595 1980
rect 28615 1960 28620 1980
rect 28590 1950 28620 1960
rect 28645 2230 28675 2240
rect 28645 2210 28650 2230
rect 28670 2210 28675 2230
rect 28645 2180 28675 2210
rect 28645 2160 28650 2180
rect 28670 2160 28675 2180
rect 28645 2130 28675 2160
rect 28645 2110 28650 2130
rect 28670 2110 28675 2130
rect 28645 2080 28675 2110
rect 28645 2060 28650 2080
rect 28670 2060 28675 2080
rect 28645 2030 28675 2060
rect 28645 2010 28650 2030
rect 28670 2010 28675 2030
rect 28645 1980 28675 2010
rect 28645 1960 28650 1980
rect 28670 1960 28675 1980
rect 28645 1950 28675 1960
rect 28700 2230 28730 2240
rect 28700 2210 28705 2230
rect 28725 2210 28730 2230
rect 28700 2180 28730 2210
rect 28700 2160 28705 2180
rect 28725 2160 28730 2180
rect 28700 2130 28730 2160
rect 28700 2110 28705 2130
rect 28725 2110 28730 2130
rect 28700 2080 28730 2110
rect 28700 2060 28705 2080
rect 28725 2060 28730 2080
rect 28700 2030 28730 2060
rect 28700 2010 28705 2030
rect 28725 2010 28730 2030
rect 28700 1980 28730 2010
rect 28700 1960 28705 1980
rect 28725 1960 28730 1980
rect 28700 1950 28730 1960
rect 28755 2230 28785 2240
rect 28755 2210 28760 2230
rect 28780 2210 28785 2230
rect 28755 2180 28785 2210
rect 28755 2160 28760 2180
rect 28780 2160 28785 2180
rect 28755 2130 28785 2160
rect 28755 2110 28760 2130
rect 28780 2110 28785 2130
rect 28755 2080 28785 2110
rect 28755 2060 28760 2080
rect 28780 2060 28785 2080
rect 28755 2030 28785 2060
rect 28755 2010 28760 2030
rect 28780 2010 28785 2030
rect 28755 1980 28785 2010
rect 28755 1960 28760 1980
rect 28780 1960 28785 1980
rect 28755 1950 28785 1960
rect 28810 2230 28845 2240
rect 28810 2210 28815 2230
rect 28835 2210 28845 2230
rect 28810 2180 28845 2210
rect 28810 2160 28815 2180
rect 28835 2160 28845 2180
rect 28810 2130 28845 2160
rect 28810 2110 28815 2130
rect 28835 2110 28845 2130
rect 28810 2080 28845 2110
rect 28810 2060 28815 2080
rect 28835 2060 28845 2080
rect 28810 2030 28845 2060
rect 28810 2010 28815 2030
rect 28835 2010 28845 2030
rect 28810 1980 28845 2010
rect 28810 1960 28815 1980
rect 28835 1960 28845 1980
rect 28810 1950 28845 1960
rect 28875 2135 28895 2320
rect 28210 1930 28230 1950
rect 28320 1930 28340 1950
rect 28430 1930 28450 1950
rect 28540 1930 28560 1950
rect 28650 1930 28670 1950
rect 28760 1930 28780 1950
rect 28200 1920 28240 1930
rect 28200 1900 28212 1920
rect 28230 1900 28240 1920
rect 28200 1890 28240 1900
rect 28310 1920 28350 1930
rect 28310 1900 28322 1920
rect 28340 1900 28350 1920
rect 28310 1890 28350 1900
rect 28420 1920 28460 1930
rect 28420 1900 28432 1920
rect 28450 1900 28460 1920
rect 28420 1890 28460 1900
rect 28530 1920 28570 1930
rect 28530 1900 28542 1920
rect 28560 1900 28570 1920
rect 28530 1890 28570 1900
rect 28640 1920 28680 1930
rect 28640 1900 28652 1920
rect 28670 1900 28680 1920
rect 28640 1890 28680 1900
rect 28750 1920 28790 1930
rect 28750 1900 28762 1920
rect 28780 1900 28790 1920
rect 28750 1890 28790 1900
rect 28875 1870 28895 2055
rect 28995 2335 29015 2665
rect 29065 2625 29280 2645
rect 29065 2605 29100 2625
rect 29245 2605 29280 2625
rect 29160 2555 29185 2605
rect 28995 1925 29015 2255
rect 29330 2335 29350 2665
rect 29065 1980 29100 1990
rect 29065 1955 29070 1980
rect 29095 1955 29100 1980
rect 29065 1945 29100 1955
rect 29125 1980 29160 1990
rect 29125 1955 29130 1980
rect 29155 1955 29160 1980
rect 29125 1945 29160 1955
rect 29185 1980 29220 1990
rect 29185 1955 29190 1980
rect 29215 1955 29220 1980
rect 29185 1945 29220 1955
rect 29245 1980 29280 1990
rect 29245 1955 29250 1980
rect 29275 1955 29280 1980
rect 29245 1945 29280 1955
rect 29330 1925 29350 2255
rect 28995 1905 29135 1925
rect 29215 1905 29350 1925
rect 28095 1850 28455 1870
rect 28535 1850 28895 1870
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4115 1785 4155 1825
rect 4205 1815 4245 1825
rect 4205 1795 4215 1815
rect 4235 1795 4245 1815
rect 4205 1785 4245 1795
rect 4445 1785 4485 1825
rect 4565 1815 4605 1825
rect 4565 1795 4575 1815
rect 4595 1795 4605 1815
rect 4565 1785 4605 1795
rect 4805 1785 4845 1825
rect 4925 1815 4965 1825
rect 4925 1795 4935 1815
rect 4955 1795 4965 1815
rect 4925 1785 4965 1795
rect 5135 1785 5175 1825
rect 5365 1790 5395 1820
rect 25940 1800 26860 1820
rect 26940 1800 27860 1820
rect 16190 1770 16230 1780
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4205 1755 4245 1765
rect 4205 1735 4215 1755
rect 4235 1735 4245 1755
rect 4205 1725 4245 1735
rect 4445 1755 4485 1765
rect 4445 1735 4455 1755
rect 4475 1735 4485 1755
rect 4445 1725 4485 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1725 4785 1735
rect 5275 1730 5305 1760
rect 16085 1755 16125 1765
rect 16085 1735 16095 1755
rect 16115 1735 16125 1755
rect 16190 1750 16200 1770
rect 16220 1750 16230 1770
rect 16410 1770 16450 1780
rect 16190 1740 16230 1750
rect 16305 1755 16345 1765
rect 16085 1725 16125 1735
rect 3165 1710 3205 1720
rect 2805 1680 2835 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4215 1660 4235 1725
rect 4325 1710 4365 1720
rect 4325 1690 4335 1710
rect 4355 1690 4365 1710
rect 4325 1680 4365 1690
rect 4335 1660 4355 1680
rect 4455 1660 4475 1725
rect 4565 1710 4605 1720
rect 4565 1690 4575 1710
rect 4595 1690 4605 1710
rect 4565 1680 4605 1690
rect 4575 1660 4595 1680
rect 4695 1660 4715 1725
rect 4805 1710 4845 1720
rect 4805 1690 4815 1710
rect 4835 1690 4845 1710
rect 4805 1680 4845 1690
rect 15105 1700 15145 1710
rect 15105 1680 15115 1700
rect 15135 1680 15145 1700
rect 4815 1660 4835 1680
rect 15105 1670 15145 1680
rect 15305 1700 15345 1710
rect 15305 1680 15315 1700
rect 15335 1680 15345 1700
rect 15305 1670 15345 1680
rect 15408 1700 15442 1710
rect 15408 1680 15416 1700
rect 15434 1680 15442 1700
rect 15408 1670 15442 1680
rect 15505 1700 15545 1710
rect 15505 1680 15515 1700
rect 15535 1680 15545 1700
rect 15505 1670 15545 1680
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 4810 1650 4840 1660
rect 15115 1650 15135 1670
rect 15315 1650 15335 1670
rect 15515 1650 15535 1670
rect 16095 1660 16115 1725
rect 16200 1660 16220 1740
rect 16305 1735 16315 1755
rect 16335 1735 16345 1755
rect 16410 1750 16420 1770
rect 16440 1750 16450 1770
rect 16640 1770 16680 1780
rect 16410 1740 16450 1750
rect 16525 1755 16565 1765
rect 16305 1725 16345 1735
rect 16237 1710 16269 1720
rect 16237 1690 16243 1710
rect 16260 1690 16269 1710
rect 16237 1680 16269 1690
rect 16315 1660 16335 1725
rect 16420 1660 16440 1740
rect 16525 1735 16535 1755
rect 16555 1735 16565 1755
rect 16640 1750 16650 1770
rect 16670 1750 16680 1770
rect 17230 1770 17270 1780
rect 16640 1740 16680 1750
rect 17125 1755 17165 1765
rect 16525 1725 16565 1735
rect 16457 1710 16489 1720
rect 16457 1690 16463 1710
rect 16480 1690 16489 1710
rect 16457 1680 16489 1690
rect 16535 1660 16555 1725
rect 16601 1710 16633 1720
rect 16601 1690 16610 1710
rect 16627 1690 16633 1710
rect 16601 1680 16633 1690
rect 16650 1660 16670 1740
rect 17125 1735 17135 1755
rect 17155 1735 17165 1755
rect 17230 1750 17240 1770
rect 17260 1750 17270 1770
rect 17450 1770 17490 1780
rect 17230 1740 17270 1750
rect 17345 1755 17385 1765
rect 17125 1725 17165 1735
rect 16820 1710 16850 1720
rect 16820 1690 16825 1710
rect 16845 1690 16850 1710
rect 16820 1680 16850 1690
rect 16867 1710 16899 1720
rect 16867 1690 16876 1710
rect 16893 1690 16899 1710
rect 16867 1680 16899 1690
rect 16950 1710 16980 1720
rect 16950 1690 16955 1710
rect 16975 1690 16980 1710
rect 16950 1680 16980 1690
rect 16830 1660 16850 1680
rect 16950 1660 16970 1680
rect 17135 1660 17155 1725
rect 17240 1660 17260 1740
rect 17345 1735 17355 1755
rect 17375 1735 17385 1755
rect 17450 1750 17460 1770
rect 17480 1750 17490 1770
rect 17680 1770 17720 1780
rect 17450 1740 17490 1750
rect 17565 1755 17605 1765
rect 17345 1725 17385 1735
rect 17277 1710 17309 1720
rect 17277 1690 17283 1710
rect 17300 1690 17309 1710
rect 17277 1680 17309 1690
rect 17355 1660 17375 1725
rect 17460 1660 17480 1740
rect 17565 1735 17575 1755
rect 17595 1735 17605 1755
rect 17680 1750 17690 1770
rect 17710 1750 17720 1770
rect 17680 1740 17720 1750
rect 17565 1725 17605 1735
rect 17497 1710 17529 1720
rect 17497 1690 17503 1710
rect 17520 1690 17529 1710
rect 17497 1680 17529 1690
rect 17575 1660 17595 1725
rect 17641 1710 17673 1720
rect 17641 1690 17650 1710
rect 17667 1690 17673 1710
rect 17641 1680 17673 1690
rect 17690 1660 17710 1740
rect 18305 1700 18345 1710
rect 18305 1680 18315 1700
rect 18335 1680 18345 1700
rect 18305 1670 18345 1680
rect 18408 1700 18442 1710
rect 18408 1680 18416 1700
rect 18434 1680 18442 1700
rect 18408 1670 18442 1680
rect 18505 1700 18545 1710
rect 18505 1680 18515 1700
rect 18535 1680 18545 1700
rect 18505 1670 18545 1680
rect 18705 1700 18745 1710
rect 18705 1680 18715 1700
rect 18735 1680 18745 1700
rect 18705 1670 18745 1680
rect 25105 1700 25145 1710
rect 25105 1680 25115 1700
rect 25135 1680 25145 1700
rect 25105 1670 25145 1680
rect 25305 1700 25345 1710
rect 25305 1680 25315 1700
rect 25335 1680 25345 1700
rect 25305 1670 25345 1680
rect 25408 1700 25442 1710
rect 25408 1680 25416 1700
rect 25434 1680 25442 1700
rect 25408 1670 25442 1680
rect 25505 1700 25545 1710
rect 25505 1680 25515 1700
rect 25535 1680 25545 1700
rect 25505 1670 25545 1680
rect 15990 1650 16065 1660
rect 4810 1630 4815 1650
rect 4835 1630 4840 1650
rect 4810 1620 4840 1630
rect 14820 1640 14855 1650
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4275 1550 4295 1620
rect 4395 1550 4415 1620
rect 4515 1550 4535 1620
rect 4635 1550 4655 1620
rect 4755 1550 4775 1620
rect 14820 1615 14825 1640
rect 14850 1615 14855 1640
rect 14820 1605 14855 1615
rect 4805 1590 4845 1600
rect 4805 1570 4815 1590
rect 4835 1570 4845 1590
rect 4805 1560 4845 1570
rect 5415 1565 5445 1595
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4265 1540 4305 1550
rect 4265 1520 4275 1540
rect 4295 1520 4305 1540
rect 4265 1510 4305 1520
rect 4385 1540 4425 1550
rect 4385 1520 4395 1540
rect 4415 1520 4425 1540
rect 4385 1510 4425 1520
rect 4505 1540 4545 1550
rect 4505 1520 4515 1540
rect 4535 1520 4545 1540
rect 4505 1510 4545 1520
rect 4625 1540 4665 1550
rect 4625 1520 4635 1540
rect 4655 1520 4665 1540
rect 4625 1510 4665 1520
rect 4745 1540 4785 1550
rect 4745 1520 4755 1540
rect 4775 1520 4785 1540
rect 4745 1510 4785 1520
rect 2925 1495 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1465 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1465 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1465 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1465 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1465 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1465 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 4205 1495 4245 1505
rect 3765 1465 3805 1475
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1465 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1465 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1465 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1465 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1465 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1465 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1465 5085 1475
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1440 2870 1450
rect 2840 1420 2845 1440
rect 2865 1420 2870 1440
rect 2840 1390 2870 1420
rect 2840 1370 2845 1390
rect 2865 1370 2870 1390
rect 2840 1340 2870 1370
rect 2840 1320 2845 1340
rect 2865 1320 2870 1340
rect 2840 1290 2870 1320
rect 2840 1270 2845 1290
rect 2865 1270 2870 1290
rect 2840 1240 2870 1270
rect 2840 1220 2845 1240
rect 2865 1220 2870 1240
rect 2840 1210 2870 1220
rect 3380 1440 3410 1450
rect 3380 1420 3385 1440
rect 3405 1420 3410 1440
rect 3380 1390 3410 1420
rect 3380 1370 3385 1390
rect 3405 1370 3410 1390
rect 3380 1340 3410 1370
rect 3380 1320 3385 1340
rect 3405 1320 3410 1340
rect 3380 1290 3410 1320
rect 3380 1270 3385 1290
rect 3405 1270 3410 1290
rect 3380 1240 3410 1270
rect 3380 1220 3385 1240
rect 3405 1220 3410 1240
rect 3380 1210 3410 1220
rect 3920 1440 3950 1450
rect 3920 1420 3925 1440
rect 3945 1420 3950 1440
rect 3920 1390 3950 1420
rect 3920 1370 3925 1390
rect 3945 1370 3950 1390
rect 3920 1340 3950 1370
rect 3920 1320 3925 1340
rect 3945 1320 3950 1340
rect 3920 1290 3950 1320
rect 3920 1270 3925 1290
rect 3945 1270 3950 1290
rect 3920 1240 3950 1270
rect 3920 1220 3925 1240
rect 3945 1220 3950 1240
rect 3920 1210 3950 1220
rect 4060 1440 4090 1450
rect 4060 1420 4065 1440
rect 4085 1420 4090 1440
rect 4060 1390 4090 1420
rect 4060 1370 4065 1390
rect 4085 1370 4090 1390
rect 4060 1340 4090 1370
rect 4060 1320 4065 1340
rect 4085 1320 4090 1340
rect 4060 1290 4090 1320
rect 4060 1270 4065 1290
rect 4085 1270 4090 1290
rect 4060 1240 4090 1270
rect 4060 1220 4065 1240
rect 4085 1220 4090 1240
rect 4060 1210 4090 1220
rect 4600 1440 4630 1450
rect 4600 1420 4605 1440
rect 4625 1420 4630 1440
rect 4600 1390 4630 1420
rect 4600 1370 4605 1390
rect 4625 1370 4630 1390
rect 4600 1340 4630 1370
rect 4600 1320 4605 1340
rect 4625 1320 4630 1340
rect 4600 1290 4630 1320
rect 4600 1270 4605 1290
rect 4625 1270 4630 1290
rect 4600 1240 4630 1270
rect 4600 1220 4605 1240
rect 4625 1220 4630 1240
rect 4600 1210 4630 1220
rect 5140 1440 5170 1450
rect 5140 1420 5145 1440
rect 5165 1420 5170 1440
rect 5140 1390 5170 1420
rect 5140 1370 5145 1390
rect 5165 1370 5170 1390
rect 14880 1640 14915 1650
rect 14880 1615 14885 1640
rect 14910 1615 14915 1640
rect 14880 1605 14915 1615
rect 14970 1640 15040 1650
rect 14970 1620 14975 1640
rect 14995 1620 15015 1640
rect 15035 1620 15040 1640
rect 14970 1590 15040 1620
rect 14970 1570 14975 1590
rect 14995 1570 15015 1590
rect 15035 1570 15040 1590
rect 14970 1540 15040 1570
rect 14970 1520 14975 1540
rect 14995 1520 15015 1540
rect 15035 1520 15040 1540
rect 14970 1490 15040 1520
rect 14970 1470 14975 1490
rect 14995 1470 15015 1490
rect 15035 1470 15040 1490
rect 14970 1440 15040 1470
rect 14970 1420 14975 1440
rect 14995 1420 15015 1440
rect 15035 1420 15040 1440
rect 14970 1390 15040 1420
rect 5140 1340 5170 1370
rect 5140 1320 5145 1340
rect 5165 1320 5170 1340
rect 5140 1290 5170 1320
rect 5140 1270 5145 1290
rect 5165 1270 5170 1290
rect 5140 1240 5170 1270
rect 5140 1220 5145 1240
rect 5165 1220 5170 1240
rect 5140 1210 5170 1220
rect 14970 1370 14975 1390
rect 14995 1370 15015 1390
rect 15035 1370 15040 1390
rect 14970 1340 15040 1370
rect 14970 1320 14975 1340
rect 14995 1320 15015 1340
rect 15035 1320 15040 1340
rect 14970 1290 15040 1320
rect 14970 1270 14975 1290
rect 14995 1270 15015 1290
rect 15035 1270 15040 1290
rect 14970 1240 15040 1270
rect 14970 1220 14975 1240
rect 14995 1220 15015 1240
rect 15035 1220 15040 1240
rect 3385 1190 3405 1210
rect 4605 1190 4625 1210
rect 14970 1190 15040 1220
rect 3375 1180 3415 1190
rect 3375 1160 3385 1180
rect 3405 1160 3415 1180
rect 3375 1150 3415 1160
rect 3990 1155 4020 1185
rect 4595 1180 4635 1190
rect 4595 1160 4605 1180
rect 4625 1160 4635 1180
rect 4595 1150 4635 1160
rect 14970 1170 14975 1190
rect 14995 1170 15015 1190
rect 15035 1170 15040 1190
rect 14970 1140 15040 1170
rect 2945 1120 2985 1130
rect 2945 1100 2955 1120
rect 2975 1100 2985 1120
rect 2945 1090 2985 1100
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 3985 1120 4025 1130
rect 3985 1100 3995 1120
rect 4015 1100 4025 1120
rect 3985 1090 4025 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2955 1070 2975 1090
rect 3995 1070 4015 1090
rect 2950 1060 2980 1070
rect 2950 1045 2955 1060
rect 2935 1040 2955 1045
rect 2975 1040 2980 1060
rect 2625 1010 2655 1040
rect 2910 1035 2980 1040
rect 2910 1015 2915 1035
rect 2935 1015 2980 1035
rect 2910 1010 2980 1015
rect 2935 1005 2955 1010
rect 2950 990 2955 1005
rect 2975 990 2980 1010
rect 2950 980 2980 990
rect 3990 1060 4020 1070
rect 3990 1040 3995 1060
rect 4015 1040 4020 1060
rect 3990 1010 4020 1040
rect 3990 990 3995 1010
rect 4015 990 4020 1010
rect 3990 980 4020 990
rect 5030 1060 5100 1070
rect 5030 1040 5035 1060
rect 5055 1040 5075 1060
rect 5095 1045 5100 1060
rect 5095 1040 5150 1045
rect 5030 1035 5150 1040
rect 5030 1015 5120 1035
rect 5140 1015 5150 1035
rect 5030 1010 5150 1015
rect 5030 990 5035 1010
rect 5055 990 5075 1010
rect 5095 1005 5150 1010
rect 5095 990 5100 1005
rect 5030 980 5100 990
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 2995 895 3035 905
rect 3175 925 3215 935
rect 3175 905 3185 925
rect 3205 905 3215 925
rect 3175 895 3215 905
rect 3355 925 3395 935
rect 3355 905 3365 925
rect 3385 905 3395 925
rect 3355 895 3395 905
rect 3535 925 3575 935
rect 3535 905 3545 925
rect 3565 905 3575 925
rect 3535 895 3575 905
rect 3715 925 3755 935
rect 3715 905 3725 925
rect 3745 905 3755 925
rect 3715 895 3755 905
rect 3895 925 3935 935
rect 3895 905 3905 925
rect 3925 905 3935 925
rect 3895 895 3935 905
rect 4075 925 4115 935
rect 4075 905 4085 925
rect 4105 905 4115 925
rect 4075 895 4115 905
rect 4255 925 4295 935
rect 4255 905 4265 925
rect 4285 905 4295 925
rect 4255 895 4295 905
rect 4435 925 4475 935
rect 4435 905 4445 925
rect 4465 905 4475 925
rect 4435 895 4475 905
rect 4615 925 4655 935
rect 4615 905 4625 925
rect 4645 905 4655 925
rect 4615 895 4655 905
rect 4795 925 4835 935
rect 4795 905 4805 925
rect 4825 905 4835 925
rect 4795 895 4835 905
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 14855 910 14880 960
rect 14970 1120 14975 1140
rect 14995 1120 15015 1140
rect 15035 1120 15040 1140
rect 14970 1090 15040 1120
rect 14970 1070 14975 1090
rect 14995 1070 15015 1090
rect 15035 1070 15040 1090
rect 14970 1040 15040 1070
rect 14970 1020 14975 1040
rect 14995 1020 15015 1040
rect 15035 1020 15040 1040
rect 14970 990 15040 1020
rect 14970 970 14975 990
rect 14995 970 15015 990
rect 15035 970 15040 990
rect 14970 960 15040 970
rect 15110 1640 15140 1650
rect 15110 1620 15115 1640
rect 15135 1620 15140 1640
rect 15110 1590 15140 1620
rect 15110 1570 15115 1590
rect 15135 1570 15140 1590
rect 15110 1540 15140 1570
rect 15110 1520 15115 1540
rect 15135 1520 15140 1540
rect 15110 1490 15140 1520
rect 15110 1470 15115 1490
rect 15135 1470 15140 1490
rect 15110 1440 15140 1470
rect 15110 1420 15115 1440
rect 15135 1420 15140 1440
rect 15110 1390 15140 1420
rect 15110 1370 15115 1390
rect 15135 1370 15140 1390
rect 15110 1340 15140 1370
rect 15110 1320 15115 1340
rect 15135 1320 15140 1340
rect 15110 1290 15140 1320
rect 15110 1270 15115 1290
rect 15135 1270 15140 1290
rect 15110 1240 15140 1270
rect 15110 1220 15115 1240
rect 15135 1220 15140 1240
rect 15110 1190 15140 1220
rect 15110 1170 15115 1190
rect 15135 1170 15140 1190
rect 15110 1140 15140 1170
rect 15110 1120 15115 1140
rect 15135 1120 15140 1140
rect 15110 1090 15140 1120
rect 15110 1070 15115 1090
rect 15135 1070 15140 1090
rect 15110 1040 15140 1070
rect 15110 1020 15115 1040
rect 15135 1020 15140 1040
rect 15110 990 15140 1020
rect 15110 970 15115 990
rect 15135 970 15140 990
rect 15110 960 15140 970
rect 15210 1640 15240 1650
rect 15210 1620 15215 1640
rect 15235 1620 15240 1640
rect 15210 1590 15240 1620
rect 15210 1570 15215 1590
rect 15235 1570 15240 1590
rect 15210 1540 15240 1570
rect 15210 1520 15215 1540
rect 15235 1520 15240 1540
rect 15210 1490 15240 1520
rect 15210 1470 15215 1490
rect 15235 1470 15240 1490
rect 15210 1440 15240 1470
rect 15210 1420 15215 1440
rect 15235 1420 15240 1440
rect 15210 1390 15240 1420
rect 15210 1370 15215 1390
rect 15235 1370 15240 1390
rect 15210 1340 15240 1370
rect 15210 1320 15215 1340
rect 15235 1320 15240 1340
rect 15210 1290 15240 1320
rect 15210 1270 15215 1290
rect 15235 1270 15240 1290
rect 15210 1240 15240 1270
rect 15210 1220 15215 1240
rect 15235 1220 15240 1240
rect 15210 1190 15240 1220
rect 15210 1170 15215 1190
rect 15235 1170 15240 1190
rect 15210 1140 15240 1170
rect 15210 1120 15215 1140
rect 15235 1120 15240 1140
rect 15210 1090 15240 1120
rect 15210 1070 15215 1090
rect 15235 1070 15240 1090
rect 15210 1040 15240 1070
rect 15210 1020 15215 1040
rect 15235 1020 15240 1040
rect 15210 990 15240 1020
rect 15210 970 15215 990
rect 15235 970 15240 990
rect 15210 960 15240 970
rect 15310 1640 15340 1650
rect 15310 1620 15315 1640
rect 15335 1620 15340 1640
rect 15310 1590 15340 1620
rect 15310 1570 15315 1590
rect 15335 1570 15340 1590
rect 15310 1540 15340 1570
rect 15310 1520 15315 1540
rect 15335 1520 15340 1540
rect 15310 1490 15340 1520
rect 15310 1470 15315 1490
rect 15335 1470 15340 1490
rect 15310 1440 15340 1470
rect 15310 1420 15315 1440
rect 15335 1420 15340 1440
rect 15310 1390 15340 1420
rect 15310 1370 15315 1390
rect 15335 1370 15340 1390
rect 15310 1340 15340 1370
rect 15310 1320 15315 1340
rect 15335 1320 15340 1340
rect 15310 1290 15340 1320
rect 15310 1270 15315 1290
rect 15335 1270 15340 1290
rect 15310 1240 15340 1270
rect 15310 1220 15315 1240
rect 15335 1220 15340 1240
rect 15310 1190 15340 1220
rect 15310 1170 15315 1190
rect 15335 1170 15340 1190
rect 15310 1140 15340 1170
rect 15310 1120 15315 1140
rect 15335 1120 15340 1140
rect 15310 1090 15340 1120
rect 15310 1070 15315 1090
rect 15335 1070 15340 1090
rect 15310 1040 15340 1070
rect 15310 1020 15315 1040
rect 15335 1020 15340 1040
rect 15310 990 15340 1020
rect 15310 970 15315 990
rect 15335 970 15340 990
rect 15310 960 15340 970
rect 15410 1640 15440 1650
rect 15410 1620 15415 1640
rect 15435 1620 15440 1640
rect 15410 1590 15440 1620
rect 15410 1570 15415 1590
rect 15435 1570 15440 1590
rect 15410 1540 15440 1570
rect 15410 1520 15415 1540
rect 15435 1520 15440 1540
rect 15410 1490 15440 1520
rect 15410 1470 15415 1490
rect 15435 1470 15440 1490
rect 15410 1440 15440 1470
rect 15410 1420 15415 1440
rect 15435 1420 15440 1440
rect 15410 1390 15440 1420
rect 15410 1370 15415 1390
rect 15435 1370 15440 1390
rect 15410 1340 15440 1370
rect 15410 1320 15415 1340
rect 15435 1320 15440 1340
rect 15410 1290 15440 1320
rect 15410 1270 15415 1290
rect 15435 1270 15440 1290
rect 15410 1240 15440 1270
rect 15410 1220 15415 1240
rect 15435 1220 15440 1240
rect 15410 1190 15440 1220
rect 15410 1170 15415 1190
rect 15435 1170 15440 1190
rect 15410 1140 15440 1170
rect 15410 1120 15415 1140
rect 15435 1120 15440 1140
rect 15410 1090 15440 1120
rect 15410 1070 15415 1090
rect 15435 1070 15440 1090
rect 15410 1040 15440 1070
rect 15410 1020 15415 1040
rect 15435 1020 15440 1040
rect 15410 990 15440 1020
rect 15410 970 15415 990
rect 15435 970 15440 990
rect 15410 960 15440 970
rect 15510 1640 15540 1650
rect 15510 1620 15515 1640
rect 15535 1620 15540 1640
rect 15510 1590 15540 1620
rect 15510 1570 15515 1590
rect 15535 1570 15540 1590
rect 15510 1540 15540 1570
rect 15510 1520 15515 1540
rect 15535 1520 15540 1540
rect 15510 1490 15540 1520
rect 15510 1470 15515 1490
rect 15535 1470 15540 1490
rect 15510 1440 15540 1470
rect 15510 1420 15515 1440
rect 15535 1420 15540 1440
rect 15510 1390 15540 1420
rect 15510 1370 15515 1390
rect 15535 1370 15540 1390
rect 15510 1340 15540 1370
rect 15510 1320 15515 1340
rect 15535 1320 15540 1340
rect 15510 1290 15540 1320
rect 15510 1270 15515 1290
rect 15535 1270 15540 1290
rect 15510 1240 15540 1270
rect 15510 1220 15515 1240
rect 15535 1220 15540 1240
rect 15510 1190 15540 1220
rect 15510 1170 15515 1190
rect 15535 1170 15540 1190
rect 15510 1140 15540 1170
rect 15510 1120 15515 1140
rect 15535 1120 15540 1140
rect 15510 1090 15540 1120
rect 15510 1070 15515 1090
rect 15535 1070 15540 1090
rect 15510 1040 15540 1070
rect 15510 1020 15515 1040
rect 15535 1020 15540 1040
rect 15510 990 15540 1020
rect 15510 970 15515 990
rect 15535 970 15540 990
rect 15510 960 15540 970
rect 15610 1640 15680 1650
rect 15610 1620 15615 1640
rect 15635 1620 15655 1640
rect 15675 1620 15680 1640
rect 15610 1590 15680 1620
rect 15610 1570 15615 1590
rect 15635 1570 15655 1590
rect 15675 1570 15680 1590
rect 15610 1540 15680 1570
rect 15610 1520 15615 1540
rect 15635 1520 15655 1540
rect 15675 1520 15680 1540
rect 15990 1630 16000 1650
rect 16020 1630 16040 1650
rect 16060 1630 16065 1650
rect 15990 1600 16065 1630
rect 15990 1580 16000 1600
rect 16020 1580 16040 1600
rect 16060 1580 16065 1600
rect 15990 1550 16065 1580
rect 15990 1530 16000 1550
rect 16020 1530 16040 1550
rect 16060 1530 16065 1550
rect 15990 1520 16065 1530
rect 16090 1650 16120 1660
rect 16090 1630 16095 1650
rect 16115 1630 16120 1650
rect 16090 1600 16120 1630
rect 16090 1580 16095 1600
rect 16115 1580 16120 1600
rect 16090 1550 16120 1580
rect 16090 1530 16095 1550
rect 16115 1530 16120 1550
rect 16090 1520 16120 1530
rect 16145 1650 16175 1660
rect 16145 1630 16150 1650
rect 16170 1630 16175 1650
rect 16145 1600 16175 1630
rect 16145 1580 16150 1600
rect 16170 1580 16175 1600
rect 16145 1550 16175 1580
rect 16145 1530 16150 1550
rect 16170 1530 16175 1550
rect 16145 1520 16175 1530
rect 16200 1650 16230 1660
rect 16200 1630 16205 1650
rect 16225 1630 16230 1650
rect 16200 1600 16230 1630
rect 16200 1580 16205 1600
rect 16225 1580 16230 1600
rect 16200 1550 16230 1580
rect 16200 1530 16205 1550
rect 16225 1530 16230 1550
rect 16200 1520 16230 1530
rect 16255 1650 16285 1660
rect 16255 1630 16260 1650
rect 16280 1630 16285 1650
rect 16255 1600 16285 1630
rect 16255 1580 16260 1600
rect 16280 1580 16285 1600
rect 16255 1550 16285 1580
rect 16255 1530 16260 1550
rect 16280 1530 16285 1550
rect 16255 1520 16285 1530
rect 16310 1650 16340 1660
rect 16310 1630 16315 1650
rect 16335 1630 16340 1650
rect 16310 1600 16340 1630
rect 16310 1580 16315 1600
rect 16335 1580 16340 1600
rect 16310 1550 16340 1580
rect 16310 1530 16315 1550
rect 16335 1530 16340 1550
rect 16310 1520 16340 1530
rect 16365 1650 16395 1660
rect 16365 1630 16370 1650
rect 16390 1630 16395 1650
rect 16365 1600 16395 1630
rect 16365 1580 16370 1600
rect 16390 1580 16395 1600
rect 16365 1550 16395 1580
rect 16365 1530 16370 1550
rect 16390 1530 16395 1550
rect 16365 1520 16395 1530
rect 16420 1650 16450 1660
rect 16420 1630 16425 1650
rect 16445 1630 16450 1650
rect 16420 1600 16450 1630
rect 16420 1580 16425 1600
rect 16445 1580 16450 1600
rect 16420 1550 16450 1580
rect 16420 1530 16425 1550
rect 16445 1530 16450 1550
rect 16420 1520 16450 1530
rect 16475 1650 16505 1660
rect 16475 1630 16480 1650
rect 16500 1630 16505 1650
rect 16475 1600 16505 1630
rect 16475 1580 16480 1600
rect 16500 1580 16505 1600
rect 16475 1550 16505 1580
rect 16475 1530 16480 1550
rect 16500 1530 16505 1550
rect 16475 1520 16505 1530
rect 16530 1650 16560 1660
rect 16530 1630 16535 1650
rect 16555 1630 16560 1650
rect 16530 1600 16560 1630
rect 16530 1580 16535 1600
rect 16555 1580 16560 1600
rect 16530 1550 16560 1580
rect 16530 1530 16535 1550
rect 16555 1530 16560 1550
rect 16530 1520 16560 1530
rect 16585 1650 16615 1660
rect 16585 1630 16590 1650
rect 16610 1630 16615 1650
rect 16585 1600 16615 1630
rect 16585 1580 16590 1600
rect 16610 1580 16615 1600
rect 16585 1550 16615 1580
rect 16585 1530 16590 1550
rect 16610 1530 16615 1550
rect 16585 1520 16615 1530
rect 16640 1650 16670 1660
rect 16640 1630 16645 1650
rect 16665 1630 16670 1650
rect 16640 1600 16670 1630
rect 16640 1580 16645 1600
rect 16665 1580 16670 1600
rect 16640 1550 16670 1580
rect 16640 1530 16645 1550
rect 16665 1530 16670 1550
rect 16640 1520 16670 1530
rect 16695 1650 16805 1660
rect 16695 1630 16700 1650
rect 16720 1630 16740 1650
rect 16760 1630 16780 1650
rect 16800 1630 16805 1650
rect 16695 1600 16805 1630
rect 16695 1580 16700 1600
rect 16720 1580 16740 1600
rect 16760 1580 16780 1600
rect 16800 1580 16805 1600
rect 16695 1550 16805 1580
rect 16695 1530 16700 1550
rect 16720 1530 16740 1550
rect 16760 1530 16780 1550
rect 16800 1530 16805 1550
rect 16695 1520 16805 1530
rect 16830 1650 16860 1660
rect 16830 1630 16835 1650
rect 16855 1630 16860 1650
rect 16830 1600 16860 1630
rect 16830 1580 16835 1600
rect 16855 1580 16860 1600
rect 16830 1550 16860 1580
rect 16830 1530 16835 1550
rect 16855 1530 16860 1550
rect 16830 1520 16860 1530
rect 16885 1650 16915 1660
rect 16885 1630 16890 1650
rect 16910 1630 16915 1650
rect 16885 1600 16915 1630
rect 16885 1580 16890 1600
rect 16910 1580 16915 1600
rect 16885 1550 16915 1580
rect 16885 1530 16890 1550
rect 16910 1530 16915 1550
rect 16885 1520 16915 1530
rect 16940 1650 16970 1660
rect 16940 1630 16945 1650
rect 16965 1630 16970 1650
rect 16940 1600 16970 1630
rect 16940 1580 16945 1600
rect 16965 1580 16970 1600
rect 16940 1550 16970 1580
rect 16940 1530 16945 1550
rect 16965 1530 16970 1550
rect 16940 1520 16970 1530
rect 16995 1650 17105 1660
rect 16995 1630 17000 1650
rect 17020 1630 17040 1650
rect 17060 1630 17080 1650
rect 17100 1630 17105 1650
rect 16995 1600 17105 1630
rect 16995 1580 17000 1600
rect 17020 1580 17040 1600
rect 17060 1580 17080 1600
rect 17100 1580 17105 1600
rect 16995 1550 17105 1580
rect 16995 1530 17000 1550
rect 17020 1530 17040 1550
rect 17060 1530 17080 1550
rect 17100 1530 17105 1550
rect 16995 1520 17105 1530
rect 17130 1650 17160 1660
rect 17130 1630 17135 1650
rect 17155 1630 17160 1650
rect 17130 1600 17160 1630
rect 17130 1580 17135 1600
rect 17155 1580 17160 1600
rect 17130 1550 17160 1580
rect 17130 1530 17135 1550
rect 17155 1530 17160 1550
rect 17130 1520 17160 1530
rect 17185 1650 17215 1660
rect 17185 1630 17190 1650
rect 17210 1630 17215 1650
rect 17185 1600 17215 1630
rect 17185 1580 17190 1600
rect 17210 1580 17215 1600
rect 17185 1550 17215 1580
rect 17185 1530 17190 1550
rect 17210 1530 17215 1550
rect 17185 1520 17215 1530
rect 17240 1650 17270 1660
rect 17240 1630 17245 1650
rect 17265 1630 17270 1650
rect 17240 1600 17270 1630
rect 17240 1580 17245 1600
rect 17265 1580 17270 1600
rect 17240 1550 17270 1580
rect 17240 1530 17245 1550
rect 17265 1530 17270 1550
rect 17240 1520 17270 1530
rect 17295 1650 17325 1660
rect 17295 1630 17300 1650
rect 17320 1630 17325 1650
rect 17295 1600 17325 1630
rect 17295 1580 17300 1600
rect 17320 1580 17325 1600
rect 17295 1550 17325 1580
rect 17295 1530 17300 1550
rect 17320 1530 17325 1550
rect 17295 1520 17325 1530
rect 17350 1650 17380 1660
rect 17350 1630 17355 1650
rect 17375 1630 17380 1650
rect 17350 1600 17380 1630
rect 17350 1580 17355 1600
rect 17375 1580 17380 1600
rect 17350 1550 17380 1580
rect 17350 1530 17355 1550
rect 17375 1530 17380 1550
rect 17350 1520 17380 1530
rect 17405 1650 17435 1660
rect 17405 1630 17410 1650
rect 17430 1630 17435 1650
rect 17405 1600 17435 1630
rect 17405 1580 17410 1600
rect 17430 1580 17435 1600
rect 17405 1550 17435 1580
rect 17405 1530 17410 1550
rect 17430 1530 17435 1550
rect 17405 1520 17435 1530
rect 17460 1650 17490 1660
rect 17460 1630 17465 1650
rect 17485 1630 17490 1650
rect 17460 1600 17490 1630
rect 17460 1580 17465 1600
rect 17485 1580 17490 1600
rect 17460 1550 17490 1580
rect 17460 1530 17465 1550
rect 17485 1530 17490 1550
rect 17460 1520 17490 1530
rect 17515 1650 17545 1660
rect 17515 1630 17520 1650
rect 17540 1630 17545 1650
rect 17515 1600 17545 1630
rect 17515 1580 17520 1600
rect 17540 1580 17545 1600
rect 17515 1550 17545 1580
rect 17515 1530 17520 1550
rect 17540 1530 17545 1550
rect 17515 1520 17545 1530
rect 17570 1650 17600 1660
rect 17570 1630 17575 1650
rect 17595 1630 17600 1650
rect 17570 1600 17600 1630
rect 17570 1580 17575 1600
rect 17595 1580 17600 1600
rect 17570 1550 17600 1580
rect 17570 1530 17575 1550
rect 17595 1530 17600 1550
rect 17570 1520 17600 1530
rect 17625 1650 17655 1660
rect 17625 1630 17630 1650
rect 17650 1630 17655 1650
rect 17625 1600 17655 1630
rect 17625 1580 17630 1600
rect 17650 1580 17655 1600
rect 17625 1550 17655 1580
rect 17625 1530 17630 1550
rect 17650 1530 17655 1550
rect 17625 1520 17655 1530
rect 17680 1650 17710 1660
rect 17680 1630 17685 1650
rect 17705 1630 17710 1650
rect 17680 1600 17710 1630
rect 17680 1580 17685 1600
rect 17705 1580 17710 1600
rect 17680 1550 17710 1580
rect 17680 1530 17685 1550
rect 17705 1530 17710 1550
rect 17680 1520 17710 1530
rect 17735 1650 17810 1660
rect 18315 1650 18335 1670
rect 18515 1650 18535 1670
rect 18715 1650 18735 1670
rect 25115 1650 25135 1670
rect 25315 1650 25335 1670
rect 25515 1650 25535 1670
rect 17735 1630 17740 1650
rect 17760 1630 17780 1650
rect 17800 1630 17810 1650
rect 17735 1600 17810 1630
rect 17735 1580 17740 1600
rect 17760 1580 17780 1600
rect 17800 1580 17810 1600
rect 17735 1550 17810 1580
rect 17735 1530 17740 1550
rect 17760 1530 17780 1550
rect 17800 1530 17810 1550
rect 17735 1520 17810 1530
rect 18170 1640 18240 1650
rect 18170 1620 18175 1640
rect 18195 1620 18215 1640
rect 18235 1620 18240 1640
rect 18170 1590 18240 1620
rect 18170 1570 18175 1590
rect 18195 1570 18215 1590
rect 18235 1570 18240 1590
rect 18170 1540 18240 1570
rect 18170 1520 18175 1540
rect 18195 1520 18215 1540
rect 18235 1520 18240 1540
rect 15610 1490 15680 1520
rect 16000 1500 16020 1520
rect 15610 1470 15615 1490
rect 15635 1470 15655 1490
rect 15675 1470 15680 1490
rect 15610 1440 15680 1470
rect 15990 1490 16030 1500
rect 15990 1470 16000 1490
rect 16020 1470 16030 1490
rect 15990 1460 16030 1470
rect 16106 1490 16138 1500
rect 16106 1470 16112 1490
rect 16129 1470 16138 1490
rect 16106 1460 16138 1470
rect 16155 1440 16175 1520
rect 16260 1440 16280 1520
rect 16305 1490 16345 1500
rect 16305 1470 16315 1490
rect 16335 1470 16345 1490
rect 16305 1460 16345 1470
rect 16370 1440 16390 1520
rect 16480 1440 16500 1520
rect 16525 1490 16565 1500
rect 16525 1470 16535 1490
rect 16555 1470 16565 1490
rect 16525 1460 16565 1470
rect 16590 1440 16610 1520
rect 16740 1500 16760 1520
rect 16830 1500 16850 1520
rect 16885 1500 16905 1520
rect 17040 1500 17060 1520
rect 16730 1490 16770 1500
rect 16730 1470 16740 1490
rect 16760 1470 16770 1490
rect 16730 1460 16770 1470
rect 16825 1490 16855 1500
rect 16825 1470 16830 1490
rect 16850 1470 16855 1490
rect 16825 1460 16855 1470
rect 16875 1490 16905 1500
rect 16875 1470 16880 1490
rect 16900 1470 16905 1490
rect 16875 1460 16905 1470
rect 16922 1490 16954 1500
rect 16922 1470 16928 1490
rect 16945 1470 16954 1490
rect 16922 1460 16954 1470
rect 17030 1490 17070 1500
rect 17030 1470 17040 1490
rect 17060 1470 17070 1490
rect 17030 1460 17070 1470
rect 17146 1490 17178 1500
rect 17146 1470 17152 1490
rect 17169 1470 17178 1490
rect 17146 1460 17178 1470
rect 17195 1440 17215 1520
rect 17300 1440 17320 1520
rect 17345 1490 17385 1500
rect 17345 1470 17355 1490
rect 17375 1470 17385 1490
rect 17345 1460 17385 1470
rect 17410 1440 17430 1520
rect 17520 1440 17540 1520
rect 17565 1490 17605 1500
rect 17565 1470 17575 1490
rect 17595 1470 17605 1490
rect 17565 1460 17605 1470
rect 17630 1440 17650 1520
rect 17780 1500 17800 1520
rect 17770 1490 17810 1500
rect 17770 1470 17780 1490
rect 17800 1470 17810 1490
rect 17770 1460 17810 1470
rect 18170 1490 18240 1520
rect 18170 1470 18175 1490
rect 18195 1470 18215 1490
rect 18235 1470 18240 1490
rect 18170 1440 18240 1470
rect 15610 1420 15615 1440
rect 15635 1420 15655 1440
rect 15675 1420 15680 1440
rect 15610 1390 15680 1420
rect 16145 1430 16185 1440
rect 16145 1410 16155 1430
rect 16175 1410 16185 1430
rect 16145 1400 16185 1410
rect 16250 1430 16290 1440
rect 16250 1410 16260 1430
rect 16280 1410 16290 1430
rect 16250 1400 16290 1410
rect 16360 1430 16400 1440
rect 16360 1410 16370 1430
rect 16390 1410 16400 1430
rect 16360 1400 16400 1410
rect 16470 1430 16510 1440
rect 16470 1410 16480 1430
rect 16500 1410 16510 1430
rect 16470 1400 16510 1410
rect 16580 1430 16620 1440
rect 16580 1410 16590 1430
rect 16610 1410 16620 1430
rect 16580 1400 16620 1410
rect 17185 1430 17225 1440
rect 17185 1410 17195 1430
rect 17215 1410 17225 1430
rect 17185 1400 17225 1410
rect 17290 1430 17330 1440
rect 17290 1410 17300 1430
rect 17320 1410 17330 1430
rect 17290 1400 17330 1410
rect 17400 1430 17440 1440
rect 17400 1410 17410 1430
rect 17430 1410 17440 1430
rect 17400 1400 17440 1410
rect 17510 1430 17550 1440
rect 17510 1410 17520 1430
rect 17540 1410 17550 1430
rect 17510 1400 17550 1410
rect 17620 1430 17660 1440
rect 17620 1410 17630 1430
rect 17650 1410 17660 1430
rect 17620 1400 17660 1410
rect 18170 1420 18175 1440
rect 18195 1420 18215 1440
rect 18235 1420 18240 1440
rect 15610 1370 15615 1390
rect 15635 1370 15655 1390
rect 15675 1370 15680 1390
rect 15610 1340 15680 1370
rect 18170 1390 18240 1420
rect 18170 1370 18175 1390
rect 18195 1370 18215 1390
rect 18235 1370 18240 1390
rect 15610 1320 15615 1340
rect 15635 1320 15655 1340
rect 15675 1320 15680 1340
rect 15610 1290 15680 1320
rect 16810 1310 16850 1350
rect 18170 1340 18240 1370
rect 18170 1320 18175 1340
rect 18195 1320 18215 1340
rect 18235 1320 18240 1340
rect 15610 1270 15615 1290
rect 15635 1270 15655 1290
rect 15675 1270 15680 1290
rect 15610 1240 15680 1270
rect 16315 1260 16355 1300
rect 16880 1260 16920 1300
rect 18170 1290 18240 1320
rect 18170 1270 18175 1290
rect 18195 1270 18215 1290
rect 18235 1270 18240 1290
rect 17595 1245 17635 1255
rect 15610 1220 15615 1240
rect 15635 1220 15655 1240
rect 15675 1220 15680 1240
rect 15610 1190 15680 1220
rect 16315 1230 16355 1240
rect 16315 1210 16325 1230
rect 16345 1210 16355 1230
rect 16315 1200 16355 1210
rect 16425 1230 16465 1240
rect 16425 1210 16435 1230
rect 16455 1210 16465 1230
rect 16425 1200 16465 1210
rect 16535 1230 16575 1240
rect 16535 1210 16545 1230
rect 16565 1210 16575 1230
rect 16535 1200 16575 1210
rect 16645 1230 16685 1240
rect 16645 1210 16655 1230
rect 16675 1210 16685 1230
rect 16645 1200 16685 1210
rect 16755 1230 16795 1240
rect 16755 1210 16765 1230
rect 16785 1210 16795 1230
rect 16755 1200 16795 1210
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 16815 1200 16845 1210
rect 16865 1230 16905 1240
rect 16865 1210 16875 1230
rect 16895 1210 16905 1230
rect 16865 1200 16905 1210
rect 16975 1230 17015 1240
rect 16975 1210 16985 1230
rect 17005 1210 17015 1230
rect 16975 1200 17015 1210
rect 17085 1230 17125 1240
rect 17085 1210 17095 1230
rect 17115 1210 17125 1230
rect 17085 1200 17125 1210
rect 17195 1230 17235 1240
rect 17195 1210 17205 1230
rect 17225 1210 17235 1230
rect 17195 1200 17235 1210
rect 17305 1230 17345 1240
rect 17305 1210 17315 1230
rect 17335 1210 17345 1230
rect 17305 1200 17345 1210
rect 17415 1230 17455 1240
rect 17415 1210 17425 1230
rect 17445 1210 17455 1230
rect 17415 1200 17455 1210
rect 17525 1230 17565 1240
rect 17525 1210 17535 1230
rect 17555 1210 17565 1230
rect 17595 1225 17605 1245
rect 17625 1225 17635 1245
rect 17595 1215 17635 1225
rect 18170 1240 18240 1270
rect 18170 1220 18175 1240
rect 18195 1220 18215 1240
rect 18235 1220 18240 1240
rect 17525 1200 17565 1210
rect 15610 1170 15615 1190
rect 15635 1170 15655 1190
rect 15675 1170 15680 1190
rect 16325 1180 16345 1200
rect 16435 1180 16455 1200
rect 16545 1180 16565 1200
rect 16655 1180 16675 1200
rect 16765 1180 16785 1200
rect 16875 1180 16895 1200
rect 16985 1180 17005 1200
rect 17095 1180 17115 1200
rect 17205 1180 17225 1200
rect 17315 1180 17335 1200
rect 17425 1180 17445 1200
rect 17535 1180 17555 1200
rect 18170 1190 18240 1220
rect 15610 1140 15680 1170
rect 15610 1120 15615 1140
rect 15635 1120 15655 1140
rect 15675 1120 15680 1140
rect 15610 1090 15680 1120
rect 15610 1070 15615 1090
rect 15635 1070 15655 1090
rect 15675 1070 15680 1090
rect 15610 1040 15680 1070
rect 15610 1020 15615 1040
rect 15635 1020 15655 1040
rect 15675 1020 15680 1040
rect 15610 990 15680 1020
rect 15610 970 15615 990
rect 15635 970 15655 990
rect 15675 970 15680 990
rect 15610 960 15680 970
rect 16170 1170 16240 1180
rect 16170 1150 16175 1170
rect 16195 1150 16215 1170
rect 16235 1150 16240 1170
rect 16170 1120 16240 1150
rect 16170 1100 16175 1120
rect 16195 1100 16215 1120
rect 16235 1100 16240 1120
rect 16170 1070 16240 1100
rect 16170 1050 16175 1070
rect 16195 1050 16215 1070
rect 16235 1050 16240 1070
rect 16170 1020 16240 1050
rect 16170 1000 16175 1020
rect 16195 1000 16215 1020
rect 16235 1000 16240 1020
rect 16170 970 16240 1000
rect 14975 940 14995 960
rect 15215 940 15235 960
rect 15415 940 15435 960
rect 15655 940 15675 960
rect 16170 950 16175 970
rect 16195 950 16215 970
rect 16235 950 16240 970
rect 16170 940 16240 950
rect 16265 1170 16295 1180
rect 16265 1150 16270 1170
rect 16290 1150 16295 1170
rect 16265 1120 16295 1150
rect 16265 1100 16270 1120
rect 16290 1100 16295 1120
rect 16265 1070 16295 1100
rect 16265 1050 16270 1070
rect 16290 1050 16295 1070
rect 16265 1020 16295 1050
rect 16265 1000 16270 1020
rect 16290 1000 16295 1020
rect 16265 970 16295 1000
rect 16265 950 16270 970
rect 16290 950 16295 970
rect 16265 940 16295 950
rect 16320 1170 16350 1180
rect 16320 1150 16325 1170
rect 16345 1150 16350 1170
rect 16320 1120 16350 1150
rect 16320 1100 16325 1120
rect 16345 1100 16350 1120
rect 16320 1070 16350 1100
rect 16320 1050 16325 1070
rect 16345 1050 16350 1070
rect 16320 1020 16350 1050
rect 16320 1000 16325 1020
rect 16345 1000 16350 1020
rect 16320 970 16350 1000
rect 16320 950 16325 970
rect 16345 950 16350 970
rect 16320 940 16350 950
rect 16375 1170 16405 1180
rect 16375 1150 16380 1170
rect 16400 1150 16405 1170
rect 16375 1120 16405 1150
rect 16375 1100 16380 1120
rect 16400 1100 16405 1120
rect 16375 1070 16405 1100
rect 16375 1050 16380 1070
rect 16400 1050 16405 1070
rect 16375 1020 16405 1050
rect 16375 1000 16380 1020
rect 16400 1000 16405 1020
rect 16375 970 16405 1000
rect 16375 950 16380 970
rect 16400 950 16405 970
rect 16375 940 16405 950
rect 16430 1170 16460 1180
rect 16430 1150 16435 1170
rect 16455 1150 16460 1170
rect 16430 1120 16460 1150
rect 16430 1100 16435 1120
rect 16455 1100 16460 1120
rect 16430 1070 16460 1100
rect 16430 1050 16435 1070
rect 16455 1050 16460 1070
rect 16430 1020 16460 1050
rect 16430 1000 16435 1020
rect 16455 1000 16460 1020
rect 16430 970 16460 1000
rect 16430 950 16435 970
rect 16455 950 16460 970
rect 16430 940 16460 950
rect 16485 1170 16515 1180
rect 16485 1150 16490 1170
rect 16510 1150 16515 1170
rect 16485 1120 16515 1150
rect 16485 1100 16490 1120
rect 16510 1100 16515 1120
rect 16485 1070 16515 1100
rect 16485 1050 16490 1070
rect 16510 1050 16515 1070
rect 16485 1020 16515 1050
rect 16485 1000 16490 1020
rect 16510 1000 16515 1020
rect 16485 970 16515 1000
rect 16485 950 16490 970
rect 16510 950 16515 970
rect 16485 940 16515 950
rect 16540 1170 16570 1180
rect 16540 1150 16545 1170
rect 16565 1150 16570 1170
rect 16540 1120 16570 1150
rect 16540 1100 16545 1120
rect 16565 1100 16570 1120
rect 16540 1070 16570 1100
rect 16540 1050 16545 1070
rect 16565 1050 16570 1070
rect 16540 1020 16570 1050
rect 16540 1000 16545 1020
rect 16565 1000 16570 1020
rect 16540 970 16570 1000
rect 16540 950 16545 970
rect 16565 950 16570 970
rect 16540 940 16570 950
rect 16595 1170 16625 1180
rect 16595 1150 16600 1170
rect 16620 1150 16625 1170
rect 16595 1120 16625 1150
rect 16595 1100 16600 1120
rect 16620 1100 16625 1120
rect 16595 1070 16625 1100
rect 16595 1050 16600 1070
rect 16620 1050 16625 1070
rect 16595 1020 16625 1050
rect 16595 1000 16600 1020
rect 16620 1000 16625 1020
rect 16595 970 16625 1000
rect 16595 950 16600 970
rect 16620 950 16625 970
rect 16595 940 16625 950
rect 16650 1170 16680 1180
rect 16650 1150 16655 1170
rect 16675 1150 16680 1170
rect 16650 1120 16680 1150
rect 16650 1100 16655 1120
rect 16675 1100 16680 1120
rect 16650 1070 16680 1100
rect 16650 1050 16655 1070
rect 16675 1050 16680 1070
rect 16650 1020 16680 1050
rect 16650 1000 16655 1020
rect 16675 1000 16680 1020
rect 16650 970 16680 1000
rect 16650 950 16655 970
rect 16675 950 16680 970
rect 16650 940 16680 950
rect 16705 1170 16735 1180
rect 16705 1150 16710 1170
rect 16730 1150 16735 1170
rect 16705 1120 16735 1150
rect 16705 1100 16710 1120
rect 16730 1100 16735 1120
rect 16705 1070 16735 1100
rect 16705 1050 16710 1070
rect 16730 1050 16735 1070
rect 16705 1020 16735 1050
rect 16705 1000 16710 1020
rect 16730 1000 16735 1020
rect 16705 970 16735 1000
rect 16705 950 16710 970
rect 16730 950 16735 970
rect 16705 940 16735 950
rect 16760 1170 16790 1180
rect 16760 1150 16765 1170
rect 16785 1150 16790 1170
rect 16760 1120 16790 1150
rect 16760 1100 16765 1120
rect 16785 1100 16790 1120
rect 16760 1070 16790 1100
rect 16760 1050 16765 1070
rect 16785 1050 16790 1070
rect 16760 1020 16790 1050
rect 16760 1000 16765 1020
rect 16785 1000 16790 1020
rect 16760 970 16790 1000
rect 16760 950 16765 970
rect 16785 950 16790 970
rect 16760 940 16790 950
rect 16815 1170 16845 1180
rect 16815 1150 16820 1170
rect 16840 1150 16845 1170
rect 16815 1120 16845 1150
rect 16815 1100 16820 1120
rect 16840 1100 16845 1120
rect 16815 1070 16845 1100
rect 16815 1050 16820 1070
rect 16840 1050 16845 1070
rect 16815 1020 16845 1050
rect 16815 1000 16820 1020
rect 16840 1000 16845 1020
rect 16815 970 16845 1000
rect 16815 950 16820 970
rect 16840 950 16845 970
rect 16815 940 16845 950
rect 16870 1170 16900 1180
rect 16870 1150 16875 1170
rect 16895 1150 16900 1170
rect 16870 1120 16900 1150
rect 16870 1100 16875 1120
rect 16895 1100 16900 1120
rect 16870 1070 16900 1100
rect 16870 1050 16875 1070
rect 16895 1050 16900 1070
rect 16870 1020 16900 1050
rect 16870 1000 16875 1020
rect 16895 1000 16900 1020
rect 16870 970 16900 1000
rect 16870 950 16875 970
rect 16895 950 16900 970
rect 16870 940 16900 950
rect 16925 1170 16955 1180
rect 16925 1150 16930 1170
rect 16950 1150 16955 1170
rect 16925 1120 16955 1150
rect 16925 1100 16930 1120
rect 16950 1100 16955 1120
rect 16925 1070 16955 1100
rect 16925 1050 16930 1070
rect 16950 1050 16955 1070
rect 16925 1020 16955 1050
rect 16925 1000 16930 1020
rect 16950 1000 16955 1020
rect 16925 970 16955 1000
rect 16925 950 16930 970
rect 16950 950 16955 970
rect 16925 940 16955 950
rect 16980 1170 17010 1180
rect 16980 1150 16985 1170
rect 17005 1150 17010 1170
rect 16980 1120 17010 1150
rect 16980 1100 16985 1120
rect 17005 1100 17010 1120
rect 16980 1070 17010 1100
rect 16980 1050 16985 1070
rect 17005 1050 17010 1070
rect 16980 1020 17010 1050
rect 16980 1000 16985 1020
rect 17005 1000 17010 1020
rect 16980 970 17010 1000
rect 16980 950 16985 970
rect 17005 950 17010 970
rect 16980 940 17010 950
rect 17035 1170 17065 1180
rect 17035 1150 17040 1170
rect 17060 1150 17065 1170
rect 17035 1120 17065 1150
rect 17035 1100 17040 1120
rect 17060 1100 17065 1120
rect 17035 1070 17065 1100
rect 17035 1050 17040 1070
rect 17060 1050 17065 1070
rect 17035 1020 17065 1050
rect 17035 1000 17040 1020
rect 17060 1000 17065 1020
rect 17035 970 17065 1000
rect 17035 950 17040 970
rect 17060 950 17065 970
rect 17035 940 17065 950
rect 17090 1170 17120 1180
rect 17090 1150 17095 1170
rect 17115 1150 17120 1170
rect 17090 1120 17120 1150
rect 17090 1100 17095 1120
rect 17115 1100 17120 1120
rect 17090 1070 17120 1100
rect 17090 1050 17095 1070
rect 17115 1050 17120 1070
rect 17090 1020 17120 1050
rect 17090 1000 17095 1020
rect 17115 1000 17120 1020
rect 17090 970 17120 1000
rect 17090 950 17095 970
rect 17115 950 17120 970
rect 17090 940 17120 950
rect 17145 1170 17175 1180
rect 17145 1150 17150 1170
rect 17170 1150 17175 1170
rect 17145 1120 17175 1150
rect 17145 1100 17150 1120
rect 17170 1100 17175 1120
rect 17145 1070 17175 1100
rect 17145 1050 17150 1070
rect 17170 1050 17175 1070
rect 17145 1020 17175 1050
rect 17145 1000 17150 1020
rect 17170 1000 17175 1020
rect 17145 970 17175 1000
rect 17145 950 17150 970
rect 17170 950 17175 970
rect 17145 940 17175 950
rect 17200 1170 17230 1180
rect 17200 1150 17205 1170
rect 17225 1150 17230 1170
rect 17200 1120 17230 1150
rect 17200 1100 17205 1120
rect 17225 1100 17230 1120
rect 17200 1070 17230 1100
rect 17200 1050 17205 1070
rect 17225 1050 17230 1070
rect 17200 1020 17230 1050
rect 17200 1000 17205 1020
rect 17225 1000 17230 1020
rect 17200 970 17230 1000
rect 17200 950 17205 970
rect 17225 950 17230 970
rect 17200 940 17230 950
rect 17255 1170 17285 1180
rect 17255 1150 17260 1170
rect 17280 1150 17285 1170
rect 17255 1120 17285 1150
rect 17255 1100 17260 1120
rect 17280 1100 17285 1120
rect 17255 1070 17285 1100
rect 17255 1050 17260 1070
rect 17280 1050 17285 1070
rect 17255 1020 17285 1050
rect 17255 1000 17260 1020
rect 17280 1000 17285 1020
rect 17255 970 17285 1000
rect 17255 950 17260 970
rect 17280 950 17285 970
rect 17255 940 17285 950
rect 17310 1170 17340 1180
rect 17310 1150 17315 1170
rect 17335 1150 17340 1170
rect 17310 1120 17340 1150
rect 17310 1100 17315 1120
rect 17335 1100 17340 1120
rect 17310 1070 17340 1100
rect 17310 1050 17315 1070
rect 17335 1050 17340 1070
rect 17310 1020 17340 1050
rect 17310 1000 17315 1020
rect 17335 1000 17340 1020
rect 17310 970 17340 1000
rect 17310 950 17315 970
rect 17335 950 17340 970
rect 17310 940 17340 950
rect 17365 1170 17395 1180
rect 17365 1150 17370 1170
rect 17390 1150 17395 1170
rect 17365 1120 17395 1150
rect 17365 1100 17370 1120
rect 17390 1100 17395 1120
rect 17365 1070 17395 1100
rect 17365 1050 17370 1070
rect 17390 1050 17395 1070
rect 17365 1020 17395 1050
rect 17365 1000 17370 1020
rect 17390 1000 17395 1020
rect 17365 970 17395 1000
rect 17365 950 17370 970
rect 17390 950 17395 970
rect 17365 940 17395 950
rect 17420 1170 17450 1180
rect 17420 1150 17425 1170
rect 17445 1150 17450 1170
rect 17420 1120 17450 1150
rect 17420 1100 17425 1120
rect 17445 1100 17450 1120
rect 17420 1070 17450 1100
rect 17420 1050 17425 1070
rect 17445 1050 17450 1070
rect 17420 1020 17450 1050
rect 17420 1000 17425 1020
rect 17445 1000 17450 1020
rect 17420 970 17450 1000
rect 17420 950 17425 970
rect 17445 950 17450 970
rect 17420 940 17450 950
rect 17475 1170 17505 1180
rect 17475 1150 17480 1170
rect 17500 1150 17505 1170
rect 17475 1120 17505 1150
rect 17475 1100 17480 1120
rect 17500 1100 17505 1120
rect 17475 1070 17505 1100
rect 17475 1050 17480 1070
rect 17500 1050 17505 1070
rect 17475 1020 17505 1050
rect 17475 1000 17480 1020
rect 17500 1000 17505 1020
rect 17475 970 17505 1000
rect 17475 950 17480 970
rect 17500 950 17505 970
rect 17475 940 17505 950
rect 17530 1170 17560 1180
rect 17530 1150 17535 1170
rect 17555 1150 17560 1170
rect 17530 1120 17560 1150
rect 17530 1100 17535 1120
rect 17555 1100 17560 1120
rect 17530 1070 17560 1100
rect 17530 1050 17535 1070
rect 17555 1050 17560 1070
rect 17530 1020 17560 1050
rect 17530 1000 17535 1020
rect 17555 1000 17560 1020
rect 17530 970 17560 1000
rect 17530 950 17535 970
rect 17555 950 17560 970
rect 17530 940 17560 950
rect 17585 1170 17655 1180
rect 17585 1150 17590 1170
rect 17610 1150 17630 1170
rect 17650 1150 17655 1170
rect 17585 1120 17655 1150
rect 17585 1100 17590 1120
rect 17610 1100 17630 1120
rect 17650 1100 17655 1120
rect 17585 1070 17655 1100
rect 17585 1050 17590 1070
rect 17610 1050 17630 1070
rect 17650 1050 17655 1070
rect 17585 1020 17655 1050
rect 17585 1000 17590 1020
rect 17610 1000 17630 1020
rect 17650 1000 17655 1020
rect 17585 970 17655 1000
rect 17585 950 17590 970
rect 17610 950 17630 970
rect 17650 950 17655 970
rect 18170 1170 18175 1190
rect 18195 1170 18215 1190
rect 18235 1170 18240 1190
rect 18170 1140 18240 1170
rect 18170 1120 18175 1140
rect 18195 1120 18215 1140
rect 18235 1120 18240 1140
rect 18170 1090 18240 1120
rect 18170 1070 18175 1090
rect 18195 1070 18215 1090
rect 18235 1070 18240 1090
rect 18170 1040 18240 1070
rect 18170 1020 18175 1040
rect 18195 1020 18215 1040
rect 18235 1020 18240 1040
rect 18170 990 18240 1020
rect 18170 970 18175 990
rect 18195 970 18215 990
rect 18235 970 18240 990
rect 18170 960 18240 970
rect 18310 1640 18340 1650
rect 18310 1620 18315 1640
rect 18335 1620 18340 1640
rect 18310 1590 18340 1620
rect 18310 1570 18315 1590
rect 18335 1570 18340 1590
rect 18310 1540 18340 1570
rect 18310 1520 18315 1540
rect 18335 1520 18340 1540
rect 18310 1490 18340 1520
rect 18310 1470 18315 1490
rect 18335 1470 18340 1490
rect 18310 1440 18340 1470
rect 18310 1420 18315 1440
rect 18335 1420 18340 1440
rect 18310 1390 18340 1420
rect 18310 1370 18315 1390
rect 18335 1370 18340 1390
rect 18310 1340 18340 1370
rect 18310 1320 18315 1340
rect 18335 1320 18340 1340
rect 18310 1290 18340 1320
rect 18310 1270 18315 1290
rect 18335 1270 18340 1290
rect 18310 1240 18340 1270
rect 18310 1220 18315 1240
rect 18335 1220 18340 1240
rect 18310 1190 18340 1220
rect 18310 1170 18315 1190
rect 18335 1170 18340 1190
rect 18310 1140 18340 1170
rect 18310 1120 18315 1140
rect 18335 1120 18340 1140
rect 18310 1090 18340 1120
rect 18310 1070 18315 1090
rect 18335 1070 18340 1090
rect 18310 1040 18340 1070
rect 18310 1020 18315 1040
rect 18335 1020 18340 1040
rect 18310 990 18340 1020
rect 18310 970 18315 990
rect 18335 970 18340 990
rect 18310 960 18340 970
rect 18410 1640 18440 1650
rect 18410 1620 18415 1640
rect 18435 1620 18440 1640
rect 18410 1590 18440 1620
rect 18410 1570 18415 1590
rect 18435 1570 18440 1590
rect 18410 1540 18440 1570
rect 18410 1520 18415 1540
rect 18435 1520 18440 1540
rect 18410 1490 18440 1520
rect 18410 1470 18415 1490
rect 18435 1470 18440 1490
rect 18410 1440 18440 1470
rect 18410 1420 18415 1440
rect 18435 1420 18440 1440
rect 18410 1390 18440 1420
rect 18410 1370 18415 1390
rect 18435 1370 18440 1390
rect 18410 1340 18440 1370
rect 18410 1320 18415 1340
rect 18435 1320 18440 1340
rect 18410 1290 18440 1320
rect 18410 1270 18415 1290
rect 18435 1270 18440 1290
rect 18410 1240 18440 1270
rect 18410 1220 18415 1240
rect 18435 1220 18440 1240
rect 18410 1190 18440 1220
rect 18410 1170 18415 1190
rect 18435 1170 18440 1190
rect 18410 1140 18440 1170
rect 18410 1120 18415 1140
rect 18435 1120 18440 1140
rect 18410 1090 18440 1120
rect 18410 1070 18415 1090
rect 18435 1070 18440 1090
rect 18410 1040 18440 1070
rect 18410 1020 18415 1040
rect 18435 1020 18440 1040
rect 18410 990 18440 1020
rect 18410 970 18415 990
rect 18435 970 18440 990
rect 18410 960 18440 970
rect 18510 1640 18540 1650
rect 18510 1620 18515 1640
rect 18535 1620 18540 1640
rect 18510 1590 18540 1620
rect 18510 1570 18515 1590
rect 18535 1570 18540 1590
rect 18510 1540 18540 1570
rect 18510 1520 18515 1540
rect 18535 1520 18540 1540
rect 18510 1490 18540 1520
rect 18510 1470 18515 1490
rect 18535 1470 18540 1490
rect 18510 1440 18540 1470
rect 18510 1420 18515 1440
rect 18535 1420 18540 1440
rect 18510 1390 18540 1420
rect 18510 1370 18515 1390
rect 18535 1370 18540 1390
rect 18510 1340 18540 1370
rect 18510 1320 18515 1340
rect 18535 1320 18540 1340
rect 18510 1290 18540 1320
rect 18510 1270 18515 1290
rect 18535 1270 18540 1290
rect 18510 1240 18540 1270
rect 18510 1220 18515 1240
rect 18535 1220 18540 1240
rect 18510 1190 18540 1220
rect 18510 1170 18515 1190
rect 18535 1170 18540 1190
rect 18510 1140 18540 1170
rect 18510 1120 18515 1140
rect 18535 1120 18540 1140
rect 18510 1090 18540 1120
rect 18510 1070 18515 1090
rect 18535 1070 18540 1090
rect 18510 1040 18540 1070
rect 18510 1020 18515 1040
rect 18535 1020 18540 1040
rect 18510 990 18540 1020
rect 18510 970 18515 990
rect 18535 970 18540 990
rect 18510 960 18540 970
rect 18610 1640 18640 1650
rect 18610 1620 18615 1640
rect 18635 1620 18640 1640
rect 18610 1590 18640 1620
rect 18610 1570 18615 1590
rect 18635 1570 18640 1590
rect 18610 1540 18640 1570
rect 18610 1520 18615 1540
rect 18635 1520 18640 1540
rect 18610 1490 18640 1520
rect 18610 1470 18615 1490
rect 18635 1470 18640 1490
rect 18610 1440 18640 1470
rect 18610 1420 18615 1440
rect 18635 1420 18640 1440
rect 18610 1390 18640 1420
rect 18610 1370 18615 1390
rect 18635 1370 18640 1390
rect 18610 1340 18640 1370
rect 18610 1320 18615 1340
rect 18635 1320 18640 1340
rect 18610 1290 18640 1320
rect 18610 1270 18615 1290
rect 18635 1270 18640 1290
rect 18610 1240 18640 1270
rect 18610 1220 18615 1240
rect 18635 1220 18640 1240
rect 18610 1190 18640 1220
rect 18610 1170 18615 1190
rect 18635 1170 18640 1190
rect 18610 1140 18640 1170
rect 18610 1120 18615 1140
rect 18635 1120 18640 1140
rect 18610 1090 18640 1120
rect 18610 1070 18615 1090
rect 18635 1070 18640 1090
rect 18610 1040 18640 1070
rect 18610 1020 18615 1040
rect 18635 1020 18640 1040
rect 18610 990 18640 1020
rect 18610 970 18615 990
rect 18635 970 18640 990
rect 18610 960 18640 970
rect 18710 1640 18740 1650
rect 18710 1620 18715 1640
rect 18735 1620 18740 1640
rect 18710 1590 18740 1620
rect 18710 1570 18715 1590
rect 18735 1570 18740 1590
rect 18710 1540 18740 1570
rect 18710 1520 18715 1540
rect 18735 1520 18740 1540
rect 18710 1490 18740 1520
rect 18710 1470 18715 1490
rect 18735 1470 18740 1490
rect 18710 1440 18740 1470
rect 18710 1420 18715 1440
rect 18735 1420 18740 1440
rect 18710 1390 18740 1420
rect 18710 1370 18715 1390
rect 18735 1370 18740 1390
rect 18710 1340 18740 1370
rect 18710 1320 18715 1340
rect 18735 1320 18740 1340
rect 18710 1290 18740 1320
rect 18710 1270 18715 1290
rect 18735 1270 18740 1290
rect 18710 1240 18740 1270
rect 18710 1220 18715 1240
rect 18735 1220 18740 1240
rect 18710 1190 18740 1220
rect 18710 1170 18715 1190
rect 18735 1170 18740 1190
rect 18710 1140 18740 1170
rect 18710 1120 18715 1140
rect 18735 1120 18740 1140
rect 18710 1090 18740 1120
rect 18710 1070 18715 1090
rect 18735 1070 18740 1090
rect 18710 1040 18740 1070
rect 18710 1020 18715 1040
rect 18735 1020 18740 1040
rect 18710 990 18740 1020
rect 18710 970 18715 990
rect 18735 970 18740 990
rect 18710 960 18740 970
rect 18810 1640 18880 1650
rect 18810 1620 18815 1640
rect 18835 1620 18855 1640
rect 18875 1620 18880 1640
rect 18810 1590 18880 1620
rect 18810 1570 18815 1590
rect 18835 1570 18855 1590
rect 18875 1570 18880 1590
rect 18810 1540 18880 1570
rect 18810 1520 18815 1540
rect 18835 1520 18855 1540
rect 18875 1520 18880 1540
rect 18810 1490 18880 1520
rect 18810 1470 18815 1490
rect 18835 1470 18855 1490
rect 18875 1470 18880 1490
rect 18810 1440 18880 1470
rect 18810 1420 18815 1440
rect 18835 1420 18855 1440
rect 18875 1420 18880 1440
rect 18810 1390 18880 1420
rect 18810 1370 18815 1390
rect 18835 1370 18855 1390
rect 18875 1370 18880 1390
rect 18935 1640 18970 1650
rect 18935 1615 18940 1640
rect 18965 1615 18970 1640
rect 18935 1605 18970 1615
rect 18995 1640 19030 1650
rect 18995 1615 19000 1640
rect 19025 1615 19030 1640
rect 18995 1605 19030 1615
rect 24820 1640 24855 1650
rect 24820 1615 24825 1640
rect 24850 1615 24855 1640
rect 24820 1605 24855 1615
rect 24880 1640 24915 1650
rect 24880 1615 24885 1640
rect 24910 1615 24915 1640
rect 24880 1605 24915 1615
rect 24970 1640 25040 1650
rect 24970 1620 24975 1640
rect 24995 1620 25015 1640
rect 25035 1620 25040 1640
rect 24970 1590 25040 1620
rect 24970 1570 24975 1590
rect 24995 1570 25015 1590
rect 25035 1570 25040 1590
rect 24970 1540 25040 1570
rect 24970 1520 24975 1540
rect 24995 1520 25015 1540
rect 25035 1520 25040 1540
rect 24970 1490 25040 1520
rect 24970 1470 24975 1490
rect 24995 1470 25015 1490
rect 25035 1470 25040 1490
rect 24970 1440 25040 1470
rect 24970 1420 24975 1440
rect 24995 1420 25015 1440
rect 25035 1420 25040 1440
rect 24970 1390 25040 1420
rect 18810 1340 18880 1370
rect 18810 1320 18815 1340
rect 18835 1320 18855 1340
rect 18875 1320 18880 1340
rect 18810 1290 18880 1320
rect 18810 1270 18815 1290
rect 18835 1270 18855 1290
rect 18875 1270 18880 1290
rect 18810 1240 18880 1270
rect 18810 1220 18815 1240
rect 18835 1220 18855 1240
rect 18875 1220 18880 1240
rect 18810 1190 18880 1220
rect 18810 1170 18815 1190
rect 18835 1170 18855 1190
rect 18875 1170 18880 1190
rect 18810 1140 18880 1170
rect 18810 1120 18815 1140
rect 18835 1120 18855 1140
rect 18875 1120 18880 1140
rect 24970 1370 24975 1390
rect 24995 1370 25015 1390
rect 25035 1370 25040 1390
rect 24970 1340 25040 1370
rect 24970 1320 24975 1340
rect 24995 1320 25015 1340
rect 25035 1320 25040 1340
rect 24970 1290 25040 1320
rect 24970 1270 24975 1290
rect 24995 1270 25015 1290
rect 25035 1270 25040 1290
rect 24970 1240 25040 1270
rect 24970 1220 24975 1240
rect 24995 1220 25015 1240
rect 25035 1220 25040 1240
rect 24970 1190 25040 1220
rect 24970 1170 24975 1190
rect 24995 1170 25015 1190
rect 25035 1170 25040 1190
rect 24970 1140 25040 1170
rect 18810 1090 18880 1120
rect 18810 1070 18815 1090
rect 18835 1070 18855 1090
rect 18875 1070 18880 1090
rect 18810 1040 18880 1070
rect 18810 1020 18815 1040
rect 18835 1020 18855 1040
rect 18875 1020 18880 1040
rect 18810 990 18880 1020
rect 18810 970 18815 990
rect 18835 970 18855 990
rect 18875 970 18880 990
rect 18810 960 18880 970
rect 17585 940 17655 950
rect 18175 940 18195 960
rect 18415 940 18435 960
rect 18615 940 18635 960
rect 18855 940 18875 960
rect 14965 930 15005 940
rect 14965 910 14975 930
rect 14995 910 15005 930
rect 4975 895 5015 905
rect 14965 900 15005 910
rect 15205 930 15245 940
rect 15205 910 15215 930
rect 15235 910 15245 930
rect 15205 900 15245 910
rect 15405 930 15445 940
rect 15405 910 15415 930
rect 15435 910 15445 930
rect 15405 900 15445 910
rect 15645 930 15685 940
rect 15645 910 15655 930
rect 15675 910 15685 930
rect 16175 920 16195 940
rect 16270 920 16290 940
rect 16380 920 16400 940
rect 16490 920 16510 940
rect 16600 920 16620 940
rect 16710 920 16730 940
rect 16820 920 16840 940
rect 16930 920 16950 940
rect 17040 920 17060 940
rect 17150 920 17170 940
rect 17260 920 17280 940
rect 17370 920 17390 940
rect 17480 920 17500 940
rect 17630 920 17650 940
rect 18165 930 18205 940
rect 15645 900 15685 910
rect 16165 910 16205 920
rect 3005 875 3025 895
rect 3185 875 3205 895
rect 3365 875 3385 895
rect 3545 875 3565 895
rect 3725 875 3745 895
rect 3905 875 3925 895
rect 4085 875 4105 895
rect 4265 875 4285 895
rect 4445 875 4465 895
rect 4625 875 4645 895
rect 4805 875 4825 895
rect 4985 875 5005 895
rect 16165 890 16175 910
rect 16195 890 16205 910
rect 16165 880 16205 890
rect 16260 910 16300 920
rect 16260 890 16270 910
rect 16290 890 16300 910
rect 16260 880 16300 890
rect 16370 910 16410 920
rect 16370 890 16380 910
rect 16400 890 16410 910
rect 16370 880 16410 890
rect 16480 910 16520 920
rect 16480 890 16490 910
rect 16510 890 16520 910
rect 16480 880 16520 890
rect 16590 910 16630 920
rect 16590 890 16600 910
rect 16620 890 16630 910
rect 16590 880 16630 890
rect 16700 910 16740 920
rect 16700 890 16710 910
rect 16730 890 16740 910
rect 16700 880 16740 890
rect 16810 910 16850 920
rect 16810 890 16820 910
rect 16840 890 16850 910
rect 16810 880 16850 890
rect 16920 910 16960 920
rect 16920 890 16930 910
rect 16950 890 16960 910
rect 16920 880 16960 890
rect 17030 910 17070 920
rect 17030 890 17040 910
rect 17060 890 17070 910
rect 17030 880 17070 890
rect 17140 910 17180 920
rect 17140 890 17150 910
rect 17170 890 17180 910
rect 17140 880 17180 890
rect 17250 910 17290 920
rect 17250 890 17260 910
rect 17280 890 17290 910
rect 17250 880 17290 890
rect 17360 910 17400 920
rect 17360 890 17370 910
rect 17390 890 17400 910
rect 17360 880 17400 890
rect 17470 910 17510 920
rect 17470 890 17480 910
rect 17500 890 17510 910
rect 17470 880 17510 890
rect 17620 910 17660 920
rect 17620 890 17630 910
rect 17650 890 17660 910
rect 18165 910 18175 930
rect 18195 910 18205 930
rect 18165 900 18205 910
rect 18405 930 18445 940
rect 18405 910 18415 930
rect 18435 910 18445 930
rect 18405 900 18445 910
rect 18605 930 18645 940
rect 18605 910 18615 930
rect 18635 910 18645 930
rect 18605 900 18645 910
rect 18845 930 18885 940
rect 18845 910 18855 930
rect 18875 910 18885 930
rect 18970 910 18995 960
rect 24855 910 24880 960
rect 24970 1120 24975 1140
rect 24995 1120 25015 1140
rect 25035 1120 25040 1140
rect 24970 1090 25040 1120
rect 24970 1070 24975 1090
rect 24995 1070 25015 1090
rect 25035 1070 25040 1090
rect 24970 1040 25040 1070
rect 24970 1020 24975 1040
rect 24995 1020 25015 1040
rect 25035 1020 25040 1040
rect 24970 990 25040 1020
rect 24970 970 24975 990
rect 24995 970 25015 990
rect 25035 970 25040 990
rect 24970 960 25040 970
rect 25110 1640 25140 1650
rect 25110 1620 25115 1640
rect 25135 1620 25140 1640
rect 25110 1590 25140 1620
rect 25110 1570 25115 1590
rect 25135 1570 25140 1590
rect 25110 1540 25140 1570
rect 25110 1520 25115 1540
rect 25135 1520 25140 1540
rect 25110 1490 25140 1520
rect 25110 1470 25115 1490
rect 25135 1470 25140 1490
rect 25110 1440 25140 1470
rect 25110 1420 25115 1440
rect 25135 1420 25140 1440
rect 25110 1390 25140 1420
rect 25110 1370 25115 1390
rect 25135 1370 25140 1390
rect 25110 1340 25140 1370
rect 25110 1320 25115 1340
rect 25135 1320 25140 1340
rect 25110 1290 25140 1320
rect 25110 1270 25115 1290
rect 25135 1270 25140 1290
rect 25110 1240 25140 1270
rect 25110 1220 25115 1240
rect 25135 1220 25140 1240
rect 25110 1190 25140 1220
rect 25110 1170 25115 1190
rect 25135 1170 25140 1190
rect 25110 1140 25140 1170
rect 25110 1120 25115 1140
rect 25135 1120 25140 1140
rect 25110 1090 25140 1120
rect 25110 1070 25115 1090
rect 25135 1070 25140 1090
rect 25110 1040 25140 1070
rect 25110 1020 25115 1040
rect 25135 1020 25140 1040
rect 25110 990 25140 1020
rect 25110 970 25115 990
rect 25135 970 25140 990
rect 25110 960 25140 970
rect 25210 1640 25240 1650
rect 25210 1620 25215 1640
rect 25235 1620 25240 1640
rect 25210 1590 25240 1620
rect 25210 1570 25215 1590
rect 25235 1570 25240 1590
rect 25210 1540 25240 1570
rect 25210 1520 25215 1540
rect 25235 1520 25240 1540
rect 25210 1490 25240 1520
rect 25210 1470 25215 1490
rect 25235 1470 25240 1490
rect 25210 1440 25240 1470
rect 25210 1420 25215 1440
rect 25235 1420 25240 1440
rect 25210 1390 25240 1420
rect 25210 1370 25215 1390
rect 25235 1370 25240 1390
rect 25210 1340 25240 1370
rect 25210 1320 25215 1340
rect 25235 1320 25240 1340
rect 25210 1290 25240 1320
rect 25210 1270 25215 1290
rect 25235 1270 25240 1290
rect 25210 1240 25240 1270
rect 25210 1220 25215 1240
rect 25235 1220 25240 1240
rect 25210 1190 25240 1220
rect 25210 1170 25215 1190
rect 25235 1170 25240 1190
rect 25210 1140 25240 1170
rect 25210 1120 25215 1140
rect 25235 1120 25240 1140
rect 25210 1090 25240 1120
rect 25210 1070 25215 1090
rect 25235 1070 25240 1090
rect 25210 1040 25240 1070
rect 25210 1020 25215 1040
rect 25235 1020 25240 1040
rect 25210 990 25240 1020
rect 25210 970 25215 990
rect 25235 970 25240 990
rect 25210 960 25240 970
rect 25310 1640 25340 1650
rect 25310 1620 25315 1640
rect 25335 1620 25340 1640
rect 25310 1590 25340 1620
rect 25310 1570 25315 1590
rect 25335 1570 25340 1590
rect 25310 1540 25340 1570
rect 25310 1520 25315 1540
rect 25335 1520 25340 1540
rect 25310 1490 25340 1520
rect 25310 1470 25315 1490
rect 25335 1470 25340 1490
rect 25310 1440 25340 1470
rect 25310 1420 25315 1440
rect 25335 1420 25340 1440
rect 25310 1390 25340 1420
rect 25310 1370 25315 1390
rect 25335 1370 25340 1390
rect 25310 1340 25340 1370
rect 25310 1320 25315 1340
rect 25335 1320 25340 1340
rect 25310 1290 25340 1320
rect 25310 1270 25315 1290
rect 25335 1270 25340 1290
rect 25310 1240 25340 1270
rect 25310 1220 25315 1240
rect 25335 1220 25340 1240
rect 25310 1190 25340 1220
rect 25310 1170 25315 1190
rect 25335 1170 25340 1190
rect 25310 1140 25340 1170
rect 25310 1120 25315 1140
rect 25335 1120 25340 1140
rect 25310 1090 25340 1120
rect 25310 1070 25315 1090
rect 25335 1070 25340 1090
rect 25310 1040 25340 1070
rect 25310 1020 25315 1040
rect 25335 1020 25340 1040
rect 25310 990 25340 1020
rect 25310 970 25315 990
rect 25335 970 25340 990
rect 25310 960 25340 970
rect 25410 1640 25440 1650
rect 25410 1620 25415 1640
rect 25435 1620 25440 1640
rect 25410 1590 25440 1620
rect 25410 1570 25415 1590
rect 25435 1570 25440 1590
rect 25410 1540 25440 1570
rect 25410 1520 25415 1540
rect 25435 1520 25440 1540
rect 25410 1490 25440 1520
rect 25410 1470 25415 1490
rect 25435 1470 25440 1490
rect 25410 1440 25440 1470
rect 25410 1420 25415 1440
rect 25435 1420 25440 1440
rect 25410 1390 25440 1420
rect 25410 1370 25415 1390
rect 25435 1370 25440 1390
rect 25410 1340 25440 1370
rect 25410 1320 25415 1340
rect 25435 1320 25440 1340
rect 25410 1290 25440 1320
rect 25410 1270 25415 1290
rect 25435 1270 25440 1290
rect 25410 1240 25440 1270
rect 25410 1220 25415 1240
rect 25435 1220 25440 1240
rect 25410 1190 25440 1220
rect 25410 1170 25415 1190
rect 25435 1170 25440 1190
rect 25410 1140 25440 1170
rect 25410 1120 25415 1140
rect 25435 1120 25440 1140
rect 25410 1090 25440 1120
rect 25410 1070 25415 1090
rect 25435 1070 25440 1090
rect 25410 1040 25440 1070
rect 25410 1020 25415 1040
rect 25435 1020 25440 1040
rect 25410 990 25440 1020
rect 25410 970 25415 990
rect 25435 970 25440 990
rect 25410 960 25440 970
rect 25510 1640 25540 1650
rect 25510 1620 25515 1640
rect 25535 1620 25540 1640
rect 25510 1590 25540 1620
rect 25510 1570 25515 1590
rect 25535 1570 25540 1590
rect 25510 1540 25540 1570
rect 25510 1520 25515 1540
rect 25535 1520 25540 1540
rect 25510 1490 25540 1520
rect 25510 1470 25515 1490
rect 25535 1470 25540 1490
rect 25510 1440 25540 1470
rect 25510 1420 25515 1440
rect 25535 1420 25540 1440
rect 25510 1390 25540 1420
rect 25510 1370 25515 1390
rect 25535 1370 25540 1390
rect 25510 1340 25540 1370
rect 25510 1320 25515 1340
rect 25535 1320 25540 1340
rect 25510 1290 25540 1320
rect 25510 1270 25515 1290
rect 25535 1270 25540 1290
rect 25510 1240 25540 1270
rect 25510 1220 25515 1240
rect 25535 1220 25540 1240
rect 25510 1190 25540 1220
rect 25510 1170 25515 1190
rect 25535 1170 25540 1190
rect 25510 1140 25540 1170
rect 25510 1120 25515 1140
rect 25535 1120 25540 1140
rect 25510 1090 25540 1120
rect 25510 1070 25515 1090
rect 25535 1070 25540 1090
rect 25510 1040 25540 1070
rect 25510 1020 25515 1040
rect 25535 1020 25540 1040
rect 25510 990 25540 1020
rect 25510 970 25515 990
rect 25535 970 25540 990
rect 25510 960 25540 970
rect 25610 1640 25680 1650
rect 25610 1620 25615 1640
rect 25635 1620 25655 1640
rect 25675 1620 25680 1640
rect 25610 1590 25680 1620
rect 25610 1570 25615 1590
rect 25635 1570 25655 1590
rect 25675 1570 25680 1590
rect 25610 1540 25680 1570
rect 25610 1520 25615 1540
rect 25635 1520 25655 1540
rect 25675 1520 25680 1540
rect 25610 1490 25680 1520
rect 25610 1470 25615 1490
rect 25635 1470 25655 1490
rect 25675 1470 25680 1490
rect 25610 1440 25680 1470
rect 25610 1420 25615 1440
rect 25635 1420 25655 1440
rect 25675 1420 25680 1440
rect 25610 1390 25680 1420
rect 25610 1370 25615 1390
rect 25635 1370 25655 1390
rect 25675 1370 25680 1390
rect 25610 1340 25680 1370
rect 25940 1630 25960 1800
rect 26190 1770 26230 1780
rect 26085 1755 26125 1765
rect 26085 1735 26095 1755
rect 26115 1735 26125 1755
rect 26190 1750 26200 1770
rect 26220 1750 26230 1770
rect 26410 1770 26450 1780
rect 26190 1740 26230 1750
rect 26305 1755 26345 1765
rect 26085 1725 26125 1735
rect 26095 1660 26115 1725
rect 26200 1660 26220 1740
rect 26305 1735 26315 1755
rect 26335 1735 26345 1755
rect 26410 1750 26420 1770
rect 26440 1750 26450 1770
rect 26640 1770 26680 1780
rect 26410 1740 26450 1750
rect 26525 1755 26565 1765
rect 26305 1725 26345 1735
rect 26237 1710 26269 1720
rect 26237 1690 26243 1710
rect 26260 1690 26269 1710
rect 26237 1680 26269 1690
rect 26315 1660 26335 1725
rect 26420 1660 26440 1740
rect 26525 1735 26535 1755
rect 26555 1735 26565 1755
rect 26640 1750 26650 1770
rect 26670 1750 26680 1770
rect 27230 1770 27270 1780
rect 26640 1740 26680 1750
rect 27125 1755 27165 1765
rect 26525 1725 26565 1735
rect 26457 1710 26489 1720
rect 26457 1690 26463 1710
rect 26480 1690 26489 1710
rect 26457 1680 26489 1690
rect 26535 1660 26555 1725
rect 26601 1710 26633 1720
rect 26601 1690 26610 1710
rect 26627 1690 26633 1710
rect 26601 1680 26633 1690
rect 26650 1660 26670 1740
rect 27125 1735 27135 1755
rect 27155 1735 27165 1755
rect 27230 1750 27240 1770
rect 27260 1750 27270 1770
rect 27450 1770 27490 1780
rect 27230 1740 27270 1750
rect 27345 1755 27385 1765
rect 27125 1725 27165 1735
rect 26820 1710 26850 1720
rect 26820 1690 26825 1710
rect 26845 1690 26850 1710
rect 26820 1680 26850 1690
rect 26867 1710 26899 1720
rect 26867 1690 26876 1710
rect 26893 1690 26899 1710
rect 26867 1680 26899 1690
rect 26950 1710 26980 1720
rect 26950 1690 26955 1710
rect 26975 1690 26980 1710
rect 26950 1680 26980 1690
rect 26830 1660 26850 1680
rect 26950 1660 26970 1680
rect 27135 1660 27155 1725
rect 27240 1660 27260 1740
rect 27345 1735 27355 1755
rect 27375 1735 27385 1755
rect 27450 1750 27460 1770
rect 27480 1750 27490 1770
rect 27680 1770 27720 1780
rect 27450 1740 27490 1750
rect 27565 1755 27605 1765
rect 27345 1725 27385 1735
rect 27277 1710 27309 1720
rect 27277 1690 27283 1710
rect 27300 1690 27309 1710
rect 27277 1680 27309 1690
rect 27355 1660 27375 1725
rect 27460 1660 27480 1740
rect 27565 1735 27575 1755
rect 27595 1735 27605 1755
rect 27680 1750 27690 1770
rect 27710 1750 27720 1770
rect 27680 1740 27720 1750
rect 27565 1725 27605 1735
rect 27497 1710 27529 1720
rect 27497 1690 27503 1710
rect 27520 1690 27529 1710
rect 27497 1680 27529 1690
rect 27575 1660 27595 1725
rect 27641 1710 27673 1720
rect 27641 1690 27650 1710
rect 27667 1690 27673 1710
rect 27641 1680 27673 1690
rect 27690 1660 27710 1740
rect 25940 1380 25960 1550
rect 26035 1650 26065 1660
rect 26035 1630 26040 1650
rect 26060 1630 26065 1650
rect 26035 1600 26065 1630
rect 26035 1580 26040 1600
rect 26060 1580 26065 1600
rect 26035 1550 26065 1580
rect 26035 1530 26040 1550
rect 26060 1530 26065 1550
rect 26035 1520 26065 1530
rect 26090 1650 26120 1660
rect 26090 1630 26095 1650
rect 26115 1630 26120 1650
rect 26090 1600 26120 1630
rect 26090 1580 26095 1600
rect 26115 1580 26120 1600
rect 26090 1550 26120 1580
rect 26090 1530 26095 1550
rect 26115 1530 26120 1550
rect 26090 1520 26120 1530
rect 26145 1650 26175 1660
rect 26145 1630 26150 1650
rect 26170 1630 26175 1650
rect 26145 1600 26175 1630
rect 26145 1580 26150 1600
rect 26170 1580 26175 1600
rect 26145 1550 26175 1580
rect 26145 1530 26150 1550
rect 26170 1530 26175 1550
rect 26145 1520 26175 1530
rect 26200 1650 26230 1660
rect 26200 1630 26205 1650
rect 26225 1630 26230 1650
rect 26200 1600 26230 1630
rect 26200 1580 26205 1600
rect 26225 1580 26230 1600
rect 26200 1550 26230 1580
rect 26200 1530 26205 1550
rect 26225 1530 26230 1550
rect 26200 1520 26230 1530
rect 26255 1650 26285 1660
rect 26255 1630 26260 1650
rect 26280 1630 26285 1650
rect 26255 1600 26285 1630
rect 26255 1580 26260 1600
rect 26280 1580 26285 1600
rect 26255 1550 26285 1580
rect 26255 1530 26260 1550
rect 26280 1530 26285 1550
rect 26255 1520 26285 1530
rect 26310 1650 26340 1660
rect 26310 1630 26315 1650
rect 26335 1630 26340 1650
rect 26310 1600 26340 1630
rect 26310 1580 26315 1600
rect 26335 1580 26340 1600
rect 26310 1550 26340 1580
rect 26310 1530 26315 1550
rect 26335 1530 26340 1550
rect 26310 1520 26340 1530
rect 26365 1650 26395 1660
rect 26365 1630 26370 1650
rect 26390 1630 26395 1650
rect 26365 1600 26395 1630
rect 26365 1580 26370 1600
rect 26390 1580 26395 1600
rect 26365 1550 26395 1580
rect 26365 1530 26370 1550
rect 26390 1530 26395 1550
rect 26365 1520 26395 1530
rect 26420 1650 26450 1660
rect 26420 1630 26425 1650
rect 26445 1630 26450 1650
rect 26420 1600 26450 1630
rect 26420 1580 26425 1600
rect 26445 1580 26450 1600
rect 26420 1550 26450 1580
rect 26420 1530 26425 1550
rect 26445 1530 26450 1550
rect 26420 1520 26450 1530
rect 26475 1650 26505 1660
rect 26475 1630 26480 1650
rect 26500 1630 26505 1650
rect 26475 1600 26505 1630
rect 26475 1580 26480 1600
rect 26500 1580 26505 1600
rect 26475 1550 26505 1580
rect 26475 1530 26480 1550
rect 26500 1530 26505 1550
rect 26475 1520 26505 1530
rect 26530 1650 26560 1660
rect 26530 1630 26535 1650
rect 26555 1630 26560 1650
rect 26530 1600 26560 1630
rect 26530 1580 26535 1600
rect 26555 1580 26560 1600
rect 26530 1550 26560 1580
rect 26530 1530 26535 1550
rect 26555 1530 26560 1550
rect 26530 1520 26560 1530
rect 26585 1650 26615 1660
rect 26585 1630 26590 1650
rect 26610 1630 26615 1650
rect 26585 1600 26615 1630
rect 26585 1580 26590 1600
rect 26610 1580 26615 1600
rect 26585 1550 26615 1580
rect 26585 1530 26590 1550
rect 26610 1530 26615 1550
rect 26585 1520 26615 1530
rect 26640 1650 26670 1660
rect 26640 1630 26645 1650
rect 26665 1630 26670 1650
rect 26640 1600 26670 1630
rect 26640 1580 26645 1600
rect 26665 1580 26670 1600
rect 26640 1550 26670 1580
rect 26640 1530 26645 1550
rect 26665 1530 26670 1550
rect 26640 1520 26670 1530
rect 26695 1650 26805 1660
rect 26695 1630 26700 1650
rect 26720 1630 26740 1650
rect 26760 1630 26780 1650
rect 26800 1630 26805 1650
rect 26695 1600 26805 1630
rect 26695 1580 26700 1600
rect 26720 1580 26740 1600
rect 26760 1580 26780 1600
rect 26800 1580 26805 1600
rect 26695 1550 26805 1580
rect 26695 1530 26700 1550
rect 26720 1530 26740 1550
rect 26760 1530 26780 1550
rect 26800 1530 26805 1550
rect 26695 1520 26805 1530
rect 26830 1650 26860 1660
rect 26830 1630 26835 1650
rect 26855 1630 26860 1650
rect 26830 1600 26860 1630
rect 26830 1580 26835 1600
rect 26855 1580 26860 1600
rect 26830 1550 26860 1580
rect 26830 1530 26835 1550
rect 26855 1530 26860 1550
rect 26830 1520 26860 1530
rect 26885 1650 26915 1660
rect 26885 1630 26890 1650
rect 26910 1630 26915 1650
rect 26885 1600 26915 1630
rect 26885 1580 26890 1600
rect 26910 1580 26915 1600
rect 26885 1550 26915 1580
rect 26885 1530 26890 1550
rect 26910 1530 26915 1550
rect 26885 1520 26915 1530
rect 26940 1650 26970 1660
rect 26940 1630 26945 1650
rect 26965 1630 26970 1650
rect 26940 1600 26970 1630
rect 26940 1580 26945 1600
rect 26965 1580 26970 1600
rect 26940 1550 26970 1580
rect 26940 1530 26945 1550
rect 26965 1530 26970 1550
rect 26940 1520 26970 1530
rect 26995 1650 27105 1660
rect 26995 1630 27000 1650
rect 27020 1630 27040 1650
rect 27060 1630 27080 1650
rect 27100 1630 27105 1650
rect 26995 1600 27105 1630
rect 26995 1580 27000 1600
rect 27020 1580 27040 1600
rect 27060 1580 27080 1600
rect 27100 1580 27105 1600
rect 26995 1550 27105 1580
rect 26995 1530 27000 1550
rect 27020 1530 27040 1550
rect 27060 1530 27080 1550
rect 27100 1530 27105 1550
rect 26995 1520 27105 1530
rect 27130 1650 27160 1660
rect 27130 1630 27135 1650
rect 27155 1630 27160 1650
rect 27130 1600 27160 1630
rect 27130 1580 27135 1600
rect 27155 1580 27160 1600
rect 27130 1550 27160 1580
rect 27130 1530 27135 1550
rect 27155 1530 27160 1550
rect 27130 1520 27160 1530
rect 27185 1650 27215 1660
rect 27185 1630 27190 1650
rect 27210 1630 27215 1650
rect 27185 1600 27215 1630
rect 27185 1580 27190 1600
rect 27210 1580 27215 1600
rect 27185 1550 27215 1580
rect 27185 1530 27190 1550
rect 27210 1530 27215 1550
rect 27185 1520 27215 1530
rect 27240 1650 27270 1660
rect 27240 1630 27245 1650
rect 27265 1630 27270 1650
rect 27240 1600 27270 1630
rect 27240 1580 27245 1600
rect 27265 1580 27270 1600
rect 27240 1550 27270 1580
rect 27240 1530 27245 1550
rect 27265 1530 27270 1550
rect 27240 1520 27270 1530
rect 27295 1650 27325 1660
rect 27295 1630 27300 1650
rect 27320 1630 27325 1650
rect 27295 1600 27325 1630
rect 27295 1580 27300 1600
rect 27320 1580 27325 1600
rect 27295 1550 27325 1580
rect 27295 1530 27300 1550
rect 27320 1530 27325 1550
rect 27295 1520 27325 1530
rect 27350 1650 27380 1660
rect 27350 1630 27355 1650
rect 27375 1630 27380 1650
rect 27350 1600 27380 1630
rect 27350 1580 27355 1600
rect 27375 1580 27380 1600
rect 27350 1550 27380 1580
rect 27350 1530 27355 1550
rect 27375 1530 27380 1550
rect 27350 1520 27380 1530
rect 27405 1650 27435 1660
rect 27405 1630 27410 1650
rect 27430 1630 27435 1650
rect 27405 1600 27435 1630
rect 27405 1580 27410 1600
rect 27430 1580 27435 1600
rect 27405 1550 27435 1580
rect 27405 1530 27410 1550
rect 27430 1530 27435 1550
rect 27405 1520 27435 1530
rect 27460 1650 27490 1660
rect 27460 1630 27465 1650
rect 27485 1630 27490 1650
rect 27460 1600 27490 1630
rect 27460 1580 27465 1600
rect 27485 1580 27490 1600
rect 27460 1550 27490 1580
rect 27460 1530 27465 1550
rect 27485 1530 27490 1550
rect 27460 1520 27490 1530
rect 27515 1650 27545 1660
rect 27515 1630 27520 1650
rect 27540 1630 27545 1650
rect 27515 1600 27545 1630
rect 27515 1580 27520 1600
rect 27540 1580 27545 1600
rect 27515 1550 27545 1580
rect 27515 1530 27520 1550
rect 27540 1530 27545 1550
rect 27515 1520 27545 1530
rect 27570 1650 27600 1660
rect 27570 1630 27575 1650
rect 27595 1630 27600 1650
rect 27570 1600 27600 1630
rect 27570 1580 27575 1600
rect 27595 1580 27600 1600
rect 27570 1550 27600 1580
rect 27570 1530 27575 1550
rect 27595 1530 27600 1550
rect 27570 1520 27600 1530
rect 27625 1650 27655 1660
rect 27625 1630 27630 1650
rect 27650 1630 27655 1650
rect 27625 1600 27655 1630
rect 27625 1580 27630 1600
rect 27650 1580 27655 1600
rect 27625 1550 27655 1580
rect 27625 1530 27630 1550
rect 27650 1530 27655 1550
rect 27625 1520 27655 1530
rect 27680 1650 27710 1660
rect 27680 1630 27685 1650
rect 27705 1630 27710 1650
rect 27680 1600 27710 1630
rect 27680 1580 27685 1600
rect 27705 1580 27710 1600
rect 27680 1550 27710 1580
rect 27680 1530 27685 1550
rect 27705 1530 27710 1550
rect 27680 1520 27710 1530
rect 27735 1650 27765 1660
rect 27735 1630 27740 1650
rect 27760 1630 27765 1650
rect 27735 1600 27765 1630
rect 27735 1580 27740 1600
rect 27760 1580 27765 1600
rect 27735 1550 27765 1580
rect 27735 1530 27740 1550
rect 27760 1530 27765 1550
rect 27735 1520 27765 1530
rect 27840 1630 27860 1800
rect 26106 1490 26138 1500
rect 26106 1470 26112 1490
rect 26129 1470 26138 1490
rect 26106 1460 26138 1470
rect 26155 1440 26175 1520
rect 26260 1440 26280 1520
rect 26305 1490 26345 1500
rect 26305 1470 26315 1490
rect 26335 1470 26345 1490
rect 26305 1460 26345 1470
rect 26370 1440 26390 1520
rect 26480 1440 26500 1520
rect 26525 1490 26565 1500
rect 26525 1470 26535 1490
rect 26555 1470 26565 1490
rect 26525 1460 26565 1470
rect 26590 1440 26610 1520
rect 26740 1500 26760 1520
rect 26830 1500 26850 1520
rect 26885 1500 26905 1520
rect 27040 1500 27060 1520
rect 26730 1490 26770 1500
rect 26730 1470 26740 1490
rect 26760 1470 26770 1490
rect 26730 1460 26770 1470
rect 26825 1490 26855 1500
rect 26825 1470 26830 1490
rect 26850 1470 26855 1490
rect 26825 1460 26855 1470
rect 26875 1490 26905 1500
rect 26875 1470 26880 1490
rect 26900 1470 26905 1490
rect 26875 1460 26905 1470
rect 26922 1490 26954 1500
rect 26922 1470 26928 1490
rect 26945 1470 26954 1490
rect 26922 1460 26954 1470
rect 27030 1490 27070 1500
rect 27030 1470 27040 1490
rect 27060 1470 27070 1490
rect 27030 1460 27070 1470
rect 27146 1490 27178 1500
rect 27146 1470 27152 1490
rect 27169 1470 27178 1490
rect 27146 1460 27178 1470
rect 27195 1440 27215 1520
rect 27300 1440 27320 1520
rect 27345 1490 27385 1500
rect 27345 1470 27355 1490
rect 27375 1470 27385 1490
rect 27345 1460 27385 1470
rect 27410 1440 27430 1520
rect 27520 1440 27540 1520
rect 27565 1490 27605 1500
rect 27565 1470 27575 1490
rect 27595 1470 27605 1490
rect 27565 1460 27605 1470
rect 27630 1440 27650 1520
rect 26145 1430 26185 1440
rect 26145 1410 26155 1430
rect 26175 1410 26185 1430
rect 26145 1400 26185 1410
rect 26250 1430 26290 1440
rect 26250 1410 26260 1430
rect 26280 1410 26290 1430
rect 26250 1400 26290 1410
rect 26360 1430 26400 1440
rect 26360 1410 26370 1430
rect 26390 1410 26400 1430
rect 26360 1400 26400 1410
rect 26470 1430 26510 1440
rect 26470 1410 26480 1430
rect 26500 1410 26510 1430
rect 26470 1400 26510 1410
rect 26580 1430 26620 1440
rect 26580 1410 26590 1430
rect 26610 1410 26620 1430
rect 26580 1400 26620 1410
rect 27185 1430 27225 1440
rect 27185 1410 27195 1430
rect 27215 1410 27225 1430
rect 27185 1400 27225 1410
rect 27290 1430 27330 1440
rect 27290 1410 27300 1430
rect 27320 1410 27330 1430
rect 27290 1400 27330 1410
rect 27400 1430 27440 1440
rect 27400 1410 27410 1430
rect 27430 1410 27440 1430
rect 27400 1400 27440 1410
rect 27510 1430 27550 1440
rect 27510 1410 27520 1430
rect 27540 1410 27550 1430
rect 27510 1400 27550 1410
rect 27620 1430 27660 1440
rect 27620 1410 27630 1430
rect 27650 1410 27660 1430
rect 27620 1400 27660 1410
rect 27840 1380 27860 1550
rect 25940 1360 26860 1380
rect 26940 1360 27860 1380
rect 28155 1730 28485 1750
rect 28565 1730 28895 1750
rect 25610 1320 25615 1340
rect 25635 1320 25655 1340
rect 25675 1320 25680 1340
rect 25610 1290 25680 1320
rect 25610 1270 25615 1290
rect 25635 1270 25655 1290
rect 25675 1270 25680 1290
rect 25610 1240 25680 1270
rect 25610 1220 25615 1240
rect 25635 1220 25655 1240
rect 25675 1220 25680 1240
rect 25610 1190 25680 1220
rect 28155 1345 28175 1730
rect 28305 1700 28345 1710
rect 28305 1680 28315 1700
rect 28335 1680 28345 1700
rect 28305 1670 28345 1680
rect 28408 1700 28442 1710
rect 28408 1680 28416 1700
rect 28434 1680 28442 1700
rect 28408 1670 28442 1680
rect 28505 1700 28545 1710
rect 28505 1680 28515 1700
rect 28535 1680 28545 1700
rect 28505 1670 28545 1680
rect 28705 1700 28745 1710
rect 28705 1680 28715 1700
rect 28735 1680 28745 1700
rect 28705 1670 28745 1680
rect 28315 1650 28335 1670
rect 28515 1650 28535 1670
rect 28715 1650 28735 1670
rect 26315 1195 26355 1200
rect 26880 1195 26920 1200
rect 25610 1170 25615 1190
rect 25635 1170 25655 1190
rect 25675 1170 25680 1190
rect 25610 1140 25680 1170
rect 25610 1120 25615 1140
rect 25635 1120 25655 1140
rect 25675 1120 25680 1140
rect 25610 1090 25680 1120
rect 25610 1070 25615 1090
rect 25635 1070 25655 1090
rect 25675 1070 25680 1090
rect 25610 1040 25680 1070
rect 25610 1020 25615 1040
rect 25635 1020 25655 1040
rect 25675 1020 25680 1040
rect 25610 990 25680 1020
rect 25610 970 25615 990
rect 25635 970 25655 990
rect 25675 970 25680 990
rect 25610 960 25680 970
rect 26155 1175 26845 1195
rect 26925 1175 27675 1195
rect 26155 980 26175 1175
rect 26315 1160 26355 1175
rect 26880 1160 26920 1175
rect 27595 1145 27635 1155
rect 26315 1130 26355 1140
rect 26315 1110 26325 1130
rect 26345 1110 26355 1130
rect 26315 1100 26355 1110
rect 26425 1130 26465 1140
rect 26425 1110 26435 1130
rect 26455 1110 26465 1130
rect 26425 1100 26465 1110
rect 26535 1130 26575 1140
rect 26535 1110 26545 1130
rect 26565 1110 26575 1130
rect 26535 1100 26575 1110
rect 26645 1130 26685 1140
rect 26645 1110 26655 1130
rect 26675 1110 26685 1130
rect 26645 1100 26685 1110
rect 26755 1130 26795 1140
rect 26755 1110 26765 1130
rect 26785 1110 26795 1130
rect 26755 1100 26795 1110
rect 26815 1130 26845 1140
rect 26815 1110 26820 1130
rect 26840 1110 26845 1130
rect 26815 1100 26845 1110
rect 26865 1130 26905 1140
rect 26865 1110 26875 1130
rect 26895 1110 26905 1130
rect 26865 1100 26905 1110
rect 26975 1130 27015 1140
rect 26975 1110 26985 1130
rect 27005 1110 27015 1130
rect 26975 1100 27015 1110
rect 27085 1130 27125 1140
rect 27085 1110 27095 1130
rect 27115 1110 27125 1130
rect 27085 1100 27125 1110
rect 27195 1130 27235 1140
rect 27195 1110 27205 1130
rect 27225 1110 27235 1130
rect 27195 1100 27235 1110
rect 27305 1130 27345 1140
rect 27305 1110 27315 1130
rect 27335 1110 27345 1130
rect 27305 1100 27345 1110
rect 27415 1130 27455 1140
rect 27415 1110 27425 1130
rect 27445 1110 27455 1130
rect 27415 1100 27455 1110
rect 27525 1130 27565 1140
rect 27525 1110 27535 1130
rect 27555 1110 27565 1130
rect 27595 1125 27605 1145
rect 27625 1125 27635 1145
rect 27595 1115 27635 1125
rect 27525 1100 27565 1110
rect 26325 1080 26345 1100
rect 26435 1080 26455 1100
rect 26545 1080 26565 1100
rect 26655 1080 26675 1100
rect 26765 1080 26785 1100
rect 26875 1080 26895 1100
rect 26985 1080 27005 1100
rect 27095 1080 27115 1100
rect 27205 1080 27225 1100
rect 27315 1080 27335 1100
rect 27425 1080 27445 1100
rect 27535 1080 27555 1100
rect 24975 940 24995 960
rect 25215 940 25235 960
rect 25415 940 25435 960
rect 25655 940 25675 960
rect 24965 930 25005 940
rect 24965 910 24975 930
rect 24995 910 25005 930
rect 18845 900 18885 910
rect 24965 900 25005 910
rect 25205 930 25245 940
rect 25205 910 25215 930
rect 25235 910 25245 930
rect 25205 900 25245 910
rect 25405 930 25445 940
rect 25405 910 25415 930
rect 25435 910 25445 930
rect 25405 900 25445 910
rect 25645 930 25685 940
rect 25645 910 25655 930
rect 25675 910 25685 930
rect 25645 900 25685 910
rect 17620 880 17660 890
rect 2960 865 3030 875
rect 2960 845 2965 865
rect 2985 845 3005 865
rect 3025 845 3030 865
rect 2960 815 3030 845
rect 2960 795 2965 815
rect 2985 795 3005 815
rect 3025 795 3030 815
rect 2960 785 3030 795
rect 3090 865 3120 875
rect 3090 845 3095 865
rect 3115 845 3120 865
rect 3090 815 3120 845
rect 3090 795 3095 815
rect 3115 795 3120 815
rect 3090 785 3120 795
rect 3180 865 3210 875
rect 3180 845 3185 865
rect 3205 845 3210 865
rect 3180 815 3210 845
rect 3180 795 3185 815
rect 3205 795 3210 815
rect 3180 785 3210 795
rect 3270 865 3300 875
rect 3270 845 3275 865
rect 3295 845 3300 865
rect 3270 815 3300 845
rect 3270 795 3275 815
rect 3295 795 3300 815
rect 3270 785 3300 795
rect 3360 865 3390 875
rect 3360 845 3365 865
rect 3385 845 3390 865
rect 3360 815 3390 845
rect 3360 795 3365 815
rect 3385 795 3390 815
rect 3360 785 3390 795
rect 3450 865 3480 875
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 815 3480 845
rect 3450 795 3455 815
rect 3475 795 3480 815
rect 3450 785 3480 795
rect 3540 865 3570 875
rect 3540 845 3545 865
rect 3565 845 3570 865
rect 3540 815 3570 845
rect 3540 795 3545 815
rect 3565 795 3570 815
rect 3540 785 3570 795
rect 3630 865 3660 875
rect 3630 845 3635 865
rect 3655 845 3660 865
rect 3630 815 3660 845
rect 3630 795 3635 815
rect 3655 795 3660 815
rect 3630 785 3660 795
rect 3720 865 3750 875
rect 3720 845 3725 865
rect 3745 845 3750 865
rect 3720 815 3750 845
rect 3720 795 3725 815
rect 3745 795 3750 815
rect 3720 785 3750 795
rect 3810 865 3840 875
rect 3810 845 3815 865
rect 3835 845 3840 865
rect 3810 815 3840 845
rect 3810 795 3815 815
rect 3835 795 3840 815
rect 3810 785 3840 795
rect 3900 865 3930 875
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 815 3930 845
rect 3900 795 3905 815
rect 3925 795 3930 815
rect 3900 785 3930 795
rect 3990 865 4020 875
rect 3990 845 3995 865
rect 4015 845 4020 865
rect 3990 815 4020 845
rect 3990 795 3995 815
rect 4015 795 4020 815
rect 3990 785 4020 795
rect 4080 865 4110 875
rect 4080 845 4085 865
rect 4105 845 4110 865
rect 4080 815 4110 845
rect 4080 795 4085 815
rect 4105 795 4110 815
rect 4080 785 4110 795
rect 4170 865 4200 875
rect 4170 845 4175 865
rect 4195 845 4200 865
rect 4170 815 4200 845
rect 4170 795 4175 815
rect 4195 795 4200 815
rect 4170 785 4200 795
rect 4260 865 4290 875
rect 4260 845 4265 865
rect 4285 845 4290 865
rect 4260 815 4290 845
rect 4260 795 4265 815
rect 4285 795 4290 815
rect 4260 785 4290 795
rect 4350 865 4380 875
rect 4350 845 4355 865
rect 4375 845 4380 865
rect 4350 815 4380 845
rect 4350 795 4355 815
rect 4375 795 4380 815
rect 4350 785 4380 795
rect 4440 865 4470 875
rect 4440 845 4445 865
rect 4465 845 4470 865
rect 4440 815 4470 845
rect 4440 795 4445 815
rect 4465 795 4470 815
rect 4440 785 4470 795
rect 4530 865 4560 875
rect 4530 845 4535 865
rect 4555 845 4560 865
rect 4530 815 4560 845
rect 4530 795 4535 815
rect 4555 795 4560 815
rect 4530 785 4560 795
rect 4620 865 4650 875
rect 4620 845 4625 865
rect 4645 845 4650 865
rect 4620 815 4650 845
rect 4620 795 4625 815
rect 4645 795 4650 815
rect 4620 785 4650 795
rect 4710 865 4740 875
rect 4710 845 4715 865
rect 4735 845 4740 865
rect 4710 815 4740 845
rect 4710 795 4715 815
rect 4735 795 4740 815
rect 4710 785 4740 795
rect 4800 865 4830 875
rect 4800 845 4805 865
rect 4825 845 4830 865
rect 4800 815 4830 845
rect 4800 795 4805 815
rect 4825 795 4830 815
rect 4800 785 4830 795
rect 4890 865 4920 875
rect 4890 845 4895 865
rect 4915 845 4920 865
rect 4890 815 4920 845
rect 4890 795 4895 815
rect 4915 795 4920 815
rect 4890 785 4920 795
rect 4980 865 5050 875
rect 4980 845 4985 865
rect 5005 845 5025 865
rect 5045 845 5050 865
rect 4980 815 5050 845
rect 16010 825 16040 855
rect 16495 820 16535 860
rect 16940 830 16970 860
rect 17160 830 17190 860
rect 17380 830 17410 860
rect 17965 830 17995 860
rect 4980 795 4985 815
rect 5005 795 5025 815
rect 5045 795 5050 815
rect 4980 785 5050 795
rect 3095 765 3115 785
rect 3275 765 3295 785
rect 3455 765 3475 785
rect 3635 765 3655 785
rect 3815 765 3835 785
rect 3995 765 4015 785
rect 4175 765 4195 785
rect 4355 765 4375 785
rect 4535 765 4555 785
rect 4715 765 4735 785
rect 4895 765 4915 785
rect 15805 770 15835 800
rect 16305 795 16345 805
rect 16305 785 16315 795
rect 16275 775 16315 785
rect 16335 775 16345 795
rect 16275 765 16345 775
rect 16375 795 16415 805
rect 16375 775 16385 795
rect 16405 775 16415 795
rect 16375 765 16415 775
rect 16445 795 16485 805
rect 16445 775 16455 795
rect 16475 775 16485 795
rect 16445 765 16485 775
rect 2525 730 2555 760
rect 3095 755 3170 765
rect 3095 745 3140 755
rect 3130 735 3140 745
rect 3160 735 3170 755
rect 3130 725 3170 735
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 755 3665 765
rect 3625 735 3635 755
rect 3655 735 3665 755
rect 3625 725 3665 735
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 755 4025 765
rect 3985 735 3995 755
rect 4015 735 4025 755
rect 3985 725 4025 735
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 755 4385 765
rect 4345 735 4355 755
rect 4375 735 4385 755
rect 4345 725 4385 735
rect 4525 755 4565 765
rect 4525 735 4535 755
rect 4555 735 4565 755
rect 4525 725 4565 735
rect 4705 755 4745 765
rect 4705 735 4715 755
rect 4735 735 4745 755
rect 4705 725 4745 735
rect 4885 755 4925 765
rect 4885 735 4895 755
rect 4915 735 4925 755
rect 16275 745 16295 765
rect 16505 745 16525 820
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 16935 765 16975 775
rect 17045 795 17085 805
rect 17045 775 17055 795
rect 17075 775 17085 795
rect 17045 765 17085 775
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17155 765 17195 775
rect 17265 795 17305 805
rect 17265 775 17275 795
rect 17295 775 17305 795
rect 17265 765 17305 775
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 17375 765 17415 775
rect 17485 795 17525 805
rect 17485 775 17495 795
rect 17515 775 17525 795
rect 17485 765 17525 775
rect 17910 770 17940 800
rect 16945 745 16965 765
rect 17055 745 17075 765
rect 17165 745 17185 765
rect 17275 745 17295 765
rect 17385 745 17405 765
rect 17495 745 17515 765
rect 26155 755 26175 900
rect 26210 1070 26240 1080
rect 26210 1050 26215 1070
rect 26235 1050 26240 1070
rect 26210 1020 26240 1050
rect 26210 1000 26215 1020
rect 26235 1000 26240 1020
rect 26210 970 26240 1000
rect 26210 950 26215 970
rect 26235 950 26240 970
rect 26210 920 26240 950
rect 26210 900 26215 920
rect 26235 900 26240 920
rect 26210 870 26240 900
rect 26210 850 26215 870
rect 26235 850 26240 870
rect 26210 840 26240 850
rect 26265 1070 26295 1080
rect 26265 1050 26270 1070
rect 26290 1050 26295 1070
rect 26265 1020 26295 1050
rect 26265 1000 26270 1020
rect 26290 1000 26295 1020
rect 26265 970 26295 1000
rect 26265 950 26270 970
rect 26290 950 26295 970
rect 26265 920 26295 950
rect 26265 900 26270 920
rect 26290 900 26295 920
rect 26265 870 26295 900
rect 26265 850 26270 870
rect 26290 850 26295 870
rect 26265 840 26295 850
rect 26320 1070 26350 1080
rect 26320 1050 26325 1070
rect 26345 1050 26350 1070
rect 26320 1020 26350 1050
rect 26320 1000 26325 1020
rect 26345 1000 26350 1020
rect 26320 970 26350 1000
rect 26320 950 26325 970
rect 26345 950 26350 970
rect 26320 920 26350 950
rect 26320 900 26325 920
rect 26345 900 26350 920
rect 26320 870 26350 900
rect 26320 850 26325 870
rect 26345 850 26350 870
rect 26320 840 26350 850
rect 26375 1070 26405 1080
rect 26375 1050 26380 1070
rect 26400 1050 26405 1070
rect 26375 1020 26405 1050
rect 26375 1000 26380 1020
rect 26400 1000 26405 1020
rect 26375 970 26405 1000
rect 26375 950 26380 970
rect 26400 950 26405 970
rect 26375 920 26405 950
rect 26375 900 26380 920
rect 26400 900 26405 920
rect 26375 870 26405 900
rect 26375 850 26380 870
rect 26400 850 26405 870
rect 26375 840 26405 850
rect 26430 1070 26460 1080
rect 26430 1050 26435 1070
rect 26455 1050 26460 1070
rect 26430 1020 26460 1050
rect 26430 1000 26435 1020
rect 26455 1000 26460 1020
rect 26430 970 26460 1000
rect 26430 950 26435 970
rect 26455 950 26460 970
rect 26430 920 26460 950
rect 26430 900 26435 920
rect 26455 900 26460 920
rect 26430 870 26460 900
rect 26430 850 26435 870
rect 26455 850 26460 870
rect 26430 840 26460 850
rect 26485 1070 26515 1080
rect 26485 1050 26490 1070
rect 26510 1050 26515 1070
rect 26485 1020 26515 1050
rect 26485 1000 26490 1020
rect 26510 1000 26515 1020
rect 26485 970 26515 1000
rect 26485 950 26490 970
rect 26510 950 26515 970
rect 26485 920 26515 950
rect 26485 900 26490 920
rect 26510 900 26515 920
rect 26485 870 26515 900
rect 26485 850 26490 870
rect 26510 850 26515 870
rect 26485 840 26515 850
rect 26540 1070 26570 1080
rect 26540 1050 26545 1070
rect 26565 1050 26570 1070
rect 26540 1020 26570 1050
rect 26540 1000 26545 1020
rect 26565 1000 26570 1020
rect 26540 970 26570 1000
rect 26540 950 26545 970
rect 26565 950 26570 970
rect 26540 920 26570 950
rect 26540 900 26545 920
rect 26565 900 26570 920
rect 26540 870 26570 900
rect 26540 850 26545 870
rect 26565 850 26570 870
rect 26540 840 26570 850
rect 26595 1070 26625 1080
rect 26595 1050 26600 1070
rect 26620 1050 26625 1070
rect 26595 1020 26625 1050
rect 26595 1000 26600 1020
rect 26620 1000 26625 1020
rect 26595 970 26625 1000
rect 26595 950 26600 970
rect 26620 950 26625 970
rect 26595 920 26625 950
rect 26595 900 26600 920
rect 26620 900 26625 920
rect 26595 870 26625 900
rect 26595 850 26600 870
rect 26620 850 26625 870
rect 26595 840 26625 850
rect 26650 1070 26680 1080
rect 26650 1050 26655 1070
rect 26675 1050 26680 1070
rect 26650 1020 26680 1050
rect 26650 1000 26655 1020
rect 26675 1000 26680 1020
rect 26650 970 26680 1000
rect 26650 950 26655 970
rect 26675 950 26680 970
rect 26650 920 26680 950
rect 26650 900 26655 920
rect 26675 900 26680 920
rect 26650 870 26680 900
rect 26650 850 26655 870
rect 26675 850 26680 870
rect 26650 840 26680 850
rect 26705 1070 26735 1080
rect 26705 1050 26710 1070
rect 26730 1050 26735 1070
rect 26705 1020 26735 1050
rect 26705 1000 26710 1020
rect 26730 1000 26735 1020
rect 26705 970 26735 1000
rect 26705 950 26710 970
rect 26730 950 26735 970
rect 26705 920 26735 950
rect 26705 900 26710 920
rect 26730 900 26735 920
rect 26705 870 26735 900
rect 26705 850 26710 870
rect 26730 850 26735 870
rect 26705 840 26735 850
rect 26760 1070 26790 1080
rect 26760 1050 26765 1070
rect 26785 1050 26790 1070
rect 26760 1020 26790 1050
rect 26760 1000 26765 1020
rect 26785 1000 26790 1020
rect 26760 970 26790 1000
rect 26760 950 26765 970
rect 26785 950 26790 970
rect 26760 920 26790 950
rect 26760 900 26765 920
rect 26785 900 26790 920
rect 26760 870 26790 900
rect 26760 850 26765 870
rect 26785 850 26790 870
rect 26760 840 26790 850
rect 26815 1070 26845 1080
rect 26815 1050 26820 1070
rect 26840 1050 26845 1070
rect 26815 1020 26845 1050
rect 26815 1000 26820 1020
rect 26840 1000 26845 1020
rect 26815 970 26845 1000
rect 26815 950 26820 970
rect 26840 950 26845 970
rect 26815 920 26845 950
rect 26815 900 26820 920
rect 26840 900 26845 920
rect 26815 870 26845 900
rect 26815 850 26820 870
rect 26840 850 26845 870
rect 26815 840 26845 850
rect 26870 1070 26900 1080
rect 26870 1050 26875 1070
rect 26895 1050 26900 1070
rect 26870 1020 26900 1050
rect 26870 1000 26875 1020
rect 26895 1000 26900 1020
rect 26870 970 26900 1000
rect 26870 950 26875 970
rect 26895 950 26900 970
rect 26870 920 26900 950
rect 26870 900 26875 920
rect 26895 900 26900 920
rect 26870 870 26900 900
rect 26870 850 26875 870
rect 26895 850 26900 870
rect 26870 840 26900 850
rect 26925 1070 26955 1080
rect 26925 1050 26930 1070
rect 26950 1050 26955 1070
rect 26925 1020 26955 1050
rect 26925 1000 26930 1020
rect 26950 1000 26955 1020
rect 26925 970 26955 1000
rect 26925 950 26930 970
rect 26950 950 26955 970
rect 26925 920 26955 950
rect 26925 900 26930 920
rect 26950 900 26955 920
rect 26925 870 26955 900
rect 26925 850 26930 870
rect 26950 850 26955 870
rect 26925 840 26955 850
rect 26980 1070 27010 1080
rect 26980 1050 26985 1070
rect 27005 1050 27010 1070
rect 26980 1020 27010 1050
rect 26980 1000 26985 1020
rect 27005 1000 27010 1020
rect 26980 970 27010 1000
rect 26980 950 26985 970
rect 27005 950 27010 970
rect 26980 920 27010 950
rect 26980 900 26985 920
rect 27005 900 27010 920
rect 26980 870 27010 900
rect 26980 850 26985 870
rect 27005 850 27010 870
rect 26980 840 27010 850
rect 27035 1070 27065 1080
rect 27035 1050 27040 1070
rect 27060 1050 27065 1070
rect 27035 1020 27065 1050
rect 27035 1000 27040 1020
rect 27060 1000 27065 1020
rect 27035 970 27065 1000
rect 27035 950 27040 970
rect 27060 950 27065 970
rect 27035 920 27065 950
rect 27035 900 27040 920
rect 27060 900 27065 920
rect 27035 870 27065 900
rect 27035 850 27040 870
rect 27060 850 27065 870
rect 27035 840 27065 850
rect 27090 1070 27120 1080
rect 27090 1050 27095 1070
rect 27115 1050 27120 1070
rect 27090 1020 27120 1050
rect 27090 1000 27095 1020
rect 27115 1000 27120 1020
rect 27090 970 27120 1000
rect 27090 950 27095 970
rect 27115 950 27120 970
rect 27090 920 27120 950
rect 27090 900 27095 920
rect 27115 900 27120 920
rect 27090 870 27120 900
rect 27090 850 27095 870
rect 27115 850 27120 870
rect 27090 840 27120 850
rect 27145 1070 27175 1080
rect 27145 1050 27150 1070
rect 27170 1050 27175 1070
rect 27145 1020 27175 1050
rect 27145 1000 27150 1020
rect 27170 1000 27175 1020
rect 27145 970 27175 1000
rect 27145 950 27150 970
rect 27170 950 27175 970
rect 27145 920 27175 950
rect 27145 900 27150 920
rect 27170 900 27175 920
rect 27145 870 27175 900
rect 27145 850 27150 870
rect 27170 850 27175 870
rect 27145 840 27175 850
rect 27200 1070 27230 1080
rect 27200 1050 27205 1070
rect 27225 1050 27230 1070
rect 27200 1020 27230 1050
rect 27200 1000 27205 1020
rect 27225 1000 27230 1020
rect 27200 970 27230 1000
rect 27200 950 27205 970
rect 27225 950 27230 970
rect 27200 920 27230 950
rect 27200 900 27205 920
rect 27225 900 27230 920
rect 27200 870 27230 900
rect 27200 850 27205 870
rect 27225 850 27230 870
rect 27200 840 27230 850
rect 27255 1070 27285 1080
rect 27255 1050 27260 1070
rect 27280 1050 27285 1070
rect 27255 1020 27285 1050
rect 27255 1000 27260 1020
rect 27280 1000 27285 1020
rect 27255 970 27285 1000
rect 27255 950 27260 970
rect 27280 950 27285 970
rect 27255 920 27285 950
rect 27255 900 27260 920
rect 27280 900 27285 920
rect 27255 870 27285 900
rect 27255 850 27260 870
rect 27280 850 27285 870
rect 27255 840 27285 850
rect 27310 1070 27340 1080
rect 27310 1050 27315 1070
rect 27335 1050 27340 1070
rect 27310 1020 27340 1050
rect 27310 1000 27315 1020
rect 27335 1000 27340 1020
rect 27310 970 27340 1000
rect 27310 950 27315 970
rect 27335 950 27340 970
rect 27310 920 27340 950
rect 27310 900 27315 920
rect 27335 900 27340 920
rect 27310 870 27340 900
rect 27310 850 27315 870
rect 27335 850 27340 870
rect 27310 840 27340 850
rect 27365 1070 27395 1080
rect 27365 1050 27370 1070
rect 27390 1050 27395 1070
rect 27365 1020 27395 1050
rect 27365 1000 27370 1020
rect 27390 1000 27395 1020
rect 27365 970 27395 1000
rect 27365 950 27370 970
rect 27390 950 27395 970
rect 27365 920 27395 950
rect 27365 900 27370 920
rect 27390 900 27395 920
rect 27365 870 27395 900
rect 27365 850 27370 870
rect 27390 850 27395 870
rect 27365 840 27395 850
rect 27420 1070 27450 1080
rect 27420 1050 27425 1070
rect 27445 1050 27450 1070
rect 27420 1020 27450 1050
rect 27420 1000 27425 1020
rect 27445 1000 27450 1020
rect 27420 970 27450 1000
rect 27420 950 27425 970
rect 27445 950 27450 970
rect 27420 920 27450 950
rect 27420 900 27425 920
rect 27445 900 27450 920
rect 27420 870 27450 900
rect 27420 850 27425 870
rect 27445 850 27450 870
rect 27420 840 27450 850
rect 27475 1070 27505 1080
rect 27475 1050 27480 1070
rect 27500 1050 27505 1070
rect 27475 1020 27505 1050
rect 27475 1000 27480 1020
rect 27500 1000 27505 1020
rect 27475 970 27505 1000
rect 27475 950 27480 970
rect 27500 950 27505 970
rect 27475 920 27505 950
rect 27475 900 27480 920
rect 27500 900 27505 920
rect 27475 870 27505 900
rect 27475 850 27480 870
rect 27500 850 27505 870
rect 27475 840 27505 850
rect 27530 1070 27560 1080
rect 27530 1050 27535 1070
rect 27555 1050 27560 1070
rect 27530 1020 27560 1050
rect 27530 1000 27535 1020
rect 27555 1000 27560 1020
rect 27530 970 27560 1000
rect 27530 950 27535 970
rect 27555 950 27560 970
rect 27530 920 27560 950
rect 27530 900 27535 920
rect 27555 900 27560 920
rect 27530 870 27560 900
rect 27530 850 27535 870
rect 27555 850 27560 870
rect 27530 840 27560 850
rect 27585 1070 27615 1080
rect 27585 1050 27590 1070
rect 27610 1050 27615 1070
rect 27585 1020 27615 1050
rect 27585 1000 27590 1020
rect 27610 1000 27615 1020
rect 27585 970 27615 1000
rect 27585 950 27590 970
rect 27610 950 27615 970
rect 27585 920 27615 950
rect 27585 900 27590 920
rect 27610 900 27615 920
rect 27585 870 27615 900
rect 27585 850 27590 870
rect 27610 850 27615 870
rect 27585 840 27615 850
rect 27655 980 27675 1175
rect 26215 820 26235 840
rect 26270 820 26290 840
rect 26380 820 26400 840
rect 26490 820 26510 840
rect 26600 820 26620 840
rect 26710 820 26730 840
rect 26820 820 26840 840
rect 26930 820 26950 840
rect 27040 820 27060 840
rect 27150 820 27170 840
rect 27260 820 27280 840
rect 27370 820 27390 840
rect 27480 820 27500 840
rect 27590 820 27610 840
rect 26195 810 26235 820
rect 26195 790 26205 810
rect 26225 790 26235 810
rect 26195 780 26235 790
rect 26260 810 26300 820
rect 26260 790 26270 810
rect 26290 790 26300 810
rect 26260 780 26300 790
rect 26370 810 26410 820
rect 26370 790 26380 810
rect 26400 790 26410 810
rect 26370 780 26410 790
rect 26480 810 26520 820
rect 26480 790 26490 810
rect 26510 790 26520 810
rect 26480 780 26520 790
rect 26590 810 26630 820
rect 26590 790 26600 810
rect 26620 790 26630 810
rect 26590 780 26630 790
rect 26700 810 26740 820
rect 26700 790 26710 810
rect 26730 790 26740 810
rect 26700 780 26740 790
rect 26810 810 26850 820
rect 26810 790 26820 810
rect 26840 790 26850 810
rect 26810 780 26850 790
rect 26920 810 26960 820
rect 26920 790 26930 810
rect 26950 790 26960 810
rect 26920 780 26960 790
rect 27030 810 27070 820
rect 27030 790 27040 810
rect 27060 790 27070 810
rect 27030 780 27070 790
rect 27140 810 27180 820
rect 27140 790 27150 810
rect 27170 790 27180 810
rect 27140 780 27180 790
rect 27250 810 27290 820
rect 27250 790 27260 810
rect 27280 790 27290 810
rect 27250 780 27290 790
rect 27360 810 27400 820
rect 27360 790 27370 810
rect 27390 790 27400 810
rect 27360 780 27400 790
rect 27470 810 27510 820
rect 27470 790 27480 810
rect 27500 790 27510 810
rect 27470 780 27510 790
rect 27585 810 27625 820
rect 27585 790 27595 810
rect 27615 790 27625 810
rect 27585 780 27625 790
rect 27655 755 27675 900
rect 28155 880 28175 1265
rect 28210 1640 28240 1650
rect 28210 1620 28215 1640
rect 28235 1620 28240 1640
rect 28210 1590 28240 1620
rect 28210 1570 28215 1590
rect 28235 1570 28240 1590
rect 28210 1540 28240 1570
rect 28210 1520 28215 1540
rect 28235 1520 28240 1540
rect 28210 1490 28240 1520
rect 28210 1470 28215 1490
rect 28235 1470 28240 1490
rect 28210 1440 28240 1470
rect 28210 1420 28215 1440
rect 28235 1420 28240 1440
rect 28210 1390 28240 1420
rect 28210 1370 28215 1390
rect 28235 1370 28240 1390
rect 28210 1340 28240 1370
rect 28210 1320 28215 1340
rect 28235 1320 28240 1340
rect 28210 1290 28240 1320
rect 28210 1270 28215 1290
rect 28235 1270 28240 1290
rect 28210 1240 28240 1270
rect 28210 1220 28215 1240
rect 28235 1220 28240 1240
rect 28210 1190 28240 1220
rect 28210 1170 28215 1190
rect 28235 1170 28240 1190
rect 28210 1140 28240 1170
rect 28210 1120 28215 1140
rect 28235 1120 28240 1140
rect 28210 1090 28240 1120
rect 28210 1070 28215 1090
rect 28235 1070 28240 1090
rect 28210 1040 28240 1070
rect 28210 1020 28215 1040
rect 28235 1020 28240 1040
rect 28210 990 28240 1020
rect 28210 970 28215 990
rect 28235 970 28240 990
rect 28210 960 28240 970
rect 28310 1640 28340 1650
rect 28310 1620 28315 1640
rect 28335 1620 28340 1640
rect 28310 1590 28340 1620
rect 28310 1570 28315 1590
rect 28335 1570 28340 1590
rect 28310 1540 28340 1570
rect 28310 1520 28315 1540
rect 28335 1520 28340 1540
rect 28310 1490 28340 1520
rect 28310 1470 28315 1490
rect 28335 1470 28340 1490
rect 28310 1440 28340 1470
rect 28310 1420 28315 1440
rect 28335 1420 28340 1440
rect 28310 1390 28340 1420
rect 28310 1370 28315 1390
rect 28335 1370 28340 1390
rect 28310 1340 28340 1370
rect 28310 1320 28315 1340
rect 28335 1320 28340 1340
rect 28310 1290 28340 1320
rect 28310 1270 28315 1290
rect 28335 1270 28340 1290
rect 28310 1240 28340 1270
rect 28310 1220 28315 1240
rect 28335 1220 28340 1240
rect 28310 1190 28340 1220
rect 28310 1170 28315 1190
rect 28335 1170 28340 1190
rect 28310 1140 28340 1170
rect 28310 1120 28315 1140
rect 28335 1120 28340 1140
rect 28310 1090 28340 1120
rect 28310 1070 28315 1090
rect 28335 1070 28340 1090
rect 28310 1040 28340 1070
rect 28310 1020 28315 1040
rect 28335 1020 28340 1040
rect 28310 990 28340 1020
rect 28310 970 28315 990
rect 28335 970 28340 990
rect 28310 960 28340 970
rect 28410 1640 28440 1650
rect 28410 1620 28415 1640
rect 28435 1620 28440 1640
rect 28410 1590 28440 1620
rect 28410 1570 28415 1590
rect 28435 1570 28440 1590
rect 28410 1540 28440 1570
rect 28410 1520 28415 1540
rect 28435 1520 28440 1540
rect 28410 1490 28440 1520
rect 28410 1470 28415 1490
rect 28435 1470 28440 1490
rect 28410 1440 28440 1470
rect 28410 1420 28415 1440
rect 28435 1420 28440 1440
rect 28410 1390 28440 1420
rect 28410 1370 28415 1390
rect 28435 1370 28440 1390
rect 28410 1340 28440 1370
rect 28410 1320 28415 1340
rect 28435 1320 28440 1340
rect 28410 1290 28440 1320
rect 28410 1270 28415 1290
rect 28435 1270 28440 1290
rect 28410 1240 28440 1270
rect 28410 1220 28415 1240
rect 28435 1220 28440 1240
rect 28410 1190 28440 1220
rect 28410 1170 28415 1190
rect 28435 1170 28440 1190
rect 28410 1140 28440 1170
rect 28410 1120 28415 1140
rect 28435 1120 28440 1140
rect 28410 1090 28440 1120
rect 28410 1070 28415 1090
rect 28435 1070 28440 1090
rect 28410 1040 28440 1070
rect 28410 1020 28415 1040
rect 28435 1020 28440 1040
rect 28410 990 28440 1020
rect 28410 970 28415 990
rect 28435 970 28440 990
rect 28410 960 28440 970
rect 28510 1640 28540 1650
rect 28510 1620 28515 1640
rect 28535 1620 28540 1640
rect 28510 1590 28540 1620
rect 28510 1570 28515 1590
rect 28535 1570 28540 1590
rect 28510 1540 28540 1570
rect 28510 1520 28515 1540
rect 28535 1520 28540 1540
rect 28510 1490 28540 1520
rect 28510 1470 28515 1490
rect 28535 1470 28540 1490
rect 28510 1440 28540 1470
rect 28510 1420 28515 1440
rect 28535 1420 28540 1440
rect 28510 1390 28540 1420
rect 28510 1370 28515 1390
rect 28535 1370 28540 1390
rect 28510 1340 28540 1370
rect 28510 1320 28515 1340
rect 28535 1320 28540 1340
rect 28510 1290 28540 1320
rect 28510 1270 28515 1290
rect 28535 1270 28540 1290
rect 28510 1240 28540 1270
rect 28510 1220 28515 1240
rect 28535 1220 28540 1240
rect 28510 1190 28540 1220
rect 28510 1170 28515 1190
rect 28535 1170 28540 1190
rect 28510 1140 28540 1170
rect 28510 1120 28515 1140
rect 28535 1120 28540 1140
rect 28510 1090 28540 1120
rect 28510 1070 28515 1090
rect 28535 1070 28540 1090
rect 28510 1040 28540 1070
rect 28510 1020 28515 1040
rect 28535 1020 28540 1040
rect 28510 990 28540 1020
rect 28510 970 28515 990
rect 28535 970 28540 990
rect 28510 960 28540 970
rect 28610 1640 28640 1650
rect 28610 1620 28615 1640
rect 28635 1620 28640 1640
rect 28610 1590 28640 1620
rect 28610 1570 28615 1590
rect 28635 1570 28640 1590
rect 28610 1540 28640 1570
rect 28610 1520 28615 1540
rect 28635 1520 28640 1540
rect 28610 1490 28640 1520
rect 28610 1470 28615 1490
rect 28635 1470 28640 1490
rect 28610 1440 28640 1470
rect 28610 1420 28615 1440
rect 28635 1420 28640 1440
rect 28610 1390 28640 1420
rect 28610 1370 28615 1390
rect 28635 1370 28640 1390
rect 28610 1340 28640 1370
rect 28610 1320 28615 1340
rect 28635 1320 28640 1340
rect 28610 1290 28640 1320
rect 28610 1270 28615 1290
rect 28635 1270 28640 1290
rect 28610 1240 28640 1270
rect 28610 1220 28615 1240
rect 28635 1220 28640 1240
rect 28610 1190 28640 1220
rect 28610 1170 28615 1190
rect 28635 1170 28640 1190
rect 28610 1140 28640 1170
rect 28610 1120 28615 1140
rect 28635 1120 28640 1140
rect 28610 1090 28640 1120
rect 28610 1070 28615 1090
rect 28635 1070 28640 1090
rect 28610 1040 28640 1070
rect 28610 1020 28615 1040
rect 28635 1020 28640 1040
rect 28610 990 28640 1020
rect 28610 970 28615 990
rect 28635 970 28640 990
rect 28610 960 28640 970
rect 28710 1640 28740 1650
rect 28710 1620 28715 1640
rect 28735 1620 28740 1640
rect 28710 1590 28740 1620
rect 28710 1570 28715 1590
rect 28735 1570 28740 1590
rect 28710 1540 28740 1570
rect 28710 1520 28715 1540
rect 28735 1520 28740 1540
rect 28710 1490 28740 1520
rect 28710 1470 28715 1490
rect 28735 1470 28740 1490
rect 28710 1440 28740 1470
rect 28710 1420 28715 1440
rect 28735 1420 28740 1440
rect 28710 1390 28740 1420
rect 28710 1370 28715 1390
rect 28735 1370 28740 1390
rect 28710 1340 28740 1370
rect 28710 1320 28715 1340
rect 28735 1320 28740 1340
rect 28710 1290 28740 1320
rect 28710 1270 28715 1290
rect 28735 1270 28740 1290
rect 28710 1240 28740 1270
rect 28710 1220 28715 1240
rect 28735 1220 28740 1240
rect 28710 1190 28740 1220
rect 28710 1170 28715 1190
rect 28735 1170 28740 1190
rect 28710 1140 28740 1170
rect 28710 1120 28715 1140
rect 28735 1120 28740 1140
rect 28710 1090 28740 1120
rect 28710 1070 28715 1090
rect 28735 1070 28740 1090
rect 28710 1040 28740 1070
rect 28710 1020 28715 1040
rect 28735 1020 28740 1040
rect 28710 990 28740 1020
rect 28710 970 28715 990
rect 28735 970 28740 990
rect 28710 960 28740 970
rect 28810 1640 28840 1650
rect 28810 1620 28815 1640
rect 28835 1620 28840 1640
rect 28810 1590 28840 1620
rect 28810 1570 28815 1590
rect 28835 1570 28840 1590
rect 28810 1540 28840 1570
rect 28810 1520 28815 1540
rect 28835 1520 28840 1540
rect 28810 1490 28840 1520
rect 28810 1470 28815 1490
rect 28835 1470 28840 1490
rect 28810 1440 28840 1470
rect 28810 1420 28815 1440
rect 28835 1420 28840 1440
rect 28810 1390 28840 1420
rect 28810 1370 28815 1390
rect 28835 1370 28840 1390
rect 28810 1340 28840 1370
rect 28810 1320 28815 1340
rect 28835 1320 28840 1340
rect 28810 1290 28840 1320
rect 28810 1270 28815 1290
rect 28835 1270 28840 1290
rect 28810 1240 28840 1270
rect 28810 1220 28815 1240
rect 28835 1220 28840 1240
rect 28810 1190 28840 1220
rect 28810 1170 28815 1190
rect 28835 1170 28840 1190
rect 28810 1140 28840 1170
rect 28810 1120 28815 1140
rect 28835 1120 28840 1140
rect 28810 1090 28840 1120
rect 28810 1070 28815 1090
rect 28835 1070 28840 1090
rect 28810 1040 28840 1070
rect 28810 1020 28815 1040
rect 28835 1020 28840 1040
rect 28810 990 28840 1020
rect 28810 970 28815 990
rect 28835 970 28840 990
rect 28810 960 28840 970
rect 28875 1345 28895 1730
rect 28415 940 28435 960
rect 28615 940 28635 960
rect 28405 930 28445 940
rect 28405 910 28415 930
rect 28435 910 28445 930
rect 28405 900 28445 910
rect 28605 930 28645 940
rect 28605 910 28615 930
rect 28635 910 28645 930
rect 28605 900 28645 910
rect 28875 880 28895 1265
rect 28155 860 28485 880
rect 28565 860 28895 880
rect 28985 1675 29065 1695
rect 29145 1675 29220 1695
rect 28985 1300 29005 1675
rect 29055 1640 29090 1650
rect 29055 1615 29060 1640
rect 29085 1615 29090 1640
rect 29055 1605 29090 1615
rect 29115 1640 29150 1650
rect 29115 1615 29120 1640
rect 29145 1615 29150 1640
rect 29115 1605 29150 1615
rect 28985 860 29005 1220
rect 29200 1300 29220 1675
rect 29090 910 29115 960
rect 29200 860 29220 1220
rect 28985 840 29065 860
rect 29145 840 29220 860
rect 4885 725 4925 735
rect 16265 735 16295 745
rect 16265 715 16270 735
rect 16290 715 16295 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 16265 685 16295 715
rect 16265 665 16270 685
rect 16290 665 16295 685
rect 16265 655 16295 665
rect 16495 735 16525 745
rect 16495 715 16500 735
rect 16520 715 16525 735
rect 16495 685 16525 715
rect 16845 735 16915 745
rect 16845 715 16850 735
rect 16870 715 16890 735
rect 16910 715 16915 735
rect 16845 705 16915 715
rect 16940 735 16970 745
rect 16940 715 16945 735
rect 16965 715 16970 735
rect 16940 705 16970 715
rect 16995 735 17025 745
rect 16995 715 17000 735
rect 17020 715 17025 735
rect 16995 705 17025 715
rect 17050 735 17080 745
rect 17050 715 17055 735
rect 17075 715 17080 735
rect 17050 705 17080 715
rect 17105 735 17135 745
rect 17105 715 17110 735
rect 17130 715 17135 735
rect 17105 705 17135 715
rect 17160 735 17190 745
rect 17160 715 17165 735
rect 17185 715 17190 735
rect 17160 705 17190 715
rect 17215 735 17245 745
rect 17215 715 17220 735
rect 17240 715 17245 735
rect 17215 705 17245 715
rect 17270 735 17300 745
rect 17270 715 17275 735
rect 17295 715 17300 735
rect 17270 705 17300 715
rect 17325 735 17355 745
rect 17325 715 17330 735
rect 17350 715 17355 735
rect 17325 705 17355 715
rect 17380 735 17410 745
rect 17380 715 17385 735
rect 17405 715 17410 735
rect 17380 705 17410 715
rect 17435 735 17465 745
rect 17435 715 17440 735
rect 17460 715 17465 735
rect 17435 705 17465 715
rect 17490 735 17520 745
rect 17490 715 17495 735
rect 17515 715 17520 735
rect 17490 705 17520 715
rect 17545 735 17615 745
rect 26155 735 26845 755
rect 26925 735 27675 755
rect 17545 715 17550 735
rect 17570 715 17590 735
rect 17610 715 17615 735
rect 17545 705 17615 715
rect 16850 685 16870 705
rect 17000 685 17020 705
rect 17110 685 17130 705
rect 17220 685 17240 705
rect 17330 685 17350 705
rect 17440 685 17460 705
rect 17590 685 17610 705
rect 16495 665 16500 685
rect 16520 665 16525 685
rect 16495 655 16525 665
rect 16840 675 16880 685
rect 16840 655 16850 675
rect 16870 655 16880 675
rect 16840 645 16880 655
rect 16990 675 17030 685
rect 16990 655 17000 675
rect 17020 655 17030 675
rect 16990 645 17030 655
rect 17100 675 17140 685
rect 17100 655 17110 675
rect 17130 655 17140 675
rect 17100 645 17140 655
rect 17210 675 17250 685
rect 17210 655 17220 675
rect 17240 655 17250 675
rect 17210 645 17250 655
rect 17320 675 17360 685
rect 17320 655 17330 675
rect 17350 655 17360 675
rect 17320 645 17360 655
rect 17430 675 17470 685
rect 17430 655 17440 675
rect 17460 655 17470 675
rect 17430 645 17470 655
rect 17580 675 17620 685
rect 17580 655 17590 675
rect 17610 655 17620 675
rect 17580 645 17620 655
rect 26010 625 26040 655
rect 26510 645 26540 655
rect 26940 645 26970 660
rect 27160 645 27190 660
rect 27380 645 27410 660
rect 26210 625 26355 645
rect 26435 625 26585 645
rect 25805 570 25835 600
rect 26210 555 26230 625
rect 26305 595 26345 605
rect 26305 585 26315 595
rect 26275 575 26315 585
rect 26335 575 26345 595
rect 26275 565 26345 575
rect 26375 595 26415 605
rect 26375 575 26385 595
rect 26405 575 26415 595
rect 26375 565 26415 575
rect 26445 595 26485 605
rect 26445 575 26455 595
rect 26475 575 26485 595
rect 26445 565 26485 575
rect 26505 595 26545 605
rect 26505 575 26515 595
rect 26535 575 26545 595
rect 26505 565 26545 575
rect 26275 545 26295 565
rect 26505 545 26525 565
rect 26210 415 26230 475
rect 26265 535 26295 545
rect 26265 515 26270 535
rect 26290 515 26295 535
rect 26265 485 26295 515
rect 26265 465 26270 485
rect 26290 465 26295 485
rect 26265 455 26295 465
rect 26495 535 26525 545
rect 26495 515 26500 535
rect 26520 515 26525 535
rect 26495 485 26525 515
rect 26495 465 26500 485
rect 26520 465 26525 485
rect 26495 455 26525 465
rect 26565 555 26585 625
rect 26565 415 26585 475
rect 26210 395 26355 415
rect 26435 395 26585 415
rect 26830 625 27190 645
rect 27270 625 27630 645
rect 27975 630 28005 660
rect 26830 555 26850 625
rect 26935 595 26975 605
rect 26935 575 26945 595
rect 26965 575 26975 595
rect 26935 565 26975 575
rect 27045 595 27085 605
rect 27045 575 27055 595
rect 27075 575 27085 595
rect 27045 565 27085 575
rect 27155 595 27195 605
rect 27155 575 27165 595
rect 27185 575 27195 595
rect 27155 565 27195 575
rect 27265 595 27305 605
rect 27265 575 27275 595
rect 27295 575 27305 595
rect 27265 565 27305 575
rect 27375 595 27415 605
rect 27375 575 27385 595
rect 27405 575 27415 595
rect 27375 565 27415 575
rect 27485 595 27525 605
rect 27485 575 27495 595
rect 27515 575 27525 595
rect 27485 565 27525 575
rect 26945 545 26965 565
rect 27055 545 27075 565
rect 27165 545 27185 565
rect 27275 545 27295 565
rect 27385 545 27405 565
rect 27495 545 27515 565
rect 27610 555 27630 625
rect 27920 570 27950 600
rect 26885 535 26915 545
rect 26885 515 26890 535
rect 26910 515 26915 535
rect 26885 505 26915 515
rect 26940 535 26970 545
rect 26940 515 26945 535
rect 26965 515 26970 535
rect 26940 505 26970 515
rect 26995 535 27025 545
rect 26995 515 27000 535
rect 27020 515 27025 535
rect 26995 505 27025 515
rect 27050 535 27080 545
rect 27050 515 27055 535
rect 27075 515 27080 535
rect 27050 505 27080 515
rect 27105 535 27135 545
rect 27105 515 27110 535
rect 27130 515 27135 535
rect 27105 505 27135 515
rect 27160 535 27190 545
rect 27160 515 27165 535
rect 27185 515 27190 535
rect 27160 505 27190 515
rect 27215 535 27245 545
rect 27215 515 27220 535
rect 27240 515 27245 535
rect 27215 505 27245 515
rect 27270 535 27300 545
rect 27270 515 27275 535
rect 27295 515 27300 535
rect 27270 505 27300 515
rect 27325 535 27355 545
rect 27325 515 27330 535
rect 27350 515 27355 535
rect 27325 505 27355 515
rect 27380 535 27410 545
rect 27380 515 27385 535
rect 27405 515 27410 535
rect 27380 505 27410 515
rect 27435 535 27465 545
rect 27435 515 27440 535
rect 27460 515 27465 535
rect 27435 505 27465 515
rect 27490 535 27520 545
rect 27490 515 27495 535
rect 27515 515 27520 535
rect 27490 505 27520 515
rect 27545 535 27580 545
rect 27545 515 27550 535
rect 27570 515 27580 535
rect 27545 505 27580 515
rect 27000 485 27020 505
rect 27110 485 27130 505
rect 27220 485 27240 505
rect 27330 485 27350 505
rect 27440 485 27460 505
rect 26830 425 26850 475
rect 26990 475 27030 485
rect 26990 455 27000 475
rect 27020 455 27030 475
rect 26990 445 27030 455
rect 27100 475 27140 485
rect 27100 455 27110 475
rect 27130 455 27140 475
rect 27100 445 27140 455
rect 27210 475 27250 485
rect 27210 455 27220 475
rect 27240 455 27250 475
rect 27210 445 27250 455
rect 27320 475 27360 485
rect 27320 455 27330 475
rect 27350 455 27360 475
rect 27320 445 27360 455
rect 27430 475 27470 485
rect 27430 455 27440 475
rect 27460 455 27470 475
rect 27430 445 27470 455
rect 27610 425 27630 475
rect 26830 405 27190 425
rect 27270 405 27630 425
<< viali >>
rect 26515 4900 26535 4920
rect 26575 4900 26595 4920
rect 26635 4900 26655 4920
rect 26695 4900 26715 4920
rect 26755 4900 26775 4920
rect 26815 4900 26835 4920
rect 26875 4900 26895 4920
rect 26355 4750 26375 4770
rect 26695 4745 26715 4765
rect 27245 4875 27265 4895
rect 27365 4875 27385 4895
rect 27485 4875 27505 4895
rect 27605 4875 27625 4895
rect 27725 4875 27745 4895
rect 27305 4745 27325 4765
rect 27366 4745 27384 4765
rect 27425 4745 27445 4765
rect 27545 4745 27565 4765
rect 27665 4745 27685 4765
rect 16605 4440 16625 4460
rect 16725 4440 16745 4460
rect 16845 4440 16865 4460
rect 26370 4455 26390 4475
rect 26480 4455 26500 4475
rect 26590 4455 26610 4475
rect 26700 4455 26720 4475
rect 26810 4455 26830 4475
rect 26920 4455 26940 4475
rect 27030 4455 27050 4475
rect 27140 4455 27160 4475
rect 27250 4455 27270 4475
rect 27360 4455 27380 4475
rect 16175 4380 16195 4400
rect 16435 4380 16455 4400
rect 16545 4395 16565 4415
rect 16665 4395 16685 4415
rect 16785 4395 16805 4415
rect 16905 4395 16925 4415
rect 17195 4370 17215 4390
rect 17315 4370 17335 4390
rect 17435 4370 17455 4390
rect 17555 4370 17575 4390
rect 17675 4370 17695 4390
rect 26315 4335 26335 4355
rect 26370 4335 26390 4355
rect 26425 4335 26445 4355
rect 26535 4335 26555 4355
rect 26645 4335 26665 4355
rect 26755 4335 26775 4355
rect 26865 4335 26885 4355
rect 26975 4335 26995 4355
rect 27085 4335 27105 4355
rect 27195 4335 27215 4355
rect 27305 4335 27325 4355
rect 27415 4335 27435 4355
rect 16305 4245 16325 4265
rect 16725 4240 16745 4260
rect 17255 4240 17275 4260
rect 17316 4240 17334 4260
rect 17375 4240 17395 4260
rect 17495 4240 17515 4260
rect 17615 4240 17635 4260
rect 16370 4130 16390 4150
rect 16480 4130 16500 4150
rect 16590 4130 16610 4150
rect 16700 4130 16720 4150
rect 16810 4130 16830 4150
rect 16920 4130 16940 4150
rect 17030 4130 17050 4150
rect 17140 4130 17160 4150
rect 17250 4130 17270 4150
rect 17360 4130 17380 4150
rect 16315 4010 16335 4030
rect 16370 4010 16390 4030
rect 16425 4010 16445 4030
rect 16535 4010 16555 4030
rect 16645 4010 16665 4030
rect 16755 4010 16775 4030
rect 16865 4010 16885 4030
rect 16975 4010 16995 4030
rect 17085 4010 17105 4030
rect 17195 4010 17215 4030
rect 17305 4010 17325 4030
rect 17415 4010 17435 4030
rect 26285 4045 26305 4065
rect 26330 4045 26350 4065
rect 26375 4045 26395 4065
rect 26430 4045 26450 4065
rect 26485 4045 26505 4065
rect 26540 4045 26560 4065
rect 26650 4045 26670 4065
rect 26760 4045 26780 4065
rect 27013 4045 27033 4065
rect 27060 4045 27080 4065
rect 27160 4045 27180 4065
rect 27215 4045 27235 4065
rect 27270 4045 27290 4065
rect 27380 4045 27400 4065
rect 27435 4045 27455 4065
rect 27490 4045 27510 4065
rect 16320 3885 16340 3905
rect 16425 3885 16445 3905
rect 16535 3885 16555 3905
rect 16645 3885 16665 3905
rect 16755 3885 16775 3905
rect 17060 3885 17080 3905
rect 17165 3885 17185 3905
rect 17275 3885 17295 3905
rect 17385 3885 17405 3905
rect 17495 3885 17515 3905
rect 26265 3925 26285 3945
rect 26360 3925 26380 3945
rect 26413 3925 26430 3945
rect 26485 3925 26505 3945
rect 26580 3925 26600 3945
rect 26633 3925 26650 3945
rect 26705 3925 26725 3945
rect 26780 3925 26797 3945
rect 26830 3925 26850 3945
rect 26995 3925 27015 3945
rect 27090 3925 27110 3945
rect 27143 3925 27160 3945
rect 27215 3925 27235 3945
rect 27310 3925 27330 3945
rect 27363 3925 27380 3945
rect 27435 3925 27455 3945
rect 27510 3925 27527 3945
rect 27560 3925 27580 3945
rect 16277 3825 16294 3845
rect 16370 3825 16390 3845
rect 16480 3825 16500 3845
rect 16700 3825 16720 3845
rect 16810 3825 16830 3845
rect 17017 3825 17034 3845
rect 17220 3825 17240 3845
rect 17440 3825 17460 3845
rect 16408 3705 16425 3725
rect 16628 3705 16645 3725
rect 16775 3705 16792 3725
rect 16260 3645 16280 3665
rect 15070 3610 15090 3630
rect 15180 3610 15200 3630
rect 15290 3610 15310 3630
rect 15400 3610 15420 3630
rect 15510 3610 15530 3630
rect 16365 3645 16385 3665
rect 16480 3645 16500 3665
rect 16585 3645 16605 3665
rect 16700 3645 16720 3665
rect 16815 3645 16835 3665
rect 17000 3655 17020 3675
rect 17148 3705 17165 3725
rect 17220 3655 17240 3675
rect 17368 3705 17385 3725
rect 17515 3705 17532 3725
rect 17440 3655 17460 3675
rect 15620 3610 15640 3630
rect 18210 3610 18230 3630
rect 18320 3610 18340 3630
rect 18430 3610 18450 3630
rect 18540 3610 18560 3630
rect 18650 3610 18670 3630
rect 18760 3610 18780 3630
rect 25070 3610 25090 3630
rect 25180 3610 25200 3630
rect 25290 3610 25310 3630
rect 25400 3610 25420 3630
rect 25510 3610 25530 3630
rect 25620 3610 25640 3630
rect 56 3175 81 3200
rect 1271 3170 1296 3195
rect 56 3115 81 3140
rect 1271 3110 1296 3135
rect 56 3035 81 3060
rect 56 2975 81 3000
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 2340 2930 2365 2955
rect 3090 2955 3110 2975
rect 3145 2955 3165 2975
rect 3275 2955 3295 2975
rect 3455 2955 3475 2975
rect 3635 2955 3655 2975
rect 3815 2955 3835 2975
rect 3995 2955 4015 2975
rect 4175 2955 4195 2975
rect 4355 2955 4375 2975
rect 4535 2955 4555 2975
rect 4715 2955 4735 2975
rect 4845 2955 4865 2975
rect 4895 2955 4915 2975
rect 16350 3550 16370 3570
rect 16470 3550 16490 3570
rect 16590 3550 16610 3570
rect 16710 3550 16730 3570
rect 16830 3550 16850 3570
rect 16950 3550 16970 3570
rect 17070 3550 17090 3570
rect 17190 3550 17210 3570
rect 17310 3550 17330 3570
rect 17430 3550 17450 3570
rect 16290 3080 16310 3100
rect 16410 3080 16430 3100
rect 16530 3080 16550 3100
rect 16650 3080 16670 3100
rect 16770 3080 16790 3100
rect 16831 3080 16849 3100
rect 16890 3080 16910 3100
rect 17010 3080 17030 3100
rect 17130 3080 17150 3100
rect 17250 3080 17270 3100
rect 17370 3080 17390 3100
rect 17490 3080 17510 3100
rect 2340 2870 2365 2895
rect 61 2825 86 2850
rect 734 2825 759 2850
rect 1271 2810 1296 2835
rect 1970 2810 1995 2835
rect 15125 2940 15145 2960
rect 15235 2940 15255 2960
rect 15345 2940 15365 2960
rect 15455 2940 15475 2960
rect 15511 2940 15529 2960
rect 15565 2940 15585 2960
rect 18265 2940 18285 2960
rect 18321 2940 18339 2960
rect 18375 2940 18395 2960
rect 18485 2940 18505 2960
rect 18595 2940 18615 2960
rect 18705 2940 18725 2960
rect 26350 3630 26370 3650
rect 26470 3630 26490 3650
rect 26590 3630 26610 3650
rect 26710 3630 26730 3650
rect 26830 3630 26850 3650
rect 26950 3630 26970 3650
rect 27070 3630 27090 3650
rect 27190 3630 27210 3650
rect 27310 3630 27330 3650
rect 27430 3630 27450 3650
rect 26290 3160 26310 3180
rect 26410 3160 26430 3180
rect 26530 3160 26550 3180
rect 26650 3160 26670 3180
rect 26770 3160 26790 3180
rect 26831 3160 26849 3180
rect 26890 3160 26910 3180
rect 27010 3160 27030 3180
rect 27130 3160 27150 3180
rect 27250 3160 27270 3180
rect 27370 3160 27390 3180
rect 27490 3160 27510 3180
rect 28210 3690 28230 3710
rect 28320 3690 28340 3710
rect 28430 3690 28450 3710
rect 28540 3690 28560 3710
rect 28650 3690 28670 3710
rect 28760 3690 28780 3710
rect 28265 3020 28285 3040
rect 28321 3020 28339 3040
rect 28375 3020 28395 3040
rect 28485 3020 28505 3040
rect 28595 3020 28615 3040
rect 28705 3020 28725 3040
rect 25125 2940 25145 2960
rect 25235 2940 25255 2960
rect 25345 2940 25365 2960
rect 25455 2940 25475 2960
rect 25511 2940 25529 2960
rect 25565 2940 25585 2960
rect 16145 2870 16165 2890
rect 16265 2870 16285 2890
rect 16385 2870 16405 2890
rect 16505 2870 16525 2890
rect 16625 2870 16645 2890
rect 17155 2870 17175 2890
rect 17275 2870 17295 2890
rect 17395 2870 17415 2890
rect 17515 2870 17535 2890
rect 17635 2870 17655 2890
rect 26145 2870 26165 2890
rect 26265 2870 26285 2890
rect 26385 2870 26405 2890
rect 26505 2870 26525 2890
rect 26625 2870 26645 2890
rect 61 2765 86 2790
rect 734 2765 759 2790
rect 3005 2785 3025 2805
rect 3185 2785 3205 2805
rect 3365 2785 3385 2805
rect 3545 2785 3565 2805
rect 3725 2785 3745 2805
rect 3905 2785 3925 2805
rect 4085 2785 4105 2805
rect 4265 2785 4285 2805
rect 4445 2785 4465 2805
rect 4625 2785 4645 2805
rect 4805 2785 4825 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 3365 2725 3385 2745
rect 3545 2725 3565 2745
rect 3725 2725 3745 2745
rect 3905 2725 3925 2745
rect 4085 2725 4105 2745
rect 4265 2725 4285 2745
rect 4445 2725 4465 2745
rect 4625 2725 4645 2745
rect 4805 2725 4825 2745
rect 15070 2680 15090 2700
rect 15180 2680 15200 2700
rect 15290 2680 15310 2700
rect 15400 2680 15420 2700
rect 15510 2680 15530 2700
rect 15620 2680 15640 2700
rect 18210 2680 18230 2700
rect 18320 2680 18340 2700
rect 18430 2680 18450 2700
rect 18540 2680 18560 2700
rect 18650 2680 18670 2700
rect 18760 2680 18780 2700
rect 25070 2680 25090 2700
rect 25180 2680 25200 2700
rect 25290 2680 25310 2700
rect 25400 2680 25420 2700
rect 25510 2680 25530 2700
rect 25620 2680 25640 2700
rect 16085 2450 16105 2470
rect 16205 2450 16225 2470
rect 16325 2450 16345 2470
rect 16386 2450 16404 2470
rect 16445 2450 16465 2470
rect 16565 2450 16585 2470
rect 16685 2450 16705 2470
rect 17095 2450 17115 2470
rect 17215 2450 17235 2470
rect 17335 2450 17355 2470
rect 17396 2450 17414 2470
rect 17455 2450 17475 2470
rect 17575 2450 17595 2470
rect 17695 2450 17715 2470
rect 3275 2355 3295 2375
rect 3365 2350 3385 2370
rect 3455 2355 3475 2375
rect 3815 2355 3835 2375
rect 3895 2355 3915 2375
rect 3995 2355 4015 2375
rect 4175 2355 4195 2375
rect 15125 2410 15145 2430
rect 15235 2410 15255 2430
rect 15345 2410 15365 2430
rect 15455 2410 15475 2430
rect 15565 2410 15585 2430
rect 18265 2410 18285 2430
rect 18375 2410 18395 2430
rect 18485 2410 18505 2430
rect 18595 2410 18615 2430
rect 18705 2410 18725 2430
rect 27165 2870 27185 2890
rect 27285 2870 27305 2890
rect 27405 2870 27425 2890
rect 27525 2870 27545 2890
rect 27645 2870 27665 2890
rect 26085 2450 26105 2470
rect 26205 2450 26225 2470
rect 26325 2450 26345 2470
rect 26386 2450 26404 2470
rect 26445 2450 26465 2470
rect 26565 2450 26585 2470
rect 26685 2450 26705 2470
rect 25125 2410 25145 2430
rect 25235 2410 25255 2430
rect 25345 2410 25365 2430
rect 25455 2410 25475 2430
rect 25565 2410 25585 2430
rect 27105 2450 27125 2470
rect 27225 2450 27245 2470
rect 27345 2450 27365 2470
rect 27406 2450 27424 2470
rect 27465 2450 27485 2470
rect 27585 2450 27605 2470
rect 27705 2450 27725 2470
rect 28210 2730 28230 2750
rect 28320 2730 28340 2750
rect 28430 2730 28450 2750
rect 28540 2730 28560 2750
rect 28650 2730 28670 2750
rect 28760 2730 28780 2750
rect 28265 2460 28285 2480
rect 28321 2460 28339 2480
rect 28375 2460 28395 2480
rect 28485 2460 28505 2480
rect 28595 2460 28615 2480
rect 28705 2460 28725 2480
rect 4535 2355 4555 2375
rect 4715 2355 4735 2375
rect 15595 2350 15615 2370
rect 18235 2350 18255 2370
rect 25595 2350 25615 2370
rect 3635 2310 3655 2330
rect 4355 2310 4375 2330
rect 3455 2265 3475 2285
rect 4535 2265 4555 2285
rect 15125 2290 15145 2310
rect 15235 2290 15255 2310
rect 15345 2290 15365 2310
rect 15455 2290 15475 2310
rect 15565 2290 15585 2310
rect 18265 2290 18285 2310
rect 18375 2290 18395 2310
rect 18485 2290 18505 2310
rect 18595 2290 18615 2310
rect 18705 2290 18725 2310
rect 25125 2290 25145 2310
rect 25235 2290 25255 2310
rect 25345 2290 25365 2310
rect 25455 2290 25475 2310
rect 25565 2290 25585 2310
rect 2755 2070 2775 2090
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 3995 2070 4015 2090
rect 4155 2070 4175 2090
rect 4275 2070 4295 2090
rect 4395 2070 4415 2090
rect 4515 2070 4535 2090
rect 4635 2070 4655 2090
rect 4755 2070 4775 2090
rect 4875 2070 4895 2090
rect 4995 2070 5015 2090
rect 5115 2070 5135 2090
rect 5235 2070 5255 2090
rect 2630 2025 2650 2045
rect -35 1695 -15 1715
rect 2815 2025 2835 2045
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4095 2025 4115 2045
rect 4455 2025 4475 2045
rect 4815 2025 4835 2045
rect 5175 2025 5195 2045
rect 14645 1975 14670 2000
rect 14705 1975 14730 2000
rect 14765 1975 14790 2000
rect 14825 1975 14850 2000
rect 16340 2155 16360 2175
rect 16450 2155 16470 2175
rect 16560 2155 16580 2175
rect 16670 2155 16690 2175
rect 16780 2155 16800 2175
rect 16836 2155 16854 2175
rect 16890 2155 16910 2175
rect 17000 2155 17020 2175
rect 17110 2155 17130 2175
rect 17220 2155 17240 2175
rect 17330 2155 17350 2175
rect 17440 2155 17460 2175
rect 19000 1975 19025 2000
rect 15070 1920 15088 1940
rect 15180 1920 15198 1940
rect 15290 1920 15308 1940
rect 15400 1920 15418 1940
rect 15510 1920 15528 1940
rect 15620 1920 15638 1940
rect 16395 1935 16415 1955
rect 16505 1935 16525 1955
rect 16615 1935 16635 1955
rect 16725 1935 16745 1955
rect 16835 1935 16855 1955
rect 16945 1935 16965 1955
rect 17055 1935 17075 1955
rect 17165 1935 17185 1955
rect 17275 1935 17295 1955
rect 17385 1935 17405 1955
rect 19060 1975 19085 2000
rect 19120 1975 19145 2000
rect 19180 1975 19205 2000
rect 24645 1975 24670 2000
rect 24705 1975 24730 2000
rect 24765 1975 24790 2000
rect 24825 1975 24850 2000
rect 26340 2155 26360 2175
rect 26450 2155 26470 2175
rect 26560 2155 26580 2175
rect 26670 2155 26690 2175
rect 26780 2155 26800 2175
rect 26836 2155 26854 2175
rect 26890 2155 26910 2175
rect 27000 2155 27020 2175
rect 27110 2155 27130 2175
rect 27220 2155 27240 2175
rect 27330 2155 27350 2175
rect 27440 2155 27460 2175
rect 18212 1920 18230 1940
rect 18322 1920 18340 1940
rect 18432 1920 18450 1940
rect 18542 1920 18560 1940
rect 18652 1920 18670 1940
rect 18762 1920 18780 1940
rect 25070 1920 25088 1940
rect 25180 1920 25198 1940
rect 25290 1920 25308 1940
rect 25400 1920 25418 1940
rect 25510 1920 25528 1940
rect 25620 1920 25638 1940
rect 26395 1935 26415 1955
rect 26505 1935 26525 1955
rect 26615 1935 26635 1955
rect 26725 1935 26745 1955
rect 26835 1935 26855 1955
rect 26945 1935 26965 1955
rect 27055 1935 27075 1955
rect 27165 1935 27185 1955
rect 27275 1935 27295 1955
rect 27385 1935 27405 1955
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 28265 2270 28285 2290
rect 28321 2270 28339 2290
rect 28375 2270 28395 2290
rect 28485 2270 28505 2290
rect 28595 2270 28615 2290
rect 28705 2270 28725 2290
rect 3865 1855 3885 1875
rect 4125 1855 4145 1875
rect 4215 1855 4235 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4575 1855 4595 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 4935 1855 4955 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 28212 1900 28230 1920
rect 28322 1900 28340 1920
rect 28432 1900 28450 1920
rect 28542 1900 28560 1920
rect 28652 1900 28670 1920
rect 28762 1900 28780 1920
rect 29070 1955 29095 1980
rect 29130 1955 29155 1980
rect 29190 1955 29215 1980
rect 29250 1955 29275 1980
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4215 1795 4235 1815
rect 4575 1795 4595 1815
rect 4935 1795 4955 1815
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4215 1735 4235 1755
rect 4455 1735 4475 1755
rect 4695 1735 4715 1755
rect 4755 1735 4775 1755
rect 16095 1735 16115 1755
rect 16200 1750 16220 1770
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4335 1690 4355 1710
rect 4575 1690 4595 1710
rect 4815 1690 4835 1710
rect 15115 1680 15135 1700
rect 15315 1680 15335 1700
rect 15416 1680 15434 1700
rect 15515 1680 15535 1700
rect 3995 1630 4015 1650
rect 16315 1735 16335 1755
rect 16420 1750 16440 1770
rect 16243 1690 16260 1710
rect 16535 1735 16555 1755
rect 16650 1750 16670 1770
rect 16463 1690 16480 1710
rect 16610 1690 16627 1710
rect 17135 1735 17155 1755
rect 17240 1750 17260 1770
rect 16825 1690 16845 1710
rect 16876 1690 16893 1710
rect 16955 1690 16975 1710
rect 17355 1735 17375 1755
rect 17460 1750 17480 1770
rect 17283 1690 17300 1710
rect 17575 1735 17595 1755
rect 17690 1750 17710 1770
rect 17503 1690 17520 1710
rect 17650 1690 17667 1710
rect 18315 1680 18335 1700
rect 18416 1680 18434 1700
rect 18515 1680 18535 1700
rect 18715 1680 18735 1700
rect 25115 1680 25135 1700
rect 25315 1680 25335 1700
rect 25416 1680 25434 1700
rect 25515 1680 25535 1700
rect 3175 1570 3195 1590
rect 14825 1615 14850 1640
rect 4815 1570 4835 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4275 1520 4295 1540
rect 4395 1520 4415 1540
rect 4515 1520 4535 1540
rect 4635 1520 4655 1540
rect 4755 1520 4775 1540
rect 2845 1460 2865 1480
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 3925 1460 3945 1480
rect 4065 1460 4085 1480
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 5145 1460 5165 1480
rect 14885 1615 14910 1640
rect 3385 1160 3405 1180
rect 4605 1160 4625 1180
rect 2955 1100 2975 1120
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 3995 1100 4015 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 2915 1015 2935 1035
rect 5120 1015 5140 1035
rect 3005 905 3025 925
rect 3185 905 3205 925
rect 3365 905 3385 925
rect 3545 905 3565 925
rect 3725 905 3745 925
rect 3905 905 3925 925
rect 4085 905 4105 925
rect 4265 905 4285 925
rect 4445 905 4465 925
rect 4625 905 4645 925
rect 4805 905 4825 925
rect 4985 905 5005 925
rect 16112 1470 16129 1490
rect 16315 1470 16335 1490
rect 16535 1470 16555 1490
rect 16830 1470 16850 1490
rect 16880 1470 16900 1490
rect 16928 1470 16945 1490
rect 17152 1470 17169 1490
rect 17355 1470 17375 1490
rect 17575 1470 17595 1490
rect 16155 1410 16175 1430
rect 16260 1410 16280 1430
rect 16370 1410 16390 1430
rect 16480 1410 16500 1430
rect 16590 1410 16610 1430
rect 17195 1410 17215 1430
rect 17300 1410 17320 1430
rect 17410 1410 17430 1430
rect 17520 1410 17540 1430
rect 17630 1410 17650 1430
rect 16325 1210 16345 1230
rect 16435 1210 16455 1230
rect 16545 1210 16565 1230
rect 16655 1210 16675 1230
rect 16765 1210 16785 1230
rect 16820 1210 16840 1230
rect 16875 1210 16895 1230
rect 16985 1210 17005 1230
rect 17095 1210 17115 1230
rect 17205 1210 17225 1230
rect 17315 1210 17335 1230
rect 17425 1210 17445 1230
rect 17535 1210 17555 1230
rect 17605 1225 17625 1245
rect 18940 1615 18965 1640
rect 19000 1615 19025 1640
rect 24825 1615 24850 1640
rect 24885 1615 24910 1640
rect 15215 910 15235 930
rect 15415 910 15435 930
rect 16175 890 16195 910
rect 16270 890 16290 910
rect 16380 890 16400 910
rect 16490 890 16510 910
rect 16600 890 16620 910
rect 16710 890 16730 910
rect 16820 890 16840 910
rect 16930 890 16950 910
rect 17040 890 17060 910
rect 17150 890 17170 910
rect 17260 890 17280 910
rect 17370 890 17390 910
rect 17480 890 17500 910
rect 17630 890 17650 910
rect 18415 910 18435 930
rect 18615 910 18635 930
rect 26095 1735 26115 1755
rect 26200 1750 26220 1770
rect 26315 1735 26335 1755
rect 26420 1750 26440 1770
rect 26243 1690 26260 1710
rect 26535 1735 26555 1755
rect 26650 1750 26670 1770
rect 26463 1690 26480 1710
rect 26610 1690 26627 1710
rect 27135 1735 27155 1755
rect 27240 1750 27260 1770
rect 26825 1690 26845 1710
rect 26876 1690 26893 1710
rect 26955 1690 26975 1710
rect 27355 1735 27375 1755
rect 27460 1750 27480 1770
rect 27283 1690 27300 1710
rect 27575 1735 27595 1755
rect 27690 1750 27710 1770
rect 27503 1690 27520 1710
rect 27650 1690 27667 1710
rect 26112 1470 26129 1490
rect 26315 1470 26335 1490
rect 26535 1470 26555 1490
rect 26830 1470 26850 1490
rect 26880 1470 26900 1490
rect 26928 1470 26945 1490
rect 27152 1470 27169 1490
rect 27355 1470 27375 1490
rect 27575 1470 27595 1490
rect 26155 1410 26175 1430
rect 26260 1410 26280 1430
rect 26370 1410 26390 1430
rect 26480 1410 26500 1430
rect 26590 1410 26610 1430
rect 27195 1410 27215 1430
rect 27300 1410 27320 1430
rect 27410 1410 27430 1430
rect 27520 1410 27540 1430
rect 27630 1410 27650 1430
rect 28315 1680 28335 1700
rect 28416 1680 28434 1700
rect 28515 1680 28535 1700
rect 28715 1680 28735 1700
rect 26325 1110 26345 1130
rect 26435 1110 26455 1130
rect 26545 1110 26565 1130
rect 26655 1110 26675 1130
rect 26765 1110 26785 1130
rect 26820 1110 26840 1130
rect 26875 1110 26895 1130
rect 26985 1110 27005 1130
rect 27095 1110 27115 1130
rect 27205 1110 27225 1130
rect 27315 1110 27335 1130
rect 27425 1110 27445 1130
rect 27535 1110 27555 1130
rect 27605 1125 27625 1145
rect 25215 910 25235 930
rect 25415 910 25435 930
rect 16315 775 16335 795
rect 16385 775 16405 795
rect 16455 775 16475 795
rect 3140 735 3160 755
rect 3275 735 3295 755
rect 3455 735 3475 755
rect 3635 735 3655 755
rect 3815 735 3835 755
rect 3995 735 4015 755
rect 4175 735 4195 755
rect 4355 735 4375 755
rect 4535 735 4555 755
rect 4715 735 4735 755
rect 4895 735 4915 755
rect 16945 775 16965 795
rect 17055 775 17075 795
rect 17165 775 17185 795
rect 17275 775 17295 795
rect 17385 775 17405 795
rect 17495 775 17515 795
rect 26205 790 26225 810
rect 26270 790 26290 810
rect 26380 790 26400 810
rect 26490 790 26510 810
rect 26600 790 26620 810
rect 26710 790 26730 810
rect 26820 790 26840 810
rect 26930 790 26950 810
rect 27040 790 27060 810
rect 27150 790 27170 810
rect 27260 790 27280 810
rect 27370 790 27390 810
rect 27480 790 27500 810
rect 27595 790 27615 810
rect 28415 910 28435 930
rect 28615 910 28635 930
rect 29060 1615 29085 1640
rect 29120 1615 29145 1640
rect 17000 655 17020 675
rect 17110 655 17130 675
rect 17220 655 17240 675
rect 17330 655 17350 675
rect 17440 655 17460 675
rect 26315 575 26335 595
rect 26385 575 26405 595
rect 26455 575 26475 595
rect 26515 575 26535 595
rect 26945 575 26965 595
rect 27055 575 27075 595
rect 27165 575 27185 595
rect 27275 575 27295 595
rect 27385 575 27405 595
rect 27495 575 27515 595
rect 27000 455 27020 475
rect 27110 455 27130 475
rect 27220 455 27240 475
rect 27330 455 27350 475
rect 27440 455 27460 475
<< metal1 >>
rect 26565 4985 26605 4990
rect 26565 4955 26570 4985
rect 26600 4955 26605 4985
rect 26565 4950 26605 4955
rect 26685 4985 26725 4990
rect 26685 4955 26690 4985
rect 26720 4955 26725 4985
rect 26685 4950 26725 4955
rect 26805 4985 26845 4990
rect 26805 4955 26810 4985
rect 26840 4955 26845 4985
rect 26805 4950 26845 4955
rect 27235 4970 27275 4975
rect 26575 4930 26595 4950
rect 26695 4930 26715 4950
rect 26815 4930 26835 4950
rect 27235 4940 27240 4970
rect 27270 4940 27275 4970
rect 27235 4935 27275 4940
rect 26505 4925 26545 4930
rect 26505 4895 26510 4925
rect 26540 4895 26545 4925
rect 26505 4890 26545 4895
rect 26572 4920 26598 4930
rect 26572 4900 26575 4920
rect 26595 4900 26598 4920
rect 26572 4890 26598 4900
rect 26625 4925 26665 4930
rect 26625 4895 26630 4925
rect 26660 4895 26665 4925
rect 26625 4890 26665 4895
rect 26692 4920 26718 4930
rect 26692 4900 26695 4920
rect 26715 4900 26718 4920
rect 26692 4890 26718 4900
rect 26745 4925 26785 4930
rect 26745 4895 26750 4925
rect 26780 4895 26785 4925
rect 26745 4890 26785 4895
rect 26812 4920 26838 4930
rect 26812 4900 26815 4920
rect 26835 4900 26838 4920
rect 26812 4890 26838 4900
rect 26865 4925 26905 4930
rect 26865 4895 26870 4925
rect 26900 4895 26905 4925
rect 27245 4905 27265 4935
rect 26865 4890 26905 4895
rect 27235 4900 27275 4905
rect 27235 4870 27240 4900
rect 27270 4870 27275 4900
rect 27235 4865 27275 4870
rect 27355 4900 27395 4905
rect 27355 4870 27360 4900
rect 27390 4870 27395 4900
rect 27355 4865 27395 4870
rect 27475 4900 27515 4905
rect 27475 4870 27480 4900
rect 27510 4870 27515 4900
rect 27475 4865 27515 4870
rect 27595 4900 27635 4905
rect 27595 4870 27600 4900
rect 27630 4870 27635 4900
rect 27595 4865 27635 4870
rect 27715 4900 27755 4905
rect 27715 4870 27720 4900
rect 27750 4870 27755 4900
rect 27715 4865 27755 4870
rect 26050 4770 26090 4775
rect 26050 4740 26055 4770
rect 26085 4740 26090 4770
rect 26345 4770 26385 4780
rect 26345 4750 26355 4770
rect 26375 4750 26385 4770
rect 26345 4740 26385 4750
rect 26685 4770 26725 4775
rect 26685 4740 26690 4770
rect 26720 4740 26725 4770
rect 26050 4735 26090 4740
rect 16597 4465 16633 4470
rect 16597 4435 16600 4465
rect 16630 4435 16633 4465
rect 16597 4430 16633 4435
rect 16717 4465 16753 4470
rect 16717 4435 16720 4465
rect 16750 4435 16753 4465
rect 16717 4430 16753 4435
rect 16837 4465 16873 4470
rect 16837 4435 16840 4465
rect 16870 4435 16873 4465
rect 16837 4430 16873 4435
rect 17185 4465 17225 4470
rect 17185 4435 17190 4465
rect 17220 4435 17225 4465
rect 17185 4430 17225 4435
rect 16535 4420 16575 4425
rect 16165 4405 16205 4410
rect 16165 4375 16170 4405
rect 16200 4375 16205 4405
rect 16165 4370 16205 4375
rect 16425 4405 16465 4410
rect 16425 4375 16430 4405
rect 16460 4375 16465 4405
rect 16535 4390 16540 4420
rect 16570 4390 16575 4420
rect 16535 4385 16575 4390
rect 16655 4420 16695 4425
rect 16655 4390 16660 4420
rect 16690 4390 16695 4420
rect 16655 4385 16695 4390
rect 16775 4420 16815 4425
rect 16775 4390 16780 4420
rect 16810 4390 16815 4420
rect 16775 4385 16815 4390
rect 16895 4420 16935 4425
rect 16895 4390 16900 4420
rect 16930 4390 16935 4420
rect 17195 4400 17215 4430
rect 16895 4385 16935 4390
rect 17185 4395 17225 4400
rect 16425 4370 16465 4375
rect 17185 4365 17190 4395
rect 17220 4365 17225 4395
rect 17185 4360 17225 4365
rect 17305 4395 17345 4400
rect 17305 4365 17310 4395
rect 17340 4365 17345 4395
rect 17305 4360 17345 4365
rect 17425 4395 17465 4400
rect 17425 4365 17430 4395
rect 17460 4365 17465 4395
rect 17425 4360 17465 4365
rect 17545 4395 17585 4400
rect 17545 4365 17550 4395
rect 17580 4365 17585 4395
rect 17545 4360 17585 4365
rect 17665 4395 17705 4400
rect 17665 4365 17670 4395
rect 17700 4365 17705 4395
rect 17665 4360 17705 4365
rect 16050 4265 16090 4270
rect 16050 4235 16055 4265
rect 16085 4235 16090 4265
rect 16295 4265 16335 4275
rect 16295 4245 16305 4265
rect 16325 4245 16335 4265
rect 16295 4235 16335 4245
rect 16715 4265 16755 4270
rect 16715 4235 16720 4265
rect 16750 4235 16755 4265
rect 16050 4230 16090 4235
rect 14605 3635 14645 3640
rect 14605 3605 14610 3635
rect 14640 3605 14645 3635
rect 14605 3600 14645 3605
rect 15060 3635 15100 3640
rect 15060 3605 15065 3635
rect 15095 3605 15100 3635
rect 15060 3600 15100 3605
rect 15170 3635 15210 3640
rect 15170 3605 15175 3635
rect 15205 3605 15210 3635
rect 15170 3600 15210 3605
rect 15280 3635 15320 3640
rect 15280 3605 15285 3635
rect 15315 3605 15320 3635
rect 15280 3600 15320 3605
rect 15390 3635 15430 3640
rect 15390 3605 15395 3635
rect 15425 3605 15430 3635
rect 15390 3600 15430 3605
rect 15500 3635 15540 3640
rect 15500 3605 15505 3635
rect 15535 3605 15540 3635
rect 15500 3600 15540 3605
rect 15610 3635 15650 3640
rect 15610 3605 15615 3635
rect 15645 3605 15650 3635
rect 15610 3600 15650 3605
rect 14615 3560 14635 3600
rect 14554 3555 14695 3560
rect 1261 3525 1301 3530
rect 1261 3495 1266 3525
rect 1296 3495 1301 3525
rect 14554 3525 14560 3555
rect 14590 3525 14610 3555
rect 14640 3525 14660 3555
rect 14690 3525 14695 3555
rect 14554 3520 14695 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3310 1245 3340
rect 1205 3305 1245 3310
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3255 1200 3285
rect 1160 3250 1200 3255
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 46 3110 51 3145
rect 86 3110 91 3145
rect 1170 3105 1190 3250
rect 1160 3100 1200 3105
rect 1160 3070 1165 3100
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 46 2970 51 3005
rect 86 2970 91 3005
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 1215 2855 1235 3305
rect 1271 3200 1291 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 1271 3140 1291 3165
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 51 2820 56 2855
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2820 769 2855
rect 1205 2850 1245 2855
rect 1205 2820 1210 2850
rect 1240 2820 1245 2850
rect 2340 2840 2360 2860
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 51 2760 56 2795
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2760 769 2795
rect 1271 2750 1291 2805
rect 2330 2800 2370 2805
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2715 1301 2745
rect 1261 2710 1301 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1330 1190 1455 1345
rect 1635 1190 1985 2200
rect 2160 1190 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3135 3340 3175 3345
rect 3135 3310 3140 3340
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 840 2180 1190
rect 2530 765 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3145 3145 3165 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5360 3335 5400 3340
rect 5360 3305 5365 3335
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 4885 3285 4925 3290
rect 4885 3255 4890 3285
rect 4920 3255 4925 3285
rect 4885 3250 4925 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3135 3140 3175 3145
rect 3135 3110 3140 3140
rect 3170 3110 3175 3140
rect 3135 3105 3175 3110
rect 4835 3140 4875 3145
rect 4835 3110 4840 3140
rect 4870 3110 4875 3140
rect 4835 3105 4875 3110
rect 3145 2985 3165 3105
rect 3985 3080 4025 3085
rect 3985 3050 3990 3080
rect 4020 3050 4025 3080
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3005 3485 3035
rect 3445 3000 3485 3005
rect 3805 3035 3845 3040
rect 3805 3005 3810 3035
rect 3840 3005 3845 3035
rect 3805 3000 3845 3005
rect 3455 2985 3475 3000
rect 3815 2985 3835 3000
rect 3995 2985 4015 3045
rect 4345 3035 4385 3040
rect 4345 3005 4350 3035
rect 4380 3005 4385 3035
rect 4345 3000 4385 3005
rect 4705 3035 4745 3040
rect 4705 3005 4710 3035
rect 4740 3005 4745 3035
rect 4705 3000 4745 3005
rect 4355 2985 4375 3000
rect 4715 2985 4735 3000
rect 4845 2985 4865 3105
rect 4895 2985 4915 3250
rect 5315 3140 5355 3145
rect 5315 3110 5320 3140
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 3080 2980 3120 2985
rect 3080 2950 3085 2980
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2950 3305 2980
rect 3265 2945 3305 2950
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2980 3665 2985
rect 3625 2950 3630 2980
rect 3660 2950 3665 2980
rect 3625 2945 3665 2950
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2980 4205 2985
rect 4165 2950 4170 2980
rect 4200 2950 4205 2980
rect 4165 2945 4205 2950
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2980 4565 2985
rect 4525 2950 4530 2980
rect 4560 2950 4565 2980
rect 4525 2945 4565 2950
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 2995 2810 3035 2815
rect 2995 2780 3000 2810
rect 3030 2780 3035 2810
rect 2995 2775 3035 2780
rect 3175 2810 3215 2815
rect 3175 2780 3180 2810
rect 3210 2780 3215 2810
rect 3175 2775 3215 2780
rect 3355 2810 3395 2815
rect 3355 2780 3360 2810
rect 3390 2780 3395 2810
rect 3355 2775 3395 2780
rect 3535 2810 3575 2815
rect 3535 2780 3540 2810
rect 3570 2780 3575 2810
rect 3535 2775 3575 2780
rect 3715 2810 3755 2815
rect 3715 2780 3720 2810
rect 3750 2780 3755 2810
rect 3715 2775 3755 2780
rect 3895 2810 3935 2815
rect 3895 2780 3900 2810
rect 3930 2780 3935 2810
rect 3895 2775 3935 2780
rect 4075 2810 4115 2815
rect 4075 2780 4080 2810
rect 4110 2780 4115 2810
rect 4075 2775 4115 2780
rect 4255 2810 4295 2815
rect 4255 2780 4260 2810
rect 4290 2780 4295 2810
rect 4255 2775 4295 2780
rect 4435 2810 4475 2815
rect 4435 2780 4440 2810
rect 4470 2780 4475 2810
rect 4435 2775 4475 2780
rect 4615 2810 4655 2815
rect 4615 2780 4620 2810
rect 4650 2780 4655 2810
rect 4615 2775 4655 2780
rect 4795 2810 4835 2815
rect 4795 2780 4800 2810
rect 4830 2780 4835 2810
rect 4795 2775 4835 2780
rect 4975 2810 5015 2815
rect 4975 2780 4980 2810
rect 5010 2780 5015 2810
rect 4975 2775 5015 2780
rect 4805 2755 4825 2775
rect 3175 2750 3215 2755
rect 3175 2720 3180 2750
rect 3210 2720 3215 2750
rect 3175 2715 3215 2720
rect 3355 2750 3395 2755
rect 3355 2720 3360 2750
rect 3390 2720 3395 2750
rect 3355 2715 3395 2720
rect 3535 2750 3575 2755
rect 3535 2720 3540 2750
rect 3570 2720 3575 2750
rect 3535 2715 3575 2720
rect 3715 2750 3755 2755
rect 3715 2720 3720 2750
rect 3750 2720 3755 2750
rect 3715 2715 3755 2720
rect 3895 2750 3935 2755
rect 3895 2720 3900 2750
rect 3930 2720 3935 2750
rect 3895 2715 3935 2720
rect 4075 2750 4115 2755
rect 4075 2720 4080 2750
rect 4110 2720 4115 2750
rect 4075 2715 4115 2720
rect 4255 2750 4295 2755
rect 4255 2720 4260 2750
rect 4290 2720 4295 2750
rect 4255 2715 4295 2720
rect 4435 2750 4475 2755
rect 4435 2720 4440 2750
rect 4470 2720 4475 2750
rect 4435 2715 4475 2720
rect 4615 2750 4655 2755
rect 4615 2720 4620 2750
rect 4650 2720 4655 2750
rect 4615 2715 4655 2720
rect 4795 2750 4835 2755
rect 4795 2720 4800 2750
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2375 3395 2380
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3805 2380 3845 2385
rect 3805 2350 3810 2380
rect 3840 2350 3845 2380
rect 3805 2345 3845 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2380 4205 2385
rect 4165 2350 4170 2380
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 3275 2205 3295 2345
rect 3355 2340 3395 2345
rect 3455 2295 3475 2345
rect 3625 2335 3665 2340
rect 3625 2305 3630 2335
rect 3660 2305 3665 2335
rect 3625 2300 3665 2305
rect 3445 2290 3485 2295
rect 3445 2260 3450 2290
rect 3480 2260 3485 2290
rect 3445 2255 3485 2260
rect 3265 2200 3305 2205
rect 3265 2170 3270 2200
rect 3300 2170 3305 2200
rect 3265 2165 3305 2170
rect 3635 2155 3655 2300
rect 3815 2250 3835 2345
rect 3805 2245 3845 2250
rect 3805 2215 3810 2245
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 3625 2150 3665 2155
rect 3625 2120 3630 2150
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2065 2785 2095
rect 2745 2060 2785 2065
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3995 2205 4015 2345
rect 4345 2335 4385 2340
rect 4345 2305 4350 2335
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 4535 2295 4555 2345
rect 4525 2290 4565 2295
rect 4525 2260 4530 2290
rect 4560 2260 4565 2290
rect 4525 2255 4565 2260
rect 4715 2205 4735 2345
rect 5270 2290 5310 2295
rect 5270 2260 5275 2290
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 3985 2200 4025 2205
rect 3985 2170 3990 2200
rect 4020 2170 4025 2200
rect 3985 2165 4025 2170
rect 4705 2200 4745 2205
rect 4705 2170 4710 2200
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2115 4125 2145
rect 4085 2110 4125 2115
rect 3985 2095 4025 2100
rect 3985 2065 3990 2095
rect 4020 2065 4025 2095
rect 3985 2060 4025 2065
rect 4095 2055 4115 2110
rect 4145 2095 4185 2100
rect 4145 2065 4150 2095
rect 4180 2065 4185 2095
rect 4145 2060 4185 2065
rect 4265 2095 4305 2100
rect 4265 2065 4270 2095
rect 4300 2065 4305 2095
rect 4265 2060 4305 2065
rect 4385 2095 4425 2100
rect 4385 2065 4390 2095
rect 4420 2065 4425 2095
rect 4385 2060 4425 2065
rect 4505 2095 4545 2100
rect 4505 2065 4510 2095
rect 4540 2065 4545 2095
rect 4505 2060 4545 2065
rect 4625 2095 4665 2100
rect 4625 2065 4630 2095
rect 4660 2065 4665 2095
rect 4625 2060 4665 2065
rect 4745 2095 4785 2100
rect 4745 2065 4750 2095
rect 4780 2065 4785 2095
rect 4745 2060 4785 2065
rect 4865 2095 4905 2100
rect 4865 2065 4870 2095
rect 4900 2065 4905 2095
rect 4865 2060 4905 2065
rect 4985 2095 5025 2100
rect 4985 2065 4990 2095
rect 5020 2065 5025 2095
rect 4985 2060 5025 2065
rect 5105 2095 5145 2100
rect 5105 2065 5110 2095
rect 5140 2065 5145 2095
rect 5105 2060 5145 2065
rect 5225 2095 5265 2100
rect 5225 2065 5230 2095
rect 5260 2065 5265 2095
rect 5225 2060 5265 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3925 2055
rect 3885 2020 3890 2050
rect 3920 2045 3925 2050
rect 4085 2050 4125 2055
rect 4085 2045 4090 2050
rect 3920 2020 3945 2045
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 2800 1765 2840 1770
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2800 1735 2805 1765
rect 2835 1735 2840 1765
rect 2800 1730 2840 1735
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 2810 1715 2830 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 2800 1710 2840 1715
rect 2800 1680 2805 1710
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2800 1675 2840 1680
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1045 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1490 2865 1510
rect 2925 1500 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1470 2930 1500
rect 2960 1470 2965 1500
rect 2925 1465 2965 1470
rect 3045 1500 3085 1505
rect 3045 1470 3050 1500
rect 3080 1470 3085 1500
rect 3045 1465 3085 1470
rect 3165 1500 3205 1505
rect 3165 1470 3170 1500
rect 3200 1470 3205 1500
rect 3165 1465 3205 1470
rect 3285 1500 3325 1505
rect 3285 1470 3290 1500
rect 3320 1470 3325 1500
rect 3285 1465 3325 1470
rect 3525 1500 3565 1505
rect 3525 1470 3530 1500
rect 3560 1470 3565 1500
rect 3525 1465 3565 1470
rect 3645 1500 3685 1505
rect 3645 1470 3650 1500
rect 3680 1470 3685 1500
rect 3645 1465 3685 1470
rect 3765 1500 3805 1505
rect 3765 1470 3770 1500
rect 3800 1470 3805 1500
rect 3925 1490 3945 2015
rect 4065 2020 4090 2045
rect 4120 2020 4125 2050
rect 4065 2015 4125 2020
rect 4445 2050 4485 2055
rect 4445 2020 4450 2050
rect 4480 2020 4485 2050
rect 4445 2015 4485 2020
rect 4805 2050 4845 2055
rect 4805 2020 4810 2050
rect 4840 2020 4845 2050
rect 4805 2015 4845 2020
rect 5165 2050 5205 2055
rect 5165 2020 5170 2050
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 3765 1465 3805 1470
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 3995 1190 4015 1620
rect 4065 1490 4085 2015
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1850 4365 1880
rect 4325 1845 4365 1850
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1880 4725 1885
rect 4685 1850 4690 1880
rect 4720 1850 4725 1880
rect 4685 1845 4725 1850
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1880 5085 1885
rect 5045 1850 5050 1880
rect 5080 1850 5085 1880
rect 5045 1845 5085 1850
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 4125 1825 4145 1845
rect 4215 1825 4235 1845
rect 4455 1825 4475 1845
rect 4575 1825 4595 1845
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1790 4155 1820
rect 4115 1785 4155 1790
rect 4205 1820 4245 1825
rect 4205 1790 4210 1820
rect 4240 1790 4245 1820
rect 4205 1785 4245 1790
rect 4445 1820 4485 1825
rect 4445 1790 4450 1820
rect 4480 1790 4485 1820
rect 4445 1785 4485 1790
rect 4565 1820 4605 1825
rect 4565 1790 4570 1820
rect 4600 1790 4605 1820
rect 4565 1785 4605 1790
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1730 4245 1760
rect 4205 1725 4245 1730
rect 4445 1760 4485 1765
rect 4445 1730 4450 1760
rect 4480 1730 4485 1760
rect 4445 1725 4485 1730
rect 4575 1720 4595 1785
rect 4695 1765 4715 1845
rect 4815 1825 4835 1845
rect 4935 1825 4955 1845
rect 5145 1825 5165 1845
rect 4805 1820 4845 1825
rect 4805 1790 4810 1820
rect 4840 1790 4845 1820
rect 4805 1785 4845 1790
rect 4925 1820 4965 1825
rect 4925 1790 4930 1820
rect 4960 1790 4965 1820
rect 4925 1785 4965 1790
rect 5135 1820 5175 1825
rect 5135 1790 5140 1820
rect 5170 1790 5175 1820
rect 5135 1785 5175 1790
rect 5280 1765 5300 2255
rect 5325 2150 5345 3105
rect 5315 2145 5355 2150
rect 5315 2115 5320 2145
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 5370 1825 5390 3300
rect 5410 3285 5450 3290
rect 5410 3255 5415 3285
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 5360 1820 5400 1825
rect 5360 1790 5365 1820
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1730 4785 1760
rect 4745 1725 4785 1730
rect 5270 1760 5310 1765
rect 5270 1730 5275 1760
rect 5305 1730 5310 1760
rect 5270 1725 5310 1730
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1685 4365 1715
rect 4325 1680 4365 1685
rect 4565 1715 4605 1720
rect 4565 1685 4570 1715
rect 4600 1685 4605 1715
rect 4565 1680 4605 1685
rect 4805 1715 4845 1720
rect 4805 1685 4810 1715
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 5420 1600 5440 3250
rect 16060 3110 16080 4230
rect 16305 4215 16325 4235
rect 16715 4230 16755 4235
rect 17245 4265 17285 4270
rect 17245 4235 17250 4265
rect 17280 4235 17285 4265
rect 17245 4230 17285 4235
rect 17308 4260 17342 4270
rect 17308 4240 17316 4260
rect 17334 4240 17342 4260
rect 17308 4230 17342 4240
rect 17365 4265 17405 4270
rect 17365 4235 17370 4265
rect 17400 4235 17405 4265
rect 17365 4230 17405 4235
rect 17485 4265 17525 4270
rect 17485 4235 17490 4265
rect 17520 4235 17525 4265
rect 17485 4230 17525 4235
rect 17605 4265 17645 4270
rect 17605 4235 17610 4265
rect 17640 4235 17645 4265
rect 17605 4230 17645 4235
rect 17315 4215 17335 4230
rect 16105 4210 16145 4215
rect 16105 4180 16110 4210
rect 16140 4180 16145 4210
rect 16105 4175 16145 4180
rect 16295 4210 16335 4215
rect 16295 4180 16300 4210
rect 16330 4180 16335 4210
rect 16295 4175 16335 4180
rect 17305 4210 17345 4215
rect 17305 4180 17310 4210
rect 17340 4180 17345 4210
rect 17305 4175 17345 4180
rect 16050 3105 16090 3110
rect 16050 3075 16055 3105
rect 16085 3075 16090 3105
rect 16050 3070 16090 3075
rect 15115 2965 15155 2970
rect 14554 2935 14695 2940
rect 14554 2905 14560 2935
rect 14590 2905 14610 2935
rect 14640 2905 14660 2935
rect 14690 2905 14695 2935
rect 15115 2935 15120 2965
rect 15150 2935 15155 2965
rect 15115 2930 15155 2935
rect 15225 2965 15265 2970
rect 15225 2935 15230 2965
rect 15260 2935 15265 2965
rect 15225 2930 15265 2935
rect 15335 2965 15375 2970
rect 15335 2935 15340 2965
rect 15370 2935 15375 2965
rect 15335 2930 15375 2935
rect 15445 2965 15485 2970
rect 15445 2935 15450 2965
rect 15480 2935 15485 2965
rect 15445 2930 15485 2935
rect 15503 2960 15537 2970
rect 15503 2940 15511 2960
rect 15529 2940 15537 2960
rect 15503 2930 15537 2940
rect 15555 2965 15595 2970
rect 15555 2935 15560 2965
rect 15590 2935 15595 2965
rect 16115 2955 16135 4175
rect 16360 4155 16400 4160
rect 16360 4125 16365 4155
rect 16395 4125 16400 4155
rect 16360 4120 16400 4125
rect 16470 4155 16510 4160
rect 16470 4125 16475 4155
rect 16505 4125 16510 4155
rect 16470 4120 16510 4125
rect 16580 4155 16620 4160
rect 16580 4125 16585 4155
rect 16615 4125 16620 4155
rect 16580 4120 16620 4125
rect 16690 4155 16730 4160
rect 16690 4125 16695 4155
rect 16725 4125 16730 4155
rect 16690 4120 16730 4125
rect 16800 4155 16840 4160
rect 16800 4125 16805 4155
rect 16835 4125 16840 4155
rect 16800 4120 16840 4125
rect 16910 4155 16950 4160
rect 16910 4125 16915 4155
rect 16945 4125 16950 4155
rect 16910 4120 16950 4125
rect 17020 4155 17060 4160
rect 17020 4125 17025 4155
rect 17055 4125 17060 4155
rect 17020 4120 17060 4125
rect 17130 4155 17170 4160
rect 17130 4125 17135 4155
rect 17165 4125 17170 4155
rect 17130 4120 17170 4125
rect 17240 4155 17280 4160
rect 17240 4125 17245 4155
rect 17275 4125 17280 4155
rect 17240 4120 17280 4125
rect 17350 4155 17390 4160
rect 17350 4125 17355 4155
rect 17385 4125 17390 4155
rect 17350 4120 17390 4125
rect 16305 4035 16345 4040
rect 16305 4005 16310 4035
rect 16340 4005 16345 4035
rect 16305 4000 16345 4005
rect 16362 4030 16398 4040
rect 16362 4010 16370 4030
rect 16390 4010 16398 4030
rect 16362 4000 16398 4010
rect 16415 4030 16455 4040
rect 16415 4010 16425 4030
rect 16445 4010 16455 4030
rect 16415 4000 16455 4010
rect 16525 4035 16565 4040
rect 16525 4005 16530 4035
rect 16560 4005 16565 4035
rect 16525 4000 16565 4005
rect 16635 4030 16675 4040
rect 16635 4010 16645 4030
rect 16665 4010 16675 4030
rect 16635 4000 16675 4010
rect 16745 4035 16785 4040
rect 16745 4005 16750 4035
rect 16780 4005 16785 4035
rect 16745 4000 16785 4005
rect 16855 4030 16895 4040
rect 16855 4010 16865 4030
rect 16885 4010 16895 4030
rect 16855 4000 16895 4010
rect 16965 4035 17005 4040
rect 16965 4005 16970 4035
rect 17000 4005 17005 4035
rect 16965 4000 17005 4005
rect 17075 4030 17115 4040
rect 17075 4010 17085 4030
rect 17105 4010 17115 4030
rect 17075 4000 17115 4010
rect 17185 4035 17225 4040
rect 17185 4005 17190 4035
rect 17220 4005 17225 4035
rect 17185 4000 17225 4005
rect 17295 4030 17335 4040
rect 17295 4010 17305 4030
rect 17325 4010 17335 4030
rect 17295 4000 17335 4010
rect 17405 4035 17445 4040
rect 17405 4005 17410 4035
rect 17440 4005 17445 4035
rect 17405 4000 17445 4005
rect 16310 3910 16350 3915
rect 16310 3880 16315 3910
rect 16345 3880 16350 3910
rect 16310 3875 16350 3880
rect 16370 3855 16390 4000
rect 16425 3980 16445 4000
rect 16645 3980 16665 4000
rect 16865 3980 16885 4000
rect 17085 3980 17105 4000
rect 17305 3980 17325 4000
rect 16415 3975 16455 3980
rect 16415 3945 16420 3975
rect 16450 3945 16455 3975
rect 16415 3940 16455 3945
rect 16635 3975 16675 3980
rect 16635 3945 16640 3975
rect 16670 3945 16675 3975
rect 16635 3940 16675 3945
rect 16855 3975 16895 3980
rect 16855 3945 16860 3975
rect 16890 3945 16895 3975
rect 16855 3940 16895 3945
rect 17075 3975 17115 3980
rect 17075 3945 17080 3975
rect 17110 3945 17115 3975
rect 17075 3940 17115 3945
rect 17295 3975 17335 3980
rect 17295 3945 17300 3975
rect 17330 3945 17335 3975
rect 17295 3940 17335 3945
rect 16425 3915 16445 3940
rect 17415 3915 17435 4000
rect 16415 3910 16455 3915
rect 16415 3880 16420 3910
rect 16450 3880 16455 3910
rect 16415 3875 16455 3880
rect 16525 3910 16565 3915
rect 16525 3880 16530 3910
rect 16560 3880 16565 3910
rect 16525 3875 16565 3880
rect 16635 3910 16675 3915
rect 16635 3880 16640 3910
rect 16670 3880 16675 3910
rect 16635 3875 16675 3880
rect 16745 3910 16785 3915
rect 16745 3880 16750 3910
rect 16780 3880 16785 3910
rect 16745 3875 16785 3880
rect 17050 3910 17090 3915
rect 17050 3880 17055 3910
rect 17085 3880 17090 3910
rect 17050 3875 17090 3880
rect 17155 3910 17195 3915
rect 17155 3880 17160 3910
rect 17190 3880 17195 3910
rect 17155 3875 17195 3880
rect 17265 3910 17305 3915
rect 17265 3880 17270 3910
rect 17300 3880 17305 3910
rect 17265 3875 17305 3880
rect 17375 3910 17435 3915
rect 17375 3880 17380 3910
rect 17410 3880 17435 3910
rect 17375 3875 17435 3880
rect 17485 3910 17525 3915
rect 17485 3880 17490 3910
rect 17520 3880 17525 3910
rect 17485 3875 17525 3880
rect 16271 3850 16303 3855
rect 16271 3820 16274 3850
rect 16300 3820 16303 3850
rect 16271 3815 16303 3820
rect 16360 3845 16400 3855
rect 16360 3825 16370 3845
rect 16390 3825 16400 3845
rect 16360 3815 16400 3825
rect 16470 3850 16510 3855
rect 16470 3820 16475 3850
rect 16505 3820 16510 3850
rect 16470 3815 16510 3820
rect 16690 3850 16730 3855
rect 16690 3820 16695 3850
rect 16725 3820 16730 3850
rect 16690 3815 16730 3820
rect 16800 3845 16840 3855
rect 16800 3825 16810 3845
rect 16830 3825 16840 3845
rect 16800 3815 16840 3825
rect 17011 3850 17043 3855
rect 17011 3820 17014 3850
rect 17040 3820 17043 3850
rect 17011 3815 17043 3820
rect 17210 3850 17250 3855
rect 17210 3820 17215 3850
rect 17245 3820 17250 3850
rect 17210 3815 17250 3820
rect 17430 3850 17470 3855
rect 17430 3820 17435 3850
rect 17465 3820 17470 3850
rect 17430 3815 17470 3820
rect 17860 3850 17900 3855
rect 17860 3820 17865 3850
rect 17895 3820 17900 3850
rect 17860 3815 17900 3820
rect 16402 3730 16434 3735
rect 16402 3700 16405 3730
rect 16431 3700 16434 3730
rect 16402 3695 16434 3700
rect 16622 3730 16654 3735
rect 16622 3700 16625 3730
rect 16651 3700 16654 3730
rect 16622 3695 16654 3700
rect 16766 3730 16798 3735
rect 16766 3700 16769 3730
rect 16795 3700 16798 3730
rect 16766 3695 16798 3700
rect 17142 3730 17174 3735
rect 17142 3700 17145 3730
rect 17171 3700 17174 3730
rect 17142 3695 17174 3700
rect 17362 3730 17394 3735
rect 17362 3700 17365 3730
rect 17391 3700 17394 3730
rect 17362 3695 17394 3700
rect 17506 3730 17538 3735
rect 17506 3700 17509 3730
rect 17535 3700 17538 3730
rect 17506 3695 17538 3700
rect 16990 3680 17030 3685
rect 16250 3670 16290 3675
rect 16250 3640 16255 3670
rect 16285 3640 16290 3670
rect 16250 3635 16290 3640
rect 16355 3670 16395 3675
rect 16355 3640 16360 3670
rect 16390 3640 16395 3670
rect 16355 3635 16395 3640
rect 16470 3670 16510 3675
rect 16470 3640 16475 3670
rect 16505 3640 16510 3670
rect 16470 3635 16510 3640
rect 16575 3670 16615 3675
rect 16575 3640 16580 3670
rect 16610 3640 16615 3670
rect 16575 3635 16615 3640
rect 16690 3670 16730 3675
rect 16690 3640 16695 3670
rect 16725 3640 16730 3670
rect 16690 3635 16730 3640
rect 16805 3670 16845 3675
rect 16805 3640 16810 3670
rect 16840 3640 16845 3670
rect 16990 3650 16995 3680
rect 17025 3650 17030 3680
rect 16990 3645 17030 3650
rect 17210 3680 17250 3685
rect 17210 3650 17215 3680
rect 17245 3650 17250 3680
rect 17210 3645 17250 3650
rect 17430 3680 17470 3685
rect 17430 3650 17435 3680
rect 17465 3650 17470 3680
rect 17430 3645 17470 3650
rect 16805 3635 16845 3640
rect 17095 3635 17135 3640
rect 17095 3605 17100 3635
rect 17130 3605 17135 3635
rect 17095 3600 17135 3605
rect 17315 3635 17355 3640
rect 17315 3605 17320 3635
rect 17350 3605 17355 3635
rect 17315 3600 17355 3605
rect 17545 3635 17585 3640
rect 17545 3605 17550 3635
rect 17580 3605 17585 3635
rect 17545 3600 17585 3605
rect 16340 3575 16380 3580
rect 16340 3545 16345 3575
rect 16375 3545 16380 3575
rect 16340 3540 16380 3545
rect 16460 3575 16500 3580
rect 16460 3545 16465 3575
rect 16495 3545 16500 3575
rect 16460 3540 16500 3545
rect 16580 3575 16620 3580
rect 16580 3545 16585 3575
rect 16615 3545 16620 3575
rect 16580 3540 16620 3545
rect 16700 3575 16740 3580
rect 16700 3545 16705 3575
rect 16735 3545 16740 3575
rect 16700 3540 16740 3545
rect 16820 3575 16860 3580
rect 16820 3545 16825 3575
rect 16855 3545 16860 3575
rect 16820 3540 16860 3545
rect 16940 3575 16980 3580
rect 16940 3545 16945 3575
rect 16975 3545 16980 3575
rect 16940 3540 16980 3545
rect 17060 3575 17100 3580
rect 17060 3545 17065 3575
rect 17095 3545 17100 3575
rect 17060 3540 17100 3545
rect 17180 3575 17220 3580
rect 17180 3545 17185 3575
rect 17215 3545 17220 3575
rect 17180 3540 17220 3545
rect 17300 3575 17340 3580
rect 17300 3545 17305 3575
rect 17335 3545 17340 3575
rect 17300 3540 17340 3545
rect 17420 3575 17460 3580
rect 17420 3545 17425 3575
rect 17455 3545 17460 3575
rect 17420 3540 17460 3545
rect 16280 3100 16320 3110
rect 16280 3080 16290 3100
rect 16310 3080 16320 3100
rect 16280 3070 16320 3080
rect 16400 3100 16440 3110
rect 16400 3080 16410 3100
rect 16430 3080 16440 3100
rect 16400 3070 16440 3080
rect 16520 3100 16560 3110
rect 16520 3080 16530 3100
rect 16550 3080 16560 3100
rect 16520 3070 16560 3080
rect 16640 3100 16680 3110
rect 16640 3080 16650 3100
rect 16670 3080 16680 3100
rect 16640 3070 16680 3080
rect 16760 3100 16800 3110
rect 16760 3080 16770 3100
rect 16790 3080 16800 3100
rect 16760 3070 16800 3080
rect 16823 3105 16857 3110
rect 16823 3075 16826 3105
rect 16854 3075 16857 3105
rect 16823 3070 16857 3075
rect 16880 3100 16920 3110
rect 16880 3080 16890 3100
rect 16910 3080 16920 3100
rect 16880 3070 16920 3080
rect 17000 3100 17040 3110
rect 17000 3080 17010 3100
rect 17030 3080 17040 3100
rect 17000 3070 17040 3080
rect 17120 3100 17160 3110
rect 17120 3080 17130 3100
rect 17150 3080 17160 3100
rect 17120 3070 17160 3080
rect 17240 3100 17280 3110
rect 17240 3080 17250 3100
rect 17270 3080 17280 3100
rect 17240 3070 17280 3080
rect 17360 3100 17400 3110
rect 17360 3080 17370 3100
rect 17390 3080 17400 3100
rect 17360 3070 17400 3080
rect 17480 3100 17520 3110
rect 17480 3080 17490 3100
rect 17510 3080 17520 3100
rect 17480 3070 17520 3080
rect 16290 3055 16310 3070
rect 16280 3050 16320 3055
rect 16280 3020 16285 3050
rect 16315 3020 16320 3050
rect 16280 3015 16320 3020
rect 16410 3010 16430 3070
rect 16530 3055 16550 3070
rect 16520 3050 16560 3055
rect 16520 3020 16525 3050
rect 16555 3020 16560 3050
rect 16520 3015 16560 3020
rect 16650 3010 16670 3070
rect 16770 3055 16790 3070
rect 16760 3050 16800 3055
rect 16760 3020 16765 3050
rect 16795 3020 16800 3050
rect 16760 3015 16800 3020
rect 16890 3010 16910 3070
rect 17010 3055 17030 3070
rect 17000 3050 17040 3055
rect 17000 3020 17005 3050
rect 17035 3020 17040 3050
rect 17000 3015 17040 3020
rect 17130 3010 17150 3070
rect 17250 3055 17270 3070
rect 17240 3050 17280 3055
rect 17240 3020 17245 3050
rect 17275 3020 17280 3050
rect 17240 3015 17280 3020
rect 17370 3010 17390 3070
rect 17490 3055 17510 3070
rect 17480 3050 17520 3055
rect 17480 3020 17485 3050
rect 17515 3020 17520 3050
rect 17480 3015 17520 3020
rect 16400 3005 16440 3010
rect 16400 2975 16405 3005
rect 16435 2975 16440 3005
rect 16400 2970 16440 2975
rect 16640 3005 16680 3010
rect 16640 2975 16645 3005
rect 16675 2975 16680 3005
rect 16640 2970 16680 2975
rect 16880 3005 16920 3010
rect 16880 2975 16885 3005
rect 16915 2975 16920 3005
rect 16880 2970 16920 2975
rect 17120 3005 17160 3010
rect 17120 2975 17125 3005
rect 17155 2975 17160 3005
rect 17120 2970 17160 2975
rect 17360 3005 17400 3010
rect 17360 2975 17365 3005
rect 17395 2975 17400 3005
rect 17360 2970 17400 2975
rect 15555 2930 15595 2935
rect 16105 2950 16145 2955
rect 14554 2900 14695 2905
rect 14615 2885 14635 2900
rect 14605 2880 14645 2885
rect 14605 2850 14610 2880
rect 14640 2850 14645 2880
rect 14605 2845 14645 2850
rect 15235 2830 15255 2930
rect 15510 2885 15530 2930
rect 16105 2920 16110 2950
rect 16140 2920 16145 2950
rect 16105 2915 16145 2920
rect 16400 2900 16415 2970
rect 16880 2950 16920 2955
rect 16880 2920 16885 2950
rect 16915 2920 16920 2950
rect 16880 2915 16920 2920
rect 16135 2895 16175 2900
rect 15500 2880 15540 2885
rect 15500 2850 15505 2880
rect 15535 2850 15540 2880
rect 15500 2845 15540 2850
rect 15780 2880 15820 2885
rect 15780 2850 15785 2880
rect 15815 2850 15820 2880
rect 16135 2865 16140 2895
rect 16170 2865 16175 2895
rect 16135 2860 16175 2865
rect 16255 2895 16295 2900
rect 16255 2865 16260 2895
rect 16290 2865 16295 2895
rect 16255 2860 16295 2865
rect 16375 2895 16415 2900
rect 16375 2865 16380 2895
rect 16410 2865 16415 2895
rect 16375 2860 16415 2865
rect 16495 2895 16535 2900
rect 16495 2865 16500 2895
rect 16530 2865 16535 2895
rect 16495 2860 16535 2865
rect 16615 2895 16655 2900
rect 16615 2865 16620 2895
rect 16650 2865 16655 2895
rect 16615 2860 16655 2865
rect 15780 2845 15820 2850
rect 14515 2825 14555 2830
rect 14515 2795 14520 2825
rect 14550 2795 14555 2825
rect 14515 2790 14555 2795
rect 15225 2825 15265 2830
rect 15225 2795 15230 2825
rect 15260 2795 15265 2825
rect 15225 2790 15265 2795
rect 14525 2120 14545 2790
rect 15060 2705 15100 2710
rect 15060 2675 15065 2705
rect 15095 2675 15100 2705
rect 15060 2670 15100 2675
rect 15170 2705 15210 2710
rect 15170 2675 15175 2705
rect 15205 2675 15210 2705
rect 15170 2670 15210 2675
rect 15280 2705 15320 2710
rect 15280 2675 15285 2705
rect 15315 2675 15320 2705
rect 15280 2670 15320 2675
rect 15390 2705 15430 2710
rect 15390 2675 15395 2705
rect 15425 2675 15430 2705
rect 15390 2670 15430 2675
rect 15500 2705 15540 2710
rect 15500 2675 15505 2705
rect 15535 2675 15540 2705
rect 15500 2670 15540 2675
rect 15610 2705 15650 2710
rect 15610 2675 15615 2705
rect 15645 2675 15650 2705
rect 15610 2670 15650 2675
rect 14870 2435 14910 2440
rect 14870 2405 14875 2435
rect 14905 2405 14910 2435
rect 14870 2400 14910 2405
rect 15115 2435 15155 2440
rect 15115 2405 15120 2435
rect 15150 2405 15155 2435
rect 15115 2400 15155 2405
rect 15225 2435 15265 2440
rect 15225 2405 15230 2435
rect 15260 2405 15265 2435
rect 15225 2400 15265 2405
rect 15335 2435 15375 2440
rect 15335 2405 15340 2435
rect 15370 2405 15375 2435
rect 15335 2400 15375 2405
rect 15445 2435 15485 2440
rect 15445 2405 15450 2435
rect 15480 2405 15485 2435
rect 15445 2400 15485 2405
rect 15555 2435 15595 2440
rect 15555 2405 15560 2435
rect 15590 2405 15595 2435
rect 15555 2400 15595 2405
rect 14510 2110 14560 2120
rect 14510 2080 14520 2110
rect 14550 2080 14560 2110
rect 14510 2070 14560 2080
rect 14525 1710 14545 2070
rect 14640 2005 14675 2011
rect 14640 1965 14675 1970
rect 14700 2005 14735 2010
rect 14700 1965 14735 1970
rect 14760 2005 14795 2011
rect 14760 1965 14795 1970
rect 14820 2005 14855 2010
rect 14880 2005 14900 2400
rect 15790 2380 15810 2845
rect 16075 2475 16115 2480
rect 16075 2445 16080 2475
rect 16110 2445 16115 2475
rect 16075 2440 16115 2445
rect 16195 2475 16235 2480
rect 16195 2445 16200 2475
rect 16230 2445 16235 2475
rect 16195 2440 16235 2445
rect 16315 2475 16355 2480
rect 16315 2445 16320 2475
rect 16350 2445 16355 2475
rect 16315 2440 16355 2445
rect 16378 2470 16412 2480
rect 16378 2450 16386 2470
rect 16404 2450 16412 2470
rect 16378 2440 16412 2450
rect 16435 2475 16475 2480
rect 16435 2445 16440 2475
rect 16470 2445 16475 2475
rect 16435 2440 16475 2445
rect 16555 2475 16595 2480
rect 16555 2445 16560 2475
rect 16590 2445 16595 2475
rect 16555 2440 16595 2445
rect 16675 2475 16715 2480
rect 16675 2445 16680 2475
rect 16710 2445 16715 2475
rect 16675 2440 16715 2445
rect 16330 2380 16350 2440
rect 16385 2425 16405 2440
rect 16890 2425 16910 2915
rect 17505 2900 17520 3015
rect 17145 2895 17185 2900
rect 17145 2865 17150 2895
rect 17180 2865 17185 2895
rect 17145 2860 17185 2865
rect 17265 2895 17305 2900
rect 17265 2865 17270 2895
rect 17300 2865 17305 2895
rect 17265 2860 17305 2865
rect 17385 2895 17425 2900
rect 17385 2865 17390 2895
rect 17420 2865 17425 2895
rect 17385 2860 17425 2865
rect 17505 2895 17545 2900
rect 17505 2865 17510 2895
rect 17540 2865 17545 2895
rect 17505 2860 17545 2865
rect 17625 2895 17665 2900
rect 17625 2865 17630 2895
rect 17660 2865 17665 2895
rect 17625 2860 17665 2865
rect 17085 2475 17125 2480
rect 17085 2445 17090 2475
rect 17120 2445 17125 2475
rect 17085 2440 17125 2445
rect 17205 2475 17245 2480
rect 17205 2445 17210 2475
rect 17240 2445 17245 2475
rect 17205 2440 17245 2445
rect 17325 2475 17365 2480
rect 17325 2445 17330 2475
rect 17360 2445 17365 2475
rect 17325 2440 17365 2445
rect 17388 2470 17422 2480
rect 17388 2450 17396 2470
rect 17414 2450 17422 2470
rect 17388 2440 17422 2450
rect 17445 2475 17485 2480
rect 17445 2445 17450 2475
rect 17480 2445 17485 2475
rect 17445 2440 17485 2445
rect 17565 2475 17605 2480
rect 17565 2445 17570 2475
rect 17600 2445 17605 2475
rect 17565 2440 17605 2445
rect 17685 2475 17725 2480
rect 17685 2445 17690 2475
rect 17720 2445 17725 2475
rect 17685 2440 17725 2445
rect 16375 2420 16415 2425
rect 16375 2390 16380 2420
rect 16410 2390 16415 2420
rect 16375 2385 16415 2390
rect 16880 2420 16920 2425
rect 16880 2390 16885 2420
rect 16915 2390 16920 2420
rect 16880 2385 16920 2390
rect 17330 2380 17350 2440
rect 17395 2425 17415 2440
rect 17385 2420 17425 2425
rect 17385 2390 17390 2420
rect 17420 2390 17425 2420
rect 17385 2385 17425 2390
rect 15585 2375 15625 2380
rect 15585 2345 15590 2375
rect 15620 2345 15625 2375
rect 15585 2340 15625 2345
rect 15780 2375 15820 2380
rect 15780 2345 15785 2375
rect 15815 2345 15820 2375
rect 15780 2340 15820 2345
rect 16320 2375 16360 2380
rect 16320 2345 16325 2375
rect 16355 2345 16360 2375
rect 16320 2340 16360 2345
rect 17320 2375 17360 2380
rect 17320 2345 17325 2375
rect 17355 2345 17360 2375
rect 17320 2340 17360 2345
rect 16000 2325 16040 2330
rect 14915 2315 14955 2320
rect 14915 2285 14920 2315
rect 14950 2285 14955 2315
rect 14915 2280 14955 2285
rect 15115 2315 15155 2320
rect 15115 2285 15120 2315
rect 15150 2285 15155 2315
rect 15115 2280 15155 2285
rect 15225 2315 15265 2320
rect 15225 2285 15230 2315
rect 15260 2285 15265 2315
rect 15225 2280 15265 2285
rect 15335 2315 15375 2320
rect 15335 2285 15340 2315
rect 15370 2285 15375 2315
rect 15335 2280 15375 2285
rect 15445 2315 15485 2320
rect 15445 2285 15450 2315
rect 15480 2285 15485 2315
rect 15445 2280 15485 2285
rect 15555 2315 15595 2320
rect 15555 2285 15560 2315
rect 15590 2285 15595 2315
rect 16000 2295 16005 2325
rect 16035 2295 16040 2325
rect 16000 2290 16040 2295
rect 15555 2280 15595 2285
rect 14820 1965 14855 1970
rect 14870 2000 14910 2005
rect 14870 1970 14875 2000
rect 14905 1970 14910 2000
rect 14870 1965 14910 1970
rect 14650 1900 14670 1965
rect 14770 1950 14790 1965
rect 14925 1950 14945 2280
rect 15800 2180 15840 2185
rect 15800 2150 15805 2180
rect 15835 2150 15840 2180
rect 15800 2145 15840 2150
rect 14760 1945 14800 1950
rect 14760 1915 14765 1945
rect 14795 1915 14800 1945
rect 14760 1910 14800 1915
rect 14915 1945 14955 1950
rect 14915 1915 14920 1945
rect 14950 1915 14955 1945
rect 14915 1910 14955 1915
rect 15060 1945 15100 1950
rect 15060 1915 15065 1945
rect 15095 1915 15100 1945
rect 15060 1910 15100 1915
rect 15170 1945 15210 1950
rect 15170 1915 15175 1945
rect 15205 1915 15210 1945
rect 15170 1910 15210 1915
rect 15280 1945 15320 1950
rect 15280 1915 15285 1945
rect 15315 1915 15320 1945
rect 15280 1910 15320 1915
rect 15390 1945 15430 1950
rect 15390 1915 15395 1945
rect 15425 1915 15430 1945
rect 15390 1910 15430 1915
rect 15500 1945 15540 1950
rect 15500 1915 15505 1945
rect 15535 1915 15540 1945
rect 15500 1910 15540 1915
rect 15610 1945 15650 1950
rect 15610 1915 15615 1945
rect 15645 1915 15650 1945
rect 15610 1910 15650 1915
rect 14640 1895 14680 1900
rect 14640 1865 14645 1895
rect 14675 1865 14680 1895
rect 14640 1860 14680 1865
rect 14815 1760 14855 1765
rect 14815 1730 14820 1760
rect 14850 1730 14855 1760
rect 14815 1725 14855 1730
rect 15405 1760 15445 1765
rect 15405 1730 15410 1760
rect 15440 1730 15445 1760
rect 15405 1725 15445 1730
rect 15735 1760 15775 1765
rect 15735 1730 15740 1760
rect 15770 1730 15775 1760
rect 15735 1725 15775 1730
rect 14515 1705 14555 1710
rect 14515 1675 14520 1705
rect 14550 1675 14555 1705
rect 14515 1670 14555 1675
rect 14825 1650 14845 1725
rect 15415 1710 15435 1725
rect 14880 1705 14920 1710
rect 14880 1675 14885 1705
rect 14915 1675 14920 1705
rect 14880 1670 14920 1675
rect 15105 1705 15145 1710
rect 15105 1675 15110 1705
rect 15140 1675 15145 1705
rect 15105 1670 15145 1675
rect 15305 1705 15345 1710
rect 15305 1675 15310 1705
rect 15340 1675 15345 1705
rect 15305 1670 15345 1675
rect 15408 1700 15442 1710
rect 15408 1680 15416 1700
rect 15434 1680 15442 1700
rect 15408 1670 15442 1680
rect 15505 1705 15545 1710
rect 15505 1675 15510 1705
rect 15540 1675 15545 1705
rect 15505 1670 15545 1675
rect 14890 1650 14910 1670
rect 14820 1645 14855 1650
rect 14820 1605 14855 1610
rect 14880 1645 14915 1650
rect 14880 1605 14915 1610
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1565 4845 1595
rect 4805 1560 4845 1565
rect 5410 1595 5450 1600
rect 5410 1565 5415 1595
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1515 4305 1545
rect 4265 1510 4305 1515
rect 4385 1545 4425 1550
rect 4385 1515 4390 1545
rect 4420 1515 4425 1545
rect 4385 1510 4425 1515
rect 4505 1545 4545 1550
rect 4505 1515 4510 1545
rect 4540 1515 4545 1545
rect 4505 1510 4545 1515
rect 4625 1545 4665 1550
rect 4625 1515 4630 1545
rect 4660 1515 4665 1545
rect 4625 1510 4665 1515
rect 4745 1545 4785 1550
rect 4745 1515 4750 1545
rect 4780 1515 4785 1545
rect 4745 1510 4785 1515
rect 5135 1545 5175 1550
rect 5135 1515 5140 1545
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 4205 1500 4245 1505
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1470 4210 1500
rect 4240 1470 4245 1500
rect 4205 1465 4245 1470
rect 4325 1500 4365 1505
rect 4325 1470 4330 1500
rect 4360 1470 4365 1500
rect 4325 1465 4365 1470
rect 4445 1500 4485 1505
rect 4445 1470 4450 1500
rect 4480 1470 4485 1500
rect 4445 1465 4485 1470
rect 4685 1500 4725 1505
rect 4685 1470 4690 1500
rect 4720 1470 4725 1500
rect 4685 1465 4725 1470
rect 4805 1500 4845 1505
rect 4805 1470 4810 1500
rect 4840 1470 4845 1500
rect 4805 1465 4845 1470
rect 4925 1500 4965 1505
rect 4925 1470 4930 1500
rect 4960 1470 4965 1500
rect 4925 1465 4965 1470
rect 5045 1500 5085 1505
rect 5045 1470 5050 1500
rect 5080 1470 5085 1500
rect 5145 1490 5165 1510
rect 5045 1465 5085 1470
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 15745 1395 15765 1725
rect 15735 1390 15775 1395
rect 15735 1360 15740 1390
rect 15770 1360 15775 1390
rect 15735 1355 15775 1360
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1155 3415 1185
rect 3375 1150 3415 1155
rect 3985 1185 4025 1190
rect 3985 1155 3990 1185
rect 4020 1155 4025 1185
rect 3985 1150 4025 1155
rect 4595 1185 4635 1190
rect 4595 1155 4600 1185
rect 4630 1155 4635 1185
rect 4595 1150 4635 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1095 2985 1125
rect 2945 1090 2985 1095
rect 3025 1125 3065 1130
rect 3025 1095 3030 1125
rect 3060 1095 3065 1125
rect 3025 1090 3065 1095
rect 3105 1125 3145 1130
rect 3105 1095 3110 1125
rect 3140 1095 3145 1125
rect 3105 1090 3145 1095
rect 3185 1125 3225 1130
rect 3185 1095 3190 1125
rect 3220 1095 3225 1125
rect 3185 1090 3225 1095
rect 3265 1125 3305 1130
rect 3265 1095 3270 1125
rect 3300 1095 3305 1125
rect 3265 1090 3305 1095
rect 3345 1125 3385 1130
rect 3345 1095 3350 1125
rect 3380 1095 3385 1125
rect 3345 1090 3385 1095
rect 3425 1125 3465 1130
rect 3425 1095 3430 1125
rect 3460 1095 3465 1125
rect 3425 1090 3465 1095
rect 3505 1125 3545 1130
rect 3505 1095 3510 1125
rect 3540 1095 3545 1125
rect 3505 1090 3545 1095
rect 3585 1125 3625 1130
rect 3585 1095 3590 1125
rect 3620 1095 3625 1125
rect 3585 1090 3625 1095
rect 3665 1125 3705 1130
rect 3665 1095 3670 1125
rect 3700 1095 3705 1125
rect 3665 1090 3705 1095
rect 3745 1125 3785 1130
rect 3745 1095 3750 1125
rect 3780 1095 3785 1125
rect 3745 1090 3785 1095
rect 3825 1125 3865 1130
rect 3825 1095 3830 1125
rect 3860 1095 3865 1125
rect 3825 1090 3865 1095
rect 3905 1125 3945 1130
rect 3905 1095 3910 1125
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1095 4025 1125
rect 3985 1090 4025 1095
rect 4065 1125 4105 1130
rect 4065 1095 4070 1125
rect 4100 1095 4105 1125
rect 4065 1090 4105 1095
rect 4145 1125 4185 1130
rect 4145 1095 4150 1125
rect 4180 1095 4185 1125
rect 4145 1090 4185 1095
rect 4225 1125 4265 1130
rect 4225 1095 4230 1125
rect 4260 1095 4265 1125
rect 4225 1090 4265 1095
rect 4305 1125 4345 1130
rect 4305 1095 4310 1125
rect 4340 1095 4345 1125
rect 4305 1090 4345 1095
rect 4385 1125 4425 1130
rect 4385 1095 4390 1125
rect 4420 1095 4425 1125
rect 4385 1090 4425 1095
rect 4465 1125 4505 1130
rect 4465 1095 4470 1125
rect 4500 1095 4505 1125
rect 4465 1090 4505 1095
rect 4545 1125 4585 1130
rect 4545 1095 4550 1125
rect 4580 1095 4585 1125
rect 4545 1090 4585 1095
rect 4625 1125 4665 1130
rect 4625 1095 4630 1125
rect 4660 1095 4665 1125
rect 4625 1090 4665 1095
rect 4705 1125 4745 1130
rect 4705 1095 4710 1125
rect 4740 1095 4745 1125
rect 4705 1090 4745 1095
rect 4785 1125 4825 1130
rect 4785 1095 4790 1125
rect 4820 1095 4825 1125
rect 4785 1090 4825 1095
rect 4865 1125 4905 1130
rect 4865 1095 4870 1125
rect 4900 1095 4905 1125
rect 4865 1090 4905 1095
rect 4945 1125 4985 1130
rect 4945 1095 4950 1125
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1010 2660 1040
rect 2620 1005 2660 1010
rect 2905 1040 2945 1045
rect 2905 1010 2910 1040
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1010 5150 1040
rect 5110 1005 5150 1010
rect 15205 935 15245 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 900 3035 930
rect 2995 895 3035 900
rect 3175 930 3215 935
rect 3175 900 3180 930
rect 3210 900 3215 930
rect 3175 895 3215 900
rect 3355 930 3395 935
rect 3355 900 3360 930
rect 3390 900 3395 930
rect 3355 895 3395 900
rect 3535 930 3575 935
rect 3535 900 3540 930
rect 3570 900 3575 930
rect 3535 895 3575 900
rect 3715 930 3755 935
rect 3715 900 3720 930
rect 3750 900 3755 930
rect 3715 895 3755 900
rect 3895 930 3935 935
rect 3895 900 3900 930
rect 3930 900 3935 930
rect 3895 895 3935 900
rect 4075 930 4115 935
rect 4075 900 4080 930
rect 4110 900 4115 930
rect 4075 895 4115 900
rect 4255 930 4295 935
rect 4255 900 4260 930
rect 4290 900 4295 930
rect 4255 895 4295 900
rect 4435 930 4475 935
rect 4435 900 4440 930
rect 4470 900 4475 930
rect 4435 895 4475 900
rect 4615 930 4655 935
rect 4615 900 4620 930
rect 4650 900 4655 930
rect 4615 895 4655 900
rect 4795 930 4835 935
rect 4795 900 4800 930
rect 4830 900 4835 930
rect 4795 895 4835 900
rect 4975 930 5015 935
rect 4975 900 4980 930
rect 5010 900 5015 930
rect 15205 905 15210 935
rect 15240 905 15245 935
rect 15205 900 15245 905
rect 15405 935 15445 940
rect 15405 905 15410 935
rect 15440 905 15445 935
rect 15405 900 15445 905
rect 4975 895 5015 900
rect 15810 805 15830 2145
rect 16010 1900 16030 2290
rect 16330 2240 16350 2340
rect 17330 2285 17350 2340
rect 17870 2330 17890 3815
rect 17960 3680 18000 3685
rect 17960 3650 17965 3680
rect 17995 3650 18000 3680
rect 17960 3645 18000 3650
rect 17905 3635 17945 3640
rect 17905 3605 17910 3635
rect 17940 3605 17945 3635
rect 17905 3600 17945 3605
rect 17860 2325 17900 2330
rect 17860 2295 17865 2325
rect 17895 2295 17900 2325
rect 17860 2290 17900 2295
rect 16440 2280 16480 2285
rect 16440 2250 16445 2280
rect 16475 2250 16480 2280
rect 16440 2245 16480 2250
rect 16660 2280 16700 2285
rect 16660 2250 16665 2280
rect 16695 2250 16700 2280
rect 16660 2245 16700 2250
rect 16880 2280 16920 2285
rect 16880 2250 16885 2280
rect 16915 2250 16920 2280
rect 16880 2245 16920 2250
rect 17100 2280 17140 2285
rect 17100 2250 17105 2280
rect 17135 2250 17140 2280
rect 17100 2245 17140 2250
rect 17320 2280 17360 2285
rect 17320 2250 17325 2280
rect 17355 2250 17360 2280
rect 17320 2245 17360 2250
rect 16330 2235 16370 2240
rect 16330 2205 16335 2235
rect 16365 2205 16370 2235
rect 16330 2200 16370 2205
rect 16340 2185 16360 2200
rect 16450 2185 16470 2245
rect 16550 2235 16590 2240
rect 16550 2205 16555 2235
rect 16585 2205 16590 2235
rect 16550 2200 16590 2205
rect 16560 2185 16580 2200
rect 16670 2185 16690 2245
rect 16770 2235 16810 2240
rect 16770 2205 16775 2235
rect 16805 2205 16810 2235
rect 16770 2200 16810 2205
rect 16780 2185 16800 2200
rect 16890 2185 16910 2245
rect 16990 2235 17030 2240
rect 16990 2205 16995 2235
rect 17025 2205 17030 2235
rect 16990 2200 17030 2205
rect 17000 2185 17020 2200
rect 17110 2185 17130 2245
rect 17210 2235 17250 2240
rect 17210 2205 17215 2235
rect 17245 2205 17250 2235
rect 17210 2200 17250 2205
rect 17220 2185 17240 2200
rect 17330 2185 17350 2245
rect 17430 2235 17470 2240
rect 17430 2205 17435 2235
rect 17465 2205 17470 2235
rect 17430 2200 17470 2205
rect 17440 2185 17460 2200
rect 16330 2175 16370 2185
rect 16330 2155 16340 2175
rect 16360 2155 16370 2175
rect 16330 2145 16370 2155
rect 16440 2175 16480 2185
rect 16440 2155 16450 2175
rect 16470 2155 16480 2175
rect 16440 2145 16480 2155
rect 16550 2175 16590 2185
rect 16550 2155 16560 2175
rect 16580 2155 16590 2175
rect 16550 2145 16590 2155
rect 16660 2175 16700 2185
rect 16660 2155 16670 2175
rect 16690 2155 16700 2175
rect 16660 2145 16700 2155
rect 16770 2175 16810 2185
rect 16770 2155 16780 2175
rect 16800 2155 16810 2175
rect 16770 2145 16810 2155
rect 16828 2180 16862 2185
rect 16828 2150 16831 2180
rect 16859 2150 16862 2180
rect 16828 2145 16862 2150
rect 16880 2175 16920 2185
rect 16880 2155 16890 2175
rect 16910 2155 16920 2175
rect 16880 2145 16920 2155
rect 16990 2175 17030 2185
rect 16990 2155 17000 2175
rect 17020 2155 17030 2175
rect 16990 2145 17030 2155
rect 17100 2175 17140 2185
rect 17100 2155 17110 2175
rect 17130 2155 17140 2175
rect 17100 2145 17140 2155
rect 17210 2175 17250 2185
rect 17210 2155 17220 2175
rect 17240 2155 17250 2175
rect 17210 2145 17250 2155
rect 17320 2175 17360 2185
rect 17320 2155 17330 2175
rect 17350 2155 17360 2175
rect 17320 2145 17360 2155
rect 17430 2175 17470 2185
rect 17430 2155 17440 2175
rect 17460 2155 17470 2175
rect 17430 2145 17470 2155
rect 16385 1960 16425 1965
rect 16385 1930 16390 1960
rect 16420 1930 16425 1960
rect 16385 1925 16425 1930
rect 16495 1955 16535 1965
rect 16495 1935 16505 1955
rect 16525 1935 16535 1955
rect 16495 1925 16535 1935
rect 16605 1960 16645 1965
rect 16605 1930 16610 1960
rect 16640 1930 16645 1960
rect 16605 1925 16645 1930
rect 16715 1955 16755 1965
rect 16715 1935 16725 1955
rect 16745 1935 16755 1955
rect 16715 1925 16755 1935
rect 16825 1960 16865 1965
rect 16825 1930 16830 1960
rect 16860 1930 16865 1960
rect 16825 1925 16865 1930
rect 16935 1955 16975 1965
rect 16935 1935 16945 1955
rect 16965 1935 16975 1955
rect 16935 1925 16975 1935
rect 17045 1960 17085 1965
rect 17045 1930 17050 1960
rect 17080 1930 17085 1960
rect 17045 1925 17085 1930
rect 17155 1955 17195 1965
rect 17155 1935 17165 1955
rect 17185 1935 17195 1955
rect 17155 1925 17195 1935
rect 17245 1960 17305 1965
rect 17245 1930 17270 1960
rect 17300 1930 17305 1960
rect 17245 1925 17305 1930
rect 17375 1955 17415 1965
rect 17375 1935 17385 1955
rect 17405 1935 17415 1955
rect 17375 1925 17415 1935
rect 16505 1910 16525 1925
rect 16725 1910 16745 1925
rect 16945 1910 16965 1925
rect 17165 1910 17185 1925
rect 16495 1905 16555 1910
rect 16000 1895 16040 1900
rect 16000 1865 16005 1895
rect 16035 1865 16040 1895
rect 16495 1875 16500 1905
rect 16530 1875 16555 1905
rect 16495 1870 16555 1875
rect 16715 1905 16755 1910
rect 16715 1875 16720 1905
rect 16750 1875 16755 1905
rect 16715 1870 16755 1875
rect 16935 1905 16975 1910
rect 16935 1875 16940 1905
rect 16970 1875 16975 1905
rect 16935 1870 16975 1875
rect 17155 1905 17195 1910
rect 17155 1875 17160 1905
rect 17190 1875 17195 1905
rect 17155 1870 17195 1875
rect 16000 1860 16040 1865
rect 16190 1850 16230 1855
rect 16190 1820 16195 1850
rect 16225 1820 16230 1850
rect 16190 1815 16230 1820
rect 16410 1850 16450 1855
rect 16410 1820 16415 1850
rect 16445 1820 16450 1850
rect 16410 1815 16450 1820
rect 16200 1780 16220 1815
rect 16420 1780 16440 1815
rect 16190 1770 16230 1780
rect 16085 1760 16125 1765
rect 16085 1730 16090 1760
rect 16120 1730 16125 1760
rect 16190 1750 16200 1770
rect 16220 1750 16230 1770
rect 16410 1770 16450 1780
rect 16190 1740 16230 1750
rect 16305 1760 16345 1765
rect 16085 1725 16125 1730
rect 16305 1730 16310 1760
rect 16340 1730 16345 1760
rect 16410 1750 16420 1770
rect 16440 1750 16450 1770
rect 16535 1765 16555 1870
rect 17245 1855 17265 1925
rect 17385 1910 17405 1925
rect 17375 1905 17415 1910
rect 17375 1875 17380 1905
rect 17410 1875 17415 1905
rect 17870 1900 17890 2290
rect 17375 1870 17415 1875
rect 17860 1895 17900 1900
rect 17860 1865 17865 1895
rect 17895 1865 17900 1895
rect 17860 1860 17900 1865
rect 16640 1850 16680 1855
rect 16640 1820 16645 1850
rect 16675 1820 16680 1850
rect 16640 1815 16680 1820
rect 17230 1850 17270 1855
rect 17230 1820 17235 1850
rect 17265 1820 17270 1850
rect 17230 1815 17270 1820
rect 17450 1850 17490 1855
rect 17450 1820 17455 1850
rect 17485 1820 17490 1850
rect 17450 1815 17490 1820
rect 17680 1850 17720 1855
rect 17680 1820 17685 1850
rect 17715 1820 17720 1850
rect 17680 1815 17720 1820
rect 16650 1780 16670 1815
rect 16820 1805 16860 1810
rect 16640 1770 16680 1780
rect 16820 1775 16825 1805
rect 16855 1775 16860 1805
rect 16820 1770 16860 1775
rect 16940 1805 16980 1810
rect 16940 1775 16945 1805
rect 16975 1775 16980 1805
rect 17240 1780 17260 1815
rect 17460 1780 17480 1815
rect 17690 1780 17710 1815
rect 16940 1770 16980 1775
rect 17230 1770 17270 1780
rect 16410 1740 16450 1750
rect 16525 1760 16565 1765
rect 16305 1725 16345 1730
rect 16525 1730 16530 1760
rect 16560 1730 16565 1760
rect 16640 1750 16650 1770
rect 16670 1750 16680 1770
rect 16640 1740 16680 1750
rect 16525 1725 16565 1730
rect 16830 1720 16850 1770
rect 16950 1720 16970 1770
rect 17125 1760 17165 1765
rect 17125 1730 17130 1760
rect 17160 1730 17165 1760
rect 17230 1750 17240 1770
rect 17260 1750 17270 1770
rect 17450 1770 17490 1780
rect 17230 1740 17270 1750
rect 17345 1760 17385 1765
rect 17125 1725 17165 1730
rect 17345 1730 17350 1760
rect 17380 1730 17385 1760
rect 17450 1750 17460 1770
rect 17480 1750 17490 1770
rect 17680 1770 17720 1780
rect 17450 1740 17490 1750
rect 17565 1760 17605 1765
rect 17345 1725 17385 1730
rect 17565 1730 17570 1760
rect 17600 1730 17605 1760
rect 17680 1750 17690 1770
rect 17710 1750 17720 1770
rect 17680 1740 17720 1750
rect 17565 1725 17605 1730
rect 16237 1715 16269 1720
rect 16237 1685 16240 1715
rect 16266 1685 16269 1715
rect 16237 1680 16269 1685
rect 16457 1715 16489 1720
rect 16457 1685 16460 1715
rect 16486 1685 16489 1715
rect 16457 1680 16489 1685
rect 16601 1715 16633 1720
rect 16601 1685 16604 1715
rect 16630 1685 16633 1715
rect 16601 1680 16633 1685
rect 16820 1710 16850 1720
rect 16820 1690 16825 1710
rect 16845 1690 16850 1710
rect 16820 1680 16850 1690
rect 16867 1715 16899 1720
rect 16867 1685 16870 1715
rect 16896 1685 16899 1715
rect 16867 1680 16899 1685
rect 16950 1710 16980 1720
rect 16950 1690 16955 1710
rect 16975 1690 16980 1710
rect 16950 1680 16980 1690
rect 17277 1715 17309 1720
rect 17277 1685 17280 1715
rect 17306 1685 17309 1715
rect 17277 1680 17309 1685
rect 17497 1715 17529 1720
rect 17497 1685 17500 1715
rect 17526 1685 17529 1715
rect 17497 1680 17529 1685
rect 17641 1715 17673 1720
rect 17641 1685 17644 1715
rect 17670 1685 17673 1715
rect 17641 1680 17673 1685
rect 16106 1495 16138 1500
rect 16106 1465 16109 1495
rect 16135 1465 16138 1495
rect 16106 1460 16138 1465
rect 16305 1495 16345 1500
rect 16305 1465 16310 1495
rect 16340 1465 16345 1495
rect 16305 1460 16345 1465
rect 16525 1495 16565 1500
rect 16525 1465 16530 1495
rect 16560 1465 16565 1495
rect 16525 1460 16565 1465
rect 16825 1490 16855 1500
rect 16825 1470 16830 1490
rect 16850 1470 16855 1490
rect 16825 1460 16855 1470
rect 16875 1490 16905 1500
rect 16875 1470 16880 1490
rect 16900 1470 16905 1490
rect 16875 1460 16905 1470
rect 16922 1495 16954 1500
rect 16922 1465 16925 1495
rect 16951 1465 16954 1495
rect 16922 1460 16954 1465
rect 17146 1495 17178 1500
rect 17146 1465 17149 1495
rect 17175 1465 17178 1495
rect 17146 1460 17178 1465
rect 17345 1495 17385 1500
rect 17345 1465 17350 1495
rect 17380 1465 17385 1495
rect 17345 1460 17385 1465
rect 17565 1495 17605 1500
rect 17565 1465 17570 1495
rect 17600 1465 17605 1495
rect 17565 1460 17605 1465
rect 16145 1435 16185 1440
rect 16145 1405 16150 1435
rect 16180 1405 16185 1435
rect 16145 1400 16185 1405
rect 16250 1435 16290 1440
rect 16250 1405 16255 1435
rect 16285 1405 16290 1435
rect 16250 1400 16290 1405
rect 16360 1435 16400 1440
rect 16360 1405 16365 1435
rect 16395 1405 16400 1435
rect 16360 1400 16400 1405
rect 16470 1435 16510 1440
rect 16470 1405 16475 1435
rect 16505 1405 16510 1435
rect 16470 1400 16510 1405
rect 16580 1435 16620 1440
rect 16580 1405 16585 1435
rect 16615 1405 16620 1435
rect 16580 1400 16620 1405
rect 16830 1350 16850 1460
rect 16005 1345 16045 1350
rect 16005 1315 16010 1345
rect 16040 1315 16045 1345
rect 16005 1310 16045 1315
rect 16810 1345 16850 1350
rect 16810 1315 16815 1345
rect 16845 1315 16850 1345
rect 16810 1310 16850 1315
rect 16015 860 16035 1310
rect 16315 1295 16355 1300
rect 16315 1265 16320 1295
rect 16350 1265 16355 1295
rect 16315 1260 16355 1265
rect 16325 1240 16345 1260
rect 16820 1240 16840 1310
rect 16880 1300 16900 1460
rect 17185 1435 17225 1440
rect 17185 1405 17190 1435
rect 17220 1405 17225 1435
rect 17185 1400 17225 1405
rect 17290 1435 17330 1440
rect 17290 1405 17295 1435
rect 17325 1405 17330 1435
rect 17290 1400 17330 1405
rect 17400 1435 17440 1440
rect 17400 1405 17405 1435
rect 17435 1405 17440 1435
rect 17400 1400 17440 1405
rect 17510 1435 17550 1440
rect 17510 1405 17515 1435
rect 17545 1405 17550 1435
rect 17510 1400 17550 1405
rect 17620 1435 17660 1440
rect 17620 1405 17625 1435
rect 17655 1405 17660 1435
rect 17620 1400 17660 1405
rect 16880 1295 16920 1300
rect 16880 1265 16885 1295
rect 16915 1265 16920 1295
rect 16880 1260 16920 1265
rect 17915 1255 17935 3600
rect 17595 1250 17635 1255
rect 16315 1230 16355 1240
rect 16315 1210 16325 1230
rect 16345 1210 16355 1230
rect 16315 1200 16355 1210
rect 16425 1235 16465 1240
rect 16425 1205 16430 1235
rect 16460 1205 16465 1235
rect 16425 1200 16465 1205
rect 16535 1235 16575 1240
rect 16535 1205 16540 1235
rect 16570 1205 16575 1235
rect 16535 1200 16575 1205
rect 16645 1235 16685 1240
rect 16645 1205 16650 1235
rect 16680 1205 16685 1235
rect 16645 1200 16685 1205
rect 16755 1235 16795 1240
rect 16755 1205 16760 1235
rect 16790 1205 16795 1235
rect 16755 1200 16795 1205
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 16815 1200 16845 1210
rect 16865 1235 16905 1240
rect 16865 1205 16870 1235
rect 16900 1205 16905 1235
rect 16865 1200 16905 1205
rect 16975 1235 17015 1240
rect 16975 1205 16980 1235
rect 17010 1205 17015 1235
rect 16975 1200 17015 1205
rect 17085 1235 17125 1240
rect 17085 1205 17090 1235
rect 17120 1205 17125 1235
rect 17085 1200 17125 1205
rect 17195 1235 17235 1240
rect 17195 1205 17200 1235
rect 17230 1205 17235 1235
rect 17195 1200 17235 1205
rect 17305 1235 17345 1240
rect 17305 1205 17310 1235
rect 17340 1205 17345 1235
rect 17305 1200 17345 1205
rect 17415 1235 17455 1240
rect 17415 1205 17420 1235
rect 17450 1205 17455 1235
rect 17415 1200 17455 1205
rect 17525 1235 17565 1240
rect 17525 1205 17530 1235
rect 17560 1205 17565 1235
rect 17595 1220 17600 1250
rect 17630 1220 17635 1250
rect 17595 1215 17635 1220
rect 17905 1250 17945 1255
rect 17905 1220 17910 1250
rect 17940 1220 17945 1250
rect 17905 1215 17945 1220
rect 17525 1200 17565 1205
rect 16165 915 16205 920
rect 16165 885 16170 915
rect 16200 885 16205 915
rect 16165 880 16205 885
rect 16260 915 16300 920
rect 16260 885 16265 915
rect 16295 885 16300 915
rect 16260 880 16300 885
rect 16370 915 16410 920
rect 16370 885 16375 915
rect 16405 885 16410 915
rect 16370 880 16410 885
rect 16480 915 16520 920
rect 16480 885 16485 915
rect 16515 885 16520 915
rect 16480 880 16520 885
rect 16590 915 16630 920
rect 16590 885 16595 915
rect 16625 885 16630 915
rect 16590 880 16630 885
rect 16700 915 16740 920
rect 16700 885 16705 915
rect 16735 885 16740 915
rect 16700 880 16740 885
rect 16810 915 16850 920
rect 16810 885 16815 915
rect 16845 885 16850 915
rect 16810 880 16850 885
rect 16920 915 16960 920
rect 16920 885 16925 915
rect 16955 885 16960 915
rect 16920 880 16960 885
rect 17030 915 17070 920
rect 17030 885 17035 915
rect 17065 885 17070 915
rect 17030 880 17070 885
rect 17140 915 17180 920
rect 17140 885 17145 915
rect 17175 885 17180 915
rect 17140 880 17180 885
rect 17250 915 17290 920
rect 17250 885 17255 915
rect 17285 885 17290 915
rect 17250 880 17290 885
rect 17360 915 17400 920
rect 17360 885 17365 915
rect 17395 885 17400 915
rect 17360 880 17400 885
rect 17470 915 17510 920
rect 17470 885 17475 915
rect 17505 885 17510 915
rect 17470 880 17510 885
rect 17620 915 17660 920
rect 17620 885 17625 915
rect 17655 885 17660 915
rect 17620 880 17660 885
rect 16935 860 16975 865
rect 16005 855 16045 860
rect 16005 825 16010 855
rect 16040 825 16045 855
rect 16005 820 16045 825
rect 16495 855 16535 860
rect 16495 825 16500 855
rect 16530 825 16535 855
rect 16935 830 16940 860
rect 16970 830 16975 860
rect 16935 825 16975 830
rect 17155 860 17195 865
rect 17155 830 17160 860
rect 17190 830 17195 860
rect 17155 825 17195 830
rect 17375 860 17415 865
rect 17375 830 17380 860
rect 17410 830 17415 860
rect 17375 825 17415 830
rect 16495 820 16535 825
rect 16945 805 16965 825
rect 17165 805 17185 825
rect 17385 805 17405 825
rect 17915 805 17935 1215
rect 17970 865 17990 3645
rect 18200 3635 18240 3640
rect 18200 3605 18205 3635
rect 18235 3605 18240 3635
rect 18200 3600 18240 3605
rect 18310 3635 18350 3640
rect 18310 3605 18315 3635
rect 18345 3605 18350 3635
rect 18310 3600 18350 3605
rect 18420 3635 18460 3640
rect 18420 3605 18425 3635
rect 18455 3605 18460 3635
rect 18420 3600 18460 3605
rect 18530 3635 18570 3640
rect 18530 3605 18535 3635
rect 18565 3605 18570 3635
rect 18530 3600 18570 3605
rect 18640 3635 18680 3640
rect 18640 3605 18645 3635
rect 18675 3605 18680 3635
rect 18640 3600 18680 3605
rect 18750 3635 18790 3640
rect 18750 3605 18755 3635
rect 18785 3605 18790 3635
rect 18750 3600 18790 3605
rect 19155 3635 19195 3640
rect 19155 3605 19160 3635
rect 19190 3605 19195 3635
rect 19155 3600 19195 3605
rect 24605 3635 24645 3640
rect 24605 3605 24610 3635
rect 24640 3605 24645 3635
rect 24605 3600 24645 3605
rect 25060 3635 25100 3640
rect 25060 3605 25065 3635
rect 25095 3605 25100 3635
rect 25060 3600 25100 3605
rect 25170 3635 25210 3640
rect 25170 3605 25175 3635
rect 25205 3605 25210 3635
rect 25170 3600 25210 3605
rect 25280 3635 25320 3640
rect 25280 3605 25285 3635
rect 25315 3605 25320 3635
rect 25280 3600 25320 3605
rect 25390 3635 25430 3640
rect 25390 3605 25395 3635
rect 25425 3605 25430 3635
rect 25390 3600 25430 3605
rect 25500 3635 25540 3640
rect 25500 3605 25505 3635
rect 25535 3605 25540 3635
rect 25500 3600 25540 3605
rect 25610 3635 25650 3640
rect 25610 3605 25615 3635
rect 25645 3605 25650 3635
rect 25610 3600 25650 3605
rect 19165 3560 19185 3600
rect 24615 3560 24635 3600
rect 19105 3555 19246 3560
rect 19105 3525 19110 3555
rect 19140 3525 19160 3555
rect 19190 3525 19210 3555
rect 19240 3525 19246 3555
rect 19105 3520 19246 3525
rect 24554 3555 24695 3560
rect 24554 3525 24560 3555
rect 24590 3525 24610 3555
rect 24640 3525 24660 3555
rect 24690 3525 24695 3555
rect 24554 3520 24695 3525
rect 26060 3190 26080 4735
rect 26355 4590 26375 4740
rect 26685 4735 26725 4740
rect 27295 4770 27335 4775
rect 27295 4740 27300 4770
rect 27330 4740 27335 4770
rect 27295 4735 27335 4740
rect 27358 4765 27392 4775
rect 27358 4745 27366 4765
rect 27384 4745 27392 4765
rect 27358 4735 27392 4745
rect 27415 4770 27455 4775
rect 27415 4740 27420 4770
rect 27450 4740 27455 4770
rect 27415 4735 27455 4740
rect 27535 4770 27575 4775
rect 27535 4740 27540 4770
rect 27570 4740 27575 4770
rect 27535 4735 27575 4740
rect 27655 4770 27695 4775
rect 27655 4740 27660 4770
rect 27690 4740 27695 4770
rect 27655 4735 27695 4740
rect 27365 4590 27385 4735
rect 26105 4585 26145 4590
rect 26105 4555 26110 4585
rect 26140 4555 26145 4585
rect 26105 4550 26145 4555
rect 26345 4585 26385 4590
rect 26345 4555 26350 4585
rect 26380 4555 26385 4585
rect 26345 4550 26385 4555
rect 27355 4585 27395 4590
rect 27355 4555 27360 4585
rect 27390 4555 27395 4585
rect 27355 4550 27395 4555
rect 26050 3185 26090 3190
rect 26050 3155 26055 3185
rect 26085 3155 26090 3185
rect 26050 3150 26090 3155
rect 18255 2965 18295 2970
rect 18255 2935 18260 2965
rect 18290 2935 18295 2965
rect 18255 2930 18295 2935
rect 18313 2960 18347 2970
rect 18313 2940 18321 2960
rect 18339 2940 18347 2960
rect 18313 2930 18347 2940
rect 18365 2965 18405 2970
rect 18365 2935 18370 2965
rect 18400 2935 18405 2965
rect 18365 2930 18405 2935
rect 18475 2965 18515 2970
rect 18475 2935 18480 2965
rect 18510 2935 18515 2965
rect 18475 2930 18515 2935
rect 18585 2965 18625 2970
rect 18585 2935 18590 2965
rect 18620 2935 18625 2965
rect 18585 2930 18625 2935
rect 18695 2965 18735 2970
rect 18695 2935 18700 2965
rect 18730 2935 18735 2965
rect 25115 2965 25155 2970
rect 18695 2930 18735 2935
rect 19105 2935 19246 2940
rect 18320 2885 18340 2930
rect 18015 2880 18055 2885
rect 18015 2850 18020 2880
rect 18050 2850 18055 2880
rect 18015 2845 18055 2850
rect 18310 2880 18350 2885
rect 18310 2850 18315 2880
rect 18345 2850 18350 2880
rect 18310 2845 18350 2850
rect 18025 2380 18045 2845
rect 18595 2830 18615 2930
rect 19105 2905 19110 2935
rect 19140 2905 19160 2935
rect 19190 2905 19210 2935
rect 19240 2905 19246 2935
rect 19105 2900 19246 2905
rect 24554 2935 24695 2940
rect 24554 2905 24560 2935
rect 24590 2905 24610 2935
rect 24640 2905 24660 2935
rect 24690 2905 24695 2935
rect 25115 2935 25120 2965
rect 25150 2935 25155 2965
rect 25115 2930 25155 2935
rect 25225 2965 25265 2970
rect 25225 2935 25230 2965
rect 25260 2935 25265 2965
rect 25225 2930 25265 2935
rect 25335 2965 25375 2970
rect 25335 2935 25340 2965
rect 25370 2935 25375 2965
rect 25335 2930 25375 2935
rect 25445 2965 25485 2970
rect 25445 2935 25450 2965
rect 25480 2935 25485 2965
rect 25445 2930 25485 2935
rect 25503 2960 25537 2970
rect 25503 2940 25511 2960
rect 25529 2940 25537 2960
rect 25503 2930 25537 2940
rect 25555 2965 25595 2970
rect 25555 2935 25560 2965
rect 25590 2935 25595 2965
rect 26115 2955 26135 4550
rect 26360 4480 26400 4485
rect 26360 4450 26365 4480
rect 26395 4450 26400 4480
rect 26360 4445 26400 4450
rect 26470 4480 26510 4485
rect 26470 4450 26475 4480
rect 26505 4450 26510 4480
rect 26470 4445 26510 4450
rect 26580 4480 26620 4485
rect 26580 4450 26585 4480
rect 26615 4450 26620 4480
rect 26580 4445 26620 4450
rect 26690 4480 26730 4485
rect 26690 4450 26695 4480
rect 26725 4450 26730 4480
rect 26690 4445 26730 4450
rect 26800 4480 26840 4485
rect 26800 4450 26805 4480
rect 26835 4450 26840 4480
rect 26800 4445 26840 4450
rect 26910 4480 26950 4485
rect 26910 4450 26915 4480
rect 26945 4450 26950 4480
rect 26910 4445 26950 4450
rect 27020 4480 27060 4485
rect 27020 4450 27025 4480
rect 27055 4450 27060 4480
rect 27020 4445 27060 4450
rect 27130 4480 27170 4485
rect 27130 4450 27135 4480
rect 27165 4450 27170 4480
rect 27130 4445 27170 4450
rect 27240 4480 27280 4485
rect 27240 4450 27245 4480
rect 27275 4450 27280 4480
rect 27240 4445 27280 4450
rect 27350 4480 27390 4485
rect 27350 4450 27355 4480
rect 27385 4450 27390 4480
rect 27350 4445 27390 4450
rect 26305 4360 26345 4365
rect 26305 4330 26310 4360
rect 26340 4330 26345 4360
rect 26305 4325 26345 4330
rect 26362 4355 26398 4365
rect 26362 4335 26370 4355
rect 26390 4335 26398 4355
rect 26362 4325 26398 4335
rect 26415 4355 26455 4365
rect 26415 4335 26425 4355
rect 26445 4335 26455 4355
rect 26415 4325 26455 4335
rect 26525 4360 26565 4365
rect 26525 4330 26530 4360
rect 26560 4330 26565 4360
rect 26525 4325 26565 4330
rect 26635 4355 26675 4365
rect 26635 4335 26645 4355
rect 26665 4335 26675 4355
rect 26635 4325 26675 4335
rect 26745 4360 26785 4365
rect 26745 4330 26750 4360
rect 26780 4330 26785 4360
rect 26745 4325 26785 4330
rect 26855 4355 26895 4365
rect 26855 4335 26865 4355
rect 26885 4335 26895 4355
rect 26855 4325 26895 4335
rect 26965 4360 27005 4365
rect 26965 4330 26970 4360
rect 27000 4330 27005 4360
rect 26965 4325 27005 4330
rect 27075 4355 27115 4365
rect 27075 4335 27085 4355
rect 27105 4335 27115 4355
rect 27075 4325 27115 4335
rect 27185 4360 27225 4365
rect 27185 4330 27190 4360
rect 27220 4330 27225 4360
rect 27185 4325 27225 4330
rect 27295 4355 27335 4365
rect 27295 4335 27305 4355
rect 27325 4335 27335 4355
rect 27295 4325 27335 4335
rect 27405 4360 27445 4365
rect 27405 4330 27410 4360
rect 27440 4330 27445 4360
rect 27405 4325 27445 4330
rect 26320 4130 26360 4135
rect 26320 4100 26325 4130
rect 26355 4100 26360 4130
rect 26320 4095 26360 4100
rect 26330 4075 26350 4095
rect 26375 4075 26395 4325
rect 26430 4250 26450 4325
rect 26645 4250 26665 4325
rect 26865 4250 26885 4325
rect 27085 4250 27105 4325
rect 27305 4250 27325 4325
rect 26420 4245 26460 4250
rect 26420 4215 26425 4245
rect 26455 4215 26460 4245
rect 26420 4210 26460 4215
rect 26635 4245 26675 4250
rect 26635 4215 26640 4245
rect 26670 4215 26675 4245
rect 26635 4210 26675 4215
rect 26855 4245 26895 4250
rect 26855 4215 26860 4245
rect 26890 4215 26895 4245
rect 26855 4210 26895 4215
rect 27075 4245 27115 4250
rect 27075 4215 27080 4245
rect 27110 4215 27115 4245
rect 27075 4210 27115 4215
rect 27295 4245 27335 4250
rect 27295 4215 27300 4245
rect 27330 4215 27335 4245
rect 27295 4210 27335 4215
rect 26430 4135 26450 4210
rect 27415 4200 27435 4325
rect 26420 4130 26460 4135
rect 26420 4100 26425 4130
rect 26455 4100 26460 4130
rect 26420 4095 26460 4100
rect 26530 4130 26570 4135
rect 26530 4100 26535 4130
rect 26565 4100 26570 4130
rect 26530 4095 26570 4100
rect 26640 4130 26680 4135
rect 26640 4100 26645 4130
rect 26675 4100 26680 4130
rect 26640 4095 26680 4100
rect 26750 4130 26790 4135
rect 26750 4100 26755 4130
rect 26785 4100 26790 4130
rect 26750 4095 26790 4100
rect 27050 4130 27090 4135
rect 27050 4100 27055 4130
rect 27085 4100 27090 4130
rect 27050 4095 27090 4100
rect 27150 4130 27190 4135
rect 27150 4100 27155 4130
rect 27185 4100 27190 4130
rect 27150 4095 27190 4100
rect 27260 4130 27300 4135
rect 27260 4100 27265 4130
rect 27295 4100 27300 4130
rect 27260 4095 27300 4100
rect 27370 4130 27410 4135
rect 27370 4100 27375 4130
rect 27405 4100 27410 4130
rect 27370 4095 27410 4100
rect 27480 4130 27520 4135
rect 27480 4100 27485 4130
rect 27515 4100 27520 4130
rect 27480 4095 27520 4100
rect 26430 4075 26450 4095
rect 26540 4075 26560 4095
rect 26650 4075 26670 4095
rect 26760 4075 26780 4095
rect 27060 4075 27080 4095
rect 27160 4075 27180 4095
rect 27270 4075 27290 4095
rect 27380 4075 27400 4095
rect 27490 4075 27510 4095
rect 26280 4069 26310 4075
rect 26280 4041 26282 4069
rect 26308 4041 26310 4069
rect 26280 4035 26310 4041
rect 26327 4065 26353 4075
rect 26327 4045 26330 4065
rect 26350 4045 26353 4065
rect 26327 4035 26353 4045
rect 26370 4065 26400 4075
rect 26370 4045 26375 4065
rect 26395 4045 26400 4065
rect 26370 4035 26400 4045
rect 26427 4065 26453 4075
rect 26427 4045 26430 4065
rect 26450 4045 26453 4065
rect 26427 4035 26453 4045
rect 26480 4069 26510 4075
rect 26480 4041 26482 4069
rect 26508 4041 26510 4069
rect 26480 4035 26510 4041
rect 26537 4065 26563 4075
rect 26537 4045 26540 4065
rect 26560 4045 26563 4065
rect 26537 4035 26563 4045
rect 26647 4065 26673 4075
rect 26647 4045 26650 4065
rect 26670 4045 26673 4065
rect 26647 4035 26673 4045
rect 26757 4065 26783 4075
rect 26757 4045 26760 4065
rect 26780 4045 26783 4065
rect 26757 4035 26783 4045
rect 27008 4069 27038 4075
rect 27008 4041 27010 4069
rect 27036 4041 27038 4069
rect 27008 4035 27038 4041
rect 27057 4065 27083 4075
rect 27057 4045 27060 4065
rect 27080 4045 27083 4065
rect 27057 4035 27083 4045
rect 27157 4065 27183 4075
rect 27157 4045 27160 4065
rect 27180 4045 27183 4065
rect 27157 4035 27183 4045
rect 27205 4070 27245 4075
rect 27205 4040 27210 4070
rect 27240 4040 27245 4070
rect 27205 4035 27245 4040
rect 27267 4065 27293 4075
rect 27267 4045 27270 4065
rect 27290 4045 27293 4065
rect 27267 4035 27293 4045
rect 27377 4065 27403 4075
rect 27377 4045 27380 4065
rect 27400 4045 27403 4065
rect 27377 4035 27403 4045
rect 27425 4070 27465 4075
rect 27425 4040 27430 4070
rect 27460 4040 27465 4070
rect 27425 4035 27465 4040
rect 27487 4065 27513 4075
rect 27487 4045 27490 4065
rect 27510 4045 27513 4065
rect 27487 4035 27513 4045
rect 27870 4070 27910 4075
rect 27870 4040 27875 4070
rect 27905 4040 27910 4070
rect 27870 4035 27910 4040
rect 26255 3945 26295 3955
rect 26255 3925 26265 3945
rect 26285 3925 26295 3945
rect 26255 3915 26295 3925
rect 26350 3945 26390 3955
rect 26350 3925 26360 3945
rect 26380 3925 26390 3945
rect 26350 3915 26390 3925
rect 26407 3950 26439 3955
rect 26407 3920 26410 3950
rect 26436 3920 26439 3950
rect 26407 3915 26439 3920
rect 26475 3945 26515 3955
rect 26475 3925 26485 3945
rect 26505 3925 26515 3945
rect 26475 3915 26515 3925
rect 26570 3945 26610 3955
rect 26570 3925 26580 3945
rect 26600 3925 26610 3945
rect 26570 3915 26610 3925
rect 26627 3950 26659 3955
rect 26627 3920 26630 3950
rect 26656 3920 26659 3950
rect 26627 3915 26659 3920
rect 26695 3945 26735 3955
rect 26695 3925 26705 3945
rect 26725 3925 26735 3945
rect 26695 3915 26735 3925
rect 26771 3950 26803 3955
rect 26771 3920 26774 3950
rect 26800 3920 26803 3950
rect 26771 3915 26803 3920
rect 26820 3945 26860 3955
rect 26820 3925 26830 3945
rect 26850 3925 26860 3945
rect 26820 3915 26860 3925
rect 26985 3945 27025 3955
rect 26985 3925 26995 3945
rect 27015 3925 27025 3945
rect 26985 3915 27025 3925
rect 27080 3945 27120 3955
rect 27080 3925 27090 3945
rect 27110 3925 27120 3945
rect 27080 3915 27120 3925
rect 27137 3950 27169 3955
rect 27137 3920 27140 3950
rect 27166 3920 27169 3950
rect 27137 3915 27169 3920
rect 27205 3945 27245 3955
rect 27205 3925 27215 3945
rect 27235 3925 27245 3945
rect 27205 3915 27245 3925
rect 27300 3945 27340 3955
rect 27300 3925 27310 3945
rect 27330 3925 27340 3945
rect 27300 3915 27340 3925
rect 27357 3950 27389 3955
rect 27357 3920 27360 3950
rect 27386 3920 27389 3950
rect 27357 3915 27389 3920
rect 27425 3945 27465 3955
rect 27425 3925 27435 3945
rect 27455 3925 27465 3945
rect 27425 3915 27465 3925
rect 27501 3950 27533 3955
rect 27501 3920 27504 3950
rect 27530 3920 27533 3950
rect 27501 3915 27533 3920
rect 27550 3945 27590 3955
rect 27550 3925 27560 3945
rect 27580 3925 27590 3945
rect 27550 3915 27590 3925
rect 26265 3895 26285 3915
rect 26370 3895 26390 3915
rect 26485 3895 26505 3915
rect 26590 3895 26610 3915
rect 26705 3895 26725 3915
rect 26820 3895 26840 3915
rect 26995 3895 27015 3915
rect 26255 3890 26295 3895
rect 26255 3860 26260 3890
rect 26290 3860 26295 3890
rect 26255 3855 26295 3860
rect 26360 3890 26400 3895
rect 26360 3860 26365 3890
rect 26395 3860 26400 3890
rect 26360 3855 26400 3860
rect 26475 3890 26515 3895
rect 26475 3860 26480 3890
rect 26510 3860 26515 3890
rect 26475 3855 26515 3860
rect 26580 3890 26620 3895
rect 26580 3860 26585 3890
rect 26615 3860 26620 3890
rect 26580 3855 26620 3860
rect 26695 3890 26735 3895
rect 26695 3860 26700 3890
rect 26730 3860 26735 3890
rect 26695 3855 26735 3860
rect 26810 3890 26850 3895
rect 26810 3860 26815 3890
rect 26845 3860 26850 3890
rect 26810 3855 26850 3860
rect 26985 3890 27025 3895
rect 26985 3860 26990 3890
rect 27020 3860 27025 3890
rect 26985 3855 27025 3860
rect 27100 3785 27120 3915
rect 27215 3895 27235 3915
rect 27205 3890 27245 3895
rect 27205 3860 27210 3890
rect 27240 3860 27245 3890
rect 27205 3855 27245 3860
rect 27320 3785 27340 3915
rect 27435 3895 27455 3915
rect 27425 3890 27465 3895
rect 27425 3860 27430 3890
rect 27460 3860 27465 3890
rect 27425 3855 27465 3860
rect 27550 3785 27570 3915
rect 27090 3780 27130 3785
rect 27090 3750 27095 3780
rect 27125 3750 27130 3780
rect 27090 3745 27130 3750
rect 27310 3780 27350 3785
rect 27310 3750 27315 3780
rect 27345 3750 27350 3780
rect 27310 3745 27350 3750
rect 27540 3780 27580 3785
rect 27540 3750 27545 3780
rect 27575 3750 27580 3780
rect 27540 3745 27580 3750
rect 26340 3655 26380 3660
rect 26340 3625 26345 3655
rect 26375 3625 26380 3655
rect 26340 3620 26380 3625
rect 26460 3655 26500 3660
rect 26460 3625 26465 3655
rect 26495 3625 26500 3655
rect 26460 3620 26500 3625
rect 26580 3655 26620 3660
rect 26580 3625 26585 3655
rect 26615 3625 26620 3655
rect 26580 3620 26620 3625
rect 26700 3655 26740 3660
rect 26700 3625 26705 3655
rect 26735 3625 26740 3655
rect 26700 3620 26740 3625
rect 26820 3655 26860 3660
rect 26820 3625 26825 3655
rect 26855 3625 26860 3655
rect 26820 3620 26860 3625
rect 26940 3655 26980 3660
rect 26940 3625 26945 3655
rect 26975 3625 26980 3655
rect 26940 3620 26980 3625
rect 27060 3655 27100 3660
rect 27060 3625 27065 3655
rect 27095 3625 27100 3655
rect 27060 3620 27100 3625
rect 27180 3655 27220 3660
rect 27180 3625 27185 3655
rect 27215 3625 27220 3655
rect 27180 3620 27220 3625
rect 27300 3655 27340 3660
rect 27300 3625 27305 3655
rect 27335 3625 27340 3655
rect 27300 3620 27340 3625
rect 27420 3655 27460 3660
rect 27420 3625 27425 3655
rect 27455 3625 27460 3655
rect 27420 3620 27460 3625
rect 26280 3180 26320 3190
rect 26280 3160 26290 3180
rect 26310 3160 26320 3180
rect 26280 3150 26320 3160
rect 26400 3180 26440 3190
rect 26400 3160 26410 3180
rect 26430 3160 26440 3180
rect 26400 3150 26440 3160
rect 26520 3180 26560 3190
rect 26520 3160 26530 3180
rect 26550 3160 26560 3180
rect 26520 3150 26560 3160
rect 26640 3180 26680 3190
rect 26640 3160 26650 3180
rect 26670 3160 26680 3180
rect 26640 3150 26680 3160
rect 26760 3180 26800 3190
rect 26760 3160 26770 3180
rect 26790 3160 26800 3180
rect 26760 3150 26800 3160
rect 26823 3185 26857 3190
rect 26823 3155 26826 3185
rect 26854 3155 26857 3185
rect 26823 3150 26857 3155
rect 26880 3180 26920 3190
rect 26880 3160 26890 3180
rect 26910 3160 26920 3180
rect 26880 3150 26920 3160
rect 27000 3180 27040 3190
rect 27000 3160 27010 3180
rect 27030 3160 27040 3180
rect 27000 3150 27040 3160
rect 27120 3180 27160 3190
rect 27120 3160 27130 3180
rect 27150 3160 27160 3180
rect 27120 3150 27160 3160
rect 27240 3180 27280 3190
rect 27240 3160 27250 3180
rect 27270 3160 27280 3180
rect 27240 3150 27280 3160
rect 27360 3180 27400 3190
rect 27360 3160 27370 3180
rect 27390 3160 27400 3180
rect 27360 3150 27400 3160
rect 27480 3180 27520 3190
rect 27480 3160 27490 3180
rect 27510 3160 27520 3180
rect 27480 3150 27520 3160
rect 26290 3135 26310 3150
rect 26280 3130 26320 3135
rect 26280 3100 26285 3130
rect 26315 3100 26320 3130
rect 26280 3095 26320 3100
rect 26410 3010 26430 3150
rect 26530 3135 26550 3150
rect 26520 3130 26560 3135
rect 26520 3100 26525 3130
rect 26555 3100 26560 3130
rect 26520 3095 26560 3100
rect 26650 3010 26670 3150
rect 26770 3135 26790 3150
rect 26760 3130 26800 3135
rect 26760 3100 26765 3130
rect 26795 3100 26800 3130
rect 26760 3095 26800 3100
rect 26890 3010 26910 3150
rect 27010 3135 27030 3150
rect 27000 3130 27040 3135
rect 27000 3100 27005 3130
rect 27035 3100 27040 3130
rect 27000 3095 27040 3100
rect 27130 3010 27150 3150
rect 27250 3135 27270 3150
rect 27240 3130 27280 3135
rect 27240 3100 27245 3130
rect 27275 3100 27280 3130
rect 27240 3095 27280 3100
rect 26400 3005 26440 3010
rect 26400 2975 26405 3005
rect 26435 2975 26440 3005
rect 26400 2970 26440 2975
rect 26640 3005 26680 3010
rect 26640 2975 26645 3005
rect 26675 2975 26680 3005
rect 26640 2970 26680 2975
rect 26880 3005 26920 3010
rect 26880 2975 26885 3005
rect 26915 2975 26920 3005
rect 26880 2970 26920 2975
rect 27120 3005 27160 3010
rect 27120 2975 27125 3005
rect 27155 2975 27160 3005
rect 27120 2970 27160 2975
rect 25555 2930 25595 2935
rect 26105 2950 26145 2955
rect 24554 2900 24695 2905
rect 19165 2885 19185 2900
rect 24615 2885 24635 2900
rect 19155 2880 19195 2885
rect 19155 2850 19160 2880
rect 19190 2850 19195 2880
rect 19155 2845 19195 2850
rect 24605 2880 24645 2885
rect 24605 2850 24610 2880
rect 24640 2850 24645 2880
rect 24605 2845 24645 2850
rect 25235 2830 25255 2930
rect 25510 2885 25530 2930
rect 26105 2920 26110 2950
rect 26140 2920 26145 2950
rect 26105 2915 26145 2920
rect 26400 2900 26415 2970
rect 26880 2950 26920 2955
rect 26880 2920 26885 2950
rect 26915 2920 26920 2950
rect 26880 2915 26920 2920
rect 26135 2895 26175 2900
rect 25500 2880 25540 2885
rect 25500 2850 25505 2880
rect 25535 2850 25540 2880
rect 25500 2845 25540 2850
rect 25780 2880 25820 2885
rect 25780 2850 25785 2880
rect 25815 2850 25820 2880
rect 26135 2865 26140 2895
rect 26170 2865 26175 2895
rect 26135 2860 26175 2865
rect 26255 2895 26295 2900
rect 26255 2865 26260 2895
rect 26290 2865 26295 2895
rect 26255 2860 26295 2865
rect 26375 2895 26415 2900
rect 26375 2865 26380 2895
rect 26410 2865 26415 2895
rect 26375 2860 26415 2865
rect 26495 2895 26535 2900
rect 26495 2865 26500 2895
rect 26530 2865 26535 2895
rect 26495 2860 26535 2865
rect 26615 2895 26655 2900
rect 26615 2865 26620 2895
rect 26650 2865 26655 2895
rect 26615 2860 26655 2865
rect 25780 2845 25820 2850
rect 18585 2825 18625 2830
rect 18585 2795 18590 2825
rect 18620 2795 18625 2825
rect 18585 2790 18625 2795
rect 19245 2825 19285 2830
rect 19245 2795 19250 2825
rect 19280 2795 19285 2825
rect 19245 2790 19285 2795
rect 24515 2825 24555 2830
rect 24515 2795 24520 2825
rect 24550 2795 24555 2825
rect 24515 2790 24555 2795
rect 25225 2825 25265 2830
rect 25225 2795 25230 2825
rect 25260 2795 25265 2825
rect 25225 2790 25265 2795
rect 18200 2705 18240 2710
rect 18200 2675 18205 2705
rect 18235 2675 18240 2705
rect 18200 2670 18240 2675
rect 18310 2705 18350 2710
rect 18310 2675 18315 2705
rect 18345 2675 18350 2705
rect 18310 2670 18350 2675
rect 18420 2705 18460 2710
rect 18420 2675 18425 2705
rect 18455 2675 18460 2705
rect 18420 2670 18460 2675
rect 18530 2705 18570 2710
rect 18530 2675 18535 2705
rect 18565 2675 18570 2705
rect 18530 2670 18570 2675
rect 18640 2705 18680 2710
rect 18640 2675 18645 2705
rect 18675 2675 18680 2705
rect 18640 2670 18680 2675
rect 18750 2705 18790 2710
rect 18750 2675 18755 2705
rect 18785 2675 18790 2705
rect 18750 2670 18790 2675
rect 18255 2435 18295 2440
rect 18255 2405 18260 2435
rect 18290 2405 18295 2435
rect 18255 2400 18295 2405
rect 18365 2435 18405 2440
rect 18365 2405 18370 2435
rect 18400 2405 18405 2435
rect 18365 2400 18405 2405
rect 18475 2435 18515 2440
rect 18475 2405 18480 2435
rect 18510 2405 18515 2435
rect 18475 2400 18515 2405
rect 18585 2435 18625 2440
rect 18585 2405 18590 2435
rect 18620 2405 18625 2435
rect 18585 2400 18625 2405
rect 18695 2435 18735 2440
rect 18695 2405 18700 2435
rect 18730 2405 18735 2435
rect 18695 2400 18735 2405
rect 18940 2435 18980 2440
rect 18940 2405 18945 2435
rect 18975 2405 18980 2435
rect 18940 2400 18980 2405
rect 18015 2375 18055 2380
rect 18015 2345 18020 2375
rect 18050 2345 18055 2375
rect 18015 2340 18055 2345
rect 18225 2375 18265 2380
rect 18225 2345 18230 2375
rect 18260 2345 18265 2375
rect 18225 2340 18265 2345
rect 18255 2315 18295 2320
rect 18255 2285 18260 2315
rect 18290 2285 18295 2315
rect 18255 2280 18295 2285
rect 18365 2315 18405 2320
rect 18365 2285 18370 2315
rect 18400 2285 18405 2315
rect 18365 2280 18405 2285
rect 18475 2315 18515 2320
rect 18475 2285 18480 2315
rect 18510 2285 18515 2315
rect 18475 2280 18515 2285
rect 18585 2315 18625 2320
rect 18585 2285 18590 2315
rect 18620 2285 18625 2315
rect 18585 2280 18625 2285
rect 18695 2315 18735 2320
rect 18695 2285 18700 2315
rect 18730 2285 18735 2315
rect 18695 2280 18735 2285
rect 18895 2315 18935 2320
rect 18895 2285 18900 2315
rect 18930 2285 18935 2315
rect 18895 2280 18935 2285
rect 18905 1950 18925 2280
rect 18950 2005 18970 2400
rect 19255 2120 19275 2790
rect 24525 2120 24545 2790
rect 25060 2705 25100 2710
rect 25060 2675 25065 2705
rect 25095 2675 25100 2705
rect 25060 2670 25100 2675
rect 25170 2705 25210 2710
rect 25170 2675 25175 2705
rect 25205 2675 25210 2705
rect 25170 2670 25210 2675
rect 25280 2705 25320 2710
rect 25280 2675 25285 2705
rect 25315 2675 25320 2705
rect 25280 2670 25320 2675
rect 25390 2705 25430 2710
rect 25390 2675 25395 2705
rect 25425 2675 25430 2705
rect 25390 2670 25430 2675
rect 25500 2705 25540 2710
rect 25500 2675 25505 2705
rect 25535 2675 25540 2705
rect 25500 2670 25540 2675
rect 25610 2705 25650 2710
rect 25610 2675 25615 2705
rect 25645 2675 25650 2705
rect 25610 2670 25650 2675
rect 24870 2435 24910 2440
rect 24870 2405 24875 2435
rect 24905 2405 24910 2435
rect 24870 2400 24910 2405
rect 25115 2435 25155 2440
rect 25115 2405 25120 2435
rect 25150 2405 25155 2435
rect 25115 2400 25155 2405
rect 25225 2435 25265 2440
rect 25225 2405 25230 2435
rect 25260 2405 25265 2435
rect 25225 2400 25265 2405
rect 25335 2435 25375 2440
rect 25335 2405 25340 2435
rect 25370 2405 25375 2435
rect 25335 2400 25375 2405
rect 25445 2435 25485 2440
rect 25445 2405 25450 2435
rect 25480 2405 25485 2435
rect 25445 2400 25485 2405
rect 25555 2435 25595 2440
rect 25555 2405 25560 2435
rect 25590 2405 25595 2435
rect 25555 2400 25595 2405
rect 19240 2110 19290 2120
rect 19240 2080 19250 2110
rect 19280 2080 19290 2110
rect 19240 2070 19290 2080
rect 24510 2110 24560 2120
rect 24510 2080 24520 2110
rect 24550 2080 24560 2110
rect 24510 2070 24560 2080
rect 18995 2005 19030 2010
rect 18940 2000 18980 2005
rect 18940 1970 18945 2000
rect 18975 1970 18980 2000
rect 18940 1965 18980 1970
rect 18995 1965 19030 1970
rect 19055 2005 19090 2011
rect 19055 1965 19090 1970
rect 19115 2005 19150 2010
rect 19115 1965 19150 1970
rect 19175 2005 19210 2011
rect 19175 1965 19210 1970
rect 19060 1950 19080 1965
rect 18200 1945 18240 1950
rect 18200 1915 18205 1945
rect 18235 1915 18240 1945
rect 18200 1910 18240 1915
rect 18310 1945 18350 1950
rect 18310 1915 18315 1945
rect 18345 1915 18350 1945
rect 18310 1910 18350 1915
rect 18420 1945 18460 1950
rect 18420 1915 18425 1945
rect 18455 1915 18460 1945
rect 18420 1910 18460 1915
rect 18530 1945 18570 1950
rect 18530 1915 18535 1945
rect 18565 1915 18570 1945
rect 18530 1910 18570 1915
rect 18640 1945 18680 1950
rect 18640 1915 18645 1945
rect 18675 1915 18680 1945
rect 18640 1910 18680 1915
rect 18750 1945 18790 1950
rect 18750 1915 18755 1945
rect 18785 1915 18790 1945
rect 18750 1910 18790 1915
rect 18895 1945 18935 1950
rect 18895 1915 18900 1945
rect 18930 1915 18935 1945
rect 18895 1910 18935 1915
rect 19050 1945 19090 1950
rect 19050 1915 19055 1945
rect 19085 1915 19090 1945
rect 19050 1910 19090 1915
rect 19180 1900 19200 1965
rect 19170 1895 19210 1900
rect 19170 1865 19175 1895
rect 19205 1865 19210 1895
rect 19170 1860 19210 1865
rect 18075 1760 18115 1765
rect 18075 1730 18080 1760
rect 18110 1730 18115 1760
rect 18075 1725 18115 1730
rect 18405 1760 18445 1765
rect 18405 1730 18410 1760
rect 18440 1730 18445 1760
rect 18405 1725 18445 1730
rect 18995 1760 19035 1765
rect 18995 1730 19000 1760
rect 19030 1730 19035 1760
rect 18995 1725 19035 1730
rect 18085 1395 18105 1725
rect 18415 1710 18435 1725
rect 18305 1705 18345 1710
rect 18305 1675 18310 1705
rect 18340 1675 18345 1705
rect 18305 1670 18345 1675
rect 18408 1700 18442 1710
rect 18408 1680 18416 1700
rect 18434 1680 18442 1700
rect 18408 1670 18442 1680
rect 18505 1705 18545 1710
rect 18505 1675 18510 1705
rect 18540 1675 18545 1705
rect 18505 1670 18545 1675
rect 18705 1705 18745 1710
rect 18705 1675 18710 1705
rect 18740 1675 18745 1705
rect 18705 1670 18745 1675
rect 18930 1705 18970 1710
rect 18930 1675 18935 1705
rect 18965 1675 18970 1705
rect 18930 1670 18970 1675
rect 18940 1650 18960 1670
rect 19005 1650 19025 1725
rect 19255 1710 19275 2070
rect 24525 1710 24545 2070
rect 24640 2005 24675 2011
rect 24640 1965 24675 1970
rect 24700 2005 24735 2010
rect 24700 1965 24735 1970
rect 24760 2005 24795 2011
rect 24760 1965 24795 1970
rect 24820 2005 24855 2010
rect 24880 2005 24900 2400
rect 25790 2380 25810 2845
rect 26075 2475 26115 2480
rect 26075 2445 26080 2475
rect 26110 2445 26115 2475
rect 26075 2440 26115 2445
rect 26195 2475 26235 2480
rect 26195 2445 26200 2475
rect 26230 2445 26235 2475
rect 26195 2440 26235 2445
rect 26315 2475 26355 2480
rect 26315 2445 26320 2475
rect 26350 2445 26355 2475
rect 26315 2440 26355 2445
rect 26378 2470 26412 2480
rect 26378 2450 26386 2470
rect 26404 2450 26412 2470
rect 26378 2440 26412 2450
rect 26435 2475 26475 2480
rect 26435 2445 26440 2475
rect 26470 2445 26475 2475
rect 26435 2440 26475 2445
rect 26555 2475 26595 2480
rect 26555 2445 26560 2475
rect 26590 2445 26595 2475
rect 26555 2440 26595 2445
rect 26675 2475 26715 2480
rect 26675 2445 26680 2475
rect 26710 2445 26715 2475
rect 26675 2440 26715 2445
rect 26330 2380 26350 2440
rect 26385 2425 26405 2440
rect 26890 2425 26910 2915
rect 27255 2900 27275 3095
rect 27370 3010 27390 3150
rect 27490 3135 27510 3150
rect 27480 3130 27520 3135
rect 27480 3100 27485 3130
rect 27515 3100 27520 3130
rect 27480 3095 27520 3100
rect 27360 3005 27400 3010
rect 27360 2975 27365 3005
rect 27395 2975 27400 3005
rect 27360 2970 27400 2975
rect 27155 2895 27195 2900
rect 27155 2865 27160 2895
rect 27190 2865 27195 2895
rect 27155 2860 27195 2865
rect 27255 2895 27315 2900
rect 27255 2865 27280 2895
rect 27310 2865 27315 2895
rect 27255 2860 27315 2865
rect 27395 2895 27435 2900
rect 27395 2865 27400 2895
rect 27430 2865 27435 2895
rect 27395 2860 27435 2865
rect 27515 2895 27555 2900
rect 27515 2865 27520 2895
rect 27550 2865 27555 2895
rect 27515 2860 27555 2865
rect 27635 2895 27675 2900
rect 27635 2865 27640 2895
rect 27670 2865 27675 2895
rect 27635 2860 27675 2865
rect 27095 2475 27135 2480
rect 27095 2445 27100 2475
rect 27130 2445 27135 2475
rect 27095 2440 27135 2445
rect 27215 2475 27255 2480
rect 27215 2445 27220 2475
rect 27250 2445 27255 2475
rect 27215 2440 27255 2445
rect 27335 2475 27375 2480
rect 27335 2445 27340 2475
rect 27370 2445 27375 2475
rect 27335 2440 27375 2445
rect 27398 2470 27432 2480
rect 27398 2450 27406 2470
rect 27424 2450 27432 2470
rect 27398 2440 27432 2450
rect 27455 2475 27495 2480
rect 27455 2445 27460 2475
rect 27490 2445 27495 2475
rect 27455 2440 27495 2445
rect 27575 2475 27615 2480
rect 27575 2445 27580 2475
rect 27610 2445 27615 2475
rect 27575 2440 27615 2445
rect 27695 2475 27735 2480
rect 27695 2445 27700 2475
rect 27730 2445 27735 2475
rect 27695 2440 27735 2445
rect 26375 2420 26415 2425
rect 26375 2390 26380 2420
rect 26410 2390 26415 2420
rect 26375 2385 26415 2390
rect 26880 2420 26920 2425
rect 26880 2390 26885 2420
rect 26915 2390 26920 2420
rect 26880 2385 26920 2390
rect 27335 2380 27355 2440
rect 27405 2425 27425 2440
rect 27395 2420 27435 2425
rect 27395 2390 27400 2420
rect 27430 2390 27435 2420
rect 27395 2385 27435 2390
rect 25585 2375 25625 2380
rect 25585 2345 25590 2375
rect 25620 2345 25625 2375
rect 25585 2340 25625 2345
rect 25780 2375 25820 2380
rect 25780 2345 25785 2375
rect 25815 2345 25820 2375
rect 25780 2340 25820 2345
rect 26320 2375 26360 2380
rect 26320 2345 26325 2375
rect 26355 2345 26360 2375
rect 26320 2340 26360 2345
rect 27320 2375 27360 2380
rect 27320 2345 27325 2375
rect 27355 2345 27360 2375
rect 27320 2340 27360 2345
rect 26000 2325 26040 2330
rect 24915 2315 24955 2320
rect 24915 2285 24920 2315
rect 24950 2285 24955 2315
rect 24915 2280 24955 2285
rect 25115 2315 25155 2320
rect 25115 2285 25120 2315
rect 25150 2285 25155 2315
rect 25115 2280 25155 2285
rect 25225 2315 25265 2320
rect 25225 2285 25230 2315
rect 25260 2285 25265 2315
rect 25225 2280 25265 2285
rect 25335 2315 25375 2320
rect 25335 2285 25340 2315
rect 25370 2285 25375 2315
rect 25335 2280 25375 2285
rect 25445 2315 25485 2320
rect 25445 2285 25450 2315
rect 25480 2285 25485 2315
rect 25445 2280 25485 2285
rect 25555 2315 25595 2320
rect 25555 2285 25560 2315
rect 25590 2285 25595 2315
rect 26000 2295 26005 2325
rect 26035 2295 26040 2325
rect 26000 2290 26040 2295
rect 25555 2280 25595 2285
rect 24820 1965 24855 1970
rect 24870 2000 24910 2005
rect 24870 1970 24875 2000
rect 24905 1970 24910 2000
rect 24870 1965 24910 1970
rect 24650 1900 24670 1965
rect 24770 1950 24790 1965
rect 24925 1950 24945 2280
rect 25800 2180 25840 2185
rect 25800 2150 25805 2180
rect 25835 2150 25840 2180
rect 25800 2145 25840 2150
rect 24760 1945 24800 1950
rect 24760 1915 24765 1945
rect 24795 1915 24800 1945
rect 24760 1910 24800 1915
rect 24915 1945 24955 1950
rect 24915 1915 24920 1945
rect 24950 1915 24955 1945
rect 24915 1910 24955 1915
rect 25060 1945 25100 1950
rect 25060 1915 25065 1945
rect 25095 1915 25100 1945
rect 25060 1910 25100 1915
rect 25170 1945 25210 1950
rect 25170 1915 25175 1945
rect 25205 1915 25210 1945
rect 25170 1910 25210 1915
rect 25280 1945 25320 1950
rect 25280 1915 25285 1945
rect 25315 1915 25320 1945
rect 25280 1910 25320 1915
rect 25390 1945 25430 1950
rect 25390 1915 25395 1945
rect 25425 1915 25430 1945
rect 25390 1910 25430 1915
rect 25500 1945 25540 1950
rect 25500 1915 25505 1945
rect 25535 1915 25540 1945
rect 25500 1910 25540 1915
rect 25610 1945 25650 1950
rect 25610 1915 25615 1945
rect 25645 1915 25650 1945
rect 25610 1910 25650 1915
rect 24640 1895 24680 1900
rect 24640 1865 24645 1895
rect 24675 1865 24680 1895
rect 24640 1860 24680 1865
rect 24815 1760 24855 1765
rect 24815 1730 24820 1760
rect 24850 1730 24855 1760
rect 24815 1725 24855 1730
rect 25405 1760 25445 1765
rect 25405 1730 25410 1760
rect 25440 1730 25445 1760
rect 25405 1725 25445 1730
rect 25735 1760 25775 1765
rect 25735 1730 25740 1760
rect 25770 1730 25775 1760
rect 25735 1725 25775 1730
rect 19245 1705 19285 1710
rect 19245 1675 19250 1705
rect 19280 1675 19285 1705
rect 19245 1670 19285 1675
rect 24515 1705 24555 1710
rect 24515 1675 24520 1705
rect 24550 1675 24555 1705
rect 24515 1670 24555 1675
rect 24825 1650 24845 1725
rect 25415 1710 25435 1725
rect 24880 1705 24920 1710
rect 24880 1675 24885 1705
rect 24915 1675 24920 1705
rect 24880 1670 24920 1675
rect 25105 1705 25145 1710
rect 25105 1675 25110 1705
rect 25140 1675 25145 1705
rect 25105 1670 25145 1675
rect 25305 1705 25345 1710
rect 25305 1675 25310 1705
rect 25340 1675 25345 1705
rect 25305 1670 25345 1675
rect 25408 1700 25442 1710
rect 25408 1680 25416 1700
rect 25434 1680 25442 1700
rect 25408 1670 25442 1680
rect 25505 1705 25545 1710
rect 25505 1675 25510 1705
rect 25540 1675 25545 1705
rect 25505 1670 25545 1675
rect 24890 1650 24910 1670
rect 18935 1645 18970 1650
rect 18935 1605 18970 1610
rect 18995 1645 19030 1650
rect 18995 1605 19030 1610
rect 24820 1645 24855 1650
rect 24820 1605 24855 1610
rect 24880 1645 24915 1650
rect 24880 1605 24915 1610
rect 25745 1395 25765 1725
rect 18075 1390 18115 1395
rect 18075 1360 18080 1390
rect 18110 1360 18115 1390
rect 18075 1355 18115 1360
rect 25735 1390 25775 1395
rect 25735 1360 25740 1390
rect 25770 1360 25775 1390
rect 25735 1355 25775 1360
rect 18405 935 18445 940
rect 18405 905 18410 935
rect 18440 905 18445 935
rect 18405 900 18445 905
rect 18605 935 18645 940
rect 18605 905 18610 935
rect 18640 905 18645 935
rect 18605 900 18645 905
rect 25205 935 25245 940
rect 25205 905 25210 935
rect 25240 905 25245 935
rect 25205 900 25245 905
rect 25405 935 25445 940
rect 25405 905 25410 935
rect 25440 905 25445 935
rect 25405 900 25445 905
rect 17960 860 18000 865
rect 17960 830 17965 860
rect 17995 830 18000 860
rect 17960 825 18000 830
rect 15800 800 15840 805
rect 15800 770 15805 800
rect 15835 770 15840 800
rect 15800 765 15840 770
rect 16305 800 16345 805
rect 16305 770 16310 800
rect 16340 770 16345 800
rect 16305 765 16345 770
rect 16375 800 16415 805
rect 16375 770 16380 800
rect 16410 770 16415 800
rect 16375 765 16415 770
rect 16445 800 16485 805
rect 16445 770 16450 800
rect 16480 770 16485 800
rect 16445 765 16485 770
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 16935 765 16975 775
rect 17045 800 17085 805
rect 17045 770 17050 800
rect 17080 770 17085 800
rect 17045 765 17085 770
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17155 765 17195 775
rect 17265 800 17305 805
rect 17265 770 17270 800
rect 17300 770 17305 800
rect 17265 765 17305 770
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 17375 765 17415 775
rect 17485 800 17525 805
rect 17485 770 17490 800
rect 17520 770 17525 800
rect 17485 765 17525 770
rect 17905 800 17945 805
rect 17905 770 17910 800
rect 17940 770 17945 800
rect 17905 765 17945 770
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 730 2560 760
rect 2520 725 2560 730
rect 3130 760 3170 765
rect 3130 730 3135 760
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 730 3665 760
rect 3625 725 3665 730
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 760 4025 765
rect 3985 730 3990 760
rect 4020 730 4025 760
rect 3985 725 4025 730
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 760 4385 765
rect 4345 730 4350 760
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 730 4565 760
rect 4525 725 4565 730
rect 4705 760 4745 765
rect 4705 730 4710 760
rect 4740 730 4745 760
rect 4705 725 4745 730
rect 4885 760 4925 765
rect 4885 730 4890 760
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3275 295 3295 725
rect 3455 710 3475 725
rect 3815 710 3835 725
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 675 3485 705
rect 3445 670 3485 675
rect 3805 705 3845 710
rect 3805 675 3810 705
rect 3840 675 3845 705
rect 3805 670 3845 675
rect 3815 295 3835 670
rect 3995 295 4015 725
rect 4175 710 4195 725
rect 4165 705 4205 710
rect 4165 675 4170 705
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 4715 295 4735 725
rect 16990 680 17030 685
rect 16990 650 16995 680
rect 17025 650 17030 680
rect 16990 645 17030 650
rect 17100 680 17140 685
rect 17100 650 17105 680
rect 17135 650 17140 680
rect 17100 645 17140 650
rect 17210 680 17250 685
rect 17210 650 17215 680
rect 17245 650 17250 680
rect 17210 645 17250 650
rect 17320 680 17360 685
rect 17320 650 17325 680
rect 17355 650 17360 680
rect 17320 645 17360 650
rect 17430 680 17470 685
rect 17430 650 17435 680
rect 17465 650 17470 680
rect 17430 645 17470 650
rect 25810 605 25830 2145
rect 26010 1900 26030 2290
rect 26330 2240 26350 2340
rect 27330 2285 27350 2340
rect 27880 2330 27900 4035
rect 27970 3825 28010 3830
rect 27970 3795 27975 3825
rect 28005 3795 28010 3825
rect 27970 3790 28010 3795
rect 27915 3780 27955 3785
rect 27915 3750 27920 3780
rect 27950 3750 27955 3780
rect 27915 3745 27955 3750
rect 27870 2325 27910 2330
rect 27870 2295 27875 2325
rect 27905 2295 27910 2325
rect 27870 2290 27910 2295
rect 26440 2280 26480 2285
rect 26440 2250 26445 2280
rect 26475 2250 26480 2280
rect 26440 2245 26480 2250
rect 26660 2280 26700 2285
rect 26660 2250 26665 2280
rect 26695 2250 26700 2280
rect 26660 2245 26700 2250
rect 26880 2280 26920 2285
rect 26880 2250 26885 2280
rect 26915 2250 26920 2280
rect 26880 2245 26920 2250
rect 27100 2280 27140 2285
rect 27100 2250 27105 2280
rect 27135 2250 27140 2280
rect 27100 2245 27140 2250
rect 27320 2280 27360 2285
rect 27320 2250 27325 2280
rect 27355 2250 27360 2280
rect 27320 2245 27360 2250
rect 26330 2235 26370 2240
rect 26330 2205 26335 2235
rect 26365 2205 26370 2235
rect 26330 2200 26370 2205
rect 26340 2185 26360 2200
rect 26450 2185 26470 2245
rect 26550 2235 26590 2240
rect 26550 2205 26555 2235
rect 26585 2205 26590 2235
rect 26550 2200 26590 2205
rect 26560 2185 26580 2200
rect 26670 2185 26690 2245
rect 26770 2235 26810 2240
rect 26770 2205 26775 2235
rect 26805 2205 26810 2235
rect 26770 2200 26810 2205
rect 26780 2185 26800 2200
rect 26890 2185 26910 2245
rect 26990 2235 27030 2240
rect 26990 2205 26995 2235
rect 27025 2205 27030 2235
rect 26990 2200 27030 2205
rect 27000 2185 27020 2200
rect 27110 2185 27130 2245
rect 27210 2235 27250 2240
rect 27210 2205 27215 2235
rect 27245 2205 27250 2235
rect 27210 2200 27250 2205
rect 27220 2185 27240 2200
rect 27330 2185 27350 2245
rect 27430 2235 27470 2240
rect 27430 2205 27435 2235
rect 27465 2205 27470 2235
rect 27430 2200 27470 2205
rect 27440 2185 27460 2200
rect 26330 2175 26370 2185
rect 26330 2155 26340 2175
rect 26360 2155 26370 2175
rect 26330 2145 26370 2155
rect 26440 2175 26480 2185
rect 26440 2155 26450 2175
rect 26470 2155 26480 2175
rect 26440 2145 26480 2155
rect 26550 2175 26590 2185
rect 26550 2155 26560 2175
rect 26580 2155 26590 2175
rect 26550 2145 26590 2155
rect 26660 2175 26700 2185
rect 26660 2155 26670 2175
rect 26690 2155 26700 2175
rect 26660 2145 26700 2155
rect 26770 2175 26810 2185
rect 26770 2155 26780 2175
rect 26800 2155 26810 2175
rect 26770 2145 26810 2155
rect 26828 2180 26862 2185
rect 26828 2150 26831 2180
rect 26859 2150 26862 2180
rect 26828 2145 26862 2150
rect 26880 2175 26920 2185
rect 26880 2155 26890 2175
rect 26910 2155 26920 2175
rect 26880 2145 26920 2155
rect 26990 2175 27030 2185
rect 26990 2155 27000 2175
rect 27020 2155 27030 2175
rect 26990 2145 27030 2155
rect 27100 2175 27140 2185
rect 27100 2155 27110 2175
rect 27130 2155 27140 2175
rect 27100 2145 27140 2155
rect 27210 2175 27250 2185
rect 27210 2155 27220 2175
rect 27240 2155 27250 2175
rect 27210 2145 27250 2155
rect 27320 2175 27360 2185
rect 27320 2155 27330 2175
rect 27350 2155 27360 2175
rect 27320 2145 27360 2155
rect 27430 2175 27470 2185
rect 27430 2155 27440 2175
rect 27460 2155 27470 2175
rect 27430 2145 27470 2155
rect 26385 1960 26425 1965
rect 26385 1930 26390 1960
rect 26420 1930 26425 1960
rect 26385 1925 26425 1930
rect 26495 1955 26535 1965
rect 26495 1935 26505 1955
rect 26525 1935 26535 1955
rect 26495 1925 26535 1935
rect 26605 1960 26645 1965
rect 26605 1930 26610 1960
rect 26640 1930 26645 1960
rect 26605 1925 26645 1930
rect 26715 1955 26755 1965
rect 26715 1935 26725 1955
rect 26745 1935 26755 1955
rect 26715 1925 26755 1935
rect 26825 1960 26865 1965
rect 26825 1930 26830 1960
rect 26860 1930 26865 1960
rect 26825 1925 26865 1930
rect 26935 1955 26975 1965
rect 26935 1935 26945 1955
rect 26965 1935 26975 1955
rect 26935 1925 26975 1935
rect 27045 1960 27085 1965
rect 27045 1930 27050 1960
rect 27080 1930 27085 1960
rect 27045 1925 27085 1930
rect 27155 1955 27195 1965
rect 27155 1935 27165 1955
rect 27185 1935 27195 1955
rect 27155 1925 27195 1935
rect 27245 1960 27305 1965
rect 27245 1930 27270 1960
rect 27300 1930 27305 1960
rect 27245 1925 27305 1930
rect 27375 1955 27415 1965
rect 27375 1935 27385 1955
rect 27405 1935 27415 1955
rect 27375 1925 27415 1935
rect 26505 1910 26525 1925
rect 26725 1910 26745 1925
rect 26945 1910 26965 1925
rect 27165 1910 27185 1925
rect 26495 1905 26555 1910
rect 26000 1895 26040 1900
rect 26000 1865 26005 1895
rect 26035 1865 26040 1895
rect 26495 1875 26500 1905
rect 26530 1875 26555 1905
rect 26495 1870 26555 1875
rect 26715 1905 26755 1910
rect 26715 1875 26720 1905
rect 26750 1875 26755 1905
rect 26715 1870 26755 1875
rect 26935 1905 26975 1910
rect 26935 1875 26940 1905
rect 26970 1875 26975 1905
rect 26935 1870 26975 1875
rect 27155 1905 27195 1910
rect 27155 1875 27160 1905
rect 27190 1875 27195 1905
rect 27155 1870 27195 1875
rect 26000 1860 26040 1865
rect 26190 1850 26230 1855
rect 26190 1820 26195 1850
rect 26225 1820 26230 1850
rect 26190 1815 26230 1820
rect 26410 1850 26450 1855
rect 26410 1820 26415 1850
rect 26445 1820 26450 1850
rect 26410 1815 26450 1820
rect 26200 1780 26220 1815
rect 26420 1780 26440 1815
rect 26190 1770 26230 1780
rect 26085 1760 26125 1765
rect 26085 1730 26090 1760
rect 26120 1730 26125 1760
rect 26190 1750 26200 1770
rect 26220 1750 26230 1770
rect 26410 1770 26450 1780
rect 26190 1740 26230 1750
rect 26305 1760 26345 1765
rect 26085 1725 26125 1730
rect 26305 1730 26310 1760
rect 26340 1730 26345 1760
rect 26410 1750 26420 1770
rect 26440 1750 26450 1770
rect 26535 1765 26555 1870
rect 27245 1855 27265 1925
rect 27385 1910 27405 1925
rect 27375 1905 27415 1910
rect 27375 1875 27380 1905
rect 27410 1875 27415 1905
rect 27880 1880 27900 2290
rect 27375 1870 27415 1875
rect 27870 1875 27910 1880
rect 26640 1850 26680 1855
rect 26640 1820 26645 1850
rect 26675 1820 26680 1850
rect 26640 1815 26680 1820
rect 27230 1850 27270 1855
rect 27230 1820 27235 1850
rect 27265 1820 27270 1850
rect 27230 1815 27270 1820
rect 27450 1850 27490 1855
rect 27450 1820 27455 1850
rect 27485 1820 27490 1850
rect 27450 1815 27490 1820
rect 27680 1850 27720 1855
rect 27680 1820 27685 1850
rect 27715 1820 27720 1850
rect 27870 1845 27875 1875
rect 27905 1845 27910 1875
rect 27870 1840 27910 1845
rect 27680 1815 27720 1820
rect 26650 1780 26670 1815
rect 26820 1805 26860 1810
rect 26640 1770 26680 1780
rect 26820 1775 26825 1805
rect 26855 1775 26860 1805
rect 26820 1770 26860 1775
rect 26940 1805 26980 1810
rect 26940 1775 26945 1805
rect 26975 1775 26980 1805
rect 27240 1780 27260 1815
rect 27460 1780 27480 1815
rect 27690 1780 27710 1815
rect 26940 1770 26980 1775
rect 27230 1770 27270 1780
rect 26410 1740 26450 1750
rect 26525 1760 26565 1765
rect 26305 1725 26345 1730
rect 26525 1730 26530 1760
rect 26560 1730 26565 1760
rect 26640 1750 26650 1770
rect 26670 1750 26680 1770
rect 26640 1740 26680 1750
rect 26525 1725 26565 1730
rect 26830 1720 26850 1770
rect 26950 1720 26970 1770
rect 27125 1760 27165 1765
rect 27125 1730 27130 1760
rect 27160 1730 27165 1760
rect 27230 1750 27240 1770
rect 27260 1750 27270 1770
rect 27450 1770 27490 1780
rect 27230 1740 27270 1750
rect 27345 1760 27385 1765
rect 27125 1725 27165 1730
rect 27345 1730 27350 1760
rect 27380 1730 27385 1760
rect 27450 1750 27460 1770
rect 27480 1750 27490 1770
rect 27680 1770 27720 1780
rect 27450 1740 27490 1750
rect 27565 1760 27605 1765
rect 27345 1725 27385 1730
rect 27565 1730 27570 1760
rect 27600 1730 27605 1760
rect 27680 1750 27690 1770
rect 27710 1750 27720 1770
rect 27680 1740 27720 1750
rect 27565 1725 27605 1730
rect 26237 1715 26269 1720
rect 26237 1685 26240 1715
rect 26266 1685 26269 1715
rect 26237 1680 26269 1685
rect 26457 1715 26489 1720
rect 26457 1685 26460 1715
rect 26486 1685 26489 1715
rect 26457 1680 26489 1685
rect 26601 1715 26633 1720
rect 26601 1685 26604 1715
rect 26630 1685 26633 1715
rect 26601 1680 26633 1685
rect 26820 1710 26850 1720
rect 26820 1690 26825 1710
rect 26845 1690 26850 1710
rect 26820 1680 26850 1690
rect 26867 1715 26899 1720
rect 26867 1685 26870 1715
rect 26896 1685 26899 1715
rect 26867 1680 26899 1685
rect 26950 1710 26980 1720
rect 26950 1690 26955 1710
rect 26975 1690 26980 1710
rect 26950 1680 26980 1690
rect 27277 1715 27309 1720
rect 27277 1685 27280 1715
rect 27306 1685 27309 1715
rect 27277 1680 27309 1685
rect 27497 1715 27529 1720
rect 27497 1685 27500 1715
rect 27526 1685 27529 1715
rect 27497 1680 27529 1685
rect 27641 1715 27673 1720
rect 27641 1685 27644 1715
rect 27670 1685 27673 1715
rect 27641 1680 27673 1685
rect 26106 1495 26138 1500
rect 26106 1465 26109 1495
rect 26135 1465 26138 1495
rect 26106 1460 26138 1465
rect 26305 1495 26345 1500
rect 26305 1465 26310 1495
rect 26340 1465 26345 1495
rect 26305 1460 26345 1465
rect 26525 1495 26565 1500
rect 26525 1465 26530 1495
rect 26560 1465 26565 1495
rect 26525 1460 26565 1465
rect 26825 1490 26855 1500
rect 26825 1470 26830 1490
rect 26850 1470 26855 1490
rect 26825 1460 26855 1470
rect 26875 1490 26905 1500
rect 26875 1470 26880 1490
rect 26900 1470 26905 1490
rect 26875 1460 26905 1470
rect 26922 1495 26954 1500
rect 26922 1465 26925 1495
rect 26951 1465 26954 1495
rect 26922 1460 26954 1465
rect 27146 1495 27178 1500
rect 27146 1465 27149 1495
rect 27175 1465 27178 1495
rect 27146 1460 27178 1465
rect 27345 1495 27385 1500
rect 27345 1465 27350 1495
rect 27380 1465 27385 1495
rect 27345 1460 27385 1465
rect 27565 1495 27605 1500
rect 27565 1465 27570 1495
rect 27600 1465 27605 1495
rect 27565 1460 27605 1465
rect 26145 1435 26185 1440
rect 26145 1405 26150 1435
rect 26180 1405 26185 1435
rect 26145 1400 26185 1405
rect 26250 1435 26290 1440
rect 26250 1405 26255 1435
rect 26285 1405 26290 1435
rect 26250 1400 26290 1405
rect 26360 1435 26400 1440
rect 26360 1405 26365 1435
rect 26395 1405 26400 1435
rect 26360 1400 26400 1405
rect 26470 1435 26510 1440
rect 26470 1405 26475 1435
rect 26505 1405 26510 1435
rect 26470 1400 26510 1405
rect 26580 1435 26620 1440
rect 26580 1405 26585 1435
rect 26615 1405 26620 1435
rect 26580 1400 26620 1405
rect 26830 1250 26850 1460
rect 26005 1245 26045 1250
rect 26005 1215 26010 1245
rect 26040 1215 26045 1245
rect 26005 1210 26045 1215
rect 26810 1245 26850 1250
rect 26810 1215 26815 1245
rect 26845 1215 26850 1245
rect 26810 1210 26850 1215
rect 26015 660 26035 1210
rect 26315 1195 26355 1200
rect 26315 1165 26320 1195
rect 26350 1165 26355 1195
rect 26315 1160 26355 1165
rect 26325 1140 26345 1160
rect 26820 1140 26840 1210
rect 26880 1200 26900 1460
rect 27185 1435 27225 1440
rect 27185 1405 27190 1435
rect 27220 1405 27225 1435
rect 27185 1400 27225 1405
rect 27290 1435 27330 1440
rect 27290 1405 27295 1435
rect 27325 1405 27330 1435
rect 27290 1400 27330 1405
rect 27400 1435 27440 1440
rect 27400 1405 27405 1435
rect 27435 1405 27440 1435
rect 27400 1400 27440 1405
rect 27510 1435 27550 1440
rect 27510 1405 27515 1435
rect 27545 1405 27550 1435
rect 27510 1400 27550 1405
rect 27620 1435 27660 1440
rect 27620 1405 27625 1435
rect 27655 1405 27660 1435
rect 27620 1400 27660 1405
rect 26880 1195 26920 1200
rect 26880 1165 26885 1195
rect 26915 1165 26920 1195
rect 26880 1160 26920 1165
rect 27925 1155 27945 3745
rect 27595 1150 27635 1155
rect 26315 1130 26355 1140
rect 26315 1110 26325 1130
rect 26345 1110 26355 1130
rect 26315 1100 26355 1110
rect 26425 1135 26465 1140
rect 26425 1105 26430 1135
rect 26460 1105 26465 1135
rect 26425 1100 26465 1105
rect 26535 1135 26575 1140
rect 26535 1105 26540 1135
rect 26570 1105 26575 1135
rect 26535 1100 26575 1105
rect 26645 1135 26685 1140
rect 26645 1105 26650 1135
rect 26680 1105 26685 1135
rect 26645 1100 26685 1105
rect 26755 1135 26795 1140
rect 26755 1105 26760 1135
rect 26790 1105 26795 1135
rect 26755 1100 26795 1105
rect 26815 1130 26845 1140
rect 26815 1110 26820 1130
rect 26840 1110 26845 1130
rect 26815 1100 26845 1110
rect 26865 1135 26905 1140
rect 26865 1105 26870 1135
rect 26900 1105 26905 1135
rect 26865 1100 26905 1105
rect 26975 1135 27015 1140
rect 26975 1105 26980 1135
rect 27010 1105 27015 1135
rect 26975 1100 27015 1105
rect 27085 1135 27125 1140
rect 27085 1105 27090 1135
rect 27120 1105 27125 1135
rect 27085 1100 27125 1105
rect 27195 1135 27235 1140
rect 27195 1105 27200 1135
rect 27230 1105 27235 1135
rect 27195 1100 27235 1105
rect 27305 1135 27345 1140
rect 27305 1105 27310 1135
rect 27340 1105 27345 1135
rect 27305 1100 27345 1105
rect 27415 1135 27455 1140
rect 27415 1105 27420 1135
rect 27450 1105 27455 1135
rect 27415 1100 27455 1105
rect 27525 1135 27565 1140
rect 27525 1105 27530 1135
rect 27560 1105 27565 1135
rect 27595 1120 27600 1150
rect 27630 1120 27635 1150
rect 27595 1115 27635 1120
rect 27915 1150 27955 1155
rect 27915 1120 27920 1150
rect 27950 1120 27955 1150
rect 27915 1115 27955 1120
rect 27525 1100 27565 1105
rect 26195 815 26235 820
rect 26195 785 26200 815
rect 26230 785 26235 815
rect 26195 780 26235 785
rect 26260 815 26300 820
rect 26260 785 26265 815
rect 26295 785 26300 815
rect 26260 780 26300 785
rect 26370 815 26410 820
rect 26370 785 26375 815
rect 26405 785 26410 815
rect 26370 780 26410 785
rect 26480 815 26520 820
rect 26480 785 26485 815
rect 26515 785 26520 815
rect 26480 780 26520 785
rect 26590 815 26630 820
rect 26590 785 26595 815
rect 26625 785 26630 815
rect 26590 780 26630 785
rect 26700 815 26740 820
rect 26700 785 26705 815
rect 26735 785 26740 815
rect 26700 780 26740 785
rect 26810 815 26850 820
rect 26810 785 26815 815
rect 26845 785 26850 815
rect 26810 780 26850 785
rect 26920 815 26960 820
rect 26920 785 26925 815
rect 26955 785 26960 815
rect 26920 780 26960 785
rect 27030 815 27070 820
rect 27030 785 27035 815
rect 27065 785 27070 815
rect 27030 780 27070 785
rect 27140 815 27180 820
rect 27140 785 27145 815
rect 27175 785 27180 815
rect 27140 780 27180 785
rect 27250 815 27290 820
rect 27250 785 27255 815
rect 27285 785 27290 815
rect 27250 780 27290 785
rect 27360 815 27400 820
rect 27360 785 27365 815
rect 27395 785 27400 815
rect 27360 780 27400 785
rect 27470 815 27510 820
rect 27470 785 27475 815
rect 27505 785 27510 815
rect 27470 780 27510 785
rect 27585 815 27625 820
rect 27585 785 27590 815
rect 27620 785 27625 815
rect 27585 780 27625 785
rect 26935 660 26975 665
rect 26005 655 26045 660
rect 26005 625 26010 655
rect 26040 625 26045 655
rect 26005 620 26045 625
rect 26505 655 26545 660
rect 26505 625 26510 655
rect 26540 625 26545 655
rect 26935 630 26940 660
rect 26970 630 26975 660
rect 26935 625 26975 630
rect 27155 660 27195 665
rect 27155 630 27160 660
rect 27190 630 27195 660
rect 27155 625 27195 630
rect 27375 660 27415 665
rect 27375 630 27380 660
rect 27410 630 27415 660
rect 27375 625 27415 630
rect 26505 620 26545 625
rect 26515 605 26535 620
rect 26945 605 26965 625
rect 27165 605 27185 625
rect 27385 605 27405 625
rect 27925 605 27945 1115
rect 27980 665 28000 3790
rect 29155 3735 29195 3740
rect 28200 3715 28240 3720
rect 28200 3685 28205 3715
rect 28235 3685 28240 3715
rect 28200 3680 28240 3685
rect 28310 3715 28350 3720
rect 28310 3685 28315 3715
rect 28345 3685 28350 3715
rect 28310 3680 28350 3685
rect 28420 3715 28460 3720
rect 28420 3685 28425 3715
rect 28455 3685 28460 3715
rect 28420 3680 28460 3685
rect 28530 3715 28570 3720
rect 28530 3685 28535 3715
rect 28565 3685 28570 3715
rect 28530 3680 28570 3685
rect 28640 3715 28680 3720
rect 28640 3685 28645 3715
rect 28675 3685 28680 3715
rect 28640 3680 28680 3685
rect 28750 3715 28790 3720
rect 28750 3685 28755 3715
rect 28785 3685 28790 3715
rect 29155 3705 29160 3735
rect 29190 3705 29195 3735
rect 29155 3700 29195 3705
rect 28750 3680 28790 3685
rect 29165 3660 29185 3700
rect 29105 3655 29246 3660
rect 29105 3625 29110 3655
rect 29140 3625 29160 3655
rect 29190 3625 29210 3655
rect 29240 3625 29246 3655
rect 29105 3620 29246 3625
rect 28255 3045 28295 3050
rect 28255 3015 28260 3045
rect 28290 3015 28295 3045
rect 28255 3010 28295 3015
rect 28313 3040 28347 3050
rect 28313 3020 28321 3040
rect 28339 3020 28347 3040
rect 28313 3010 28347 3020
rect 28365 3045 28405 3050
rect 28365 3015 28370 3045
rect 28400 3015 28405 3045
rect 28365 3010 28405 3015
rect 28475 3045 28515 3050
rect 28475 3015 28480 3045
rect 28510 3015 28515 3045
rect 28475 3010 28515 3015
rect 28585 3045 28625 3050
rect 28585 3015 28590 3045
rect 28620 3015 28625 3045
rect 28585 3010 28625 3015
rect 28695 3045 28735 3050
rect 28695 3015 28700 3045
rect 28730 3015 28735 3045
rect 28695 3010 28735 3015
rect 29105 3035 29246 3040
rect 28320 2885 28340 3010
rect 28015 2880 28055 2885
rect 28015 2850 28020 2880
rect 28050 2850 28055 2880
rect 28015 2845 28055 2850
rect 28310 2880 28350 2885
rect 28310 2850 28315 2880
rect 28345 2850 28350 2880
rect 28310 2845 28350 2850
rect 28025 2380 28045 2845
rect 28595 2840 28615 3010
rect 29105 3005 29110 3035
rect 29140 3005 29160 3035
rect 29190 3005 29210 3035
rect 29240 3005 29246 3035
rect 29105 3000 29246 3005
rect 29165 2885 29185 3000
rect 29155 2880 29195 2885
rect 29155 2850 29160 2880
rect 29190 2850 29195 2880
rect 29155 2845 29195 2850
rect 28585 2835 28625 2840
rect 28585 2805 28590 2835
rect 28620 2805 28625 2835
rect 28585 2800 28625 2805
rect 29395 2835 29435 2840
rect 29395 2805 29400 2835
rect 29430 2805 29435 2835
rect 29395 2800 29435 2805
rect 28200 2755 28240 2760
rect 28200 2725 28205 2755
rect 28235 2725 28240 2755
rect 28200 2720 28240 2725
rect 28310 2755 28350 2760
rect 28310 2725 28315 2755
rect 28345 2725 28350 2755
rect 28310 2720 28350 2725
rect 28420 2755 28460 2760
rect 28420 2725 28425 2755
rect 28455 2725 28460 2755
rect 28420 2720 28460 2725
rect 28530 2755 28570 2760
rect 28530 2725 28535 2755
rect 28565 2725 28570 2755
rect 28530 2720 28570 2725
rect 28640 2755 28680 2760
rect 28640 2725 28645 2755
rect 28675 2725 28680 2755
rect 28640 2720 28680 2725
rect 28750 2755 28790 2760
rect 28750 2725 28755 2755
rect 28785 2725 28790 2755
rect 28750 2720 28790 2725
rect 28255 2485 28295 2490
rect 28255 2455 28260 2485
rect 28290 2455 28295 2485
rect 28255 2450 28295 2455
rect 28313 2480 28347 2490
rect 28313 2460 28321 2480
rect 28339 2460 28347 2480
rect 28313 2450 28347 2460
rect 28365 2485 28405 2490
rect 28365 2455 28370 2485
rect 28400 2455 28405 2485
rect 28365 2450 28405 2455
rect 28475 2485 28515 2490
rect 28475 2455 28480 2485
rect 28510 2455 28515 2485
rect 28475 2450 28515 2455
rect 28585 2485 28625 2490
rect 28585 2455 28590 2485
rect 28620 2455 28625 2485
rect 28585 2450 28625 2455
rect 28695 2485 28735 2490
rect 28695 2455 28700 2485
rect 28730 2455 28735 2485
rect 28695 2450 28735 2455
rect 28940 2485 28980 2490
rect 28940 2455 28945 2485
rect 28975 2455 28980 2485
rect 28940 2450 28980 2455
rect 28320 2380 28340 2450
rect 28015 2375 28055 2380
rect 28015 2345 28020 2375
rect 28050 2345 28055 2375
rect 28015 2340 28055 2345
rect 28310 2375 28350 2380
rect 28310 2345 28315 2375
rect 28345 2345 28350 2375
rect 28310 2340 28350 2345
rect 28320 2300 28340 2340
rect 28255 2295 28295 2300
rect 28255 2265 28260 2295
rect 28290 2265 28295 2295
rect 28255 2260 28295 2265
rect 28313 2290 28347 2300
rect 28313 2270 28321 2290
rect 28339 2270 28347 2290
rect 28313 2260 28347 2270
rect 28365 2295 28405 2300
rect 28365 2265 28370 2295
rect 28400 2265 28405 2295
rect 28365 2260 28405 2265
rect 28475 2295 28515 2300
rect 28475 2265 28480 2295
rect 28510 2265 28515 2295
rect 28475 2260 28515 2265
rect 28585 2295 28625 2300
rect 28585 2265 28590 2295
rect 28620 2265 28625 2295
rect 28585 2260 28625 2265
rect 28695 2295 28735 2300
rect 28695 2265 28700 2295
rect 28730 2265 28735 2295
rect 28695 2260 28735 2265
rect 28895 2295 28935 2300
rect 28895 2265 28900 2295
rect 28930 2265 28935 2295
rect 28895 2260 28935 2265
rect 28905 1930 28925 2260
rect 28950 1985 28970 2450
rect 29405 2120 29425 2800
rect 29390 2110 29440 2120
rect 29390 2080 29400 2110
rect 29430 2080 29440 2110
rect 29390 2070 29440 2080
rect 29065 1985 29100 1990
rect 28940 1980 28980 1985
rect 28940 1950 28945 1980
rect 28975 1950 28980 1980
rect 28940 1945 28980 1950
rect 29065 1945 29100 1950
rect 29125 1985 29160 1991
rect 29125 1945 29160 1950
rect 29185 1985 29220 1990
rect 29185 1945 29220 1950
rect 29245 1985 29280 1991
rect 29245 1945 29280 1950
rect 29130 1930 29150 1945
rect 28200 1925 28240 1930
rect 28200 1895 28205 1925
rect 28235 1895 28240 1925
rect 28200 1890 28240 1895
rect 28310 1925 28350 1930
rect 28310 1895 28315 1925
rect 28345 1895 28350 1925
rect 28310 1890 28350 1895
rect 28420 1925 28460 1930
rect 28420 1895 28425 1925
rect 28455 1895 28460 1925
rect 28420 1890 28460 1895
rect 28530 1925 28570 1930
rect 28530 1895 28535 1925
rect 28565 1895 28570 1925
rect 28530 1890 28570 1895
rect 28640 1925 28680 1930
rect 28640 1895 28645 1925
rect 28675 1895 28680 1925
rect 28640 1890 28680 1895
rect 28750 1925 28790 1930
rect 28750 1895 28755 1925
rect 28785 1895 28790 1925
rect 28750 1890 28790 1895
rect 28895 1925 28935 1930
rect 28895 1895 28900 1925
rect 28930 1895 28935 1925
rect 28895 1890 28935 1895
rect 29120 1925 29160 1930
rect 29120 1895 29125 1925
rect 29155 1895 29160 1925
rect 29120 1890 29160 1895
rect 29250 1880 29270 1945
rect 29240 1875 29280 1880
rect 29240 1845 29245 1875
rect 29275 1845 29280 1875
rect 29240 1840 29280 1845
rect 28025 1760 28065 1765
rect 28025 1730 28030 1760
rect 28060 1730 28065 1760
rect 28025 1725 28065 1730
rect 28405 1760 28445 1765
rect 28405 1730 28410 1760
rect 28440 1730 28445 1760
rect 28405 1725 28445 1730
rect 29115 1760 29155 1765
rect 29115 1730 29120 1760
rect 29150 1730 29155 1760
rect 29115 1725 29155 1730
rect 28035 1395 28055 1725
rect 28415 1710 28435 1725
rect 28305 1705 28345 1710
rect 28305 1675 28310 1705
rect 28340 1675 28345 1705
rect 28305 1670 28345 1675
rect 28408 1700 28442 1710
rect 28408 1680 28416 1700
rect 28434 1680 28442 1700
rect 28408 1670 28442 1680
rect 28505 1705 28545 1710
rect 28505 1675 28510 1705
rect 28540 1675 28545 1705
rect 28505 1670 28545 1675
rect 28705 1705 28745 1710
rect 28705 1675 28710 1705
rect 28740 1675 28745 1705
rect 28705 1670 28745 1675
rect 29050 1705 29090 1710
rect 29050 1675 29055 1705
rect 29085 1675 29090 1705
rect 29050 1670 29090 1675
rect 29060 1650 29080 1670
rect 29125 1650 29145 1725
rect 29405 1710 29425 2070
rect 29395 1705 29435 1710
rect 29395 1675 29400 1705
rect 29430 1675 29435 1705
rect 29395 1670 29435 1675
rect 29055 1645 29090 1650
rect 29055 1605 29090 1610
rect 29115 1645 29150 1650
rect 29115 1605 29150 1610
rect 28025 1390 28065 1395
rect 28025 1360 28030 1390
rect 28060 1360 28065 1390
rect 28025 1355 28065 1360
rect 28405 935 28445 940
rect 28405 905 28410 935
rect 28440 905 28445 935
rect 28405 900 28445 905
rect 28605 935 28645 940
rect 28605 905 28610 935
rect 28640 905 28645 935
rect 28605 900 28645 905
rect 27970 660 28010 665
rect 27970 630 27975 660
rect 28005 630 28010 660
rect 27970 625 28010 630
rect 25800 600 25840 605
rect 25800 570 25805 600
rect 25835 570 25840 600
rect 25800 565 25840 570
rect 26305 600 26345 605
rect 26305 570 26310 600
rect 26340 570 26345 600
rect 26305 565 26345 570
rect 26375 600 26415 605
rect 26375 570 26380 600
rect 26410 570 26415 600
rect 26375 565 26415 570
rect 26445 600 26485 605
rect 26445 570 26450 600
rect 26480 570 26485 600
rect 26445 565 26485 570
rect 26505 595 26545 605
rect 26505 575 26515 595
rect 26535 575 26545 595
rect 26505 565 26545 575
rect 26935 595 26975 605
rect 26935 575 26945 595
rect 26965 575 26975 595
rect 26935 565 26975 575
rect 27045 600 27085 605
rect 27045 570 27050 600
rect 27080 570 27085 600
rect 27045 565 27085 570
rect 27155 595 27195 605
rect 27155 575 27165 595
rect 27185 575 27195 595
rect 27155 565 27195 575
rect 27265 600 27305 605
rect 27265 570 27270 600
rect 27300 570 27305 600
rect 27265 565 27305 570
rect 27375 595 27415 605
rect 27375 575 27385 595
rect 27405 575 27415 595
rect 27375 565 27415 575
rect 27485 600 27525 605
rect 27485 570 27490 600
rect 27520 570 27525 600
rect 27485 565 27525 570
rect 27915 600 27955 605
rect 27915 570 27920 600
rect 27950 570 27955 600
rect 27915 565 27955 570
rect 26990 480 27030 485
rect 26990 450 26995 480
rect 27025 450 27030 480
rect 26990 445 27030 450
rect 27100 480 27140 485
rect 27100 450 27105 480
rect 27135 450 27140 480
rect 27100 445 27140 450
rect 27210 480 27250 485
rect 27210 450 27215 480
rect 27245 450 27250 480
rect 27210 445 27250 450
rect 27320 480 27360 485
rect 27320 450 27325 480
rect 27355 450 27360 480
rect 27320 445 27360 450
rect 27430 480 27470 485
rect 27430 450 27435 480
rect 27465 450 27470 480
rect 27430 445 27470 450
<< via1 >>
rect 26570 4955 26600 4985
rect 26690 4955 26720 4985
rect 26810 4955 26840 4985
rect 27240 4940 27270 4970
rect 26510 4920 26540 4925
rect 26510 4900 26515 4920
rect 26515 4900 26535 4920
rect 26535 4900 26540 4920
rect 26510 4895 26540 4900
rect 26630 4920 26660 4925
rect 26630 4900 26635 4920
rect 26635 4900 26655 4920
rect 26655 4900 26660 4920
rect 26630 4895 26660 4900
rect 26750 4920 26780 4925
rect 26750 4900 26755 4920
rect 26755 4900 26775 4920
rect 26775 4900 26780 4920
rect 26750 4895 26780 4900
rect 26870 4920 26900 4925
rect 26870 4900 26875 4920
rect 26875 4900 26895 4920
rect 26895 4900 26900 4920
rect 26870 4895 26900 4900
rect 27240 4895 27270 4900
rect 27240 4875 27245 4895
rect 27245 4875 27265 4895
rect 27265 4875 27270 4895
rect 27240 4870 27270 4875
rect 27360 4895 27390 4900
rect 27360 4875 27365 4895
rect 27365 4875 27385 4895
rect 27385 4875 27390 4895
rect 27360 4870 27390 4875
rect 27480 4895 27510 4900
rect 27480 4875 27485 4895
rect 27485 4875 27505 4895
rect 27505 4875 27510 4895
rect 27480 4870 27510 4875
rect 27600 4895 27630 4900
rect 27600 4875 27605 4895
rect 27605 4875 27625 4895
rect 27625 4875 27630 4895
rect 27600 4870 27630 4875
rect 27720 4895 27750 4900
rect 27720 4875 27725 4895
rect 27725 4875 27745 4895
rect 27745 4875 27750 4895
rect 27720 4870 27750 4875
rect 26055 4740 26085 4770
rect 26690 4765 26720 4770
rect 26690 4745 26695 4765
rect 26695 4745 26715 4765
rect 26715 4745 26720 4765
rect 26690 4740 26720 4745
rect 16600 4460 16630 4465
rect 16600 4440 16605 4460
rect 16605 4440 16625 4460
rect 16625 4440 16630 4460
rect 16600 4435 16630 4440
rect 16720 4460 16750 4465
rect 16720 4440 16725 4460
rect 16725 4440 16745 4460
rect 16745 4440 16750 4460
rect 16720 4435 16750 4440
rect 16840 4460 16870 4465
rect 16840 4440 16845 4460
rect 16845 4440 16865 4460
rect 16865 4440 16870 4460
rect 16840 4435 16870 4440
rect 17190 4435 17220 4465
rect 16170 4400 16200 4405
rect 16170 4380 16175 4400
rect 16175 4380 16195 4400
rect 16195 4380 16200 4400
rect 16170 4375 16200 4380
rect 16430 4400 16460 4405
rect 16430 4380 16435 4400
rect 16435 4380 16455 4400
rect 16455 4380 16460 4400
rect 16430 4375 16460 4380
rect 16540 4415 16570 4420
rect 16540 4395 16545 4415
rect 16545 4395 16565 4415
rect 16565 4395 16570 4415
rect 16540 4390 16570 4395
rect 16660 4415 16690 4420
rect 16660 4395 16665 4415
rect 16665 4395 16685 4415
rect 16685 4395 16690 4415
rect 16660 4390 16690 4395
rect 16780 4415 16810 4420
rect 16780 4395 16785 4415
rect 16785 4395 16805 4415
rect 16805 4395 16810 4415
rect 16780 4390 16810 4395
rect 16900 4415 16930 4420
rect 16900 4395 16905 4415
rect 16905 4395 16925 4415
rect 16925 4395 16930 4415
rect 16900 4390 16930 4395
rect 17190 4390 17220 4395
rect 17190 4370 17195 4390
rect 17195 4370 17215 4390
rect 17215 4370 17220 4390
rect 17190 4365 17220 4370
rect 17310 4390 17340 4395
rect 17310 4370 17315 4390
rect 17315 4370 17335 4390
rect 17335 4370 17340 4390
rect 17310 4365 17340 4370
rect 17430 4390 17460 4395
rect 17430 4370 17435 4390
rect 17435 4370 17455 4390
rect 17455 4370 17460 4390
rect 17430 4365 17460 4370
rect 17550 4390 17580 4395
rect 17550 4370 17555 4390
rect 17555 4370 17575 4390
rect 17575 4370 17580 4390
rect 17550 4365 17580 4370
rect 17670 4390 17700 4395
rect 17670 4370 17675 4390
rect 17675 4370 17695 4390
rect 17695 4370 17700 4390
rect 17670 4365 17700 4370
rect 16055 4235 16085 4265
rect 16720 4260 16750 4265
rect 16720 4240 16725 4260
rect 16725 4240 16745 4260
rect 16745 4240 16750 4260
rect 16720 4235 16750 4240
rect 14610 3605 14640 3635
rect 15065 3630 15095 3635
rect 15065 3610 15070 3630
rect 15070 3610 15090 3630
rect 15090 3610 15095 3630
rect 15065 3605 15095 3610
rect 15175 3630 15205 3635
rect 15175 3610 15180 3630
rect 15180 3610 15200 3630
rect 15200 3610 15205 3630
rect 15175 3605 15205 3610
rect 15285 3630 15315 3635
rect 15285 3610 15290 3630
rect 15290 3610 15310 3630
rect 15310 3610 15315 3630
rect 15285 3605 15315 3610
rect 15395 3630 15425 3635
rect 15395 3610 15400 3630
rect 15400 3610 15420 3630
rect 15420 3610 15425 3630
rect 15395 3605 15425 3610
rect 15505 3630 15535 3635
rect 15505 3610 15510 3630
rect 15510 3610 15530 3630
rect 15530 3610 15535 3630
rect 15505 3605 15535 3610
rect 15615 3630 15645 3635
rect 15615 3610 15620 3630
rect 15620 3610 15640 3630
rect 15640 3610 15645 3630
rect 15615 3605 15645 3610
rect 1266 3495 1296 3525
rect 14560 3525 14590 3555
rect 14610 3525 14640 3555
rect 14660 3525 14690 3555
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1210 3310 1240 3340
rect 1165 3255 1195 3285
rect 51 3200 86 3205
rect 51 3175 56 3200
rect 56 3175 81 3200
rect 81 3175 86 3200
rect 51 3170 86 3175
rect 51 3140 86 3145
rect 51 3115 56 3140
rect 56 3115 81 3140
rect 81 3115 86 3140
rect 51 3110 86 3115
rect 1165 3070 1195 3100
rect 51 3060 86 3065
rect 51 3035 56 3060
rect 56 3035 81 3060
rect 81 3035 86 3060
rect 51 3030 86 3035
rect 51 3000 86 3005
rect 51 2975 56 3000
rect 56 2975 81 3000
rect 81 2975 86 3000
rect 51 2970 86 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1266 3195 1301 3200
rect 1266 3170 1271 3195
rect 1271 3170 1296 3195
rect 1296 3170 1301 3195
rect 1266 3165 1301 3170
rect 1266 3135 1301 3140
rect 1266 3110 1271 3135
rect 1271 3110 1296 3135
rect 1296 3110 1301 3135
rect 1266 3105 1301 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 56 2850 91 2855
rect 56 2825 61 2850
rect 61 2825 86 2850
rect 86 2825 91 2850
rect 56 2820 91 2825
rect 729 2850 764 2855
rect 729 2825 734 2850
rect 734 2825 759 2850
rect 759 2825 764 2850
rect 729 2820 764 2825
rect 1210 2820 1240 2850
rect 1266 2835 1301 2840
rect 1266 2810 1271 2835
rect 1271 2810 1296 2835
rect 1296 2810 1301 2835
rect 1266 2805 1301 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 56 2790 91 2795
rect 56 2765 61 2790
rect 61 2765 86 2790
rect 86 2765 91 2790
rect 56 2760 91 2765
rect 729 2790 764 2795
rect 729 2765 734 2790
rect 734 2765 759 2790
rect 759 2765 764 2790
rect 729 2760 764 2765
rect 1266 2715 1296 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5365 3305 5395 3335
rect 4890 3255 4920 3285
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 3990 3050 4020 3080
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 5320 3110 5350 3140
rect 3085 2975 3115 2980
rect 3085 2955 3090 2975
rect 3090 2955 3110 2975
rect 3110 2955 3115 2975
rect 3085 2950 3115 2955
rect 3270 2975 3300 2980
rect 3270 2955 3275 2975
rect 3275 2955 3295 2975
rect 3295 2955 3300 2975
rect 3270 2950 3300 2955
rect 3630 2975 3660 2980
rect 3630 2955 3635 2975
rect 3635 2955 3655 2975
rect 3655 2955 3660 2975
rect 3630 2950 3660 2955
rect 4170 2975 4200 2980
rect 4170 2955 4175 2975
rect 4175 2955 4195 2975
rect 4195 2955 4200 2975
rect 4170 2950 4200 2955
rect 4530 2975 4560 2980
rect 4530 2955 4535 2975
rect 4535 2955 4555 2975
rect 4555 2955 4560 2975
rect 4530 2950 4560 2955
rect 3000 2805 3030 2810
rect 3000 2785 3005 2805
rect 3005 2785 3025 2805
rect 3025 2785 3030 2805
rect 3000 2780 3030 2785
rect 3180 2805 3210 2810
rect 3180 2785 3185 2805
rect 3185 2785 3205 2805
rect 3205 2785 3210 2805
rect 3180 2780 3210 2785
rect 3360 2805 3390 2810
rect 3360 2785 3365 2805
rect 3365 2785 3385 2805
rect 3385 2785 3390 2805
rect 3360 2780 3390 2785
rect 3540 2805 3570 2810
rect 3540 2785 3545 2805
rect 3545 2785 3565 2805
rect 3565 2785 3570 2805
rect 3540 2780 3570 2785
rect 3720 2805 3750 2810
rect 3720 2785 3725 2805
rect 3725 2785 3745 2805
rect 3745 2785 3750 2805
rect 3720 2780 3750 2785
rect 3900 2805 3930 2810
rect 3900 2785 3905 2805
rect 3905 2785 3925 2805
rect 3925 2785 3930 2805
rect 3900 2780 3930 2785
rect 4080 2805 4110 2810
rect 4080 2785 4085 2805
rect 4085 2785 4105 2805
rect 4105 2785 4110 2805
rect 4080 2780 4110 2785
rect 4260 2805 4290 2810
rect 4260 2785 4265 2805
rect 4265 2785 4285 2805
rect 4285 2785 4290 2805
rect 4260 2780 4290 2785
rect 4440 2805 4470 2810
rect 4440 2785 4445 2805
rect 4445 2785 4465 2805
rect 4465 2785 4470 2805
rect 4440 2780 4470 2785
rect 4620 2805 4650 2810
rect 4620 2785 4625 2805
rect 4625 2785 4645 2805
rect 4645 2785 4650 2805
rect 4620 2780 4650 2785
rect 4800 2805 4830 2810
rect 4800 2785 4805 2805
rect 4805 2785 4825 2805
rect 4825 2785 4830 2805
rect 4800 2780 4830 2785
rect 4980 2805 5010 2810
rect 4980 2785 4985 2805
rect 4985 2785 5005 2805
rect 5005 2785 5010 2805
rect 4980 2780 5010 2785
rect 3180 2745 3210 2750
rect 3180 2725 3185 2745
rect 3185 2725 3205 2745
rect 3205 2725 3210 2745
rect 3180 2720 3210 2725
rect 3360 2745 3390 2750
rect 3360 2725 3365 2745
rect 3365 2725 3385 2745
rect 3385 2725 3390 2745
rect 3360 2720 3390 2725
rect 3540 2745 3570 2750
rect 3540 2725 3545 2745
rect 3545 2725 3565 2745
rect 3565 2725 3570 2745
rect 3540 2720 3570 2725
rect 3720 2745 3750 2750
rect 3720 2725 3725 2745
rect 3725 2725 3745 2745
rect 3745 2725 3750 2745
rect 3720 2720 3750 2725
rect 3900 2745 3930 2750
rect 3900 2725 3905 2745
rect 3905 2725 3925 2745
rect 3925 2725 3930 2745
rect 3900 2720 3930 2725
rect 4080 2745 4110 2750
rect 4080 2725 4085 2745
rect 4085 2725 4105 2745
rect 4105 2725 4110 2745
rect 4080 2720 4110 2725
rect 4260 2745 4290 2750
rect 4260 2725 4265 2745
rect 4265 2725 4285 2745
rect 4285 2725 4290 2745
rect 4260 2720 4290 2725
rect 4440 2745 4470 2750
rect 4440 2725 4445 2745
rect 4445 2725 4465 2745
rect 4465 2725 4470 2745
rect 4440 2720 4470 2725
rect 4620 2745 4650 2750
rect 4620 2725 4625 2745
rect 4625 2725 4645 2745
rect 4645 2725 4650 2745
rect 4620 2720 4650 2725
rect 4800 2745 4830 2750
rect 4800 2725 4805 2745
rect 4805 2725 4825 2745
rect 4825 2725 4830 2745
rect 4800 2720 4830 2725
rect 3360 2370 3390 2375
rect 3360 2350 3365 2370
rect 3365 2350 3385 2370
rect 3385 2350 3390 2370
rect 3360 2345 3390 2350
rect 3810 2375 3840 2380
rect 3810 2355 3815 2375
rect 3815 2355 3835 2375
rect 3835 2355 3840 2375
rect 3810 2350 3840 2355
rect 4170 2375 4200 2380
rect 4170 2355 4175 2375
rect 4175 2355 4195 2375
rect 4195 2355 4200 2375
rect 4170 2350 4200 2355
rect 2740 2260 2770 2290
rect 3630 2330 3660 2335
rect 3630 2310 3635 2330
rect 3635 2310 3655 2330
rect 3655 2310 3660 2330
rect 3630 2305 3660 2310
rect 3450 2285 3480 2290
rect 3450 2265 3455 2285
rect 3455 2265 3475 2285
rect 3475 2265 3480 2285
rect 3450 2260 3480 2265
rect 3270 2170 3300 2200
rect 3810 2215 3840 2245
rect 3630 2120 3660 2150
rect 2750 2090 2780 2095
rect 2750 2070 2755 2090
rect 2755 2070 2775 2090
rect 2775 2070 2780 2090
rect 2750 2065 2780 2070
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4350 2330 4380 2335
rect 4350 2310 4355 2330
rect 4355 2310 4375 2330
rect 4375 2310 4380 2330
rect 4350 2305 4380 2310
rect 4530 2285 4560 2290
rect 4530 2265 4535 2285
rect 4535 2265 4555 2285
rect 4555 2265 4560 2285
rect 4530 2260 4560 2265
rect 5275 2260 5305 2290
rect 3990 2170 4020 2200
rect 4710 2170 4740 2200
rect 4090 2115 4120 2145
rect 3990 2090 4020 2095
rect 3990 2070 3995 2090
rect 3995 2070 4015 2090
rect 4015 2070 4020 2090
rect 3990 2065 4020 2070
rect 4150 2090 4180 2095
rect 4150 2070 4155 2090
rect 4155 2070 4175 2090
rect 4175 2070 4180 2090
rect 4150 2065 4180 2070
rect 4270 2090 4300 2095
rect 4270 2070 4275 2090
rect 4275 2070 4295 2090
rect 4295 2070 4300 2090
rect 4270 2065 4300 2070
rect 4390 2090 4420 2095
rect 4390 2070 4395 2090
rect 4395 2070 4415 2090
rect 4415 2070 4420 2090
rect 4390 2065 4420 2070
rect 4510 2090 4540 2095
rect 4510 2070 4515 2090
rect 4515 2070 4535 2090
rect 4535 2070 4540 2090
rect 4510 2065 4540 2070
rect 4630 2090 4660 2095
rect 4630 2070 4635 2090
rect 4635 2070 4655 2090
rect 4655 2070 4660 2090
rect 4630 2065 4660 2070
rect 4750 2090 4780 2095
rect 4750 2070 4755 2090
rect 4755 2070 4775 2090
rect 4775 2070 4780 2090
rect 4750 2065 4780 2070
rect 4870 2090 4900 2095
rect 4870 2070 4875 2090
rect 4875 2070 4895 2090
rect 4895 2070 4900 2090
rect 4870 2065 4900 2070
rect 4990 2090 5020 2095
rect 4990 2070 4995 2090
rect 4995 2070 5015 2090
rect 5015 2070 5020 2090
rect 4990 2065 5020 2070
rect 5110 2090 5140 2095
rect 5110 2070 5115 2090
rect 5115 2070 5135 2090
rect 5135 2070 5140 2090
rect 5110 2065 5140 2070
rect 5230 2090 5260 2095
rect 5230 2070 5235 2090
rect 5235 2070 5255 2090
rect 5255 2070 5260 2090
rect 5230 2065 5260 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 4090 2045 4120 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 2805 1680 2835 1710
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 2930 1495 2960 1500
rect 2930 1475 2935 1495
rect 2935 1475 2955 1495
rect 2955 1475 2960 1495
rect 2930 1470 2960 1475
rect 3050 1495 3080 1500
rect 3050 1475 3055 1495
rect 3055 1475 3075 1495
rect 3075 1475 3080 1495
rect 3050 1470 3080 1475
rect 3170 1495 3200 1500
rect 3170 1475 3175 1495
rect 3175 1475 3195 1495
rect 3195 1475 3200 1495
rect 3170 1470 3200 1475
rect 3290 1495 3320 1500
rect 3290 1475 3295 1495
rect 3295 1475 3315 1495
rect 3315 1475 3320 1495
rect 3290 1470 3320 1475
rect 3530 1495 3560 1500
rect 3530 1475 3535 1495
rect 3535 1475 3555 1495
rect 3555 1475 3560 1495
rect 3530 1470 3560 1475
rect 3650 1495 3680 1500
rect 3650 1475 3655 1495
rect 3655 1475 3675 1495
rect 3675 1475 3680 1495
rect 3650 1470 3680 1475
rect 3770 1495 3800 1500
rect 3770 1475 3775 1495
rect 3775 1475 3795 1495
rect 3795 1475 3800 1495
rect 3770 1470 3800 1475
rect 4090 2025 4095 2045
rect 4095 2025 4115 2045
rect 4115 2025 4120 2045
rect 4090 2020 4120 2025
rect 4450 2045 4480 2050
rect 4450 2025 4455 2045
rect 4455 2025 4475 2045
rect 4475 2025 4480 2045
rect 4450 2020 4480 2025
rect 4810 2045 4840 2050
rect 4810 2025 4815 2045
rect 4815 2025 4835 2045
rect 4835 2025 4840 2045
rect 4810 2020 4840 2025
rect 5170 2045 5200 2050
rect 5170 2025 5175 2045
rect 5175 2025 5195 2045
rect 5195 2025 5200 2045
rect 5170 2020 5200 2025
rect 4330 1875 4360 1880
rect 4330 1855 4335 1875
rect 4335 1855 4355 1875
rect 4355 1855 4360 1875
rect 4330 1850 4360 1855
rect 4690 1875 4720 1880
rect 4690 1855 4695 1875
rect 4695 1855 4715 1875
rect 4715 1855 4720 1875
rect 4690 1850 4720 1855
rect 5050 1875 5080 1880
rect 5050 1855 5055 1875
rect 5055 1855 5075 1875
rect 5075 1855 5080 1875
rect 5050 1850 5080 1855
rect 4120 1790 4150 1820
rect 4210 1815 4240 1820
rect 4210 1795 4215 1815
rect 4215 1795 4235 1815
rect 4235 1795 4240 1815
rect 4210 1790 4240 1795
rect 4450 1790 4480 1820
rect 4570 1815 4600 1820
rect 4570 1795 4575 1815
rect 4575 1795 4595 1815
rect 4595 1795 4600 1815
rect 4570 1790 4600 1795
rect 4210 1755 4240 1760
rect 4210 1735 4215 1755
rect 4215 1735 4235 1755
rect 4235 1735 4240 1755
rect 4210 1730 4240 1735
rect 4450 1755 4480 1760
rect 4450 1735 4455 1755
rect 4455 1735 4475 1755
rect 4475 1735 4480 1755
rect 4450 1730 4480 1735
rect 4810 1790 4840 1820
rect 4930 1815 4960 1820
rect 4930 1795 4935 1815
rect 4935 1795 4955 1815
rect 4955 1795 4960 1815
rect 4930 1790 4960 1795
rect 5140 1790 5170 1820
rect 5320 2115 5350 2145
rect 5415 3255 5445 3285
rect 5365 1790 5395 1820
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 4750 1755 4780 1760
rect 4750 1735 4755 1755
rect 4755 1735 4775 1755
rect 4775 1735 4780 1755
rect 4750 1730 4780 1735
rect 5275 1730 5305 1760
rect 4330 1710 4360 1715
rect 4330 1690 4335 1710
rect 4335 1690 4355 1710
rect 4355 1690 4360 1710
rect 4330 1685 4360 1690
rect 4570 1710 4600 1715
rect 4570 1690 4575 1710
rect 4575 1690 4595 1710
rect 4595 1690 4600 1710
rect 4570 1685 4600 1690
rect 4810 1710 4840 1715
rect 4810 1690 4815 1710
rect 4815 1690 4835 1710
rect 4835 1690 4840 1710
rect 4810 1685 4840 1690
rect 17250 4260 17280 4265
rect 17250 4240 17255 4260
rect 17255 4240 17275 4260
rect 17275 4240 17280 4260
rect 17250 4235 17280 4240
rect 17370 4260 17400 4265
rect 17370 4240 17375 4260
rect 17375 4240 17395 4260
rect 17395 4240 17400 4260
rect 17370 4235 17400 4240
rect 17490 4260 17520 4265
rect 17490 4240 17495 4260
rect 17495 4240 17515 4260
rect 17515 4240 17520 4260
rect 17490 4235 17520 4240
rect 17610 4260 17640 4265
rect 17610 4240 17615 4260
rect 17615 4240 17635 4260
rect 17635 4240 17640 4260
rect 17610 4235 17640 4240
rect 16110 4180 16140 4210
rect 16300 4180 16330 4210
rect 17310 4180 17340 4210
rect 16055 3075 16085 3105
rect 14560 2905 14590 2935
rect 14610 2905 14640 2935
rect 14660 2905 14690 2935
rect 15120 2960 15150 2965
rect 15120 2940 15125 2960
rect 15125 2940 15145 2960
rect 15145 2940 15150 2960
rect 15120 2935 15150 2940
rect 15230 2960 15260 2965
rect 15230 2940 15235 2960
rect 15235 2940 15255 2960
rect 15255 2940 15260 2960
rect 15230 2935 15260 2940
rect 15340 2960 15370 2965
rect 15340 2940 15345 2960
rect 15345 2940 15365 2960
rect 15365 2940 15370 2960
rect 15340 2935 15370 2940
rect 15450 2960 15480 2965
rect 15450 2940 15455 2960
rect 15455 2940 15475 2960
rect 15475 2940 15480 2960
rect 15450 2935 15480 2940
rect 15560 2960 15590 2965
rect 15560 2940 15565 2960
rect 15565 2940 15585 2960
rect 15585 2940 15590 2960
rect 15560 2935 15590 2940
rect 16365 4150 16395 4155
rect 16365 4130 16370 4150
rect 16370 4130 16390 4150
rect 16390 4130 16395 4150
rect 16365 4125 16395 4130
rect 16475 4150 16505 4155
rect 16475 4130 16480 4150
rect 16480 4130 16500 4150
rect 16500 4130 16505 4150
rect 16475 4125 16505 4130
rect 16585 4150 16615 4155
rect 16585 4130 16590 4150
rect 16590 4130 16610 4150
rect 16610 4130 16615 4150
rect 16585 4125 16615 4130
rect 16695 4150 16725 4155
rect 16695 4130 16700 4150
rect 16700 4130 16720 4150
rect 16720 4130 16725 4150
rect 16695 4125 16725 4130
rect 16805 4150 16835 4155
rect 16805 4130 16810 4150
rect 16810 4130 16830 4150
rect 16830 4130 16835 4150
rect 16805 4125 16835 4130
rect 16915 4150 16945 4155
rect 16915 4130 16920 4150
rect 16920 4130 16940 4150
rect 16940 4130 16945 4150
rect 16915 4125 16945 4130
rect 17025 4150 17055 4155
rect 17025 4130 17030 4150
rect 17030 4130 17050 4150
rect 17050 4130 17055 4150
rect 17025 4125 17055 4130
rect 17135 4150 17165 4155
rect 17135 4130 17140 4150
rect 17140 4130 17160 4150
rect 17160 4130 17165 4150
rect 17135 4125 17165 4130
rect 17245 4150 17275 4155
rect 17245 4130 17250 4150
rect 17250 4130 17270 4150
rect 17270 4130 17275 4150
rect 17245 4125 17275 4130
rect 17355 4150 17385 4155
rect 17355 4130 17360 4150
rect 17360 4130 17380 4150
rect 17380 4130 17385 4150
rect 17355 4125 17385 4130
rect 16310 4030 16340 4035
rect 16310 4010 16315 4030
rect 16315 4010 16335 4030
rect 16335 4010 16340 4030
rect 16310 4005 16340 4010
rect 16530 4030 16560 4035
rect 16530 4010 16535 4030
rect 16535 4010 16555 4030
rect 16555 4010 16560 4030
rect 16530 4005 16560 4010
rect 16750 4030 16780 4035
rect 16750 4010 16755 4030
rect 16755 4010 16775 4030
rect 16775 4010 16780 4030
rect 16750 4005 16780 4010
rect 16970 4030 17000 4035
rect 16970 4010 16975 4030
rect 16975 4010 16995 4030
rect 16995 4010 17000 4030
rect 16970 4005 17000 4010
rect 17190 4030 17220 4035
rect 17190 4010 17195 4030
rect 17195 4010 17215 4030
rect 17215 4010 17220 4030
rect 17190 4005 17220 4010
rect 17410 4030 17440 4035
rect 17410 4010 17415 4030
rect 17415 4010 17435 4030
rect 17435 4010 17440 4030
rect 17410 4005 17440 4010
rect 16315 3905 16345 3910
rect 16315 3885 16320 3905
rect 16320 3885 16340 3905
rect 16340 3885 16345 3905
rect 16315 3880 16345 3885
rect 16420 3945 16450 3975
rect 16640 3945 16670 3975
rect 16860 3945 16890 3975
rect 17080 3945 17110 3975
rect 17300 3945 17330 3975
rect 16420 3905 16450 3910
rect 16420 3885 16425 3905
rect 16425 3885 16445 3905
rect 16445 3885 16450 3905
rect 16420 3880 16450 3885
rect 16530 3905 16560 3910
rect 16530 3885 16535 3905
rect 16535 3885 16555 3905
rect 16555 3885 16560 3905
rect 16530 3880 16560 3885
rect 16640 3905 16670 3910
rect 16640 3885 16645 3905
rect 16645 3885 16665 3905
rect 16665 3885 16670 3905
rect 16640 3880 16670 3885
rect 16750 3905 16780 3910
rect 16750 3885 16755 3905
rect 16755 3885 16775 3905
rect 16775 3885 16780 3905
rect 16750 3880 16780 3885
rect 17055 3905 17085 3910
rect 17055 3885 17060 3905
rect 17060 3885 17080 3905
rect 17080 3885 17085 3905
rect 17055 3880 17085 3885
rect 17160 3905 17190 3910
rect 17160 3885 17165 3905
rect 17165 3885 17185 3905
rect 17185 3885 17190 3905
rect 17160 3880 17190 3885
rect 17270 3905 17300 3910
rect 17270 3885 17275 3905
rect 17275 3885 17295 3905
rect 17295 3885 17300 3905
rect 17270 3880 17300 3885
rect 17380 3905 17410 3910
rect 17380 3885 17385 3905
rect 17385 3885 17405 3905
rect 17405 3885 17410 3905
rect 17380 3880 17410 3885
rect 17490 3905 17520 3910
rect 17490 3885 17495 3905
rect 17495 3885 17515 3905
rect 17515 3885 17520 3905
rect 17490 3880 17520 3885
rect 16274 3845 16300 3850
rect 16274 3825 16277 3845
rect 16277 3825 16294 3845
rect 16294 3825 16300 3845
rect 16274 3820 16300 3825
rect 16475 3845 16505 3850
rect 16475 3825 16480 3845
rect 16480 3825 16500 3845
rect 16500 3825 16505 3845
rect 16475 3820 16505 3825
rect 16695 3845 16725 3850
rect 16695 3825 16700 3845
rect 16700 3825 16720 3845
rect 16720 3825 16725 3845
rect 16695 3820 16725 3825
rect 17014 3845 17040 3850
rect 17014 3825 17017 3845
rect 17017 3825 17034 3845
rect 17034 3825 17040 3845
rect 17014 3820 17040 3825
rect 17215 3845 17245 3850
rect 17215 3825 17220 3845
rect 17220 3825 17240 3845
rect 17240 3825 17245 3845
rect 17215 3820 17245 3825
rect 17435 3845 17465 3850
rect 17435 3825 17440 3845
rect 17440 3825 17460 3845
rect 17460 3825 17465 3845
rect 17435 3820 17465 3825
rect 17865 3820 17895 3850
rect 16405 3725 16431 3730
rect 16405 3705 16408 3725
rect 16408 3705 16425 3725
rect 16425 3705 16431 3725
rect 16405 3700 16431 3705
rect 16625 3725 16651 3730
rect 16625 3705 16628 3725
rect 16628 3705 16645 3725
rect 16645 3705 16651 3725
rect 16625 3700 16651 3705
rect 16769 3725 16795 3730
rect 16769 3705 16775 3725
rect 16775 3705 16792 3725
rect 16792 3705 16795 3725
rect 16769 3700 16795 3705
rect 17145 3725 17171 3730
rect 17145 3705 17148 3725
rect 17148 3705 17165 3725
rect 17165 3705 17171 3725
rect 17145 3700 17171 3705
rect 17365 3725 17391 3730
rect 17365 3705 17368 3725
rect 17368 3705 17385 3725
rect 17385 3705 17391 3725
rect 17365 3700 17391 3705
rect 17509 3725 17535 3730
rect 17509 3705 17515 3725
rect 17515 3705 17532 3725
rect 17532 3705 17535 3725
rect 17509 3700 17535 3705
rect 16255 3665 16285 3670
rect 16255 3645 16260 3665
rect 16260 3645 16280 3665
rect 16280 3645 16285 3665
rect 16255 3640 16285 3645
rect 16360 3665 16390 3670
rect 16360 3645 16365 3665
rect 16365 3645 16385 3665
rect 16385 3645 16390 3665
rect 16360 3640 16390 3645
rect 16475 3665 16505 3670
rect 16475 3645 16480 3665
rect 16480 3645 16500 3665
rect 16500 3645 16505 3665
rect 16475 3640 16505 3645
rect 16580 3665 16610 3670
rect 16580 3645 16585 3665
rect 16585 3645 16605 3665
rect 16605 3645 16610 3665
rect 16580 3640 16610 3645
rect 16695 3665 16725 3670
rect 16695 3645 16700 3665
rect 16700 3645 16720 3665
rect 16720 3645 16725 3665
rect 16695 3640 16725 3645
rect 16810 3665 16840 3670
rect 16810 3645 16815 3665
rect 16815 3645 16835 3665
rect 16835 3645 16840 3665
rect 16810 3640 16840 3645
rect 16995 3675 17025 3680
rect 16995 3655 17000 3675
rect 17000 3655 17020 3675
rect 17020 3655 17025 3675
rect 16995 3650 17025 3655
rect 17215 3675 17245 3680
rect 17215 3655 17220 3675
rect 17220 3655 17240 3675
rect 17240 3655 17245 3675
rect 17215 3650 17245 3655
rect 17435 3675 17465 3680
rect 17435 3655 17440 3675
rect 17440 3655 17460 3675
rect 17460 3655 17465 3675
rect 17435 3650 17465 3655
rect 17100 3605 17130 3635
rect 17320 3605 17350 3635
rect 17550 3605 17580 3635
rect 16345 3570 16375 3575
rect 16345 3550 16350 3570
rect 16350 3550 16370 3570
rect 16370 3550 16375 3570
rect 16345 3545 16375 3550
rect 16465 3570 16495 3575
rect 16465 3550 16470 3570
rect 16470 3550 16490 3570
rect 16490 3550 16495 3570
rect 16465 3545 16495 3550
rect 16585 3570 16615 3575
rect 16585 3550 16590 3570
rect 16590 3550 16610 3570
rect 16610 3550 16615 3570
rect 16585 3545 16615 3550
rect 16705 3570 16735 3575
rect 16705 3550 16710 3570
rect 16710 3550 16730 3570
rect 16730 3550 16735 3570
rect 16705 3545 16735 3550
rect 16825 3570 16855 3575
rect 16825 3550 16830 3570
rect 16830 3550 16850 3570
rect 16850 3550 16855 3570
rect 16825 3545 16855 3550
rect 16945 3570 16975 3575
rect 16945 3550 16950 3570
rect 16950 3550 16970 3570
rect 16970 3550 16975 3570
rect 16945 3545 16975 3550
rect 17065 3570 17095 3575
rect 17065 3550 17070 3570
rect 17070 3550 17090 3570
rect 17090 3550 17095 3570
rect 17065 3545 17095 3550
rect 17185 3570 17215 3575
rect 17185 3550 17190 3570
rect 17190 3550 17210 3570
rect 17210 3550 17215 3570
rect 17185 3545 17215 3550
rect 17305 3570 17335 3575
rect 17305 3550 17310 3570
rect 17310 3550 17330 3570
rect 17330 3550 17335 3570
rect 17305 3545 17335 3550
rect 17425 3570 17455 3575
rect 17425 3550 17430 3570
rect 17430 3550 17450 3570
rect 17450 3550 17455 3570
rect 17425 3545 17455 3550
rect 16826 3100 16854 3105
rect 16826 3080 16831 3100
rect 16831 3080 16849 3100
rect 16849 3080 16854 3100
rect 16826 3075 16854 3080
rect 16285 3020 16315 3050
rect 16525 3020 16555 3050
rect 16765 3020 16795 3050
rect 17005 3020 17035 3050
rect 17245 3020 17275 3050
rect 17485 3020 17515 3050
rect 16405 2975 16435 3005
rect 16645 2975 16675 3005
rect 16885 2975 16915 3005
rect 17125 2975 17155 3005
rect 17365 2975 17395 3005
rect 14610 2850 14640 2880
rect 16110 2920 16140 2950
rect 16885 2920 16915 2950
rect 15505 2850 15535 2880
rect 15785 2850 15815 2880
rect 16140 2890 16170 2895
rect 16140 2870 16145 2890
rect 16145 2870 16165 2890
rect 16165 2870 16170 2890
rect 16140 2865 16170 2870
rect 16260 2890 16290 2895
rect 16260 2870 16265 2890
rect 16265 2870 16285 2890
rect 16285 2870 16290 2890
rect 16260 2865 16290 2870
rect 16380 2890 16410 2895
rect 16380 2870 16385 2890
rect 16385 2870 16405 2890
rect 16405 2870 16410 2890
rect 16380 2865 16410 2870
rect 16500 2890 16530 2895
rect 16500 2870 16505 2890
rect 16505 2870 16525 2890
rect 16525 2870 16530 2890
rect 16500 2865 16530 2870
rect 16620 2890 16650 2895
rect 16620 2870 16625 2890
rect 16625 2870 16645 2890
rect 16645 2870 16650 2890
rect 16620 2865 16650 2870
rect 14520 2795 14550 2825
rect 15230 2795 15260 2825
rect 15065 2700 15095 2705
rect 15065 2680 15070 2700
rect 15070 2680 15090 2700
rect 15090 2680 15095 2700
rect 15065 2675 15095 2680
rect 15175 2700 15205 2705
rect 15175 2680 15180 2700
rect 15180 2680 15200 2700
rect 15200 2680 15205 2700
rect 15175 2675 15205 2680
rect 15285 2700 15315 2705
rect 15285 2680 15290 2700
rect 15290 2680 15310 2700
rect 15310 2680 15315 2700
rect 15285 2675 15315 2680
rect 15395 2700 15425 2705
rect 15395 2680 15400 2700
rect 15400 2680 15420 2700
rect 15420 2680 15425 2700
rect 15395 2675 15425 2680
rect 15505 2700 15535 2705
rect 15505 2680 15510 2700
rect 15510 2680 15530 2700
rect 15530 2680 15535 2700
rect 15505 2675 15535 2680
rect 15615 2700 15645 2705
rect 15615 2680 15620 2700
rect 15620 2680 15640 2700
rect 15640 2680 15645 2700
rect 15615 2675 15645 2680
rect 14875 2405 14905 2435
rect 15120 2430 15150 2435
rect 15120 2410 15125 2430
rect 15125 2410 15145 2430
rect 15145 2410 15150 2430
rect 15120 2405 15150 2410
rect 15230 2430 15260 2435
rect 15230 2410 15235 2430
rect 15235 2410 15255 2430
rect 15255 2410 15260 2430
rect 15230 2405 15260 2410
rect 15340 2430 15370 2435
rect 15340 2410 15345 2430
rect 15345 2410 15365 2430
rect 15365 2410 15370 2430
rect 15340 2405 15370 2410
rect 15450 2430 15480 2435
rect 15450 2410 15455 2430
rect 15455 2410 15475 2430
rect 15475 2410 15480 2430
rect 15450 2405 15480 2410
rect 15560 2430 15590 2435
rect 15560 2410 15565 2430
rect 15565 2410 15585 2430
rect 15585 2410 15590 2430
rect 15560 2405 15590 2410
rect 14520 2080 14550 2110
rect 14640 2000 14675 2005
rect 14640 1975 14645 2000
rect 14645 1975 14670 2000
rect 14670 1975 14675 2000
rect 14640 1970 14675 1975
rect 14700 2000 14735 2005
rect 14700 1975 14705 2000
rect 14705 1975 14730 2000
rect 14730 1975 14735 2000
rect 14700 1970 14735 1975
rect 14760 2000 14795 2005
rect 14760 1975 14765 2000
rect 14765 1975 14790 2000
rect 14790 1975 14795 2000
rect 14760 1970 14795 1975
rect 16080 2470 16110 2475
rect 16080 2450 16085 2470
rect 16085 2450 16105 2470
rect 16105 2450 16110 2470
rect 16080 2445 16110 2450
rect 16200 2470 16230 2475
rect 16200 2450 16205 2470
rect 16205 2450 16225 2470
rect 16225 2450 16230 2470
rect 16200 2445 16230 2450
rect 16320 2470 16350 2475
rect 16320 2450 16325 2470
rect 16325 2450 16345 2470
rect 16345 2450 16350 2470
rect 16320 2445 16350 2450
rect 16440 2470 16470 2475
rect 16440 2450 16445 2470
rect 16445 2450 16465 2470
rect 16465 2450 16470 2470
rect 16440 2445 16470 2450
rect 16560 2470 16590 2475
rect 16560 2450 16565 2470
rect 16565 2450 16585 2470
rect 16585 2450 16590 2470
rect 16560 2445 16590 2450
rect 16680 2470 16710 2475
rect 16680 2450 16685 2470
rect 16685 2450 16705 2470
rect 16705 2450 16710 2470
rect 16680 2445 16710 2450
rect 17150 2890 17180 2895
rect 17150 2870 17155 2890
rect 17155 2870 17175 2890
rect 17175 2870 17180 2890
rect 17150 2865 17180 2870
rect 17270 2890 17300 2895
rect 17270 2870 17275 2890
rect 17275 2870 17295 2890
rect 17295 2870 17300 2890
rect 17270 2865 17300 2870
rect 17390 2890 17420 2895
rect 17390 2870 17395 2890
rect 17395 2870 17415 2890
rect 17415 2870 17420 2890
rect 17390 2865 17420 2870
rect 17510 2890 17540 2895
rect 17510 2870 17515 2890
rect 17515 2870 17535 2890
rect 17535 2870 17540 2890
rect 17510 2865 17540 2870
rect 17630 2890 17660 2895
rect 17630 2870 17635 2890
rect 17635 2870 17655 2890
rect 17655 2870 17660 2890
rect 17630 2865 17660 2870
rect 17090 2470 17120 2475
rect 17090 2450 17095 2470
rect 17095 2450 17115 2470
rect 17115 2450 17120 2470
rect 17090 2445 17120 2450
rect 17210 2470 17240 2475
rect 17210 2450 17215 2470
rect 17215 2450 17235 2470
rect 17235 2450 17240 2470
rect 17210 2445 17240 2450
rect 17330 2470 17360 2475
rect 17330 2450 17335 2470
rect 17335 2450 17355 2470
rect 17355 2450 17360 2470
rect 17330 2445 17360 2450
rect 17450 2470 17480 2475
rect 17450 2450 17455 2470
rect 17455 2450 17475 2470
rect 17475 2450 17480 2470
rect 17450 2445 17480 2450
rect 17570 2470 17600 2475
rect 17570 2450 17575 2470
rect 17575 2450 17595 2470
rect 17595 2450 17600 2470
rect 17570 2445 17600 2450
rect 17690 2470 17720 2475
rect 17690 2450 17695 2470
rect 17695 2450 17715 2470
rect 17715 2450 17720 2470
rect 17690 2445 17720 2450
rect 16380 2390 16410 2420
rect 16885 2390 16915 2420
rect 17390 2390 17420 2420
rect 15590 2370 15620 2375
rect 15590 2350 15595 2370
rect 15595 2350 15615 2370
rect 15615 2350 15620 2370
rect 15590 2345 15620 2350
rect 15785 2345 15815 2375
rect 16325 2345 16355 2375
rect 17325 2345 17355 2375
rect 14920 2285 14950 2315
rect 15120 2310 15150 2315
rect 15120 2290 15125 2310
rect 15125 2290 15145 2310
rect 15145 2290 15150 2310
rect 15120 2285 15150 2290
rect 15230 2310 15260 2315
rect 15230 2290 15235 2310
rect 15235 2290 15255 2310
rect 15255 2290 15260 2310
rect 15230 2285 15260 2290
rect 15340 2310 15370 2315
rect 15340 2290 15345 2310
rect 15345 2290 15365 2310
rect 15365 2290 15370 2310
rect 15340 2285 15370 2290
rect 15450 2310 15480 2315
rect 15450 2290 15455 2310
rect 15455 2290 15475 2310
rect 15475 2290 15480 2310
rect 15450 2285 15480 2290
rect 15560 2310 15590 2315
rect 15560 2290 15565 2310
rect 15565 2290 15585 2310
rect 15585 2290 15590 2310
rect 15560 2285 15590 2290
rect 16005 2295 16035 2325
rect 14820 2000 14855 2005
rect 14820 1975 14825 2000
rect 14825 1975 14850 2000
rect 14850 1975 14855 2000
rect 14820 1970 14855 1975
rect 14875 1970 14905 2000
rect 15805 2150 15835 2180
rect 14765 1915 14795 1945
rect 14920 1915 14950 1945
rect 15065 1940 15095 1945
rect 15065 1920 15070 1940
rect 15070 1920 15088 1940
rect 15088 1920 15095 1940
rect 15065 1915 15095 1920
rect 15175 1940 15205 1945
rect 15175 1920 15180 1940
rect 15180 1920 15198 1940
rect 15198 1920 15205 1940
rect 15175 1915 15205 1920
rect 15285 1940 15315 1945
rect 15285 1920 15290 1940
rect 15290 1920 15308 1940
rect 15308 1920 15315 1940
rect 15285 1915 15315 1920
rect 15395 1940 15425 1945
rect 15395 1920 15400 1940
rect 15400 1920 15418 1940
rect 15418 1920 15425 1940
rect 15395 1915 15425 1920
rect 15505 1940 15535 1945
rect 15505 1920 15510 1940
rect 15510 1920 15528 1940
rect 15528 1920 15535 1940
rect 15505 1915 15535 1920
rect 15615 1940 15645 1945
rect 15615 1920 15620 1940
rect 15620 1920 15638 1940
rect 15638 1920 15645 1940
rect 15615 1915 15645 1920
rect 14645 1865 14675 1895
rect 14820 1730 14850 1760
rect 15410 1730 15440 1760
rect 15740 1730 15770 1760
rect 14520 1675 14550 1705
rect 14885 1675 14915 1705
rect 15110 1700 15140 1705
rect 15110 1680 15115 1700
rect 15115 1680 15135 1700
rect 15135 1680 15140 1700
rect 15110 1675 15140 1680
rect 15310 1700 15340 1705
rect 15310 1680 15315 1700
rect 15315 1680 15335 1700
rect 15335 1680 15340 1700
rect 15310 1675 15340 1680
rect 15510 1700 15540 1705
rect 15510 1680 15515 1700
rect 15515 1680 15535 1700
rect 15535 1680 15540 1700
rect 15510 1675 15540 1680
rect 14820 1640 14855 1645
rect 14820 1615 14825 1640
rect 14825 1615 14850 1640
rect 14850 1615 14855 1640
rect 14820 1610 14855 1615
rect 14880 1640 14915 1645
rect 14880 1615 14885 1640
rect 14885 1615 14910 1640
rect 14910 1615 14915 1640
rect 14880 1610 14915 1615
rect 4810 1590 4840 1595
rect 4810 1570 4815 1590
rect 4815 1570 4835 1590
rect 4835 1570 4840 1590
rect 4810 1565 4840 1570
rect 5415 1565 5445 1595
rect 4270 1540 4300 1545
rect 4270 1520 4275 1540
rect 4275 1520 4295 1540
rect 4295 1520 4300 1540
rect 4270 1515 4300 1520
rect 4390 1540 4420 1545
rect 4390 1520 4395 1540
rect 4395 1520 4415 1540
rect 4415 1520 4420 1540
rect 4390 1515 4420 1520
rect 4510 1540 4540 1545
rect 4510 1520 4515 1540
rect 4515 1520 4535 1540
rect 4535 1520 4540 1540
rect 4510 1515 4540 1520
rect 4630 1540 4660 1545
rect 4630 1520 4635 1540
rect 4635 1520 4655 1540
rect 4655 1520 4660 1540
rect 4630 1515 4660 1520
rect 4750 1540 4780 1545
rect 4750 1520 4755 1540
rect 4755 1520 4775 1540
rect 4775 1520 4780 1540
rect 4750 1515 4780 1520
rect 5140 1515 5170 1545
rect 4210 1495 4240 1500
rect 4210 1475 4215 1495
rect 4215 1475 4235 1495
rect 4235 1475 4240 1495
rect 4210 1470 4240 1475
rect 4330 1495 4360 1500
rect 4330 1475 4335 1495
rect 4335 1475 4355 1495
rect 4355 1475 4360 1495
rect 4330 1470 4360 1475
rect 4450 1495 4480 1500
rect 4450 1475 4455 1495
rect 4455 1475 4475 1495
rect 4475 1475 4480 1495
rect 4450 1470 4480 1475
rect 4690 1495 4720 1500
rect 4690 1475 4695 1495
rect 4695 1475 4715 1495
rect 4715 1475 4720 1495
rect 4690 1470 4720 1475
rect 4810 1495 4840 1500
rect 4810 1475 4815 1495
rect 4815 1475 4835 1495
rect 4835 1475 4840 1495
rect 4810 1470 4840 1475
rect 4930 1495 4960 1500
rect 4930 1475 4935 1495
rect 4935 1475 4955 1495
rect 4955 1475 4960 1495
rect 4930 1470 4960 1475
rect 5050 1495 5080 1500
rect 5050 1475 5055 1495
rect 5055 1475 5075 1495
rect 5075 1475 5080 1495
rect 5050 1470 5080 1475
rect 15740 1360 15770 1390
rect 3380 1180 3410 1185
rect 3380 1160 3385 1180
rect 3385 1160 3405 1180
rect 3405 1160 3410 1180
rect 3380 1155 3410 1160
rect 3990 1155 4020 1185
rect 4600 1180 4630 1185
rect 4600 1160 4605 1180
rect 4605 1160 4625 1180
rect 4625 1160 4630 1180
rect 4600 1155 4630 1160
rect 2950 1120 2980 1125
rect 2950 1100 2955 1120
rect 2955 1100 2975 1120
rect 2975 1100 2980 1120
rect 2950 1095 2980 1100
rect 3030 1120 3060 1125
rect 3030 1100 3035 1120
rect 3035 1100 3055 1120
rect 3055 1100 3060 1120
rect 3030 1095 3060 1100
rect 3110 1120 3140 1125
rect 3110 1100 3115 1120
rect 3115 1100 3135 1120
rect 3135 1100 3140 1120
rect 3110 1095 3140 1100
rect 3190 1120 3220 1125
rect 3190 1100 3195 1120
rect 3195 1100 3215 1120
rect 3215 1100 3220 1120
rect 3190 1095 3220 1100
rect 3270 1120 3300 1125
rect 3270 1100 3275 1120
rect 3275 1100 3295 1120
rect 3295 1100 3300 1120
rect 3270 1095 3300 1100
rect 3350 1120 3380 1125
rect 3350 1100 3355 1120
rect 3355 1100 3375 1120
rect 3375 1100 3380 1120
rect 3350 1095 3380 1100
rect 3430 1120 3460 1125
rect 3430 1100 3435 1120
rect 3435 1100 3455 1120
rect 3455 1100 3460 1120
rect 3430 1095 3460 1100
rect 3510 1120 3540 1125
rect 3510 1100 3515 1120
rect 3515 1100 3535 1120
rect 3535 1100 3540 1120
rect 3510 1095 3540 1100
rect 3590 1120 3620 1125
rect 3590 1100 3595 1120
rect 3595 1100 3615 1120
rect 3615 1100 3620 1120
rect 3590 1095 3620 1100
rect 3670 1120 3700 1125
rect 3670 1100 3675 1120
rect 3675 1100 3695 1120
rect 3695 1100 3700 1120
rect 3670 1095 3700 1100
rect 3750 1120 3780 1125
rect 3750 1100 3755 1120
rect 3755 1100 3775 1120
rect 3775 1100 3780 1120
rect 3750 1095 3780 1100
rect 3830 1120 3860 1125
rect 3830 1100 3835 1120
rect 3835 1100 3855 1120
rect 3855 1100 3860 1120
rect 3830 1095 3860 1100
rect 3910 1120 3940 1125
rect 3910 1100 3915 1120
rect 3915 1100 3935 1120
rect 3935 1100 3940 1120
rect 3910 1095 3940 1100
rect 3990 1120 4020 1125
rect 3990 1100 3995 1120
rect 3995 1100 4015 1120
rect 4015 1100 4020 1120
rect 3990 1095 4020 1100
rect 4070 1120 4100 1125
rect 4070 1100 4075 1120
rect 4075 1100 4095 1120
rect 4095 1100 4100 1120
rect 4070 1095 4100 1100
rect 4150 1120 4180 1125
rect 4150 1100 4155 1120
rect 4155 1100 4175 1120
rect 4175 1100 4180 1120
rect 4150 1095 4180 1100
rect 4230 1120 4260 1125
rect 4230 1100 4235 1120
rect 4235 1100 4255 1120
rect 4255 1100 4260 1120
rect 4230 1095 4260 1100
rect 4310 1120 4340 1125
rect 4310 1100 4315 1120
rect 4315 1100 4335 1120
rect 4335 1100 4340 1120
rect 4310 1095 4340 1100
rect 4390 1120 4420 1125
rect 4390 1100 4395 1120
rect 4395 1100 4415 1120
rect 4415 1100 4420 1120
rect 4390 1095 4420 1100
rect 4470 1120 4500 1125
rect 4470 1100 4475 1120
rect 4475 1100 4495 1120
rect 4495 1100 4500 1120
rect 4470 1095 4500 1100
rect 4550 1120 4580 1125
rect 4550 1100 4555 1120
rect 4555 1100 4575 1120
rect 4575 1100 4580 1120
rect 4550 1095 4580 1100
rect 4630 1120 4660 1125
rect 4630 1100 4635 1120
rect 4635 1100 4655 1120
rect 4655 1100 4660 1120
rect 4630 1095 4660 1100
rect 4710 1120 4740 1125
rect 4710 1100 4715 1120
rect 4715 1100 4735 1120
rect 4735 1100 4740 1120
rect 4710 1095 4740 1100
rect 4790 1120 4820 1125
rect 4790 1100 4795 1120
rect 4795 1100 4815 1120
rect 4815 1100 4820 1120
rect 4790 1095 4820 1100
rect 4870 1120 4900 1125
rect 4870 1100 4875 1120
rect 4875 1100 4895 1120
rect 4895 1100 4900 1120
rect 4870 1095 4900 1100
rect 4950 1120 4980 1125
rect 4950 1100 4955 1120
rect 4955 1100 4975 1120
rect 4975 1100 4980 1120
rect 4950 1095 4980 1100
rect 2625 1010 2655 1040
rect 2910 1035 2940 1040
rect 2910 1015 2915 1035
rect 2915 1015 2935 1035
rect 2935 1015 2940 1035
rect 2910 1010 2940 1015
rect 5115 1035 5145 1040
rect 5115 1015 5120 1035
rect 5120 1015 5140 1035
rect 5140 1015 5145 1035
rect 5115 1010 5145 1015
rect 3000 925 3030 930
rect 3000 905 3005 925
rect 3005 905 3025 925
rect 3025 905 3030 925
rect 3000 900 3030 905
rect 3180 925 3210 930
rect 3180 905 3185 925
rect 3185 905 3205 925
rect 3205 905 3210 925
rect 3180 900 3210 905
rect 3360 925 3390 930
rect 3360 905 3365 925
rect 3365 905 3385 925
rect 3385 905 3390 925
rect 3360 900 3390 905
rect 3540 925 3570 930
rect 3540 905 3545 925
rect 3545 905 3565 925
rect 3565 905 3570 925
rect 3540 900 3570 905
rect 3720 925 3750 930
rect 3720 905 3725 925
rect 3725 905 3745 925
rect 3745 905 3750 925
rect 3720 900 3750 905
rect 3900 925 3930 930
rect 3900 905 3905 925
rect 3905 905 3925 925
rect 3925 905 3930 925
rect 3900 900 3930 905
rect 4080 925 4110 930
rect 4080 905 4085 925
rect 4085 905 4105 925
rect 4105 905 4110 925
rect 4080 900 4110 905
rect 4260 925 4290 930
rect 4260 905 4265 925
rect 4265 905 4285 925
rect 4285 905 4290 925
rect 4260 900 4290 905
rect 4440 925 4470 930
rect 4440 905 4445 925
rect 4445 905 4465 925
rect 4465 905 4470 925
rect 4440 900 4470 905
rect 4620 925 4650 930
rect 4620 905 4625 925
rect 4625 905 4645 925
rect 4645 905 4650 925
rect 4620 900 4650 905
rect 4800 925 4830 930
rect 4800 905 4805 925
rect 4805 905 4825 925
rect 4825 905 4830 925
rect 4800 900 4830 905
rect 4980 925 5010 930
rect 4980 905 4985 925
rect 4985 905 5005 925
rect 5005 905 5010 925
rect 4980 900 5010 905
rect 15210 930 15240 935
rect 15210 910 15215 930
rect 15215 910 15235 930
rect 15235 910 15240 930
rect 15210 905 15240 910
rect 15410 930 15440 935
rect 15410 910 15415 930
rect 15415 910 15435 930
rect 15435 910 15440 930
rect 15410 905 15440 910
rect 17965 3650 17995 3680
rect 17910 3605 17940 3635
rect 17865 2295 17895 2325
rect 16445 2250 16475 2280
rect 16665 2250 16695 2280
rect 16885 2250 16915 2280
rect 17105 2250 17135 2280
rect 17325 2250 17355 2280
rect 16335 2205 16365 2235
rect 16555 2205 16585 2235
rect 16775 2205 16805 2235
rect 16995 2205 17025 2235
rect 17215 2205 17245 2235
rect 17435 2205 17465 2235
rect 16831 2175 16859 2180
rect 16831 2155 16836 2175
rect 16836 2155 16854 2175
rect 16854 2155 16859 2175
rect 16831 2150 16859 2155
rect 16390 1955 16420 1960
rect 16390 1935 16395 1955
rect 16395 1935 16415 1955
rect 16415 1935 16420 1955
rect 16390 1930 16420 1935
rect 16610 1955 16640 1960
rect 16610 1935 16615 1955
rect 16615 1935 16635 1955
rect 16635 1935 16640 1955
rect 16610 1930 16640 1935
rect 16830 1955 16860 1960
rect 16830 1935 16835 1955
rect 16835 1935 16855 1955
rect 16855 1935 16860 1955
rect 16830 1930 16860 1935
rect 17050 1955 17080 1960
rect 17050 1935 17055 1955
rect 17055 1935 17075 1955
rect 17075 1935 17080 1955
rect 17050 1930 17080 1935
rect 17270 1955 17300 1960
rect 17270 1935 17275 1955
rect 17275 1935 17295 1955
rect 17295 1935 17300 1955
rect 17270 1930 17300 1935
rect 16005 1865 16035 1895
rect 16500 1875 16530 1905
rect 16720 1875 16750 1905
rect 16940 1875 16970 1905
rect 17160 1875 17190 1905
rect 16195 1820 16225 1850
rect 16415 1820 16445 1850
rect 16090 1755 16120 1760
rect 16090 1735 16095 1755
rect 16095 1735 16115 1755
rect 16115 1735 16120 1755
rect 16090 1730 16120 1735
rect 16310 1755 16340 1760
rect 16310 1735 16315 1755
rect 16315 1735 16335 1755
rect 16335 1735 16340 1755
rect 16310 1730 16340 1735
rect 17380 1875 17410 1905
rect 17865 1865 17895 1895
rect 16645 1820 16675 1850
rect 17235 1820 17265 1850
rect 17455 1820 17485 1850
rect 17685 1820 17715 1850
rect 16825 1775 16855 1805
rect 16945 1775 16975 1805
rect 16530 1755 16560 1760
rect 16530 1735 16535 1755
rect 16535 1735 16555 1755
rect 16555 1735 16560 1755
rect 16530 1730 16560 1735
rect 17130 1755 17160 1760
rect 17130 1735 17135 1755
rect 17135 1735 17155 1755
rect 17155 1735 17160 1755
rect 17130 1730 17160 1735
rect 17350 1755 17380 1760
rect 17350 1735 17355 1755
rect 17355 1735 17375 1755
rect 17375 1735 17380 1755
rect 17350 1730 17380 1735
rect 17570 1755 17600 1760
rect 17570 1735 17575 1755
rect 17575 1735 17595 1755
rect 17595 1735 17600 1755
rect 17570 1730 17600 1735
rect 16240 1710 16266 1715
rect 16240 1690 16243 1710
rect 16243 1690 16260 1710
rect 16260 1690 16266 1710
rect 16240 1685 16266 1690
rect 16460 1710 16486 1715
rect 16460 1690 16463 1710
rect 16463 1690 16480 1710
rect 16480 1690 16486 1710
rect 16460 1685 16486 1690
rect 16604 1710 16630 1715
rect 16604 1690 16610 1710
rect 16610 1690 16627 1710
rect 16627 1690 16630 1710
rect 16604 1685 16630 1690
rect 16870 1710 16896 1715
rect 16870 1690 16876 1710
rect 16876 1690 16893 1710
rect 16893 1690 16896 1710
rect 16870 1685 16896 1690
rect 17280 1710 17306 1715
rect 17280 1690 17283 1710
rect 17283 1690 17300 1710
rect 17300 1690 17306 1710
rect 17280 1685 17306 1690
rect 17500 1710 17526 1715
rect 17500 1690 17503 1710
rect 17503 1690 17520 1710
rect 17520 1690 17526 1710
rect 17500 1685 17526 1690
rect 17644 1710 17670 1715
rect 17644 1690 17650 1710
rect 17650 1690 17667 1710
rect 17667 1690 17670 1710
rect 17644 1685 17670 1690
rect 16109 1490 16135 1495
rect 16109 1470 16112 1490
rect 16112 1470 16129 1490
rect 16129 1470 16135 1490
rect 16109 1465 16135 1470
rect 16310 1490 16340 1495
rect 16310 1470 16315 1490
rect 16315 1470 16335 1490
rect 16335 1470 16340 1490
rect 16310 1465 16340 1470
rect 16530 1490 16560 1495
rect 16530 1470 16535 1490
rect 16535 1470 16555 1490
rect 16555 1470 16560 1490
rect 16530 1465 16560 1470
rect 16925 1490 16951 1495
rect 16925 1470 16928 1490
rect 16928 1470 16945 1490
rect 16945 1470 16951 1490
rect 16925 1465 16951 1470
rect 17149 1490 17175 1495
rect 17149 1470 17152 1490
rect 17152 1470 17169 1490
rect 17169 1470 17175 1490
rect 17149 1465 17175 1470
rect 17350 1490 17380 1495
rect 17350 1470 17355 1490
rect 17355 1470 17375 1490
rect 17375 1470 17380 1490
rect 17350 1465 17380 1470
rect 17570 1490 17600 1495
rect 17570 1470 17575 1490
rect 17575 1470 17595 1490
rect 17595 1470 17600 1490
rect 17570 1465 17600 1470
rect 16150 1430 16180 1435
rect 16150 1410 16155 1430
rect 16155 1410 16175 1430
rect 16175 1410 16180 1430
rect 16150 1405 16180 1410
rect 16255 1430 16285 1435
rect 16255 1410 16260 1430
rect 16260 1410 16280 1430
rect 16280 1410 16285 1430
rect 16255 1405 16285 1410
rect 16365 1430 16395 1435
rect 16365 1410 16370 1430
rect 16370 1410 16390 1430
rect 16390 1410 16395 1430
rect 16365 1405 16395 1410
rect 16475 1430 16505 1435
rect 16475 1410 16480 1430
rect 16480 1410 16500 1430
rect 16500 1410 16505 1430
rect 16475 1405 16505 1410
rect 16585 1430 16615 1435
rect 16585 1410 16590 1430
rect 16590 1410 16610 1430
rect 16610 1410 16615 1430
rect 16585 1405 16615 1410
rect 16010 1315 16040 1345
rect 16815 1315 16845 1345
rect 16320 1265 16350 1295
rect 17190 1430 17220 1435
rect 17190 1410 17195 1430
rect 17195 1410 17215 1430
rect 17215 1410 17220 1430
rect 17190 1405 17220 1410
rect 17295 1430 17325 1435
rect 17295 1410 17300 1430
rect 17300 1410 17320 1430
rect 17320 1410 17325 1430
rect 17295 1405 17325 1410
rect 17405 1430 17435 1435
rect 17405 1410 17410 1430
rect 17410 1410 17430 1430
rect 17430 1410 17435 1430
rect 17405 1405 17435 1410
rect 17515 1430 17545 1435
rect 17515 1410 17520 1430
rect 17520 1410 17540 1430
rect 17540 1410 17545 1430
rect 17515 1405 17545 1410
rect 17625 1430 17655 1435
rect 17625 1410 17630 1430
rect 17630 1410 17650 1430
rect 17650 1410 17655 1430
rect 17625 1405 17655 1410
rect 16885 1265 16915 1295
rect 16430 1230 16460 1235
rect 16430 1210 16435 1230
rect 16435 1210 16455 1230
rect 16455 1210 16460 1230
rect 16430 1205 16460 1210
rect 16540 1230 16570 1235
rect 16540 1210 16545 1230
rect 16545 1210 16565 1230
rect 16565 1210 16570 1230
rect 16540 1205 16570 1210
rect 16650 1230 16680 1235
rect 16650 1210 16655 1230
rect 16655 1210 16675 1230
rect 16675 1210 16680 1230
rect 16650 1205 16680 1210
rect 16760 1230 16790 1235
rect 16760 1210 16765 1230
rect 16765 1210 16785 1230
rect 16785 1210 16790 1230
rect 16760 1205 16790 1210
rect 16870 1230 16900 1235
rect 16870 1210 16875 1230
rect 16875 1210 16895 1230
rect 16895 1210 16900 1230
rect 16870 1205 16900 1210
rect 16980 1230 17010 1235
rect 16980 1210 16985 1230
rect 16985 1210 17005 1230
rect 17005 1210 17010 1230
rect 16980 1205 17010 1210
rect 17090 1230 17120 1235
rect 17090 1210 17095 1230
rect 17095 1210 17115 1230
rect 17115 1210 17120 1230
rect 17090 1205 17120 1210
rect 17200 1230 17230 1235
rect 17200 1210 17205 1230
rect 17205 1210 17225 1230
rect 17225 1210 17230 1230
rect 17200 1205 17230 1210
rect 17310 1230 17340 1235
rect 17310 1210 17315 1230
rect 17315 1210 17335 1230
rect 17335 1210 17340 1230
rect 17310 1205 17340 1210
rect 17420 1230 17450 1235
rect 17420 1210 17425 1230
rect 17425 1210 17445 1230
rect 17445 1210 17450 1230
rect 17420 1205 17450 1210
rect 17530 1230 17560 1235
rect 17530 1210 17535 1230
rect 17535 1210 17555 1230
rect 17555 1210 17560 1230
rect 17530 1205 17560 1210
rect 17600 1245 17630 1250
rect 17600 1225 17605 1245
rect 17605 1225 17625 1245
rect 17625 1225 17630 1245
rect 17600 1220 17630 1225
rect 17910 1220 17940 1250
rect 16170 910 16200 915
rect 16170 890 16175 910
rect 16175 890 16195 910
rect 16195 890 16200 910
rect 16170 885 16200 890
rect 16265 910 16295 915
rect 16265 890 16270 910
rect 16270 890 16290 910
rect 16290 890 16295 910
rect 16265 885 16295 890
rect 16375 910 16405 915
rect 16375 890 16380 910
rect 16380 890 16400 910
rect 16400 890 16405 910
rect 16375 885 16405 890
rect 16485 910 16515 915
rect 16485 890 16490 910
rect 16490 890 16510 910
rect 16510 890 16515 910
rect 16485 885 16515 890
rect 16595 910 16625 915
rect 16595 890 16600 910
rect 16600 890 16620 910
rect 16620 890 16625 910
rect 16595 885 16625 890
rect 16705 910 16735 915
rect 16705 890 16710 910
rect 16710 890 16730 910
rect 16730 890 16735 910
rect 16705 885 16735 890
rect 16815 910 16845 915
rect 16815 890 16820 910
rect 16820 890 16840 910
rect 16840 890 16845 910
rect 16815 885 16845 890
rect 16925 910 16955 915
rect 16925 890 16930 910
rect 16930 890 16950 910
rect 16950 890 16955 910
rect 16925 885 16955 890
rect 17035 910 17065 915
rect 17035 890 17040 910
rect 17040 890 17060 910
rect 17060 890 17065 910
rect 17035 885 17065 890
rect 17145 910 17175 915
rect 17145 890 17150 910
rect 17150 890 17170 910
rect 17170 890 17175 910
rect 17145 885 17175 890
rect 17255 910 17285 915
rect 17255 890 17260 910
rect 17260 890 17280 910
rect 17280 890 17285 910
rect 17255 885 17285 890
rect 17365 910 17395 915
rect 17365 890 17370 910
rect 17370 890 17390 910
rect 17390 890 17395 910
rect 17365 885 17395 890
rect 17475 910 17505 915
rect 17475 890 17480 910
rect 17480 890 17500 910
rect 17500 890 17505 910
rect 17475 885 17505 890
rect 17625 910 17655 915
rect 17625 890 17630 910
rect 17630 890 17650 910
rect 17650 890 17655 910
rect 17625 885 17655 890
rect 16010 825 16040 855
rect 16500 825 16530 855
rect 16940 830 16970 860
rect 17160 830 17190 860
rect 17380 830 17410 860
rect 18205 3630 18235 3635
rect 18205 3610 18210 3630
rect 18210 3610 18230 3630
rect 18230 3610 18235 3630
rect 18205 3605 18235 3610
rect 18315 3630 18345 3635
rect 18315 3610 18320 3630
rect 18320 3610 18340 3630
rect 18340 3610 18345 3630
rect 18315 3605 18345 3610
rect 18425 3630 18455 3635
rect 18425 3610 18430 3630
rect 18430 3610 18450 3630
rect 18450 3610 18455 3630
rect 18425 3605 18455 3610
rect 18535 3630 18565 3635
rect 18535 3610 18540 3630
rect 18540 3610 18560 3630
rect 18560 3610 18565 3630
rect 18535 3605 18565 3610
rect 18645 3630 18675 3635
rect 18645 3610 18650 3630
rect 18650 3610 18670 3630
rect 18670 3610 18675 3630
rect 18645 3605 18675 3610
rect 18755 3630 18785 3635
rect 18755 3610 18760 3630
rect 18760 3610 18780 3630
rect 18780 3610 18785 3630
rect 18755 3605 18785 3610
rect 19160 3605 19190 3635
rect 24610 3605 24640 3635
rect 25065 3630 25095 3635
rect 25065 3610 25070 3630
rect 25070 3610 25090 3630
rect 25090 3610 25095 3630
rect 25065 3605 25095 3610
rect 25175 3630 25205 3635
rect 25175 3610 25180 3630
rect 25180 3610 25200 3630
rect 25200 3610 25205 3630
rect 25175 3605 25205 3610
rect 25285 3630 25315 3635
rect 25285 3610 25290 3630
rect 25290 3610 25310 3630
rect 25310 3610 25315 3630
rect 25285 3605 25315 3610
rect 25395 3630 25425 3635
rect 25395 3610 25400 3630
rect 25400 3610 25420 3630
rect 25420 3610 25425 3630
rect 25395 3605 25425 3610
rect 25505 3630 25535 3635
rect 25505 3610 25510 3630
rect 25510 3610 25530 3630
rect 25530 3610 25535 3630
rect 25505 3605 25535 3610
rect 25615 3630 25645 3635
rect 25615 3610 25620 3630
rect 25620 3610 25640 3630
rect 25640 3610 25645 3630
rect 25615 3605 25645 3610
rect 19110 3525 19140 3555
rect 19160 3525 19190 3555
rect 19210 3525 19240 3555
rect 24560 3525 24590 3555
rect 24610 3525 24640 3555
rect 24660 3525 24690 3555
rect 27300 4765 27330 4770
rect 27300 4745 27305 4765
rect 27305 4745 27325 4765
rect 27325 4745 27330 4765
rect 27300 4740 27330 4745
rect 27420 4765 27450 4770
rect 27420 4745 27425 4765
rect 27425 4745 27445 4765
rect 27445 4745 27450 4765
rect 27420 4740 27450 4745
rect 27540 4765 27570 4770
rect 27540 4745 27545 4765
rect 27545 4745 27565 4765
rect 27565 4745 27570 4765
rect 27540 4740 27570 4745
rect 27660 4765 27690 4770
rect 27660 4745 27665 4765
rect 27665 4745 27685 4765
rect 27685 4745 27690 4765
rect 27660 4740 27690 4745
rect 26110 4555 26140 4585
rect 26350 4555 26380 4585
rect 27360 4555 27390 4585
rect 26055 3155 26085 3185
rect 18260 2960 18290 2965
rect 18260 2940 18265 2960
rect 18265 2940 18285 2960
rect 18285 2940 18290 2960
rect 18260 2935 18290 2940
rect 18370 2960 18400 2965
rect 18370 2940 18375 2960
rect 18375 2940 18395 2960
rect 18395 2940 18400 2960
rect 18370 2935 18400 2940
rect 18480 2960 18510 2965
rect 18480 2940 18485 2960
rect 18485 2940 18505 2960
rect 18505 2940 18510 2960
rect 18480 2935 18510 2940
rect 18590 2960 18620 2965
rect 18590 2940 18595 2960
rect 18595 2940 18615 2960
rect 18615 2940 18620 2960
rect 18590 2935 18620 2940
rect 18700 2960 18730 2965
rect 18700 2940 18705 2960
rect 18705 2940 18725 2960
rect 18725 2940 18730 2960
rect 18700 2935 18730 2940
rect 18020 2850 18050 2880
rect 18315 2850 18345 2880
rect 19110 2905 19140 2935
rect 19160 2905 19190 2935
rect 19210 2905 19240 2935
rect 24560 2905 24590 2935
rect 24610 2905 24640 2935
rect 24660 2905 24690 2935
rect 25120 2960 25150 2965
rect 25120 2940 25125 2960
rect 25125 2940 25145 2960
rect 25145 2940 25150 2960
rect 25120 2935 25150 2940
rect 25230 2960 25260 2965
rect 25230 2940 25235 2960
rect 25235 2940 25255 2960
rect 25255 2940 25260 2960
rect 25230 2935 25260 2940
rect 25340 2960 25370 2965
rect 25340 2940 25345 2960
rect 25345 2940 25365 2960
rect 25365 2940 25370 2960
rect 25340 2935 25370 2940
rect 25450 2960 25480 2965
rect 25450 2940 25455 2960
rect 25455 2940 25475 2960
rect 25475 2940 25480 2960
rect 25450 2935 25480 2940
rect 25560 2960 25590 2965
rect 25560 2940 25565 2960
rect 25565 2940 25585 2960
rect 25585 2940 25590 2960
rect 25560 2935 25590 2940
rect 26365 4475 26395 4480
rect 26365 4455 26370 4475
rect 26370 4455 26390 4475
rect 26390 4455 26395 4475
rect 26365 4450 26395 4455
rect 26475 4475 26505 4480
rect 26475 4455 26480 4475
rect 26480 4455 26500 4475
rect 26500 4455 26505 4475
rect 26475 4450 26505 4455
rect 26585 4475 26615 4480
rect 26585 4455 26590 4475
rect 26590 4455 26610 4475
rect 26610 4455 26615 4475
rect 26585 4450 26615 4455
rect 26695 4475 26725 4480
rect 26695 4455 26700 4475
rect 26700 4455 26720 4475
rect 26720 4455 26725 4475
rect 26695 4450 26725 4455
rect 26805 4475 26835 4480
rect 26805 4455 26810 4475
rect 26810 4455 26830 4475
rect 26830 4455 26835 4475
rect 26805 4450 26835 4455
rect 26915 4475 26945 4480
rect 26915 4455 26920 4475
rect 26920 4455 26940 4475
rect 26940 4455 26945 4475
rect 26915 4450 26945 4455
rect 27025 4475 27055 4480
rect 27025 4455 27030 4475
rect 27030 4455 27050 4475
rect 27050 4455 27055 4475
rect 27025 4450 27055 4455
rect 27135 4475 27165 4480
rect 27135 4455 27140 4475
rect 27140 4455 27160 4475
rect 27160 4455 27165 4475
rect 27135 4450 27165 4455
rect 27245 4475 27275 4480
rect 27245 4455 27250 4475
rect 27250 4455 27270 4475
rect 27270 4455 27275 4475
rect 27245 4450 27275 4455
rect 27355 4475 27385 4480
rect 27355 4455 27360 4475
rect 27360 4455 27380 4475
rect 27380 4455 27385 4475
rect 27355 4450 27385 4455
rect 26310 4355 26340 4360
rect 26310 4335 26315 4355
rect 26315 4335 26335 4355
rect 26335 4335 26340 4355
rect 26310 4330 26340 4335
rect 26530 4355 26560 4360
rect 26530 4335 26535 4355
rect 26535 4335 26555 4355
rect 26555 4335 26560 4355
rect 26530 4330 26560 4335
rect 26750 4355 26780 4360
rect 26750 4335 26755 4355
rect 26755 4335 26775 4355
rect 26775 4335 26780 4355
rect 26750 4330 26780 4335
rect 26970 4355 27000 4360
rect 26970 4335 26975 4355
rect 26975 4335 26995 4355
rect 26995 4335 27000 4355
rect 26970 4330 27000 4335
rect 27190 4355 27220 4360
rect 27190 4335 27195 4355
rect 27195 4335 27215 4355
rect 27215 4335 27220 4355
rect 27190 4330 27220 4335
rect 27410 4355 27440 4360
rect 27410 4335 27415 4355
rect 27415 4335 27435 4355
rect 27435 4335 27440 4355
rect 27410 4330 27440 4335
rect 26325 4100 26355 4130
rect 26425 4215 26455 4245
rect 26640 4215 26670 4245
rect 26860 4215 26890 4245
rect 27080 4215 27110 4245
rect 27300 4215 27330 4245
rect 26425 4100 26455 4130
rect 26535 4100 26565 4130
rect 26645 4100 26675 4130
rect 26755 4100 26785 4130
rect 27055 4100 27085 4130
rect 27155 4100 27185 4130
rect 27265 4100 27295 4130
rect 27375 4100 27405 4130
rect 27485 4100 27515 4130
rect 26282 4065 26308 4069
rect 26282 4045 26285 4065
rect 26285 4045 26305 4065
rect 26305 4045 26308 4065
rect 26282 4041 26308 4045
rect 26482 4065 26508 4069
rect 26482 4045 26485 4065
rect 26485 4045 26505 4065
rect 26505 4045 26508 4065
rect 26482 4041 26508 4045
rect 27010 4065 27036 4069
rect 27010 4045 27013 4065
rect 27013 4045 27033 4065
rect 27033 4045 27036 4065
rect 27010 4041 27036 4045
rect 27210 4065 27240 4070
rect 27210 4045 27215 4065
rect 27215 4045 27235 4065
rect 27235 4045 27240 4065
rect 27210 4040 27240 4045
rect 27430 4065 27460 4070
rect 27430 4045 27435 4065
rect 27435 4045 27455 4065
rect 27455 4045 27460 4065
rect 27430 4040 27460 4045
rect 27875 4040 27905 4070
rect 26410 3945 26436 3950
rect 26410 3925 26413 3945
rect 26413 3925 26430 3945
rect 26430 3925 26436 3945
rect 26410 3920 26436 3925
rect 26630 3945 26656 3950
rect 26630 3925 26633 3945
rect 26633 3925 26650 3945
rect 26650 3925 26656 3945
rect 26630 3920 26656 3925
rect 26774 3945 26800 3950
rect 26774 3925 26780 3945
rect 26780 3925 26797 3945
rect 26797 3925 26800 3945
rect 26774 3920 26800 3925
rect 27140 3945 27166 3950
rect 27140 3925 27143 3945
rect 27143 3925 27160 3945
rect 27160 3925 27166 3945
rect 27140 3920 27166 3925
rect 27360 3945 27386 3950
rect 27360 3925 27363 3945
rect 27363 3925 27380 3945
rect 27380 3925 27386 3945
rect 27360 3920 27386 3925
rect 27504 3945 27530 3950
rect 27504 3925 27510 3945
rect 27510 3925 27527 3945
rect 27527 3925 27530 3945
rect 27504 3920 27530 3925
rect 26260 3860 26290 3890
rect 26365 3860 26395 3890
rect 26480 3860 26510 3890
rect 26585 3860 26615 3890
rect 26700 3860 26730 3890
rect 26815 3860 26845 3890
rect 26990 3860 27020 3890
rect 27210 3860 27240 3890
rect 27430 3860 27460 3890
rect 27095 3750 27125 3780
rect 27315 3750 27345 3780
rect 27545 3750 27575 3780
rect 26345 3650 26375 3655
rect 26345 3630 26350 3650
rect 26350 3630 26370 3650
rect 26370 3630 26375 3650
rect 26345 3625 26375 3630
rect 26465 3650 26495 3655
rect 26465 3630 26470 3650
rect 26470 3630 26490 3650
rect 26490 3630 26495 3650
rect 26465 3625 26495 3630
rect 26585 3650 26615 3655
rect 26585 3630 26590 3650
rect 26590 3630 26610 3650
rect 26610 3630 26615 3650
rect 26585 3625 26615 3630
rect 26705 3650 26735 3655
rect 26705 3630 26710 3650
rect 26710 3630 26730 3650
rect 26730 3630 26735 3650
rect 26705 3625 26735 3630
rect 26825 3650 26855 3655
rect 26825 3630 26830 3650
rect 26830 3630 26850 3650
rect 26850 3630 26855 3650
rect 26825 3625 26855 3630
rect 26945 3650 26975 3655
rect 26945 3630 26950 3650
rect 26950 3630 26970 3650
rect 26970 3630 26975 3650
rect 26945 3625 26975 3630
rect 27065 3650 27095 3655
rect 27065 3630 27070 3650
rect 27070 3630 27090 3650
rect 27090 3630 27095 3650
rect 27065 3625 27095 3630
rect 27185 3650 27215 3655
rect 27185 3630 27190 3650
rect 27190 3630 27210 3650
rect 27210 3630 27215 3650
rect 27185 3625 27215 3630
rect 27305 3650 27335 3655
rect 27305 3630 27310 3650
rect 27310 3630 27330 3650
rect 27330 3630 27335 3650
rect 27305 3625 27335 3630
rect 27425 3650 27455 3655
rect 27425 3630 27430 3650
rect 27430 3630 27450 3650
rect 27450 3630 27455 3650
rect 27425 3625 27455 3630
rect 26826 3180 26854 3185
rect 26826 3160 26831 3180
rect 26831 3160 26849 3180
rect 26849 3160 26854 3180
rect 26826 3155 26854 3160
rect 26285 3100 26315 3130
rect 26525 3100 26555 3130
rect 26765 3100 26795 3130
rect 27005 3100 27035 3130
rect 27245 3100 27275 3130
rect 26405 2975 26435 3005
rect 26645 2975 26675 3005
rect 26885 2975 26915 3005
rect 27125 2975 27155 3005
rect 19160 2850 19190 2880
rect 24610 2850 24640 2880
rect 26110 2920 26140 2950
rect 26885 2920 26915 2950
rect 25505 2850 25535 2880
rect 25785 2850 25815 2880
rect 26140 2890 26170 2895
rect 26140 2870 26145 2890
rect 26145 2870 26165 2890
rect 26165 2870 26170 2890
rect 26140 2865 26170 2870
rect 26260 2890 26290 2895
rect 26260 2870 26265 2890
rect 26265 2870 26285 2890
rect 26285 2870 26290 2890
rect 26260 2865 26290 2870
rect 26380 2890 26410 2895
rect 26380 2870 26385 2890
rect 26385 2870 26405 2890
rect 26405 2870 26410 2890
rect 26380 2865 26410 2870
rect 26500 2890 26530 2895
rect 26500 2870 26505 2890
rect 26505 2870 26525 2890
rect 26525 2870 26530 2890
rect 26500 2865 26530 2870
rect 26620 2890 26650 2895
rect 26620 2870 26625 2890
rect 26625 2870 26645 2890
rect 26645 2870 26650 2890
rect 26620 2865 26650 2870
rect 18590 2795 18620 2825
rect 19250 2795 19280 2825
rect 24520 2795 24550 2825
rect 25230 2795 25260 2825
rect 18205 2700 18235 2705
rect 18205 2680 18210 2700
rect 18210 2680 18230 2700
rect 18230 2680 18235 2700
rect 18205 2675 18235 2680
rect 18315 2700 18345 2705
rect 18315 2680 18320 2700
rect 18320 2680 18340 2700
rect 18340 2680 18345 2700
rect 18315 2675 18345 2680
rect 18425 2700 18455 2705
rect 18425 2680 18430 2700
rect 18430 2680 18450 2700
rect 18450 2680 18455 2700
rect 18425 2675 18455 2680
rect 18535 2700 18565 2705
rect 18535 2680 18540 2700
rect 18540 2680 18560 2700
rect 18560 2680 18565 2700
rect 18535 2675 18565 2680
rect 18645 2700 18675 2705
rect 18645 2680 18650 2700
rect 18650 2680 18670 2700
rect 18670 2680 18675 2700
rect 18645 2675 18675 2680
rect 18755 2700 18785 2705
rect 18755 2680 18760 2700
rect 18760 2680 18780 2700
rect 18780 2680 18785 2700
rect 18755 2675 18785 2680
rect 18260 2430 18290 2435
rect 18260 2410 18265 2430
rect 18265 2410 18285 2430
rect 18285 2410 18290 2430
rect 18260 2405 18290 2410
rect 18370 2430 18400 2435
rect 18370 2410 18375 2430
rect 18375 2410 18395 2430
rect 18395 2410 18400 2430
rect 18370 2405 18400 2410
rect 18480 2430 18510 2435
rect 18480 2410 18485 2430
rect 18485 2410 18505 2430
rect 18505 2410 18510 2430
rect 18480 2405 18510 2410
rect 18590 2430 18620 2435
rect 18590 2410 18595 2430
rect 18595 2410 18615 2430
rect 18615 2410 18620 2430
rect 18590 2405 18620 2410
rect 18700 2430 18730 2435
rect 18700 2410 18705 2430
rect 18705 2410 18725 2430
rect 18725 2410 18730 2430
rect 18700 2405 18730 2410
rect 18945 2405 18975 2435
rect 18020 2345 18050 2375
rect 18230 2370 18260 2375
rect 18230 2350 18235 2370
rect 18235 2350 18255 2370
rect 18255 2350 18260 2370
rect 18230 2345 18260 2350
rect 18260 2310 18290 2315
rect 18260 2290 18265 2310
rect 18265 2290 18285 2310
rect 18285 2290 18290 2310
rect 18260 2285 18290 2290
rect 18370 2310 18400 2315
rect 18370 2290 18375 2310
rect 18375 2290 18395 2310
rect 18395 2290 18400 2310
rect 18370 2285 18400 2290
rect 18480 2310 18510 2315
rect 18480 2290 18485 2310
rect 18485 2290 18505 2310
rect 18505 2290 18510 2310
rect 18480 2285 18510 2290
rect 18590 2310 18620 2315
rect 18590 2290 18595 2310
rect 18595 2290 18615 2310
rect 18615 2290 18620 2310
rect 18590 2285 18620 2290
rect 18700 2310 18730 2315
rect 18700 2290 18705 2310
rect 18705 2290 18725 2310
rect 18725 2290 18730 2310
rect 18700 2285 18730 2290
rect 18900 2285 18930 2315
rect 25065 2700 25095 2705
rect 25065 2680 25070 2700
rect 25070 2680 25090 2700
rect 25090 2680 25095 2700
rect 25065 2675 25095 2680
rect 25175 2700 25205 2705
rect 25175 2680 25180 2700
rect 25180 2680 25200 2700
rect 25200 2680 25205 2700
rect 25175 2675 25205 2680
rect 25285 2700 25315 2705
rect 25285 2680 25290 2700
rect 25290 2680 25310 2700
rect 25310 2680 25315 2700
rect 25285 2675 25315 2680
rect 25395 2700 25425 2705
rect 25395 2680 25400 2700
rect 25400 2680 25420 2700
rect 25420 2680 25425 2700
rect 25395 2675 25425 2680
rect 25505 2700 25535 2705
rect 25505 2680 25510 2700
rect 25510 2680 25530 2700
rect 25530 2680 25535 2700
rect 25505 2675 25535 2680
rect 25615 2700 25645 2705
rect 25615 2680 25620 2700
rect 25620 2680 25640 2700
rect 25640 2680 25645 2700
rect 25615 2675 25645 2680
rect 24875 2405 24905 2435
rect 25120 2430 25150 2435
rect 25120 2410 25125 2430
rect 25125 2410 25145 2430
rect 25145 2410 25150 2430
rect 25120 2405 25150 2410
rect 25230 2430 25260 2435
rect 25230 2410 25235 2430
rect 25235 2410 25255 2430
rect 25255 2410 25260 2430
rect 25230 2405 25260 2410
rect 25340 2430 25370 2435
rect 25340 2410 25345 2430
rect 25345 2410 25365 2430
rect 25365 2410 25370 2430
rect 25340 2405 25370 2410
rect 25450 2430 25480 2435
rect 25450 2410 25455 2430
rect 25455 2410 25475 2430
rect 25475 2410 25480 2430
rect 25450 2405 25480 2410
rect 25560 2430 25590 2435
rect 25560 2410 25565 2430
rect 25565 2410 25585 2430
rect 25585 2410 25590 2430
rect 25560 2405 25590 2410
rect 19250 2080 19280 2110
rect 24520 2080 24550 2110
rect 18945 1970 18975 2000
rect 18995 2000 19030 2005
rect 18995 1975 19000 2000
rect 19000 1975 19025 2000
rect 19025 1975 19030 2000
rect 18995 1970 19030 1975
rect 19055 2000 19090 2005
rect 19055 1975 19060 2000
rect 19060 1975 19085 2000
rect 19085 1975 19090 2000
rect 19055 1970 19090 1975
rect 19115 2000 19150 2005
rect 19115 1975 19120 2000
rect 19120 1975 19145 2000
rect 19145 1975 19150 2000
rect 19115 1970 19150 1975
rect 19175 2000 19210 2005
rect 19175 1975 19180 2000
rect 19180 1975 19205 2000
rect 19205 1975 19210 2000
rect 19175 1970 19210 1975
rect 18205 1940 18235 1945
rect 18205 1920 18212 1940
rect 18212 1920 18230 1940
rect 18230 1920 18235 1940
rect 18205 1915 18235 1920
rect 18315 1940 18345 1945
rect 18315 1920 18322 1940
rect 18322 1920 18340 1940
rect 18340 1920 18345 1940
rect 18315 1915 18345 1920
rect 18425 1940 18455 1945
rect 18425 1920 18432 1940
rect 18432 1920 18450 1940
rect 18450 1920 18455 1940
rect 18425 1915 18455 1920
rect 18535 1940 18565 1945
rect 18535 1920 18542 1940
rect 18542 1920 18560 1940
rect 18560 1920 18565 1940
rect 18535 1915 18565 1920
rect 18645 1940 18675 1945
rect 18645 1920 18652 1940
rect 18652 1920 18670 1940
rect 18670 1920 18675 1940
rect 18645 1915 18675 1920
rect 18755 1940 18785 1945
rect 18755 1920 18762 1940
rect 18762 1920 18780 1940
rect 18780 1920 18785 1940
rect 18755 1915 18785 1920
rect 18900 1915 18930 1945
rect 19055 1915 19085 1945
rect 19175 1865 19205 1895
rect 18080 1730 18110 1760
rect 18410 1730 18440 1760
rect 19000 1730 19030 1760
rect 18310 1700 18340 1705
rect 18310 1680 18315 1700
rect 18315 1680 18335 1700
rect 18335 1680 18340 1700
rect 18310 1675 18340 1680
rect 18510 1700 18540 1705
rect 18510 1680 18515 1700
rect 18515 1680 18535 1700
rect 18535 1680 18540 1700
rect 18510 1675 18540 1680
rect 18710 1700 18740 1705
rect 18710 1680 18715 1700
rect 18715 1680 18735 1700
rect 18735 1680 18740 1700
rect 18710 1675 18740 1680
rect 18935 1675 18965 1705
rect 24640 2000 24675 2005
rect 24640 1975 24645 2000
rect 24645 1975 24670 2000
rect 24670 1975 24675 2000
rect 24640 1970 24675 1975
rect 24700 2000 24735 2005
rect 24700 1975 24705 2000
rect 24705 1975 24730 2000
rect 24730 1975 24735 2000
rect 24700 1970 24735 1975
rect 24760 2000 24795 2005
rect 24760 1975 24765 2000
rect 24765 1975 24790 2000
rect 24790 1975 24795 2000
rect 24760 1970 24795 1975
rect 26080 2470 26110 2475
rect 26080 2450 26085 2470
rect 26085 2450 26105 2470
rect 26105 2450 26110 2470
rect 26080 2445 26110 2450
rect 26200 2470 26230 2475
rect 26200 2450 26205 2470
rect 26205 2450 26225 2470
rect 26225 2450 26230 2470
rect 26200 2445 26230 2450
rect 26320 2470 26350 2475
rect 26320 2450 26325 2470
rect 26325 2450 26345 2470
rect 26345 2450 26350 2470
rect 26320 2445 26350 2450
rect 26440 2470 26470 2475
rect 26440 2450 26445 2470
rect 26445 2450 26465 2470
rect 26465 2450 26470 2470
rect 26440 2445 26470 2450
rect 26560 2470 26590 2475
rect 26560 2450 26565 2470
rect 26565 2450 26585 2470
rect 26585 2450 26590 2470
rect 26560 2445 26590 2450
rect 26680 2470 26710 2475
rect 26680 2450 26685 2470
rect 26685 2450 26705 2470
rect 26705 2450 26710 2470
rect 26680 2445 26710 2450
rect 27485 3100 27515 3130
rect 27365 2975 27395 3005
rect 27160 2890 27190 2895
rect 27160 2870 27165 2890
rect 27165 2870 27185 2890
rect 27185 2870 27190 2890
rect 27160 2865 27190 2870
rect 27280 2890 27310 2895
rect 27280 2870 27285 2890
rect 27285 2870 27305 2890
rect 27305 2870 27310 2890
rect 27280 2865 27310 2870
rect 27400 2890 27430 2895
rect 27400 2870 27405 2890
rect 27405 2870 27425 2890
rect 27425 2870 27430 2890
rect 27400 2865 27430 2870
rect 27520 2890 27550 2895
rect 27520 2870 27525 2890
rect 27525 2870 27545 2890
rect 27545 2870 27550 2890
rect 27520 2865 27550 2870
rect 27640 2890 27670 2895
rect 27640 2870 27645 2890
rect 27645 2870 27665 2890
rect 27665 2870 27670 2890
rect 27640 2865 27670 2870
rect 27100 2470 27130 2475
rect 27100 2450 27105 2470
rect 27105 2450 27125 2470
rect 27125 2450 27130 2470
rect 27100 2445 27130 2450
rect 27220 2470 27250 2475
rect 27220 2450 27225 2470
rect 27225 2450 27245 2470
rect 27245 2450 27250 2470
rect 27220 2445 27250 2450
rect 27340 2470 27370 2475
rect 27340 2450 27345 2470
rect 27345 2450 27365 2470
rect 27365 2450 27370 2470
rect 27340 2445 27370 2450
rect 27460 2470 27490 2475
rect 27460 2450 27465 2470
rect 27465 2450 27485 2470
rect 27485 2450 27490 2470
rect 27460 2445 27490 2450
rect 27580 2470 27610 2475
rect 27580 2450 27585 2470
rect 27585 2450 27605 2470
rect 27605 2450 27610 2470
rect 27580 2445 27610 2450
rect 27700 2470 27730 2475
rect 27700 2450 27705 2470
rect 27705 2450 27725 2470
rect 27725 2450 27730 2470
rect 27700 2445 27730 2450
rect 26380 2390 26410 2420
rect 26885 2390 26915 2420
rect 27400 2390 27430 2420
rect 25590 2370 25620 2375
rect 25590 2350 25595 2370
rect 25595 2350 25615 2370
rect 25615 2350 25620 2370
rect 25590 2345 25620 2350
rect 25785 2345 25815 2375
rect 26325 2345 26355 2375
rect 27325 2345 27355 2375
rect 24920 2285 24950 2315
rect 25120 2310 25150 2315
rect 25120 2290 25125 2310
rect 25125 2290 25145 2310
rect 25145 2290 25150 2310
rect 25120 2285 25150 2290
rect 25230 2310 25260 2315
rect 25230 2290 25235 2310
rect 25235 2290 25255 2310
rect 25255 2290 25260 2310
rect 25230 2285 25260 2290
rect 25340 2310 25370 2315
rect 25340 2290 25345 2310
rect 25345 2290 25365 2310
rect 25365 2290 25370 2310
rect 25340 2285 25370 2290
rect 25450 2310 25480 2315
rect 25450 2290 25455 2310
rect 25455 2290 25475 2310
rect 25475 2290 25480 2310
rect 25450 2285 25480 2290
rect 25560 2310 25590 2315
rect 25560 2290 25565 2310
rect 25565 2290 25585 2310
rect 25585 2290 25590 2310
rect 25560 2285 25590 2290
rect 26005 2295 26035 2325
rect 24820 2000 24855 2005
rect 24820 1975 24825 2000
rect 24825 1975 24850 2000
rect 24850 1975 24855 2000
rect 24820 1970 24855 1975
rect 24875 1970 24905 2000
rect 25805 2150 25835 2180
rect 24765 1915 24795 1945
rect 24920 1915 24950 1945
rect 25065 1940 25095 1945
rect 25065 1920 25070 1940
rect 25070 1920 25088 1940
rect 25088 1920 25095 1940
rect 25065 1915 25095 1920
rect 25175 1940 25205 1945
rect 25175 1920 25180 1940
rect 25180 1920 25198 1940
rect 25198 1920 25205 1940
rect 25175 1915 25205 1920
rect 25285 1940 25315 1945
rect 25285 1920 25290 1940
rect 25290 1920 25308 1940
rect 25308 1920 25315 1940
rect 25285 1915 25315 1920
rect 25395 1940 25425 1945
rect 25395 1920 25400 1940
rect 25400 1920 25418 1940
rect 25418 1920 25425 1940
rect 25395 1915 25425 1920
rect 25505 1940 25535 1945
rect 25505 1920 25510 1940
rect 25510 1920 25528 1940
rect 25528 1920 25535 1940
rect 25505 1915 25535 1920
rect 25615 1940 25645 1945
rect 25615 1920 25620 1940
rect 25620 1920 25638 1940
rect 25638 1920 25645 1940
rect 25615 1915 25645 1920
rect 24645 1865 24675 1895
rect 24820 1730 24850 1760
rect 25410 1730 25440 1760
rect 25740 1730 25770 1760
rect 19250 1675 19280 1705
rect 24520 1675 24550 1705
rect 24885 1675 24915 1705
rect 25110 1700 25140 1705
rect 25110 1680 25115 1700
rect 25115 1680 25135 1700
rect 25135 1680 25140 1700
rect 25110 1675 25140 1680
rect 25310 1700 25340 1705
rect 25310 1680 25315 1700
rect 25315 1680 25335 1700
rect 25335 1680 25340 1700
rect 25310 1675 25340 1680
rect 25510 1700 25540 1705
rect 25510 1680 25515 1700
rect 25515 1680 25535 1700
rect 25535 1680 25540 1700
rect 25510 1675 25540 1680
rect 18935 1640 18970 1645
rect 18935 1615 18940 1640
rect 18940 1615 18965 1640
rect 18965 1615 18970 1640
rect 18935 1610 18970 1615
rect 18995 1640 19030 1645
rect 18995 1615 19000 1640
rect 19000 1615 19025 1640
rect 19025 1615 19030 1640
rect 18995 1610 19030 1615
rect 24820 1640 24855 1645
rect 24820 1615 24825 1640
rect 24825 1615 24850 1640
rect 24850 1615 24855 1640
rect 24820 1610 24855 1615
rect 24880 1640 24915 1645
rect 24880 1615 24885 1640
rect 24885 1615 24910 1640
rect 24910 1615 24915 1640
rect 24880 1610 24915 1615
rect 18080 1360 18110 1390
rect 25740 1360 25770 1390
rect 18410 930 18440 935
rect 18410 910 18415 930
rect 18415 910 18435 930
rect 18435 910 18440 930
rect 18410 905 18440 910
rect 18610 930 18640 935
rect 18610 910 18615 930
rect 18615 910 18635 930
rect 18635 910 18640 930
rect 18610 905 18640 910
rect 25210 930 25240 935
rect 25210 910 25215 930
rect 25215 910 25235 930
rect 25235 910 25240 930
rect 25210 905 25240 910
rect 25410 930 25440 935
rect 25410 910 25415 930
rect 25415 910 25435 930
rect 25435 910 25440 930
rect 25410 905 25440 910
rect 17965 830 17995 860
rect 15805 770 15835 800
rect 16310 795 16340 800
rect 16310 775 16315 795
rect 16315 775 16335 795
rect 16335 775 16340 795
rect 16310 770 16340 775
rect 16380 795 16410 800
rect 16380 775 16385 795
rect 16385 775 16405 795
rect 16405 775 16410 795
rect 16380 770 16410 775
rect 16450 795 16480 800
rect 16450 775 16455 795
rect 16455 775 16475 795
rect 16475 775 16480 795
rect 16450 770 16480 775
rect 17050 795 17080 800
rect 17050 775 17055 795
rect 17055 775 17075 795
rect 17075 775 17080 795
rect 17050 770 17080 775
rect 17270 795 17300 800
rect 17270 775 17275 795
rect 17275 775 17295 795
rect 17295 775 17300 795
rect 17270 770 17300 775
rect 17490 795 17520 800
rect 17490 775 17495 795
rect 17495 775 17515 795
rect 17515 775 17520 795
rect 17490 770 17520 775
rect 17910 770 17940 800
rect 2525 730 2555 760
rect 3135 755 3165 760
rect 3135 735 3140 755
rect 3140 735 3160 755
rect 3160 735 3165 755
rect 3135 730 3165 735
rect 3630 755 3660 760
rect 3630 735 3635 755
rect 3635 735 3655 755
rect 3655 735 3660 755
rect 3630 730 3660 735
rect 3990 755 4020 760
rect 3990 735 3995 755
rect 3995 735 4015 755
rect 4015 735 4020 755
rect 3990 730 4020 735
rect 4350 755 4380 760
rect 4350 735 4355 755
rect 4355 735 4375 755
rect 4375 735 4380 755
rect 4350 730 4380 735
rect 4530 755 4560 760
rect 4530 735 4535 755
rect 4535 735 4555 755
rect 4555 735 4560 755
rect 4530 730 4560 735
rect 4710 755 4740 760
rect 4710 735 4715 755
rect 4715 735 4735 755
rect 4735 735 4740 755
rect 4710 730 4740 735
rect 4890 755 4920 760
rect 4890 735 4895 755
rect 4895 735 4915 755
rect 4915 735 4920 755
rect 4890 730 4920 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 16995 675 17025 680
rect 16995 655 17000 675
rect 17000 655 17020 675
rect 17020 655 17025 675
rect 16995 650 17025 655
rect 17105 675 17135 680
rect 17105 655 17110 675
rect 17110 655 17130 675
rect 17130 655 17135 675
rect 17105 650 17135 655
rect 17215 675 17245 680
rect 17215 655 17220 675
rect 17220 655 17240 675
rect 17240 655 17245 675
rect 17215 650 17245 655
rect 17325 675 17355 680
rect 17325 655 17330 675
rect 17330 655 17350 675
rect 17350 655 17355 675
rect 17325 650 17355 655
rect 17435 675 17465 680
rect 17435 655 17440 675
rect 17440 655 17460 675
rect 17460 655 17465 675
rect 17435 650 17465 655
rect 27975 3795 28005 3825
rect 27920 3750 27950 3780
rect 27875 2295 27905 2325
rect 26445 2250 26475 2280
rect 26665 2250 26695 2280
rect 26885 2250 26915 2280
rect 27105 2250 27135 2280
rect 27325 2250 27355 2280
rect 26335 2205 26365 2235
rect 26555 2205 26585 2235
rect 26775 2205 26805 2235
rect 26995 2205 27025 2235
rect 27215 2205 27245 2235
rect 27435 2205 27465 2235
rect 26831 2175 26859 2180
rect 26831 2155 26836 2175
rect 26836 2155 26854 2175
rect 26854 2155 26859 2175
rect 26831 2150 26859 2155
rect 26390 1955 26420 1960
rect 26390 1935 26395 1955
rect 26395 1935 26415 1955
rect 26415 1935 26420 1955
rect 26390 1930 26420 1935
rect 26610 1955 26640 1960
rect 26610 1935 26615 1955
rect 26615 1935 26635 1955
rect 26635 1935 26640 1955
rect 26610 1930 26640 1935
rect 26830 1955 26860 1960
rect 26830 1935 26835 1955
rect 26835 1935 26855 1955
rect 26855 1935 26860 1955
rect 26830 1930 26860 1935
rect 27050 1955 27080 1960
rect 27050 1935 27055 1955
rect 27055 1935 27075 1955
rect 27075 1935 27080 1955
rect 27050 1930 27080 1935
rect 27270 1955 27300 1960
rect 27270 1935 27275 1955
rect 27275 1935 27295 1955
rect 27295 1935 27300 1955
rect 27270 1930 27300 1935
rect 26005 1865 26035 1895
rect 26500 1875 26530 1905
rect 26720 1875 26750 1905
rect 26940 1875 26970 1905
rect 27160 1875 27190 1905
rect 26195 1820 26225 1850
rect 26415 1820 26445 1850
rect 26090 1755 26120 1760
rect 26090 1735 26095 1755
rect 26095 1735 26115 1755
rect 26115 1735 26120 1755
rect 26090 1730 26120 1735
rect 26310 1755 26340 1760
rect 26310 1735 26315 1755
rect 26315 1735 26335 1755
rect 26335 1735 26340 1755
rect 26310 1730 26340 1735
rect 27380 1875 27410 1905
rect 26645 1820 26675 1850
rect 27235 1820 27265 1850
rect 27455 1820 27485 1850
rect 27685 1820 27715 1850
rect 27875 1845 27905 1875
rect 26825 1775 26855 1805
rect 26945 1775 26975 1805
rect 26530 1755 26560 1760
rect 26530 1735 26535 1755
rect 26535 1735 26555 1755
rect 26555 1735 26560 1755
rect 26530 1730 26560 1735
rect 27130 1755 27160 1760
rect 27130 1735 27135 1755
rect 27135 1735 27155 1755
rect 27155 1735 27160 1755
rect 27130 1730 27160 1735
rect 27350 1755 27380 1760
rect 27350 1735 27355 1755
rect 27355 1735 27375 1755
rect 27375 1735 27380 1755
rect 27350 1730 27380 1735
rect 27570 1755 27600 1760
rect 27570 1735 27575 1755
rect 27575 1735 27595 1755
rect 27595 1735 27600 1755
rect 27570 1730 27600 1735
rect 26240 1710 26266 1715
rect 26240 1690 26243 1710
rect 26243 1690 26260 1710
rect 26260 1690 26266 1710
rect 26240 1685 26266 1690
rect 26460 1710 26486 1715
rect 26460 1690 26463 1710
rect 26463 1690 26480 1710
rect 26480 1690 26486 1710
rect 26460 1685 26486 1690
rect 26604 1710 26630 1715
rect 26604 1690 26610 1710
rect 26610 1690 26627 1710
rect 26627 1690 26630 1710
rect 26604 1685 26630 1690
rect 26870 1710 26896 1715
rect 26870 1690 26876 1710
rect 26876 1690 26893 1710
rect 26893 1690 26896 1710
rect 26870 1685 26896 1690
rect 27280 1710 27306 1715
rect 27280 1690 27283 1710
rect 27283 1690 27300 1710
rect 27300 1690 27306 1710
rect 27280 1685 27306 1690
rect 27500 1710 27526 1715
rect 27500 1690 27503 1710
rect 27503 1690 27520 1710
rect 27520 1690 27526 1710
rect 27500 1685 27526 1690
rect 27644 1710 27670 1715
rect 27644 1690 27650 1710
rect 27650 1690 27667 1710
rect 27667 1690 27670 1710
rect 27644 1685 27670 1690
rect 26109 1490 26135 1495
rect 26109 1470 26112 1490
rect 26112 1470 26129 1490
rect 26129 1470 26135 1490
rect 26109 1465 26135 1470
rect 26310 1490 26340 1495
rect 26310 1470 26315 1490
rect 26315 1470 26335 1490
rect 26335 1470 26340 1490
rect 26310 1465 26340 1470
rect 26530 1490 26560 1495
rect 26530 1470 26535 1490
rect 26535 1470 26555 1490
rect 26555 1470 26560 1490
rect 26530 1465 26560 1470
rect 26925 1490 26951 1495
rect 26925 1470 26928 1490
rect 26928 1470 26945 1490
rect 26945 1470 26951 1490
rect 26925 1465 26951 1470
rect 27149 1490 27175 1495
rect 27149 1470 27152 1490
rect 27152 1470 27169 1490
rect 27169 1470 27175 1490
rect 27149 1465 27175 1470
rect 27350 1490 27380 1495
rect 27350 1470 27355 1490
rect 27355 1470 27375 1490
rect 27375 1470 27380 1490
rect 27350 1465 27380 1470
rect 27570 1490 27600 1495
rect 27570 1470 27575 1490
rect 27575 1470 27595 1490
rect 27595 1470 27600 1490
rect 27570 1465 27600 1470
rect 26150 1430 26180 1435
rect 26150 1410 26155 1430
rect 26155 1410 26175 1430
rect 26175 1410 26180 1430
rect 26150 1405 26180 1410
rect 26255 1430 26285 1435
rect 26255 1410 26260 1430
rect 26260 1410 26280 1430
rect 26280 1410 26285 1430
rect 26255 1405 26285 1410
rect 26365 1430 26395 1435
rect 26365 1410 26370 1430
rect 26370 1410 26390 1430
rect 26390 1410 26395 1430
rect 26365 1405 26395 1410
rect 26475 1430 26505 1435
rect 26475 1410 26480 1430
rect 26480 1410 26500 1430
rect 26500 1410 26505 1430
rect 26475 1405 26505 1410
rect 26585 1430 26615 1435
rect 26585 1410 26590 1430
rect 26590 1410 26610 1430
rect 26610 1410 26615 1430
rect 26585 1405 26615 1410
rect 26010 1215 26040 1245
rect 26815 1215 26845 1245
rect 26320 1165 26350 1195
rect 27190 1430 27220 1435
rect 27190 1410 27195 1430
rect 27195 1410 27215 1430
rect 27215 1410 27220 1430
rect 27190 1405 27220 1410
rect 27295 1430 27325 1435
rect 27295 1410 27300 1430
rect 27300 1410 27320 1430
rect 27320 1410 27325 1430
rect 27295 1405 27325 1410
rect 27405 1430 27435 1435
rect 27405 1410 27410 1430
rect 27410 1410 27430 1430
rect 27430 1410 27435 1430
rect 27405 1405 27435 1410
rect 27515 1430 27545 1435
rect 27515 1410 27520 1430
rect 27520 1410 27540 1430
rect 27540 1410 27545 1430
rect 27515 1405 27545 1410
rect 27625 1430 27655 1435
rect 27625 1410 27630 1430
rect 27630 1410 27650 1430
rect 27650 1410 27655 1430
rect 27625 1405 27655 1410
rect 26885 1165 26915 1195
rect 26430 1130 26460 1135
rect 26430 1110 26435 1130
rect 26435 1110 26455 1130
rect 26455 1110 26460 1130
rect 26430 1105 26460 1110
rect 26540 1130 26570 1135
rect 26540 1110 26545 1130
rect 26545 1110 26565 1130
rect 26565 1110 26570 1130
rect 26540 1105 26570 1110
rect 26650 1130 26680 1135
rect 26650 1110 26655 1130
rect 26655 1110 26675 1130
rect 26675 1110 26680 1130
rect 26650 1105 26680 1110
rect 26760 1130 26790 1135
rect 26760 1110 26765 1130
rect 26765 1110 26785 1130
rect 26785 1110 26790 1130
rect 26760 1105 26790 1110
rect 26870 1130 26900 1135
rect 26870 1110 26875 1130
rect 26875 1110 26895 1130
rect 26895 1110 26900 1130
rect 26870 1105 26900 1110
rect 26980 1130 27010 1135
rect 26980 1110 26985 1130
rect 26985 1110 27005 1130
rect 27005 1110 27010 1130
rect 26980 1105 27010 1110
rect 27090 1130 27120 1135
rect 27090 1110 27095 1130
rect 27095 1110 27115 1130
rect 27115 1110 27120 1130
rect 27090 1105 27120 1110
rect 27200 1130 27230 1135
rect 27200 1110 27205 1130
rect 27205 1110 27225 1130
rect 27225 1110 27230 1130
rect 27200 1105 27230 1110
rect 27310 1130 27340 1135
rect 27310 1110 27315 1130
rect 27315 1110 27335 1130
rect 27335 1110 27340 1130
rect 27310 1105 27340 1110
rect 27420 1130 27450 1135
rect 27420 1110 27425 1130
rect 27425 1110 27445 1130
rect 27445 1110 27450 1130
rect 27420 1105 27450 1110
rect 27530 1130 27560 1135
rect 27530 1110 27535 1130
rect 27535 1110 27555 1130
rect 27555 1110 27560 1130
rect 27530 1105 27560 1110
rect 27600 1145 27630 1150
rect 27600 1125 27605 1145
rect 27605 1125 27625 1145
rect 27625 1125 27630 1145
rect 27600 1120 27630 1125
rect 27920 1120 27950 1150
rect 26200 810 26230 815
rect 26200 790 26205 810
rect 26205 790 26225 810
rect 26225 790 26230 810
rect 26200 785 26230 790
rect 26265 810 26295 815
rect 26265 790 26270 810
rect 26270 790 26290 810
rect 26290 790 26295 810
rect 26265 785 26295 790
rect 26375 810 26405 815
rect 26375 790 26380 810
rect 26380 790 26400 810
rect 26400 790 26405 810
rect 26375 785 26405 790
rect 26485 810 26515 815
rect 26485 790 26490 810
rect 26490 790 26510 810
rect 26510 790 26515 810
rect 26485 785 26515 790
rect 26595 810 26625 815
rect 26595 790 26600 810
rect 26600 790 26620 810
rect 26620 790 26625 810
rect 26595 785 26625 790
rect 26705 810 26735 815
rect 26705 790 26710 810
rect 26710 790 26730 810
rect 26730 790 26735 810
rect 26705 785 26735 790
rect 26815 810 26845 815
rect 26815 790 26820 810
rect 26820 790 26840 810
rect 26840 790 26845 810
rect 26815 785 26845 790
rect 26925 810 26955 815
rect 26925 790 26930 810
rect 26930 790 26950 810
rect 26950 790 26955 810
rect 26925 785 26955 790
rect 27035 810 27065 815
rect 27035 790 27040 810
rect 27040 790 27060 810
rect 27060 790 27065 810
rect 27035 785 27065 790
rect 27145 810 27175 815
rect 27145 790 27150 810
rect 27150 790 27170 810
rect 27170 790 27175 810
rect 27145 785 27175 790
rect 27255 810 27285 815
rect 27255 790 27260 810
rect 27260 790 27280 810
rect 27280 790 27285 810
rect 27255 785 27285 790
rect 27365 810 27395 815
rect 27365 790 27370 810
rect 27370 790 27390 810
rect 27390 790 27395 810
rect 27365 785 27395 790
rect 27475 810 27505 815
rect 27475 790 27480 810
rect 27480 790 27500 810
rect 27500 790 27505 810
rect 27475 785 27505 790
rect 27590 810 27620 815
rect 27590 790 27595 810
rect 27595 790 27615 810
rect 27615 790 27620 810
rect 27590 785 27620 790
rect 26010 625 26040 655
rect 26510 625 26540 655
rect 26940 630 26970 660
rect 27160 630 27190 660
rect 27380 630 27410 660
rect 28205 3710 28235 3715
rect 28205 3690 28210 3710
rect 28210 3690 28230 3710
rect 28230 3690 28235 3710
rect 28205 3685 28235 3690
rect 28315 3710 28345 3715
rect 28315 3690 28320 3710
rect 28320 3690 28340 3710
rect 28340 3690 28345 3710
rect 28315 3685 28345 3690
rect 28425 3710 28455 3715
rect 28425 3690 28430 3710
rect 28430 3690 28450 3710
rect 28450 3690 28455 3710
rect 28425 3685 28455 3690
rect 28535 3710 28565 3715
rect 28535 3690 28540 3710
rect 28540 3690 28560 3710
rect 28560 3690 28565 3710
rect 28535 3685 28565 3690
rect 28645 3710 28675 3715
rect 28645 3690 28650 3710
rect 28650 3690 28670 3710
rect 28670 3690 28675 3710
rect 28645 3685 28675 3690
rect 28755 3710 28785 3715
rect 28755 3690 28760 3710
rect 28760 3690 28780 3710
rect 28780 3690 28785 3710
rect 28755 3685 28785 3690
rect 29160 3705 29190 3735
rect 29110 3625 29140 3655
rect 29160 3625 29190 3655
rect 29210 3625 29240 3655
rect 28260 3040 28290 3045
rect 28260 3020 28265 3040
rect 28265 3020 28285 3040
rect 28285 3020 28290 3040
rect 28260 3015 28290 3020
rect 28370 3040 28400 3045
rect 28370 3020 28375 3040
rect 28375 3020 28395 3040
rect 28395 3020 28400 3040
rect 28370 3015 28400 3020
rect 28480 3040 28510 3045
rect 28480 3020 28485 3040
rect 28485 3020 28505 3040
rect 28505 3020 28510 3040
rect 28480 3015 28510 3020
rect 28590 3040 28620 3045
rect 28590 3020 28595 3040
rect 28595 3020 28615 3040
rect 28615 3020 28620 3040
rect 28590 3015 28620 3020
rect 28700 3040 28730 3045
rect 28700 3020 28705 3040
rect 28705 3020 28725 3040
rect 28725 3020 28730 3040
rect 28700 3015 28730 3020
rect 28020 2850 28050 2880
rect 28315 2850 28345 2880
rect 29110 3005 29140 3035
rect 29160 3005 29190 3035
rect 29210 3005 29240 3035
rect 29160 2850 29190 2880
rect 28590 2805 28620 2835
rect 29400 2805 29430 2835
rect 28205 2750 28235 2755
rect 28205 2730 28210 2750
rect 28210 2730 28230 2750
rect 28230 2730 28235 2750
rect 28205 2725 28235 2730
rect 28315 2750 28345 2755
rect 28315 2730 28320 2750
rect 28320 2730 28340 2750
rect 28340 2730 28345 2750
rect 28315 2725 28345 2730
rect 28425 2750 28455 2755
rect 28425 2730 28430 2750
rect 28430 2730 28450 2750
rect 28450 2730 28455 2750
rect 28425 2725 28455 2730
rect 28535 2750 28565 2755
rect 28535 2730 28540 2750
rect 28540 2730 28560 2750
rect 28560 2730 28565 2750
rect 28535 2725 28565 2730
rect 28645 2750 28675 2755
rect 28645 2730 28650 2750
rect 28650 2730 28670 2750
rect 28670 2730 28675 2750
rect 28645 2725 28675 2730
rect 28755 2750 28785 2755
rect 28755 2730 28760 2750
rect 28760 2730 28780 2750
rect 28780 2730 28785 2750
rect 28755 2725 28785 2730
rect 28260 2480 28290 2485
rect 28260 2460 28265 2480
rect 28265 2460 28285 2480
rect 28285 2460 28290 2480
rect 28260 2455 28290 2460
rect 28370 2480 28400 2485
rect 28370 2460 28375 2480
rect 28375 2460 28395 2480
rect 28395 2460 28400 2480
rect 28370 2455 28400 2460
rect 28480 2480 28510 2485
rect 28480 2460 28485 2480
rect 28485 2460 28505 2480
rect 28505 2460 28510 2480
rect 28480 2455 28510 2460
rect 28590 2480 28620 2485
rect 28590 2460 28595 2480
rect 28595 2460 28615 2480
rect 28615 2460 28620 2480
rect 28590 2455 28620 2460
rect 28700 2480 28730 2485
rect 28700 2460 28705 2480
rect 28705 2460 28725 2480
rect 28725 2460 28730 2480
rect 28700 2455 28730 2460
rect 28945 2455 28975 2485
rect 28020 2345 28050 2375
rect 28315 2345 28345 2375
rect 28260 2290 28290 2295
rect 28260 2270 28265 2290
rect 28265 2270 28285 2290
rect 28285 2270 28290 2290
rect 28260 2265 28290 2270
rect 28370 2290 28400 2295
rect 28370 2270 28375 2290
rect 28375 2270 28395 2290
rect 28395 2270 28400 2290
rect 28370 2265 28400 2270
rect 28480 2290 28510 2295
rect 28480 2270 28485 2290
rect 28485 2270 28505 2290
rect 28505 2270 28510 2290
rect 28480 2265 28510 2270
rect 28590 2290 28620 2295
rect 28590 2270 28595 2290
rect 28595 2270 28615 2290
rect 28615 2270 28620 2290
rect 28590 2265 28620 2270
rect 28700 2290 28730 2295
rect 28700 2270 28705 2290
rect 28705 2270 28725 2290
rect 28725 2270 28730 2290
rect 28700 2265 28730 2270
rect 28900 2265 28930 2295
rect 29400 2080 29430 2110
rect 28945 1950 28975 1980
rect 29065 1980 29100 1985
rect 29065 1955 29070 1980
rect 29070 1955 29095 1980
rect 29095 1955 29100 1980
rect 29065 1950 29100 1955
rect 29125 1980 29160 1985
rect 29125 1955 29130 1980
rect 29130 1955 29155 1980
rect 29155 1955 29160 1980
rect 29125 1950 29160 1955
rect 29185 1980 29220 1985
rect 29185 1955 29190 1980
rect 29190 1955 29215 1980
rect 29215 1955 29220 1980
rect 29185 1950 29220 1955
rect 29245 1980 29280 1985
rect 29245 1955 29250 1980
rect 29250 1955 29275 1980
rect 29275 1955 29280 1980
rect 29245 1950 29280 1955
rect 28205 1920 28235 1925
rect 28205 1900 28212 1920
rect 28212 1900 28230 1920
rect 28230 1900 28235 1920
rect 28205 1895 28235 1900
rect 28315 1920 28345 1925
rect 28315 1900 28322 1920
rect 28322 1900 28340 1920
rect 28340 1900 28345 1920
rect 28315 1895 28345 1900
rect 28425 1920 28455 1925
rect 28425 1900 28432 1920
rect 28432 1900 28450 1920
rect 28450 1900 28455 1920
rect 28425 1895 28455 1900
rect 28535 1920 28565 1925
rect 28535 1900 28542 1920
rect 28542 1900 28560 1920
rect 28560 1900 28565 1920
rect 28535 1895 28565 1900
rect 28645 1920 28675 1925
rect 28645 1900 28652 1920
rect 28652 1900 28670 1920
rect 28670 1900 28675 1920
rect 28645 1895 28675 1900
rect 28755 1920 28785 1925
rect 28755 1900 28762 1920
rect 28762 1900 28780 1920
rect 28780 1900 28785 1920
rect 28755 1895 28785 1900
rect 28900 1895 28930 1925
rect 29125 1895 29155 1925
rect 29245 1845 29275 1875
rect 28030 1730 28060 1760
rect 28410 1730 28440 1760
rect 29120 1730 29150 1760
rect 28310 1700 28340 1705
rect 28310 1680 28315 1700
rect 28315 1680 28335 1700
rect 28335 1680 28340 1700
rect 28310 1675 28340 1680
rect 28510 1700 28540 1705
rect 28510 1680 28515 1700
rect 28515 1680 28535 1700
rect 28535 1680 28540 1700
rect 28510 1675 28540 1680
rect 28710 1700 28740 1705
rect 28710 1680 28715 1700
rect 28715 1680 28735 1700
rect 28735 1680 28740 1700
rect 28710 1675 28740 1680
rect 29055 1675 29085 1705
rect 29400 1675 29430 1705
rect 29055 1640 29090 1645
rect 29055 1615 29060 1640
rect 29060 1615 29085 1640
rect 29085 1615 29090 1640
rect 29055 1610 29090 1615
rect 29115 1640 29150 1645
rect 29115 1615 29120 1640
rect 29120 1615 29145 1640
rect 29145 1615 29150 1640
rect 29115 1610 29150 1615
rect 28030 1360 28060 1390
rect 28410 930 28440 935
rect 28410 910 28415 930
rect 28415 910 28435 930
rect 28435 910 28440 930
rect 28410 905 28440 910
rect 28610 930 28640 935
rect 28610 910 28615 930
rect 28615 910 28635 930
rect 28635 910 28640 930
rect 28610 905 28640 910
rect 27975 630 28005 660
rect 25805 570 25835 600
rect 26310 595 26340 600
rect 26310 575 26315 595
rect 26315 575 26335 595
rect 26335 575 26340 595
rect 26310 570 26340 575
rect 26380 595 26410 600
rect 26380 575 26385 595
rect 26385 575 26405 595
rect 26405 575 26410 595
rect 26380 570 26410 575
rect 26450 595 26480 600
rect 26450 575 26455 595
rect 26455 575 26475 595
rect 26475 575 26480 595
rect 26450 570 26480 575
rect 27050 595 27080 600
rect 27050 575 27055 595
rect 27055 575 27075 595
rect 27075 575 27080 595
rect 27050 570 27080 575
rect 27270 595 27300 600
rect 27270 575 27275 595
rect 27275 575 27295 595
rect 27295 575 27300 595
rect 27270 570 27300 575
rect 27490 595 27520 600
rect 27490 575 27495 595
rect 27495 575 27515 595
rect 27515 575 27520 595
rect 27490 570 27520 575
rect 27920 570 27950 600
rect 26995 475 27025 480
rect 26995 455 27000 475
rect 27000 455 27020 475
rect 27020 455 27025 475
rect 26995 450 27025 455
rect 27105 475 27135 480
rect 27105 455 27110 475
rect 27110 455 27130 475
rect 27130 455 27135 475
rect 27105 450 27135 455
rect 27215 475 27245 480
rect 27215 455 27220 475
rect 27220 455 27240 475
rect 27240 455 27245 475
rect 27215 450 27245 455
rect 27325 475 27355 480
rect 27325 455 27330 475
rect 27330 455 27350 475
rect 27350 455 27355 475
rect 27325 450 27355 455
rect 27435 475 27465 480
rect 27435 455 27440 475
rect 27440 455 27460 475
rect 27460 455 27465 475
rect 27435 450 27465 455
<< metal2 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect 26565 4985 26605 4990
rect 26565 4955 26570 4985
rect 26600 4980 26605 4985
rect 26685 4985 26725 4990
rect 26685 4980 26690 4985
rect 26600 4960 26690 4980
rect 26600 4955 26605 4960
rect 26565 4950 26605 4955
rect 26685 4955 26690 4960
rect 26720 4980 26725 4985
rect 26805 4985 26845 4990
rect 26805 4980 26810 4985
rect 26720 4960 26810 4980
rect 26720 4955 26725 4960
rect 26685 4950 26725 4955
rect 26805 4955 26810 4960
rect 26840 4970 26845 4985
rect 27235 4970 27275 4975
rect 26840 4955 27240 4970
rect 26805 4950 27240 4955
rect 27235 4940 27240 4950
rect 27270 4940 27275 4970
rect 27235 4935 27275 4940
rect 26505 4925 26545 4930
rect 26505 4895 26510 4925
rect 26540 4920 26545 4925
rect 26625 4925 26665 4930
rect 26625 4920 26630 4925
rect 26540 4900 26630 4920
rect 26540 4895 26545 4900
rect 26505 4890 26545 4895
rect 26625 4895 26630 4900
rect 26660 4920 26665 4925
rect 26745 4925 26785 4930
rect 26745 4920 26750 4925
rect 26660 4900 26750 4920
rect 26660 4895 26665 4900
rect 26625 4890 26665 4895
rect 26745 4895 26750 4900
rect 26780 4920 26785 4925
rect 26865 4925 26905 4930
rect 26865 4920 26870 4925
rect 26780 4900 26870 4920
rect 26780 4895 26785 4900
rect 26745 4890 26785 4895
rect 26865 4895 26870 4900
rect 26900 4895 26905 4925
rect 26865 4890 26905 4895
rect 27235 4900 27275 4905
rect 27235 4870 27240 4900
rect 27270 4895 27275 4900
rect 27355 4900 27395 4905
rect 27355 4895 27360 4900
rect 27270 4875 27360 4895
rect 27270 4870 27275 4875
rect 27235 4865 27275 4870
rect 27355 4870 27360 4875
rect 27390 4895 27395 4900
rect 27475 4900 27515 4905
rect 27475 4895 27480 4900
rect 27390 4875 27480 4895
rect 27390 4870 27395 4875
rect 27355 4865 27395 4870
rect 27475 4870 27480 4875
rect 27510 4895 27515 4900
rect 27595 4900 27635 4905
rect 27595 4895 27600 4900
rect 27510 4875 27600 4895
rect 27510 4870 27515 4875
rect 27475 4865 27515 4870
rect 27595 4870 27600 4875
rect 27630 4895 27635 4900
rect 27715 4900 27755 4905
rect 27715 4895 27720 4900
rect 27630 4875 27720 4895
rect 27630 4870 27635 4875
rect 27595 4865 27635 4870
rect 27715 4870 27720 4875
rect 27750 4870 27755 4900
rect 27715 4865 27755 4870
rect 26050 4770 26090 4775
rect 26050 4740 26055 4770
rect 26085 4765 26090 4770
rect 26685 4770 26725 4775
rect 26685 4765 26690 4770
rect 26085 4745 26690 4765
rect 26085 4740 26090 4745
rect 26050 4735 26090 4740
rect 26685 4740 26690 4745
rect 26720 4765 26725 4770
rect 27295 4770 27335 4775
rect 27295 4765 27300 4770
rect 26720 4745 27300 4765
rect 26720 4740 26725 4745
rect 26685 4735 26725 4740
rect 27295 4740 27300 4745
rect 27330 4765 27335 4770
rect 27415 4770 27455 4775
rect 27415 4765 27420 4770
rect 27330 4745 27420 4765
rect 27330 4740 27335 4745
rect 27295 4735 27335 4740
rect 27415 4740 27420 4745
rect 27450 4765 27455 4770
rect 27535 4770 27575 4775
rect 27535 4765 27540 4770
rect 27450 4745 27540 4765
rect 27450 4740 27455 4745
rect 27415 4735 27455 4740
rect 27535 4740 27540 4745
rect 27570 4765 27575 4770
rect 27655 4770 27695 4775
rect 27655 4765 27660 4770
rect 27570 4745 27660 4765
rect 27570 4740 27575 4745
rect 27535 4735 27575 4740
rect 27655 4740 27660 4745
rect 27690 4740 27695 4770
rect 27655 4735 27695 4740
rect 26105 4585 26145 4590
rect 26105 4555 26110 4585
rect 26140 4580 26145 4585
rect 26345 4585 26385 4590
rect 26345 4580 26350 4585
rect 26140 4560 26350 4580
rect 26140 4555 26145 4560
rect 26105 4550 26145 4555
rect 26345 4555 26350 4560
rect 26380 4580 26385 4585
rect 27355 4585 27395 4590
rect 27355 4580 27360 4585
rect 26380 4560 27360 4580
rect 26380 4555 26385 4560
rect 26345 4550 26385 4555
rect 27355 4555 27360 4560
rect 27390 4555 27395 4585
rect 27355 4550 27395 4555
rect 26360 4480 26400 4485
rect 16597 4465 16633 4470
rect 16597 4435 16600 4465
rect 16630 4460 16633 4465
rect 16717 4465 16753 4470
rect 16717 4460 16720 4465
rect 16630 4440 16720 4460
rect 16630 4435 16633 4440
rect 16597 4430 16633 4435
rect 16717 4435 16720 4440
rect 16750 4460 16753 4465
rect 16837 4465 16873 4470
rect 16837 4460 16840 4465
rect 16750 4440 16840 4460
rect 16750 4435 16753 4440
rect 16717 4430 16753 4435
rect 16837 4435 16840 4440
rect 16870 4460 16873 4465
rect 17185 4465 17225 4470
rect 17185 4460 17190 4465
rect 16870 4440 17190 4460
rect 16870 4435 16873 4440
rect 16837 4430 16873 4435
rect 17185 4435 17190 4440
rect 17220 4435 17225 4465
rect 26360 4450 26365 4480
rect 26395 4475 26400 4480
rect 26470 4480 26510 4485
rect 26470 4475 26475 4480
rect 26395 4455 26475 4475
rect 26395 4450 26400 4455
rect 26360 4445 26400 4450
rect 26470 4450 26475 4455
rect 26505 4475 26510 4480
rect 26580 4480 26620 4485
rect 26580 4475 26585 4480
rect 26505 4455 26585 4475
rect 26505 4450 26510 4455
rect 26470 4445 26510 4450
rect 26580 4450 26585 4455
rect 26615 4475 26620 4480
rect 26690 4480 26730 4485
rect 26690 4475 26695 4480
rect 26615 4455 26695 4475
rect 26615 4450 26620 4455
rect 26580 4445 26620 4450
rect 26690 4450 26695 4455
rect 26725 4475 26730 4480
rect 26800 4480 26840 4485
rect 26800 4475 26805 4480
rect 26725 4455 26805 4475
rect 26725 4450 26730 4455
rect 26690 4445 26730 4450
rect 26800 4450 26805 4455
rect 26835 4475 26840 4480
rect 26910 4480 26950 4485
rect 26910 4475 26915 4480
rect 26835 4455 26915 4475
rect 26835 4450 26840 4455
rect 26800 4445 26840 4450
rect 26910 4450 26915 4455
rect 26945 4475 26950 4480
rect 27020 4480 27060 4485
rect 27020 4475 27025 4480
rect 26945 4455 27025 4475
rect 26945 4450 26950 4455
rect 26910 4445 26950 4450
rect 27020 4450 27025 4455
rect 27055 4475 27060 4480
rect 27130 4480 27170 4485
rect 27130 4475 27135 4480
rect 27055 4455 27135 4475
rect 27055 4450 27060 4455
rect 27020 4445 27060 4450
rect 27130 4450 27135 4455
rect 27165 4475 27170 4480
rect 27240 4480 27280 4485
rect 27240 4475 27245 4480
rect 27165 4455 27245 4475
rect 27165 4450 27170 4455
rect 27130 4445 27170 4450
rect 27240 4450 27245 4455
rect 27275 4475 27280 4480
rect 27350 4480 27390 4485
rect 27350 4475 27355 4480
rect 27275 4455 27355 4475
rect 27275 4450 27280 4455
rect 27240 4445 27280 4450
rect 27350 4450 27355 4455
rect 27385 4450 27390 4480
rect 27350 4445 27390 4450
rect 17185 4430 17225 4435
rect 16535 4420 16575 4425
rect 16535 4410 16540 4420
rect 16165 4405 16205 4410
rect 16165 4375 16170 4405
rect 16200 4375 16205 4405
rect 16165 4370 16205 4375
rect 16425 4405 16540 4410
rect 16425 4375 16430 4405
rect 16460 4390 16540 4405
rect 16570 4415 16575 4420
rect 16655 4420 16695 4425
rect 16655 4415 16660 4420
rect 16570 4395 16660 4415
rect 16570 4390 16575 4395
rect 16460 4375 16465 4390
rect 16535 4385 16575 4390
rect 16655 4390 16660 4395
rect 16690 4415 16695 4420
rect 16775 4420 16815 4425
rect 16775 4415 16780 4420
rect 16690 4395 16780 4415
rect 16690 4390 16695 4395
rect 16655 4385 16695 4390
rect 16775 4390 16780 4395
rect 16810 4415 16815 4420
rect 16895 4420 16935 4425
rect 16895 4415 16900 4420
rect 16810 4395 16900 4415
rect 16810 4390 16815 4395
rect 16775 4385 16815 4390
rect 16895 4390 16900 4395
rect 16930 4390 16935 4420
rect 16895 4385 16935 4390
rect 17185 4395 17225 4400
rect 16425 4370 16465 4375
rect 17185 4365 17190 4395
rect 17220 4390 17225 4395
rect 17305 4395 17345 4400
rect 17305 4390 17310 4395
rect 17220 4370 17310 4390
rect 17220 4365 17225 4370
rect 17185 4360 17225 4365
rect 17305 4365 17310 4370
rect 17340 4390 17345 4395
rect 17425 4395 17465 4400
rect 17425 4390 17430 4395
rect 17340 4370 17430 4390
rect 17340 4365 17345 4370
rect 17305 4360 17345 4365
rect 17425 4365 17430 4370
rect 17460 4390 17465 4395
rect 17545 4395 17585 4400
rect 17545 4390 17550 4395
rect 17460 4370 17550 4390
rect 17460 4365 17465 4370
rect 17425 4360 17465 4365
rect 17545 4365 17550 4370
rect 17580 4390 17585 4395
rect 17665 4395 17705 4400
rect 17665 4390 17670 4395
rect 17580 4370 17670 4390
rect 17580 4365 17585 4370
rect 17545 4360 17585 4365
rect 17665 4365 17670 4370
rect 17700 4365 17705 4395
rect 17665 4360 17705 4365
rect 26305 4360 26345 4365
rect 26305 4330 26310 4360
rect 26340 4355 26345 4360
rect 26525 4360 26565 4365
rect 26525 4355 26530 4360
rect 26340 4335 26530 4355
rect 26340 4330 26345 4335
rect 26305 4325 26345 4330
rect 26525 4330 26530 4335
rect 26560 4355 26565 4360
rect 26745 4360 26785 4365
rect 26745 4355 26750 4360
rect 26560 4335 26750 4355
rect 26560 4330 26565 4335
rect 26525 4325 26565 4330
rect 26745 4330 26750 4335
rect 26780 4355 26785 4360
rect 26965 4360 27005 4365
rect 26965 4355 26970 4360
rect 26780 4335 26970 4355
rect 26780 4330 26785 4335
rect 26745 4325 26785 4330
rect 26965 4330 26970 4335
rect 27000 4355 27005 4360
rect 27185 4360 27225 4365
rect 27185 4355 27190 4360
rect 27000 4335 27190 4355
rect 27000 4330 27005 4335
rect 26965 4325 27005 4330
rect 27185 4330 27190 4335
rect 27220 4355 27225 4360
rect 27405 4360 27445 4365
rect 27405 4355 27410 4360
rect 27220 4335 27410 4355
rect 27220 4330 27225 4335
rect 27185 4325 27225 4330
rect 27405 4330 27410 4335
rect 27440 4330 27445 4360
rect 27405 4325 27445 4330
rect 16050 4265 16090 4270
rect 16050 4235 16055 4265
rect 16085 4260 16090 4265
rect 16715 4265 16755 4270
rect 16715 4260 16720 4265
rect 16085 4240 16720 4260
rect 16085 4235 16090 4240
rect 16050 4230 16090 4235
rect 16715 4235 16720 4240
rect 16750 4260 16755 4265
rect 17245 4265 17285 4270
rect 17245 4260 17250 4265
rect 16750 4240 17250 4260
rect 16750 4235 16755 4240
rect 16715 4230 16755 4235
rect 17245 4235 17250 4240
rect 17280 4260 17285 4265
rect 17365 4265 17405 4270
rect 17365 4260 17370 4265
rect 17280 4240 17370 4260
rect 17280 4235 17285 4240
rect 17245 4230 17285 4235
rect 17365 4235 17370 4240
rect 17400 4260 17405 4265
rect 17485 4265 17525 4270
rect 17485 4260 17490 4265
rect 17400 4240 17490 4260
rect 17400 4235 17405 4240
rect 17365 4230 17405 4235
rect 17485 4235 17490 4240
rect 17520 4260 17525 4265
rect 17605 4265 17645 4270
rect 17605 4260 17610 4265
rect 17520 4240 17610 4260
rect 17520 4235 17525 4240
rect 17485 4230 17525 4235
rect 17605 4235 17610 4240
rect 17640 4235 17645 4265
rect 17605 4230 17645 4235
rect 26420 4245 26460 4250
rect 26420 4215 26425 4245
rect 26455 4240 26460 4245
rect 26635 4245 26675 4250
rect 26635 4240 26640 4245
rect 26455 4220 26640 4240
rect 26455 4215 26460 4220
rect 16105 4210 16145 4215
rect 16105 4180 16110 4210
rect 16140 4205 16145 4210
rect 16295 4210 16335 4215
rect 16295 4205 16300 4210
rect 16140 4185 16300 4205
rect 16140 4180 16145 4185
rect 16105 4175 16145 4180
rect 16295 4180 16300 4185
rect 16330 4205 16335 4210
rect 17305 4210 17345 4215
rect 26420 4210 26460 4215
rect 26635 4215 26640 4220
rect 26670 4240 26675 4245
rect 26855 4245 26895 4250
rect 26855 4240 26860 4245
rect 26670 4220 26860 4240
rect 26670 4215 26675 4220
rect 26635 4210 26675 4215
rect 26855 4215 26860 4220
rect 26890 4240 26895 4245
rect 27075 4245 27115 4250
rect 27075 4240 27080 4245
rect 26890 4220 27080 4240
rect 26890 4215 26895 4220
rect 26855 4210 26895 4215
rect 27075 4215 27080 4220
rect 27110 4240 27115 4245
rect 27295 4245 27335 4250
rect 27295 4240 27300 4245
rect 27110 4220 27300 4240
rect 27110 4215 27115 4220
rect 27075 4210 27115 4215
rect 27295 4215 27300 4220
rect 27330 4215 27335 4245
rect 27295 4210 27335 4215
rect 17305 4205 17310 4210
rect 16330 4185 17310 4205
rect 16330 4180 16335 4185
rect 16295 4175 16335 4180
rect 17305 4180 17310 4185
rect 17340 4180 17345 4210
rect 17305 4175 17345 4180
rect 16360 4155 16400 4160
rect 16360 4125 16365 4155
rect 16395 4150 16400 4155
rect 16470 4155 16510 4160
rect 16470 4150 16475 4155
rect 16395 4130 16475 4150
rect 16395 4125 16400 4130
rect 16360 4120 16400 4125
rect 16470 4125 16475 4130
rect 16505 4150 16510 4155
rect 16580 4155 16620 4160
rect 16580 4150 16585 4155
rect 16505 4130 16585 4150
rect 16505 4125 16510 4130
rect 16470 4120 16510 4125
rect 16580 4125 16585 4130
rect 16615 4150 16620 4155
rect 16690 4155 16730 4160
rect 16690 4150 16695 4155
rect 16615 4130 16695 4150
rect 16615 4125 16620 4130
rect 16580 4120 16620 4125
rect 16690 4125 16695 4130
rect 16725 4150 16730 4155
rect 16800 4155 16840 4160
rect 16800 4150 16805 4155
rect 16725 4130 16805 4150
rect 16725 4125 16730 4130
rect 16690 4120 16730 4125
rect 16800 4125 16805 4130
rect 16835 4150 16840 4155
rect 16910 4155 16950 4160
rect 16910 4150 16915 4155
rect 16835 4130 16915 4150
rect 16835 4125 16840 4130
rect 16800 4120 16840 4125
rect 16910 4125 16915 4130
rect 16945 4150 16950 4155
rect 17020 4155 17060 4160
rect 17020 4150 17025 4155
rect 16945 4130 17025 4150
rect 16945 4125 16950 4130
rect 16910 4120 16950 4125
rect 17020 4125 17025 4130
rect 17055 4150 17060 4155
rect 17130 4155 17170 4160
rect 17130 4150 17135 4155
rect 17055 4130 17135 4150
rect 17055 4125 17060 4130
rect 17020 4120 17060 4125
rect 17130 4125 17135 4130
rect 17165 4150 17170 4155
rect 17240 4155 17280 4160
rect 17240 4150 17245 4155
rect 17165 4130 17245 4150
rect 17165 4125 17170 4130
rect 17130 4120 17170 4125
rect 17240 4125 17245 4130
rect 17275 4150 17280 4155
rect 17350 4155 17390 4160
rect 17350 4150 17355 4155
rect 17275 4130 17355 4150
rect 17275 4125 17280 4130
rect 17240 4120 17280 4125
rect 17350 4125 17355 4130
rect 17385 4125 17390 4155
rect 17350 4120 17390 4125
rect 26320 4130 26360 4135
rect 26320 4100 26325 4130
rect 26355 4125 26360 4130
rect 26420 4130 26460 4135
rect 26420 4125 26425 4130
rect 26355 4105 26425 4125
rect 26355 4100 26360 4105
rect 26320 4095 26360 4100
rect 26420 4100 26425 4105
rect 26455 4125 26460 4130
rect 26530 4130 26570 4135
rect 26530 4125 26535 4130
rect 26455 4105 26535 4125
rect 26455 4100 26460 4105
rect 26420 4095 26460 4100
rect 26530 4100 26535 4105
rect 26565 4125 26570 4130
rect 26640 4130 26680 4135
rect 26640 4125 26645 4130
rect 26565 4105 26645 4125
rect 26565 4100 26570 4105
rect 26530 4095 26570 4100
rect 26640 4100 26645 4105
rect 26675 4125 26680 4130
rect 26750 4130 26790 4135
rect 26750 4125 26755 4130
rect 26675 4105 26755 4125
rect 26675 4100 26680 4105
rect 26640 4095 26680 4100
rect 26750 4100 26755 4105
rect 26785 4100 26790 4130
rect 26750 4095 26790 4100
rect 27050 4130 27090 4135
rect 27050 4100 27055 4130
rect 27085 4125 27090 4130
rect 27150 4130 27190 4135
rect 27150 4125 27155 4130
rect 27085 4105 27155 4125
rect 27085 4100 27090 4105
rect 27050 4095 27090 4100
rect 27150 4100 27155 4105
rect 27185 4125 27190 4130
rect 27260 4130 27300 4135
rect 27260 4125 27265 4130
rect 27185 4105 27265 4125
rect 27185 4100 27190 4105
rect 27150 4095 27190 4100
rect 27260 4100 27265 4105
rect 27295 4125 27300 4130
rect 27370 4130 27410 4135
rect 27370 4125 27375 4130
rect 27295 4105 27375 4125
rect 27295 4100 27300 4105
rect 27260 4095 27300 4100
rect 27370 4100 27375 4105
rect 27405 4125 27410 4130
rect 27480 4130 27520 4135
rect 27480 4125 27485 4130
rect 27405 4105 27485 4125
rect 27405 4100 27410 4105
rect 27370 4095 27410 4100
rect 27480 4100 27485 4105
rect 27515 4100 27520 4130
rect 27480 4095 27520 4100
rect 26280 4069 26310 4075
rect 26280 4041 26282 4069
rect 26308 4065 26310 4069
rect 26480 4069 26510 4075
rect 26480 4065 26482 4069
rect 26308 4045 26482 4065
rect 26308 4041 26310 4045
rect 16305 4035 16345 4040
rect 16305 4005 16310 4035
rect 16340 4030 16345 4035
rect 16525 4035 16565 4040
rect 16525 4030 16530 4035
rect 16340 4010 16530 4030
rect 16340 4005 16345 4010
rect 16305 4000 16345 4005
rect 16525 4005 16530 4010
rect 16560 4030 16565 4035
rect 16745 4035 16785 4040
rect 16745 4030 16750 4035
rect 16560 4010 16750 4030
rect 16560 4005 16565 4010
rect 16525 4000 16565 4005
rect 16745 4005 16750 4010
rect 16780 4030 16785 4035
rect 16965 4035 17005 4040
rect 16965 4030 16970 4035
rect 16780 4010 16970 4030
rect 16780 4005 16785 4010
rect 16745 4000 16785 4005
rect 16965 4005 16970 4010
rect 17000 4030 17005 4035
rect 17185 4035 17225 4040
rect 17185 4030 17190 4035
rect 17000 4010 17190 4030
rect 17000 4005 17005 4010
rect 16965 4000 17005 4005
rect 17185 4005 17190 4010
rect 17220 4030 17225 4035
rect 17405 4035 17445 4040
rect 26280 4035 26310 4041
rect 26480 4041 26482 4045
rect 26508 4065 26510 4069
rect 27008 4069 27038 4075
rect 27008 4065 27010 4069
rect 26508 4045 27010 4065
rect 26508 4041 26510 4045
rect 26480 4035 26510 4041
rect 27008 4041 27010 4045
rect 27036 4065 27038 4069
rect 27205 4070 27245 4075
rect 27205 4065 27210 4070
rect 27036 4045 27210 4065
rect 27036 4041 27038 4045
rect 27008 4035 27038 4041
rect 27205 4040 27210 4045
rect 27240 4065 27245 4070
rect 27425 4070 27465 4075
rect 27425 4065 27430 4070
rect 27240 4045 27430 4065
rect 27240 4040 27245 4045
rect 27205 4035 27245 4040
rect 27425 4040 27430 4045
rect 27460 4065 27465 4070
rect 27870 4070 27910 4075
rect 27870 4065 27875 4070
rect 27460 4045 27875 4065
rect 27460 4040 27465 4045
rect 27425 4035 27465 4040
rect 27870 4040 27875 4045
rect 27905 4040 27910 4070
rect 27870 4035 27910 4040
rect 17405 4030 17410 4035
rect 17220 4010 17410 4030
rect 17220 4005 17225 4010
rect 17185 4000 17225 4005
rect 17405 4005 17410 4010
rect 17440 4005 17445 4035
rect 17405 4000 17445 4005
rect 16415 3975 16455 3980
rect 16415 3945 16420 3975
rect 16450 3970 16455 3975
rect 16635 3975 16675 3980
rect 16635 3970 16640 3975
rect 16450 3950 16640 3970
rect 16450 3945 16455 3950
rect 16415 3940 16455 3945
rect 16635 3945 16640 3950
rect 16670 3970 16675 3975
rect 16855 3975 16895 3980
rect 16855 3970 16860 3975
rect 16670 3950 16860 3970
rect 16670 3945 16675 3950
rect 16635 3940 16675 3945
rect 16855 3945 16860 3950
rect 16890 3970 16895 3975
rect 17075 3975 17115 3980
rect 17075 3970 17080 3975
rect 16890 3950 17080 3970
rect 16890 3945 16895 3950
rect 16855 3940 16895 3945
rect 17075 3945 17080 3950
rect 17110 3970 17115 3975
rect 17295 3975 17335 3980
rect 17295 3970 17300 3975
rect 17110 3950 17300 3970
rect 17110 3945 17115 3950
rect 17075 3940 17115 3945
rect 17295 3945 17300 3950
rect 17330 3945 17335 3975
rect 26407 3950 26439 3955
rect 26407 3945 26410 3950
rect 17295 3940 17335 3945
rect 26185 3925 26410 3945
rect 26407 3920 26410 3925
rect 26436 3945 26439 3950
rect 26627 3950 26659 3955
rect 26627 3945 26630 3950
rect 26436 3925 26630 3945
rect 26436 3920 26439 3925
rect 26407 3915 26439 3920
rect 26627 3920 26630 3925
rect 26656 3945 26659 3950
rect 26771 3950 26803 3955
rect 26771 3945 26774 3950
rect 26656 3925 26774 3945
rect 26656 3920 26659 3925
rect 26627 3915 26659 3920
rect 26771 3920 26774 3925
rect 26800 3945 26803 3950
rect 27137 3950 27169 3955
rect 27137 3945 27140 3950
rect 26800 3925 27140 3945
rect 26800 3920 26803 3925
rect 26771 3915 26803 3920
rect 27137 3920 27140 3925
rect 27166 3945 27169 3950
rect 27357 3950 27389 3955
rect 27357 3945 27360 3950
rect 27166 3925 27360 3945
rect 27166 3920 27169 3925
rect 27137 3915 27169 3920
rect 27357 3920 27360 3925
rect 27386 3945 27389 3950
rect 27501 3950 27533 3955
rect 27501 3945 27504 3950
rect 27386 3925 27504 3945
rect 27386 3920 27389 3925
rect 27357 3915 27389 3920
rect 27501 3920 27504 3925
rect 27530 3920 27533 3950
rect 27501 3915 27533 3920
rect 16310 3910 16350 3915
rect 16310 3880 16315 3910
rect 16345 3905 16350 3910
rect 16415 3910 16455 3915
rect 16415 3905 16420 3910
rect 16345 3885 16420 3905
rect 16345 3880 16350 3885
rect 16310 3875 16350 3880
rect 16415 3880 16420 3885
rect 16450 3905 16455 3910
rect 16525 3910 16565 3915
rect 16525 3905 16530 3910
rect 16450 3885 16530 3905
rect 16450 3880 16455 3885
rect 16415 3875 16455 3880
rect 16525 3880 16530 3885
rect 16560 3905 16565 3910
rect 16635 3910 16675 3915
rect 16635 3905 16640 3910
rect 16560 3885 16640 3905
rect 16560 3880 16565 3885
rect 16525 3875 16565 3880
rect 16635 3880 16640 3885
rect 16670 3905 16675 3910
rect 16745 3910 16785 3915
rect 16745 3905 16750 3910
rect 16670 3885 16750 3905
rect 16670 3880 16675 3885
rect 16635 3875 16675 3880
rect 16745 3880 16750 3885
rect 16780 3880 16785 3910
rect 16745 3875 16785 3880
rect 17050 3910 17090 3915
rect 17050 3880 17055 3910
rect 17085 3905 17090 3910
rect 17155 3910 17195 3915
rect 17155 3905 17160 3910
rect 17085 3885 17160 3905
rect 17085 3880 17090 3885
rect 17050 3875 17090 3880
rect 17155 3880 17160 3885
rect 17190 3905 17195 3910
rect 17265 3910 17305 3915
rect 17265 3905 17270 3910
rect 17190 3885 17270 3905
rect 17190 3880 17195 3885
rect 17155 3875 17195 3880
rect 17265 3880 17270 3885
rect 17300 3905 17305 3910
rect 17375 3910 17415 3915
rect 17375 3905 17380 3910
rect 17300 3885 17380 3905
rect 17300 3880 17305 3885
rect 17265 3875 17305 3880
rect 17375 3880 17380 3885
rect 17410 3905 17415 3910
rect 17485 3910 17525 3915
rect 17485 3905 17490 3910
rect 17410 3885 17490 3905
rect 17410 3880 17415 3885
rect 17375 3875 17415 3880
rect 17485 3880 17490 3885
rect 17520 3880 17525 3910
rect 17485 3875 17525 3880
rect 26255 3890 26295 3895
rect 26255 3860 26260 3890
rect 26290 3885 26295 3890
rect 26360 3890 26400 3895
rect 26360 3885 26365 3890
rect 26290 3865 26365 3885
rect 26290 3860 26295 3865
rect 26255 3855 26295 3860
rect 26360 3860 26365 3865
rect 26395 3885 26400 3890
rect 26475 3890 26515 3895
rect 26475 3885 26480 3890
rect 26395 3865 26480 3885
rect 26395 3860 26400 3865
rect 26360 3855 26400 3860
rect 26475 3860 26480 3865
rect 26510 3885 26515 3890
rect 26580 3890 26620 3895
rect 26580 3885 26585 3890
rect 26510 3865 26585 3885
rect 26510 3860 26515 3865
rect 26475 3855 26515 3860
rect 26580 3860 26585 3865
rect 26615 3885 26620 3890
rect 26695 3890 26735 3895
rect 26695 3885 26700 3890
rect 26615 3865 26700 3885
rect 26615 3860 26620 3865
rect 26580 3855 26620 3860
rect 26695 3860 26700 3865
rect 26730 3885 26735 3890
rect 26810 3890 26850 3895
rect 26810 3885 26815 3890
rect 26730 3865 26815 3885
rect 26730 3860 26735 3865
rect 26695 3855 26735 3860
rect 26810 3860 26815 3865
rect 26845 3860 26850 3890
rect 26810 3855 26850 3860
rect 26985 3890 27025 3895
rect 26985 3860 26990 3890
rect 27020 3885 27025 3890
rect 27205 3890 27245 3895
rect 27205 3885 27210 3890
rect 27020 3865 27210 3885
rect 27020 3860 27025 3865
rect 26985 3855 27025 3860
rect 27205 3860 27210 3865
rect 27240 3885 27245 3890
rect 27425 3890 27465 3895
rect 27425 3885 27430 3890
rect 27240 3865 27430 3885
rect 27240 3860 27245 3865
rect 27205 3855 27245 3860
rect 27425 3860 27430 3865
rect 27460 3885 27465 3890
rect 27460 3865 27955 3885
rect 27460 3860 27465 3865
rect 27425 3855 27465 3860
rect 16271 3850 16303 3855
rect 16271 3820 16274 3850
rect 16300 3845 16303 3850
rect 16470 3850 16510 3855
rect 16470 3845 16475 3850
rect 16300 3825 16475 3845
rect 16300 3820 16303 3825
rect 16271 3815 16303 3820
rect 16470 3820 16475 3825
rect 16505 3845 16510 3850
rect 16690 3850 16730 3855
rect 16690 3845 16695 3850
rect 16505 3825 16695 3845
rect 16505 3820 16510 3825
rect 16470 3815 16510 3820
rect 16690 3820 16695 3825
rect 16725 3845 16730 3850
rect 17011 3850 17043 3855
rect 17011 3845 17014 3850
rect 16725 3825 17014 3845
rect 16725 3820 16730 3825
rect 16690 3815 16730 3820
rect 17011 3820 17014 3825
rect 17040 3845 17043 3850
rect 17210 3850 17250 3855
rect 17210 3845 17215 3850
rect 17040 3825 17215 3845
rect 17040 3820 17043 3825
rect 17011 3815 17043 3820
rect 17210 3820 17215 3825
rect 17245 3845 17250 3850
rect 17430 3850 17470 3855
rect 17430 3845 17435 3850
rect 17245 3825 17435 3845
rect 17245 3820 17250 3825
rect 17210 3815 17250 3820
rect 17430 3820 17435 3825
rect 17465 3845 17470 3850
rect 17860 3850 17900 3855
rect 17860 3845 17865 3850
rect 17465 3825 17865 3845
rect 17465 3820 17470 3825
rect 17430 3815 17470 3820
rect 17860 3820 17865 3825
rect 17895 3820 17900 3850
rect 27970 3825 28010 3830
rect 27970 3820 27975 3825
rect 17860 3815 17900 3820
rect 27955 3800 27975 3820
rect 27970 3795 27975 3800
rect 28005 3795 28010 3825
rect 27970 3790 28010 3795
rect 27090 3780 27130 3785
rect 27090 3750 27095 3780
rect 27125 3775 27130 3780
rect 27310 3780 27350 3785
rect 27310 3775 27315 3780
rect 27125 3755 27315 3775
rect 27125 3750 27130 3755
rect 27090 3745 27130 3750
rect 27310 3750 27315 3755
rect 27345 3775 27350 3780
rect 27540 3780 27580 3785
rect 27540 3775 27545 3780
rect 27345 3755 27545 3775
rect 27345 3750 27350 3755
rect 27310 3745 27350 3750
rect 27540 3750 27545 3755
rect 27575 3775 27580 3780
rect 27915 3780 27955 3785
rect 27915 3775 27920 3780
rect 27575 3755 27920 3775
rect 27575 3750 27580 3755
rect 27540 3745 27580 3750
rect 27915 3750 27920 3755
rect 27950 3750 27955 3780
rect 27915 3745 27955 3750
rect 29155 3735 29195 3740
rect 16402 3730 16434 3735
rect 16402 3725 16405 3730
rect 15915 3705 16405 3725
rect 16402 3700 16405 3705
rect 16431 3725 16434 3730
rect 16622 3730 16654 3735
rect 16622 3725 16625 3730
rect 16431 3705 16625 3725
rect 16431 3700 16434 3705
rect 16402 3695 16434 3700
rect 16622 3700 16625 3705
rect 16651 3725 16654 3730
rect 16766 3730 16798 3735
rect 16766 3725 16769 3730
rect 16651 3705 16769 3725
rect 16651 3700 16654 3705
rect 16622 3695 16654 3700
rect 16766 3700 16769 3705
rect 16795 3725 16798 3730
rect 17142 3730 17174 3735
rect 17142 3725 17145 3730
rect 16795 3705 17145 3725
rect 16795 3700 16798 3705
rect 16766 3695 16798 3700
rect 17142 3700 17145 3705
rect 17171 3725 17174 3730
rect 17362 3730 17394 3735
rect 17362 3725 17365 3730
rect 17171 3705 17365 3725
rect 17171 3700 17174 3705
rect 17142 3695 17174 3700
rect 17362 3700 17365 3705
rect 17391 3725 17394 3730
rect 17506 3730 17538 3735
rect 17506 3725 17509 3730
rect 17391 3705 17509 3725
rect 17391 3700 17394 3705
rect 17362 3695 17394 3700
rect 17506 3700 17509 3705
rect 17535 3700 17538 3730
rect 17506 3695 17538 3700
rect 28200 3715 28240 3720
rect 28200 3685 28205 3715
rect 28235 3710 28240 3715
rect 28310 3715 28350 3720
rect 28310 3710 28315 3715
rect 28235 3690 28315 3710
rect 28235 3685 28240 3690
rect 16990 3680 17030 3685
rect 16250 3670 16290 3675
rect 16250 3640 16255 3670
rect 16285 3665 16290 3670
rect 16355 3670 16395 3675
rect 16355 3665 16360 3670
rect 16285 3645 16360 3665
rect 16285 3640 16290 3645
rect 14605 3635 14645 3640
rect 14605 3605 14610 3635
rect 14640 3605 14645 3635
rect 14605 3600 14645 3605
rect 15060 3635 15100 3640
rect 15060 3605 15065 3635
rect 15095 3630 15100 3635
rect 15170 3635 15210 3640
rect 15170 3630 15175 3635
rect 15095 3610 15175 3630
rect 15095 3605 15100 3610
rect 15060 3600 15100 3605
rect 15170 3605 15175 3610
rect 15205 3630 15210 3635
rect 15280 3635 15320 3640
rect 15280 3630 15285 3635
rect 15205 3610 15285 3630
rect 15205 3605 15210 3610
rect 15170 3600 15210 3605
rect 15280 3605 15285 3610
rect 15315 3630 15320 3635
rect 15390 3635 15430 3640
rect 15390 3630 15395 3635
rect 15315 3610 15395 3630
rect 15315 3605 15320 3610
rect 15280 3600 15320 3605
rect 15390 3605 15395 3610
rect 15425 3630 15430 3635
rect 15500 3635 15540 3640
rect 15500 3630 15505 3635
rect 15425 3610 15505 3630
rect 15425 3605 15430 3610
rect 15390 3600 15430 3605
rect 15500 3605 15505 3610
rect 15535 3630 15540 3635
rect 15610 3635 15650 3640
rect 16250 3635 16290 3640
rect 16355 3640 16360 3645
rect 16390 3665 16395 3670
rect 16470 3670 16510 3675
rect 16470 3665 16475 3670
rect 16390 3645 16475 3665
rect 16390 3640 16395 3645
rect 16355 3635 16395 3640
rect 16470 3640 16475 3645
rect 16505 3665 16510 3670
rect 16575 3670 16615 3675
rect 16575 3665 16580 3670
rect 16505 3645 16580 3665
rect 16505 3640 16510 3645
rect 16470 3635 16510 3640
rect 16575 3640 16580 3645
rect 16610 3665 16615 3670
rect 16690 3670 16730 3675
rect 16690 3665 16695 3670
rect 16610 3645 16695 3665
rect 16610 3640 16615 3645
rect 16575 3635 16615 3640
rect 16690 3640 16695 3645
rect 16725 3665 16730 3670
rect 16805 3670 16845 3675
rect 16805 3665 16810 3670
rect 16725 3645 16810 3665
rect 16725 3640 16730 3645
rect 16690 3635 16730 3640
rect 16805 3640 16810 3645
rect 16840 3640 16845 3670
rect 16990 3650 16995 3680
rect 17025 3675 17030 3680
rect 17210 3680 17250 3685
rect 17210 3675 17215 3680
rect 17025 3655 17215 3675
rect 17025 3650 17030 3655
rect 16990 3645 17030 3650
rect 17210 3650 17215 3655
rect 17245 3675 17250 3680
rect 17430 3680 17470 3685
rect 17430 3675 17435 3680
rect 17245 3655 17435 3675
rect 17245 3650 17250 3655
rect 17210 3645 17250 3650
rect 17430 3650 17435 3655
rect 17465 3675 17470 3680
rect 17960 3680 18000 3685
rect 28200 3680 28240 3685
rect 28310 3685 28315 3690
rect 28345 3710 28350 3715
rect 28420 3715 28460 3720
rect 28420 3710 28425 3715
rect 28345 3690 28425 3710
rect 28345 3685 28350 3690
rect 28310 3680 28350 3685
rect 28420 3685 28425 3690
rect 28455 3710 28460 3715
rect 28530 3715 28570 3720
rect 28530 3710 28535 3715
rect 28455 3690 28535 3710
rect 28455 3685 28460 3690
rect 28420 3680 28460 3685
rect 28530 3685 28535 3690
rect 28565 3710 28570 3715
rect 28640 3715 28680 3720
rect 28640 3710 28645 3715
rect 28565 3690 28645 3710
rect 28565 3685 28570 3690
rect 28530 3680 28570 3685
rect 28640 3685 28645 3690
rect 28675 3710 28680 3715
rect 28750 3715 28790 3720
rect 28750 3710 28755 3715
rect 28675 3690 28755 3710
rect 28675 3685 28680 3690
rect 28640 3680 28680 3685
rect 28750 3685 28755 3690
rect 28785 3685 28790 3715
rect 29155 3705 29160 3735
rect 29190 3705 29195 3735
rect 29155 3700 29195 3705
rect 28750 3680 28790 3685
rect 17960 3675 17965 3680
rect 17465 3655 17965 3675
rect 17465 3650 17470 3655
rect 17430 3645 17470 3650
rect 17960 3650 17965 3655
rect 17995 3650 18000 3680
rect 17960 3645 18000 3650
rect 26340 3655 26380 3660
rect 16805 3635 16845 3640
rect 17095 3635 17135 3640
rect 15610 3630 15615 3635
rect 15535 3610 15615 3630
rect 15535 3605 15540 3610
rect 15500 3600 15540 3605
rect 15610 3605 15615 3610
rect 15645 3605 15650 3635
rect 15610 3600 15650 3605
rect 17095 3605 17100 3635
rect 17130 3630 17135 3635
rect 17315 3635 17355 3640
rect 17315 3630 17320 3635
rect 17130 3610 17320 3630
rect 17130 3605 17135 3610
rect 17095 3600 17135 3605
rect 17315 3605 17320 3610
rect 17350 3630 17355 3635
rect 17545 3635 17585 3640
rect 17545 3630 17550 3635
rect 17350 3610 17550 3630
rect 17350 3605 17355 3610
rect 17315 3600 17355 3605
rect 17545 3605 17550 3610
rect 17580 3630 17585 3635
rect 17905 3635 17945 3640
rect 17905 3630 17910 3635
rect 17580 3610 17910 3630
rect 17580 3605 17585 3610
rect 17545 3600 17585 3605
rect 17905 3605 17910 3610
rect 17940 3605 17945 3635
rect 17905 3600 17945 3605
rect 18200 3635 18240 3640
rect 18200 3605 18205 3635
rect 18235 3630 18240 3635
rect 18310 3635 18350 3640
rect 18310 3630 18315 3635
rect 18235 3610 18315 3630
rect 18235 3605 18240 3610
rect 18200 3600 18240 3605
rect 18310 3605 18315 3610
rect 18345 3630 18350 3635
rect 18420 3635 18460 3640
rect 18420 3630 18425 3635
rect 18345 3610 18425 3630
rect 18345 3605 18350 3610
rect 18310 3600 18350 3605
rect 18420 3605 18425 3610
rect 18455 3630 18460 3635
rect 18530 3635 18570 3640
rect 18530 3630 18535 3635
rect 18455 3610 18535 3630
rect 18455 3605 18460 3610
rect 18420 3600 18460 3605
rect 18530 3605 18535 3610
rect 18565 3630 18570 3635
rect 18640 3635 18680 3640
rect 18640 3630 18645 3635
rect 18565 3610 18645 3630
rect 18565 3605 18570 3610
rect 18530 3600 18570 3605
rect 18640 3605 18645 3610
rect 18675 3630 18680 3635
rect 18750 3635 18790 3640
rect 18750 3630 18755 3635
rect 18675 3610 18755 3630
rect 18675 3605 18680 3610
rect 18640 3600 18680 3605
rect 18750 3605 18755 3610
rect 18785 3605 18790 3635
rect 18750 3600 18790 3605
rect 19155 3635 19195 3640
rect 19155 3605 19160 3635
rect 19190 3605 19195 3635
rect 19155 3600 19195 3605
rect 24605 3635 24645 3640
rect 24605 3605 24610 3635
rect 24640 3605 24645 3635
rect 24605 3600 24645 3605
rect 25060 3635 25100 3640
rect 25060 3605 25065 3635
rect 25095 3630 25100 3635
rect 25170 3635 25210 3640
rect 25170 3630 25175 3635
rect 25095 3610 25175 3630
rect 25095 3605 25100 3610
rect 25060 3600 25100 3605
rect 25170 3605 25175 3610
rect 25205 3630 25210 3635
rect 25280 3635 25320 3640
rect 25280 3630 25285 3635
rect 25205 3610 25285 3630
rect 25205 3605 25210 3610
rect 25170 3600 25210 3605
rect 25280 3605 25285 3610
rect 25315 3630 25320 3635
rect 25390 3635 25430 3640
rect 25390 3630 25395 3635
rect 25315 3610 25395 3630
rect 25315 3605 25320 3610
rect 25280 3600 25320 3605
rect 25390 3605 25395 3610
rect 25425 3630 25430 3635
rect 25500 3635 25540 3640
rect 25500 3630 25505 3635
rect 25425 3610 25505 3630
rect 25425 3605 25430 3610
rect 25390 3600 25430 3605
rect 25500 3605 25505 3610
rect 25535 3630 25540 3635
rect 25610 3635 25650 3640
rect 25610 3630 25615 3635
rect 25535 3610 25615 3630
rect 25535 3605 25540 3610
rect 25500 3600 25540 3605
rect 25610 3605 25615 3610
rect 25645 3605 25650 3635
rect 26340 3625 26345 3655
rect 26375 3650 26380 3655
rect 26460 3655 26500 3660
rect 26460 3650 26465 3655
rect 26375 3630 26465 3650
rect 26375 3625 26380 3630
rect 26340 3620 26380 3625
rect 26460 3625 26465 3630
rect 26495 3650 26500 3655
rect 26580 3655 26620 3660
rect 26580 3650 26585 3655
rect 26495 3630 26585 3650
rect 26495 3625 26500 3630
rect 26460 3620 26500 3625
rect 26580 3625 26585 3630
rect 26615 3650 26620 3655
rect 26700 3655 26740 3660
rect 26700 3650 26705 3655
rect 26615 3630 26705 3650
rect 26615 3625 26620 3630
rect 26580 3620 26620 3625
rect 26700 3625 26705 3630
rect 26735 3650 26740 3655
rect 26820 3655 26860 3660
rect 26820 3650 26825 3655
rect 26735 3630 26825 3650
rect 26735 3625 26740 3630
rect 26700 3620 26740 3625
rect 26820 3625 26825 3630
rect 26855 3650 26860 3655
rect 26940 3655 26980 3660
rect 26940 3650 26945 3655
rect 26855 3630 26945 3650
rect 26855 3625 26860 3630
rect 26820 3620 26860 3625
rect 26940 3625 26945 3630
rect 26975 3650 26980 3655
rect 27060 3655 27100 3660
rect 27060 3650 27065 3655
rect 26975 3630 27065 3650
rect 26975 3625 26980 3630
rect 26940 3620 26980 3625
rect 27060 3625 27065 3630
rect 27095 3650 27100 3655
rect 27180 3655 27220 3660
rect 27180 3650 27185 3655
rect 27095 3630 27185 3650
rect 27095 3625 27100 3630
rect 27060 3620 27100 3625
rect 27180 3625 27185 3630
rect 27215 3650 27220 3655
rect 27300 3655 27340 3660
rect 27300 3650 27305 3655
rect 27215 3630 27305 3650
rect 27215 3625 27220 3630
rect 27180 3620 27220 3625
rect 27300 3625 27305 3630
rect 27335 3650 27340 3655
rect 27420 3655 27460 3660
rect 27420 3650 27425 3655
rect 27335 3630 27425 3650
rect 27335 3625 27340 3630
rect 27300 3620 27340 3625
rect 27420 3625 27425 3630
rect 27455 3625 27460 3655
rect 27420 3620 27460 3625
rect 29105 3655 29246 3660
rect 29105 3625 29110 3655
rect 29140 3625 29160 3655
rect 29190 3625 29210 3655
rect 29240 3625 29246 3655
rect 29105 3620 29246 3625
rect 25610 3600 25650 3605
rect 16340 3575 16380 3580
rect 14554 3555 14695 3560
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1261 3525 1301 3530
rect 1261 3520 1266 3525
rect -75 3500 1266 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1261 3495 1266 3500
rect 1296 3495 1301 3525
rect 14554 3525 14560 3555
rect 14590 3525 14610 3555
rect 14640 3525 14660 3555
rect 14690 3525 14695 3555
rect 16340 3545 16345 3575
rect 16375 3570 16380 3575
rect 16460 3575 16500 3580
rect 16460 3570 16465 3575
rect 16375 3550 16465 3570
rect 16375 3545 16380 3550
rect 16340 3540 16380 3545
rect 16460 3545 16465 3550
rect 16495 3570 16500 3575
rect 16580 3575 16620 3580
rect 16580 3570 16585 3575
rect 16495 3550 16585 3570
rect 16495 3545 16500 3550
rect 16460 3540 16500 3545
rect 16580 3545 16585 3550
rect 16615 3570 16620 3575
rect 16700 3575 16740 3580
rect 16700 3570 16705 3575
rect 16615 3550 16705 3570
rect 16615 3545 16620 3550
rect 16580 3540 16620 3545
rect 16700 3545 16705 3550
rect 16735 3570 16740 3575
rect 16820 3575 16860 3580
rect 16820 3570 16825 3575
rect 16735 3550 16825 3570
rect 16735 3545 16740 3550
rect 16700 3540 16740 3545
rect 16820 3545 16825 3550
rect 16855 3570 16860 3575
rect 16940 3575 16980 3580
rect 16940 3570 16945 3575
rect 16855 3550 16945 3570
rect 16855 3545 16860 3550
rect 16820 3540 16860 3545
rect 16940 3545 16945 3550
rect 16975 3570 16980 3575
rect 17060 3575 17100 3580
rect 17060 3570 17065 3575
rect 16975 3550 17065 3570
rect 16975 3545 16980 3550
rect 16940 3540 16980 3545
rect 17060 3545 17065 3550
rect 17095 3570 17100 3575
rect 17180 3575 17220 3580
rect 17180 3570 17185 3575
rect 17095 3550 17185 3570
rect 17095 3545 17100 3550
rect 17060 3540 17100 3545
rect 17180 3545 17185 3550
rect 17215 3570 17220 3575
rect 17300 3575 17340 3580
rect 17300 3570 17305 3575
rect 17215 3550 17305 3570
rect 17215 3545 17220 3550
rect 17180 3540 17220 3545
rect 17300 3545 17305 3550
rect 17335 3570 17340 3575
rect 17420 3575 17460 3580
rect 17420 3570 17425 3575
rect 17335 3550 17425 3570
rect 17335 3545 17340 3550
rect 17300 3540 17340 3545
rect 17420 3545 17425 3550
rect 17455 3545 17460 3575
rect 17420 3540 17460 3545
rect 19105 3555 19246 3560
rect 14554 3520 14695 3525
rect 19105 3525 19110 3555
rect 19140 3525 19160 3555
rect 19190 3525 19210 3555
rect 19240 3525 19246 3555
rect 19105 3520 19246 3525
rect 24554 3555 24695 3560
rect 24554 3525 24560 3555
rect 24590 3525 24610 3555
rect 24640 3525 24660 3555
rect 24690 3525 24695 3555
rect 24554 3520 24695 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5550 3445 5590 3450
rect 5550 3440 5555 3445
rect 5175 3420 5555 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5550 3415 5555 3420
rect 5585 3415 5590 3445
rect 5550 3410 5590 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3335 1245 3340
rect 3135 3340 3175 3345
rect 3135 3335 3140 3340
rect 1240 3315 3140 3335
rect 1240 3310 1245 3315
rect 1205 3305 1245 3310
rect 3135 3310 3140 3315
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5360 3335 5400 3340
rect 5360 3330 5365 3335
rect 3425 3310 5365 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5360 3305 5365 3310
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3280 1200 3285
rect 4885 3285 4925 3290
rect 4885 3280 4890 3285
rect 1195 3260 4890 3280
rect 1195 3255 1200 3260
rect 1160 3250 1200 3255
rect 4885 3255 4890 3260
rect 4920 3280 4925 3285
rect 5410 3285 5450 3290
rect 5410 3280 5415 3285
rect 4920 3260 5415 3280
rect 4920 3255 4925 3260
rect 4885 3250 4925 3255
rect 5410 3255 5415 3260
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 46 3215 2740 3235
rect 46 3205 91 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 26050 3185 26090 3190
rect 26050 3155 26055 3185
rect 26085 3180 26090 3185
rect 26823 3185 26857 3190
rect 26823 3180 26826 3185
rect 26085 3160 26826 3180
rect 26085 3155 26090 3160
rect 26050 3150 26090 3155
rect 26823 3155 26826 3160
rect 26854 3155 26857 3185
rect 26823 3150 26857 3155
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 46 3135 51 3145
rect -75 3115 51 3135
rect -75 3110 -70 3115
rect 46 3110 51 3115
rect 86 3110 91 3145
rect 3135 3140 3175 3145
rect -110 3105 -70 3110
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 3135 3110 3140 3140
rect 3170 3135 3175 3140
rect 4835 3140 4875 3145
rect 4835 3135 4840 3140
rect 3170 3115 4840 3135
rect 3170 3110 3175 3115
rect 3135 3105 3175 3110
rect 4835 3110 4840 3115
rect 4870 3135 4875 3140
rect 5315 3140 5355 3145
rect 5315 3135 5320 3140
rect 4870 3115 5320 3135
rect 4870 3110 4875 3115
rect 4835 3105 4875 3110
rect 5315 3110 5320 3115
rect 5350 3110 5355 3140
rect 26280 3130 26320 3135
rect 5315 3105 5355 3110
rect 16050 3105 16090 3110
rect 1160 3100 1200 3105
rect 1160 3095 1165 3100
rect 46 3075 1165 3095
rect 46 3065 91 3075
rect 1160 3070 1165 3075
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 3985 3080 4025 3085
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 3985 3050 3990 3080
rect 4020 3075 4025 3080
rect 16050 3075 16055 3105
rect 16085 3100 16090 3105
rect 16823 3105 16857 3110
rect 16823 3100 16826 3105
rect 16085 3080 16826 3100
rect 16085 3075 16090 3080
rect 4020 3055 6100 3075
rect 16050 3070 16090 3075
rect 16823 3075 16826 3080
rect 16854 3075 16857 3105
rect 26280 3100 26285 3130
rect 26315 3125 26320 3130
rect 26520 3130 26560 3135
rect 26520 3125 26525 3130
rect 26315 3105 26525 3125
rect 26315 3100 26320 3105
rect 26280 3095 26320 3100
rect 26520 3100 26525 3105
rect 26555 3125 26560 3130
rect 26760 3130 26800 3135
rect 26760 3125 26765 3130
rect 26555 3105 26765 3125
rect 26555 3100 26560 3105
rect 26520 3095 26560 3100
rect 26760 3100 26765 3105
rect 26795 3125 26800 3130
rect 27000 3130 27040 3135
rect 27000 3125 27005 3130
rect 26795 3105 27005 3125
rect 26795 3100 26800 3105
rect 26760 3095 26800 3100
rect 27000 3100 27005 3105
rect 27035 3125 27040 3130
rect 27240 3130 27280 3135
rect 27240 3125 27245 3130
rect 27035 3105 27245 3125
rect 27035 3100 27040 3105
rect 27000 3095 27040 3100
rect 27240 3100 27245 3105
rect 27275 3125 27280 3130
rect 27480 3130 27520 3135
rect 27480 3125 27485 3130
rect 27275 3105 27485 3125
rect 27275 3100 27280 3105
rect 27240 3095 27280 3100
rect 27480 3100 27485 3105
rect 27515 3100 27520 3130
rect 27480 3095 27520 3100
rect 16823 3070 16857 3075
rect 4020 3050 4025 3055
rect 3985 3045 4025 3050
rect 16280 3050 16320 3055
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3030 3485 3035
rect 3805 3035 3845 3040
rect 3805 3030 3810 3035
rect 3480 3010 3810 3030
rect 3480 3005 3485 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 46 2995 51 3005
rect -75 2975 51 2995
rect -75 2970 -70 2975
rect 46 2970 51 2975
rect 86 2970 91 3005
rect 3445 3000 3485 3005
rect 3805 3005 3810 3010
rect 3840 3030 3845 3035
rect 4345 3035 4385 3040
rect 4345 3030 4350 3035
rect 3840 3010 4350 3030
rect 3840 3005 3845 3010
rect 3805 3000 3845 3005
rect 4345 3005 4350 3010
rect 4380 3030 4385 3035
rect 4705 3035 4745 3040
rect 4705 3030 4710 3035
rect 4380 3010 4710 3030
rect 4380 3005 4385 3010
rect 4345 3000 4385 3005
rect 4705 3005 4710 3010
rect 4740 3030 4745 3035
rect 4740 3010 6100 3030
rect 16280 3020 16285 3050
rect 16315 3045 16320 3050
rect 16520 3050 16560 3055
rect 16520 3045 16525 3050
rect 16315 3025 16525 3045
rect 16315 3020 16320 3025
rect 16280 3015 16320 3020
rect 16520 3020 16525 3025
rect 16555 3045 16560 3050
rect 16760 3050 16800 3055
rect 16760 3045 16765 3050
rect 16555 3025 16765 3045
rect 16555 3020 16560 3025
rect 16520 3015 16560 3020
rect 16760 3020 16765 3025
rect 16795 3045 16800 3050
rect 17000 3050 17040 3055
rect 17000 3045 17005 3050
rect 16795 3025 17005 3045
rect 16795 3020 16800 3025
rect 16760 3015 16800 3020
rect 17000 3020 17005 3025
rect 17035 3045 17040 3050
rect 17240 3050 17280 3055
rect 17240 3045 17245 3050
rect 17035 3025 17245 3045
rect 17035 3020 17040 3025
rect 17000 3015 17040 3020
rect 17240 3020 17245 3025
rect 17275 3045 17280 3050
rect 17480 3050 17520 3055
rect 17480 3045 17485 3050
rect 17275 3025 17485 3045
rect 17275 3020 17280 3025
rect 17240 3015 17280 3020
rect 17480 3020 17485 3025
rect 17515 3020 17520 3050
rect 17480 3015 17520 3020
rect 28255 3045 28295 3050
rect 28255 3015 28260 3045
rect 28290 3040 28295 3045
rect 28365 3045 28405 3050
rect 28365 3040 28370 3045
rect 28290 3020 28370 3040
rect 28290 3015 28295 3020
rect 28255 3010 28295 3015
rect 28365 3015 28370 3020
rect 28400 3040 28405 3045
rect 28475 3045 28515 3050
rect 28475 3040 28480 3045
rect 28400 3020 28480 3040
rect 28400 3015 28405 3020
rect 28365 3010 28405 3015
rect 28475 3015 28480 3020
rect 28510 3040 28515 3045
rect 28585 3045 28625 3050
rect 28585 3040 28590 3045
rect 28510 3020 28590 3040
rect 28510 3015 28515 3020
rect 28475 3010 28515 3015
rect 28585 3015 28590 3020
rect 28620 3040 28625 3045
rect 28695 3045 28735 3050
rect 28695 3040 28700 3045
rect 28620 3020 28700 3040
rect 28620 3015 28625 3020
rect 28585 3010 28625 3015
rect 28695 3015 28700 3020
rect 28730 3015 28735 3045
rect 28695 3010 28735 3015
rect 29105 3035 29246 3040
rect 4740 3005 4745 3010
rect 4705 3000 4745 3005
rect 16400 3005 16440 3010
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3080 2980 3120 2985
rect 3080 2975 3085 2980
rect 2555 2955 3085 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3080 2950 3085 2955
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2975 3305 2980
rect 3625 2980 3665 2985
rect 3625 2975 3630 2980
rect 3300 2955 3630 2975
rect 3300 2950 3305 2955
rect 3265 2945 3305 2950
rect 3625 2950 3630 2955
rect 3660 2975 3665 2980
rect 4165 2980 4205 2985
rect 4165 2975 4170 2980
rect 3660 2955 4170 2975
rect 3660 2950 3665 2955
rect 3625 2945 3665 2950
rect 4165 2950 4170 2955
rect 4200 2975 4205 2980
rect 4525 2980 4565 2985
rect 4525 2975 4530 2980
rect 4200 2955 4530 2975
rect 4200 2950 4205 2955
rect 4165 2945 4205 2950
rect 4525 2950 4530 2955
rect 4560 2975 4565 2980
rect 16400 2975 16405 3005
rect 16435 3000 16440 3005
rect 16640 3005 16680 3010
rect 16640 3000 16645 3005
rect 16435 2980 16645 3000
rect 16435 2975 16440 2980
rect 4560 2955 6100 2975
rect 16400 2970 16440 2975
rect 16640 2975 16645 2980
rect 16675 3000 16680 3005
rect 16880 3005 16920 3010
rect 16880 3000 16885 3005
rect 16675 2980 16885 3000
rect 16675 2975 16680 2980
rect 16640 2970 16680 2975
rect 16880 2975 16885 2980
rect 16915 3000 16920 3005
rect 17120 3005 17160 3010
rect 17120 3000 17125 3005
rect 16915 2980 17125 3000
rect 16915 2975 16920 2980
rect 16880 2970 16920 2975
rect 17120 2975 17125 2980
rect 17155 3000 17160 3005
rect 17360 3005 17400 3010
rect 17360 3000 17365 3005
rect 17155 2980 17365 3000
rect 17155 2975 17160 2980
rect 17120 2970 17160 2975
rect 17360 2975 17365 2980
rect 17395 2975 17400 3005
rect 17360 2970 17400 2975
rect 26400 3005 26440 3010
rect 26400 2975 26405 3005
rect 26435 3000 26440 3005
rect 26640 3005 26680 3010
rect 26640 3000 26645 3005
rect 26435 2980 26645 3000
rect 26435 2975 26440 2980
rect 26400 2970 26440 2975
rect 26640 2975 26645 2980
rect 26675 3000 26680 3005
rect 26880 3005 26920 3010
rect 26880 3000 26885 3005
rect 26675 2980 26885 3000
rect 26675 2975 26680 2980
rect 26640 2970 26680 2975
rect 26880 2975 26885 2980
rect 26915 3000 26920 3005
rect 27120 3005 27160 3010
rect 27120 3000 27125 3005
rect 26915 2980 27125 3000
rect 26915 2975 26920 2980
rect 26880 2970 26920 2975
rect 27120 2975 27125 2980
rect 27155 3000 27160 3005
rect 27360 3005 27400 3010
rect 27360 3000 27365 3005
rect 27155 2980 27365 3000
rect 27155 2975 27160 2980
rect 27120 2970 27160 2975
rect 27360 2975 27365 2980
rect 27395 2975 27400 3005
rect 29105 3005 29110 3035
rect 29140 3005 29160 3035
rect 29190 3005 29210 3035
rect 29240 3005 29246 3035
rect 29105 3000 29246 3005
rect 27360 2970 27400 2975
rect 15115 2965 15155 2970
rect 4560 2950 4565 2955
rect 4525 2945 4565 2950
rect 2425 2920 2465 2925
rect 14554 2935 14695 2940
rect -110 2910 -70 2915
rect -110 2880 -105 2910
rect -75 2905 -70 2910
rect 905 2910 1125 2920
rect 905 2905 920 2910
rect -75 2885 920 2905
rect -75 2880 -70 2885
rect -110 2875 -70 2880
rect 905 2880 920 2885
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 14554 2905 14560 2935
rect 14590 2905 14610 2935
rect 14640 2905 14660 2935
rect 14690 2905 14695 2935
rect 15115 2935 15120 2965
rect 15150 2960 15155 2965
rect 15225 2965 15265 2970
rect 15225 2960 15230 2965
rect 15150 2940 15230 2960
rect 15150 2935 15155 2940
rect 15115 2930 15155 2935
rect 15225 2935 15230 2940
rect 15260 2960 15265 2965
rect 15335 2965 15375 2970
rect 15335 2960 15340 2965
rect 15260 2940 15340 2960
rect 15260 2935 15265 2940
rect 15225 2930 15265 2935
rect 15335 2935 15340 2940
rect 15370 2960 15375 2965
rect 15445 2965 15485 2970
rect 15445 2960 15450 2965
rect 15370 2940 15450 2960
rect 15370 2935 15375 2940
rect 15335 2930 15375 2935
rect 15445 2935 15450 2940
rect 15480 2960 15485 2965
rect 15555 2965 15595 2970
rect 15555 2960 15560 2965
rect 15480 2940 15560 2960
rect 15480 2935 15485 2940
rect 15445 2930 15485 2935
rect 15555 2935 15560 2940
rect 15590 2935 15595 2965
rect 18255 2965 18295 2970
rect 15555 2930 15595 2935
rect 16105 2950 16145 2955
rect 16105 2920 16110 2950
rect 16140 2945 16145 2950
rect 16880 2950 16920 2955
rect 16880 2945 16885 2950
rect 16140 2925 16885 2945
rect 16140 2920 16145 2925
rect 16105 2915 16145 2920
rect 16880 2920 16885 2925
rect 16915 2920 16920 2950
rect 18255 2935 18260 2965
rect 18290 2960 18295 2965
rect 18365 2965 18405 2970
rect 18365 2960 18370 2965
rect 18290 2940 18370 2960
rect 18290 2935 18295 2940
rect 18255 2930 18295 2935
rect 18365 2935 18370 2940
rect 18400 2960 18405 2965
rect 18475 2965 18515 2970
rect 18475 2960 18480 2965
rect 18400 2940 18480 2960
rect 18400 2935 18405 2940
rect 18365 2930 18405 2935
rect 18475 2935 18480 2940
rect 18510 2960 18515 2965
rect 18585 2965 18625 2970
rect 18585 2960 18590 2965
rect 18510 2940 18590 2960
rect 18510 2935 18515 2940
rect 18475 2930 18515 2935
rect 18585 2935 18590 2940
rect 18620 2960 18625 2965
rect 18695 2965 18735 2970
rect 18695 2960 18700 2965
rect 18620 2940 18700 2960
rect 18620 2935 18625 2940
rect 18585 2930 18625 2935
rect 18695 2935 18700 2940
rect 18730 2935 18735 2965
rect 25115 2965 25155 2970
rect 18695 2930 18735 2935
rect 19105 2935 19246 2940
rect 16880 2915 16920 2920
rect 905 2870 1125 2880
rect 2330 2900 2375 2905
rect 14554 2900 14695 2905
rect 19105 2905 19110 2935
rect 19140 2905 19160 2935
rect 19190 2905 19210 2935
rect 19240 2905 19246 2935
rect 19105 2900 19246 2905
rect 24554 2935 24695 2940
rect 24554 2905 24560 2935
rect 24590 2905 24610 2935
rect 24640 2905 24660 2935
rect 24690 2905 24695 2935
rect 25115 2935 25120 2965
rect 25150 2960 25155 2965
rect 25225 2965 25265 2970
rect 25225 2960 25230 2965
rect 25150 2940 25230 2960
rect 25150 2935 25155 2940
rect 25115 2930 25155 2935
rect 25225 2935 25230 2940
rect 25260 2960 25265 2965
rect 25335 2965 25375 2970
rect 25335 2960 25340 2965
rect 25260 2940 25340 2960
rect 25260 2935 25265 2940
rect 25225 2930 25265 2935
rect 25335 2935 25340 2940
rect 25370 2960 25375 2965
rect 25445 2965 25485 2970
rect 25445 2960 25450 2965
rect 25370 2940 25450 2960
rect 25370 2935 25375 2940
rect 25335 2930 25375 2935
rect 25445 2935 25450 2940
rect 25480 2960 25485 2965
rect 25555 2965 25595 2970
rect 25555 2960 25560 2965
rect 25480 2940 25560 2960
rect 25480 2935 25485 2940
rect 25445 2930 25485 2935
rect 25555 2935 25560 2940
rect 25590 2935 25595 2965
rect 25555 2930 25595 2935
rect 26105 2950 26145 2955
rect 26105 2920 26110 2950
rect 26140 2945 26145 2950
rect 26880 2950 26920 2955
rect 26880 2945 26885 2950
rect 26140 2925 26885 2945
rect 26140 2920 26145 2925
rect 26105 2915 26145 2920
rect 26880 2920 26885 2925
rect 26915 2920 26920 2950
rect 26880 2915 26920 2920
rect 24554 2900 24695 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 16135 2895 16175 2900
rect 2330 2860 2375 2865
rect 14605 2880 14645 2885
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 51 2850 56 2855
rect -25 2830 56 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 51 2820 56 2830
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2845 769 2855
rect 1205 2850 1245 2855
rect 1205 2845 1210 2850
rect 764 2825 1210 2845
rect 764 2820 769 2825
rect 1205 2820 1210 2825
rect 1240 2820 1245 2850
rect 14605 2850 14610 2880
rect 14640 2875 14645 2880
rect 15500 2880 15540 2885
rect 15500 2875 15505 2880
rect 14640 2855 15505 2875
rect 14640 2850 14645 2855
rect 14605 2845 14645 2850
rect 15500 2850 15505 2855
rect 15535 2875 15540 2880
rect 15780 2880 15820 2885
rect 15780 2875 15785 2880
rect 15535 2855 15785 2875
rect 15535 2850 15540 2855
rect 15500 2845 15540 2850
rect 15780 2850 15785 2855
rect 15815 2850 15820 2880
rect 16135 2865 16140 2895
rect 16170 2890 16175 2895
rect 16255 2895 16295 2900
rect 16255 2890 16260 2895
rect 16170 2870 16260 2890
rect 16170 2865 16175 2870
rect 16135 2860 16175 2865
rect 16255 2865 16260 2870
rect 16290 2890 16295 2895
rect 16375 2895 16415 2900
rect 16375 2890 16380 2895
rect 16290 2870 16380 2890
rect 16290 2865 16295 2870
rect 16255 2860 16295 2865
rect 16375 2865 16380 2870
rect 16410 2890 16415 2895
rect 16495 2895 16535 2900
rect 16495 2890 16500 2895
rect 16410 2870 16500 2890
rect 16410 2865 16415 2870
rect 16375 2860 16415 2865
rect 16495 2865 16500 2870
rect 16530 2890 16535 2895
rect 16615 2895 16655 2900
rect 16615 2890 16620 2895
rect 16530 2870 16620 2890
rect 16530 2865 16535 2870
rect 16495 2860 16535 2865
rect 16615 2865 16620 2870
rect 16650 2865 16655 2895
rect 16615 2860 16655 2865
rect 17145 2895 17185 2900
rect 17145 2865 17150 2895
rect 17180 2890 17185 2895
rect 17265 2895 17305 2900
rect 17265 2890 17270 2895
rect 17180 2870 17270 2890
rect 17180 2865 17185 2870
rect 17145 2860 17185 2865
rect 17265 2865 17270 2870
rect 17300 2890 17305 2895
rect 17385 2895 17425 2900
rect 17385 2890 17390 2895
rect 17300 2870 17390 2890
rect 17300 2865 17305 2870
rect 17265 2860 17305 2865
rect 17385 2865 17390 2870
rect 17420 2890 17425 2895
rect 17505 2895 17545 2900
rect 17505 2890 17510 2895
rect 17420 2870 17510 2890
rect 17420 2865 17425 2870
rect 17385 2860 17425 2865
rect 17505 2865 17510 2870
rect 17540 2890 17545 2895
rect 17625 2895 17665 2900
rect 17625 2890 17630 2895
rect 17540 2870 17630 2890
rect 17540 2865 17545 2870
rect 17505 2860 17545 2865
rect 17625 2865 17630 2870
rect 17660 2865 17665 2895
rect 26135 2895 26175 2900
rect 17625 2860 17665 2865
rect 18015 2880 18055 2885
rect 15780 2845 15820 2850
rect 18015 2850 18020 2880
rect 18050 2875 18055 2880
rect 18310 2880 18350 2885
rect 18310 2875 18315 2880
rect 18050 2855 18315 2875
rect 18050 2850 18055 2855
rect 18015 2845 18055 2850
rect 18310 2850 18315 2855
rect 18345 2875 18350 2880
rect 19155 2880 19195 2885
rect 19155 2875 19160 2880
rect 18345 2855 19160 2875
rect 18345 2850 18350 2855
rect 18310 2845 18350 2850
rect 19155 2850 19160 2855
rect 19190 2850 19195 2880
rect 19155 2845 19195 2850
rect 24605 2880 24645 2885
rect 24605 2850 24610 2880
rect 24640 2875 24645 2880
rect 25500 2880 25540 2885
rect 25500 2875 25505 2880
rect 24640 2855 25505 2875
rect 24640 2850 24645 2855
rect 24605 2845 24645 2850
rect 25500 2850 25505 2855
rect 25535 2875 25540 2880
rect 25780 2880 25820 2885
rect 25780 2875 25785 2880
rect 25535 2855 25785 2875
rect 25535 2850 25540 2855
rect 25500 2845 25540 2850
rect 25780 2850 25785 2855
rect 25815 2850 25820 2880
rect 26135 2865 26140 2895
rect 26170 2890 26175 2895
rect 26255 2895 26295 2900
rect 26255 2890 26260 2895
rect 26170 2870 26260 2890
rect 26170 2865 26175 2870
rect 26135 2860 26175 2865
rect 26255 2865 26260 2870
rect 26290 2890 26295 2895
rect 26375 2895 26415 2900
rect 26375 2890 26380 2895
rect 26290 2870 26380 2890
rect 26290 2865 26295 2870
rect 26255 2860 26295 2865
rect 26375 2865 26380 2870
rect 26410 2890 26415 2895
rect 26495 2895 26535 2900
rect 26495 2890 26500 2895
rect 26410 2870 26500 2890
rect 26410 2865 26415 2870
rect 26375 2860 26415 2865
rect 26495 2865 26500 2870
rect 26530 2890 26535 2895
rect 26615 2895 26655 2900
rect 26615 2890 26620 2895
rect 26530 2870 26620 2890
rect 26530 2865 26535 2870
rect 26495 2860 26535 2865
rect 26615 2865 26620 2870
rect 26650 2865 26655 2895
rect 26615 2860 26655 2865
rect 27155 2895 27195 2900
rect 27155 2865 27160 2895
rect 27190 2890 27195 2895
rect 27275 2895 27315 2900
rect 27275 2890 27280 2895
rect 27190 2870 27280 2890
rect 27190 2865 27195 2870
rect 27155 2860 27195 2865
rect 27275 2865 27280 2870
rect 27310 2890 27315 2895
rect 27395 2895 27435 2900
rect 27395 2890 27400 2895
rect 27310 2870 27400 2890
rect 27310 2865 27315 2870
rect 27275 2860 27315 2865
rect 27395 2865 27400 2870
rect 27430 2890 27435 2895
rect 27515 2895 27555 2900
rect 27515 2890 27520 2895
rect 27430 2870 27520 2890
rect 27430 2865 27435 2870
rect 27395 2860 27435 2865
rect 27515 2865 27520 2870
rect 27550 2890 27555 2895
rect 27635 2895 27675 2900
rect 27635 2890 27640 2895
rect 27550 2870 27640 2890
rect 27550 2865 27555 2870
rect 27515 2860 27555 2865
rect 27635 2865 27640 2870
rect 27670 2865 27675 2895
rect 27635 2860 27675 2865
rect 28015 2880 28055 2885
rect 25780 2845 25820 2850
rect 28015 2850 28020 2880
rect 28050 2875 28055 2880
rect 28310 2880 28350 2885
rect 28310 2875 28315 2880
rect 28050 2855 28315 2875
rect 28050 2850 28055 2855
rect 28015 2845 28055 2850
rect 28310 2850 28315 2855
rect 28345 2875 28350 2880
rect 29155 2880 29195 2885
rect 29155 2875 29160 2880
rect 28345 2855 29160 2875
rect 28345 2850 28350 2855
rect 28310 2845 28350 2850
rect 29155 2850 29160 2855
rect 29190 2850 29195 2880
rect 29155 2845 29195 2850
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 28585 2835 28625 2840
rect 14515 2825 14555 2830
rect 2330 2800 2370 2805
rect 2995 2810 3035 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 51 2785 56 2795
rect 20 2765 56 2785
rect -15 2760 25 2765
rect 51 2760 56 2765
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2785 769 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 764 2765 2625 2785
rect 764 2760 769 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2995 2780 3000 2810
rect 3030 2805 3035 2810
rect 3175 2810 3215 2815
rect 3175 2805 3180 2810
rect 3030 2785 3180 2805
rect 3030 2780 3035 2785
rect 2995 2775 3035 2780
rect 3175 2780 3180 2785
rect 3210 2805 3215 2810
rect 3355 2810 3395 2815
rect 3355 2805 3360 2810
rect 3210 2785 3360 2805
rect 3210 2780 3215 2785
rect 3175 2775 3215 2780
rect 3355 2780 3360 2785
rect 3390 2805 3395 2810
rect 3535 2810 3575 2815
rect 3535 2805 3540 2810
rect 3390 2785 3540 2805
rect 3390 2780 3395 2785
rect 3355 2775 3395 2780
rect 3535 2780 3540 2785
rect 3570 2805 3575 2810
rect 3715 2810 3755 2815
rect 3715 2805 3720 2810
rect 3570 2785 3720 2805
rect 3570 2780 3575 2785
rect 3535 2775 3575 2780
rect 3715 2780 3720 2785
rect 3750 2805 3755 2810
rect 3895 2810 3935 2815
rect 3895 2805 3900 2810
rect 3750 2785 3900 2805
rect 3750 2780 3755 2785
rect 3715 2775 3755 2780
rect 3895 2780 3900 2785
rect 3930 2805 3935 2810
rect 4075 2810 4115 2815
rect 4075 2805 4080 2810
rect 3930 2785 4080 2805
rect 3930 2780 3935 2785
rect 3895 2775 3935 2780
rect 4075 2780 4080 2785
rect 4110 2805 4115 2810
rect 4255 2810 4295 2815
rect 4255 2805 4260 2810
rect 4110 2785 4260 2805
rect 4110 2780 4115 2785
rect 4075 2775 4115 2780
rect 4255 2780 4260 2785
rect 4290 2805 4295 2810
rect 4435 2810 4475 2815
rect 4435 2805 4440 2810
rect 4290 2785 4440 2805
rect 4290 2780 4295 2785
rect 4255 2775 4295 2780
rect 4435 2780 4440 2785
rect 4470 2805 4475 2810
rect 4615 2810 4655 2815
rect 4615 2805 4620 2810
rect 4470 2785 4620 2805
rect 4470 2780 4475 2785
rect 4435 2775 4475 2780
rect 4615 2780 4620 2785
rect 4650 2805 4655 2810
rect 4795 2810 4835 2815
rect 4795 2805 4800 2810
rect 4650 2785 4800 2805
rect 4650 2780 4655 2785
rect 4615 2775 4655 2780
rect 4795 2780 4800 2785
rect 4830 2805 4835 2810
rect 4975 2810 5015 2815
rect 4975 2805 4980 2810
rect 4830 2785 4980 2805
rect 4830 2780 4835 2785
rect 4795 2775 4835 2780
rect 4975 2780 4980 2785
rect 5010 2805 5015 2810
rect 5550 2810 5590 2815
rect 5550 2805 5555 2810
rect 5010 2785 5555 2805
rect 5010 2780 5015 2785
rect 4975 2775 5015 2780
rect 5550 2780 5555 2785
rect 5585 2780 5590 2810
rect 14515 2795 14520 2825
rect 14550 2820 14555 2825
rect 15225 2825 15265 2830
rect 15225 2820 15230 2825
rect 14550 2800 15230 2820
rect 14550 2795 14555 2800
rect 14515 2790 14555 2795
rect 15225 2795 15230 2800
rect 15260 2795 15265 2825
rect 15225 2790 15265 2795
rect 18585 2825 18625 2830
rect 18585 2795 18590 2825
rect 18620 2820 18625 2825
rect 19245 2825 19285 2830
rect 19245 2820 19250 2825
rect 18620 2800 19250 2820
rect 18620 2795 18625 2800
rect 18585 2790 18625 2795
rect 19245 2795 19250 2800
rect 19280 2795 19285 2825
rect 19245 2790 19285 2795
rect 24515 2825 24555 2830
rect 24515 2795 24520 2825
rect 24550 2820 24555 2825
rect 25225 2825 25265 2830
rect 25225 2820 25230 2825
rect 24550 2800 25230 2820
rect 24550 2795 24555 2800
rect 24515 2790 24555 2795
rect 25225 2795 25230 2800
rect 25260 2795 25265 2825
rect 28585 2805 28590 2835
rect 28620 2830 28625 2835
rect 29395 2835 29435 2840
rect 29395 2830 29400 2835
rect 28620 2810 29400 2830
rect 28620 2805 28625 2810
rect 28585 2800 28625 2805
rect 29395 2805 29400 2810
rect 29430 2805 29435 2835
rect 29395 2800 29435 2805
rect 25225 2790 25265 2795
rect 5550 2775 5590 2780
rect 2620 2755 2660 2760
rect 28200 2755 28240 2760
rect 3175 2750 3215 2755
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2740 1301 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1296 2720 2155 2740
rect 1296 2715 1301 2720
rect 1261 2710 1301 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 3175 2720 3180 2750
rect 3210 2745 3215 2750
rect 3355 2750 3395 2755
rect 3355 2745 3360 2750
rect 3210 2725 3360 2745
rect 3210 2720 3215 2725
rect 3175 2715 3215 2720
rect 3355 2720 3360 2725
rect 3390 2745 3395 2750
rect 3535 2750 3575 2755
rect 3535 2745 3540 2750
rect 3390 2725 3540 2745
rect 3390 2720 3395 2725
rect 3355 2715 3395 2720
rect 3535 2720 3540 2725
rect 3570 2745 3575 2750
rect 3715 2750 3755 2755
rect 3715 2745 3720 2750
rect 3570 2725 3720 2745
rect 3570 2720 3575 2725
rect 3535 2715 3575 2720
rect 3715 2720 3720 2725
rect 3750 2745 3755 2750
rect 3895 2750 3935 2755
rect 3895 2745 3900 2750
rect 3750 2725 3900 2745
rect 3750 2720 3755 2725
rect 3715 2715 3755 2720
rect 3895 2720 3900 2725
rect 3930 2745 3935 2750
rect 4075 2750 4115 2755
rect 4075 2745 4080 2750
rect 3930 2725 4080 2745
rect 3930 2720 3935 2725
rect 3895 2715 3935 2720
rect 4075 2720 4080 2725
rect 4110 2745 4115 2750
rect 4255 2750 4295 2755
rect 4255 2745 4260 2750
rect 4110 2725 4260 2745
rect 4110 2720 4115 2725
rect 4075 2715 4115 2720
rect 4255 2720 4260 2725
rect 4290 2745 4295 2750
rect 4435 2750 4475 2755
rect 4435 2745 4440 2750
rect 4290 2725 4440 2745
rect 4290 2720 4295 2725
rect 4255 2715 4295 2720
rect 4435 2720 4440 2725
rect 4470 2745 4475 2750
rect 4615 2750 4655 2755
rect 4615 2745 4620 2750
rect 4470 2725 4620 2745
rect 4470 2720 4475 2725
rect 4435 2715 4475 2720
rect 4615 2720 4620 2725
rect 4650 2745 4655 2750
rect 4795 2750 4835 2755
rect 4795 2745 4800 2750
rect 4650 2725 4800 2745
rect 4650 2720 4655 2725
rect 4615 2715 4655 2720
rect 4795 2720 4800 2725
rect 4830 2720 4835 2750
rect 28200 2725 28205 2755
rect 28235 2750 28240 2755
rect 28310 2755 28350 2760
rect 28310 2750 28315 2755
rect 28235 2730 28315 2750
rect 28235 2725 28240 2730
rect 28200 2720 28240 2725
rect 28310 2725 28315 2730
rect 28345 2750 28350 2755
rect 28420 2755 28460 2760
rect 28420 2750 28425 2755
rect 28345 2730 28425 2750
rect 28345 2725 28350 2730
rect 28310 2720 28350 2725
rect 28420 2725 28425 2730
rect 28455 2750 28460 2755
rect 28530 2755 28570 2760
rect 28530 2750 28535 2755
rect 28455 2730 28535 2750
rect 28455 2725 28460 2730
rect 28420 2720 28460 2725
rect 28530 2725 28535 2730
rect 28565 2750 28570 2755
rect 28640 2755 28680 2760
rect 28640 2750 28645 2755
rect 28565 2730 28645 2750
rect 28565 2725 28570 2730
rect 28530 2720 28570 2725
rect 28640 2725 28645 2730
rect 28675 2750 28680 2755
rect 28750 2755 28790 2760
rect 28750 2750 28755 2755
rect 28675 2730 28755 2750
rect 28675 2725 28680 2730
rect 28640 2720 28680 2725
rect 28750 2725 28755 2730
rect 28785 2725 28790 2755
rect 28750 2720 28790 2725
rect 4795 2715 4835 2720
rect 2150 2710 2190 2715
rect 15060 2705 15100 2710
rect 15060 2675 15065 2705
rect 15095 2700 15100 2705
rect 15170 2705 15210 2710
rect 15170 2700 15175 2705
rect 15095 2680 15175 2700
rect 15095 2675 15100 2680
rect 15060 2670 15100 2675
rect 15170 2675 15175 2680
rect 15205 2700 15210 2705
rect 15280 2705 15320 2710
rect 15280 2700 15285 2705
rect 15205 2680 15285 2700
rect 15205 2675 15210 2680
rect 15170 2670 15210 2675
rect 15280 2675 15285 2680
rect 15315 2700 15320 2705
rect 15390 2705 15430 2710
rect 15390 2700 15395 2705
rect 15315 2680 15395 2700
rect 15315 2675 15320 2680
rect 15280 2670 15320 2675
rect 15390 2675 15395 2680
rect 15425 2700 15430 2705
rect 15500 2705 15540 2710
rect 15500 2700 15505 2705
rect 15425 2680 15505 2700
rect 15425 2675 15430 2680
rect 15390 2670 15430 2675
rect 15500 2675 15505 2680
rect 15535 2700 15540 2705
rect 15610 2705 15650 2710
rect 15610 2700 15615 2705
rect 15535 2680 15615 2700
rect 15535 2675 15540 2680
rect 15500 2670 15540 2675
rect 15610 2675 15615 2680
rect 15645 2675 15650 2705
rect 15610 2670 15650 2675
rect 18200 2705 18240 2710
rect 18200 2675 18205 2705
rect 18235 2700 18240 2705
rect 18310 2705 18350 2710
rect 18310 2700 18315 2705
rect 18235 2680 18315 2700
rect 18235 2675 18240 2680
rect 18200 2670 18240 2675
rect 18310 2675 18315 2680
rect 18345 2700 18350 2705
rect 18420 2705 18460 2710
rect 18420 2700 18425 2705
rect 18345 2680 18425 2700
rect 18345 2675 18350 2680
rect 18310 2670 18350 2675
rect 18420 2675 18425 2680
rect 18455 2700 18460 2705
rect 18530 2705 18570 2710
rect 18530 2700 18535 2705
rect 18455 2680 18535 2700
rect 18455 2675 18460 2680
rect 18420 2670 18460 2675
rect 18530 2675 18535 2680
rect 18565 2700 18570 2705
rect 18640 2705 18680 2710
rect 18640 2700 18645 2705
rect 18565 2680 18645 2700
rect 18565 2675 18570 2680
rect 18530 2670 18570 2675
rect 18640 2675 18645 2680
rect 18675 2700 18680 2705
rect 18750 2705 18790 2710
rect 18750 2700 18755 2705
rect 18675 2680 18755 2700
rect 18675 2675 18680 2680
rect 18640 2670 18680 2675
rect 18750 2675 18755 2680
rect 18785 2675 18790 2705
rect 18750 2670 18790 2675
rect 25060 2705 25100 2710
rect 25060 2675 25065 2705
rect 25095 2700 25100 2705
rect 25170 2705 25210 2710
rect 25170 2700 25175 2705
rect 25095 2680 25175 2700
rect 25095 2675 25100 2680
rect 25060 2670 25100 2675
rect 25170 2675 25175 2680
rect 25205 2700 25210 2705
rect 25280 2705 25320 2710
rect 25280 2700 25285 2705
rect 25205 2680 25285 2700
rect 25205 2675 25210 2680
rect 25170 2670 25210 2675
rect 25280 2675 25285 2680
rect 25315 2700 25320 2705
rect 25390 2705 25430 2710
rect 25390 2700 25395 2705
rect 25315 2680 25395 2700
rect 25315 2675 25320 2680
rect 25280 2670 25320 2675
rect 25390 2675 25395 2680
rect 25425 2700 25430 2705
rect 25500 2705 25540 2710
rect 25500 2700 25505 2705
rect 25425 2680 25505 2700
rect 25425 2675 25430 2680
rect 25390 2670 25430 2675
rect 25500 2675 25505 2680
rect 25535 2700 25540 2705
rect 25610 2705 25650 2710
rect 25610 2700 25615 2705
rect 25535 2680 25615 2700
rect 25535 2675 25540 2680
rect 25500 2670 25540 2675
rect 25610 2675 25615 2680
rect 25645 2675 25650 2705
rect 25610 2670 25650 2675
rect 28255 2485 28295 2490
rect 16075 2475 16115 2480
rect 16075 2445 16080 2475
rect 16110 2470 16115 2475
rect 16195 2475 16235 2480
rect 16195 2470 16200 2475
rect 16110 2450 16200 2470
rect 16110 2445 16115 2450
rect 16075 2440 16115 2445
rect 16195 2445 16200 2450
rect 16230 2470 16235 2475
rect 16315 2475 16355 2480
rect 16315 2470 16320 2475
rect 16230 2450 16320 2470
rect 16230 2445 16235 2450
rect 16195 2440 16235 2445
rect 16315 2445 16320 2450
rect 16350 2470 16355 2475
rect 16435 2475 16475 2480
rect 16435 2470 16440 2475
rect 16350 2450 16440 2470
rect 16350 2445 16355 2450
rect 16315 2440 16355 2445
rect 16435 2445 16440 2450
rect 16470 2470 16475 2475
rect 16555 2475 16595 2480
rect 16555 2470 16560 2475
rect 16470 2450 16560 2470
rect 16470 2445 16475 2450
rect 16435 2440 16475 2445
rect 16555 2445 16560 2450
rect 16590 2470 16595 2475
rect 16675 2475 16715 2480
rect 16675 2470 16680 2475
rect 16590 2450 16680 2470
rect 16590 2445 16595 2450
rect 16555 2440 16595 2445
rect 16675 2445 16680 2450
rect 16710 2445 16715 2475
rect 16675 2440 16715 2445
rect 17085 2475 17125 2480
rect 17085 2445 17090 2475
rect 17120 2470 17125 2475
rect 17205 2475 17245 2480
rect 17205 2470 17210 2475
rect 17120 2450 17210 2470
rect 17120 2445 17125 2450
rect 17085 2440 17125 2445
rect 17205 2445 17210 2450
rect 17240 2470 17245 2475
rect 17325 2475 17365 2480
rect 17325 2470 17330 2475
rect 17240 2450 17330 2470
rect 17240 2445 17245 2450
rect 17205 2440 17245 2445
rect 17325 2445 17330 2450
rect 17360 2470 17365 2475
rect 17445 2475 17485 2480
rect 17445 2470 17450 2475
rect 17360 2450 17450 2470
rect 17360 2445 17365 2450
rect 17325 2440 17365 2445
rect 17445 2445 17450 2450
rect 17480 2470 17485 2475
rect 17565 2475 17605 2480
rect 17565 2470 17570 2475
rect 17480 2450 17570 2470
rect 17480 2445 17485 2450
rect 17445 2440 17485 2445
rect 17565 2445 17570 2450
rect 17600 2470 17605 2475
rect 17685 2475 17725 2480
rect 17685 2470 17690 2475
rect 17600 2450 17690 2470
rect 17600 2445 17605 2450
rect 17565 2440 17605 2445
rect 17685 2445 17690 2450
rect 17720 2445 17725 2475
rect 17685 2440 17725 2445
rect 26075 2475 26115 2480
rect 26075 2445 26080 2475
rect 26110 2470 26115 2475
rect 26195 2475 26235 2480
rect 26195 2470 26200 2475
rect 26110 2450 26200 2470
rect 26110 2445 26115 2450
rect 26075 2440 26115 2445
rect 26195 2445 26200 2450
rect 26230 2470 26235 2475
rect 26315 2475 26355 2480
rect 26315 2470 26320 2475
rect 26230 2450 26320 2470
rect 26230 2445 26235 2450
rect 26195 2440 26235 2445
rect 26315 2445 26320 2450
rect 26350 2470 26355 2475
rect 26435 2475 26475 2480
rect 26435 2470 26440 2475
rect 26350 2450 26440 2470
rect 26350 2445 26355 2450
rect 26315 2440 26355 2445
rect 26435 2445 26440 2450
rect 26470 2470 26475 2475
rect 26555 2475 26595 2480
rect 26555 2470 26560 2475
rect 26470 2450 26560 2470
rect 26470 2445 26475 2450
rect 26435 2440 26475 2445
rect 26555 2445 26560 2450
rect 26590 2470 26595 2475
rect 26675 2475 26715 2480
rect 26675 2470 26680 2475
rect 26590 2450 26680 2470
rect 26590 2445 26595 2450
rect 26555 2440 26595 2445
rect 26675 2445 26680 2450
rect 26710 2445 26715 2475
rect 26675 2440 26715 2445
rect 27095 2475 27135 2480
rect 27095 2445 27100 2475
rect 27130 2470 27135 2475
rect 27215 2475 27255 2480
rect 27215 2470 27220 2475
rect 27130 2450 27220 2470
rect 27130 2445 27135 2450
rect 27095 2440 27135 2445
rect 27215 2445 27220 2450
rect 27250 2470 27255 2475
rect 27335 2475 27375 2480
rect 27335 2470 27340 2475
rect 27250 2450 27340 2470
rect 27250 2445 27255 2450
rect 27215 2440 27255 2445
rect 27335 2445 27340 2450
rect 27370 2470 27375 2475
rect 27455 2475 27495 2480
rect 27455 2470 27460 2475
rect 27370 2450 27460 2470
rect 27370 2445 27375 2450
rect 27335 2440 27375 2445
rect 27455 2445 27460 2450
rect 27490 2470 27495 2475
rect 27575 2475 27615 2480
rect 27575 2470 27580 2475
rect 27490 2450 27580 2470
rect 27490 2445 27495 2450
rect 27455 2440 27495 2445
rect 27575 2445 27580 2450
rect 27610 2470 27615 2475
rect 27695 2475 27735 2480
rect 27695 2470 27700 2475
rect 27610 2450 27700 2470
rect 27610 2445 27615 2450
rect 27575 2440 27615 2445
rect 27695 2445 27700 2450
rect 27730 2445 27735 2475
rect 28255 2455 28260 2485
rect 28290 2480 28295 2485
rect 28365 2485 28405 2490
rect 28365 2480 28370 2485
rect 28290 2460 28370 2480
rect 28290 2455 28295 2460
rect 28255 2450 28295 2455
rect 28365 2455 28370 2460
rect 28400 2480 28405 2485
rect 28475 2485 28515 2490
rect 28475 2480 28480 2485
rect 28400 2460 28480 2480
rect 28400 2455 28405 2460
rect 28365 2450 28405 2455
rect 28475 2455 28480 2460
rect 28510 2480 28515 2485
rect 28585 2485 28625 2490
rect 28585 2480 28590 2485
rect 28510 2460 28590 2480
rect 28510 2455 28515 2460
rect 28475 2450 28515 2455
rect 28585 2455 28590 2460
rect 28620 2480 28625 2485
rect 28695 2485 28735 2490
rect 28695 2480 28700 2485
rect 28620 2460 28700 2480
rect 28620 2455 28625 2460
rect 28585 2450 28625 2455
rect 28695 2455 28700 2460
rect 28730 2480 28735 2485
rect 28940 2485 28980 2490
rect 28940 2480 28945 2485
rect 28730 2460 28945 2480
rect 28730 2455 28735 2460
rect 28695 2450 28735 2455
rect 28940 2455 28945 2460
rect 28975 2455 28980 2485
rect 28940 2450 28980 2455
rect 27695 2440 27735 2445
rect 14870 2435 14910 2440
rect 14870 2405 14875 2435
rect 14905 2430 14910 2435
rect 15115 2435 15155 2440
rect 15115 2430 15120 2435
rect 14905 2410 15120 2430
rect 14905 2405 14910 2410
rect 14870 2400 14910 2405
rect 15115 2405 15120 2410
rect 15150 2430 15155 2435
rect 15225 2435 15265 2440
rect 15225 2430 15230 2435
rect 15150 2410 15230 2430
rect 15150 2405 15155 2410
rect 15115 2400 15155 2405
rect 15225 2405 15230 2410
rect 15260 2430 15265 2435
rect 15335 2435 15375 2440
rect 15335 2430 15340 2435
rect 15260 2410 15340 2430
rect 15260 2405 15265 2410
rect 15225 2400 15265 2405
rect 15335 2405 15340 2410
rect 15370 2430 15375 2435
rect 15445 2435 15485 2440
rect 15445 2430 15450 2435
rect 15370 2410 15450 2430
rect 15370 2405 15375 2410
rect 15335 2400 15375 2405
rect 15445 2405 15450 2410
rect 15480 2430 15485 2435
rect 15555 2435 15595 2440
rect 15555 2430 15560 2435
rect 15480 2410 15560 2430
rect 15480 2405 15485 2410
rect 15445 2400 15485 2405
rect 15555 2405 15560 2410
rect 15590 2405 15595 2435
rect 18255 2435 18295 2440
rect 15555 2400 15595 2405
rect 16375 2420 16415 2425
rect 16375 2390 16380 2420
rect 16410 2415 16415 2420
rect 16880 2420 16920 2425
rect 16880 2415 16885 2420
rect 16410 2395 16885 2415
rect 16410 2390 16415 2395
rect 16375 2385 16415 2390
rect 16880 2390 16885 2395
rect 16915 2415 16920 2420
rect 17385 2420 17425 2425
rect 17385 2415 17390 2420
rect 16915 2395 17390 2415
rect 16915 2390 16920 2395
rect 16880 2385 16920 2390
rect 17385 2390 17390 2395
rect 17420 2390 17425 2420
rect 18255 2405 18260 2435
rect 18290 2430 18295 2435
rect 18365 2435 18405 2440
rect 18365 2430 18370 2435
rect 18290 2410 18370 2430
rect 18290 2405 18295 2410
rect 18255 2400 18295 2405
rect 18365 2405 18370 2410
rect 18400 2430 18405 2435
rect 18475 2435 18515 2440
rect 18475 2430 18480 2435
rect 18400 2410 18480 2430
rect 18400 2405 18405 2410
rect 18365 2400 18405 2405
rect 18475 2405 18480 2410
rect 18510 2430 18515 2435
rect 18585 2435 18625 2440
rect 18585 2430 18590 2435
rect 18510 2410 18590 2430
rect 18510 2405 18515 2410
rect 18475 2400 18515 2405
rect 18585 2405 18590 2410
rect 18620 2430 18625 2435
rect 18695 2435 18735 2440
rect 18695 2430 18700 2435
rect 18620 2410 18700 2430
rect 18620 2405 18625 2410
rect 18585 2400 18625 2405
rect 18695 2405 18700 2410
rect 18730 2430 18735 2435
rect 18940 2435 18980 2440
rect 18940 2430 18945 2435
rect 18730 2410 18945 2430
rect 18730 2405 18735 2410
rect 18695 2400 18735 2405
rect 18940 2405 18945 2410
rect 18975 2405 18980 2435
rect 18940 2400 18980 2405
rect 24870 2435 24910 2440
rect 24870 2405 24875 2435
rect 24905 2430 24910 2435
rect 25115 2435 25155 2440
rect 25115 2430 25120 2435
rect 24905 2410 25120 2430
rect 24905 2405 24910 2410
rect 24870 2400 24910 2405
rect 25115 2405 25120 2410
rect 25150 2430 25155 2435
rect 25225 2435 25265 2440
rect 25225 2430 25230 2435
rect 25150 2410 25230 2430
rect 25150 2405 25155 2410
rect 25115 2400 25155 2405
rect 25225 2405 25230 2410
rect 25260 2430 25265 2435
rect 25335 2435 25375 2440
rect 25335 2430 25340 2435
rect 25260 2410 25340 2430
rect 25260 2405 25265 2410
rect 25225 2400 25265 2405
rect 25335 2405 25340 2410
rect 25370 2430 25375 2435
rect 25445 2435 25485 2440
rect 25445 2430 25450 2435
rect 25370 2410 25450 2430
rect 25370 2405 25375 2410
rect 25335 2400 25375 2405
rect 25445 2405 25450 2410
rect 25480 2430 25485 2435
rect 25555 2435 25595 2440
rect 25555 2430 25560 2435
rect 25480 2410 25560 2430
rect 25480 2405 25485 2410
rect 25445 2400 25485 2405
rect 25555 2405 25560 2410
rect 25590 2405 25595 2435
rect 25555 2400 25595 2405
rect 26375 2420 26415 2425
rect 17385 2385 17425 2390
rect 26375 2390 26380 2420
rect 26410 2415 26415 2420
rect 26880 2420 26920 2425
rect 26880 2415 26885 2420
rect 26410 2395 26885 2415
rect 26410 2390 26415 2395
rect 26375 2385 26415 2390
rect 26880 2390 26885 2395
rect 26915 2415 26920 2420
rect 27395 2420 27435 2425
rect 27395 2415 27400 2420
rect 26915 2395 27400 2415
rect 26915 2390 26920 2395
rect 26880 2385 26920 2390
rect 27395 2390 27400 2395
rect 27430 2390 27435 2420
rect 27395 2385 27435 2390
rect 3805 2380 3845 2385
rect 3355 2375 3395 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3805 2350 3810 2380
rect 3840 2375 3845 2380
rect 4165 2380 4205 2385
rect 4165 2375 4170 2380
rect 3840 2355 4170 2375
rect 3840 2350 3845 2355
rect 3805 2345 3845 2350
rect 4165 2350 4170 2355
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 15585 2375 15625 2380
rect 15585 2345 15590 2375
rect 15620 2370 15625 2375
rect 15780 2375 15820 2380
rect 15780 2370 15785 2375
rect 15620 2350 15785 2370
rect 15620 2345 15625 2350
rect 3355 2340 3395 2345
rect 15585 2340 15625 2345
rect 15780 2345 15785 2350
rect 15815 2370 15820 2375
rect 16320 2375 16360 2380
rect 16320 2370 16325 2375
rect 15815 2350 16325 2370
rect 15815 2345 15820 2350
rect 15780 2340 15820 2345
rect 16320 2345 16325 2350
rect 16355 2345 16360 2375
rect 16320 2340 16360 2345
rect 17320 2375 17360 2380
rect 17320 2345 17325 2375
rect 17355 2370 17360 2375
rect 18015 2375 18055 2380
rect 18015 2370 18020 2375
rect 17355 2350 18020 2370
rect 17355 2345 17360 2350
rect 17320 2340 17360 2345
rect 18015 2345 18020 2350
rect 18050 2370 18055 2375
rect 18225 2375 18265 2380
rect 18225 2370 18230 2375
rect 18050 2350 18230 2370
rect 18050 2345 18055 2350
rect 18015 2340 18055 2345
rect 18225 2345 18230 2350
rect 18260 2345 18265 2375
rect 18225 2340 18265 2345
rect 25585 2375 25625 2380
rect 25585 2345 25590 2375
rect 25620 2370 25625 2375
rect 25780 2375 25820 2380
rect 25780 2370 25785 2375
rect 25620 2350 25785 2370
rect 25620 2345 25625 2350
rect 25585 2340 25625 2345
rect 25780 2345 25785 2350
rect 25815 2370 25820 2375
rect 26320 2375 26360 2380
rect 26320 2370 26325 2375
rect 25815 2350 26325 2370
rect 25815 2345 25820 2350
rect 25780 2340 25820 2345
rect 26320 2345 26325 2350
rect 26355 2345 26360 2375
rect 26320 2340 26360 2345
rect 27320 2375 27360 2380
rect 27320 2345 27325 2375
rect 27355 2370 27360 2375
rect 28015 2375 28055 2380
rect 28015 2370 28020 2375
rect 27355 2350 28020 2370
rect 27355 2345 27360 2350
rect 27320 2340 27360 2345
rect 28015 2345 28020 2350
rect 28050 2370 28055 2375
rect 28310 2375 28350 2380
rect 28310 2370 28315 2375
rect 28050 2350 28315 2370
rect 28050 2345 28055 2350
rect 28015 2340 28055 2345
rect 28310 2345 28315 2350
rect 28345 2345 28350 2375
rect 28310 2340 28350 2345
rect 2655 2320 3395 2340
rect 3625 2335 3665 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3625 2305 3630 2335
rect 3660 2330 3665 2335
rect 4345 2335 4385 2340
rect 4345 2330 4350 2335
rect 3660 2310 4350 2330
rect 3660 2305 3665 2310
rect 3625 2300 3665 2305
rect 4345 2305 4350 2310
rect 4380 2305 4385 2335
rect 16000 2325 16040 2330
rect 4345 2300 4385 2305
rect 14915 2315 14955 2320
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3445 2290 3485 2295
rect 3445 2285 3450 2290
rect 2770 2265 3450 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3445 2260 3450 2265
rect 3480 2285 3485 2290
rect 4525 2290 4565 2295
rect 4525 2285 4530 2290
rect 3480 2265 4530 2285
rect 3480 2260 3485 2265
rect 3445 2255 3485 2260
rect 4525 2260 4530 2265
rect 4560 2285 4565 2290
rect 5270 2290 5310 2295
rect 5270 2285 5275 2290
rect 4560 2265 5275 2285
rect 4560 2260 4565 2265
rect 4525 2255 4565 2260
rect 5270 2260 5275 2265
rect 5305 2260 5310 2290
rect 14915 2285 14920 2315
rect 14950 2310 14955 2315
rect 15115 2315 15155 2320
rect 15115 2310 15120 2315
rect 14950 2290 15120 2310
rect 14950 2285 14955 2290
rect 14915 2280 14955 2285
rect 15115 2285 15120 2290
rect 15150 2310 15155 2315
rect 15225 2315 15265 2320
rect 15225 2310 15230 2315
rect 15150 2290 15230 2310
rect 15150 2285 15155 2290
rect 15115 2280 15155 2285
rect 15225 2285 15230 2290
rect 15260 2310 15265 2315
rect 15335 2315 15375 2320
rect 15335 2310 15340 2315
rect 15260 2290 15340 2310
rect 15260 2285 15265 2290
rect 15225 2280 15265 2285
rect 15335 2285 15340 2290
rect 15370 2310 15375 2315
rect 15445 2315 15485 2320
rect 15445 2310 15450 2315
rect 15370 2290 15450 2310
rect 15370 2285 15375 2290
rect 15335 2280 15375 2285
rect 15445 2285 15450 2290
rect 15480 2310 15485 2315
rect 15555 2315 15595 2320
rect 15555 2310 15560 2315
rect 15480 2290 15560 2310
rect 15480 2285 15485 2290
rect 15445 2280 15485 2285
rect 15555 2285 15560 2290
rect 15590 2285 15595 2315
rect 16000 2295 16005 2325
rect 16035 2320 16040 2325
rect 17860 2325 17900 2330
rect 17860 2320 17865 2325
rect 16035 2300 17865 2320
rect 16035 2295 16040 2300
rect 16000 2290 16040 2295
rect 17860 2295 17865 2300
rect 17895 2295 17900 2325
rect 26000 2325 26040 2330
rect 17860 2290 17900 2295
rect 18255 2315 18295 2320
rect 18255 2285 18260 2315
rect 18290 2310 18295 2315
rect 18365 2315 18405 2320
rect 18365 2310 18370 2315
rect 18290 2290 18370 2310
rect 18290 2285 18295 2290
rect 15555 2280 15595 2285
rect 16440 2280 16480 2285
rect 5270 2255 5310 2260
rect 16440 2250 16445 2280
rect 16475 2275 16480 2280
rect 16660 2280 16700 2285
rect 16660 2275 16665 2280
rect 16475 2255 16665 2275
rect 16475 2250 16480 2255
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3805 2245 3845 2250
rect 16440 2245 16480 2250
rect 16660 2250 16665 2255
rect 16695 2275 16700 2280
rect 16880 2280 16920 2285
rect 16880 2275 16885 2280
rect 16695 2255 16885 2275
rect 16695 2250 16700 2255
rect 16660 2245 16700 2250
rect 16880 2250 16885 2255
rect 16915 2275 16920 2280
rect 17100 2280 17140 2285
rect 17100 2275 17105 2280
rect 16915 2255 17105 2275
rect 16915 2250 16920 2255
rect 16880 2245 16920 2250
rect 17100 2250 17105 2255
rect 17135 2275 17140 2280
rect 17320 2280 17360 2285
rect 18255 2280 18295 2285
rect 18365 2285 18370 2290
rect 18400 2310 18405 2315
rect 18475 2315 18515 2320
rect 18475 2310 18480 2315
rect 18400 2290 18480 2310
rect 18400 2285 18405 2290
rect 18365 2280 18405 2285
rect 18475 2285 18480 2290
rect 18510 2310 18515 2315
rect 18585 2315 18625 2320
rect 18585 2310 18590 2315
rect 18510 2290 18590 2310
rect 18510 2285 18515 2290
rect 18475 2280 18515 2285
rect 18585 2285 18590 2290
rect 18620 2310 18625 2315
rect 18695 2315 18735 2320
rect 18695 2310 18700 2315
rect 18620 2290 18700 2310
rect 18620 2285 18625 2290
rect 18585 2280 18625 2285
rect 18695 2285 18700 2290
rect 18730 2310 18735 2315
rect 18895 2315 18935 2320
rect 18895 2310 18900 2315
rect 18730 2290 18900 2310
rect 18730 2285 18735 2290
rect 18695 2280 18735 2285
rect 18895 2285 18900 2290
rect 18930 2285 18935 2315
rect 18895 2280 18935 2285
rect 24915 2315 24955 2320
rect 24915 2285 24920 2315
rect 24950 2310 24955 2315
rect 25115 2315 25155 2320
rect 25115 2310 25120 2315
rect 24950 2290 25120 2310
rect 24950 2285 24955 2290
rect 24915 2280 24955 2285
rect 25115 2285 25120 2290
rect 25150 2310 25155 2315
rect 25225 2315 25265 2320
rect 25225 2310 25230 2315
rect 25150 2290 25230 2310
rect 25150 2285 25155 2290
rect 25115 2280 25155 2285
rect 25225 2285 25230 2290
rect 25260 2310 25265 2315
rect 25335 2315 25375 2320
rect 25335 2310 25340 2315
rect 25260 2290 25340 2310
rect 25260 2285 25265 2290
rect 25225 2280 25265 2285
rect 25335 2285 25340 2290
rect 25370 2310 25375 2315
rect 25445 2315 25485 2320
rect 25445 2310 25450 2315
rect 25370 2290 25450 2310
rect 25370 2285 25375 2290
rect 25335 2280 25375 2285
rect 25445 2285 25450 2290
rect 25480 2310 25485 2315
rect 25555 2315 25595 2320
rect 25555 2310 25560 2315
rect 25480 2290 25560 2310
rect 25480 2285 25485 2290
rect 25445 2280 25485 2285
rect 25555 2285 25560 2290
rect 25590 2285 25595 2315
rect 26000 2295 26005 2325
rect 26035 2320 26040 2325
rect 27870 2325 27910 2330
rect 27870 2320 27875 2325
rect 26035 2300 27875 2320
rect 26035 2295 26040 2300
rect 26000 2290 26040 2295
rect 27870 2295 27875 2300
rect 27905 2295 27910 2325
rect 27870 2290 27910 2295
rect 28255 2295 28295 2300
rect 25555 2280 25595 2285
rect 26440 2280 26480 2285
rect 17320 2275 17325 2280
rect 17135 2255 17325 2275
rect 17135 2250 17140 2255
rect 17100 2245 17140 2250
rect 17320 2250 17325 2255
rect 17355 2250 17360 2280
rect 17320 2245 17360 2250
rect 26440 2250 26445 2280
rect 26475 2275 26480 2280
rect 26660 2280 26700 2285
rect 26660 2275 26665 2280
rect 26475 2255 26665 2275
rect 26475 2250 26480 2255
rect 26440 2245 26480 2250
rect 26660 2250 26665 2255
rect 26695 2275 26700 2280
rect 26880 2280 26920 2285
rect 26880 2275 26885 2280
rect 26695 2255 26885 2275
rect 26695 2250 26700 2255
rect 26660 2245 26700 2250
rect 26880 2250 26885 2255
rect 26915 2275 26920 2280
rect 27100 2280 27140 2285
rect 27100 2275 27105 2280
rect 26915 2255 27105 2275
rect 26915 2250 26920 2255
rect 26880 2245 26920 2250
rect 27100 2250 27105 2255
rect 27135 2275 27140 2280
rect 27320 2280 27360 2285
rect 27320 2275 27325 2280
rect 27135 2255 27325 2275
rect 27135 2250 27140 2255
rect 27100 2245 27140 2250
rect 27320 2250 27325 2255
rect 27355 2250 27360 2280
rect 28255 2265 28260 2295
rect 28290 2290 28295 2295
rect 28365 2295 28405 2300
rect 28365 2290 28370 2295
rect 28290 2270 28370 2290
rect 28290 2265 28295 2270
rect 28255 2260 28295 2265
rect 28365 2265 28370 2270
rect 28400 2290 28405 2295
rect 28475 2295 28515 2300
rect 28475 2290 28480 2295
rect 28400 2270 28480 2290
rect 28400 2265 28405 2270
rect 28365 2260 28405 2265
rect 28475 2265 28480 2270
rect 28510 2290 28515 2295
rect 28585 2295 28625 2300
rect 28585 2290 28590 2295
rect 28510 2270 28590 2290
rect 28510 2265 28515 2270
rect 28475 2260 28515 2265
rect 28585 2265 28590 2270
rect 28620 2290 28625 2295
rect 28695 2295 28735 2300
rect 28695 2290 28700 2295
rect 28620 2270 28700 2290
rect 28620 2265 28625 2270
rect 28585 2260 28625 2265
rect 28695 2265 28700 2270
rect 28730 2290 28735 2295
rect 28895 2295 28935 2300
rect 28895 2290 28900 2295
rect 28730 2270 28900 2290
rect 28730 2265 28735 2270
rect 28695 2260 28735 2265
rect 28895 2265 28900 2270
rect 28930 2265 28935 2295
rect 28895 2260 28935 2265
rect 27320 2245 27360 2250
rect 3805 2240 3810 2245
rect 2460 2220 3810 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3805 2215 3810 2220
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 16330 2235 16370 2240
rect 16330 2205 16335 2235
rect 16365 2230 16370 2235
rect 16550 2235 16590 2240
rect 16550 2230 16555 2235
rect 16365 2210 16555 2230
rect 16365 2205 16370 2210
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 3265 2200 3305 2205
rect 3265 2195 3270 2200
rect 2365 2175 3270 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 3265 2170 3270 2175
rect 3300 2195 3305 2200
rect 3985 2200 4025 2205
rect 3985 2195 3990 2200
rect 3300 2175 3990 2195
rect 3300 2170 3305 2175
rect 3265 2165 3305 2170
rect 3985 2170 3990 2175
rect 4020 2195 4025 2200
rect 4705 2200 4745 2205
rect 16330 2200 16370 2205
rect 16550 2205 16555 2210
rect 16585 2230 16590 2235
rect 16770 2235 16810 2240
rect 16770 2230 16775 2235
rect 16585 2210 16775 2230
rect 16585 2205 16590 2210
rect 16550 2200 16590 2205
rect 16770 2205 16775 2210
rect 16805 2230 16810 2235
rect 16990 2235 17030 2240
rect 16990 2230 16995 2235
rect 16805 2210 16995 2230
rect 16805 2205 16810 2210
rect 16770 2200 16810 2205
rect 16990 2205 16995 2210
rect 17025 2230 17030 2235
rect 17210 2235 17250 2240
rect 17210 2230 17215 2235
rect 17025 2210 17215 2230
rect 17025 2205 17030 2210
rect 16990 2200 17030 2205
rect 17210 2205 17215 2210
rect 17245 2230 17250 2235
rect 17430 2235 17470 2240
rect 17430 2230 17435 2235
rect 17245 2210 17435 2230
rect 17245 2205 17250 2210
rect 17210 2200 17250 2205
rect 17430 2205 17435 2210
rect 17465 2205 17470 2235
rect 17430 2200 17470 2205
rect 26330 2235 26370 2240
rect 26330 2205 26335 2235
rect 26365 2230 26370 2235
rect 26550 2235 26590 2240
rect 26550 2230 26555 2235
rect 26365 2210 26555 2230
rect 26365 2205 26370 2210
rect 26330 2200 26370 2205
rect 26550 2205 26555 2210
rect 26585 2230 26590 2235
rect 26770 2235 26810 2240
rect 26770 2230 26775 2235
rect 26585 2210 26775 2230
rect 26585 2205 26590 2210
rect 26550 2200 26590 2205
rect 26770 2205 26775 2210
rect 26805 2230 26810 2235
rect 26990 2235 27030 2240
rect 26990 2230 26995 2235
rect 26805 2210 26995 2230
rect 26805 2205 26810 2210
rect 26770 2200 26810 2205
rect 26990 2205 26995 2210
rect 27025 2230 27030 2235
rect 27210 2235 27250 2240
rect 27210 2230 27215 2235
rect 27025 2210 27215 2230
rect 27025 2205 27030 2210
rect 26990 2200 27030 2205
rect 27210 2205 27215 2210
rect 27245 2230 27250 2235
rect 27430 2235 27470 2240
rect 27430 2230 27435 2235
rect 27245 2210 27435 2230
rect 27245 2205 27250 2210
rect 27210 2200 27250 2205
rect 27430 2205 27435 2210
rect 27465 2205 27470 2235
rect 27430 2200 27470 2205
rect 4705 2195 4710 2200
rect 4020 2175 4710 2195
rect 4020 2170 4025 2175
rect 3985 2165 4025 2170
rect 4705 2170 4710 2175
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 15800 2180 15840 2185
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3625 2150 3665 2155
rect 15800 2150 15805 2180
rect 15835 2175 15840 2180
rect 16828 2180 16862 2185
rect 16828 2175 16831 2180
rect 15835 2155 16831 2175
rect 15835 2150 15840 2155
rect 3625 2145 3630 2150
rect 2415 2125 3630 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3625 2120 3630 2125
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2140 4125 2145
rect 5315 2145 5355 2150
rect 15800 2145 15840 2150
rect 16828 2150 16831 2155
rect 16859 2150 16862 2180
rect 16828 2145 16862 2150
rect 25800 2180 25840 2185
rect 25800 2150 25805 2180
rect 25835 2175 25840 2180
rect 26828 2180 26862 2185
rect 26828 2175 26831 2180
rect 25835 2155 26831 2175
rect 25835 2150 25840 2155
rect 25800 2145 25840 2150
rect 26828 2150 26831 2155
rect 26859 2150 26862 2180
rect 26828 2145 26862 2150
rect 5315 2140 5320 2145
rect 4120 2120 5320 2140
rect 4120 2115 4125 2120
rect 4085 2110 4125 2115
rect 5315 2115 5320 2120
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 14510 2110 14560 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2090 2785 2095
rect 2865 2095 2905 2100
rect 2865 2090 2870 2095
rect 2780 2070 2870 2090
rect 2780 2065 2785 2070
rect 2745 2060 2785 2065
rect 2865 2065 2870 2070
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2090 3865 2095
rect 3985 2095 4025 2100
rect 3985 2090 3990 2095
rect 3860 2070 3990 2090
rect 3860 2065 3865 2070
rect 3825 2060 3865 2065
rect 3985 2065 3990 2070
rect 4020 2090 4025 2095
rect 4145 2095 4185 2100
rect 4145 2090 4150 2095
rect 4020 2070 4150 2090
rect 4020 2065 4025 2070
rect 3985 2060 4025 2065
rect 4145 2065 4150 2070
rect 4180 2090 4185 2095
rect 4265 2095 4305 2100
rect 4265 2090 4270 2095
rect 4180 2070 4270 2090
rect 4180 2065 4185 2070
rect 4145 2060 4185 2065
rect 4265 2065 4270 2070
rect 4300 2090 4305 2095
rect 4385 2095 4425 2100
rect 4385 2090 4390 2095
rect 4300 2070 4390 2090
rect 4300 2065 4305 2070
rect 4265 2060 4305 2065
rect 4385 2065 4390 2070
rect 4420 2090 4425 2095
rect 4505 2095 4545 2100
rect 4505 2090 4510 2095
rect 4420 2070 4510 2090
rect 4420 2065 4425 2070
rect 4385 2060 4425 2065
rect 4505 2065 4510 2070
rect 4540 2090 4545 2095
rect 4625 2095 4665 2100
rect 4625 2090 4630 2095
rect 4540 2070 4630 2090
rect 4540 2065 4545 2070
rect 4505 2060 4545 2065
rect 4625 2065 4630 2070
rect 4660 2090 4665 2095
rect 4745 2095 4785 2100
rect 4745 2090 4750 2095
rect 4660 2070 4750 2090
rect 4660 2065 4665 2070
rect 4625 2060 4665 2065
rect 4745 2065 4750 2070
rect 4780 2090 4785 2095
rect 4865 2095 4905 2100
rect 4865 2090 4870 2095
rect 4780 2070 4870 2090
rect 4780 2065 4785 2070
rect 4745 2060 4785 2065
rect 4865 2065 4870 2070
rect 4900 2090 4905 2095
rect 4985 2095 5025 2100
rect 4985 2090 4990 2095
rect 4900 2070 4990 2090
rect 4900 2065 4905 2070
rect 4865 2060 4905 2065
rect 4985 2065 4990 2070
rect 5020 2090 5025 2095
rect 5105 2095 5145 2100
rect 5105 2090 5110 2095
rect 5020 2070 5110 2090
rect 5020 2065 5025 2070
rect 4985 2060 5025 2065
rect 5105 2065 5110 2070
rect 5140 2090 5145 2095
rect 5225 2095 5265 2100
rect 5225 2090 5230 2095
rect 5140 2070 5230 2090
rect 5140 2065 5145 2070
rect 5105 2060 5145 2065
rect 5225 2065 5230 2070
rect 5260 2090 5265 2095
rect 5550 2095 5590 2100
rect 5550 2090 5555 2095
rect 5260 2070 5555 2090
rect 5260 2065 5265 2070
rect 5225 2060 5265 2065
rect 5550 2065 5555 2070
rect 5585 2065 5590 2095
rect 14510 2080 14520 2110
rect 14550 2080 14560 2110
rect 14510 2070 14560 2080
rect 19240 2110 19290 2120
rect 19240 2080 19250 2110
rect 19280 2080 19290 2110
rect 19240 2070 19290 2080
rect 24510 2110 24560 2120
rect 24510 2080 24520 2110
rect 24550 2080 24560 2110
rect 24510 2070 24560 2080
rect 29390 2110 29440 2120
rect 29390 2080 29400 2110
rect 29430 2080 29440 2110
rect 29390 2070 29440 2080
rect 5550 2060 5590 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4085 2050 4125 2055
rect 4085 2020 4090 2050
rect 4120 2045 4125 2050
rect 4445 2050 4485 2055
rect 4445 2045 4450 2050
rect 4120 2025 4450 2045
rect 4120 2020 4125 2025
rect 4085 2015 4125 2020
rect 4445 2020 4450 2025
rect 4480 2045 4485 2050
rect 4805 2050 4845 2055
rect 4805 2045 4810 2050
rect 4480 2025 4810 2045
rect 4480 2020 4485 2025
rect 4445 2015 4485 2020
rect 4805 2020 4810 2025
rect 4840 2045 4845 2050
rect 5165 2050 5205 2055
rect 5165 2045 5170 2050
rect 4840 2025 5170 2045
rect 4840 2020 4845 2025
rect 4805 2015 4845 2020
rect 5165 2020 5170 2025
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 14640 2010 14675 2011
rect 14640 2005 14735 2010
rect 14675 1970 14700 2005
rect 14640 1965 14735 1970
rect 14760 2005 14795 2011
rect 14760 1965 14795 1970
rect 14820 2005 14855 2010
rect 18995 2005 19030 2010
rect 14870 2000 14910 2005
rect 14870 1995 14875 2000
rect 14855 1975 14875 1995
rect 14820 1965 14855 1970
rect 14870 1970 14875 1975
rect 14905 1970 14910 2000
rect 14870 1965 14910 1970
rect 18940 2000 18980 2005
rect 18940 1970 18945 2000
rect 18975 1995 18980 2000
rect 18975 1975 18995 1995
rect 18975 1970 18980 1975
rect 18940 1965 18980 1970
rect 18995 1965 19030 1970
rect 19055 2005 19090 2011
rect 19175 2010 19210 2011
rect 19055 1965 19090 1970
rect 19115 2005 19210 2010
rect 19150 1970 19175 2005
rect 19115 1965 19210 1970
rect 24640 2010 24675 2011
rect 24640 2005 24735 2010
rect 24675 1970 24700 2005
rect 24640 1965 24735 1970
rect 24760 2005 24795 2011
rect 24760 1965 24795 1970
rect 24820 2005 24855 2010
rect 24870 2000 24910 2005
rect 24870 1995 24875 2000
rect 24855 1975 24875 1995
rect 24820 1965 24855 1970
rect 24870 1970 24875 1975
rect 24905 1970 24910 2000
rect 29065 1985 29100 1990
rect 24870 1965 24910 1970
rect 28940 1980 28980 1985
rect 16385 1960 16425 1965
rect 14760 1945 14800 1950
rect 14760 1915 14765 1945
rect 14795 1940 14800 1945
rect 14915 1945 14955 1950
rect 14915 1940 14920 1945
rect 14795 1920 14920 1940
rect 14795 1915 14800 1920
rect 14760 1910 14800 1915
rect 14915 1915 14920 1920
rect 14950 1915 14955 1945
rect 14915 1910 14955 1915
rect 15060 1945 15100 1950
rect 15060 1915 15065 1945
rect 15095 1940 15100 1945
rect 15170 1945 15210 1950
rect 15170 1940 15175 1945
rect 15095 1920 15175 1940
rect 15095 1915 15100 1920
rect 15060 1910 15100 1915
rect 15170 1915 15175 1920
rect 15205 1940 15210 1945
rect 15280 1945 15320 1950
rect 15280 1940 15285 1945
rect 15205 1920 15285 1940
rect 15205 1915 15210 1920
rect 15170 1910 15210 1915
rect 15280 1915 15285 1920
rect 15315 1940 15320 1945
rect 15390 1945 15430 1950
rect 15390 1940 15395 1945
rect 15315 1920 15395 1940
rect 15315 1915 15320 1920
rect 15280 1910 15320 1915
rect 15390 1915 15395 1920
rect 15425 1940 15430 1945
rect 15500 1945 15540 1950
rect 15500 1940 15505 1945
rect 15425 1920 15505 1940
rect 15425 1915 15430 1920
rect 15390 1910 15430 1915
rect 15500 1915 15505 1920
rect 15535 1940 15540 1945
rect 15610 1945 15650 1950
rect 15610 1940 15615 1945
rect 15535 1920 15615 1940
rect 15535 1915 15540 1920
rect 15500 1910 15540 1915
rect 15610 1915 15615 1920
rect 15645 1915 15650 1945
rect 16385 1930 16390 1960
rect 16420 1955 16425 1960
rect 16605 1960 16645 1965
rect 16605 1955 16610 1960
rect 16420 1935 16610 1955
rect 16420 1930 16425 1935
rect 16385 1925 16425 1930
rect 16605 1930 16610 1935
rect 16640 1955 16645 1960
rect 16825 1960 16865 1965
rect 16825 1955 16830 1960
rect 16640 1935 16830 1955
rect 16640 1930 16645 1935
rect 16605 1925 16645 1930
rect 16825 1930 16830 1935
rect 16860 1955 16865 1960
rect 17045 1960 17085 1965
rect 17045 1955 17050 1960
rect 16860 1935 17050 1955
rect 16860 1930 16865 1935
rect 16825 1925 16865 1930
rect 17045 1930 17050 1935
rect 17080 1955 17085 1960
rect 17265 1960 17305 1965
rect 17265 1955 17270 1960
rect 17080 1935 17270 1955
rect 17080 1930 17085 1935
rect 17045 1925 17085 1930
rect 17265 1930 17270 1935
rect 17300 1930 17305 1960
rect 26385 1960 26425 1965
rect 17265 1925 17305 1930
rect 18200 1945 18240 1950
rect 15610 1910 15650 1915
rect 18200 1915 18205 1945
rect 18235 1940 18240 1945
rect 18310 1945 18350 1950
rect 18310 1940 18315 1945
rect 18235 1920 18315 1940
rect 18235 1915 18240 1920
rect 18200 1910 18240 1915
rect 18310 1915 18315 1920
rect 18345 1940 18350 1945
rect 18420 1945 18460 1950
rect 18420 1940 18425 1945
rect 18345 1920 18425 1940
rect 18345 1915 18350 1920
rect 18310 1910 18350 1915
rect 18420 1915 18425 1920
rect 18455 1940 18460 1945
rect 18530 1945 18570 1950
rect 18530 1940 18535 1945
rect 18455 1920 18535 1940
rect 18455 1915 18460 1920
rect 18420 1910 18460 1915
rect 18530 1915 18535 1920
rect 18565 1940 18570 1945
rect 18640 1945 18680 1950
rect 18640 1940 18645 1945
rect 18565 1920 18645 1940
rect 18565 1915 18570 1920
rect 18530 1910 18570 1915
rect 18640 1915 18645 1920
rect 18675 1940 18680 1945
rect 18750 1945 18790 1950
rect 18750 1940 18755 1945
rect 18675 1920 18755 1940
rect 18675 1915 18680 1920
rect 18640 1910 18680 1915
rect 18750 1915 18755 1920
rect 18785 1915 18790 1945
rect 18750 1910 18790 1915
rect 18895 1945 18935 1950
rect 18895 1915 18900 1945
rect 18930 1940 18935 1945
rect 19050 1945 19090 1950
rect 19050 1940 19055 1945
rect 18930 1920 19055 1940
rect 18930 1915 18935 1920
rect 18895 1910 18935 1915
rect 19050 1915 19055 1920
rect 19085 1915 19090 1945
rect 19050 1910 19090 1915
rect 24760 1945 24800 1950
rect 24760 1915 24765 1945
rect 24795 1940 24800 1945
rect 24915 1945 24955 1950
rect 24915 1940 24920 1945
rect 24795 1920 24920 1940
rect 24795 1915 24800 1920
rect 24760 1910 24800 1915
rect 24915 1915 24920 1920
rect 24950 1915 24955 1945
rect 24915 1910 24955 1915
rect 25060 1945 25100 1950
rect 25060 1915 25065 1945
rect 25095 1940 25100 1945
rect 25170 1945 25210 1950
rect 25170 1940 25175 1945
rect 25095 1920 25175 1940
rect 25095 1915 25100 1920
rect 25060 1910 25100 1915
rect 25170 1915 25175 1920
rect 25205 1940 25210 1945
rect 25280 1945 25320 1950
rect 25280 1940 25285 1945
rect 25205 1920 25285 1940
rect 25205 1915 25210 1920
rect 25170 1910 25210 1915
rect 25280 1915 25285 1920
rect 25315 1940 25320 1945
rect 25390 1945 25430 1950
rect 25390 1940 25395 1945
rect 25315 1920 25395 1940
rect 25315 1915 25320 1920
rect 25280 1910 25320 1915
rect 25390 1915 25395 1920
rect 25425 1940 25430 1945
rect 25500 1945 25540 1950
rect 25500 1940 25505 1945
rect 25425 1920 25505 1940
rect 25425 1915 25430 1920
rect 25390 1910 25430 1915
rect 25500 1915 25505 1920
rect 25535 1940 25540 1945
rect 25610 1945 25650 1950
rect 25610 1940 25615 1945
rect 25535 1920 25615 1940
rect 25535 1915 25540 1920
rect 25500 1910 25540 1915
rect 25610 1915 25615 1920
rect 25645 1915 25650 1945
rect 26385 1930 26390 1960
rect 26420 1955 26425 1960
rect 26605 1960 26645 1965
rect 26605 1955 26610 1960
rect 26420 1935 26610 1955
rect 26420 1930 26425 1935
rect 26385 1925 26425 1930
rect 26605 1930 26610 1935
rect 26640 1955 26645 1960
rect 26825 1960 26865 1965
rect 26825 1955 26830 1960
rect 26640 1935 26830 1955
rect 26640 1930 26645 1935
rect 26605 1925 26645 1930
rect 26825 1930 26830 1935
rect 26860 1955 26865 1960
rect 27045 1960 27085 1965
rect 27045 1955 27050 1960
rect 26860 1935 27050 1955
rect 26860 1930 26865 1935
rect 26825 1925 26865 1930
rect 27045 1930 27050 1935
rect 27080 1955 27085 1960
rect 27265 1960 27305 1965
rect 27265 1955 27270 1960
rect 27080 1935 27270 1955
rect 27080 1930 27085 1935
rect 27045 1925 27085 1930
rect 27265 1930 27270 1935
rect 27300 1930 27305 1960
rect 28940 1950 28945 1980
rect 28975 1975 28980 1980
rect 28975 1955 29065 1975
rect 28975 1950 28980 1955
rect 28940 1945 28980 1950
rect 29065 1945 29100 1950
rect 29125 1985 29160 1991
rect 29245 1990 29280 1991
rect 29125 1945 29160 1950
rect 29185 1985 29280 1990
rect 29220 1950 29245 1985
rect 29185 1945 29280 1950
rect 27265 1925 27305 1930
rect 28200 1925 28240 1930
rect 25610 1910 25650 1915
rect 16495 1905 16535 1910
rect 14640 1895 14680 1900
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4205 1845 4245 1885
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1875 4365 1880
rect 4565 1875 4605 1885
rect 4685 1880 4725 1885
rect 4685 1875 4690 1880
rect 4360 1855 4690 1875
rect 4360 1850 4365 1855
rect 4325 1845 4365 1850
rect 4565 1845 4605 1855
rect 4685 1850 4690 1855
rect 4720 1875 4725 1880
rect 4925 1875 4965 1885
rect 5045 1880 5085 1885
rect 5045 1875 5050 1880
rect 4720 1855 5050 1875
rect 4720 1850 4725 1855
rect 4685 1845 4725 1850
rect 4925 1845 4965 1855
rect 5045 1850 5050 1855
rect 5080 1875 5085 1880
rect 5080 1855 5175 1875
rect 14640 1865 14645 1895
rect 14675 1890 14680 1895
rect 16000 1895 16040 1900
rect 16000 1890 16005 1895
rect 14675 1870 16005 1890
rect 14675 1865 14680 1870
rect 14640 1860 14680 1865
rect 16000 1865 16005 1870
rect 16035 1865 16040 1895
rect 16495 1875 16500 1905
rect 16530 1900 16535 1905
rect 16715 1905 16755 1910
rect 16715 1900 16720 1905
rect 16530 1880 16720 1900
rect 16530 1875 16535 1880
rect 16495 1870 16535 1875
rect 16715 1875 16720 1880
rect 16750 1900 16755 1905
rect 16935 1905 16975 1910
rect 16935 1900 16940 1905
rect 16750 1880 16940 1900
rect 16750 1875 16755 1880
rect 16715 1870 16755 1875
rect 16935 1875 16940 1880
rect 16970 1900 16975 1905
rect 17155 1905 17195 1910
rect 17155 1900 17160 1905
rect 16970 1880 17160 1900
rect 16970 1875 16975 1880
rect 16935 1870 16975 1875
rect 17155 1875 17160 1880
rect 17190 1900 17195 1905
rect 17375 1905 17415 1910
rect 17375 1900 17380 1905
rect 17190 1880 17380 1900
rect 17190 1875 17195 1880
rect 17155 1870 17195 1875
rect 17375 1875 17380 1880
rect 17410 1875 17415 1905
rect 26495 1905 26535 1910
rect 17375 1870 17415 1875
rect 17860 1895 17900 1900
rect 16000 1860 16040 1865
rect 17860 1865 17865 1895
rect 17895 1890 17900 1895
rect 19170 1895 19210 1900
rect 19170 1890 19175 1895
rect 17895 1870 19175 1890
rect 17895 1865 17900 1870
rect 17860 1860 17900 1865
rect 19170 1865 19175 1870
rect 19205 1865 19210 1895
rect 19170 1860 19210 1865
rect 24640 1895 24680 1900
rect 24640 1865 24645 1895
rect 24675 1890 24680 1895
rect 26000 1895 26040 1900
rect 26000 1890 26005 1895
rect 24675 1870 26005 1890
rect 24675 1865 24680 1870
rect 24640 1860 24680 1865
rect 26000 1865 26005 1870
rect 26035 1865 26040 1895
rect 26495 1875 26500 1905
rect 26530 1900 26535 1905
rect 26715 1905 26755 1910
rect 26715 1900 26720 1905
rect 26530 1880 26720 1900
rect 26530 1875 26535 1880
rect 26495 1870 26535 1875
rect 26715 1875 26720 1880
rect 26750 1900 26755 1905
rect 26935 1905 26975 1910
rect 26935 1900 26940 1905
rect 26750 1880 26940 1900
rect 26750 1875 26755 1880
rect 26715 1870 26755 1875
rect 26935 1875 26940 1880
rect 26970 1900 26975 1905
rect 27155 1905 27195 1910
rect 27155 1900 27160 1905
rect 26970 1880 27160 1900
rect 26970 1875 26975 1880
rect 26935 1870 26975 1875
rect 27155 1875 27160 1880
rect 27190 1900 27195 1905
rect 27375 1905 27415 1910
rect 27375 1900 27380 1905
rect 27190 1880 27380 1900
rect 27190 1875 27195 1880
rect 27155 1870 27195 1875
rect 27375 1875 27380 1880
rect 27410 1875 27415 1905
rect 28200 1895 28205 1925
rect 28235 1920 28240 1925
rect 28310 1925 28350 1930
rect 28310 1920 28315 1925
rect 28235 1900 28315 1920
rect 28235 1895 28240 1900
rect 28200 1890 28240 1895
rect 28310 1895 28315 1900
rect 28345 1920 28350 1925
rect 28420 1925 28460 1930
rect 28420 1920 28425 1925
rect 28345 1900 28425 1920
rect 28345 1895 28350 1900
rect 28310 1890 28350 1895
rect 28420 1895 28425 1900
rect 28455 1920 28460 1925
rect 28530 1925 28570 1930
rect 28530 1920 28535 1925
rect 28455 1900 28535 1920
rect 28455 1895 28460 1900
rect 28420 1890 28460 1895
rect 28530 1895 28535 1900
rect 28565 1920 28570 1925
rect 28640 1925 28680 1930
rect 28640 1920 28645 1925
rect 28565 1900 28645 1920
rect 28565 1895 28570 1900
rect 28530 1890 28570 1895
rect 28640 1895 28645 1900
rect 28675 1920 28680 1925
rect 28750 1925 28790 1930
rect 28750 1920 28755 1925
rect 28675 1900 28755 1920
rect 28675 1895 28680 1900
rect 28640 1890 28680 1895
rect 28750 1895 28755 1900
rect 28785 1895 28790 1925
rect 28750 1890 28790 1895
rect 28895 1925 28935 1930
rect 28895 1895 28900 1925
rect 28930 1920 28935 1925
rect 29120 1925 29160 1930
rect 29120 1920 29125 1925
rect 28930 1900 29125 1920
rect 28930 1895 28935 1900
rect 28895 1890 28935 1895
rect 29120 1895 29125 1900
rect 29155 1895 29160 1925
rect 29120 1890 29160 1895
rect 27375 1870 27415 1875
rect 27870 1875 27910 1880
rect 26000 1860 26040 1865
rect 5080 1850 5085 1855
rect 5045 1845 5085 1850
rect 16190 1850 16230 1855
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1815 4155 1820
rect 4205 1820 4245 1825
rect 4205 1815 4210 1820
rect 4150 1795 4210 1815
rect 4150 1790 4155 1795
rect 4115 1785 4155 1790
rect 4205 1790 4210 1795
rect 4240 1815 4245 1820
rect 4445 1820 4485 1825
rect 4445 1815 4450 1820
rect 4240 1795 4450 1815
rect 4240 1790 4245 1795
rect 4205 1785 4245 1790
rect 4445 1790 4450 1795
rect 4480 1815 4485 1820
rect 4565 1820 4605 1825
rect 4565 1815 4570 1820
rect 4480 1795 4570 1815
rect 4480 1790 4485 1795
rect 4445 1785 4485 1790
rect 4565 1790 4570 1795
rect 4600 1815 4605 1820
rect 4805 1820 4845 1825
rect 4805 1815 4810 1820
rect 4600 1795 4810 1815
rect 4600 1790 4605 1795
rect 4565 1785 4605 1790
rect 4805 1790 4810 1795
rect 4840 1815 4845 1820
rect 4925 1820 4965 1825
rect 4925 1815 4930 1820
rect 4840 1795 4930 1815
rect 4840 1790 4845 1795
rect 4805 1785 4845 1790
rect 4925 1790 4930 1795
rect 4960 1815 4965 1820
rect 5135 1820 5175 1825
rect 5135 1815 5140 1820
rect 4960 1795 5140 1815
rect 4960 1790 4965 1795
rect 4925 1785 4965 1790
rect 5135 1790 5140 1795
rect 5170 1815 5175 1820
rect 5360 1820 5400 1825
rect 5360 1815 5365 1820
rect 5170 1795 5365 1815
rect 5170 1790 5175 1795
rect 5135 1785 5175 1790
rect 5360 1790 5365 1795
rect 5395 1790 5400 1820
rect 16190 1820 16195 1850
rect 16225 1845 16230 1850
rect 16410 1850 16450 1855
rect 16410 1845 16415 1850
rect 16225 1825 16415 1845
rect 16225 1820 16230 1825
rect 16190 1815 16230 1820
rect 16410 1820 16415 1825
rect 16445 1845 16450 1850
rect 16640 1850 16680 1855
rect 16640 1845 16645 1850
rect 16445 1825 16645 1845
rect 16445 1820 16450 1825
rect 16410 1815 16450 1820
rect 16640 1820 16645 1825
rect 16675 1845 16680 1850
rect 17230 1850 17270 1855
rect 17230 1845 17235 1850
rect 16675 1825 17235 1845
rect 16675 1820 16680 1825
rect 16640 1815 16680 1820
rect 17230 1820 17235 1825
rect 17265 1845 17270 1850
rect 17450 1850 17490 1855
rect 17450 1845 17455 1850
rect 17265 1825 17455 1845
rect 17265 1820 17270 1825
rect 17230 1815 17270 1820
rect 17450 1820 17455 1825
rect 17485 1845 17490 1850
rect 17680 1850 17720 1855
rect 17680 1845 17685 1850
rect 17485 1825 17685 1845
rect 17485 1820 17490 1825
rect 17450 1815 17490 1820
rect 17680 1820 17685 1825
rect 17715 1820 17720 1850
rect 17680 1815 17720 1820
rect 26190 1850 26230 1855
rect 26190 1820 26195 1850
rect 26225 1845 26230 1850
rect 26410 1850 26450 1855
rect 26410 1845 26415 1850
rect 26225 1825 26415 1845
rect 26225 1820 26230 1825
rect 26190 1815 26230 1820
rect 26410 1820 26415 1825
rect 26445 1845 26450 1850
rect 26640 1850 26680 1855
rect 26640 1845 26645 1850
rect 26445 1825 26645 1845
rect 26445 1820 26450 1825
rect 26410 1815 26450 1820
rect 26640 1820 26645 1825
rect 26675 1845 26680 1850
rect 27230 1850 27270 1855
rect 27230 1845 27235 1850
rect 26675 1825 27235 1845
rect 26675 1820 26680 1825
rect 26640 1815 26680 1820
rect 27230 1820 27235 1825
rect 27265 1845 27270 1850
rect 27450 1850 27490 1855
rect 27450 1845 27455 1850
rect 27265 1825 27455 1845
rect 27265 1820 27270 1825
rect 27230 1815 27270 1820
rect 27450 1820 27455 1825
rect 27485 1845 27490 1850
rect 27680 1850 27720 1855
rect 27680 1845 27685 1850
rect 27485 1825 27685 1845
rect 27485 1820 27490 1825
rect 27450 1815 27490 1820
rect 27680 1820 27685 1825
rect 27715 1820 27720 1850
rect 27870 1845 27875 1875
rect 27905 1870 27910 1875
rect 29240 1875 29280 1880
rect 29240 1870 29245 1875
rect 27905 1850 29245 1870
rect 27905 1845 27910 1850
rect 27870 1840 27910 1845
rect 29240 1845 29245 1850
rect 29275 1845 29280 1875
rect 29240 1840 29280 1845
rect 27680 1815 27720 1820
rect 5360 1785 5400 1790
rect 16820 1805 16860 1810
rect 16820 1775 16825 1805
rect 16855 1800 16860 1805
rect 16940 1805 16980 1810
rect 16940 1800 16945 1805
rect 16855 1780 16945 1800
rect 16855 1775 16860 1780
rect 16820 1770 16860 1775
rect 16940 1775 16945 1780
rect 16975 1775 16980 1805
rect 16940 1770 16980 1775
rect 26820 1805 26860 1810
rect 26820 1775 26825 1805
rect 26855 1800 26860 1805
rect 26940 1805 26980 1810
rect 26940 1800 26945 1805
rect 26855 1780 26945 1800
rect 26855 1775 26860 1780
rect 26820 1770 26860 1775
rect 26940 1775 26945 1780
rect 26975 1775 26980 1805
rect 26940 1770 26980 1775
rect 2800 1765 2840 1770
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 2800 1755 2805 1765
rect 2710 1735 2805 1755
rect 2835 1755 2840 1765
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2835 1735 3230 1755
rect 2710 1730 2715 1735
rect 2800 1730 2840 1735
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1755 4245 1760
rect 4445 1760 4485 1765
rect 4445 1755 4450 1760
rect 4240 1735 4450 1755
rect 4240 1730 4245 1735
rect 4205 1725 4245 1730
rect 4445 1730 4450 1735
rect 4480 1755 4485 1760
rect 4685 1760 4725 1765
rect 4685 1755 4690 1760
rect 4480 1735 4690 1755
rect 4480 1730 4485 1735
rect 4445 1725 4485 1730
rect 4685 1730 4690 1735
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1755 4785 1760
rect 5270 1760 5310 1765
rect 5270 1755 5275 1760
rect 4780 1735 5275 1755
rect 4780 1730 4785 1735
rect 4745 1725 4785 1730
rect 5270 1730 5275 1735
rect 5305 1755 5310 1760
rect 14815 1760 14855 1765
rect 5305 1735 6100 1755
rect 5305 1730 5310 1735
rect 5270 1725 5310 1730
rect 14815 1730 14820 1760
rect 14850 1755 14855 1760
rect 15405 1760 15445 1765
rect 15405 1755 15410 1760
rect 14850 1735 15410 1755
rect 14850 1730 14855 1735
rect 14815 1725 14855 1730
rect 15405 1730 15410 1735
rect 15440 1755 15445 1760
rect 15735 1760 15775 1765
rect 15735 1755 15740 1760
rect 15440 1735 15740 1755
rect 15440 1730 15445 1735
rect 15405 1725 15445 1730
rect 15735 1730 15740 1735
rect 15770 1730 15775 1760
rect 15735 1725 15775 1730
rect 16085 1760 16125 1765
rect 16085 1730 16090 1760
rect 16120 1755 16125 1760
rect 16305 1760 16345 1765
rect 16305 1755 16310 1760
rect 16120 1735 16310 1755
rect 16120 1730 16125 1735
rect 16085 1725 16125 1730
rect 16305 1730 16310 1735
rect 16340 1755 16345 1760
rect 16525 1760 16565 1765
rect 16525 1755 16530 1760
rect 16340 1735 16530 1755
rect 16340 1730 16345 1735
rect 16305 1725 16345 1730
rect 16525 1730 16530 1735
rect 16560 1755 16565 1760
rect 17125 1760 17165 1765
rect 17125 1755 17130 1760
rect 16560 1735 17130 1755
rect 16560 1730 16565 1735
rect 16525 1725 16565 1730
rect 17125 1730 17130 1735
rect 17160 1755 17165 1760
rect 17345 1760 17385 1765
rect 17345 1755 17350 1760
rect 17160 1735 17350 1755
rect 17160 1730 17165 1735
rect 17125 1725 17165 1730
rect 17345 1730 17350 1735
rect 17380 1755 17385 1760
rect 17565 1760 17605 1765
rect 17565 1755 17570 1760
rect 17380 1735 17570 1755
rect 17380 1730 17385 1735
rect 17345 1725 17385 1730
rect 17565 1730 17570 1735
rect 17600 1730 17605 1760
rect 17565 1725 17605 1730
rect 18075 1760 18115 1765
rect 18075 1730 18080 1760
rect 18110 1755 18115 1760
rect 18405 1760 18445 1765
rect 18405 1755 18410 1760
rect 18110 1735 18410 1755
rect 18110 1730 18115 1735
rect 18075 1725 18115 1730
rect 18405 1730 18410 1735
rect 18440 1755 18445 1760
rect 18995 1760 19035 1765
rect 18995 1755 19000 1760
rect 18440 1735 19000 1755
rect 18440 1730 18445 1735
rect 18405 1725 18445 1730
rect 18995 1730 19000 1735
rect 19030 1730 19035 1760
rect 18995 1725 19035 1730
rect 24815 1760 24855 1765
rect 24815 1730 24820 1760
rect 24850 1755 24855 1760
rect 25405 1760 25445 1765
rect 25405 1755 25410 1760
rect 24850 1735 25410 1755
rect 24850 1730 24855 1735
rect 24815 1725 24855 1730
rect 25405 1730 25410 1735
rect 25440 1755 25445 1760
rect 25735 1760 25775 1765
rect 25735 1755 25740 1760
rect 25440 1735 25740 1755
rect 25440 1730 25445 1735
rect 25405 1725 25445 1730
rect 25735 1730 25740 1735
rect 25770 1730 25775 1760
rect 25735 1725 25775 1730
rect 26085 1760 26125 1765
rect 26085 1730 26090 1760
rect 26120 1755 26125 1760
rect 26305 1760 26345 1765
rect 26305 1755 26310 1760
rect 26120 1735 26310 1755
rect 26120 1730 26125 1735
rect 26085 1725 26125 1730
rect 26305 1730 26310 1735
rect 26340 1755 26345 1760
rect 26525 1760 26565 1765
rect 26525 1755 26530 1760
rect 26340 1735 26530 1755
rect 26340 1730 26345 1735
rect 26305 1725 26345 1730
rect 26525 1730 26530 1735
rect 26560 1755 26565 1760
rect 27125 1760 27165 1765
rect 27125 1755 27130 1760
rect 26560 1735 27130 1755
rect 26560 1730 26565 1735
rect 26525 1725 26565 1730
rect 27125 1730 27130 1735
rect 27160 1755 27165 1760
rect 27345 1760 27385 1765
rect 27345 1755 27350 1760
rect 27160 1735 27350 1755
rect 27160 1730 27165 1735
rect 27125 1725 27165 1730
rect 27345 1730 27350 1735
rect 27380 1755 27385 1760
rect 27565 1760 27605 1765
rect 27565 1755 27570 1760
rect 27380 1735 27570 1755
rect 27380 1730 27385 1735
rect 27345 1725 27385 1730
rect 27565 1730 27570 1735
rect 27600 1730 27605 1760
rect 27565 1725 27605 1730
rect 28025 1760 28065 1765
rect 28025 1730 28030 1760
rect 28060 1755 28065 1760
rect 28405 1760 28445 1765
rect 28405 1755 28410 1760
rect 28060 1735 28410 1755
rect 28060 1730 28065 1735
rect 28025 1725 28065 1730
rect 28405 1730 28410 1735
rect 28440 1755 28445 1760
rect 29115 1760 29155 1765
rect 29115 1755 29120 1760
rect 28440 1735 29120 1755
rect 28440 1730 28445 1735
rect 28405 1725 28445 1730
rect 29115 1730 29120 1735
rect 29150 1730 29155 1760
rect 29115 1725 29155 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2800 1710 2840 1715
rect 2800 1705 2805 1710
rect 1297 1685 2805 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2800 1680 2805 1685
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1710 4365 1715
rect 4565 1715 4605 1720
rect 4565 1710 4570 1715
rect 4360 1690 4570 1710
rect 4360 1685 4365 1690
rect 4325 1680 4365 1685
rect 4565 1685 4570 1690
rect 4600 1710 4605 1715
rect 4805 1715 4845 1720
rect 4805 1710 4810 1715
rect 4600 1690 4810 1710
rect 4600 1685 4605 1690
rect 4565 1680 4605 1685
rect 4805 1685 4810 1690
rect 4840 1685 4845 1715
rect 16237 1715 16269 1720
rect 16237 1710 16240 1715
rect 4805 1680 4845 1685
rect 14515 1705 14555 1710
rect 2800 1675 2840 1680
rect 14515 1675 14520 1705
rect 14550 1700 14555 1705
rect 14880 1705 14920 1710
rect 14880 1700 14885 1705
rect 14550 1680 14885 1700
rect 14550 1675 14555 1680
rect 14515 1670 14555 1675
rect 14880 1675 14885 1680
rect 14915 1700 14920 1705
rect 15105 1705 15145 1710
rect 15105 1700 15110 1705
rect 14915 1680 15110 1700
rect 14915 1675 14920 1680
rect 14880 1670 14920 1675
rect 15105 1675 15110 1680
rect 15140 1700 15145 1705
rect 15305 1705 15345 1710
rect 15305 1700 15310 1705
rect 15140 1680 15310 1700
rect 15140 1675 15145 1680
rect 15105 1670 15145 1675
rect 15305 1675 15310 1680
rect 15340 1700 15345 1705
rect 15505 1705 15545 1710
rect 15505 1700 15510 1705
rect 15340 1680 15510 1700
rect 15340 1675 15345 1680
rect 15305 1670 15345 1675
rect 15505 1675 15510 1680
rect 15540 1675 15545 1705
rect 15940 1690 16240 1710
rect 16237 1685 16240 1690
rect 16266 1710 16269 1715
rect 16457 1715 16489 1720
rect 16457 1710 16460 1715
rect 16266 1690 16460 1710
rect 16266 1685 16269 1690
rect 16237 1680 16269 1685
rect 16457 1685 16460 1690
rect 16486 1710 16489 1715
rect 16601 1715 16633 1720
rect 16601 1710 16604 1715
rect 16486 1690 16604 1710
rect 16486 1685 16489 1690
rect 16457 1680 16489 1685
rect 16601 1685 16604 1690
rect 16630 1710 16633 1715
rect 16867 1715 16899 1720
rect 16867 1710 16870 1715
rect 16630 1690 16870 1710
rect 16630 1685 16633 1690
rect 16601 1680 16633 1685
rect 16867 1685 16870 1690
rect 16896 1710 16899 1715
rect 17277 1715 17309 1720
rect 17277 1710 17280 1715
rect 16896 1690 17280 1710
rect 16896 1685 16899 1690
rect 16867 1680 16899 1685
rect 17277 1685 17280 1690
rect 17306 1710 17309 1715
rect 17497 1715 17529 1720
rect 17497 1710 17500 1715
rect 17306 1690 17500 1710
rect 17306 1685 17309 1690
rect 17277 1680 17309 1685
rect 17497 1685 17500 1690
rect 17526 1710 17529 1715
rect 17641 1715 17673 1720
rect 17641 1710 17644 1715
rect 17526 1690 17644 1710
rect 17526 1685 17529 1690
rect 17497 1680 17529 1685
rect 17641 1685 17644 1690
rect 17670 1685 17673 1715
rect 26237 1715 26269 1720
rect 26237 1710 26240 1715
rect 17641 1680 17673 1685
rect 18305 1705 18345 1710
rect 15505 1670 15545 1675
rect 18305 1675 18310 1705
rect 18340 1700 18345 1705
rect 18505 1705 18545 1710
rect 18505 1700 18510 1705
rect 18340 1680 18510 1700
rect 18340 1675 18345 1680
rect 18305 1670 18345 1675
rect 18505 1675 18510 1680
rect 18540 1700 18545 1705
rect 18705 1705 18745 1710
rect 18705 1700 18710 1705
rect 18540 1680 18710 1700
rect 18540 1675 18545 1680
rect 18505 1670 18545 1675
rect 18705 1675 18710 1680
rect 18740 1700 18745 1705
rect 18930 1705 18970 1710
rect 18930 1700 18935 1705
rect 18740 1680 18935 1700
rect 18740 1675 18745 1680
rect 18705 1670 18745 1675
rect 18930 1675 18935 1680
rect 18965 1700 18970 1705
rect 19245 1705 19285 1710
rect 19245 1700 19250 1705
rect 18965 1680 19250 1700
rect 18965 1675 18970 1680
rect 18930 1670 18970 1675
rect 19245 1675 19250 1680
rect 19280 1675 19285 1705
rect 19245 1670 19285 1675
rect 24515 1705 24555 1710
rect 24515 1675 24520 1705
rect 24550 1700 24555 1705
rect 24880 1705 24920 1710
rect 24880 1700 24885 1705
rect 24550 1680 24885 1700
rect 24550 1675 24555 1680
rect 24515 1670 24555 1675
rect 24880 1675 24885 1680
rect 24915 1700 24920 1705
rect 25105 1705 25145 1710
rect 25105 1700 25110 1705
rect 24915 1680 25110 1700
rect 24915 1675 24920 1680
rect 24880 1670 24920 1675
rect 25105 1675 25110 1680
rect 25140 1700 25145 1705
rect 25305 1705 25345 1710
rect 25305 1700 25310 1705
rect 25140 1680 25310 1700
rect 25140 1675 25145 1680
rect 25105 1670 25145 1675
rect 25305 1675 25310 1680
rect 25340 1700 25345 1705
rect 25505 1705 25545 1710
rect 25505 1700 25510 1705
rect 25340 1680 25510 1700
rect 25340 1675 25345 1680
rect 25305 1670 25345 1675
rect 25505 1675 25510 1680
rect 25540 1675 25545 1705
rect 25940 1690 26240 1710
rect 26237 1685 26240 1690
rect 26266 1710 26269 1715
rect 26457 1715 26489 1720
rect 26457 1710 26460 1715
rect 26266 1690 26460 1710
rect 26266 1685 26269 1690
rect 26237 1680 26269 1685
rect 26457 1685 26460 1690
rect 26486 1710 26489 1715
rect 26601 1715 26633 1720
rect 26601 1710 26604 1715
rect 26486 1690 26604 1710
rect 26486 1685 26489 1690
rect 26457 1680 26489 1685
rect 26601 1685 26604 1690
rect 26630 1710 26633 1715
rect 26867 1715 26899 1720
rect 26867 1710 26870 1715
rect 26630 1690 26870 1710
rect 26630 1685 26633 1690
rect 26601 1680 26633 1685
rect 26867 1685 26870 1690
rect 26896 1710 26899 1715
rect 27277 1715 27309 1720
rect 27277 1710 27280 1715
rect 26896 1690 27280 1710
rect 26896 1685 26899 1690
rect 26867 1680 26899 1685
rect 27277 1685 27280 1690
rect 27306 1710 27309 1715
rect 27497 1715 27529 1720
rect 27497 1710 27500 1715
rect 27306 1690 27500 1710
rect 27306 1685 27309 1690
rect 27277 1680 27309 1685
rect 27497 1685 27500 1690
rect 27526 1710 27529 1715
rect 27641 1715 27673 1720
rect 27641 1710 27644 1715
rect 27526 1690 27644 1710
rect 27526 1685 27529 1690
rect 27497 1680 27529 1685
rect 27641 1685 27644 1690
rect 27670 1685 27673 1715
rect 27641 1680 27673 1685
rect 28305 1705 28345 1710
rect 25505 1670 25545 1675
rect 28305 1675 28310 1705
rect 28340 1700 28345 1705
rect 28505 1705 28545 1710
rect 28505 1700 28510 1705
rect 28340 1680 28510 1700
rect 28340 1675 28345 1680
rect 28305 1670 28345 1675
rect 28505 1675 28510 1680
rect 28540 1700 28545 1705
rect 28705 1705 28745 1710
rect 28705 1700 28710 1705
rect 28540 1680 28710 1700
rect 28540 1675 28545 1680
rect 28505 1670 28545 1675
rect 28705 1675 28710 1680
rect 28740 1700 28745 1705
rect 29050 1705 29090 1710
rect 29050 1700 29055 1705
rect 28740 1680 29055 1700
rect 28740 1675 28745 1680
rect 28705 1670 28745 1675
rect 29050 1675 29055 1680
rect 29085 1700 29090 1705
rect 29395 1705 29435 1710
rect 29395 1700 29400 1705
rect 29085 1680 29400 1700
rect 29085 1675 29090 1680
rect 29050 1670 29090 1675
rect 29395 1675 29400 1680
rect 29430 1675 29435 1705
rect 29395 1670 29435 1675
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 14820 1645 14855 1650
rect 14820 1605 14855 1610
rect 14880 1645 14915 1650
rect 14880 1605 14915 1610
rect 18935 1645 18970 1650
rect 18935 1605 18970 1610
rect 18995 1645 19030 1650
rect 18995 1605 19030 1610
rect 24820 1645 24855 1650
rect 24820 1605 24855 1610
rect 24880 1645 24915 1650
rect 24880 1605 24915 1610
rect 29055 1645 29090 1650
rect 29055 1605 29090 1610
rect 29115 1645 29150 1650
rect 29115 1605 29150 1610
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1590 4845 1595
rect 5410 1595 5450 1600
rect 5410 1590 5415 1595
rect 4840 1570 5415 1590
rect 4840 1565 4845 1570
rect 4805 1560 4845 1565
rect 5410 1565 5415 1570
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1540 4305 1545
rect 4385 1545 4425 1550
rect 4385 1540 4390 1545
rect 4300 1520 4390 1540
rect 4300 1515 4305 1520
rect 4265 1510 4305 1515
rect 4385 1515 4390 1520
rect 4420 1540 4425 1545
rect 4505 1545 4545 1550
rect 4505 1540 4510 1545
rect 4420 1520 4510 1540
rect 4420 1515 4425 1520
rect 4385 1510 4425 1515
rect 4505 1515 4510 1520
rect 4540 1540 4545 1545
rect 4625 1545 4665 1550
rect 4625 1540 4630 1545
rect 4540 1520 4630 1540
rect 4540 1515 4545 1520
rect 4505 1510 4545 1515
rect 4625 1515 4630 1520
rect 4660 1540 4665 1545
rect 4745 1545 4785 1550
rect 4745 1540 4750 1545
rect 4660 1520 4750 1540
rect 4660 1515 4665 1520
rect 4625 1510 4665 1515
rect 4745 1515 4750 1520
rect 4780 1540 4785 1545
rect 5135 1545 5175 1550
rect 5135 1540 5140 1545
rect 4780 1520 5140 1540
rect 4780 1515 4785 1520
rect 4745 1510 4785 1515
rect 5135 1515 5140 1520
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 2925 1500 2965 1505
rect 2925 1470 2930 1500
rect 2960 1495 2965 1500
rect 3045 1500 3085 1505
rect 3045 1495 3050 1500
rect 2960 1475 3050 1495
rect 2960 1470 2965 1475
rect 2925 1465 2965 1470
rect 3045 1470 3050 1475
rect 3080 1495 3085 1500
rect 3165 1500 3205 1505
rect 3165 1495 3170 1500
rect 3080 1475 3170 1495
rect 3080 1470 3085 1475
rect 3045 1465 3085 1470
rect 3165 1470 3170 1475
rect 3200 1495 3205 1500
rect 3285 1500 3325 1505
rect 3285 1495 3290 1500
rect 3200 1475 3290 1495
rect 3200 1470 3205 1475
rect 3165 1465 3205 1470
rect 3285 1470 3290 1475
rect 3320 1495 3325 1500
rect 3525 1500 3565 1505
rect 3525 1495 3530 1500
rect 3320 1475 3530 1495
rect 3320 1470 3325 1475
rect 3285 1465 3325 1470
rect 3525 1470 3530 1475
rect 3560 1495 3565 1500
rect 3645 1500 3685 1505
rect 3645 1495 3650 1500
rect 3560 1475 3650 1495
rect 3560 1470 3565 1475
rect 3525 1465 3565 1470
rect 3645 1470 3650 1475
rect 3680 1495 3685 1500
rect 3765 1500 3805 1505
rect 3765 1495 3770 1500
rect 3680 1475 3770 1495
rect 3680 1470 3685 1475
rect 3645 1465 3685 1470
rect 3765 1470 3770 1475
rect 3800 1495 3805 1500
rect 4205 1500 4245 1505
rect 4205 1495 4210 1500
rect 3800 1475 4210 1495
rect 3800 1470 3805 1475
rect 3765 1465 3805 1470
rect 4205 1470 4210 1475
rect 4240 1495 4245 1500
rect 4325 1500 4365 1505
rect 4325 1495 4330 1500
rect 4240 1475 4330 1495
rect 4240 1470 4245 1475
rect 4205 1465 4245 1470
rect 4325 1470 4330 1475
rect 4360 1495 4365 1500
rect 4445 1500 4485 1505
rect 4445 1495 4450 1500
rect 4360 1475 4450 1495
rect 4360 1470 4365 1475
rect 4325 1465 4365 1470
rect 4445 1470 4450 1475
rect 4480 1495 4485 1500
rect 4685 1500 4725 1505
rect 4685 1495 4690 1500
rect 4480 1475 4690 1495
rect 4480 1470 4485 1475
rect 4445 1465 4485 1470
rect 4685 1470 4690 1475
rect 4720 1495 4725 1500
rect 4805 1500 4845 1505
rect 4805 1495 4810 1500
rect 4720 1475 4810 1495
rect 4720 1470 4725 1475
rect 4685 1465 4725 1470
rect 4805 1470 4810 1475
rect 4840 1495 4845 1500
rect 4925 1500 4965 1505
rect 4925 1495 4930 1500
rect 4840 1475 4930 1495
rect 4840 1470 4845 1475
rect 4805 1465 4845 1470
rect 4925 1470 4930 1475
rect 4960 1495 4965 1500
rect 5045 1500 5085 1505
rect 5045 1495 5050 1500
rect 4960 1475 5050 1495
rect 4960 1470 4965 1475
rect 4925 1465 4965 1470
rect 5045 1470 5050 1475
rect 5080 1495 5085 1500
rect 5550 1500 5590 1505
rect 5550 1495 5555 1500
rect 5080 1475 5555 1495
rect 5080 1470 5085 1475
rect 5045 1465 5085 1470
rect 5550 1470 5555 1475
rect 5585 1470 5590 1500
rect 16106 1495 16138 1500
rect 16106 1490 16109 1495
rect 15940 1470 16109 1490
rect 5550 1465 5590 1470
rect 16106 1465 16109 1470
rect 16135 1490 16138 1495
rect 16305 1495 16345 1500
rect 16305 1490 16310 1495
rect 16135 1470 16310 1490
rect 16135 1465 16138 1470
rect 16106 1460 16138 1465
rect 16305 1465 16310 1470
rect 16340 1490 16345 1495
rect 16525 1495 16565 1500
rect 16525 1490 16530 1495
rect 16340 1470 16530 1490
rect 16340 1465 16345 1470
rect 16305 1460 16345 1465
rect 16525 1465 16530 1470
rect 16560 1490 16565 1495
rect 16922 1495 16954 1500
rect 16922 1490 16925 1495
rect 16560 1470 16925 1490
rect 16560 1465 16565 1470
rect 16525 1460 16565 1465
rect 16922 1465 16925 1470
rect 16951 1490 16954 1495
rect 17146 1495 17178 1500
rect 17146 1490 17149 1495
rect 16951 1470 17149 1490
rect 16951 1465 16954 1470
rect 16922 1460 16954 1465
rect 17146 1465 17149 1470
rect 17175 1490 17178 1495
rect 17345 1495 17385 1500
rect 17345 1490 17350 1495
rect 17175 1470 17350 1490
rect 17175 1465 17178 1470
rect 17146 1460 17178 1465
rect 17345 1465 17350 1470
rect 17380 1490 17385 1495
rect 17565 1495 17605 1500
rect 17565 1490 17570 1495
rect 17380 1470 17570 1490
rect 17380 1465 17385 1470
rect 17345 1460 17385 1465
rect 17565 1465 17570 1470
rect 17600 1465 17605 1495
rect 26106 1495 26138 1500
rect 26106 1490 26109 1495
rect 25940 1470 26109 1490
rect 17565 1460 17605 1465
rect 26106 1465 26109 1470
rect 26135 1490 26138 1495
rect 26305 1495 26345 1500
rect 26305 1490 26310 1495
rect 26135 1470 26310 1490
rect 26135 1465 26138 1470
rect 26106 1460 26138 1465
rect 26305 1465 26310 1470
rect 26340 1490 26345 1495
rect 26525 1495 26565 1500
rect 26525 1490 26530 1495
rect 26340 1470 26530 1490
rect 26340 1465 26345 1470
rect 26305 1460 26345 1465
rect 26525 1465 26530 1470
rect 26560 1490 26565 1495
rect 26922 1495 26954 1500
rect 26922 1490 26925 1495
rect 26560 1470 26925 1490
rect 26560 1465 26565 1470
rect 26525 1460 26565 1465
rect 26922 1465 26925 1470
rect 26951 1490 26954 1495
rect 27146 1495 27178 1500
rect 27146 1490 27149 1495
rect 26951 1470 27149 1490
rect 26951 1465 26954 1470
rect 26922 1460 26954 1465
rect 27146 1465 27149 1470
rect 27175 1490 27178 1495
rect 27345 1495 27385 1500
rect 27345 1490 27350 1495
rect 27175 1470 27350 1490
rect 27175 1465 27178 1470
rect 27146 1460 27178 1465
rect 27345 1465 27350 1470
rect 27380 1490 27385 1495
rect 27565 1495 27605 1500
rect 27565 1490 27570 1495
rect 27380 1470 27570 1490
rect 27380 1465 27385 1470
rect 27345 1460 27385 1465
rect 27565 1465 27570 1470
rect 27600 1465 27605 1495
rect 27565 1460 27605 1465
rect 16145 1435 16185 1440
rect 16145 1405 16150 1435
rect 16180 1430 16185 1435
rect 16250 1435 16290 1440
rect 16250 1430 16255 1435
rect 16180 1410 16255 1430
rect 16180 1405 16185 1410
rect 16145 1400 16185 1405
rect 16250 1405 16255 1410
rect 16285 1430 16290 1435
rect 16360 1435 16400 1440
rect 16360 1430 16365 1435
rect 16285 1410 16365 1430
rect 16285 1405 16290 1410
rect 16250 1400 16290 1405
rect 16360 1405 16365 1410
rect 16395 1430 16400 1435
rect 16470 1435 16510 1440
rect 16470 1430 16475 1435
rect 16395 1410 16475 1430
rect 16395 1405 16400 1410
rect 16360 1400 16400 1405
rect 16470 1405 16475 1410
rect 16505 1430 16510 1435
rect 16580 1435 16620 1440
rect 16580 1430 16585 1435
rect 16505 1410 16585 1430
rect 16505 1405 16510 1410
rect 16470 1400 16510 1405
rect 16580 1405 16585 1410
rect 16615 1430 16620 1435
rect 17185 1435 17225 1440
rect 17185 1430 17190 1435
rect 16615 1410 17190 1430
rect 16615 1405 16620 1410
rect 16580 1400 16620 1405
rect 17185 1405 17190 1410
rect 17220 1430 17225 1435
rect 17290 1435 17330 1440
rect 17290 1430 17295 1435
rect 17220 1410 17295 1430
rect 17220 1405 17225 1410
rect 17185 1400 17225 1405
rect 17290 1405 17295 1410
rect 17325 1430 17330 1435
rect 17400 1435 17440 1440
rect 17400 1430 17405 1435
rect 17325 1410 17405 1430
rect 17325 1405 17330 1410
rect 17290 1400 17330 1405
rect 17400 1405 17405 1410
rect 17435 1430 17440 1435
rect 17510 1435 17550 1440
rect 17510 1430 17515 1435
rect 17435 1410 17515 1430
rect 17435 1405 17440 1410
rect 17400 1400 17440 1405
rect 17510 1405 17515 1410
rect 17545 1430 17550 1435
rect 17620 1435 17660 1440
rect 17620 1430 17625 1435
rect 17545 1410 17625 1430
rect 17545 1405 17550 1410
rect 17510 1400 17550 1405
rect 17620 1405 17625 1410
rect 17655 1405 17660 1435
rect 17620 1400 17660 1405
rect 26145 1435 26185 1440
rect 26145 1405 26150 1435
rect 26180 1430 26185 1435
rect 26250 1435 26290 1440
rect 26250 1430 26255 1435
rect 26180 1410 26255 1430
rect 26180 1405 26185 1410
rect 26145 1400 26185 1405
rect 26250 1405 26255 1410
rect 26285 1430 26290 1435
rect 26360 1435 26400 1440
rect 26360 1430 26365 1435
rect 26285 1410 26365 1430
rect 26285 1405 26290 1410
rect 26250 1400 26290 1405
rect 26360 1405 26365 1410
rect 26395 1430 26400 1435
rect 26470 1435 26510 1440
rect 26470 1430 26475 1435
rect 26395 1410 26475 1430
rect 26395 1405 26400 1410
rect 26360 1400 26400 1405
rect 26470 1405 26475 1410
rect 26505 1430 26510 1435
rect 26580 1435 26620 1440
rect 26580 1430 26585 1435
rect 26505 1410 26585 1430
rect 26505 1405 26510 1410
rect 26470 1400 26510 1405
rect 26580 1405 26585 1410
rect 26615 1430 26620 1435
rect 27185 1435 27225 1440
rect 27185 1430 27190 1435
rect 26615 1410 27190 1430
rect 26615 1405 26620 1410
rect 26580 1400 26620 1405
rect 27185 1405 27190 1410
rect 27220 1430 27225 1435
rect 27290 1435 27330 1440
rect 27290 1430 27295 1435
rect 27220 1410 27295 1430
rect 27220 1405 27225 1410
rect 27185 1400 27225 1405
rect 27290 1405 27295 1410
rect 27325 1430 27330 1435
rect 27400 1435 27440 1440
rect 27400 1430 27405 1435
rect 27325 1410 27405 1430
rect 27325 1405 27330 1410
rect 27290 1400 27330 1405
rect 27400 1405 27405 1410
rect 27435 1430 27440 1435
rect 27510 1435 27550 1440
rect 27510 1430 27515 1435
rect 27435 1410 27515 1430
rect 27435 1405 27440 1410
rect 27400 1400 27440 1405
rect 27510 1405 27515 1410
rect 27545 1430 27550 1435
rect 27620 1435 27660 1440
rect 27620 1430 27625 1435
rect 27545 1410 27625 1430
rect 27545 1405 27550 1410
rect 27510 1400 27550 1405
rect 27620 1405 27625 1410
rect 27655 1405 27660 1435
rect 27620 1400 27660 1405
rect 15735 1390 15775 1395
rect 15735 1360 15740 1390
rect 15770 1385 15775 1390
rect 18075 1390 18115 1395
rect 18075 1385 18080 1390
rect 15770 1365 18080 1385
rect 15770 1360 15775 1365
rect 15735 1355 15775 1360
rect 18075 1360 18080 1365
rect 18110 1360 18115 1390
rect 18075 1355 18115 1360
rect 25735 1390 25775 1395
rect 25735 1360 25740 1390
rect 25770 1385 25775 1390
rect 28025 1390 28065 1395
rect 28025 1385 28030 1390
rect 25770 1365 28030 1385
rect 25770 1360 25775 1365
rect 25735 1355 25775 1360
rect 28025 1360 28030 1365
rect 28060 1360 28065 1390
rect 28025 1355 28065 1360
rect 16005 1345 16045 1350
rect 16005 1315 16010 1345
rect 16040 1340 16045 1345
rect 16810 1345 16850 1350
rect 16810 1340 16815 1345
rect 16040 1320 16815 1340
rect 16040 1315 16045 1320
rect 16005 1310 16045 1315
rect 16810 1315 16815 1320
rect 16845 1315 16850 1345
rect 16810 1310 16850 1315
rect 16315 1295 16355 1300
rect 16315 1265 16320 1295
rect 16350 1290 16355 1295
rect 16880 1295 16920 1300
rect 16880 1290 16885 1295
rect 16350 1270 16885 1290
rect 16350 1265 16355 1270
rect 16315 1260 16355 1265
rect 16880 1265 16885 1270
rect 16915 1265 16920 1295
rect 16880 1260 16920 1265
rect 17595 1250 17635 1255
rect 16425 1235 16465 1240
rect 16425 1205 16430 1235
rect 16460 1230 16465 1235
rect 16535 1235 16575 1240
rect 16535 1230 16540 1235
rect 16460 1210 16540 1230
rect 16460 1205 16465 1210
rect 16425 1200 16465 1205
rect 16535 1205 16540 1210
rect 16570 1230 16575 1235
rect 16645 1235 16685 1240
rect 16645 1230 16650 1235
rect 16570 1210 16650 1230
rect 16570 1205 16575 1210
rect 16535 1200 16575 1205
rect 16645 1205 16650 1210
rect 16680 1230 16685 1235
rect 16755 1235 16795 1240
rect 16755 1230 16760 1235
rect 16680 1210 16760 1230
rect 16680 1205 16685 1210
rect 16645 1200 16685 1205
rect 16755 1205 16760 1210
rect 16790 1230 16795 1235
rect 16865 1235 16905 1240
rect 16865 1230 16870 1235
rect 16790 1210 16870 1230
rect 16790 1205 16795 1210
rect 16755 1200 16795 1205
rect 16865 1205 16870 1210
rect 16900 1230 16905 1235
rect 16975 1235 17015 1240
rect 16975 1230 16980 1235
rect 16900 1210 16980 1230
rect 16900 1205 16905 1210
rect 16865 1200 16905 1205
rect 16975 1205 16980 1210
rect 17010 1230 17015 1235
rect 17085 1235 17125 1240
rect 17085 1230 17090 1235
rect 17010 1210 17090 1230
rect 17010 1205 17015 1210
rect 16975 1200 17015 1205
rect 17085 1205 17090 1210
rect 17120 1230 17125 1235
rect 17195 1235 17235 1240
rect 17195 1230 17200 1235
rect 17120 1210 17200 1230
rect 17120 1205 17125 1210
rect 17085 1200 17125 1205
rect 17195 1205 17200 1210
rect 17230 1230 17235 1235
rect 17305 1235 17345 1240
rect 17305 1230 17310 1235
rect 17230 1210 17310 1230
rect 17230 1205 17235 1210
rect 17195 1200 17235 1205
rect 17305 1205 17310 1210
rect 17340 1230 17345 1235
rect 17415 1235 17455 1240
rect 17415 1230 17420 1235
rect 17340 1210 17420 1230
rect 17340 1205 17345 1210
rect 17305 1200 17345 1205
rect 17415 1205 17420 1210
rect 17450 1230 17455 1235
rect 17525 1235 17565 1240
rect 17525 1230 17530 1235
rect 17450 1210 17530 1230
rect 17450 1205 17455 1210
rect 17415 1200 17455 1205
rect 17525 1205 17530 1210
rect 17560 1205 17565 1235
rect 17595 1220 17600 1250
rect 17630 1245 17635 1250
rect 17905 1250 17945 1255
rect 17905 1245 17910 1250
rect 17630 1225 17910 1245
rect 17630 1220 17635 1225
rect 17595 1215 17635 1220
rect 17905 1220 17910 1225
rect 17940 1220 17945 1250
rect 17905 1215 17945 1220
rect 26005 1245 26045 1250
rect 26005 1215 26010 1245
rect 26040 1240 26045 1245
rect 26810 1245 26850 1250
rect 26810 1240 26815 1245
rect 26040 1220 26815 1240
rect 26040 1215 26045 1220
rect 26005 1210 26045 1215
rect 26810 1215 26815 1220
rect 26845 1215 26850 1245
rect 26810 1210 26850 1215
rect 17525 1200 17565 1205
rect 26315 1195 26355 1200
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1180 3415 1185
rect 3985 1185 4025 1190
rect 3985 1180 3990 1185
rect 3410 1160 3990 1180
rect 3410 1155 3415 1160
rect 3375 1150 3415 1155
rect 3985 1155 3990 1160
rect 4020 1180 4025 1185
rect 4595 1185 4635 1190
rect 4595 1180 4600 1185
rect 4020 1160 4600 1180
rect 4020 1155 4025 1160
rect 3985 1150 4025 1155
rect 4595 1155 4600 1160
rect 4630 1180 4635 1185
rect 5465 1185 5505 1190
rect 5465 1180 5470 1185
rect 4630 1160 5470 1180
rect 4630 1155 4635 1160
rect 4595 1150 4635 1155
rect 5465 1155 5470 1160
rect 5500 1155 5505 1185
rect 26315 1165 26320 1195
rect 26350 1190 26355 1195
rect 26880 1195 26920 1200
rect 26880 1190 26885 1195
rect 26350 1170 26885 1190
rect 26350 1165 26355 1170
rect 26315 1160 26355 1165
rect 26880 1165 26885 1170
rect 26915 1165 26920 1195
rect 26880 1160 26920 1165
rect 5465 1150 5505 1155
rect 27595 1150 27635 1155
rect 26425 1135 26465 1140
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1120 2985 1125
rect 3025 1125 3065 1130
rect 3025 1120 3030 1125
rect 2980 1100 3030 1120
rect 2980 1095 2985 1100
rect 2945 1090 2985 1095
rect 3025 1095 3030 1100
rect 3060 1120 3065 1125
rect 3105 1125 3145 1130
rect 3105 1120 3110 1125
rect 3060 1100 3110 1120
rect 3060 1095 3065 1100
rect 3025 1090 3065 1095
rect 3105 1095 3110 1100
rect 3140 1120 3145 1125
rect 3185 1125 3225 1130
rect 3185 1120 3190 1125
rect 3140 1100 3190 1120
rect 3140 1095 3145 1100
rect 3105 1090 3145 1095
rect 3185 1095 3190 1100
rect 3220 1120 3225 1125
rect 3265 1125 3305 1130
rect 3265 1120 3270 1125
rect 3220 1100 3270 1120
rect 3220 1095 3225 1100
rect 3185 1090 3225 1095
rect 3265 1095 3270 1100
rect 3300 1120 3305 1125
rect 3345 1125 3385 1130
rect 3345 1120 3350 1125
rect 3300 1100 3350 1120
rect 3300 1095 3305 1100
rect 3265 1090 3305 1095
rect 3345 1095 3350 1100
rect 3380 1120 3385 1125
rect 3425 1125 3465 1130
rect 3425 1120 3430 1125
rect 3380 1100 3430 1120
rect 3380 1095 3385 1100
rect 3345 1090 3385 1095
rect 3425 1095 3430 1100
rect 3460 1120 3465 1125
rect 3505 1125 3545 1130
rect 3505 1120 3510 1125
rect 3460 1100 3510 1120
rect 3460 1095 3465 1100
rect 3425 1090 3465 1095
rect 3505 1095 3510 1100
rect 3540 1120 3545 1125
rect 3585 1125 3625 1130
rect 3585 1120 3590 1125
rect 3540 1100 3590 1120
rect 3540 1095 3545 1100
rect 3505 1090 3545 1095
rect 3585 1095 3590 1100
rect 3620 1120 3625 1125
rect 3665 1125 3705 1130
rect 3665 1120 3670 1125
rect 3620 1100 3670 1120
rect 3620 1095 3625 1100
rect 3585 1090 3625 1095
rect 3665 1095 3670 1100
rect 3700 1120 3705 1125
rect 3745 1125 3785 1130
rect 3745 1120 3750 1125
rect 3700 1100 3750 1120
rect 3700 1095 3705 1100
rect 3665 1090 3705 1095
rect 3745 1095 3750 1100
rect 3780 1120 3785 1125
rect 3825 1125 3865 1130
rect 3825 1120 3830 1125
rect 3780 1100 3830 1120
rect 3780 1095 3785 1100
rect 3745 1090 3785 1095
rect 3825 1095 3830 1100
rect 3860 1120 3865 1125
rect 3905 1125 3945 1130
rect 3905 1120 3910 1125
rect 3860 1100 3910 1120
rect 3860 1095 3865 1100
rect 3825 1090 3865 1095
rect 3905 1095 3910 1100
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1120 4025 1125
rect 4065 1125 4105 1130
rect 4065 1120 4070 1125
rect 4020 1100 4070 1120
rect 4020 1095 4025 1100
rect 3985 1090 4025 1095
rect 4065 1095 4070 1100
rect 4100 1120 4105 1125
rect 4145 1125 4185 1130
rect 4145 1120 4150 1125
rect 4100 1100 4150 1120
rect 4100 1095 4105 1100
rect 4065 1090 4105 1095
rect 4145 1095 4150 1100
rect 4180 1120 4185 1125
rect 4225 1125 4265 1130
rect 4225 1120 4230 1125
rect 4180 1100 4230 1120
rect 4180 1095 4185 1100
rect 4145 1090 4185 1095
rect 4225 1095 4230 1100
rect 4260 1120 4265 1125
rect 4305 1125 4345 1130
rect 4305 1120 4310 1125
rect 4260 1100 4310 1120
rect 4260 1095 4265 1100
rect 4225 1090 4265 1095
rect 4305 1095 4310 1100
rect 4340 1120 4345 1125
rect 4385 1125 4425 1130
rect 4385 1120 4390 1125
rect 4340 1100 4390 1120
rect 4340 1095 4345 1100
rect 4305 1090 4345 1095
rect 4385 1095 4390 1100
rect 4420 1120 4425 1125
rect 4465 1125 4505 1130
rect 4465 1120 4470 1125
rect 4420 1100 4470 1120
rect 4420 1095 4425 1100
rect 4385 1090 4425 1095
rect 4465 1095 4470 1100
rect 4500 1120 4505 1125
rect 4545 1125 4585 1130
rect 4545 1120 4550 1125
rect 4500 1100 4550 1120
rect 4500 1095 4505 1100
rect 4465 1090 4505 1095
rect 4545 1095 4550 1100
rect 4580 1120 4585 1125
rect 4625 1125 4665 1130
rect 4625 1120 4630 1125
rect 4580 1100 4630 1120
rect 4580 1095 4585 1100
rect 4545 1090 4585 1095
rect 4625 1095 4630 1100
rect 4660 1120 4665 1125
rect 4705 1125 4745 1130
rect 4705 1120 4710 1125
rect 4660 1100 4710 1120
rect 4660 1095 4665 1100
rect 4625 1090 4665 1095
rect 4705 1095 4710 1100
rect 4740 1120 4745 1125
rect 4785 1125 4825 1130
rect 4785 1120 4790 1125
rect 4740 1100 4790 1120
rect 4740 1095 4745 1100
rect 4705 1090 4745 1095
rect 4785 1095 4790 1100
rect 4820 1120 4825 1125
rect 4865 1125 4905 1130
rect 4865 1120 4870 1125
rect 4820 1100 4870 1120
rect 4820 1095 4825 1100
rect 4785 1090 4825 1095
rect 4865 1095 4870 1100
rect 4900 1120 4905 1125
rect 4945 1125 4985 1130
rect 4945 1120 4950 1125
rect 4900 1100 4950 1120
rect 4900 1095 4905 1100
rect 4865 1090 4905 1095
rect 4945 1095 4950 1100
rect 4980 1095 4985 1125
rect 26425 1105 26430 1135
rect 26460 1130 26465 1135
rect 26535 1135 26575 1140
rect 26535 1130 26540 1135
rect 26460 1110 26540 1130
rect 26460 1105 26465 1110
rect 26425 1100 26465 1105
rect 26535 1105 26540 1110
rect 26570 1130 26575 1135
rect 26645 1135 26685 1140
rect 26645 1130 26650 1135
rect 26570 1110 26650 1130
rect 26570 1105 26575 1110
rect 26535 1100 26575 1105
rect 26645 1105 26650 1110
rect 26680 1130 26685 1135
rect 26755 1135 26795 1140
rect 26755 1130 26760 1135
rect 26680 1110 26760 1130
rect 26680 1105 26685 1110
rect 26645 1100 26685 1105
rect 26755 1105 26760 1110
rect 26790 1130 26795 1135
rect 26865 1135 26905 1140
rect 26865 1130 26870 1135
rect 26790 1110 26870 1130
rect 26790 1105 26795 1110
rect 26755 1100 26795 1105
rect 26865 1105 26870 1110
rect 26900 1130 26905 1135
rect 26975 1135 27015 1140
rect 26975 1130 26980 1135
rect 26900 1110 26980 1130
rect 26900 1105 26905 1110
rect 26865 1100 26905 1105
rect 26975 1105 26980 1110
rect 27010 1130 27015 1135
rect 27085 1135 27125 1140
rect 27085 1130 27090 1135
rect 27010 1110 27090 1130
rect 27010 1105 27015 1110
rect 26975 1100 27015 1105
rect 27085 1105 27090 1110
rect 27120 1130 27125 1135
rect 27195 1135 27235 1140
rect 27195 1130 27200 1135
rect 27120 1110 27200 1130
rect 27120 1105 27125 1110
rect 27085 1100 27125 1105
rect 27195 1105 27200 1110
rect 27230 1130 27235 1135
rect 27305 1135 27345 1140
rect 27305 1130 27310 1135
rect 27230 1110 27310 1130
rect 27230 1105 27235 1110
rect 27195 1100 27235 1105
rect 27305 1105 27310 1110
rect 27340 1130 27345 1135
rect 27415 1135 27455 1140
rect 27415 1130 27420 1135
rect 27340 1110 27420 1130
rect 27340 1105 27345 1110
rect 27305 1100 27345 1105
rect 27415 1105 27420 1110
rect 27450 1130 27455 1135
rect 27525 1135 27565 1140
rect 27525 1130 27530 1135
rect 27450 1110 27530 1130
rect 27450 1105 27455 1110
rect 27415 1100 27455 1105
rect 27525 1105 27530 1110
rect 27560 1105 27565 1135
rect 27595 1120 27600 1150
rect 27630 1145 27635 1150
rect 27915 1150 27955 1155
rect 27915 1145 27920 1150
rect 27630 1125 27920 1145
rect 27630 1120 27635 1125
rect 27595 1115 27635 1120
rect 27915 1120 27920 1125
rect 27950 1120 27955 1150
rect 27915 1115 27955 1120
rect 27525 1100 27565 1105
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1035 2660 1040
rect 2905 1040 2945 1045
rect 2905 1035 2910 1040
rect 2655 1015 2910 1035
rect 2655 1010 2660 1015
rect 2620 1005 2660 1010
rect 2905 1010 2910 1015
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1035 5150 1040
rect 5465 1040 5505 1045
rect 5465 1035 5470 1040
rect 5145 1015 5470 1035
rect 5145 1010 5150 1015
rect 5110 1005 5150 1010
rect 5465 1010 5470 1015
rect 5500 1010 5505 1040
rect 5465 1005 5505 1010
rect 15205 935 15245 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 925 3035 930
rect 3175 930 3215 935
rect 3175 925 3180 930
rect 3030 905 3180 925
rect 3030 900 3035 905
rect 2995 895 3035 900
rect 3175 900 3180 905
rect 3210 925 3215 930
rect 3355 930 3395 935
rect 3355 925 3360 930
rect 3210 905 3360 925
rect 3210 900 3215 905
rect 3175 895 3215 900
rect 3355 900 3360 905
rect 3390 925 3395 930
rect 3535 930 3575 935
rect 3535 925 3540 930
rect 3390 905 3540 925
rect 3390 900 3395 905
rect 3355 895 3395 900
rect 3535 900 3540 905
rect 3570 925 3575 930
rect 3715 930 3755 935
rect 3715 925 3720 930
rect 3570 905 3720 925
rect 3570 900 3575 905
rect 3535 895 3575 900
rect 3715 900 3720 905
rect 3750 925 3755 930
rect 3895 930 3935 935
rect 3895 925 3900 930
rect 3750 905 3900 925
rect 3750 900 3755 905
rect 3715 895 3755 900
rect 3895 900 3900 905
rect 3930 925 3935 930
rect 4075 930 4115 935
rect 4075 925 4080 930
rect 3930 905 4080 925
rect 3930 900 3935 905
rect 3895 895 3935 900
rect 4075 900 4080 905
rect 4110 925 4115 930
rect 4255 930 4295 935
rect 4255 925 4260 930
rect 4110 905 4260 925
rect 4110 900 4115 905
rect 4075 895 4115 900
rect 4255 900 4260 905
rect 4290 925 4295 930
rect 4435 930 4475 935
rect 4435 925 4440 930
rect 4290 905 4440 925
rect 4290 900 4295 905
rect 4255 895 4295 900
rect 4435 900 4440 905
rect 4470 925 4475 930
rect 4615 930 4655 935
rect 4615 925 4620 930
rect 4470 905 4620 925
rect 4470 900 4475 905
rect 4435 895 4475 900
rect 4615 900 4620 905
rect 4650 925 4655 930
rect 4795 930 4835 935
rect 4795 925 4800 930
rect 4650 905 4800 925
rect 4650 900 4655 905
rect 4615 895 4655 900
rect 4795 900 4800 905
rect 4830 925 4835 930
rect 4975 930 5015 935
rect 4975 925 4980 930
rect 4830 905 4980 925
rect 4830 900 4835 905
rect 4795 895 4835 900
rect 4975 900 4980 905
rect 5010 925 5015 930
rect 5465 930 5505 935
rect 5465 925 5470 930
rect 5010 905 5470 925
rect 5010 900 5015 905
rect 4975 895 5015 900
rect 5465 900 5470 905
rect 5500 900 5505 930
rect 15205 905 15210 935
rect 15240 930 15245 935
rect 15405 935 15445 940
rect 15405 930 15410 935
rect 15240 910 15410 930
rect 15240 905 15245 910
rect 15205 900 15245 905
rect 15405 905 15410 910
rect 15440 905 15445 935
rect 18405 935 18445 940
rect 15405 900 15445 905
rect 16165 915 16205 920
rect 5465 895 5505 900
rect 16165 885 16170 915
rect 16200 910 16205 915
rect 16260 915 16300 920
rect 16260 910 16265 915
rect 16200 890 16265 910
rect 16200 885 16205 890
rect 16165 880 16205 885
rect 16260 885 16265 890
rect 16295 910 16300 915
rect 16370 915 16410 920
rect 16370 910 16375 915
rect 16295 890 16375 910
rect 16295 885 16300 890
rect 16260 880 16300 885
rect 16370 885 16375 890
rect 16405 910 16410 915
rect 16480 915 16520 920
rect 16480 910 16485 915
rect 16405 890 16485 910
rect 16405 885 16410 890
rect 16370 880 16410 885
rect 16480 885 16485 890
rect 16515 910 16520 915
rect 16590 915 16630 920
rect 16590 910 16595 915
rect 16515 890 16595 910
rect 16515 885 16520 890
rect 16480 880 16520 885
rect 16590 885 16595 890
rect 16625 910 16630 915
rect 16700 915 16740 920
rect 16700 910 16705 915
rect 16625 890 16705 910
rect 16625 885 16630 890
rect 16590 880 16630 885
rect 16700 885 16705 890
rect 16735 910 16740 915
rect 16810 915 16850 920
rect 16810 910 16815 915
rect 16735 890 16815 910
rect 16735 885 16740 890
rect 16700 880 16740 885
rect 16810 885 16815 890
rect 16845 910 16850 915
rect 16920 915 16960 920
rect 16920 910 16925 915
rect 16845 890 16925 910
rect 16845 885 16850 890
rect 16810 880 16850 885
rect 16920 885 16925 890
rect 16955 910 16960 915
rect 17030 915 17070 920
rect 17030 910 17035 915
rect 16955 890 17035 910
rect 16955 885 16960 890
rect 16920 880 16960 885
rect 17030 885 17035 890
rect 17065 910 17070 915
rect 17140 915 17180 920
rect 17140 910 17145 915
rect 17065 890 17145 910
rect 17065 885 17070 890
rect 17030 880 17070 885
rect 17140 885 17145 890
rect 17175 910 17180 915
rect 17250 915 17290 920
rect 17250 910 17255 915
rect 17175 890 17255 910
rect 17175 885 17180 890
rect 17140 880 17180 885
rect 17250 885 17255 890
rect 17285 910 17290 915
rect 17360 915 17400 920
rect 17360 910 17365 915
rect 17285 890 17365 910
rect 17285 885 17290 890
rect 17250 880 17290 885
rect 17360 885 17365 890
rect 17395 910 17400 915
rect 17470 915 17510 920
rect 17470 910 17475 915
rect 17395 890 17475 910
rect 17395 885 17400 890
rect 17360 880 17400 885
rect 17470 885 17475 890
rect 17505 910 17510 915
rect 17620 915 17660 920
rect 17620 910 17625 915
rect 17505 890 17625 910
rect 17505 885 17510 890
rect 17470 880 17510 885
rect 17620 885 17625 890
rect 17655 885 17660 915
rect 18405 905 18410 935
rect 18440 930 18445 935
rect 18605 935 18645 940
rect 18605 930 18610 935
rect 18440 910 18610 930
rect 18440 905 18445 910
rect 18405 900 18445 905
rect 18605 905 18610 910
rect 18640 905 18645 935
rect 18605 900 18645 905
rect 25205 935 25245 940
rect 25205 905 25210 935
rect 25240 930 25245 935
rect 25405 935 25445 940
rect 25405 930 25410 935
rect 25240 910 25410 930
rect 25240 905 25245 910
rect 25205 900 25245 905
rect 25405 905 25410 910
rect 25440 905 25445 935
rect 25405 900 25445 905
rect 28405 935 28445 940
rect 28405 905 28410 935
rect 28440 930 28445 935
rect 28605 935 28645 940
rect 28605 930 28610 935
rect 28440 910 28610 930
rect 28440 905 28445 910
rect 28405 900 28445 905
rect 28605 905 28610 910
rect 28640 905 28645 935
rect 28605 900 28645 905
rect 17620 880 17660 885
rect 16935 860 16975 865
rect 16005 855 16045 860
rect 16005 825 16010 855
rect 16040 850 16045 855
rect 16495 855 16535 860
rect 16495 850 16500 855
rect 16040 830 16500 850
rect 16040 825 16045 830
rect 16005 820 16045 825
rect 16495 825 16500 830
rect 16530 825 16535 855
rect 16935 830 16940 860
rect 16970 855 16975 860
rect 17155 860 17195 865
rect 17155 855 17160 860
rect 16970 835 17160 855
rect 16970 830 16975 835
rect 16935 825 16975 830
rect 17155 830 17160 835
rect 17190 855 17195 860
rect 17375 860 17415 865
rect 17375 855 17380 860
rect 17190 835 17380 855
rect 17190 830 17195 835
rect 17155 825 17195 830
rect 17375 830 17380 835
rect 17410 855 17415 860
rect 17960 860 18000 865
rect 17960 855 17965 860
rect 17410 835 17965 855
rect 17410 830 17415 835
rect 17375 825 17415 830
rect 17960 830 17965 835
rect 17995 830 18000 860
rect 17960 825 18000 830
rect 16495 820 16535 825
rect 26195 815 26235 820
rect 15800 800 15840 805
rect 15800 770 15805 800
rect 15835 795 15840 800
rect 16305 800 16345 805
rect 16305 795 16310 800
rect 15835 775 16310 795
rect 15835 770 15840 775
rect 15800 765 15840 770
rect 16305 770 16310 775
rect 16340 795 16345 800
rect 16375 800 16415 805
rect 16375 795 16380 800
rect 16340 775 16380 795
rect 16340 770 16345 775
rect 16305 765 16345 770
rect 16375 770 16380 775
rect 16410 795 16415 800
rect 16445 800 16485 805
rect 16445 795 16450 800
rect 16410 775 16450 795
rect 16410 770 16415 775
rect 16375 765 16415 770
rect 16445 770 16450 775
rect 16480 770 16485 800
rect 16445 765 16485 770
rect 17045 800 17085 805
rect 17045 770 17050 800
rect 17080 795 17085 800
rect 17265 800 17305 805
rect 17265 795 17270 800
rect 17080 775 17270 795
rect 17080 770 17085 775
rect 17045 765 17085 770
rect 17265 770 17270 775
rect 17300 795 17305 800
rect 17485 800 17525 805
rect 17485 795 17490 800
rect 17300 775 17490 795
rect 17300 770 17305 775
rect 17265 765 17305 770
rect 17485 770 17490 775
rect 17520 795 17525 800
rect 17905 800 17945 805
rect 17905 795 17910 800
rect 17520 775 17910 795
rect 17520 770 17525 775
rect 17485 765 17525 770
rect 17905 770 17910 775
rect 17940 770 17945 800
rect 26195 785 26200 815
rect 26230 810 26235 815
rect 26260 815 26300 820
rect 26260 810 26265 815
rect 26230 790 26265 810
rect 26230 785 26235 790
rect 26195 780 26235 785
rect 26260 785 26265 790
rect 26295 810 26300 815
rect 26370 815 26410 820
rect 26370 810 26375 815
rect 26295 790 26375 810
rect 26295 785 26300 790
rect 26260 780 26300 785
rect 26370 785 26375 790
rect 26405 810 26410 815
rect 26480 815 26520 820
rect 26480 810 26485 815
rect 26405 790 26485 810
rect 26405 785 26410 790
rect 26370 780 26410 785
rect 26480 785 26485 790
rect 26515 810 26520 815
rect 26590 815 26630 820
rect 26590 810 26595 815
rect 26515 790 26595 810
rect 26515 785 26520 790
rect 26480 780 26520 785
rect 26590 785 26595 790
rect 26625 810 26630 815
rect 26700 815 26740 820
rect 26700 810 26705 815
rect 26625 790 26705 810
rect 26625 785 26630 790
rect 26590 780 26630 785
rect 26700 785 26705 790
rect 26735 810 26740 815
rect 26810 815 26850 820
rect 26810 810 26815 815
rect 26735 790 26815 810
rect 26735 785 26740 790
rect 26700 780 26740 785
rect 26810 785 26815 790
rect 26845 810 26850 815
rect 26920 815 26960 820
rect 26920 810 26925 815
rect 26845 790 26925 810
rect 26845 785 26850 790
rect 26810 780 26850 785
rect 26920 785 26925 790
rect 26955 810 26960 815
rect 27030 815 27070 820
rect 27030 810 27035 815
rect 26955 790 27035 810
rect 26955 785 26960 790
rect 26920 780 26960 785
rect 27030 785 27035 790
rect 27065 810 27070 815
rect 27140 815 27180 820
rect 27140 810 27145 815
rect 27065 790 27145 810
rect 27065 785 27070 790
rect 27030 780 27070 785
rect 27140 785 27145 790
rect 27175 810 27180 815
rect 27250 815 27290 820
rect 27250 810 27255 815
rect 27175 790 27255 810
rect 27175 785 27180 790
rect 27140 780 27180 785
rect 27250 785 27255 790
rect 27285 810 27290 815
rect 27360 815 27400 820
rect 27360 810 27365 815
rect 27285 790 27365 810
rect 27285 785 27290 790
rect 27250 780 27290 785
rect 27360 785 27365 790
rect 27395 810 27400 815
rect 27470 815 27510 820
rect 27470 810 27475 815
rect 27395 790 27475 810
rect 27395 785 27400 790
rect 27360 780 27400 785
rect 27470 785 27475 790
rect 27505 810 27510 815
rect 27585 815 27625 820
rect 27585 810 27590 815
rect 27505 790 27590 810
rect 27505 785 27510 790
rect 27470 780 27510 785
rect 27585 785 27590 790
rect 27620 785 27625 815
rect 27585 780 27625 785
rect 17905 765 17945 770
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 755 2560 760
rect 3130 760 3170 765
rect 3130 755 3135 760
rect 2555 735 3135 755
rect 2555 730 2560 735
rect 2520 725 2560 730
rect 3130 730 3135 735
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 755 3665 760
rect 3985 760 4025 765
rect 3985 755 3990 760
rect 3660 735 3990 755
rect 3660 730 3665 735
rect 3625 725 3665 730
rect 3985 730 3990 735
rect 4020 755 4025 760
rect 4345 760 4385 765
rect 4345 755 4350 760
rect 4020 735 4350 755
rect 4020 730 4025 735
rect 3985 725 4025 730
rect 4345 730 4350 735
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 755 4565 760
rect 4705 760 4745 765
rect 4705 755 4710 760
rect 4560 735 4710 755
rect 4560 730 4565 735
rect 4525 725 4565 730
rect 4705 730 4710 735
rect 4740 755 4745 760
rect 4885 760 4925 765
rect 4885 755 4890 760
rect 4740 735 4890 755
rect 4740 730 4745 735
rect 4705 725 4745 730
rect 4885 730 4890 735
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 700 3485 705
rect 3805 705 3845 710
rect 3805 700 3810 705
rect 3480 680 3810 700
rect 3480 675 3485 680
rect 3445 670 3485 675
rect 3805 675 3810 680
rect 3840 700 3845 705
rect 4165 705 4205 710
rect 4165 700 4170 705
rect 3840 680 4170 700
rect 3840 675 3845 680
rect 3805 670 3845 675
rect 4165 675 4170 680
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 16990 680 17030 685
rect 16990 650 16995 680
rect 17025 675 17030 680
rect 17100 680 17140 685
rect 17100 675 17105 680
rect 17025 655 17105 675
rect 17025 650 17030 655
rect 16990 645 17030 650
rect 17100 650 17105 655
rect 17135 675 17140 680
rect 17210 680 17250 685
rect 17210 675 17215 680
rect 17135 655 17215 675
rect 17135 650 17140 655
rect 17100 645 17140 650
rect 17210 650 17215 655
rect 17245 675 17250 680
rect 17320 680 17360 685
rect 17320 675 17325 680
rect 17245 655 17325 675
rect 17245 650 17250 655
rect 17210 645 17250 650
rect 17320 650 17325 655
rect 17355 675 17360 680
rect 17430 680 17470 685
rect 17430 675 17435 680
rect 17355 655 17435 675
rect 17355 650 17360 655
rect 17320 645 17360 650
rect 17430 650 17435 655
rect 17465 650 17470 680
rect 26935 660 26975 665
rect 17430 645 17470 650
rect 26005 655 26045 660
rect 26005 625 26010 655
rect 26040 650 26045 655
rect 26505 655 26545 660
rect 26505 650 26510 655
rect 26040 630 26510 650
rect 26040 625 26045 630
rect 26005 620 26045 625
rect 26505 625 26510 630
rect 26540 625 26545 655
rect 26935 630 26940 660
rect 26970 655 26975 660
rect 27155 660 27195 665
rect 27155 655 27160 660
rect 26970 635 27160 655
rect 26970 630 26975 635
rect 26935 625 26975 630
rect 27155 630 27160 635
rect 27190 655 27195 660
rect 27375 660 27415 665
rect 27375 655 27380 660
rect 27190 635 27380 655
rect 27190 630 27195 635
rect 27155 625 27195 630
rect 27375 630 27380 635
rect 27410 655 27415 660
rect 27970 660 28010 665
rect 27970 655 27975 660
rect 27410 635 27975 655
rect 27410 630 27415 635
rect 27375 625 27415 630
rect 27970 630 27975 635
rect 28005 630 28010 660
rect 27970 625 28010 630
rect 26505 620 26545 625
rect 25800 600 25840 605
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect 25800 570 25805 600
rect 25835 595 25840 600
rect 26305 600 26345 605
rect 26305 595 26310 600
rect 25835 575 26310 595
rect 25835 570 25840 575
rect 25800 565 25840 570
rect 26305 570 26310 575
rect 26340 595 26345 600
rect 26375 600 26415 605
rect 26375 595 26380 600
rect 26340 575 26380 595
rect 26340 570 26345 575
rect 26305 565 26345 570
rect 26375 570 26380 575
rect 26410 595 26415 600
rect 26445 600 26485 605
rect 26445 595 26450 600
rect 26410 575 26450 595
rect 26410 570 26415 575
rect 26375 565 26415 570
rect 26445 570 26450 575
rect 26480 570 26485 600
rect 26445 565 26485 570
rect 27045 600 27085 605
rect 27045 570 27050 600
rect 27080 595 27085 600
rect 27265 600 27305 605
rect 27265 595 27270 600
rect 27080 575 27270 595
rect 27080 570 27085 575
rect 27045 565 27085 570
rect 27265 570 27270 575
rect 27300 595 27305 600
rect 27485 600 27525 605
rect 27485 595 27490 600
rect 27300 575 27490 595
rect 27300 570 27305 575
rect 27265 565 27305 570
rect 27485 570 27490 575
rect 27520 595 27525 600
rect 27915 600 27955 605
rect 27915 595 27920 600
rect 27520 575 27920 595
rect 27520 570 27525 575
rect 27485 565 27525 570
rect 27915 570 27920 575
rect 27950 570 27955 600
rect 27915 565 27955 570
rect -195 540 -155 545
rect 26990 480 27030 485
rect 26990 450 26995 480
rect 27025 475 27030 480
rect 27100 480 27140 485
rect 27100 475 27105 480
rect 27025 455 27105 475
rect 27025 450 27030 455
rect 26990 445 27030 450
rect 27100 450 27105 455
rect 27135 475 27140 480
rect 27210 480 27250 485
rect 27210 475 27215 480
rect 27135 455 27215 475
rect 27135 450 27140 455
rect 27100 445 27140 450
rect 27210 450 27215 455
rect 27245 475 27250 480
rect 27320 480 27360 485
rect 27320 475 27325 480
rect 27245 455 27325 475
rect 27245 450 27250 455
rect 27210 445 27250 450
rect 27320 450 27325 455
rect 27355 475 27360 480
rect 27430 480 27470 485
rect 27430 475 27435 480
rect 27355 455 27435 475
rect 27355 450 27360 455
rect 27320 445 27360 450
rect 27430 450 27435 455
rect 27465 450 27470 480
rect 27430 445 27470 450
<< via2 >>
rect -190 4960 -160 4990
rect 5555 4960 5585 4990
rect 14610 3605 14640 3635
rect 29160 3705 29190 3735
rect 19160 3605 19190 3635
rect 24610 3605 24640 3635
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5555 3415 5585 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect -105 2880 -75 2910
rect 5555 2780 5585 2810
rect 5555 2065 5585 2095
rect 14520 2080 14550 2110
rect 19250 2080 19280 2110
rect 24520 2080 24550 2110
rect 29400 2080 29430 2110
rect -105 1690 -75 1720
rect 5555 1470 5585 1500
rect 5470 1155 5500 1185
rect 5470 1010 5500 1040
rect 5470 900 5500 930
rect -190 545 -160 575
<< metal3 >>
rect 12760 5620 12990 5705
rect 13110 5620 13340 5705
rect 13460 5620 13690 5705
rect 12760 5570 13690 5620
rect 12760 5475 12990 5570
rect 13110 5475 13340 5570
rect 13460 5475 13690 5570
rect 13810 5475 14040 5705
rect 14160 5475 14390 5705
rect 14510 5475 14740 5705
rect 14860 5475 15090 5705
rect 15210 5475 15440 5705
rect 15560 5475 15790 5705
rect 15910 5475 16140 5705
rect 16260 5475 16490 5705
rect 16610 5475 16840 5705
rect 16960 5475 17190 5705
rect 17310 5475 17540 5705
rect 17660 5475 17890 5705
rect 18010 5475 18240 5705
rect 18360 5475 18590 5705
rect 18710 5475 18940 5705
rect 19060 5475 19290 5705
rect 19410 5475 19640 5705
rect 19760 5475 19990 5705
rect 20110 5620 20340 5705
rect 20460 5620 20690 5705
rect 20810 5620 21040 5705
rect 20110 5570 21040 5620
rect 20110 5475 20340 5570
rect 20460 5475 20690 5570
rect 20810 5475 21040 5570
rect 13550 5355 13600 5475
rect 13900 5355 13950 5475
rect 14250 5355 14300 5475
rect 14600 5355 14650 5475
rect 14950 5355 15000 5475
rect 15300 5355 15350 5475
rect 15650 5355 15700 5475
rect 16000 5355 16050 5475
rect 16350 5355 16400 5475
rect 16700 5355 16750 5475
rect 17050 5355 17100 5475
rect 17400 5355 17450 5475
rect 17750 5355 17800 5475
rect 18100 5355 18150 5475
rect 18450 5355 18500 5475
rect 18800 5355 18850 5475
rect 19150 5355 19200 5475
rect 19500 5355 19550 5475
rect 19850 5355 19900 5475
rect 20200 5355 20250 5475
rect 12760 5270 12990 5355
rect 13110 5270 13340 5355
rect 13460 5270 13690 5355
rect 13810 5270 14040 5355
rect 14160 5270 14390 5355
rect 14510 5270 14740 5355
rect 14860 5270 15090 5355
rect 15210 5270 15440 5355
rect 15560 5270 15790 5355
rect 15910 5270 16140 5355
rect 16260 5270 16490 5355
rect 16610 5270 16840 5355
rect 12760 5220 16840 5270
rect 12760 5125 12990 5220
rect 13110 5125 13340 5220
rect 13460 5125 13690 5220
rect 13810 5125 14040 5220
rect 14160 5125 14390 5220
rect 14510 5125 14740 5220
rect 14860 5125 15090 5220
rect 15210 5125 15440 5220
rect 15560 5125 15790 5220
rect 15910 5125 16140 5220
rect 16260 5125 16490 5220
rect 16610 5125 16840 5220
rect 16960 5270 17190 5355
rect 17310 5270 17540 5355
rect 17660 5270 17890 5355
rect 18010 5270 18240 5355
rect 18360 5270 18590 5355
rect 18710 5270 18940 5355
rect 19060 5270 19290 5355
rect 19410 5270 19640 5355
rect 19760 5270 19990 5355
rect 20110 5270 20340 5355
rect 20460 5270 20690 5355
rect 20810 5270 21040 5355
rect 16960 5220 21040 5270
rect 16960 5125 17190 5220
rect 17310 5125 17540 5220
rect 17660 5125 17890 5220
rect 18010 5125 18240 5220
rect 18360 5125 18590 5220
rect 18710 5125 18940 5220
rect 19060 5125 19290 5220
rect 19410 5125 19640 5220
rect 19760 5125 19990 5220
rect 20110 5125 20340 5220
rect 20460 5125 20690 5220
rect 20810 5125 21040 5220
rect 13550 5005 13600 5125
rect 14600 5005 14650 5125
rect 14950 5005 15000 5125
rect 15300 5005 15350 5125
rect 15650 5005 15700 5125
rect 16000 5005 16050 5125
rect 16350 5005 16400 5125
rect 16700 5005 16750 5125
rect 17050 5005 17100 5125
rect 17400 5005 17450 5125
rect 17750 5005 17800 5125
rect 18100 5005 18150 5125
rect 18450 5005 18500 5125
rect 18800 5005 18850 5125
rect 19150 5005 19200 5125
rect 20200 5005 20250 5125
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5545 4995 5595 5000
rect 5545 4955 5550 4995
rect 5590 4955 5595 4995
rect 5545 4950 5595 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5460 4910 5510 4915
rect 5460 4870 5465 4910
rect 5505 4870 5510 4910
rect 5460 4865 5510 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 2910 -70 2970
rect -110 2880 -105 2910
rect -75 2880 -70 2910
rect -110 1720 -70 2880
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5465 1185 5505 4865
rect 5465 1155 5470 1185
rect 5500 1155 5505 1185
rect 5465 1040 5505 1155
rect 5465 1010 5470 1040
rect 5500 1010 5505 1040
rect 5465 930 5505 1010
rect 5465 900 5470 930
rect 5500 900 5505 930
rect 5465 665 5505 900
rect 5550 3445 5590 4950
rect 12760 4920 12990 5005
rect 13110 4920 13340 5005
rect 13460 4920 13690 5005
rect 13810 4920 14040 5005
rect 14160 4920 14390 5005
rect 12760 4870 14390 4920
rect 12760 4775 12990 4870
rect 13110 4775 13340 4870
rect 13460 4775 13690 4870
rect 13810 4775 14040 4870
rect 14160 4775 14390 4870
rect 14510 4775 14740 5005
rect 14860 4775 15090 5005
rect 15210 4775 15440 5005
rect 15560 4775 15790 5005
rect 15910 4775 16140 5005
rect 16260 4775 16490 5005
rect 16610 4775 16840 5005
rect 16960 4775 17190 5005
rect 17310 4775 17540 5005
rect 17660 4775 17890 5005
rect 18010 4775 18240 5005
rect 18360 4775 18590 5005
rect 18710 4775 18940 5005
rect 19060 4775 19290 5005
rect 19410 4920 19640 5005
rect 19760 4920 19990 5005
rect 20110 4920 20340 5005
rect 20460 4920 20690 5005
rect 20810 4920 21040 5005
rect 19410 4870 21040 4920
rect 19410 4775 19640 4870
rect 19760 4775 19990 4870
rect 20110 4775 20340 4870
rect 20460 4775 20690 4870
rect 20810 4775 21040 4870
rect 13550 4655 13600 4775
rect 14600 4655 14650 4775
rect 14950 4655 15000 4775
rect 15300 4655 15350 4775
rect 15650 4655 15700 4775
rect 18100 4655 18150 4775
rect 18450 4655 18500 4775
rect 18800 4655 18850 4775
rect 19150 4655 19200 4775
rect 20200 4655 20250 4775
rect 12760 4570 12990 4655
rect 13110 4570 13340 4655
rect 13460 4570 13690 4655
rect 13810 4570 14040 4655
rect 14160 4570 14390 4655
rect 12760 4520 14390 4570
rect 12760 4425 12990 4520
rect 13110 4425 13340 4520
rect 13460 4425 13690 4520
rect 13810 4425 14040 4520
rect 14160 4425 14390 4520
rect 14510 4425 14740 4655
rect 14860 4425 15090 4655
rect 15210 4425 15440 4655
rect 15560 4425 15790 4655
rect 18010 4425 18240 4655
rect 18360 4425 18590 4655
rect 18710 4425 18940 4655
rect 19060 4425 19290 4655
rect 19410 4570 19640 4655
rect 19760 4570 19990 4655
rect 20110 4570 20340 4655
rect 20460 4570 20690 4655
rect 20810 4570 21040 4655
rect 19410 4520 21040 4570
rect 19410 4425 19640 4520
rect 19760 4425 19990 4520
rect 20110 4425 20340 4520
rect 20460 4425 20690 4520
rect 20810 4425 21040 4520
rect 13550 4305 13600 4425
rect 14600 4305 14650 4425
rect 14950 4305 15000 4425
rect 15300 4305 15350 4425
rect 15650 4305 15700 4425
rect 18100 4305 18150 4425
rect 18450 4305 18500 4425
rect 18800 4305 18850 4425
rect 19150 4305 19200 4425
rect 20200 4305 20250 4425
rect 12760 4220 12990 4305
rect 13110 4220 13340 4305
rect 13460 4220 13690 4305
rect 13810 4220 14040 4305
rect 14160 4220 14390 4305
rect 12760 4170 14390 4220
rect 12760 4075 12990 4170
rect 13110 4075 13340 4170
rect 13460 4075 13690 4170
rect 13810 4075 14040 4170
rect 14160 4075 14390 4170
rect 14510 4075 14740 4305
rect 14860 4075 15090 4305
rect 15210 4075 15440 4305
rect 15560 4075 15790 4305
rect 18010 4075 18240 4305
rect 18360 4075 18590 4305
rect 18710 4075 18940 4305
rect 19060 4075 19290 4305
rect 19410 4220 19640 4305
rect 19760 4220 19990 4305
rect 20110 4220 20340 4305
rect 20460 4220 20690 4305
rect 20810 4220 21040 4305
rect 19410 4170 21040 4220
rect 19410 4075 19640 4170
rect 19760 4075 19990 4170
rect 20110 4075 20340 4170
rect 20460 4075 20690 4170
rect 20810 4075 21040 4170
rect 13550 3955 13600 4075
rect 14600 3955 14650 4075
rect 14950 3955 15000 4075
rect 15300 3955 15350 4075
rect 15650 3955 15700 4075
rect 18100 3955 18150 4075
rect 18450 3955 18500 4075
rect 18800 3955 18850 4075
rect 19150 3955 19200 4075
rect 20200 3955 20250 4075
rect 12760 3870 12990 3955
rect 13110 3870 13340 3955
rect 13460 3870 13690 3955
rect 13810 3870 14040 3955
rect 14160 3870 14390 3955
rect 12760 3820 14390 3870
rect 12760 3725 12990 3820
rect 13110 3725 13340 3820
rect 13460 3725 13690 3820
rect 13810 3725 14040 3820
rect 14160 3725 14390 3820
rect 14510 3725 14740 3955
rect 14860 3725 15090 3955
rect 15210 3725 15440 3955
rect 15560 3725 15790 3955
rect 18010 3725 18240 3955
rect 18360 3725 18590 3955
rect 18710 3725 18940 3955
rect 19060 3725 19290 3955
rect 19410 3870 19640 3955
rect 19760 3870 19990 3955
rect 20110 3870 20340 3955
rect 20460 3870 20690 3955
rect 20810 3870 21040 3955
rect 19410 3820 21040 3870
rect 19410 3725 19640 3820
rect 19760 3725 19990 3820
rect 20110 3725 20340 3820
rect 20460 3725 20690 3820
rect 20810 3725 21040 3820
rect 29155 3735 29195 3800
rect 13550 3605 13600 3725
rect 14605 3635 14645 3725
rect 14605 3605 14610 3635
rect 14640 3605 14645 3635
rect 5550 3415 5555 3445
rect 5585 3415 5590 3445
rect 5550 2810 5590 3415
rect 12760 3520 12990 3605
rect 13110 3520 13340 3605
rect 13460 3520 13690 3605
rect 13810 3520 14040 3605
rect 14160 3520 14390 3605
rect 14605 3600 14645 3605
rect 19155 3635 19195 3725
rect 19155 3605 19160 3635
rect 19190 3605 19195 3635
rect 20200 3605 20250 3725
rect 29155 3705 29160 3735
rect 29190 3705 29195 3735
rect 29155 3700 29195 3705
rect 24605 3635 24645 3680
rect 24605 3605 24610 3635
rect 24640 3605 24645 3635
rect 19155 3600 19195 3605
rect 12760 3470 14390 3520
rect 12760 3375 12990 3470
rect 13110 3375 13340 3470
rect 13460 3375 13690 3470
rect 13810 3375 14040 3470
rect 14160 3375 14390 3470
rect 19410 3520 19640 3605
rect 19760 3520 19990 3605
rect 20110 3520 20340 3605
rect 20460 3520 20690 3605
rect 20810 3520 21040 3605
rect 24605 3600 24645 3605
rect 19410 3470 21040 3520
rect 19410 3375 19640 3470
rect 19760 3375 19990 3470
rect 20110 3375 20340 3470
rect 20460 3375 20690 3470
rect 20810 3375 21040 3470
rect 13550 3255 13600 3375
rect 20200 3255 20250 3375
rect 12760 3170 12990 3255
rect 13110 3170 13340 3255
rect 13460 3170 13690 3255
rect 13810 3170 14040 3255
rect 14160 3170 14390 3255
rect 12760 3120 14390 3170
rect 12760 3025 12990 3120
rect 13110 3025 13340 3120
rect 13460 3025 13690 3120
rect 13810 3025 14040 3120
rect 14160 3025 14390 3120
rect 19410 3170 19640 3255
rect 19760 3170 19990 3255
rect 20110 3170 20340 3255
rect 20460 3170 20690 3255
rect 20810 3170 21040 3255
rect 19410 3120 21040 3170
rect 19410 3025 19640 3120
rect 19760 3025 19990 3120
rect 20110 3025 20340 3120
rect 20460 3025 20690 3120
rect 20810 3025 21040 3120
rect 13550 2905 13600 3025
rect 20200 2905 20250 3025
rect 5550 2780 5555 2810
rect 5585 2780 5590 2810
rect 5550 2095 5590 2780
rect 12760 2820 12990 2905
rect 13110 2820 13340 2905
rect 13460 2820 13690 2905
rect 13810 2820 14040 2905
rect 14160 2820 14390 2905
rect 12760 2770 14390 2820
rect 12760 2675 12990 2770
rect 13110 2675 13340 2770
rect 13460 2675 13690 2770
rect 13810 2675 14040 2770
rect 14160 2675 14390 2770
rect 19410 2820 19640 2905
rect 19760 2820 19990 2905
rect 20110 2820 20340 2905
rect 20460 2820 20690 2905
rect 20810 2820 21040 2905
rect 19410 2770 21040 2820
rect 19410 2675 19640 2770
rect 19760 2675 19990 2770
rect 20110 2675 20340 2770
rect 20460 2675 20690 2770
rect 20810 2675 21040 2770
rect 13550 2555 13600 2675
rect 20200 2555 20250 2675
rect 12760 2470 12990 2555
rect 13110 2470 13340 2555
rect 13460 2470 13690 2555
rect 13810 2470 14040 2555
rect 14160 2470 14390 2555
rect 12760 2420 14390 2470
rect 12760 2325 12990 2420
rect 13110 2325 13340 2420
rect 13460 2325 13690 2420
rect 13810 2325 14040 2420
rect 14160 2325 14390 2420
rect 19410 2470 19640 2555
rect 19760 2470 19990 2555
rect 20110 2470 20340 2555
rect 20460 2470 20690 2555
rect 20810 2470 21040 2555
rect 19410 2420 21040 2470
rect 19410 2325 19640 2420
rect 19760 2325 19990 2420
rect 20110 2325 20340 2420
rect 20460 2325 20690 2420
rect 20810 2325 21040 2420
rect 13550 2205 13600 2325
rect 20200 2205 20250 2325
rect 5550 2065 5555 2095
rect 5585 2065 5590 2095
rect 5550 1500 5590 2065
rect 12760 2120 12990 2205
rect 13110 2120 13340 2205
rect 13460 2120 13690 2205
rect 13810 2120 14040 2205
rect 14160 2120 14390 2205
rect 19410 2120 19640 2205
rect 19760 2120 19990 2205
rect 20110 2120 20340 2205
rect 20460 2120 20690 2205
rect 20810 2120 21040 2205
rect 12760 2070 14390 2120
rect 14510 2115 14560 2120
rect 14510 2075 14515 2115
rect 14555 2075 14560 2115
rect 14510 2070 14560 2075
rect 19240 2115 19290 2120
rect 19240 2075 19245 2115
rect 19285 2075 19290 2115
rect 19240 2070 19290 2075
rect 19410 2070 21040 2120
rect 24510 2115 24560 2120
rect 24510 2075 24515 2115
rect 24555 2075 24560 2115
rect 24510 2070 24560 2075
rect 29390 2115 29440 2120
rect 29390 2075 29395 2115
rect 29435 2075 29440 2115
rect 29390 2070 29440 2075
rect 12760 1975 12990 2070
rect 13110 1975 13340 2070
rect 13460 1975 13690 2070
rect 13810 1975 14040 2070
rect 14160 1975 14390 2070
rect 19410 1975 19640 2070
rect 19760 1975 19990 2070
rect 20110 1975 20340 2070
rect 20460 1975 20690 2070
rect 20810 1975 21040 2070
rect 13550 1855 13600 1975
rect 20200 1855 20250 1975
rect 12760 1770 12990 1855
rect 13110 1770 13340 1855
rect 13460 1770 13690 1855
rect 13810 1770 14040 1855
rect 14160 1770 14390 1855
rect 12760 1720 14390 1770
rect 12760 1625 12990 1720
rect 13110 1625 13340 1720
rect 13460 1625 13690 1720
rect 13810 1625 14040 1720
rect 14160 1625 14390 1720
rect 19410 1770 19640 1855
rect 19760 1770 19990 1855
rect 20110 1770 20340 1855
rect 20460 1770 20690 1855
rect 20810 1770 21040 1855
rect 19410 1720 21040 1770
rect 19410 1625 19640 1720
rect 19760 1625 19990 1720
rect 20110 1625 20340 1720
rect 20460 1625 20690 1720
rect 20810 1625 21040 1720
rect 13550 1505 13600 1625
rect 20200 1505 20250 1625
rect 5550 1470 5555 1500
rect 5585 1470 5590 1500
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5460 660 5510 665
rect 5460 620 5465 660
rect 5505 620 5510 660
rect 5460 615 5510 620
rect 5550 585 5590 1470
rect 12760 1420 12990 1505
rect 13110 1420 13340 1505
rect 13460 1420 13690 1505
rect 13810 1420 14040 1505
rect 14160 1420 14390 1505
rect 12760 1370 14390 1420
rect 12760 1275 12990 1370
rect 13110 1275 13340 1370
rect 13460 1275 13690 1370
rect 13810 1275 14040 1370
rect 14160 1275 14390 1370
rect 19410 1420 19640 1505
rect 19760 1420 19990 1505
rect 20110 1420 20340 1505
rect 20460 1420 20690 1505
rect 20810 1420 21040 1505
rect 19410 1370 21040 1420
rect 19410 1275 19640 1370
rect 19760 1275 19990 1370
rect 20110 1275 20340 1370
rect 20460 1275 20690 1370
rect 20810 1275 21040 1370
rect 13550 1155 13600 1275
rect 20200 1155 20250 1275
rect 12760 1070 12990 1155
rect 13110 1070 13340 1155
rect 13460 1070 13690 1155
rect 13810 1070 14040 1155
rect 14160 1070 14390 1155
rect 12760 1020 14390 1070
rect 12760 925 12990 1020
rect 13110 925 13340 1020
rect 13460 925 13690 1020
rect 13810 925 14040 1020
rect 14160 925 14390 1020
rect 19410 1070 19640 1155
rect 19760 1070 19990 1155
rect 20110 1070 20340 1155
rect 20460 1070 20690 1155
rect 20810 1070 21040 1155
rect 19410 1020 21040 1070
rect 19410 925 19640 1020
rect 19760 925 19990 1020
rect 20110 925 20340 1020
rect 20460 925 20690 1020
rect 20810 925 21040 1020
rect 13550 805 13600 925
rect 20200 805 20250 925
rect 12760 720 12990 805
rect 13110 720 13340 805
rect 13460 720 13690 805
rect 13810 720 14040 805
rect 14160 720 14390 805
rect 12760 670 14390 720
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5545 580 5595 585
rect 5545 540 5550 580
rect 5590 540 5595 580
rect 12760 575 12990 670
rect 13110 575 13340 670
rect 13460 575 13690 670
rect 13810 575 14040 670
rect 14160 575 14390 670
rect 19410 720 19640 805
rect 19760 720 19990 805
rect 20110 720 20340 805
rect 20460 720 20690 805
rect 20810 720 21040 805
rect 19410 670 21040 720
rect 19410 575 19640 670
rect 19760 575 19990 670
rect 20110 575 20340 670
rect 20460 575 20690 670
rect 20810 575 21040 670
rect 5545 535 5595 540
rect 13550 455 13600 575
rect 20200 455 20250 575
rect 12760 370 12990 455
rect 13110 370 13340 455
rect 13460 370 13690 455
rect 12760 320 13690 370
rect 12760 225 12990 320
rect 13110 225 13340 320
rect 13460 225 13690 320
rect 13810 225 14040 455
rect 14160 225 14390 455
rect 14510 225 14740 455
rect 14860 225 15090 455
rect 15210 225 15440 455
rect 15560 225 15790 455
rect 15910 225 16140 455
rect 16260 225 16490 455
rect 16610 225 16840 455
rect 16960 225 17190 455
rect 17310 225 17540 455
rect 17660 225 17890 455
rect 18010 225 18240 455
rect 18360 225 18590 455
rect 18710 225 18940 455
rect 19060 225 19290 455
rect 19410 225 19640 455
rect 19760 225 19990 455
rect 20110 370 20340 455
rect 20460 370 20690 455
rect 20810 370 21040 455
rect 20110 320 21040 370
rect 20110 225 20340 320
rect 20460 225 20690 320
rect 20810 225 21040 320
rect 13550 105 13600 225
rect 13900 105 13950 225
rect 14250 105 14300 225
rect 14600 105 14650 225
rect 14950 105 15000 225
rect 15300 105 15350 225
rect 15650 105 15700 225
rect 16000 105 16050 225
rect 16350 105 16400 225
rect 16700 105 16750 225
rect 17050 105 17100 225
rect 17400 105 17450 225
rect 17750 105 17800 225
rect 18100 105 18150 225
rect 18450 105 18500 225
rect 18800 105 18850 225
rect 19150 105 19200 225
rect 19500 105 19550 225
rect 19850 105 19900 225
rect 20200 105 20250 225
rect 12760 20 12990 105
rect 13110 20 13340 105
rect 13460 20 13690 105
rect 13810 20 14040 105
rect 14160 20 14390 105
rect 14510 20 14740 105
rect 14860 20 15090 105
rect 15210 20 15440 105
rect 15560 20 15790 105
rect 15910 20 16140 105
rect 16260 20 16490 105
rect 16610 20 16840 105
rect 12760 -30 16840 20
rect 12760 -125 12990 -30
rect 13110 -125 13340 -30
rect 13460 -125 13690 -30
rect 13810 -125 14040 -30
rect 14160 -125 14390 -30
rect 14510 -125 14740 -30
rect 14860 -125 15090 -30
rect 15210 -125 15440 -30
rect 15560 -125 15790 -30
rect 15910 -125 16140 -30
rect 16260 -125 16490 -30
rect 16610 -125 16840 -30
rect 16960 20 17190 105
rect 17310 20 17540 105
rect 17660 20 17890 105
rect 18010 20 18240 105
rect 18360 20 18590 105
rect 18710 20 18940 105
rect 19060 20 19290 105
rect 19410 20 19640 105
rect 19760 20 19990 105
rect 20110 20 20340 105
rect 20460 20 20690 105
rect 20810 20 21040 105
rect 16960 -30 21040 20
rect 16960 -125 17190 -30
rect 17310 -125 17540 -30
rect 17660 -125 17890 -30
rect 18010 -125 18240 -30
rect 18360 -125 18590 -30
rect 18710 -125 18940 -30
rect 19060 -125 19290 -30
rect 19410 -125 19640 -30
rect 19760 -125 19990 -30
rect 20110 -125 20340 -30
rect 20460 -125 20690 -30
rect 20810 -125 21040 -30
rect 13550 -245 13600 -125
rect 13900 -245 13950 -125
rect 14250 -245 14300 -125
rect 14600 -245 14650 -125
rect 14950 -245 15000 -125
rect 15300 -245 15350 -125
rect 15650 -245 15700 -125
rect 16000 -245 16050 -125
rect 16350 -245 16400 -125
rect 16700 -245 16750 -125
rect 17050 -245 17100 -125
rect 17400 -245 17450 -125
rect 17750 -245 17800 -125
rect 18100 -245 18150 -125
rect 18450 -245 18500 -125
rect 18800 -245 18850 -125
rect 19150 -245 19200 -125
rect 19500 -245 19550 -125
rect 19850 -245 19900 -125
rect 20200 -245 20250 -125
rect 12760 -330 12990 -245
rect 13110 -330 13340 -245
rect 13460 -330 13690 -245
rect 12760 -380 13690 -330
rect 12760 -475 12990 -380
rect 13110 -475 13340 -380
rect 13460 -475 13690 -380
rect 13810 -475 14040 -245
rect 14160 -475 14390 -245
rect 14510 -475 14740 -245
rect 14860 -475 15090 -245
rect 15210 -475 15440 -245
rect 15560 -475 15790 -245
rect 15910 -475 16140 -245
rect 16260 -475 16490 -245
rect 16610 -475 16840 -245
rect 16960 -475 17190 -245
rect 17310 -475 17540 -245
rect 17660 -475 17890 -245
rect 18010 -475 18240 -245
rect 18360 -475 18590 -245
rect 18710 -475 18940 -245
rect 19060 -475 19290 -245
rect 19410 -475 19640 -245
rect 19760 -475 19990 -245
rect 20110 -330 20340 -245
rect 20460 -330 20690 -245
rect 20810 -330 21040 -245
rect 20110 -380 21040 -330
rect 20110 -475 20340 -380
rect 20460 -475 20690 -380
rect 20810 -475 21040 -380
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5555 4960 5585 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 4870 -70 4910
rect 5465 4870 5505 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect 14515 2110 14555 2115
rect 14515 2080 14520 2110
rect 14520 2080 14550 2110
rect 14550 2080 14555 2110
rect 14515 2075 14555 2080
rect 19245 2110 19285 2115
rect 19245 2080 19250 2110
rect 19250 2080 19280 2110
rect 19280 2080 19285 2110
rect 19245 2075 19285 2080
rect 24515 2110 24555 2115
rect 24515 2080 24520 2110
rect 24520 2080 24550 2110
rect 24550 2080 24555 2110
rect 24515 2075 24555 2080
rect 29395 2110 29435 2115
rect 29395 2080 29400 2110
rect 29400 2080 29430 2110
rect 29430 2080 29435 2110
rect 29395 2075 29435 2080
rect -110 620 -70 660
rect 5465 620 5505 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5550 540 5590 580
<< mimcap >>
rect 12775 5615 12975 5690
rect 12775 5575 12855 5615
rect 12895 5575 12975 5615
rect 12775 5490 12975 5575
rect 13125 5615 13325 5690
rect 13125 5575 13205 5615
rect 13245 5575 13325 5615
rect 13125 5490 13325 5575
rect 13475 5615 13675 5690
rect 13475 5575 13555 5615
rect 13595 5575 13675 5615
rect 13475 5490 13675 5575
rect 13825 5615 14025 5690
rect 13825 5575 13905 5615
rect 13945 5575 14025 5615
rect 13825 5490 14025 5575
rect 14175 5615 14375 5690
rect 14175 5575 14255 5615
rect 14295 5575 14375 5615
rect 14175 5490 14375 5575
rect 14525 5615 14725 5690
rect 14525 5575 14605 5615
rect 14645 5575 14725 5615
rect 14525 5490 14725 5575
rect 14875 5615 15075 5690
rect 14875 5575 14955 5615
rect 14995 5575 15075 5615
rect 14875 5490 15075 5575
rect 15225 5615 15425 5690
rect 15225 5575 15305 5615
rect 15345 5575 15425 5615
rect 15225 5490 15425 5575
rect 15575 5615 15775 5690
rect 15575 5575 15655 5615
rect 15695 5575 15775 5615
rect 15575 5490 15775 5575
rect 15925 5615 16125 5690
rect 15925 5575 16005 5615
rect 16045 5575 16125 5615
rect 15925 5490 16125 5575
rect 16275 5615 16475 5690
rect 16275 5575 16355 5615
rect 16395 5575 16475 5615
rect 16275 5490 16475 5575
rect 16625 5615 16825 5690
rect 16625 5575 16705 5615
rect 16745 5575 16825 5615
rect 16625 5490 16825 5575
rect 16975 5615 17175 5690
rect 16975 5575 17055 5615
rect 17095 5575 17175 5615
rect 16975 5490 17175 5575
rect 17325 5615 17525 5690
rect 17325 5575 17405 5615
rect 17445 5575 17525 5615
rect 17325 5490 17525 5575
rect 17675 5615 17875 5690
rect 17675 5575 17755 5615
rect 17795 5575 17875 5615
rect 17675 5490 17875 5575
rect 18025 5615 18225 5690
rect 18025 5575 18105 5615
rect 18145 5575 18225 5615
rect 18025 5490 18225 5575
rect 18375 5615 18575 5690
rect 18375 5575 18455 5615
rect 18495 5575 18575 5615
rect 18375 5490 18575 5575
rect 18725 5615 18925 5690
rect 18725 5575 18805 5615
rect 18845 5575 18925 5615
rect 18725 5490 18925 5575
rect 19075 5615 19275 5690
rect 19075 5575 19155 5615
rect 19195 5575 19275 5615
rect 19075 5490 19275 5575
rect 19425 5615 19625 5690
rect 19425 5575 19505 5615
rect 19545 5575 19625 5615
rect 19425 5490 19625 5575
rect 19775 5615 19975 5690
rect 19775 5575 19855 5615
rect 19895 5575 19975 5615
rect 19775 5490 19975 5575
rect 20125 5615 20325 5690
rect 20125 5575 20205 5615
rect 20245 5575 20325 5615
rect 20125 5490 20325 5575
rect 20475 5615 20675 5690
rect 20475 5575 20555 5615
rect 20595 5575 20675 5615
rect 20475 5490 20675 5575
rect 20825 5615 21025 5690
rect 20825 5575 20905 5615
rect 20945 5575 21025 5615
rect 20825 5490 21025 5575
rect 12775 5265 12975 5340
rect 12775 5225 12855 5265
rect 12895 5225 12975 5265
rect 12775 5140 12975 5225
rect 13125 5265 13325 5340
rect 13125 5225 13205 5265
rect 13245 5225 13325 5265
rect 13125 5140 13325 5225
rect 13475 5265 13675 5340
rect 13475 5225 13555 5265
rect 13595 5225 13675 5265
rect 13475 5140 13675 5225
rect 13825 5265 14025 5340
rect 13825 5225 13905 5265
rect 13945 5225 14025 5265
rect 13825 5140 14025 5225
rect 14175 5265 14375 5340
rect 14175 5225 14255 5265
rect 14295 5225 14375 5265
rect 14175 5140 14375 5225
rect 14525 5265 14725 5340
rect 14525 5225 14605 5265
rect 14645 5225 14725 5265
rect 14525 5140 14725 5225
rect 14875 5265 15075 5340
rect 14875 5225 14955 5265
rect 14995 5225 15075 5265
rect 14875 5140 15075 5225
rect 15225 5265 15425 5340
rect 15225 5225 15305 5265
rect 15345 5225 15425 5265
rect 15225 5140 15425 5225
rect 15575 5265 15775 5340
rect 15575 5225 15655 5265
rect 15695 5225 15775 5265
rect 15575 5140 15775 5225
rect 15925 5265 16125 5340
rect 15925 5225 16005 5265
rect 16045 5225 16125 5265
rect 15925 5140 16125 5225
rect 16275 5265 16475 5340
rect 16275 5225 16355 5265
rect 16395 5225 16475 5265
rect 16275 5140 16475 5225
rect 16625 5265 16825 5340
rect 16625 5225 16705 5265
rect 16745 5225 16825 5265
rect 16625 5140 16825 5225
rect 16975 5265 17175 5340
rect 16975 5225 17055 5265
rect 17095 5225 17175 5265
rect 16975 5140 17175 5225
rect 17325 5265 17525 5340
rect 17325 5225 17405 5265
rect 17445 5225 17525 5265
rect 17325 5140 17525 5225
rect 17675 5265 17875 5340
rect 17675 5225 17755 5265
rect 17795 5225 17875 5265
rect 17675 5140 17875 5225
rect 18025 5265 18225 5340
rect 18025 5225 18105 5265
rect 18145 5225 18225 5265
rect 18025 5140 18225 5225
rect 18375 5265 18575 5340
rect 18375 5225 18455 5265
rect 18495 5225 18575 5265
rect 18375 5140 18575 5225
rect 18725 5265 18925 5340
rect 18725 5225 18805 5265
rect 18845 5225 18925 5265
rect 18725 5140 18925 5225
rect 19075 5265 19275 5340
rect 19075 5225 19155 5265
rect 19195 5225 19275 5265
rect 19075 5140 19275 5225
rect 19425 5265 19625 5340
rect 19425 5225 19505 5265
rect 19545 5225 19625 5265
rect 19425 5140 19625 5225
rect 19775 5265 19975 5340
rect 19775 5225 19855 5265
rect 19895 5225 19975 5265
rect 19775 5140 19975 5225
rect 20125 5265 20325 5340
rect 20125 5225 20205 5265
rect 20245 5225 20325 5265
rect 20125 5140 20325 5225
rect 20475 5265 20675 5340
rect 20475 5225 20555 5265
rect 20595 5225 20675 5265
rect 20475 5140 20675 5225
rect 20825 5265 21025 5340
rect 20825 5225 20905 5265
rect 20945 5225 21025 5265
rect 20825 5140 21025 5225
rect 12775 4915 12975 4990
rect 12775 4875 12855 4915
rect 12895 4875 12975 4915
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 12775 4790 12975 4875
rect 13125 4915 13325 4990
rect 13125 4875 13205 4915
rect 13245 4875 13325 4915
rect 13125 4790 13325 4875
rect 13475 4915 13675 4990
rect 13475 4875 13555 4915
rect 13595 4875 13675 4915
rect 13475 4790 13675 4875
rect 13825 4915 14025 4990
rect 13825 4875 13905 4915
rect 13945 4875 14025 4915
rect 13825 4790 14025 4875
rect 14175 4915 14375 4990
rect 14175 4875 14255 4915
rect 14295 4875 14375 4915
rect 14175 4790 14375 4875
rect 14525 4915 14725 4990
rect 14525 4875 14605 4915
rect 14645 4875 14725 4915
rect 14525 4790 14725 4875
rect 14875 4915 15075 4990
rect 14875 4875 14955 4915
rect 14995 4875 15075 4915
rect 14875 4790 15075 4875
rect 15225 4915 15425 4990
rect 15225 4875 15305 4915
rect 15345 4875 15425 4915
rect 15225 4790 15425 4875
rect 15575 4915 15775 4990
rect 15575 4875 15655 4915
rect 15695 4875 15775 4915
rect 15575 4790 15775 4875
rect 15925 4915 16125 4990
rect 15925 4875 16005 4915
rect 16045 4875 16125 4915
rect 15925 4790 16125 4875
rect 16275 4915 16475 4990
rect 16275 4875 16355 4915
rect 16395 4875 16475 4915
rect 16275 4790 16475 4875
rect 16625 4915 16825 4990
rect 16625 4875 16705 4915
rect 16745 4875 16825 4915
rect 16625 4790 16825 4875
rect 16975 4915 17175 4990
rect 16975 4875 17055 4915
rect 17095 4875 17175 4915
rect 16975 4790 17175 4875
rect 17325 4915 17525 4990
rect 17325 4875 17405 4915
rect 17445 4875 17525 4915
rect 17325 4790 17525 4875
rect 17675 4915 17875 4990
rect 17675 4875 17755 4915
rect 17795 4875 17875 4915
rect 17675 4790 17875 4875
rect 18025 4915 18225 4990
rect 18025 4875 18105 4915
rect 18145 4875 18225 4915
rect 18025 4790 18225 4875
rect 18375 4915 18575 4990
rect 18375 4875 18455 4915
rect 18495 4875 18575 4915
rect 18375 4790 18575 4875
rect 18725 4915 18925 4990
rect 18725 4875 18805 4915
rect 18845 4875 18925 4915
rect 18725 4790 18925 4875
rect 19075 4915 19275 4990
rect 19075 4875 19155 4915
rect 19195 4875 19275 4915
rect 19075 4790 19275 4875
rect 19425 4915 19625 4990
rect 19425 4875 19505 4915
rect 19545 4875 19625 4915
rect 19425 4790 19625 4875
rect 19775 4915 19975 4990
rect 19775 4875 19855 4915
rect 19895 4875 19975 4915
rect 19775 4790 19975 4875
rect 20125 4915 20325 4990
rect 20125 4875 20205 4915
rect 20245 4875 20325 4915
rect 20125 4790 20325 4875
rect 20475 4915 20675 4990
rect 20475 4875 20555 4915
rect 20595 4875 20675 4915
rect 20475 4790 20675 4875
rect 20825 4915 21025 4990
rect 20825 4875 20905 4915
rect 20945 4875 21025 4915
rect 20825 4790 21025 4875
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 12775 4565 12975 4640
rect 12775 4525 12855 4565
rect 12895 4525 12975 4565
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 12775 4440 12975 4525
rect 13125 4565 13325 4640
rect 13125 4525 13205 4565
rect 13245 4525 13325 4565
rect 13125 4440 13325 4525
rect 13475 4565 13675 4640
rect 13475 4525 13555 4565
rect 13595 4525 13675 4565
rect 13475 4440 13675 4525
rect 13825 4565 14025 4640
rect 13825 4525 13905 4565
rect 13945 4525 14025 4565
rect 13825 4440 14025 4525
rect 14175 4565 14375 4640
rect 14175 4525 14255 4565
rect 14295 4525 14375 4565
rect 14175 4440 14375 4525
rect 14525 4565 14725 4640
rect 14525 4525 14605 4565
rect 14645 4525 14725 4565
rect 14525 4440 14725 4525
rect 14875 4565 15075 4640
rect 14875 4525 14955 4565
rect 14995 4525 15075 4565
rect 14875 4440 15075 4525
rect 15225 4565 15425 4640
rect 15225 4525 15305 4565
rect 15345 4525 15425 4565
rect 15225 4440 15425 4525
rect 15575 4565 15775 4640
rect 15575 4525 15655 4565
rect 15695 4525 15775 4565
rect 15575 4440 15775 4525
rect 18025 4565 18225 4640
rect 18025 4525 18105 4565
rect 18145 4525 18225 4565
rect 18025 4440 18225 4525
rect 18375 4565 18575 4640
rect 18375 4525 18455 4565
rect 18495 4525 18575 4565
rect 18375 4440 18575 4525
rect 18725 4565 18925 4640
rect 18725 4525 18805 4565
rect 18845 4525 18925 4565
rect 18725 4440 18925 4525
rect 19075 4565 19275 4640
rect 19075 4525 19155 4565
rect 19195 4525 19275 4565
rect 19075 4440 19275 4525
rect 19425 4565 19625 4640
rect 19425 4525 19505 4565
rect 19545 4525 19625 4565
rect 19425 4440 19625 4525
rect 19775 4565 19975 4640
rect 19775 4525 19855 4565
rect 19895 4525 19975 4565
rect 19775 4440 19975 4525
rect 20125 4565 20325 4640
rect 20125 4525 20205 4565
rect 20245 4525 20325 4565
rect 20125 4440 20325 4525
rect 20475 4565 20675 4640
rect 20475 4525 20555 4565
rect 20595 4525 20675 4565
rect 20475 4440 20675 4525
rect 20825 4565 21025 4640
rect 20825 4525 20905 4565
rect 20945 4525 21025 4565
rect 20825 4440 21025 4525
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 12775 4215 12975 4290
rect 12775 4175 12855 4215
rect 12895 4175 12975 4215
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 12775 4090 12975 4175
rect 13125 4215 13325 4290
rect 13125 4175 13205 4215
rect 13245 4175 13325 4215
rect 13125 4090 13325 4175
rect 13475 4215 13675 4290
rect 13475 4175 13555 4215
rect 13595 4175 13675 4215
rect 13475 4090 13675 4175
rect 13825 4215 14025 4290
rect 13825 4175 13905 4215
rect 13945 4175 14025 4215
rect 13825 4090 14025 4175
rect 14175 4215 14375 4290
rect 14175 4175 14255 4215
rect 14295 4175 14375 4215
rect 14175 4090 14375 4175
rect 14525 4215 14725 4290
rect 14525 4175 14605 4215
rect 14645 4175 14725 4215
rect 14525 4090 14725 4175
rect 14875 4215 15075 4290
rect 14875 4175 14955 4215
rect 14995 4175 15075 4215
rect 14875 4090 15075 4175
rect 15225 4215 15425 4290
rect 15225 4175 15305 4215
rect 15345 4175 15425 4215
rect 15225 4090 15425 4175
rect 15575 4215 15775 4290
rect 15575 4175 15655 4215
rect 15695 4175 15775 4215
rect 15575 4090 15775 4175
rect 18025 4215 18225 4290
rect 18025 4175 18105 4215
rect 18145 4175 18225 4215
rect 18025 4090 18225 4175
rect 18375 4215 18575 4290
rect 18375 4175 18455 4215
rect 18495 4175 18575 4215
rect 18375 4090 18575 4175
rect 18725 4215 18925 4290
rect 18725 4175 18805 4215
rect 18845 4175 18925 4215
rect 18725 4090 18925 4175
rect 19075 4215 19275 4290
rect 19075 4175 19155 4215
rect 19195 4175 19275 4215
rect 19075 4090 19275 4175
rect 19425 4215 19625 4290
rect 19425 4175 19505 4215
rect 19545 4175 19625 4215
rect 19425 4090 19625 4175
rect 19775 4215 19975 4290
rect 19775 4175 19855 4215
rect 19895 4175 19975 4215
rect 19775 4090 19975 4175
rect 20125 4215 20325 4290
rect 20125 4175 20205 4215
rect 20245 4175 20325 4215
rect 20125 4090 20325 4175
rect 20475 4215 20675 4290
rect 20475 4175 20555 4215
rect 20595 4175 20675 4215
rect 20475 4090 20675 4175
rect 20825 4215 21025 4290
rect 20825 4175 20905 4215
rect 20945 4175 21025 4215
rect 20825 4090 21025 4175
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 12775 3865 12975 3940
rect 12775 3825 12855 3865
rect 12895 3825 12975 3865
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 12775 3740 12975 3825
rect 13125 3865 13325 3940
rect 13125 3825 13205 3865
rect 13245 3825 13325 3865
rect 13125 3740 13325 3825
rect 13475 3865 13675 3940
rect 13475 3825 13555 3865
rect 13595 3825 13675 3865
rect 13475 3740 13675 3825
rect 13825 3865 14025 3940
rect 13825 3825 13905 3865
rect 13945 3825 14025 3865
rect 13825 3740 14025 3825
rect 14175 3865 14375 3940
rect 14175 3825 14255 3865
rect 14295 3825 14375 3865
rect 14175 3740 14375 3825
rect 14525 3865 14725 3940
rect 14525 3825 14605 3865
rect 14645 3825 14725 3865
rect 14525 3740 14725 3825
rect 14875 3865 15075 3940
rect 14875 3825 14955 3865
rect 14995 3825 15075 3865
rect 14875 3740 15075 3825
rect 15225 3865 15425 3940
rect 15225 3825 15305 3865
rect 15345 3825 15425 3865
rect 15225 3740 15425 3825
rect 15575 3865 15775 3940
rect 15575 3825 15655 3865
rect 15695 3825 15775 3865
rect 15575 3740 15775 3825
rect 18025 3865 18225 3940
rect 18025 3825 18105 3865
rect 18145 3825 18225 3865
rect 18025 3740 18225 3825
rect 18375 3865 18575 3940
rect 18375 3825 18455 3865
rect 18495 3825 18575 3865
rect 18375 3740 18575 3825
rect 18725 3865 18925 3940
rect 18725 3825 18805 3865
rect 18845 3825 18925 3865
rect 18725 3740 18925 3825
rect 19075 3865 19275 3940
rect 19075 3825 19155 3865
rect 19195 3825 19275 3865
rect 19075 3740 19275 3825
rect 19425 3865 19625 3940
rect 19425 3825 19505 3865
rect 19545 3825 19625 3865
rect 19425 3740 19625 3825
rect 19775 3865 19975 3940
rect 19775 3825 19855 3865
rect 19895 3825 19975 3865
rect 19775 3740 19975 3825
rect 20125 3865 20325 3940
rect 20125 3825 20205 3865
rect 20245 3825 20325 3865
rect 20125 3740 20325 3825
rect 20475 3865 20675 3940
rect 20475 3825 20555 3865
rect 20595 3825 20675 3865
rect 20475 3740 20675 3825
rect 20825 3865 21025 3940
rect 20825 3825 20905 3865
rect 20945 3825 21025 3865
rect 20825 3740 21025 3825
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
rect 12775 3515 12975 3590
rect 12775 3475 12855 3515
rect 12895 3475 12975 3515
rect 12775 3390 12975 3475
rect 13125 3515 13325 3590
rect 13125 3475 13205 3515
rect 13245 3475 13325 3515
rect 13125 3390 13325 3475
rect 13475 3515 13675 3590
rect 13475 3475 13555 3515
rect 13595 3475 13675 3515
rect 13475 3390 13675 3475
rect 13825 3515 14025 3590
rect 13825 3475 13905 3515
rect 13945 3475 14025 3515
rect 13825 3390 14025 3475
rect 14175 3515 14375 3590
rect 14175 3475 14255 3515
rect 14295 3475 14375 3515
rect 14175 3390 14375 3475
rect 19425 3515 19625 3590
rect 19425 3475 19505 3515
rect 19545 3475 19625 3515
rect 19425 3390 19625 3475
rect 19775 3515 19975 3590
rect 19775 3475 19855 3515
rect 19895 3475 19975 3515
rect 19775 3390 19975 3475
rect 20125 3515 20325 3590
rect 20125 3475 20205 3515
rect 20245 3475 20325 3515
rect 20125 3390 20325 3475
rect 20475 3515 20675 3590
rect 20475 3475 20555 3515
rect 20595 3475 20675 3515
rect 20475 3390 20675 3475
rect 20825 3515 21025 3590
rect 20825 3475 20905 3515
rect 20945 3475 21025 3515
rect 20825 3390 21025 3475
rect 12775 3165 12975 3240
rect 12775 3125 12855 3165
rect 12895 3125 12975 3165
rect 12775 3040 12975 3125
rect 13125 3165 13325 3240
rect 13125 3125 13205 3165
rect 13245 3125 13325 3165
rect 13125 3040 13325 3125
rect 13475 3165 13675 3240
rect 13475 3125 13555 3165
rect 13595 3125 13675 3165
rect 13475 3040 13675 3125
rect 13825 3165 14025 3240
rect 13825 3125 13905 3165
rect 13945 3125 14025 3165
rect 13825 3040 14025 3125
rect 14175 3165 14375 3240
rect 14175 3125 14255 3165
rect 14295 3125 14375 3165
rect 14175 3040 14375 3125
rect 19425 3165 19625 3240
rect 19425 3125 19505 3165
rect 19545 3125 19625 3165
rect 19425 3040 19625 3125
rect 19775 3165 19975 3240
rect 19775 3125 19855 3165
rect 19895 3125 19975 3165
rect 19775 3040 19975 3125
rect 20125 3165 20325 3240
rect 20125 3125 20205 3165
rect 20245 3125 20325 3165
rect 20125 3040 20325 3125
rect 20475 3165 20675 3240
rect 20475 3125 20555 3165
rect 20595 3125 20675 3165
rect 20475 3040 20675 3125
rect 20825 3165 21025 3240
rect 20825 3125 20905 3165
rect 20945 3125 21025 3165
rect 20825 3040 21025 3125
rect 12775 2815 12975 2890
rect 12775 2775 12855 2815
rect 12895 2775 12975 2815
rect 12775 2690 12975 2775
rect 13125 2815 13325 2890
rect 13125 2775 13205 2815
rect 13245 2775 13325 2815
rect 13125 2690 13325 2775
rect 13475 2815 13675 2890
rect 13475 2775 13555 2815
rect 13595 2775 13675 2815
rect 13475 2690 13675 2775
rect 13825 2815 14025 2890
rect 13825 2775 13905 2815
rect 13945 2775 14025 2815
rect 13825 2690 14025 2775
rect 14175 2815 14375 2890
rect 14175 2775 14255 2815
rect 14295 2775 14375 2815
rect 14175 2690 14375 2775
rect 19425 2815 19625 2890
rect 19425 2775 19505 2815
rect 19545 2775 19625 2815
rect 19425 2690 19625 2775
rect 19775 2815 19975 2890
rect 19775 2775 19855 2815
rect 19895 2775 19975 2815
rect 19775 2690 19975 2775
rect 20125 2815 20325 2890
rect 20125 2775 20205 2815
rect 20245 2775 20325 2815
rect 20125 2690 20325 2775
rect 20475 2815 20675 2890
rect 20475 2775 20555 2815
rect 20595 2775 20675 2815
rect 20475 2690 20675 2775
rect 20825 2815 21025 2890
rect 20825 2775 20905 2815
rect 20945 2775 21025 2815
rect 20825 2690 21025 2775
rect 12775 2465 12975 2540
rect 12775 2425 12855 2465
rect 12895 2425 12975 2465
rect 12775 2340 12975 2425
rect 13125 2465 13325 2540
rect 13125 2425 13205 2465
rect 13245 2425 13325 2465
rect 13125 2340 13325 2425
rect 13475 2465 13675 2540
rect 13475 2425 13555 2465
rect 13595 2425 13675 2465
rect 13475 2340 13675 2425
rect 13825 2465 14025 2540
rect 13825 2425 13905 2465
rect 13945 2425 14025 2465
rect 13825 2340 14025 2425
rect 14175 2465 14375 2540
rect 14175 2425 14255 2465
rect 14295 2425 14375 2465
rect 14175 2340 14375 2425
rect 19425 2465 19625 2540
rect 19425 2425 19505 2465
rect 19545 2425 19625 2465
rect 19425 2340 19625 2425
rect 19775 2465 19975 2540
rect 19775 2425 19855 2465
rect 19895 2425 19975 2465
rect 19775 2340 19975 2425
rect 20125 2465 20325 2540
rect 20125 2425 20205 2465
rect 20245 2425 20325 2465
rect 20125 2340 20325 2425
rect 20475 2465 20675 2540
rect 20475 2425 20555 2465
rect 20595 2425 20675 2465
rect 20475 2340 20675 2425
rect 20825 2465 21025 2540
rect 20825 2425 20905 2465
rect 20945 2425 21025 2465
rect 20825 2340 21025 2425
rect 12775 2115 12975 2190
rect 12775 2075 12855 2115
rect 12895 2075 12975 2115
rect 12775 1990 12975 2075
rect 13125 2115 13325 2190
rect 13125 2075 13205 2115
rect 13245 2075 13325 2115
rect 13125 1990 13325 2075
rect 13475 2115 13675 2190
rect 13475 2075 13555 2115
rect 13595 2075 13675 2115
rect 13475 1990 13675 2075
rect 13825 2115 14025 2190
rect 13825 2075 13905 2115
rect 13945 2075 14025 2115
rect 13825 1990 14025 2075
rect 14175 2115 14375 2190
rect 14175 2075 14255 2115
rect 14295 2075 14375 2115
rect 14175 1990 14375 2075
rect 19425 2115 19625 2190
rect 19425 2075 19505 2115
rect 19545 2075 19625 2115
rect 19425 1990 19625 2075
rect 19775 2115 19975 2190
rect 19775 2075 19855 2115
rect 19895 2075 19975 2115
rect 19775 1990 19975 2075
rect 20125 2115 20325 2190
rect 20125 2075 20205 2115
rect 20245 2075 20325 2115
rect 20125 1990 20325 2075
rect 20475 2115 20675 2190
rect 20475 2075 20555 2115
rect 20595 2075 20675 2115
rect 20475 1990 20675 2075
rect 20825 2115 21025 2190
rect 20825 2075 20905 2115
rect 20945 2075 21025 2115
rect 20825 1990 21025 2075
rect 12775 1765 12975 1840
rect 12775 1725 12855 1765
rect 12895 1725 12975 1765
rect 12775 1640 12975 1725
rect 13125 1765 13325 1840
rect 13125 1725 13205 1765
rect 13245 1725 13325 1765
rect 13125 1640 13325 1725
rect 13475 1765 13675 1840
rect 13475 1725 13555 1765
rect 13595 1725 13675 1765
rect 13475 1640 13675 1725
rect 13825 1765 14025 1840
rect 13825 1725 13905 1765
rect 13945 1725 14025 1765
rect 13825 1640 14025 1725
rect 14175 1765 14375 1840
rect 14175 1725 14255 1765
rect 14295 1725 14375 1765
rect 14175 1640 14375 1725
rect 19425 1765 19625 1840
rect 19425 1725 19505 1765
rect 19545 1725 19625 1765
rect 19425 1640 19625 1725
rect 19775 1765 19975 1840
rect 19775 1725 19855 1765
rect 19895 1725 19975 1765
rect 19775 1640 19975 1725
rect 20125 1765 20325 1840
rect 20125 1725 20205 1765
rect 20245 1725 20325 1765
rect 20125 1640 20325 1725
rect 20475 1765 20675 1840
rect 20475 1725 20555 1765
rect 20595 1725 20675 1765
rect 20475 1640 20675 1725
rect 20825 1765 21025 1840
rect 20825 1725 20905 1765
rect 20945 1725 21025 1765
rect 20825 1640 21025 1725
rect 12775 1415 12975 1490
rect 12775 1375 12855 1415
rect 12895 1375 12975 1415
rect 12775 1290 12975 1375
rect 13125 1415 13325 1490
rect 13125 1375 13205 1415
rect 13245 1375 13325 1415
rect 13125 1290 13325 1375
rect 13475 1415 13675 1490
rect 13475 1375 13555 1415
rect 13595 1375 13675 1415
rect 13475 1290 13675 1375
rect 13825 1415 14025 1490
rect 13825 1375 13905 1415
rect 13945 1375 14025 1415
rect 13825 1290 14025 1375
rect 14175 1415 14375 1490
rect 14175 1375 14255 1415
rect 14295 1375 14375 1415
rect 14175 1290 14375 1375
rect 19425 1415 19625 1490
rect 19425 1375 19505 1415
rect 19545 1375 19625 1415
rect 19425 1290 19625 1375
rect 19775 1415 19975 1490
rect 19775 1375 19855 1415
rect 19895 1375 19975 1415
rect 19775 1290 19975 1375
rect 20125 1415 20325 1490
rect 20125 1375 20205 1415
rect 20245 1375 20325 1415
rect 20125 1290 20325 1375
rect 20475 1415 20675 1490
rect 20475 1375 20555 1415
rect 20595 1375 20675 1415
rect 20475 1290 20675 1375
rect 20825 1415 21025 1490
rect 20825 1375 20905 1415
rect 20945 1375 21025 1415
rect 20825 1290 21025 1375
rect 12775 1065 12975 1140
rect 12775 1025 12855 1065
rect 12895 1025 12975 1065
rect 12775 940 12975 1025
rect 13125 1065 13325 1140
rect 13125 1025 13205 1065
rect 13245 1025 13325 1065
rect 13125 940 13325 1025
rect 13475 1065 13675 1140
rect 13475 1025 13555 1065
rect 13595 1025 13675 1065
rect 13475 940 13675 1025
rect 13825 1065 14025 1140
rect 13825 1025 13905 1065
rect 13945 1025 14025 1065
rect 13825 940 14025 1025
rect 14175 1065 14375 1140
rect 14175 1025 14255 1065
rect 14295 1025 14375 1065
rect 14175 940 14375 1025
rect 19425 1065 19625 1140
rect 19425 1025 19505 1065
rect 19545 1025 19625 1065
rect 19425 940 19625 1025
rect 19775 1065 19975 1140
rect 19775 1025 19855 1065
rect 19895 1025 19975 1065
rect 19775 940 19975 1025
rect 20125 1065 20325 1140
rect 20125 1025 20205 1065
rect 20245 1025 20325 1065
rect 20125 940 20325 1025
rect 20475 1065 20675 1140
rect 20475 1025 20555 1065
rect 20595 1025 20675 1065
rect 20475 940 20675 1025
rect 20825 1065 21025 1140
rect 20825 1025 20905 1065
rect 20945 1025 21025 1065
rect 20825 940 21025 1025
rect 12775 715 12975 790
rect 12775 675 12855 715
rect 12895 675 12975 715
rect 12775 590 12975 675
rect 13125 715 13325 790
rect 13125 675 13205 715
rect 13245 675 13325 715
rect 13125 590 13325 675
rect 13475 715 13675 790
rect 13475 675 13555 715
rect 13595 675 13675 715
rect 13475 590 13675 675
rect 13825 715 14025 790
rect 13825 675 13905 715
rect 13945 675 14025 715
rect 13825 590 14025 675
rect 14175 715 14375 790
rect 14175 675 14255 715
rect 14295 675 14375 715
rect 14175 590 14375 675
rect 19425 715 19625 790
rect 19425 675 19505 715
rect 19545 675 19625 715
rect 19425 590 19625 675
rect 19775 715 19975 790
rect 19775 675 19855 715
rect 19895 675 19975 715
rect 19775 590 19975 675
rect 20125 715 20325 790
rect 20125 675 20205 715
rect 20245 675 20325 715
rect 20125 590 20325 675
rect 20475 715 20675 790
rect 20475 675 20555 715
rect 20595 675 20675 715
rect 20475 590 20675 675
rect 20825 715 21025 790
rect 20825 675 20905 715
rect 20945 675 21025 715
rect 20825 590 21025 675
rect 12775 365 12975 440
rect 12775 325 12855 365
rect 12895 325 12975 365
rect 12775 240 12975 325
rect 13125 365 13325 440
rect 13125 325 13205 365
rect 13245 325 13325 365
rect 13125 240 13325 325
rect 13475 365 13675 440
rect 13475 325 13555 365
rect 13595 325 13675 365
rect 13475 240 13675 325
rect 13825 365 14025 440
rect 13825 325 13905 365
rect 13945 325 14025 365
rect 13825 240 14025 325
rect 14175 365 14375 440
rect 14175 325 14255 365
rect 14295 325 14375 365
rect 14175 240 14375 325
rect 14525 365 14725 440
rect 14525 325 14605 365
rect 14645 325 14725 365
rect 14525 240 14725 325
rect 14875 365 15075 440
rect 14875 325 14955 365
rect 14995 325 15075 365
rect 14875 240 15075 325
rect 15225 365 15425 440
rect 15225 325 15305 365
rect 15345 325 15425 365
rect 15225 240 15425 325
rect 15575 365 15775 440
rect 15575 325 15655 365
rect 15695 325 15775 365
rect 15575 240 15775 325
rect 15925 365 16125 440
rect 15925 325 16005 365
rect 16045 325 16125 365
rect 15925 240 16125 325
rect 16275 365 16475 440
rect 16275 325 16355 365
rect 16395 325 16475 365
rect 16275 240 16475 325
rect 16625 365 16825 440
rect 16625 325 16705 365
rect 16745 325 16825 365
rect 16625 240 16825 325
rect 16975 365 17175 440
rect 16975 325 17055 365
rect 17095 325 17175 365
rect 16975 240 17175 325
rect 17325 365 17525 440
rect 17325 325 17405 365
rect 17445 325 17525 365
rect 17325 240 17525 325
rect 17675 365 17875 440
rect 17675 325 17755 365
rect 17795 325 17875 365
rect 17675 240 17875 325
rect 18025 365 18225 440
rect 18025 325 18105 365
rect 18145 325 18225 365
rect 18025 240 18225 325
rect 18375 365 18575 440
rect 18375 325 18455 365
rect 18495 325 18575 365
rect 18375 240 18575 325
rect 18725 365 18925 440
rect 18725 325 18805 365
rect 18845 325 18925 365
rect 18725 240 18925 325
rect 19075 365 19275 440
rect 19075 325 19155 365
rect 19195 325 19275 365
rect 19075 240 19275 325
rect 19425 365 19625 440
rect 19425 325 19505 365
rect 19545 325 19625 365
rect 19425 240 19625 325
rect 19775 365 19975 440
rect 19775 325 19855 365
rect 19895 325 19975 365
rect 19775 240 19975 325
rect 20125 365 20325 440
rect 20125 325 20205 365
rect 20245 325 20325 365
rect 20125 240 20325 325
rect 20475 365 20675 440
rect 20475 325 20555 365
rect 20595 325 20675 365
rect 20475 240 20675 325
rect 20825 365 21025 440
rect 20825 325 20905 365
rect 20945 325 21025 365
rect 20825 240 21025 325
rect 12775 15 12975 90
rect 12775 -25 12855 15
rect 12895 -25 12975 15
rect 12775 -110 12975 -25
rect 13125 15 13325 90
rect 13125 -25 13205 15
rect 13245 -25 13325 15
rect 13125 -110 13325 -25
rect 13475 15 13675 90
rect 13475 -25 13555 15
rect 13595 -25 13675 15
rect 13475 -110 13675 -25
rect 13825 15 14025 90
rect 13825 -25 13905 15
rect 13945 -25 14025 15
rect 13825 -110 14025 -25
rect 14175 15 14375 90
rect 14175 -25 14255 15
rect 14295 -25 14375 15
rect 14175 -110 14375 -25
rect 14525 15 14725 90
rect 14525 -25 14605 15
rect 14645 -25 14725 15
rect 14525 -110 14725 -25
rect 14875 15 15075 90
rect 14875 -25 14955 15
rect 14995 -25 15075 15
rect 14875 -110 15075 -25
rect 15225 15 15425 90
rect 15225 -25 15305 15
rect 15345 -25 15425 15
rect 15225 -110 15425 -25
rect 15575 15 15775 90
rect 15575 -25 15655 15
rect 15695 -25 15775 15
rect 15575 -110 15775 -25
rect 15925 15 16125 90
rect 15925 -25 16005 15
rect 16045 -25 16125 15
rect 15925 -110 16125 -25
rect 16275 15 16475 90
rect 16275 -25 16355 15
rect 16395 -25 16475 15
rect 16275 -110 16475 -25
rect 16625 15 16825 90
rect 16625 -25 16705 15
rect 16745 -25 16825 15
rect 16625 -110 16825 -25
rect 16975 15 17175 90
rect 16975 -25 17055 15
rect 17095 -25 17175 15
rect 16975 -110 17175 -25
rect 17325 15 17525 90
rect 17325 -25 17405 15
rect 17445 -25 17525 15
rect 17325 -110 17525 -25
rect 17675 15 17875 90
rect 17675 -25 17755 15
rect 17795 -25 17875 15
rect 17675 -110 17875 -25
rect 18025 15 18225 90
rect 18025 -25 18105 15
rect 18145 -25 18225 15
rect 18025 -110 18225 -25
rect 18375 15 18575 90
rect 18375 -25 18455 15
rect 18495 -25 18575 15
rect 18375 -110 18575 -25
rect 18725 15 18925 90
rect 18725 -25 18805 15
rect 18845 -25 18925 15
rect 18725 -110 18925 -25
rect 19075 15 19275 90
rect 19075 -25 19155 15
rect 19195 -25 19275 15
rect 19075 -110 19275 -25
rect 19425 15 19625 90
rect 19425 -25 19505 15
rect 19545 -25 19625 15
rect 19425 -110 19625 -25
rect 19775 15 19975 90
rect 19775 -25 19855 15
rect 19895 -25 19975 15
rect 19775 -110 19975 -25
rect 20125 15 20325 90
rect 20125 -25 20205 15
rect 20245 -25 20325 15
rect 20125 -110 20325 -25
rect 20475 15 20675 90
rect 20475 -25 20555 15
rect 20595 -25 20675 15
rect 20475 -110 20675 -25
rect 20825 15 21025 90
rect 20825 -25 20905 15
rect 20945 -25 21025 15
rect 20825 -110 21025 -25
rect 12775 -335 12975 -260
rect 12775 -375 12855 -335
rect 12895 -375 12975 -335
rect 12775 -460 12975 -375
rect 13125 -335 13325 -260
rect 13125 -375 13205 -335
rect 13245 -375 13325 -335
rect 13125 -460 13325 -375
rect 13475 -335 13675 -260
rect 13475 -375 13555 -335
rect 13595 -375 13675 -335
rect 13475 -460 13675 -375
rect 13825 -335 14025 -260
rect 13825 -375 13905 -335
rect 13945 -375 14025 -335
rect 13825 -460 14025 -375
rect 14175 -335 14375 -260
rect 14175 -375 14255 -335
rect 14295 -375 14375 -335
rect 14175 -460 14375 -375
rect 14525 -335 14725 -260
rect 14525 -375 14605 -335
rect 14645 -375 14725 -335
rect 14525 -460 14725 -375
rect 14875 -335 15075 -260
rect 14875 -375 14955 -335
rect 14995 -375 15075 -335
rect 14875 -460 15075 -375
rect 15225 -335 15425 -260
rect 15225 -375 15305 -335
rect 15345 -375 15425 -335
rect 15225 -460 15425 -375
rect 15575 -335 15775 -260
rect 15575 -375 15655 -335
rect 15695 -375 15775 -335
rect 15575 -460 15775 -375
rect 15925 -335 16125 -260
rect 15925 -375 16005 -335
rect 16045 -375 16125 -335
rect 15925 -460 16125 -375
rect 16275 -335 16475 -260
rect 16275 -375 16355 -335
rect 16395 -375 16475 -335
rect 16275 -460 16475 -375
rect 16625 -335 16825 -260
rect 16625 -375 16705 -335
rect 16745 -375 16825 -335
rect 16625 -460 16825 -375
rect 16975 -335 17175 -260
rect 16975 -375 17055 -335
rect 17095 -375 17175 -335
rect 16975 -460 17175 -375
rect 17325 -335 17525 -260
rect 17325 -375 17405 -335
rect 17445 -375 17525 -335
rect 17325 -460 17525 -375
rect 17675 -335 17875 -260
rect 17675 -375 17755 -335
rect 17795 -375 17875 -335
rect 17675 -460 17875 -375
rect 18025 -335 18225 -260
rect 18025 -375 18105 -335
rect 18145 -375 18225 -335
rect 18025 -460 18225 -375
rect 18375 -335 18575 -260
rect 18375 -375 18455 -335
rect 18495 -375 18575 -335
rect 18375 -460 18575 -375
rect 18725 -335 18925 -260
rect 18725 -375 18805 -335
rect 18845 -375 18925 -335
rect 18725 -460 18925 -375
rect 19075 -335 19275 -260
rect 19075 -375 19155 -335
rect 19195 -375 19275 -335
rect 19075 -460 19275 -375
rect 19425 -335 19625 -260
rect 19425 -375 19505 -335
rect 19545 -375 19625 -335
rect 19425 -460 19625 -375
rect 19775 -335 19975 -260
rect 19775 -375 19855 -335
rect 19895 -375 19975 -335
rect 19775 -460 19975 -375
rect 20125 -335 20325 -260
rect 20125 -375 20205 -335
rect 20245 -375 20325 -335
rect 20125 -460 20325 -375
rect 20475 -335 20675 -260
rect 20475 -375 20555 -335
rect 20595 -375 20675 -335
rect 20475 -460 20675 -375
rect 20825 -335 21025 -260
rect 20825 -375 20905 -335
rect 20945 -375 21025 -335
rect 20825 -460 21025 -375
<< mimcapcontact >>
rect 12855 5575 12895 5615
rect 13205 5575 13245 5615
rect 13555 5575 13595 5615
rect 13905 5575 13945 5615
rect 14255 5575 14295 5615
rect 14605 5575 14645 5615
rect 14955 5575 14995 5615
rect 15305 5575 15345 5615
rect 15655 5575 15695 5615
rect 16005 5575 16045 5615
rect 16355 5575 16395 5615
rect 16705 5575 16745 5615
rect 17055 5575 17095 5615
rect 17405 5575 17445 5615
rect 17755 5575 17795 5615
rect 18105 5575 18145 5615
rect 18455 5575 18495 5615
rect 18805 5575 18845 5615
rect 19155 5575 19195 5615
rect 19505 5575 19545 5615
rect 19855 5575 19895 5615
rect 20205 5575 20245 5615
rect 20555 5575 20595 5615
rect 20905 5575 20945 5615
rect 12855 5225 12895 5265
rect 13205 5225 13245 5265
rect 13555 5225 13595 5265
rect 13905 5225 13945 5265
rect 14255 5225 14295 5265
rect 14605 5225 14645 5265
rect 14955 5225 14995 5265
rect 15305 5225 15345 5265
rect 15655 5225 15695 5265
rect 16005 5225 16045 5265
rect 16355 5225 16395 5265
rect 16705 5225 16745 5265
rect 17055 5225 17095 5265
rect 17405 5225 17445 5265
rect 17755 5225 17795 5265
rect 18105 5225 18145 5265
rect 18455 5225 18495 5265
rect 18805 5225 18845 5265
rect 19155 5225 19195 5265
rect 19505 5225 19545 5265
rect 19855 5225 19895 5265
rect 20205 5225 20245 5265
rect 20555 5225 20595 5265
rect 20905 5225 20945 5265
rect 12855 4875 12895 4915
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 13205 4875 13245 4915
rect 13555 4875 13595 4915
rect 13905 4875 13945 4915
rect 14255 4875 14295 4915
rect 14605 4875 14645 4915
rect 14955 4875 14995 4915
rect 15305 4875 15345 4915
rect 15655 4875 15695 4915
rect 16005 4875 16045 4915
rect 16355 4875 16395 4915
rect 16705 4875 16745 4915
rect 17055 4875 17095 4915
rect 17405 4875 17445 4915
rect 17755 4875 17795 4915
rect 18105 4875 18145 4915
rect 18455 4875 18495 4915
rect 18805 4875 18845 4915
rect 19155 4875 19195 4915
rect 19505 4875 19545 4915
rect 19855 4875 19895 4915
rect 20205 4875 20245 4915
rect 20555 4875 20595 4915
rect 20905 4875 20945 4915
rect 5140 4725 5180 4765
rect 12855 4525 12895 4565
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 13205 4525 13245 4565
rect 13555 4525 13595 4565
rect 13905 4525 13945 4565
rect 14255 4525 14295 4565
rect 14605 4525 14645 4565
rect 14955 4525 14995 4565
rect 15305 4525 15345 4565
rect 15655 4525 15695 4565
rect 18105 4525 18145 4565
rect 18455 4525 18495 4565
rect 18805 4525 18845 4565
rect 19155 4525 19195 4565
rect 19505 4525 19545 4565
rect 19855 4525 19895 4565
rect 20205 4525 20245 4565
rect 20555 4525 20595 4565
rect 20905 4525 20945 4565
rect 5140 4375 5180 4415
rect 12855 4175 12895 4215
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 13205 4175 13245 4215
rect 13555 4175 13595 4215
rect 13905 4175 13945 4215
rect 14255 4175 14295 4215
rect 14605 4175 14645 4215
rect 14955 4175 14995 4215
rect 15305 4175 15345 4215
rect 15655 4175 15695 4215
rect 18105 4175 18145 4215
rect 18455 4175 18495 4215
rect 18805 4175 18845 4215
rect 19155 4175 19195 4215
rect 19505 4175 19545 4215
rect 19855 4175 19895 4215
rect 20205 4175 20245 4215
rect 20555 4175 20595 4215
rect 20905 4175 20945 4215
rect 5140 4025 5180 4065
rect 12855 3825 12895 3865
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 13205 3825 13245 3865
rect 13555 3825 13595 3865
rect 13905 3825 13945 3865
rect 14255 3825 14295 3865
rect 14605 3825 14645 3865
rect 14955 3825 14995 3865
rect 15305 3825 15345 3865
rect 15655 3825 15695 3865
rect 18105 3825 18145 3865
rect 18455 3825 18495 3865
rect 18805 3825 18845 3865
rect 19155 3825 19195 3865
rect 19505 3825 19545 3865
rect 19855 3825 19895 3865
rect 20205 3825 20245 3865
rect 20555 3825 20595 3865
rect 20905 3825 20945 3865
rect 5140 3675 5180 3715
rect 12855 3475 12895 3515
rect 13205 3475 13245 3515
rect 13555 3475 13595 3515
rect 13905 3475 13945 3515
rect 14255 3475 14295 3515
rect 19505 3475 19545 3515
rect 19855 3475 19895 3515
rect 20205 3475 20245 3515
rect 20555 3475 20595 3515
rect 20905 3475 20945 3515
rect 12855 3125 12895 3165
rect 13205 3125 13245 3165
rect 13555 3125 13595 3165
rect 13905 3125 13945 3165
rect 14255 3125 14295 3165
rect 19505 3125 19545 3165
rect 19855 3125 19895 3165
rect 20205 3125 20245 3165
rect 20555 3125 20595 3165
rect 20905 3125 20945 3165
rect 12855 2775 12895 2815
rect 13205 2775 13245 2815
rect 13555 2775 13595 2815
rect 13905 2775 13945 2815
rect 14255 2775 14295 2815
rect 19505 2775 19545 2815
rect 19855 2775 19895 2815
rect 20205 2775 20245 2815
rect 20555 2775 20595 2815
rect 20905 2775 20945 2815
rect 12855 2425 12895 2465
rect 13205 2425 13245 2465
rect 13555 2425 13595 2465
rect 13905 2425 13945 2465
rect 14255 2425 14295 2465
rect 19505 2425 19545 2465
rect 19855 2425 19895 2465
rect 20205 2425 20245 2465
rect 20555 2425 20595 2465
rect 20905 2425 20945 2465
rect 12855 2075 12895 2115
rect 13205 2075 13245 2115
rect 13555 2075 13595 2115
rect 13905 2075 13945 2115
rect 14255 2075 14295 2115
rect 19505 2075 19545 2115
rect 19855 2075 19895 2115
rect 20205 2075 20245 2115
rect 20555 2075 20595 2115
rect 20905 2075 20945 2115
rect 12855 1725 12895 1765
rect 13205 1725 13245 1765
rect 13555 1725 13595 1765
rect 13905 1725 13945 1765
rect 14255 1725 14295 1765
rect 19505 1725 19545 1765
rect 19855 1725 19895 1765
rect 20205 1725 20245 1765
rect 20555 1725 20595 1765
rect 20905 1725 20945 1765
rect 12855 1375 12895 1415
rect 13205 1375 13245 1415
rect 13555 1375 13595 1415
rect 13905 1375 13945 1415
rect 14255 1375 14295 1415
rect 19505 1375 19545 1415
rect 19855 1375 19895 1415
rect 20205 1375 20245 1415
rect 20555 1375 20595 1415
rect 20905 1375 20945 1415
rect 12855 1025 12895 1065
rect 13205 1025 13245 1065
rect 13555 1025 13595 1065
rect 13905 1025 13945 1065
rect 14255 1025 14295 1065
rect 19505 1025 19545 1065
rect 19855 1025 19895 1065
rect 20205 1025 20245 1065
rect 20555 1025 20595 1065
rect 20905 1025 20945 1065
rect 12855 675 12895 715
rect 13205 675 13245 715
rect 13555 675 13595 715
rect 13905 675 13945 715
rect 14255 675 14295 715
rect 19505 675 19545 715
rect 19855 675 19895 715
rect 20205 675 20245 715
rect 20555 675 20595 715
rect 20905 675 20945 715
rect 12855 325 12895 365
rect 13205 325 13245 365
rect 13555 325 13595 365
rect 13905 325 13945 365
rect 14255 325 14295 365
rect 14605 325 14645 365
rect 14955 325 14995 365
rect 15305 325 15345 365
rect 15655 325 15695 365
rect 16005 325 16045 365
rect 16355 325 16395 365
rect 16705 325 16745 365
rect 17055 325 17095 365
rect 17405 325 17445 365
rect 17755 325 17795 365
rect 18105 325 18145 365
rect 18455 325 18495 365
rect 18805 325 18845 365
rect 19155 325 19195 365
rect 19505 325 19545 365
rect 19855 325 19895 365
rect 20205 325 20245 365
rect 20555 325 20595 365
rect 20905 325 20945 365
rect 12855 -25 12895 15
rect 13205 -25 13245 15
rect 13555 -25 13595 15
rect 13905 -25 13945 15
rect 14255 -25 14295 15
rect 14605 -25 14645 15
rect 14955 -25 14995 15
rect 15305 -25 15345 15
rect 15655 -25 15695 15
rect 16005 -25 16045 15
rect 16355 -25 16395 15
rect 16705 -25 16745 15
rect 17055 -25 17095 15
rect 17405 -25 17445 15
rect 17755 -25 17795 15
rect 18105 -25 18145 15
rect 18455 -25 18495 15
rect 18805 -25 18845 15
rect 19155 -25 19195 15
rect 19505 -25 19545 15
rect 19855 -25 19895 15
rect 20205 -25 20245 15
rect 20555 -25 20595 15
rect 20905 -25 20945 15
rect 12855 -375 12895 -335
rect 13205 -375 13245 -335
rect 13555 -375 13595 -335
rect 13905 -375 13945 -335
rect 14255 -375 14295 -335
rect 14605 -375 14645 -335
rect 14955 -375 14995 -335
rect 15305 -375 15345 -335
rect 15655 -375 15695 -335
rect 16005 -375 16045 -335
rect 16355 -375 16395 -335
rect 16705 -375 16745 -335
rect 17055 -375 17095 -335
rect 17405 -375 17445 -335
rect 17755 -375 17795 -335
rect 18105 -375 18145 -335
rect 18455 -375 18495 -335
rect 18805 -375 18845 -335
rect 19155 -375 19195 -335
rect 19505 -375 19545 -335
rect 19855 -375 19895 -335
rect 20205 -375 20245 -335
rect 20555 -375 20595 -335
rect 20905 -375 20945 -335
<< metal4 >>
rect 12850 5615 13600 5620
rect 12850 5575 12855 5615
rect 12895 5575 13205 5615
rect 13245 5575 13555 5615
rect 13595 5575 13600 5615
rect 12850 5570 13600 5575
rect 13550 5270 13600 5570
rect 13900 5615 13950 5620
rect 13900 5575 13905 5615
rect 13945 5575 13950 5615
rect 13900 5270 13950 5575
rect 14250 5615 14300 5620
rect 14250 5575 14255 5615
rect 14295 5575 14300 5615
rect 14250 5270 14300 5575
rect 14600 5615 14650 5620
rect 14600 5575 14605 5615
rect 14645 5575 14650 5615
rect 14600 5270 14650 5575
rect 14950 5615 15000 5620
rect 14950 5575 14955 5615
rect 14995 5575 15000 5615
rect 14950 5270 15000 5575
rect 15300 5615 15350 5620
rect 15300 5575 15305 5615
rect 15345 5575 15350 5615
rect 15300 5270 15350 5575
rect 15650 5615 15700 5620
rect 15650 5575 15655 5615
rect 15695 5575 15700 5615
rect 15650 5270 15700 5575
rect 16000 5615 16050 5620
rect 16000 5575 16005 5615
rect 16045 5575 16050 5615
rect 16000 5270 16050 5575
rect 16350 5615 16400 5620
rect 16350 5575 16355 5615
rect 16395 5575 16400 5615
rect 16350 5270 16400 5575
rect 16700 5615 16750 5620
rect 16700 5575 16705 5615
rect 16745 5575 16750 5615
rect 16700 5270 16750 5575
rect 12850 5265 16750 5270
rect 12850 5225 12855 5265
rect 12895 5225 13205 5265
rect 13245 5225 13555 5265
rect 13595 5225 13905 5265
rect 13945 5225 14255 5265
rect 14295 5225 14605 5265
rect 14645 5225 14955 5265
rect 14995 5225 15305 5265
rect 15345 5225 15655 5265
rect 15695 5225 16005 5265
rect 16045 5225 16355 5265
rect 16395 5225 16705 5265
rect 16745 5225 16750 5265
rect 12850 5220 16750 5225
rect -200 4995 5595 5000
rect -200 4955 -195 4995
rect -155 4955 5550 4995
rect 5590 4955 5595 4995
rect -200 4950 5595 4955
rect 13550 4920 13600 5220
rect 12850 4915 14300 4920
rect -115 4910 5510 4915
rect -115 4870 -110 4910
rect -70 4870 5465 4910
rect 5505 4870 5510 4910
rect 12850 4875 12855 4915
rect 12895 4875 13205 4915
rect 13245 4875 13555 4915
rect 13595 4875 13905 4915
rect 13945 4875 14255 4915
rect 14295 4875 14300 4915
rect 12850 4870 14300 4875
rect 14600 4915 14650 5220
rect 14600 4875 14605 4915
rect 14645 4875 14650 4915
rect -115 4865 5510 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 13550 4570 13600 4870
rect 12850 4565 14300 4570
rect 12850 4525 12855 4565
rect 12895 4525 13205 4565
rect 13245 4525 13555 4565
rect 13595 4525 13905 4565
rect 13945 4525 14255 4565
rect 14295 4525 14300 4565
rect 12850 4520 14300 4525
rect 14600 4565 14650 4875
rect 14600 4525 14605 4565
rect 14645 4525 14650 4565
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 13550 4220 13600 4520
rect 12850 4215 14300 4220
rect 12850 4175 12855 4215
rect 12895 4175 13205 4215
rect 13245 4175 13555 4215
rect 13595 4175 13905 4215
rect 13945 4175 14255 4215
rect 14295 4175 14300 4215
rect 12850 4170 14300 4175
rect 14600 4215 14650 4525
rect 14600 4175 14605 4215
rect 14645 4175 14650 4215
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 13550 3870 13600 4170
rect 12850 3865 14300 3870
rect 12850 3825 12855 3865
rect 12895 3825 13205 3865
rect 13245 3825 13555 3865
rect 13595 3825 13905 3865
rect 13945 3825 14255 3865
rect 14295 3825 14300 3865
rect 12850 3820 14300 3825
rect 14600 3865 14650 4175
rect 14600 3825 14605 3865
rect 14645 3825 14650 3865
rect 14600 3820 14650 3825
rect 14950 4915 15000 5220
rect 14950 4875 14955 4915
rect 14995 4875 15000 4915
rect 14950 4565 15000 4875
rect 14950 4525 14955 4565
rect 14995 4525 15000 4565
rect 14950 4215 15000 4525
rect 14950 4175 14955 4215
rect 14995 4175 15000 4215
rect 14950 3865 15000 4175
rect 14950 3825 14955 3865
rect 14995 3825 15000 3865
rect 14950 3820 15000 3825
rect 15300 4915 15350 5220
rect 15300 4875 15305 4915
rect 15345 4875 15350 4915
rect 15300 4565 15350 4875
rect 15300 4525 15305 4565
rect 15345 4525 15350 4565
rect 15300 4215 15350 4525
rect 15300 4175 15305 4215
rect 15345 4175 15350 4215
rect 15300 3865 15350 4175
rect 15300 3825 15305 3865
rect 15345 3825 15350 3865
rect 15300 3820 15350 3825
rect 15650 4915 15700 5220
rect 15650 4875 15655 4915
rect 15695 4875 15700 4915
rect 15650 4565 15700 4875
rect 16000 4915 16050 5220
rect 16000 4875 16005 4915
rect 16045 4875 16050 4915
rect 16000 4870 16050 4875
rect 16350 4915 16400 5220
rect 16350 4875 16355 4915
rect 16395 4875 16400 4915
rect 16350 4870 16400 4875
rect 16700 4915 16750 5220
rect 16700 4875 16705 4915
rect 16745 4875 16750 4915
rect 16700 4870 16750 4875
rect 17050 5615 17100 5620
rect 17050 5575 17055 5615
rect 17095 5575 17100 5615
rect 17050 5270 17100 5575
rect 17400 5615 17450 5620
rect 17400 5575 17405 5615
rect 17445 5575 17450 5615
rect 17400 5270 17450 5575
rect 17750 5615 17800 5620
rect 17750 5575 17755 5615
rect 17795 5575 17800 5615
rect 17750 5270 17800 5575
rect 18100 5615 18150 5620
rect 18100 5575 18105 5615
rect 18145 5575 18150 5615
rect 18100 5270 18150 5575
rect 18450 5615 18500 5620
rect 18450 5575 18455 5615
rect 18495 5575 18500 5615
rect 18450 5270 18500 5575
rect 18800 5615 18850 5620
rect 18800 5575 18805 5615
rect 18845 5575 18850 5615
rect 18800 5270 18850 5575
rect 19150 5615 19200 5620
rect 19150 5575 19155 5615
rect 19195 5575 19200 5615
rect 19150 5270 19200 5575
rect 19500 5615 19550 5620
rect 19500 5575 19505 5615
rect 19545 5575 19550 5615
rect 19500 5270 19550 5575
rect 19850 5615 19900 5620
rect 19850 5575 19855 5615
rect 19895 5575 19900 5615
rect 19850 5270 19900 5575
rect 20200 5615 20950 5620
rect 20200 5575 20205 5615
rect 20245 5575 20555 5615
rect 20595 5575 20905 5615
rect 20945 5575 20950 5615
rect 20200 5570 20950 5575
rect 20200 5270 20250 5570
rect 17050 5265 20950 5270
rect 17050 5225 17055 5265
rect 17095 5225 17405 5265
rect 17445 5225 17755 5265
rect 17795 5225 18105 5265
rect 18145 5225 18455 5265
rect 18495 5225 18805 5265
rect 18845 5225 19155 5265
rect 19195 5225 19505 5265
rect 19545 5225 19855 5265
rect 19895 5225 20205 5265
rect 20245 5225 20555 5265
rect 20595 5225 20905 5265
rect 20945 5225 20950 5265
rect 17050 5220 20950 5225
rect 17050 4915 17100 5220
rect 17050 4875 17055 4915
rect 17095 4875 17100 4915
rect 17050 4870 17100 4875
rect 17400 4915 17450 5220
rect 17400 4875 17405 4915
rect 17445 4875 17450 4915
rect 17400 4870 17450 4875
rect 17750 4915 17800 5220
rect 17750 4875 17755 4915
rect 17795 4875 17800 4915
rect 17750 4870 17800 4875
rect 18100 4915 18150 5220
rect 18100 4875 18105 4915
rect 18145 4875 18150 4915
rect 15650 4525 15655 4565
rect 15695 4525 15700 4565
rect 15650 4215 15700 4525
rect 15650 4175 15655 4215
rect 15695 4175 15700 4215
rect 15650 3865 15700 4175
rect 15650 3825 15655 3865
rect 15695 3825 15700 3865
rect 15650 3820 15700 3825
rect 18100 4565 18150 4875
rect 18100 4525 18105 4565
rect 18145 4525 18150 4565
rect 18100 4215 18150 4525
rect 18100 4175 18105 4215
rect 18145 4175 18150 4215
rect 18100 3865 18150 4175
rect 18100 3825 18105 3865
rect 18145 3825 18150 3865
rect 18100 3820 18150 3825
rect 18450 4915 18500 5220
rect 18450 4875 18455 4915
rect 18495 4875 18500 4915
rect 18450 4565 18500 4875
rect 18450 4525 18455 4565
rect 18495 4525 18500 4565
rect 18450 4215 18500 4525
rect 18450 4175 18455 4215
rect 18495 4175 18500 4215
rect 18450 3865 18500 4175
rect 18450 3825 18455 3865
rect 18495 3825 18500 3865
rect 18450 3820 18500 3825
rect 18800 4915 18850 5220
rect 18800 4875 18805 4915
rect 18845 4875 18850 4915
rect 18800 4565 18850 4875
rect 18800 4525 18805 4565
rect 18845 4525 18850 4565
rect 18800 4215 18850 4525
rect 18800 4175 18805 4215
rect 18845 4175 18850 4215
rect 18800 3865 18850 4175
rect 18800 3825 18805 3865
rect 18845 3825 18850 3865
rect 18800 3820 18850 3825
rect 19150 4915 19200 5220
rect 20200 4920 20250 5220
rect 19150 4875 19155 4915
rect 19195 4875 19200 4915
rect 19150 4565 19200 4875
rect 19500 4915 20950 4920
rect 19500 4875 19505 4915
rect 19545 4875 19855 4915
rect 19895 4875 20205 4915
rect 20245 4875 20555 4915
rect 20595 4875 20905 4915
rect 20945 4875 20950 4915
rect 19500 4870 20950 4875
rect 20200 4570 20250 4870
rect 19150 4525 19155 4565
rect 19195 4525 19200 4565
rect 19150 4215 19200 4525
rect 19500 4565 20950 4570
rect 19500 4525 19505 4565
rect 19545 4525 19855 4565
rect 19895 4525 20205 4565
rect 20245 4525 20555 4565
rect 20595 4525 20905 4565
rect 20945 4525 20950 4565
rect 19500 4520 20950 4525
rect 20200 4220 20250 4520
rect 19150 4175 19155 4215
rect 19195 4175 19200 4215
rect 19150 3865 19200 4175
rect 19500 4215 20950 4220
rect 19500 4175 19505 4215
rect 19545 4175 19855 4215
rect 19895 4175 20205 4215
rect 20245 4175 20555 4215
rect 20595 4175 20905 4215
rect 20945 4175 20950 4215
rect 19500 4170 20950 4175
rect 20200 3870 20250 4170
rect 19150 3825 19155 3865
rect 19195 3825 19200 3865
rect 19150 3820 19200 3825
rect 19500 3865 20950 3870
rect 19500 3825 19505 3865
rect 19545 3825 19855 3865
rect 19895 3825 20205 3865
rect 20245 3825 20555 3865
rect 20595 3825 20905 3865
rect 20945 3825 20950 3865
rect 19500 3820 20950 3825
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 13550 3520 13600 3820
rect 20200 3520 20250 3820
rect 12850 3515 14300 3520
rect 12850 3475 12855 3515
rect 12895 3475 13205 3515
rect 13245 3475 13555 3515
rect 13595 3475 13905 3515
rect 13945 3475 14255 3515
rect 14295 3475 14300 3515
rect 12850 3470 14300 3475
rect 19500 3515 20950 3520
rect 19500 3475 19505 3515
rect 19545 3475 19855 3515
rect 19895 3475 20205 3515
rect 20245 3475 20555 3515
rect 20595 3475 20905 3515
rect 20945 3475 20950 3515
rect 19500 3470 20950 3475
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect 13550 3170 13600 3470
rect 20200 3170 20250 3470
rect 12850 3165 14300 3170
rect 12850 3125 12855 3165
rect 12895 3125 13205 3165
rect 13245 3125 13555 3165
rect 13595 3125 13905 3165
rect 13945 3125 14255 3165
rect 14295 3125 14300 3165
rect 12850 3120 14300 3125
rect 19500 3165 20950 3170
rect 19500 3125 19505 3165
rect 19545 3125 19855 3165
rect 19895 3125 20205 3165
rect 20245 3125 20555 3165
rect 20595 3125 20905 3165
rect 20945 3125 20950 3165
rect 19500 3120 20950 3125
rect 13550 2820 13600 3120
rect 20200 2820 20250 3120
rect 12850 2815 14300 2820
rect 12850 2775 12855 2815
rect 12895 2775 13205 2815
rect 13245 2775 13555 2815
rect 13595 2775 13905 2815
rect 13945 2775 14255 2815
rect 14295 2775 14300 2815
rect 12850 2770 14300 2775
rect 19500 2815 20950 2820
rect 19500 2775 19505 2815
rect 19545 2775 19855 2815
rect 19895 2775 20205 2815
rect 20245 2775 20555 2815
rect 20595 2775 20905 2815
rect 20945 2775 20950 2815
rect 19500 2770 20950 2775
rect 13550 2470 13600 2770
rect 20200 2470 20250 2770
rect 12850 2465 14300 2470
rect 12850 2425 12855 2465
rect 12895 2425 13205 2465
rect 13245 2425 13555 2465
rect 13595 2425 13905 2465
rect 13945 2425 14255 2465
rect 14295 2425 14300 2465
rect 12850 2420 14300 2425
rect 19500 2465 20950 2470
rect 19500 2425 19505 2465
rect 19545 2425 19855 2465
rect 19895 2425 20205 2465
rect 20245 2425 20555 2465
rect 20595 2425 20905 2465
rect 20945 2425 20950 2465
rect 19500 2420 20950 2425
rect 13550 2120 13600 2420
rect 20200 2120 20250 2420
rect 12850 2115 14560 2120
rect 12850 2075 12855 2115
rect 12895 2075 13205 2115
rect 13245 2075 13555 2115
rect 13595 2075 13905 2115
rect 13945 2075 14255 2115
rect 14295 2075 14515 2115
rect 14555 2075 14560 2115
rect 12850 2070 14560 2075
rect 19240 2115 20950 2120
rect 19240 2075 19245 2115
rect 19285 2075 19505 2115
rect 19545 2075 19855 2115
rect 19895 2075 20205 2115
rect 20245 2075 20555 2115
rect 20595 2075 20905 2115
rect 20945 2075 20950 2115
rect 19240 2070 20950 2075
rect 24460 2115 24560 2120
rect 24460 2075 24515 2115
rect 24555 2075 24560 2115
rect 24460 2070 24560 2075
rect 29390 2115 29480 2120
rect 29390 2075 29395 2115
rect 29435 2075 29480 2115
rect 29390 2070 29480 2075
rect 13550 1770 13600 2070
rect 20200 1770 20250 2070
rect 12850 1765 14300 1770
rect 12850 1725 12855 1765
rect 12895 1725 13205 1765
rect 13245 1725 13555 1765
rect 13595 1725 13905 1765
rect 13945 1725 14255 1765
rect 14295 1725 14300 1765
rect 12850 1720 14300 1725
rect 19500 1765 20950 1770
rect 19500 1725 19505 1765
rect 19545 1725 19855 1765
rect 19895 1725 20205 1765
rect 20245 1725 20555 1765
rect 20595 1725 20905 1765
rect 20945 1725 20950 1765
rect 19500 1720 20950 1725
rect 13550 1420 13600 1720
rect 20200 1420 20250 1720
rect 12850 1415 14300 1420
rect 12850 1375 12855 1415
rect 12895 1375 13205 1415
rect 13245 1375 13555 1415
rect 13595 1375 13905 1415
rect 13945 1375 14255 1415
rect 14295 1375 14300 1415
rect 12850 1370 14300 1375
rect 19500 1415 20950 1420
rect 19500 1375 19505 1415
rect 19545 1375 19855 1415
rect 19895 1375 20205 1415
rect 20245 1375 20555 1415
rect 20595 1375 20905 1415
rect 20945 1375 20950 1415
rect 19500 1370 20950 1375
rect 13550 1070 13600 1370
rect 20200 1070 20250 1370
rect 12850 1065 14300 1070
rect 12850 1025 12855 1065
rect 12895 1025 13205 1065
rect 13245 1025 13555 1065
rect 13595 1025 13905 1065
rect 13945 1025 14255 1065
rect 14295 1025 14300 1065
rect 12850 1020 14300 1025
rect 19500 1065 20950 1070
rect 19500 1025 19505 1065
rect 19545 1025 19855 1065
rect 19895 1025 20205 1065
rect 20245 1025 20555 1065
rect 20595 1025 20905 1065
rect 20945 1025 20950 1065
rect 19500 1020 20950 1025
rect 13550 720 13600 1020
rect 20200 720 20250 1020
rect 12850 715 14300 720
rect 12850 675 12855 715
rect 12895 675 13205 715
rect 13245 675 13555 715
rect 13595 675 13905 715
rect 13945 675 14255 715
rect 14295 675 14300 715
rect 12850 670 14300 675
rect 19500 715 20950 720
rect 19500 675 19505 715
rect 19545 675 19855 715
rect 19895 675 20205 715
rect 20245 675 20555 715
rect 20595 675 20905 715
rect 20945 675 20950 715
rect 19500 670 20950 675
rect -115 660 5510 665
rect -115 620 -110 660
rect -70 620 5465 660
rect 5505 620 5510 660
rect -115 615 5510 620
rect -200 580 5595 585
rect -200 540 -195 580
rect -155 540 5550 580
rect 5590 540 5595 580
rect -200 535 5595 540
rect 13550 370 13600 670
rect 20200 370 20250 670
rect 12850 365 13600 370
rect 12850 325 12855 365
rect 12895 325 13205 365
rect 13245 325 13555 365
rect 13595 325 13600 365
rect 12850 320 13600 325
rect 13550 20 13600 320
rect 13900 365 13950 370
rect 13900 325 13905 365
rect 13945 325 13950 365
rect 13900 20 13950 325
rect 14250 365 14300 370
rect 14250 325 14255 365
rect 14295 325 14300 365
rect 14250 20 14300 325
rect 14600 365 14650 370
rect 14600 325 14605 365
rect 14645 325 14650 365
rect 14600 20 14650 325
rect 14950 365 15000 370
rect 14950 325 14955 365
rect 14995 325 15000 365
rect 14950 20 15000 325
rect 15300 365 15350 370
rect 15300 325 15305 365
rect 15345 325 15350 365
rect 15300 20 15350 325
rect 15650 365 15700 370
rect 15650 325 15655 365
rect 15695 325 15700 365
rect 15650 20 15700 325
rect 16000 365 16050 370
rect 16000 325 16005 365
rect 16045 325 16050 365
rect 16000 20 16050 325
rect 16350 365 16400 370
rect 16350 325 16355 365
rect 16395 325 16400 365
rect 16350 20 16400 325
rect 16700 365 16750 370
rect 16700 325 16705 365
rect 16745 325 16750 365
rect 16700 20 16750 325
rect 12850 15 16750 20
rect 12850 -25 12855 15
rect 12895 -25 13205 15
rect 13245 -25 13555 15
rect 13595 -25 13905 15
rect 13945 -25 14255 15
rect 14295 -25 14605 15
rect 14645 -25 14955 15
rect 14995 -25 15305 15
rect 15345 -25 15655 15
rect 15695 -25 16005 15
rect 16045 -25 16355 15
rect 16395 -25 16705 15
rect 16745 -25 16750 15
rect 12850 -30 16750 -25
rect 13550 -330 13600 -30
rect 12850 -335 13600 -330
rect 12850 -375 12855 -335
rect 12895 -375 13205 -335
rect 13245 -375 13555 -335
rect 13595 -375 13600 -335
rect 12850 -380 13600 -375
rect 13900 -335 13950 -30
rect 13900 -375 13905 -335
rect 13945 -375 13950 -335
rect 13900 -380 13950 -375
rect 14250 -335 14300 -30
rect 14250 -375 14255 -335
rect 14295 -375 14300 -335
rect 14250 -380 14300 -375
rect 14600 -335 14650 -30
rect 14600 -375 14605 -335
rect 14645 -375 14650 -335
rect 14600 -380 14650 -375
rect 14950 -335 15000 -30
rect 14950 -375 14955 -335
rect 14995 -375 15000 -335
rect 14950 -380 15000 -375
rect 15300 -335 15350 -30
rect 15300 -375 15305 -335
rect 15345 -375 15350 -335
rect 15300 -380 15350 -375
rect 15650 -335 15700 -30
rect 15650 -375 15655 -335
rect 15695 -375 15700 -335
rect 15650 -380 15700 -375
rect 16000 -335 16050 -30
rect 16000 -375 16005 -335
rect 16045 -375 16050 -335
rect 16000 -380 16050 -375
rect 16350 -335 16400 -30
rect 16350 -375 16355 -335
rect 16395 -375 16400 -335
rect 16350 -380 16400 -375
rect 16700 -335 16750 -30
rect 16700 -375 16705 -335
rect 16745 -375 16750 -335
rect 16700 -380 16750 -375
rect 17050 365 17100 370
rect 17050 325 17055 365
rect 17095 325 17100 365
rect 17050 20 17100 325
rect 17400 365 17450 370
rect 17400 325 17405 365
rect 17445 325 17450 365
rect 17400 20 17450 325
rect 17750 365 17800 370
rect 17750 325 17755 365
rect 17795 325 17800 365
rect 17750 20 17800 325
rect 18100 365 18150 370
rect 18100 325 18105 365
rect 18145 325 18150 365
rect 18100 20 18150 325
rect 18450 365 18500 370
rect 18450 325 18455 365
rect 18495 325 18500 365
rect 18450 20 18500 325
rect 18800 365 18850 370
rect 18800 325 18805 365
rect 18845 325 18850 365
rect 18800 20 18850 325
rect 19150 365 19200 370
rect 19150 325 19155 365
rect 19195 325 19200 365
rect 19150 20 19200 325
rect 19500 365 19550 370
rect 19500 325 19505 365
rect 19545 325 19550 365
rect 19500 20 19550 325
rect 19850 365 19900 370
rect 19850 325 19855 365
rect 19895 325 19900 365
rect 19850 20 19900 325
rect 20200 365 20950 370
rect 20200 325 20205 365
rect 20245 325 20555 365
rect 20595 325 20905 365
rect 20945 325 20950 365
rect 20200 320 20950 325
rect 20200 20 20250 320
rect 17050 15 20950 20
rect 17050 -25 17055 15
rect 17095 -25 17405 15
rect 17445 -25 17755 15
rect 17795 -25 18105 15
rect 18145 -25 18455 15
rect 18495 -25 18805 15
rect 18845 -25 19155 15
rect 19195 -25 19505 15
rect 19545 -25 19855 15
rect 19895 -25 20205 15
rect 20245 -25 20555 15
rect 20595 -25 20905 15
rect 20945 -25 20950 15
rect 17050 -30 20950 -25
rect 17050 -335 17100 -30
rect 17050 -375 17055 -335
rect 17095 -375 17100 -335
rect 17050 -380 17100 -375
rect 17400 -335 17450 -30
rect 17400 -375 17405 -335
rect 17445 -375 17450 -335
rect 17400 -380 17450 -375
rect 17750 -335 17800 -30
rect 17750 -375 17755 -335
rect 17795 -375 17800 -335
rect 17750 -380 17800 -375
rect 18100 -335 18150 -30
rect 18100 -375 18105 -335
rect 18145 -375 18150 -335
rect 18100 -380 18150 -375
rect 18450 -335 18500 -30
rect 18450 -375 18455 -335
rect 18495 -375 18500 -335
rect 18450 -380 18500 -375
rect 18800 -335 18850 -30
rect 18800 -375 18805 -335
rect 18845 -375 18850 -335
rect 18800 -380 18850 -375
rect 19150 -335 19200 -30
rect 19150 -375 19155 -335
rect 19195 -375 19200 -335
rect 19150 -380 19200 -375
rect 19500 -335 19550 -30
rect 19500 -375 19505 -335
rect 19545 -375 19550 -335
rect 19500 -380 19550 -375
rect 19850 -335 19900 -30
rect 19850 -375 19855 -335
rect 19895 -375 19900 -335
rect 19850 -380 19900 -375
rect 20200 -330 20250 -30
rect 20200 -335 20950 -330
rect 20200 -375 20205 -335
rect 20245 -375 20555 -335
rect 20595 -375 20905 -335
rect 20945 -375 20950 -335
rect 20200 -380 20950 -375
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 2950 1735 2950 1735 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2955 1590 2955 1590 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 1845 2945 1845 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3745 1530 3745 1530 3 FreeSans 400 0 40 0 V_p1
flabel metal1 2650 1155 2650 1155 3 FreeSans 400 0 200 0 START_UP
flabel metal2 3785 1785 3785 1785 5 FreeSans 400 0 0 -40 1st_Vout1
flabel metal2 455 3440 455 3440 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3375 2730 3375 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 2550 845 2550 845 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal2 5120 1590 5120 1590 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 4225 1785 4225 1785 5 FreeSans 400 0 0 -40 1st_Vout2
flabel metal2 5065 1845 5065 1845 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 4265 1530 4265 1530 7 FreeSans 400 0 -40 0 V_p2
flabel metal1 3275 350 3275 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3825 295 3825 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4015 350 4015 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4725 295 4725 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal1 4985 1110 4985 1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 4115 3135 4115 3135 1 FreeSans 400 0 0 40 PFET_GATE_10uA
flabel metal2 6080 3075 6080 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6100 3020 6100 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6080 2955 6080 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6100 1745 6100 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5590 4400 5590 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5505 4175 5505 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 2180 1010 2180 1010 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4635 2375 4635 2375 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
