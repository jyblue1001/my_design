* PEX produced on Mon Feb 24 09:44:57 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_cp_lf_magic_3.ext - technology: sky130A

.subckt pfd_cp_lf_magic_3 V_OUT VDDA F_REF F_VCO
X0 V_OUT.t99 a_6200_5250.t2 a_6200_5250.t3 V_OUT.t98 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X1 a_5970_4630.t10 opamp_cell_4_0.VIN- a_6200_5250.t5 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 pfd_8_0.DOWN_b.t0 VDDA.t130 pfd_8_0.DOWN_PFD_b.t1 V_OUT.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X3 a_870_1400.t1 pfd_8_0.QA_b.t3 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X4 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t2 VDDA.t108 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X5 V_OUT.t143 V_OUT.t141 V_OUT.t143 V_OUT.t142 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X6 VDDA.t8 pfd_8_0.UP_input.t13 opamp_cell_4_0.VIN+.t5 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X7 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.VIN+.t6 a_6320_5840.t1 V_OUT.t152 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X8 opamp_cell_4_0.n_right.t3 opamp_cell_4_0.n_left.t6 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X9 pfd_8_0.UP_input.t7 opamp_cell_4_0.n_right.t5 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 pfd_8_0.UP_input.t11 a_6490_4630.t5 V_OUT.t78 V_OUT.t77 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 a_2350_1400.t1 pfd_8_0.before_Reset.t3 V_OUT.t80 V_OUT.t79 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X12 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t3 V_OUT.t160 V_OUT.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X13 VDDA.t5 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t7 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X14 a_n30_1400.t1 F_REF.t0 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X15 V_OUT.t29 pfd_8_0.QA.t3 pfd_8_0.QA_b.t1 V_OUT.t28 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X16 a_6200_5250.t1 a_6200_5250.t0 V_OUT.t97 V_OUT.t96 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X17 a_6200_5250.t4 opamp_cell_4_0.VIN- a_5970_4630.t9 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X18 VDDA.t16 opamp_cell_4_0.p_bias.t9 a_5970_4630.t2 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 VDDA.t77 VDDA.t74 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X20 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN_b.t4 pfd_8_0.I_IN.t4 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X21 VDDA.t73 VDDA.t71 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X22 VDDA.t3 pfd_8_0.UP_input.t14 V_OUT.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X23 a_1910_2020.t0 pfd_8_0.QB.t3 V_OUT.t65 V_OUT.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 a_6220_5810.t7 a_6220_5810.t6 V_OUT.t62 V_OUT.t61 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X25 V_OUT.t14 pfd_8_0.DOWN_input.t3 V_OUT.t14 V_OUT.t13 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X26 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t2 VDDA.t129 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 a_6320_5840.t12 a_6220_5810.t9 V_OUT.t147 V_OUT.t146 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X28 pfd_8_0.UP_input.t3 pfd_8_0.UP.t2 pfd_8_0.UP_input.t2 V_OUT.t46 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X29 pfd_8_0.QA.t2 pfd_8_0.QA_b.t4 V_OUT.t19 V_OUT.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X30 a_5970_4630.t8 opamp_cell_4_0.p_bias.t10 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X31 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN.t2 pfd_8_0.I_IN.t5 V_OUT.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X32 V_OUT.t12 pfd_8_0.I_IN.t6 opamp_cell_4_0.VIN+.t0 V_OUT.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X33 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t1 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X34 a_870_640.t1 pfd_8_0.QB_b.t3 VDDA.t18 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X35 VDDA.t70 VDDA.t67 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X36 V_OUT.t9 loop_filter_2_0.R1_C1.t0 V_OUT.t8 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X37 VDDA.t110 a_2530_190.t2 a_2200_190.t0 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X38 V_OUT.t140 V_OUT.t138 V_OUT.t140 V_OUT.t139 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X39 V_OUT.t137 V_OUT.t134 V_OUT.t136 V_OUT.t135 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X40 opamp_cell_4_0.p_bias.t5 opamp_cell_4_0.p_bias.t4 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X41 VDDA.t66 VDDA.t64 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X42 V_OUT.t70 pfd_8_0.UP_input.t15 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X43 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t5 V_OUT.t33 V_OUT.t32 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X44 V_OUT.t162 a_2530_190.t3 a_2200_190.t1 V_OUT.t161 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X45 pfd_8_0.F.t1 pfd_8_0.QB_b.t4 V_OUT.t59 V_OUT.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X46 V_OUT.t133 V_OUT.t130 V_OUT.t132 V_OUT.t131 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X47 pfd_8_0.UP_input.t16 a_9360_6440.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X48 V_OUT.t31 pfd_8_0.DOWN_input.t4 V_OUT.t31 V_OUT.t30 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X49 pfd_8_0.UP_b.t1 pfd_8_0.UP.t3 V_OUT.t149 V_OUT.t148 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X50 V_OUT.t151 pfd_8_0.E_b.t3 pfd_8_0.E.t2 V_OUT.t150 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X51 V_OUT.t50 a_6220_5810.t10 a_6320_5840.t4 V_OUT.t49 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X52 a_1390_640.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t1 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X53 a_2350_1400.t0 pfd_8_0.before_Reset.t4 VDDA.t107 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X54 opamp_cell_4_0.VIN+.t1 pfd_8_0.I_IN.t7 V_OUT.t45 V_OUT.t44 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X55 V_OUT.t17 a_6220_5810.t4 a_6220_5810.t5 V_OUT.t16 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X56 V_OUT.t129 V_OUT.t127 V_OUT.t129 V_OUT.t128 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X57 a_5970_4630.t7 a_5970_4630.t6 a_5970_4630.t7 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X58 pfd_8_0.F_b.t2 pfd_8_0.F.t4 V_OUT.t84 V_OUT.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X59 VDDA.t83 pfd_8_0.UP_input.t17 V_OUT.t63 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 V_OUT.t163 loop_filter_2_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X61 VDDA.t27 pfd_8_0.F.t5 a_490_640.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X62 VDDA.t63 VDDA.t61 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X63 V_OUT.t126 V_OUT.t124 V_OUT.t126 V_OUT.t125 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X64 pfd_8_0.QA_b.t0 pfd_8_0.QA.t4 a_n30_1400.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X65 V_OUT.t123 V_OUT.t121 V_OUT.t123 V_OUT.t122 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X66 pfd_8_0.UP_input.t18 charge_pump_cell_6_0.UP_b.t0 sky130_fd_pr__cap_mim_m3_1 l=16 w=13.9
X67 V_OUT.t27 pfd_8_0.F.t6 pfd_8_0.QB.t0 V_OUT.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X68 V_OUT.t120 V_OUT.t118 V_OUT.t120 V_OUT.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X69 pfd_8_0.before_Reset.t1 pfd_8_0.QB.t4 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X70 V_OUT.t76 a_6490_4630.t6 pfd_8_0.UP_input.t10 V_OUT.t75 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X71 VDDA.t93 opamp_cell_4_0.n_right.t6 pfd_8_0.UP_input.t6 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X72 opamp_cell_4_0.VIN+.t4 pfd_8_0.UP_input.t19 VDDA.t99 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X73 pfd_8_0.UP_input.t1 pfd_8_0.UP_b.t2 pfd_8_0.UP_input.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.15
X74 a_490_1400.t1 pfd_8_0.QA_b.t5 pfd_8_0.QA.t1 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X75 V_OUT.t55 pfd_8_0.UP_input.t20 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X76 V_OUT.t21 pfd_8_0.Reset.t2 pfd_8_0.E_b.t0 V_OUT.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X77 a_2530_190.t1 a_2350_1400.t2 V_OUT.t69 V_OUT.t68 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X78 VDDA.t42 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X79 a_6320_5840.t11 opamp_cell_4_0.VIN- opamp_cell_4_0.n_left.t5 V_OUT.t145 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X80 V_OUT.t89 pfd_8_0.I_IN.t2 pfd_8_0.I_IN.t3 V_OUT.t88 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X81 pfd_8_0.E.t0 pfd_8_0.E_b.t4 a_870_1400.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X82 pfd_8_0.UP_b.t0 pfd_8_0.UP.t4 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X83 a_5970_4630.t5 a_5970_4630.t3 a_5970_4630.t4 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X84 V_OUT.t117 V_OUT.t114 V_OUT.t116 V_OUT.t115 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X85 pfd_8_0.DOWN_input.t5 charge_pump_cell_6_0.DOWN.t0 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.8
X86 VDDA.t23 a_1870_190.t2 pfd_8_0.Reset.t0 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X87 pfd_8_0.UP_input.t9 a_6490_4630.t7 V_OUT.t74 V_OUT.t73 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X88 pfd_8_0.UP_input.t5 opamp_cell_4_0.n_right.t7 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X89 V_OUT.t42 a_1870_190.t3 pfd_8_0.Reset.t1 V_OUT.t41 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X90 VDDA.t60 VDDA.t57 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X91 opamp_cell_4_0.p_bias.t3 opamp_cell_4_0.p_bias.t2 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X92 pfd_8_0.I_IN.t1 pfd_8_0.I_IN.t0 V_OUT.t67 V_OUT.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X93 opamp_cell_4_0.p_bias.t8 a_6220_5810.t8 V_OUT.t156 sky130_fd_pr__res_xhigh_po_5p73 l=1
X94 opamp_cell_4_0.n_left.t1 opamp_cell_4_0.n_left.t0 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X95 V_OUT.t108 V_OUT.t109 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X96 opamp_cell_4_0.n_left.t4 opamp_cell_4_0.VIN- a_6320_5840.t10 V_OUT.t144 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X97 a_5970_4630.t1 opamp_cell_4_0.p_bias.t11 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X98 pfd_8_0.before_Reset.t0 pfd_8_0.QA.t5 a_1910_2020.t1 V_OUT.t10 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X99 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t6 V_OUT.t35 V_OUT.t34 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X100 V_OUT.t113 V_OUT.t110 V_OUT.t112 V_OUT.t111 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X101 V_OUT.t57 pfd_8_0.E.t4 pfd_8_0.QA.t0 V_OUT.t56 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X102 a_9360_6440.t0 a_6490_4630.t2 V_OUT.t60 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X103 pfd_8_0.F.t0 pfd_8_0.F_b.t3 a_870_640.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X104 VDDA.t21 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X105 VDDA.t56 VDDA.t54 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X106 V_OUT.t107 V_OUT.t104 V_OUT.t106 V_OUT.t105 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X107 a_2530_190.t0 a_2350_1400.t3 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X108 V_OUT.t91 a_6220_5810.t2 a_6220_5810.t3 V_OUT.t90 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X109 V_OUT.t72 a_6490_4630.t8 pfd_8_0.UP_input.t8 V_OUT.t71 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X110 VDDA.t89 opamp_cell_4_0.n_right.t8 pfd_8_0.UP_input.t4 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X111 VDDA.t53 VDDA.t50 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X112 V_OUT.t86 pfd_8_0.F_b.t4 pfd_8_0.F.t2 V_OUT.t85 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X113 V_OUT.t103 V_OUT.t100 V_OUT.t102 V_OUT.t101 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X114 V_OUT.t5 a_6220_5810.t11 a_6320_5840.t0 V_OUT.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X115 pfd_8_0.QB_b.t0 pfd_8_0.QB.t5 a_n30_640.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X116 V_OUT.t95 a_6200_5250.t6 a_6490_4630.t4 V_OUT.t94 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X117 a_5970_4630.t12 opamp_cell_4_0.VIN+.t7 a_6490_4630.t1 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X118 VDDA.t12 opamp_cell_4_0.p_bias.t12 a_5970_4630.t0 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X119 VDDA.t36 pfd_8_0.Reset.t4 a_1390_640.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X120 VDDA.t33 opamp_cell_4_0.p_bias.t0 opamp_cell_4_0.p_bias.t1 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X121 pfd_8_0.UP_input.t12 pfd_8_0.UP.t5 VDDA.t122 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X122 opamp_cell_4_0.n_right.t4 charge_pump_cell_6_0.UP_b.t1 V_OUT.t87 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X123 VDDA.t49 VDDA.t46 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X124 a_6320_5840.t9 a_6320_5840.t7 a_6320_5840.t8 V_OUT.t43 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X125 V_OUT.t3 pfd_8_0.QB.t6 pfd_8_0.QB_b.t1 V_OUT.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X126 a_6320_5840.t3 a_6220_5810.t12 V_OUT.t48 V_OUT.t47 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X127 V_OUT.t7 pfd_8_0.Reset.t5 pfd_8_0.F_b.t0 V_OUT.t6 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X128 a_6320_5840.t6 a_6320_5840.t5 a_6320_5840.t6 V_OUT.t40 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X129 VDDA.t45 VDDA.t43 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X130 a_6220_5810.t1 a_6220_5810.t0 V_OUT.t39 V_OUT.t38 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X131 pfd_8_0.E.t1 pfd_8_0.QA_b.t6 V_OUT.t154 V_OUT.t153 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X132 VDDA.t120 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t2 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X133 a_n30_640.t1 F_VCO.t0 VDDA.t111 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X134 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t8 VDDA.t118 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X135 a_6490_4630.t3 a_6200_5250.t7 V_OUT.t93 V_OUT.t92 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X136 a_6490_4630.t0 opamp_cell_4_0.VIN+.t8 a_5970_4630.t11 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X137 VDDA.t123 pfd_8_0.E.t5 a_490_1400.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X138 VDDA.t128 a_2200_190.t2 a_1870_190.t0 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X139 pfd_8_0.QA_b.t2 F_REF.t1 V_OUT.t82 V_OUT.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X140 pfd_8_0.QB_b.t2 F_VCO.t1 V_OUT.t23 V_OUT.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X141 a_490_640.t1 pfd_8_0.QB_b.t5 pfd_8_0.QB.t2 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X142 VDDA.t1 pfd_8_0.UP_input.t21 opamp_cell_4_0.VIN+.t3 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X143 V_OUT.t25 a_2200_190.t3 a_1870_190.t1 V_OUT.t24 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X144 a_6320_5840.t2 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t0 V_OUT.t155 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X145 VDDA.t81 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t2 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X146 pfd_8_0.QB.t1 pfd_8_0.QB_b.t6 V_OUT.t54 V_OUT.t53 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X147 pfd_8_0.DOWN_PFD_b.t2 pfd_8_0.QB.t7 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X148 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t3 V_OUT.t158 V_OUT.t157 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X149 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 V_OUT.t37 V_OUT.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X150 pfd_8_0.E_b.t2 pfd_8_0.E.t6 V_OUT.t52 V_OUT.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X151 opamp_cell_4_0.VIN+.t2 pfd_8_0.UP_input.t22 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X152 pfd_8_0.DOWN_b.t1 V_OUT.t164 pfd_8_0.DOWN_PFD_b.t3 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
R0 a_6200_5250.n5 a_6200_5250.n4 427.647
R1 a_6200_5250.n1 a_6200_5250.t6 321.334
R2 a_6200_5250.n4 a_6200_5250.n0 210.601
R3 a_6200_5250.n2 a_6200_5250.n1 208.868
R4 a_6200_5250.n3 a_6200_5250.t0 174.056
R5 a_6200_5250.n4 a_6200_5250.n3 152
R6 a_6200_5250.n1 a_6200_5250.t7 112.468
R7 a_6200_5250.n2 a_6200_5250.t2 112.468
R8 a_6200_5250.n3 a_6200_5250.n2 61.5894
R9 a_6200_5250.n0 a_6200_5250.t3 60.0005
R10 a_6200_5250.n0 a_6200_5250.t1 60.0005
R11 a_6200_5250.n5 a_6200_5250.t5 49.2505
R12 a_6200_5250.t4 a_6200_5250.n5 49.2505
R13 V_OUT.n384 V_OUT.n383 348175
R14 V_OUT.n383 V_OUT.n382 292776
R15 V_OUT.n280 V_OUT.t46 25257.7
R16 V_OUT.n286 V_OUT.n280 15376.3
R17 V_OUT.n382 V_OUT.t32 2083.03
R18 V_OUT.t83 V_OUT.t85 1939.79
R19 V_OUT.t53 V_OUT.t2 1939.79
R20 V_OUT.n224 V_OUT.n36 1860.65
R21 V_OUT.t1 V_OUT.t36 1845.16
R22 V_OUT.t15 V_OUT.t159 1372.04
R23 V_OUT.t41 V_OUT.n371 1253.76
R24 V_OUT.n378 V_OUT.n377 1230.11
R25 V_OUT.n270 V_OUT.n269 1186
R26 V_OUT.n223 V_OUT.n222 1186
R27 V_OUT.n216 V_OUT.n215 1186
R28 V_OUT.n277 V_OUT.n276 1186
R29 V_OUT.n279 V_OUT.n278 1170
R30 V_OUT.n381 V_OUT.t15 1064.52
R31 V_OUT.n379 V_OUT.t1 1064.52
R32 V_OUT.n382 V_OUT.n366 1052.76
R33 V_OUT.t161 V_OUT.n375 922.582
R34 V_OUT.t24 V_OUT.n373 922.582
R35 V_OUT.n118 V_OUT.t81 783.001
R36 V_OUT.t32 V_OUT.n381 780.645
R37 V_OUT.t159 V_OUT.n379 780.645
R38 V_OUT.t36 V_OUT.n378 780.645
R39 V_OUT.n338 V_OUT.n337 669.307
R40 V_OUT.n340 V_OUT.n48 669.307
R41 V_OUT.n333 V_OUT.n332 669.307
R42 V_OUT.n330 V_OUT.n52 669.307
R43 V_OUT.n285 V_OUT.n284 669.307
R44 V_OUT.n288 V_OUT.n287 669.307
R45 V_OUT.n377 V_OUT.t161 638.711
R46 V_OUT.n375 V_OUT.t24 638.711
R47 V_OUT.n373 V_OUT.t41 638.711
R48 V_OUT.n371 V_OUT.t6 638.711
R49 V_OUT.t58 V_OUT.n369 638.711
R50 V_OUT.n369 V_OUT.t26 638.711
R51 V_OUT.n384 V_OUT.t22 638.711
R52 V_OUT.t150 V_OUT.t51 601.333
R53 V_OUT.t28 V_OUT.t18 601.333
R54 V_OUT.t142 V_OUT.t13 593.865
R55 V_OUT.t13 V_OUT.t30 593.865
R56 V_OUT.t30 V_OUT.t111 593.865
R57 V_OUT.t11 V_OUT.t125 593.865
R58 V_OUT.t44 V_OUT.t11 593.865
R59 V_OUT.t105 V_OUT.t44 593.865
R60 V_OUT.t119 V_OUT.t88 593.865
R61 V_OUT.t88 V_OUT.t66 593.865
R62 V_OUT.t66 V_OUT.t101 593.865
R63 V_OUT.n369 V_OUT.n368 585.003
R64 V_OUT.n117 V_OUT.n116 585.003
R65 V_OUT.n114 V_OUT.n113 585.001
R66 V_OUT.n112 V_OUT.n111 585.001
R67 V_OUT.n110 V_OUT.n109 585.001
R68 V_OUT.n89 V_OUT.n37 585.001
R69 V_OUT.n268 V_OUT.n267 585.001
R70 V_OUT.n225 V_OUT.n224 585.001
R71 V_OUT.n186 V_OUT.n185 585.001
R72 V_OUT.n86 V_OUT.n85 585.001
R73 V_OUT.n84 V_OUT.n81 585.001
R74 V_OUT.n381 V_OUT.n380 585.001
R75 V_OUT.n379 V_OUT.n8 585.001
R76 V_OUT.n378 V_OUT.n14 585.001
R77 V_OUT.n377 V_OUT.n376 585.001
R78 V_OUT.n375 V_OUT.n374 585.001
R79 V_OUT.n373 V_OUT.n372 585.001
R80 V_OUT.n371 V_OUT.n370 585.001
R81 V_OUT.n385 V_OUT.n384 585.001
R82 V_OUT.n283 V_OUT.n281 585
R83 V_OUT.n78 V_OUT.n76 585
R84 V_OUT.n56 V_OUT.n53 585
R85 V_OUT.n59 V_OUT.n58 585
R86 V_OUT.n51 V_OUT.n50 585
R87 V_OUT.n342 V_OUT.n341 585
R88 V_OUT.n365 V_OUT.n364 585
R89 V_OUT.n366 V_OUT.n365 585
R90 V_OUT.n363 V_OUT.n40 585
R91 V_OUT.n361 V_OUT.n360 585
R92 V_OUT.n359 V_OUT.n39 585
R93 V_OUT.n366 V_OUT.n39 585
R94 V_OUT.n12 V_OUT.t164 566.966
R95 V_OUT.n286 V_OUT.t142 566.871
R96 V_OUT.n334 V_OUT.t111 566.871
R97 V_OUT.t125 V_OUT.n334 566.871
R98 V_OUT.n339 V_OUT.t105 566.871
R99 V_OUT.n339 V_OUT.t119 566.871
R100 V_OUT.n366 V_OUT.t101 566.871
R101 V_OUT.t60 V_OUT.n277 564.696
R102 V_OUT.n280 V_OUT.t87 534.24
R103 V_OUT.t6 V_OUT.t83 520.431
R104 V_OUT.t85 V_OUT.t58 520.431
R105 V_OUT.t26 V_OUT.t53 520.431
R106 V_OUT.t2 V_OUT.t22 520.431
R107 V_OUT.t87 V_OUT.t60 509.197
R108 V_OUT.t46 V_OUT.t148 425.334
R109 V_OUT.n85 V_OUT.t68 418
R110 V_OUT.n186 V_OUT.t157 344.668
R111 V_OUT.t34 V_OUT.n84 344.668
R112 V_OUT.n335 V_OUT.t118 336.329
R113 V_OUT.n335 V_OUT.t104 336.329
R114 V_OUT.n54 V_OUT.t124 336.329
R115 V_OUT.n54 V_OUT.t110 336.329
R116 V_OUT.n358 V_OUT.t100 320.7
R117 V_OUT.n289 V_OUT.t141 320.7
R118 V_OUT.n280 V_OUT.n279 309.736
R119 V_OUT.n187 V_OUT.t121 304.634
R120 V_OUT.n271 V_OUT.t134 304.634
R121 V_OUT.n221 V_OUT.t114 304.634
R122 V_OUT.n217 V_OUT.t127 304.634
R123 V_OUT.n266 V_OUT.t138 292.584
R124 V_OUT.n226 V_OUT.t130 292.584
R125 V_OUT.t79 V_OUT.n37 286
R126 V_OUT.t10 V_OUT.n110 286
R127 V_OUT.n286 V_OUT.n285 250.349
R128 V_OUT.n287 V_OUT.n286 250.349
R129 V_OUT.n334 V_OUT.n333 250.349
R130 V_OUT.n334 V_OUT.n52 250.349
R131 V_OUT.n339 V_OUT.n338 250.349
R132 V_OUT.n340 V_OUT.n339 250.349
R133 V_OUT.n366 V_OUT.n38 250.349
R134 V_OUT.n276 V_OUT.t123 245
R135 V_OUT.n270 V_OUT.t137 245
R136 V_OUT.n222 V_OUT.t117 245
R137 V_OUT.n216 V_OUT.t129 245
R138 V_OUT.n69 V_OUT.n68 242.903
R139 V_OUT.t148 V_OUT.n186 227.333
R140 V_OUT.n84 V_OUT.t157 227.333
R141 V_OUT.n85 V_OUT.t34 227.333
R142 V_OUT.n114 V_OUT.n112 205.333
R143 V_OUT.n273 V_OUT.n189 204.201
R144 V_OUT.n219 V_OUT.n213 204.201
R145 V_OUT.n220 V_OUT.n212 204.201
R146 V_OUT.n218 V_OUT.n214 204.201
R147 V_OUT.n272 V_OUT.n190 204.201
R148 V_OUT.n275 V_OUT.n274 204.201
R149 V_OUT.n391 V_OUT.t3 198.058
R150 V_OUT.n32 V_OUT.t54 198.058
R151 V_OUT.n405 V_OUT.t86 198.058
R152 V_OUT.n410 V_OUT.t84 198.058
R153 V_OUT.n143 V_OUT.t52 198.058
R154 V_OUT.n138 V_OUT.t151 198.058
R155 V_OUT.n105 V_OUT.t19 198.058
R156 V_OUT.n124 V_OUT.t29 198.058
R157 V_OUT.n110 V_OUT.t79 198
R158 V_OUT.n112 V_OUT.t64 198
R159 V_OUT.t20 V_OUT.n114 198
R160 V_OUT.n117 V_OUT.t153 198
R161 V_OUT.t56 V_OUT.n117 198
R162 V_OUT.n341 V_OUT.n51 197
R163 V_OUT.n58 V_OUT.n53 197
R164 V_OUT.n281 V_OUT.n78 197
R165 V_OUT.n365 V_OUT.n40 197
R166 V_OUT.n360 V_OUT.n39 197
R167 V_OUT.n337 V_OUT.n336 185
R168 V_OUT.n336 V_OUT.n48 185
R169 V_OUT.n332 V_OUT.n331 185
R170 V_OUT.n331 V_OUT.n330 185
R171 V_OUT.n284 V_OUT.n77 185
R172 V_OUT.n288 V_OUT.n77 185
R173 V_OUT.n364 V_OUT.n41 185
R174 V_OUT.n359 V_OUT.n41 185
R175 V_OUT.n69 V_OUT.n67 172.502
R176 V_OUT.n337 V_OUT.n335 166.63
R177 V_OUT.n332 V_OUT.n54 166.63
R178 V_OUT.t64 V_OUT.t10 161.333
R179 V_OUT.t51 V_OUT.t20 161.333
R180 V_OUT.t153 V_OUT.t150 161.333
R181 V_OUT.t18 V_OUT.t56 161.333
R182 V_OUT.t81 V_OUT.t28 161.333
R183 V_OUT.n3 V_OUT.t9 158.893
R184 V_OUT.n267 V_OUT.t140 134.501
R185 V_OUT.n225 V_OUT.t133 134.501
R186 V_OUT.n31 V_OUT.t27 130.713
R187 V_OUT.n385 V_OUT.t23 130.001
R188 V_OUT.n370 V_OUT.t7 130.001
R189 V_OUT.n372 V_OUT.t42 130.001
R190 V_OUT.n374 V_OUT.t25 130.001
R191 V_OUT.n376 V_OUT.t162 130.001
R192 V_OUT.n118 V_OUT.t82 130.001
R193 V_OUT.n113 V_OUT.t21 130.001
R194 V_OUT.n111 V_OUT.t65 130.001
R195 V_OUT.n109 V_OUT.t80 130.001
R196 V_OUT.n89 V_OUT.t69 130.001
R197 V_OUT.n115 V_OUT.t154 130.001
R198 V_OUT.n104 V_OUT.t57 130.001
R199 V_OUT.n367 V_OUT.t59 130.001
R200 V_OUT.n14 V_OUT.t37 122.501
R201 V_OUT.n8 V_OUT.t160 122.501
R202 V_OUT.n380 V_OUT.t33 122.501
R203 V_OUT.n86 V_OUT.t35 122.501
R204 V_OUT.n185 V_OUT.t149 122.501
R205 V_OUT.n81 V_OUT.t158 122.501
R206 V_OUT.n73 V_OUT.n72 118.35
R207 V_OUT.n268 V_OUT.t40 112.157
R208 V_OUT.n74 V_OUT.n73 106.662
R209 V_OUT.n194 V_OUT.n193 97.8707
R210 V_OUT.n198 V_OUT.n197 97.8707
R211 V_OUT.n202 V_OUT.n201 97.8707
R212 V_OUT.n206 V_OUT.n205 97.8707
R213 V_OUT.n211 V_OUT.n210 97.8707
R214 V_OUT.n215 V_OUT.t61 97.7783
R215 V_OUT.n277 V_OUT.t122 94.9025
R216 V_OUT.n269 V_OUT.t135 94.9025
R217 V_OUT.n298 V_OUT.n64 92.2612
R218 V_OUT.n291 V_OUT.n75 92.2612
R219 V_OUT.n324 V_OUT.n304 92.2612
R220 V_OUT.n318 V_OUT.n307 92.2612
R221 V_OUT.n346 V_OUT.n345 92.2612
R222 V_OUT.n353 V_OUT.n352 92.2612
R223 V_OUT.n336 V_OUT.n49 91.3721
R224 V_OUT.n344 V_OUT.n47 91.3721
R225 V_OUT.n344 V_OUT.n343 91.3721
R226 V_OUT.n331 V_OUT.n57 91.3721
R227 V_OUT.n303 V_OUT.n55 91.3721
R228 V_OUT.n303 V_OUT.n60 91.3721
R229 V_OUT.n282 V_OUT.n77 90.7567
R230 V_OUT.n362 V_OUT.n41 90.7567
R231 V_OUT.t61 V_OUT.t43 89.1508
R232 V_OUT.n223 V_OUT.t131 86.275
R233 V_OUT.n285 V_OUT.n281 84.306
R234 V_OUT.n287 V_OUT.n78 84.306
R235 V_OUT.n333 V_OUT.n53 84.306
R236 V_OUT.n58 V_OUT.n52 84.306
R237 V_OUT.n338 V_OUT.n51 84.306
R238 V_OUT.n341 V_OUT.n340 84.306
R239 V_OUT.n40 V_OUT.n38 84.306
R240 V_OUT.n360 V_OUT.n38 84.306
R241 V_OUT.n278 V_OUT.t108 84.2543
R242 V_OUT.n219 V_OUT.n218 83.2005
R243 V_OUT.n220 V_OUT.n219 83.2005
R244 V_OUT.n278 V_OUT.t163 81.0543
R245 V_OUT.n383 V_OUT.n36 80.6672
R246 V_OUT.t16 V_OUT.t128 77.6476
R247 V_OUT.t75 V_OUT.t122 74.7717
R248 V_OUT.t73 V_OUT.t75 74.7717
R249 V_OUT.t71 V_OUT.t73 74.7717
R250 V_OUT.t77 V_OUT.t71 74.7717
R251 V_OUT.t135 V_OUT.t77 74.7717
R252 V_OUT.n269 V_OUT.n268 74.7717
R253 V_OUT.t145 V_OUT.t152 74.7717
R254 V_OUT.t94 V_OUT.t92 74.7717
R255 V_OUT.t96 V_OUT.t115 74.7717
R256 V_OUT.n383 V_OUT.n37 73.3338
R257 V_OUT.t155 V_OUT.t139 71.8959
R258 V_OUT.t49 V_OUT.t98 71.8959
R259 V_OUT.n274 V_OUT.n273 66.5605
R260 V_OUT.n273 V_OUT.n272 66.5605
R261 V_OUT.t144 V_OUT.t146 66.1443
R262 V_OUT.n273 V_OUT.n188 65.9634
R263 V_OUT.n119 V_OUT.n118 60.29
R264 V_OUT.n113 V_OUT.n97 60.29
R265 V_OUT.n111 V_OUT.n96 60.29
R266 V_OUT.n109 V_OUT.n92 60.29
R267 V_OUT.n90 V_OUT.n89 60.29
R268 V_OUT.n376 V_OUT.n17 60.29
R269 V_OUT.n374 V_OUT.n19 60.29
R270 V_OUT.n372 V_OUT.n21 60.29
R271 V_OUT.n370 V_OUT.n25 60.29
R272 V_OUT.n386 V_OUT.n385 60.29
R273 V_OUT.n189 V_OUT.t74 60.0005
R274 V_OUT.n189 V_OUT.t72 60.0005
R275 V_OUT.n213 V_OUT.t93 60.0005
R276 V_OUT.n213 V_OUT.t99 60.0005
R277 V_OUT.n212 V_OUT.t97 60.0005
R278 V_OUT.n212 V_OUT.t116 60.0005
R279 V_OUT.t129 V_OUT.n214 60.0005
R280 V_OUT.n214 V_OUT.t95 60.0005
R281 V_OUT.n190 V_OUT.t78 60.0005
R282 V_OUT.n190 V_OUT.t136 60.0005
R283 V_OUT.t123 V_OUT.n275 60.0005
R284 V_OUT.n275 V_OUT.t76 60.0005
R285 V_OUT.n171 V_OUT.n86 59.5478
R286 V_OUT.n185 V_OUT.n184 59.5478
R287 V_OUT.n178 V_OUT.n81 59.5478
R288 V_OUT.n450 V_OUT.n8 58.9809
R289 V_OUT.n438 V_OUT.n14 58.9809
R290 V_OUT.n380 V_OUT.n4 58.9809
R291 V_OUT.n279 V_OUT.t8 56.0165
R292 V_OUT.n132 V_OUT.n104 54.4005
R293 V_OUT.n115 V_OUT.n103 54.4005
R294 V_OUT.n367 V_OUT.n30 54.4005
R295 V_OUT.n399 V_OUT.n31 54.4005
R296 V_OUT.t90 V_OUT.t144 48.8894
R297 V_OUT.t68 V_OUT.n36 44.0005
R298 V_OUT.t4 V_OUT.t155 43.1378
R299 V_OUT.t98 V_OUT.t47 43.1378
R300 V_OUT.n219 V_OUT.n208 41.6005
R301 V_OUT.n463 V_OUT.n1 41.3005
R302 V_OUT.n263 V_OUT.n188 39.4985
R303 V_OUT.t128 V_OUT.t38 37.3861
R304 V_OUT.t38 V_OUT.t94 37.3861
R305 V_OUT.n119 V_OUT.n108 33.0991
R306 V_OUT.n386 V_OUT.n35 33.0991
R307 V_OUT.n299 V_OUT.n298 32.0005
R308 V_OUT.n299 V_OUT.n61 32.0005
R309 V_OUT.n293 V_OUT.n292 32.0005
R310 V_OUT.n293 V_OUT.n65 32.0005
R311 V_OUT.n297 V_OUT.n65 32.0005
R312 V_OUT.n325 V_OUT.n62 32.0005
R313 V_OUT.n323 V_OUT.n305 32.0005
R314 V_OUT.n319 V_OUT.n305 32.0005
R315 V_OUT.n319 V_OUT.n318 32.0005
R316 V_OUT.n317 V_OUT.n308 32.0005
R317 V_OUT.n313 V_OUT.n308 32.0005
R318 V_OUT.n312 V_OUT.n311 32.0005
R319 V_OUT.n311 V_OUT.n46 32.0005
R320 V_OUT.n350 V_OUT.n44 32.0005
R321 V_OUT.n351 V_OUT.n350 32.0005
R322 V_OUT.n357 V_OUT.n42 32.0005
R323 V_OUT.n263 V_OUT.n262 32.0005
R324 V_OUT.n262 V_OUT.n261 32.0005
R325 V_OUT.n261 V_OUT.n192 32.0005
R326 V_OUT.n257 V_OUT.n192 32.0005
R327 V_OUT.n257 V_OUT.n256 32.0005
R328 V_OUT.n256 V_OUT.n255 32.0005
R329 V_OUT.n255 V_OUT.n196 32.0005
R330 V_OUT.n251 V_OUT.n196 32.0005
R331 V_OUT.n251 V_OUT.n250 32.0005
R332 V_OUT.n250 V_OUT.n249 32.0005
R333 V_OUT.n249 V_OUT.n200 32.0005
R334 V_OUT.n245 V_OUT.n200 32.0005
R335 V_OUT.n245 V_OUT.n244 32.0005
R336 V_OUT.n244 V_OUT.n243 32.0005
R337 V_OUT.n243 V_OUT.n204 32.0005
R338 V_OUT.n239 V_OUT.n238 32.0005
R339 V_OUT.n238 V_OUT.n237 32.0005
R340 V_OUT.n237 V_OUT.n209 32.0005
R341 V_OUT.n232 V_OUT.n209 32.0005
R342 V_OUT.n232 V_OUT.n231 32.0005
R343 V_OUT.n231 V_OUT.n230 32.0005
R344 V_OUT.n184 V_OUT.n79 32.0005
R345 V_OUT.n180 V_OUT.n79 32.0005
R346 V_OUT.n180 V_OUT.n179 32.0005
R347 V_OUT.n177 V_OUT.n82 32.0005
R348 V_OUT.n173 V_OUT.n82 32.0005
R349 V_OUT.n173 V_OUT.n172 32.0005
R350 V_OUT.n170 V_OUT.n87 32.0005
R351 V_OUT.n166 V_OUT.n87 32.0005
R352 V_OUT.n166 V_OUT.n165 32.0005
R353 V_OUT.n165 V_OUT.n164 32.0005
R354 V_OUT.n161 V_OUT.n160 32.0005
R355 V_OUT.n160 V_OUT.n159 32.0005
R356 V_OUT.n156 V_OUT.n155 32.0005
R357 V_OUT.n155 V_OUT.n154 32.0005
R358 V_OUT.n154 V_OUT.n94 32.0005
R359 V_OUT.n150 V_OUT.n149 32.0005
R360 V_OUT.n149 V_OUT.n148 32.0005
R361 V_OUT.n145 V_OUT.n144 32.0005
R362 V_OUT.n144 V_OUT.n143 32.0005
R363 V_OUT.n143 V_OUT.n99 32.0005
R364 V_OUT.n139 V_OUT.n99 32.0005
R365 V_OUT.n139 V_OUT.n138 32.0005
R366 V_OUT.n138 V_OUT.n137 32.0005
R367 V_OUT.n137 V_OUT.n101 32.0005
R368 V_OUT.n131 V_OUT.n130 32.0005
R369 V_OUT.n130 V_OUT.n105 32.0005
R370 V_OUT.n126 V_OUT.n105 32.0005
R371 V_OUT.n126 V_OUT.n125 32.0005
R372 V_OUT.n125 V_OUT.n124 32.0005
R373 V_OUT.n124 V_OUT.n107 32.0005
R374 V_OUT.n120 V_OUT.n107 32.0005
R375 V_OUT.n458 V_OUT.n457 32.0005
R376 V_OUT.n457 V_OUT.n456 32.0005
R377 V_OUT.n456 V_OUT.n6 32.0005
R378 V_OUT.n452 V_OUT.n6 32.0005
R379 V_OUT.n452 V_OUT.n451 32.0005
R380 V_OUT.n451 V_OUT.n450 32.0005
R381 V_OUT.n450 V_OUT.n9 32.0005
R382 V_OUT.n446 V_OUT.n9 32.0005
R383 V_OUT.n446 V_OUT.n445 32.0005
R384 V_OUT.n445 V_OUT.n444 32.0005
R385 V_OUT.n444 V_OUT.n11 32.0005
R386 V_OUT.n440 V_OUT.n11 32.0005
R387 V_OUT.n440 V_OUT.n439 32.0005
R388 V_OUT.n437 V_OUT.n15 32.0005
R389 V_OUT.n433 V_OUT.n15 32.0005
R390 V_OUT.n433 V_OUT.n432 32.0005
R391 V_OUT.n432 V_OUT.n431 32.0005
R392 V_OUT.n428 V_OUT.n427 32.0005
R393 V_OUT.n427 V_OUT.n426 32.0005
R394 V_OUT.n423 V_OUT.n422 32.0005
R395 V_OUT.n422 V_OUT.n421 32.0005
R396 V_OUT.n418 V_OUT.n417 32.0005
R397 V_OUT.n417 V_OUT.n416 32.0005
R398 V_OUT.n416 V_OUT.n23 32.0005
R399 V_OUT.n412 V_OUT.n411 32.0005
R400 V_OUT.n411 V_OUT.n410 32.0005
R401 V_OUT.n410 V_OUT.n26 32.0005
R402 V_OUT.n406 V_OUT.n26 32.0005
R403 V_OUT.n406 V_OUT.n405 32.0005
R404 V_OUT.n405 V_OUT.n404 32.0005
R405 V_OUT.n404 V_OUT.n28 32.0005
R406 V_OUT.n398 V_OUT.n397 32.0005
R407 V_OUT.n397 V_OUT.n32 32.0005
R408 V_OUT.n393 V_OUT.n32 32.0005
R409 V_OUT.n393 V_OUT.n392 32.0005
R410 V_OUT.n392 V_OUT.n391 32.0005
R411 V_OUT.n391 V_OUT.n34 32.0005
R412 V_OUT.n387 V_OUT.n34 32.0005
R413 V_OUT.t152 V_OUT.t4 31.6345
R414 V_OUT.n312 V_OUT.n48 29.0291
R415 V_OUT.n330 V_OUT.n329 29.0291
R416 V_OUT.n179 V_OUT.n178 28.8005
R417 V_OUT.n161 V_OUT.n90 28.8005
R418 V_OUT.n224 V_OUT.n223 28.7587
R419 V_OUT.n461 V_OUT.n3 28.1154
R420 V_OUT.n271 V_OUT.n270 27.2005
R421 V_OUT.n276 V_OUT.n187 27.2005
R422 V_OUT.t43 V_OUT.t90 25.8829
R423 V_OUT.n329 V_OUT.n62 25.6005
R424 V_OUT.n346 V_OUT.n44 25.6005
R425 V_OUT.n353 V_OUT.n351 25.6005
R426 V_OUT.n222 V_OUT.n221 25.6005
R427 V_OUT.n217 V_OUT.n216 25.6005
R428 V_OUT.n239 V_OUT.n208 25.6005
R429 V_OUT.n230 V_OUT 25.6005
R430 V_OUT.n172 V_OUT.n171 25.6005
R431 V_OUT.n96 V_OUT.n94 25.6005
R432 V_OUT.n148 V_OUT.n97 25.6005
R433 V_OUT.n133 V_OUT.n103 25.6005
R434 V_OUT.n133 V_OUT.n132 25.6005
R435 V_OUT.n458 V_OUT.n4 25.6005
R436 V_OUT.n439 V_OUT.n438 25.6005
R437 V_OUT.n428 V_OUT.n17 25.6005
R438 V_OUT.n421 V_OUT.n21 25.6005
R439 V_OUT.n25 V_OUT.n23 25.6005
R440 V_OUT.n400 V_OUT.n30 25.6005
R441 V_OUT.n267 V_OUT.n266 24.8279
R442 V_OUT.n226 V_OUT.n225 24.8279
R443 V_OUT.n67 V_OUT.t63 24.6255
R444 V_OUT.n67 V_OUT.t55 24.6255
R445 V_OUT.n68 V_OUT.t0 24.6255
R446 V_OUT.n68 V_OUT.t70 24.6255
R447 V_OUT.n193 V_OUT.t140 24.0005
R448 V_OUT.n193 V_OUT.t5 24.0005
R449 V_OUT.n197 V_OUT.t147 24.0005
R450 V_OUT.n197 V_OUT.t91 24.0005
R451 V_OUT.n201 V_OUT.t62 24.0005
R452 V_OUT.n201 V_OUT.t17 24.0005
R453 V_OUT.n205 V_OUT.t39 24.0005
R454 V_OUT.n205 V_OUT.t50 24.0005
R455 V_OUT.n210 V_OUT.t48 24.0005
R456 V_OUT.n210 V_OUT.t132 24.0005
R457 V_OUT.n400 V_OUT.n399 22.4005
R458 V_OUT.n290 V_OUT.n289 20.9665
R459 V_OUT.n73 V_OUT.n69 19.2005
R460 V_OUT.n325 V_OUT.n324 19.2005
R461 V_OUT.n324 V_OUT.n323 19.2005
R462 V_OUT.n156 V_OUT.n92 19.2005
R463 V_OUT.t156 V_OUT.t96 17.8306
R464 V_OUT.n215 V_OUT.t16 17.2554
R465 V_OUT.n426 V_OUT.n19 16.0005
R466 V_OUT.n423 V_OUT.n19 16.0005
R467 V_OUT.n228 V_OUT 15.7005
R468 V_OUT.n289 V_OUT.n288 15.6449
R469 V_OUT.n359 V_OUT.n358 15.6449
R470 V_OUT.t14 V_OUT.n74 15.0005
R471 V_OUT.n74 V_OUT.t31 15.0005
R472 V_OUT.t31 V_OUT.n64 15.0005
R473 V_OUT.n64 V_OUT.t112 15.0005
R474 V_OUT.t143 V_OUT.n75 15.0005
R475 V_OUT.n75 V_OUT.t14 15.0005
R476 V_OUT.n304 V_OUT.t126 15.0005
R477 V_OUT.n304 V_OUT.t12 15.0005
R478 V_OUT.n307 V_OUT.t45 15.0005
R479 V_OUT.n307 V_OUT.t106 15.0005
R480 V_OUT.n345 V_OUT.t120 15.0005
R481 V_OUT.n345 V_OUT.t89 15.0005
R482 V_OUT.n352 V_OUT.t67 15.0005
R483 V_OUT.n352 V_OUT.t102 15.0005
R484 V_OUT.t120 V_OUT.n344 15.0005
R485 V_OUT.n336 V_OUT.t107 15.0005
R486 V_OUT.t126 V_OUT.n303 15.0005
R487 V_OUT.n331 V_OUT.t113 15.0005
R488 V_OUT.n77 V_OUT.t143 15.0005
R489 V_OUT.n41 V_OUT.t103 15.0005
R490 V_OUT.n358 V_OUT.n357 14.4005
R491 V_OUT.n272 V_OUT.n271 14.0805
R492 V_OUT.n274 V_OUT.n187 14.0805
R493 V_OUT.n460 V_OUT.n4 13.9181
R494 V_OUT.t47 V_OUT.t156 13.8044
R495 V_OUT.n228 V_OUT.n2 13.1958
R496 V_OUT.n183 V_OUT.n2 12.8163
R497 V_OUT.n329 V_OUT.n61 12.8005
R498 V_OUT.n292 V_OUT.n291 12.8005
R499 V_OUT.n346 V_OUT.n46 12.8005
R500 V_OUT.n353 V_OUT.n42 12.8005
R501 V_OUT.n221 V_OUT.n220 12.8005
R502 V_OUT.n218 V_OUT.n217 12.8005
R503 V_OUT.n159 V_OUT.n92 12.8005
R504 V_OUT.n108 V_OUT 12.7806
R505 V_OUT V_OUT.n35 11.8876
R506 V_OUT.n461 V_OUT.n460 11.7212
R507 V_OUT.n463 V_OUT.n462 11.6542
R508 V_OUT.n72 V_OUT.n71 9.91717
R509 V_OUT.n399 V_OUT.n398 9.6005
R510 V_OUT.n266 V_OUT.n265 9.58175
R511 V_OUT.n234 V_OUT.n226 9.58175
R512 V_OUT.n264 V_OUT.n263 9.3005
R513 V_OUT.n262 V_OUT.n191 9.3005
R514 V_OUT.n261 V_OUT.n260 9.3005
R515 V_OUT.n259 V_OUT.n192 9.3005
R516 V_OUT.n258 V_OUT.n257 9.3005
R517 V_OUT.n256 V_OUT.n195 9.3005
R518 V_OUT.n255 V_OUT.n254 9.3005
R519 V_OUT.n253 V_OUT.n196 9.3005
R520 V_OUT.n252 V_OUT.n251 9.3005
R521 V_OUT.n250 V_OUT.n199 9.3005
R522 V_OUT.n249 V_OUT.n248 9.3005
R523 V_OUT.n247 V_OUT.n200 9.3005
R524 V_OUT.n246 V_OUT.n245 9.3005
R525 V_OUT.n244 V_OUT.n203 9.3005
R526 V_OUT.n243 V_OUT.n242 9.3005
R527 V_OUT.n241 V_OUT.n204 9.3005
R528 V_OUT.n240 V_OUT.n239 9.3005
R529 V_OUT.n238 V_OUT.n207 9.3005
R530 V_OUT.n237 V_OUT.n236 9.3005
R531 V_OUT.n235 V_OUT.n209 9.3005
R532 V_OUT.n233 V_OUT.n232 9.3005
R533 V_OUT.n231 V_OUT.n227 9.3005
R534 V_OUT.n230 V_OUT.n229 9.3005
R535 V_OUT.n134 V_OUT.n133 9.3005
R536 V_OUT.n121 V_OUT.n120 9.3005
R537 V_OUT.n122 V_OUT.n107 9.3005
R538 V_OUT.n124 V_OUT.n123 9.3005
R539 V_OUT.n125 V_OUT.n106 9.3005
R540 V_OUT.n127 V_OUT.n126 9.3005
R541 V_OUT.n128 V_OUT.n105 9.3005
R542 V_OUT.n130 V_OUT.n129 9.3005
R543 V_OUT.n131 V_OUT.n102 9.3005
R544 V_OUT.n135 V_OUT.n101 9.3005
R545 V_OUT.n137 V_OUT.n136 9.3005
R546 V_OUT.n138 V_OUT.n100 9.3005
R547 V_OUT.n140 V_OUT.n139 9.3005
R548 V_OUT.n141 V_OUT.n99 9.3005
R549 V_OUT.n143 V_OUT.n142 9.3005
R550 V_OUT.n144 V_OUT.n98 9.3005
R551 V_OUT.n146 V_OUT.n145 9.3005
R552 V_OUT.n148 V_OUT.n147 9.3005
R553 V_OUT.n149 V_OUT.n95 9.3005
R554 V_OUT.n151 V_OUT.n150 9.3005
R555 V_OUT.n152 V_OUT.n94 9.3005
R556 V_OUT.n154 V_OUT.n153 9.3005
R557 V_OUT.n155 V_OUT.n93 9.3005
R558 V_OUT.n157 V_OUT.n156 9.3005
R559 V_OUT.n159 V_OUT.n158 9.3005
R560 V_OUT.n160 V_OUT.n91 9.3005
R561 V_OUT.n162 V_OUT.n161 9.3005
R562 V_OUT.n164 V_OUT.n163 9.3005
R563 V_OUT.n165 V_OUT.n88 9.3005
R564 V_OUT.n167 V_OUT.n166 9.3005
R565 V_OUT.n168 V_OUT.n87 9.3005
R566 V_OUT.n170 V_OUT.n169 9.3005
R567 V_OUT.n172 V_OUT.n83 9.3005
R568 V_OUT.n174 V_OUT.n173 9.3005
R569 V_OUT.n175 V_OUT.n82 9.3005
R570 V_OUT.n177 V_OUT.n176 9.3005
R571 V_OUT.n179 V_OUT.n80 9.3005
R572 V_OUT.n181 V_OUT.n180 9.3005
R573 V_OUT.n182 V_OUT.n79 9.3005
R574 V_OUT.n459 V_OUT.n458 9.3005
R575 V_OUT.n457 V_OUT.n5 9.3005
R576 V_OUT.n456 V_OUT.n455 9.3005
R577 V_OUT.n454 V_OUT.n6 9.3005
R578 V_OUT.n453 V_OUT.n452 9.3005
R579 V_OUT.n451 V_OUT.n7 9.3005
R580 V_OUT.n450 V_OUT.n449 9.3005
R581 V_OUT.n448 V_OUT.n9 9.3005
R582 V_OUT.n447 V_OUT.n446 9.3005
R583 V_OUT.n445 V_OUT.n10 9.3005
R584 V_OUT.n444 V_OUT.n443 9.3005
R585 V_OUT.n442 V_OUT.n11 9.3005
R586 V_OUT.n441 V_OUT.n440 9.3005
R587 V_OUT.n439 V_OUT.n13 9.3005
R588 V_OUT.n437 V_OUT.n436 9.3005
R589 V_OUT.n435 V_OUT.n15 9.3005
R590 V_OUT.n434 V_OUT.n433 9.3005
R591 V_OUT.n432 V_OUT.n16 9.3005
R592 V_OUT.n431 V_OUT.n430 9.3005
R593 V_OUT.n429 V_OUT.n428 9.3005
R594 V_OUT.n427 V_OUT.n18 9.3005
R595 V_OUT.n426 V_OUT.n425 9.3005
R596 V_OUT.n424 V_OUT.n423 9.3005
R597 V_OUT.n422 V_OUT.n20 9.3005
R598 V_OUT.n421 V_OUT.n420 9.3005
R599 V_OUT.n419 V_OUT.n418 9.3005
R600 V_OUT.n417 V_OUT.n22 9.3005
R601 V_OUT.n416 V_OUT.n415 9.3005
R602 V_OUT.n414 V_OUT.n23 9.3005
R603 V_OUT.n413 V_OUT.n412 9.3005
R604 V_OUT.n411 V_OUT.n24 9.3005
R605 V_OUT.n410 V_OUT.n409 9.3005
R606 V_OUT.n408 V_OUT.n26 9.3005
R607 V_OUT.n407 V_OUT.n406 9.3005
R608 V_OUT.n405 V_OUT.n27 9.3005
R609 V_OUT.n404 V_OUT.n403 9.3005
R610 V_OUT.n402 V_OUT.n28 9.3005
R611 V_OUT.n401 V_OUT.n400 9.3005
R612 V_OUT.n398 V_OUT.n29 9.3005
R613 V_OUT.n397 V_OUT.n396 9.3005
R614 V_OUT.n395 V_OUT.n32 9.3005
R615 V_OUT.n394 V_OUT.n393 9.3005
R616 V_OUT.n392 V_OUT.n33 9.3005
R617 V_OUT.n391 V_OUT.n390 9.3005
R618 V_OUT.n389 V_OUT.n34 9.3005
R619 V_OUT.n388 V_OUT.n387 9.3005
R620 V_OUT.n1 V_OUT.n0 9.3005
R621 V_OUT.n357 V_OUT.n356 9.3005
R622 V_OUT.n355 V_OUT.n42 9.3005
R623 V_OUT.n354 V_OUT.n353 9.3005
R624 V_OUT.n351 V_OUT.n43 9.3005
R625 V_OUT.n350 V_OUT.n349 9.3005
R626 V_OUT.n348 V_OUT.n44 9.3005
R627 V_OUT.n347 V_OUT.n346 9.3005
R628 V_OUT.n46 V_OUT.n45 9.3005
R629 V_OUT.n311 V_OUT.n310 9.3005
R630 V_OUT.n312 V_OUT.n309 9.3005
R631 V_OUT.n292 V_OUT.n66 9.3005
R632 V_OUT.n294 V_OUT.n293 9.3005
R633 V_OUT.n295 V_OUT.n65 9.3005
R634 V_OUT.n297 V_OUT.n296 9.3005
R635 V_OUT.n298 V_OUT.n63 9.3005
R636 V_OUT.n300 V_OUT.n299 9.3005
R637 V_OUT.n301 V_OUT.n61 9.3005
R638 V_OUT.n329 V_OUT.n328 9.3005
R639 V_OUT.n327 V_OUT.n62 9.3005
R640 V_OUT.n326 V_OUT.n325 9.3005
R641 V_OUT.n324 V_OUT.n302 9.3005
R642 V_OUT.n323 V_OUT.n322 9.3005
R643 V_OUT.n321 V_OUT.n305 9.3005
R644 V_OUT.n320 V_OUT.n319 9.3005
R645 V_OUT.n318 V_OUT.n306 9.3005
R646 V_OUT.n317 V_OUT.n316 9.3005
R647 V_OUT.n315 V_OUT.n308 9.3005
R648 V_OUT.n314 V_OUT.n313 9.3005
R649 V_OUT.t146 V_OUT.t145 8.62795
R650 V_OUT.t115 V_OUT.t131 8.62795
R651 V_OUT.n71 V_OUT.t109 8.246
R652 V_OUT.n184 V_OUT.n183 7.49888
R653 V_OUT.n284 V_OUT.n283 7.11161
R654 V_OUT.n288 V_OUT.n76 7.11161
R655 V_OUT.n364 V_OUT.n363 7.11161
R656 V_OUT.n361 V_OUT.n359 7.11161
R657 V_OUT.n291 V_OUT.n290 6.69883
R658 V_OUT.n298 V_OUT.n297 6.4005
R659 V_OUT.n318 V_OUT.n317 6.4005
R660 V_OUT.n313 V_OUT.n312 6.4005
R661 V_OUT.n208 V_OUT.n204 6.4005
R662 V_OUT.n171 V_OUT.n170 6.4005
R663 V_OUT.n150 V_OUT.n96 6.4005
R664 V_OUT.n145 V_OUT.n97 6.4005
R665 V_OUT.n103 V_OUT.n101 6.4005
R666 V_OUT.n132 V_OUT.n131 6.4005
R667 V_OUT.n120 V_OUT.n119 6.4005
R668 V_OUT.n438 V_OUT.n437 6.4005
R669 V_OUT.n431 V_OUT.n17 6.4005
R670 V_OUT.n418 V_OUT.n21 6.4005
R671 V_OUT.n412 V_OUT.n25 6.4005
R672 V_OUT.n30 V_OUT.n28 6.4005
R673 V_OUT.n387 V_OUT.n386 6.4005
R674 V_OUT.n357 V_OUT.n1 6.4005
R675 V_OUT.n116 V_OUT.n115 5.68939
R676 V_OUT.n116 V_OUT.n104 5.68939
R677 V_OUT.n368 V_OUT.n367 5.68939
R678 V_OUT.n71 V_OUT.n3 5.22371
R679 V_OUT.n368 V_OUT.n31 4.97828
R680 V_OUT.n283 V_OUT.n282 3.48951
R681 V_OUT.n282 V_OUT.n76 3.48951
R682 V_OUT.n363 V_OUT.n362 3.48951
R683 V_OUT.n362 V_OUT.n361 3.48951
R684 V_OUT.n178 V_OUT.n177 3.2005
R685 V_OUT.n164 V_OUT.n90 3.2005
R686 V_OUT.t139 V_OUT.t40 2.87632
R687 V_OUT.t92 V_OUT.t49 2.87632
R688 V_OUT.n50 V_OUT.n47 2.25882
R689 V_OUT.n50 V_OUT.n49 2.25882
R690 V_OUT.n343 V_OUT.n48 2.25882
R691 V_OUT.n342 V_OUT.n49 2.25882
R692 V_OUT.n337 V_OUT.n47 2.25882
R693 V_OUT.n343 V_OUT.n342 2.25882
R694 V_OUT.n56 V_OUT.n55 2.25882
R695 V_OUT.n57 V_OUT.n56 2.25882
R696 V_OUT.n330 V_OUT.n60 2.25882
R697 V_OUT.n59 V_OUT.n57 2.25882
R698 V_OUT.n332 V_OUT.n55 2.25882
R699 V_OUT.n60 V_OUT.n59 2.25882
R700 V_OUT.n462 V_OUT.n2 0.9875
R701 V_OUT.n290 V_OUT.n66 0.703977
R702 V_OUT.n183 V_OUT.n182 0.193977
R703 V_OUT.n121 V_OUT.n108 0.193881
R704 V_OUT.n388 V_OUT.n35 0.193881
R705 V_OUT.n460 V_OUT.n459 0.193695
R706 V_OUT.n229 V_OUT.n228 0.188
R707 V_OUT.n264 V_OUT.n191 0.15675
R708 V_OUT.n260 V_OUT.n259 0.15675
R709 V_OUT.n259 V_OUT.n258 0.15675
R710 V_OUT.n258 V_OUT.n195 0.15675
R711 V_OUT.n254 V_OUT.n253 0.15675
R712 V_OUT.n253 V_OUT.n252 0.15675
R713 V_OUT.n252 V_OUT.n199 0.15675
R714 V_OUT.n248 V_OUT.n247 0.15675
R715 V_OUT.n247 V_OUT.n246 0.15675
R716 V_OUT.n246 V_OUT.n203 0.15675
R717 V_OUT.n242 V_OUT.n241 0.15675
R718 V_OUT.n241 V_OUT.n240 0.15675
R719 V_OUT.n240 V_OUT.n207 0.15675
R720 V_OUT.n236 V_OUT.n235 0.15675
R721 V_OUT.n233 V_OUT.n227 0.15675
R722 V_OUT.n229 V_OUT.n227 0.15675
R723 V_OUT.n182 V_OUT.n181 0.15675
R724 V_OUT.n181 V_OUT.n80 0.15675
R725 V_OUT.n176 V_OUT.n80 0.15675
R726 V_OUT.n176 V_OUT.n175 0.15675
R727 V_OUT.n175 V_OUT.n174 0.15675
R728 V_OUT.n174 V_OUT.n83 0.15675
R729 V_OUT.n169 V_OUT.n83 0.15675
R730 V_OUT.n169 V_OUT.n168 0.15675
R731 V_OUT.n168 V_OUT.n167 0.15675
R732 V_OUT.n167 V_OUT.n88 0.15675
R733 V_OUT.n163 V_OUT.n88 0.15675
R734 V_OUT.n163 V_OUT.n162 0.15675
R735 V_OUT.n162 V_OUT.n91 0.15675
R736 V_OUT.n158 V_OUT.n91 0.15675
R737 V_OUT.n158 V_OUT.n157 0.15675
R738 V_OUT.n157 V_OUT.n93 0.15675
R739 V_OUT.n153 V_OUT.n93 0.15675
R740 V_OUT.n153 V_OUT.n152 0.15675
R741 V_OUT.n152 V_OUT.n151 0.15675
R742 V_OUT.n151 V_OUT.n95 0.15675
R743 V_OUT.n147 V_OUT.n95 0.15675
R744 V_OUT.n147 V_OUT.n146 0.15675
R745 V_OUT.n146 V_OUT.n98 0.15675
R746 V_OUT.n142 V_OUT.n98 0.15675
R747 V_OUT.n142 V_OUT.n141 0.15675
R748 V_OUT.n141 V_OUT.n140 0.15675
R749 V_OUT.n140 V_OUT.n100 0.15675
R750 V_OUT.n136 V_OUT.n100 0.15675
R751 V_OUT.n136 V_OUT.n135 0.15675
R752 V_OUT.n135 V_OUT.n134 0.15675
R753 V_OUT.n134 V_OUT.n102 0.15675
R754 V_OUT.n129 V_OUT.n102 0.15675
R755 V_OUT.n129 V_OUT.n128 0.15675
R756 V_OUT.n128 V_OUT.n127 0.15675
R757 V_OUT.n127 V_OUT.n106 0.15675
R758 V_OUT.n123 V_OUT.n106 0.15675
R759 V_OUT.n123 V_OUT.n122 0.15675
R760 V_OUT.n122 V_OUT.n121 0.15675
R761 V_OUT.n459 V_OUT.n5 0.15675
R762 V_OUT.n455 V_OUT.n5 0.15675
R763 V_OUT.n455 V_OUT.n454 0.15675
R764 V_OUT.n454 V_OUT.n453 0.15675
R765 V_OUT.n453 V_OUT.n7 0.15675
R766 V_OUT.n449 V_OUT.n7 0.15675
R767 V_OUT.n449 V_OUT.n448 0.15675
R768 V_OUT.n448 V_OUT.n447 0.15675
R769 V_OUT.n447 V_OUT.n10 0.15675
R770 V_OUT.n443 V_OUT.n442 0.15675
R771 V_OUT.n442 V_OUT.n441 0.15675
R772 V_OUT.n441 V_OUT.n13 0.15675
R773 V_OUT.n436 V_OUT.n13 0.15675
R774 V_OUT.n436 V_OUT.n435 0.15675
R775 V_OUT.n435 V_OUT.n434 0.15675
R776 V_OUT.n434 V_OUT.n16 0.15675
R777 V_OUT.n430 V_OUT.n16 0.15675
R778 V_OUT.n430 V_OUT.n429 0.15675
R779 V_OUT.n429 V_OUT.n18 0.15675
R780 V_OUT.n425 V_OUT.n18 0.15675
R781 V_OUT.n425 V_OUT.n424 0.15675
R782 V_OUT.n424 V_OUT.n20 0.15675
R783 V_OUT.n420 V_OUT.n20 0.15675
R784 V_OUT.n420 V_OUT.n419 0.15675
R785 V_OUT.n419 V_OUT.n22 0.15675
R786 V_OUT.n415 V_OUT.n22 0.15675
R787 V_OUT.n415 V_OUT.n414 0.15675
R788 V_OUT.n414 V_OUT.n413 0.15675
R789 V_OUT.n413 V_OUT.n24 0.15675
R790 V_OUT.n409 V_OUT.n24 0.15675
R791 V_OUT.n409 V_OUT.n408 0.15675
R792 V_OUT.n408 V_OUT.n407 0.15675
R793 V_OUT.n407 V_OUT.n27 0.15675
R794 V_OUT.n403 V_OUT.n27 0.15675
R795 V_OUT.n403 V_OUT.n402 0.15675
R796 V_OUT.n402 V_OUT.n401 0.15675
R797 V_OUT.n401 V_OUT.n29 0.15675
R798 V_OUT.n396 V_OUT.n29 0.15675
R799 V_OUT.n396 V_OUT.n395 0.15675
R800 V_OUT.n395 V_OUT.n394 0.15675
R801 V_OUT.n394 V_OUT.n33 0.15675
R802 V_OUT.n390 V_OUT.n33 0.15675
R803 V_OUT.n390 V_OUT.n389 0.15675
R804 V_OUT.n389 V_OUT.n388 0.15675
R805 V_OUT.n294 V_OUT.n66 0.15675
R806 V_OUT.n295 V_OUT.n294 0.15675
R807 V_OUT.n296 V_OUT.n295 0.15675
R808 V_OUT.n296 V_OUT.n63 0.15675
R809 V_OUT.n300 V_OUT.n63 0.15675
R810 V_OUT.n301 V_OUT.n300 0.15675
R811 V_OUT.n328 V_OUT.n301 0.15675
R812 V_OUT.n328 V_OUT.n327 0.15675
R813 V_OUT.n327 V_OUT.n326 0.15675
R814 V_OUT.n326 V_OUT.n302 0.15675
R815 V_OUT.n322 V_OUT.n302 0.15675
R816 V_OUT.n322 V_OUT.n321 0.15675
R817 V_OUT.n321 V_OUT.n320 0.15675
R818 V_OUT.n320 V_OUT.n306 0.15675
R819 V_OUT.n316 V_OUT.n306 0.15675
R820 V_OUT.n316 V_OUT.n315 0.15675
R821 V_OUT.n315 V_OUT.n314 0.15675
R822 V_OUT.n314 V_OUT.n309 0.15675
R823 V_OUT.n310 V_OUT.n309 0.15675
R824 V_OUT.n310 V_OUT.n45 0.15675
R825 V_OUT.n347 V_OUT.n45 0.15675
R826 V_OUT.n348 V_OUT.n347 0.15675
R827 V_OUT.n349 V_OUT.n348 0.15675
R828 V_OUT.n349 V_OUT.n43 0.15675
R829 V_OUT.n354 V_OUT.n43 0.15675
R830 V_OUT.n355 V_OUT.n354 0.15675
R831 V_OUT.n356 V_OUT.n355 0.15675
R832 V_OUT.n356 V_OUT.n0 0.15675
R833 V_OUT.n462 V_OUT.n461 0.1321
R834 V_OUT.n265 V_OUT.n188 0.131895
R835 V_OUT V_OUT.n0 0.1255
R836 V_OUT.n12 V_OUT.n10 0.109875
R837 V_OUT.n194 V_OUT.n191 0.09425
R838 V_OUT.n198 V_OUT.n195 0.09425
R839 V_OUT.n202 V_OUT.n199 0.09425
R840 V_OUT.n206 V_OUT.n203 0.09425
R841 V_OUT.n211 V_OUT.n207 0.09425
R842 V_OUT.n235 V_OUT.n234 0.09425
R843 V_OUT.n72 V_OUT.n70 0.0838333
R844 V_OUT.n72 V_OUT 0.063
R845 V_OUT.n265 V_OUT.n264 0.063
R846 V_OUT.n260 V_OUT.n194 0.063
R847 V_OUT.n254 V_OUT.n198 0.063
R848 V_OUT.n248 V_OUT.n202 0.063
R849 V_OUT.n242 V_OUT.n206 0.063
R850 V_OUT.n236 V_OUT.n211 0.063
R851 V_OUT.n234 V_OUT.n233 0.063
R852 V_OUT V_OUT.n463 0.063
R853 V_OUT.n443 V_OUT.n12 0.047375
R854 a_5970_4630.n8 a_5970_4630.n6 522.322
R855 a_5970_4630.n3 a_5970_4630.t3 384.967
R856 a_5970_4630.n0 a_5970_4630.t6 384.967
R857 a_5970_4630.n3 a_5970_4630.t5 379.166
R858 a_5970_4630.t7 a_5970_4630.n0 376.56
R859 a_5970_4630.n5 a_5970_4630.n1 315.647
R860 a_5970_4630.n4 a_5970_4630.n2 315.647
R861 a_5970_4630.n11 a_5970_4630.n10 314.502
R862 a_5970_4630.n8 a_5970_4630.n7 160.721
R863 a_5970_4630.n5 a_5970_4630.n4 83.2005
R864 a_5970_4630.n1 a_5970_4630.t11 49.2505
R865 a_5970_4630.n1 a_5970_4630.t10 49.2505
R866 a_5970_4630.n2 a_5970_4630.t9 49.2505
R867 a_5970_4630.n2 a_5970_4630.t4 49.2505
R868 a_5970_4630.t7 a_5970_4630.n11 49.2505
R869 a_5970_4630.n11 a_5970_4630.t12 49.2505
R870 a_5970_4630.n10 a_5970_4630.n9 42.6672
R871 a_5970_4630.n9 a_5970_4630.n8 37.763
R872 a_5970_4630.n9 a_5970_4630.n5 23.4672
R873 a_5970_4630.n6 a_5970_4630.t2 19.7005
R874 a_5970_4630.n6 a_5970_4630.t1 19.7005
R875 a_5970_4630.n7 a_5970_4630.t0 19.7005
R876 a_5970_4630.n7 a_5970_4630.t8 19.7005
R877 a_5970_4630.n4 a_5970_4630.n3 16.0005
R878 a_5970_4630.n10 a_5970_4630.n0 16.0005
R879 VDDA.n468 VDDA.n460 831.25
R880 VDDA.n463 VDDA.n462 831.25
R881 VDDA.n457 VDDA.n449 831.25
R882 VDDA.n452 VDDA.n451 831.25
R883 VDDA.n461 VDDA.n460 585
R884 VDDA.n465 VDDA.n463 585
R885 VDDA.n361 VDDA.n355 585
R886 VDDA.n356 VDDA.n355 585
R887 VDDA.n367 VDDA.n44 585
R888 VDDA.n371 VDDA.n44 585
R889 VDDA.n312 VDDA.n50 585
R890 VDDA.n307 VDDA.n50 585
R891 VDDA.n288 VDDA.n283 585
R892 VDDA.n292 VDDA.n283 585
R893 VDDA.n450 VDDA.n449 585
R894 VDDA.n454 VDDA.n452 585
R895 VDDA.n352 VDDA.n346 585
R896 VDDA.n347 VDDA.n346 585
R897 VDDA.n58 VDDA.n51 585
R898 VDDA.n53 VDDA.n51 585
R899 VDDA.n123 VDDA.n116 585
R900 VDDA.n105 VDDA.n97 585
R901 VDDA.n271 VDDA.n175 585
R902 VDDA.n264 VDDA.n175 585
R903 VDDA.n261 VDDA.n260 585
R904 VDDA.n260 VDDA.n259 585
R905 VDDA.n230 VDDA.n229 585
R906 VDDA.n230 VDDA.n219 585
R907 VDDA.n467 VDDA.t10 465.079
R908 VDDA.t10 VDDA.n466 465.079
R909 VDDA.n456 VDDA.t18 465.079
R910 VDDA.t18 VDDA.n455 465.079
R911 VDDA.t110 VDDA.n336 464.281
R912 VDDA.n338 VDDA.t110 464.281
R913 VDDA.n444 VDDA.t97 464.281
R914 VDDA.t97 VDDA.n443 464.281
R915 VDDA.n481 VDDA.t21 464.281
R916 VDDA.t21 VDDA.n480 464.281
R917 VDDA.n425 VDDA.t87 464.281
R918 VDDA.t87 VDDA.n424 464.281
R919 VDDA.n403 VDDA.t107 464.281
R920 VDDA.t107 VDDA.n402 464.281
R921 VDDA.n333 VDDA.t25 464.281
R922 VDDA.t25 VDDA.n332 464.281
R923 VDDA.t111 VDDA.n433 464.281
R924 VDDA.n434 VDDA.t111 464.281
R925 VDDA.t36 VDDA.n17 464.281
R926 VDDA.n471 VDDA.t36 464.281
R927 VDDA.t23 VDDA.n25 464.281
R928 VDDA.n406 VDDA.t23 464.281
R929 VDDA.t128 VDDA.n321 464.281
R930 VDDA.n322 VDDA.t128 464.281
R931 VDDA.n41 VDDA.t130 415.336
R932 VDDA.n86 VDDA.t61 384.967
R933 VDDA.n128 VDDA.t67 384.967
R934 VDDA.n91 VDDA.t46 384.967
R935 VDDA.n111 VDDA.t43 384.967
R936 VDDA.n123 VDDA.t54 374.878
R937 VDDA.t65 VDDA.t82 360.346
R938 VDDA.t82 VDDA.t39 360.346
R939 VDDA.t39 VDDA.t2 360.346
R940 VDDA.t2 VDDA.t100 360.346
R941 VDDA.t100 VDDA.t58 360.346
R942 VDDA.t0 VDDA.t72 360.346
R943 VDDA.t37 VDDA.t0 360.346
R944 VDDA.t7 VDDA.t37 360.346
R945 VDDA.t98 VDDA.t7 360.346
R946 VDDA.t75 VDDA.t98 360.346
R947 VDDA.n96 VDDA.t50 352.834
R948 VDDA.n225 VDDA.t65 343.966
R949 VDDA.n263 VDDA.t58 343.966
R950 VDDA.t72 VDDA.n263 343.966
R951 VDDA.n269 VDDA.t75 343.966
R952 VDDA.n112 VDDA.t45 341.752
R953 VDDA.n127 VDDA.t70 341.752
R954 VDDA.n87 VDDA.t63 341.752
R955 VDDA.n92 VDDA.t49 341.752
R956 VDDA.n258 VDDA.t71 336.329
R957 VDDA.n258 VDDA.t57 336.329
R958 VDDA.n220 VDDA.t64 320.7
R959 VDDA.n272 VDDA.t74 320.7
R960 VDDA.n85 VDDA.n83 315.647
R961 VDDA.n79 VDDA.n78 315.647
R962 VDDA.n110 VDDA.n109 315.647
R963 VDDA.n90 VDDA.n89 315.647
R964 VDDA.n130 VDDA.n82 315.647
R965 VDDA.n129 VDDA.n84 315.647
R966 VDDA.n24 VDDA.t120 315.25
R967 VDDA.t112 VDDA.t6 314.113
R968 VDDA.t124 VDDA.t17 314.113
R969 VDDA.t62 VDDA.n87 304.659
R970 VDDA.n260 VDDA.n183 291.363
R971 VDDA.n256 VDDA.n181 291.363
R972 VDDA.n257 VDDA.n256 291.363
R973 VDDA.n359 VDDA.n355 290.733
R974 VDDA.n365 VDDA.n44 290.733
R975 VDDA.n310 VDDA.n50 290.733
R976 VDDA.n286 VDDA.n283 290.733
R977 VDDA.n350 VDDA.n346 290.733
R978 VDDA.n52 VDDA.n51 290.733
R979 VDDA.n121 VDDA.n116 290.733
R980 VDDA.n117 VDDA.n116 290.733
R981 VDDA.n103 VDDA.n97 290.733
R982 VDDA.n98 VDDA.n97 290.733
R983 VDDA.n265 VDDA.n175 290.733
R984 VDDA.n230 VDDA.n218 290.733
R985 VDDA.n445 VDDA.n444 243.698
R986 VDDA.n482 VDDA.n481 243.698
R987 VDDA.n426 VDDA.n425 243.698
R988 VDDA.n404 VDDA.n403 243.698
R989 VDDA.n334 VDDA.n333 243.698
R990 VDDA.n434 VDDA.n431 243.698
R991 VDDA.n475 VDDA.n471 243.698
R992 VDDA.n410 VDDA.n406 243.698
R993 VDDA.n322 VDDA.n319 243.698
R994 VDDA.n430 VDDA.n1 238.367
R995 VDDA.n469 VDDA.n468 238.367
R996 VDDA.n462 VDDA.n429 238.367
R997 VDDA.n428 VDDA.n16 238.367
R998 VDDA.n421 VDDA.n19 238.367
R999 VDDA.n399 VDDA.n27 238.367
R1000 VDDA.n318 VDDA.n35 238.367
R1001 VDDA.n438 VDDA.n2 238.367
R1002 VDDA.n458 VDDA.n457 238.367
R1003 VDDA.n485 VDDA.n484 238.367
R1004 VDDA.n413 VDDA.n412 238.367
R1005 VDDA.n326 VDDA.n31 238.367
R1006 VDDA.n451 VDDA.n447 238.367
R1007 VDDA.n117 VDDA.n88 233.841
R1008 VDDA.n98 VDDA.n94 233.841
R1009 VDDA.n362 VDDA.n361 230.308
R1010 VDDA.n356 VDDA.n315 230.308
R1011 VDDA.n368 VDDA.n367 230.308
R1012 VDDA.n371 VDDA.n370 230.308
R1013 VDDA.n313 VDDA.n312 230.308
R1014 VDDA.n307 VDDA.n46 230.308
R1015 VDDA.n289 VDDA.n288 230.308
R1016 VDDA.n292 VDDA.n291 230.308
R1017 VDDA.n353 VDDA.n352 230.308
R1018 VDDA.n58 VDDA.n48 230.308
R1019 VDDA.n53 VDDA.n47 230.308
R1020 VDDA.n347 VDDA.n344 230.308
R1021 VDDA.n124 VDDA.n123 230.308
R1022 VDDA.n271 VDDA.n270 230.308
R1023 VDDA.n268 VDDA.n264 230.308
R1024 VDDA.n262 VDDA.n261 230.308
R1025 VDDA.n259 VDDA.n178 230.308
R1026 VDDA.t19 VDDA.t30 222.178
R1027 VDDA.n363 VDDA.n343 199.195
R1028 VDDA.n192 VDDA.n191 196.502
R1029 VDDA.n189 VDDA.n188 196.502
R1030 VDDA.n255 VDDA.n254 196.502
R1031 VDDA.n246 VDDA.n211 196.502
R1032 VDDA.n239 VDDA.n214 196.502
R1033 VDDA.n232 VDDA.n231 196.502
R1034 VDDA.n338 VDDA.n317 190.333
R1035 VDDA.n127 VDDA.n126 185.001
R1036 VDDA.n113 VDDA.n112 185.001
R1037 VDDA.n108 VDDA.n92 185.001
R1038 VDDA.n57 VDDA.n56 185
R1039 VDDA.n55 VDDA.n54 185
R1040 VDDA.n351 VDDA.n345 185
R1041 VDDA.n349 VDDA.n348 185
R1042 VDDA.n325 VDDA.n324 185
R1043 VDDA.n323 VDDA.n320 185
R1044 VDDA.n407 VDDA.n26 185
R1045 VDDA.n409 VDDA.n408 185
R1046 VDDA.n472 VDDA.n18 185
R1047 VDDA.n474 VDDA.n473 185
R1048 VDDA.n450 VDDA.n448 185
R1049 VDDA.n454 VDDA.n453 185
R1050 VDDA.n437 VDDA.n436 185
R1051 VDDA.n435 VDDA.n432 185
R1052 VDDA.n287 VDDA.n285 185
R1053 VDDA.n284 VDDA.n282 185
R1054 VDDA.n311 VDDA.n49 185
R1055 VDDA.n309 VDDA.n308 185
R1056 VDDA.n366 VDDA.n364 185
R1057 VDDA.n45 VDDA.n43 185
R1058 VDDA.n360 VDDA.n354 185
R1059 VDDA.n358 VDDA.n357 185
R1060 VDDA.n329 VDDA.n328 185
R1061 VDDA.n331 VDDA.n330 185
R1062 VDDA.n29 VDDA.n28 185
R1063 VDDA.n401 VDDA.n400 185
R1064 VDDA.n21 VDDA.n20 185
R1065 VDDA.n423 VDDA.n422 185
R1066 VDDA.n477 VDDA.n476 185
R1067 VDDA.n479 VDDA.n478 185
R1068 VDDA.n461 VDDA.n459 185
R1069 VDDA.n465 VDDA.n464 185
R1070 VDDA.n440 VDDA.n439 185
R1071 VDDA.n442 VDDA.n441 185
R1072 VDDA.n342 VDDA.n34 185
R1073 VDDA.n343 VDDA.n342 185
R1074 VDDA.n341 VDDA.n340 185
R1075 VDDA.n339 VDDA.n337 185
R1076 VDDA.n343 VDDA.n317 185
R1077 VDDA.n122 VDDA.n115 185
R1078 VDDA.n120 VDDA.n114 185
R1079 VDDA.n125 VDDA.n114 185
R1080 VDDA.n119 VDDA.n118 185
R1081 VDDA.n106 VDDA.n105 185
R1082 VDDA.n107 VDDA.n106 185
R1083 VDDA.n104 VDDA.n95 185
R1084 VDDA.n102 VDDA.n101 185
R1085 VDDA.n100 VDDA.n99 185
R1086 VDDA.n182 VDDA.n179 185
R1087 VDDA.n185 VDDA.n184 185
R1088 VDDA.n177 VDDA.n176 185
R1089 VDDA.n267 VDDA.n266 185
R1090 VDDA.n229 VDDA.n221 185
R1091 VDDA.n225 VDDA.n221 185
R1092 VDDA.n228 VDDA.n227 185
R1093 VDDA.n223 VDDA.n222 185
R1094 VDDA.n224 VDDA.n219 185
R1095 VDDA.n225 VDDA.n224 185
R1096 VDDA.n290 VDDA.t19 172.38
R1097 VDDA.t115 VDDA.n314 172.38
R1098 VDDA.n369 VDDA.t113 172.38
R1099 VDDA.n259 VDDA.n258 166.63
R1100 VDDA.n441 VDDA.n439 150
R1101 VDDA.n464 VDDA.n459 150
R1102 VDDA.n478 VDDA.n476 150
R1103 VDDA.n422 VDDA.n20 150
R1104 VDDA.n400 VDDA.n28 150
R1105 VDDA.n330 VDDA.n328 150
R1106 VDDA.n437 VDDA.n432 150
R1107 VDDA.n453 VDDA.n448 150
R1108 VDDA.n474 VDDA.n18 150
R1109 VDDA.n409 VDDA.n26 150
R1110 VDDA.n325 VDDA.n320 150
R1111 VDDA.n342 VDDA.n341 150
R1112 VDDA.n337 VDDA.n317 150
R1113 VDDA.t32 VDDA.t84 145.038
R1114 VDDA.n335 VDDA.n327 137.904
R1115 VDDA.n411 VDDA.n405 137.904
R1116 VDDA.n290 VDDA.t121 126.412
R1117 VDDA.n314 VDDA.t30 126.412
R1118 VDDA.n369 VDDA.t115 126.412
R1119 VDDA.t113 VDDA.n363 126.412
R1120 VDDA.t123 VDDA.n460 123.126
R1121 VDDA.n463 VDDA.t123 123.126
R1122 VDDA.t27 VDDA.n449 123.126
R1123 VDDA.n452 VDDA.t27 123.126
R1124 VDDA.n357 VDDA.n354 120.001
R1125 VDDA.n364 VDDA.n45 120.001
R1126 VDDA.n308 VDDA.n49 120.001
R1127 VDDA.n285 VDDA.n284 120.001
R1128 VDDA.n348 VDDA.n345 120.001
R1129 VDDA.n56 VDDA.n55 120.001
R1130 VDDA.n115 VDDA.n114 120.001
R1131 VDDA.n118 VDDA.n114 120.001
R1132 VDDA.n106 VDDA.n95 120.001
R1133 VDDA.n101 VDDA.n100 120.001
R1134 VDDA.n267 VDDA.n177 120.001
R1135 VDDA.n184 VDDA.n179 120.001
R1136 VDDA.n227 VDDA.n221 120.001
R1137 VDDA.n224 VDDA.n223 120.001
R1138 VDDA.n161 VDDA.n67 119.737
R1139 VDDA.n154 VDDA.n70 119.737
R1140 VDDA.n147 VDDA.n73 119.737
R1141 VDDA.n140 VDDA.n76 119.737
R1142 VDDA.n132 VDDA.n81 119.737
R1143 VDDA.n126 VDDA.t68 119.656
R1144 VDDA.n125 VDDA.n113 108.779
R1145 VDDA.n483 VDDA.n427 107.258
R1146 VDDA.n483 VDDA.t20 103.427
R1147 VDDA.t9 VDDA.n470 103.427
R1148 VDDA.n470 VDDA.t26 103.427
R1149 VDDA.t96 VDDA.n446 103.427
R1150 VDDA.n427 VDDA.t22 95.7666
R1151 VDDA.t92 VDDA.t62 94.2753
R1152 VDDA.t90 VDDA.t92 94.2753
R1153 VDDA.t88 VDDA.t90 94.2753
R1154 VDDA.t94 VDDA.t88 94.2753
R1155 VDDA.t68 VDDA.t94 94.2753
R1156 VDDA.t80 VDDA.t104 94.2753
R1157 VDDA.t102 VDDA.t47 94.2753
R1158 VDDA.t28 VDDA.n108 94.2753
R1159 VDDA.t35 VDDA.t126 94.2753
R1160 VDDA.t117 VDDA.t116 94.2753
R1161 VDDA.t24 VDDA.t109 91.936
R1162 VDDA.t106 VDDA.t127 91.936
R1163 VDDA.t119 VDDA.t86 84.2747
R1164 VDDA.t20 VDDA.t112 84.2747
R1165 VDDA.t6 VDDA.t9 84.2747
R1166 VDDA.t26 VDDA.t124 84.2747
R1167 VDDA.t17 VDDA.t96 84.2747
R1168 VDDA.t55 VDDA.t44 83.3974
R1169 VDDA.t11 VDDA.t125 83.3974
R1170 VDDA.n110 VDDA.n79 83.2005
R1171 VDDA.n90 VDDA.n79 83.2005
R1172 VDDA.n130 VDDA.n83 83.2005
R1173 VDDA.n130 VDDA.n129 83.2005
R1174 VDDA.t13 VDDA.t41 76.1455
R1175 VDDA.t51 VDDA.t34 76.1455
R1176 VDDA.n314 VDDA.n48 69.8479
R1177 VDDA.n314 VDDA.n47 69.8479
R1178 VDDA.n363 VDDA.n353 69.8479
R1179 VDDA.n363 VDDA.n344 69.8479
R1180 VDDA.n290 VDDA.n289 69.8479
R1181 VDDA.n291 VDDA.n290 69.8479
R1182 VDDA.n314 VDDA.n313 69.8479
R1183 VDDA.n314 VDDA.n46 69.8479
R1184 VDDA.n369 VDDA.n368 69.8479
R1185 VDDA.n370 VDDA.n369 69.8479
R1186 VDDA.n363 VDDA.n362 69.8479
R1187 VDDA.n363 VDDA.n315 69.8479
R1188 VDDA.n125 VDDA.n124 69.8479
R1189 VDDA.n125 VDDA.n88 69.8479
R1190 VDDA.n107 VDDA.n93 69.8479
R1191 VDDA.n107 VDDA.n94 69.8479
R1192 VDDA.n263 VDDA.n262 69.8479
R1193 VDDA.n263 VDDA.n178 69.8479
R1194 VDDA.n270 VDDA.n269 69.8479
R1195 VDDA.n269 VDDA.n268 69.8479
R1196 VDDA.n226 VDDA.n225 69.8479
R1197 VDDA.n131 VDDA.n130 69.3203
R1198 VDDA.t41 VDDA.t4 68.8936
R1199 VDDA.t34 VDDA.n107 68.8936
R1200 VDDA.n327 VDDA.n326 65.8183
R1201 VDDA.n327 VDDA.n319 65.8183
R1202 VDDA.n412 VDDA.n411 65.8183
R1203 VDDA.n411 VDDA.n410 65.8183
R1204 VDDA.n484 VDDA.n483 65.8183
R1205 VDDA.n483 VDDA.n475 65.8183
R1206 VDDA.n470 VDDA.n458 65.8183
R1207 VDDA.n470 VDDA.n447 65.8183
R1208 VDDA.n446 VDDA.n438 65.8183
R1209 VDDA.n446 VDDA.n431 65.8183
R1210 VDDA.n335 VDDA.n334 65.8183
R1211 VDDA.n335 VDDA.n318 65.8183
R1212 VDDA.n405 VDDA.n404 65.8183
R1213 VDDA.n405 VDDA.n27 65.8183
R1214 VDDA.n427 VDDA.n426 65.8183
R1215 VDDA.n427 VDDA.n19 65.8183
R1216 VDDA.n483 VDDA.n482 65.8183
R1217 VDDA.n483 VDDA.n428 65.8183
R1218 VDDA.n470 VDDA.n469 65.8183
R1219 VDDA.n470 VDDA.n429 65.8183
R1220 VDDA.n446 VDDA.n445 65.8183
R1221 VDDA.n446 VDDA.n430 65.8183
R1222 VDDA.n343 VDDA.n316 65.8183
R1223 VDDA.t44 VDDA.t15 61.6417
R1224 VDDA.t125 VDDA.t78 61.6417
R1225 VDDA.n516 VDDA.n1 58.0576
R1226 VDDA.n486 VDDA.n16 58.0576
R1227 VDDA.n421 VDDA.n420 58.0576
R1228 VDDA.n399 VDDA.n398 58.0576
R1229 VDDA.n389 VDDA.n35 58.0576
R1230 VDDA.n516 VDDA.n2 58.0576
R1231 VDDA.n486 VDDA.n485 58.0576
R1232 VDDA.n414 VDDA.n413 58.0576
R1233 VDDA.n397 VDDA.n31 58.0576
R1234 VDDA.n390 VDDA.n34 58.0576
R1235 VDDA.n356 VDDA.n38 57.2449
R1236 VDDA.n372 VDDA.n371 57.2449
R1237 VDDA.n307 VDDA.n306 57.2449
R1238 VDDA.n293 VDDA.n292 57.2449
R1239 VDDA.n352 VDDA.n38 57.2449
R1240 VDDA.n306 VDDA.n58 57.2449
R1241 VDDA.n503 VDDA.n7 54.4005
R1242 VDDA.n9 VDDA.n7 54.4005
R1243 VDDA.n9 VDDA.n8 54.4005
R1244 VDDA.n503 VDDA.n8 54.4005
R1245 VDDA.n432 VDDA.n431 53.3664
R1246 VDDA.n453 VDDA.n447 53.3664
R1247 VDDA.n475 VDDA.n474 53.3664
R1248 VDDA.n326 VDDA.n325 53.3664
R1249 VDDA.n320 VDDA.n319 53.3664
R1250 VDDA.n412 VDDA.n26 53.3664
R1251 VDDA.n410 VDDA.n409 53.3664
R1252 VDDA.n484 VDDA.n18 53.3664
R1253 VDDA.n458 VDDA.n448 53.3664
R1254 VDDA.n438 VDDA.n437 53.3664
R1255 VDDA.n334 VDDA.n328 53.3664
R1256 VDDA.n330 VDDA.n318 53.3664
R1257 VDDA.n404 VDDA.n28 53.3664
R1258 VDDA.n400 VDDA.n27 53.3664
R1259 VDDA.n426 VDDA.n20 53.3664
R1260 VDDA.n422 VDDA.n19 53.3664
R1261 VDDA.n482 VDDA.n476 53.3664
R1262 VDDA.n478 VDDA.n428 53.3664
R1263 VDDA.n469 VDDA.n459 53.3664
R1264 VDDA.n464 VDDA.n429 53.3664
R1265 VDDA.n445 VDDA.n439 53.3664
R1266 VDDA.n441 VDDA.n430 53.3664
R1267 VDDA.n341 VDDA.n316 53.3664
R1268 VDDA.n337 VDDA.n316 53.3664
R1269 VDDA.n108 VDDA.t32 50.7639
R1270 VDDA.t63 VDDA.n85 49.2505
R1271 VDDA.n85 VDDA.t93 49.2505
R1272 VDDA.n78 VDDA.t105 49.2505
R1273 VDDA.n78 VDDA.t42 49.2505
R1274 VDDA.n109 VDDA.t45 49.2505
R1275 VDDA.n109 VDDA.t81 49.2505
R1276 VDDA.n89 VDDA.t103 49.2505
R1277 VDDA.n89 VDDA.t48 49.2505
R1278 VDDA.n82 VDDA.t91 49.2505
R1279 VDDA.n82 VDDA.t89 49.2505
R1280 VDDA.n84 VDDA.t95 49.2505
R1281 VDDA.n84 VDDA.t69 49.2505
R1282 VDDA VDDA.n517 47.763
R1283 VDDA.n348 VDDA.n344 45.3071
R1284 VDDA.n55 VDDA.n47 45.3071
R1285 VDDA.n56 VDDA.n48 45.3071
R1286 VDDA.n353 VDDA.n345 45.3071
R1287 VDDA.n289 VDDA.n285 45.3071
R1288 VDDA.n291 VDDA.n284 45.3071
R1289 VDDA.n313 VDDA.n49 45.3071
R1290 VDDA.n308 VDDA.n46 45.3071
R1291 VDDA.n368 VDDA.n364 45.3071
R1292 VDDA.n370 VDDA.n45 45.3071
R1293 VDDA.n362 VDDA.n354 45.3071
R1294 VDDA.n357 VDDA.n315 45.3071
R1295 VDDA.n118 VDDA.n88 45.3071
R1296 VDDA.n124 VDDA.n115 45.3071
R1297 VDDA.n95 VDDA.n93 45.3071
R1298 VDDA.n100 VDDA.n94 45.3071
R1299 VDDA.n101 VDDA.n93 45.3071
R1300 VDDA.n262 VDDA.n179 45.3071
R1301 VDDA.n184 VDDA.n178 45.3071
R1302 VDDA.n270 VDDA.n177 45.3071
R1303 VDDA.n268 VDDA.n267 45.3071
R1304 VDDA.n227 VDDA.n226 45.3071
R1305 VDDA.n226 VDDA.n223 45.3071
R1306 VDDA.n137 VDDA.n79 41.6005
R1307 VDDA.t84 VDDA.t35 39.886
R1308 VDDA.n131 VDDA.n80 39.4988
R1309 VDDA.n279 VDDA.n278 38.1005
R1310 VDDA.n113 VDDA.t55 36.26
R1311 VDDA.t15 VDDA.t80 32.6341
R1312 VDDA.t78 VDDA.t117 32.6341
R1313 VDDA.n261 VDDA.n180 32.2291
R1314 VDDA.n294 VDDA.n62 32.0005
R1315 VDDA.n298 VDDA.n62 32.0005
R1316 VDDA.n299 VDDA.n298 32.0005
R1317 VDDA.n300 VDDA.n299 32.0005
R1318 VDDA.n300 VDDA.n59 32.0005
R1319 VDDA.n306 VDDA.n59 32.0005
R1320 VDDA.n306 VDDA.n60 32.0005
R1321 VDDA.n60 VDDA.n42 32.0005
R1322 VDDA.n373 VDDA.n42 32.0005
R1323 VDDA.n377 VDDA.n40 32.0005
R1324 VDDA.n378 VDDA.n377 32.0005
R1325 VDDA.n379 VDDA.n378 32.0005
R1326 VDDA.n383 VDDA.n382 32.0005
R1327 VDDA.n384 VDDA.n383 32.0005
R1328 VDDA.n384 VDDA.n36 32.0005
R1329 VDDA.n388 VDDA.n36 32.0005
R1330 VDDA.n392 VDDA.n391 32.0005
R1331 VDDA.n392 VDDA.n30 32.0005
R1332 VDDA.n396 VDDA.n32 32.0005
R1333 VDDA.n419 VDDA.n22 32.0005
R1334 VDDA.n487 VDDA.n15 32.0005
R1335 VDDA.n491 VDDA.n13 32.0005
R1336 VDDA.n492 VDDA.n491 32.0005
R1337 VDDA.n493 VDDA.n492 32.0005
R1338 VDDA.n493 VDDA.n11 32.0005
R1339 VDDA.n497 VDDA.n11 32.0005
R1340 VDDA.n498 VDDA.n497 32.0005
R1341 VDDA.n499 VDDA.n498 32.0005
R1342 VDDA.n505 VDDA.n504 32.0005
R1343 VDDA.n505 VDDA.n5 32.0005
R1344 VDDA.n509 VDDA.n5 32.0005
R1345 VDDA.n510 VDDA.n509 32.0005
R1346 VDDA.n511 VDDA.n510 32.0005
R1347 VDDA.n511 VDDA.n3 32.0005
R1348 VDDA.n515 VDDA.n3 32.0005
R1349 VDDA.n135 VDDA.n80 32.0005
R1350 VDDA.n136 VDDA.n135 32.0005
R1351 VDDA.n138 VDDA.n75 32.0005
R1352 VDDA.n143 VDDA.n75 32.0005
R1353 VDDA.n144 VDDA.n143 32.0005
R1354 VDDA.n145 VDDA.n144 32.0005
R1355 VDDA.n145 VDDA.n72 32.0005
R1356 VDDA.n150 VDDA.n72 32.0005
R1357 VDDA.n151 VDDA.n150 32.0005
R1358 VDDA.n152 VDDA.n151 32.0005
R1359 VDDA.n152 VDDA.n69 32.0005
R1360 VDDA.n157 VDDA.n69 32.0005
R1361 VDDA.n158 VDDA.n157 32.0005
R1362 VDDA.n159 VDDA.n158 32.0005
R1363 VDDA.n159 VDDA.n66 32.0005
R1364 VDDA.n164 VDDA.n66 32.0005
R1365 VDDA.n165 VDDA.n164 32.0005
R1366 VDDA.n165 VDDA.n64 32.0005
R1367 VDDA.n169 VDDA.n64 32.0005
R1368 VDDA.n170 VDDA.n169 32.0005
R1369 VDDA.n274 VDDA.n172 32.0005
R1370 VDDA.n278 VDDA.n172 32.0005
R1371 VDDA.n198 VDDA.n197 32.0005
R1372 VDDA.n197 VDDA.n196 32.0005
R1373 VDDA.n204 VDDA.n186 32.0005
R1374 VDDA.n204 VDDA.n203 32.0005
R1375 VDDA.n203 VDDA.n202 32.0005
R1376 VDDA.n253 VDDA.n208 32.0005
R1377 VDDA.n248 VDDA.n247 32.0005
R1378 VDDA.n241 VDDA.n240 32.0005
R1379 VDDA.n241 VDDA.n212 32.0005
R1380 VDDA.n245 VDDA.n212 32.0005
R1381 VDDA.n234 VDDA.n233 32.0005
R1382 VDDA.n234 VDDA.n215 32.0005
R1383 VDDA.n238 VDDA.n215 32.0005
R1384 VDDA.n128 VDDA.n127 30.754
R1385 VDDA.n92 VDDA.n91 30.754
R1386 VDDA.n112 VDDA.n111 30.186
R1387 VDDA.n87 VDDA.n86 30.186
R1388 VDDA.n373 VDDA.n372 28.8005
R1389 VDDA.n273 VDDA.n174 28.8005
R1390 VDDA.n198 VDDA.n189 28.8005
R1391 VDDA.n254 VDDA.n253 28.8005
R1392 VDDA.n294 VDDA.n293 25.6005
R1393 VDDA.n379 VDDA.n38 25.6005
R1394 VDDA.n391 VDDA.n390 25.6005
R1395 VDDA.n415 VDDA.n414 25.6005
R1396 VDDA.n420 VDDA.n15 25.6005
R1397 VDDA.n487 VDDA.n486 25.6005
R1398 VDDA.n502 VDDA.n9 25.6005
R1399 VDDA.n503 VDDA.n502 25.6005
R1400 VDDA.n517 VDDA.n516 25.6005
R1401 VDDA.n137 VDDA.n136 25.6005
R1402 VDDA VDDA.n170 25.6005
R1403 VDDA.t4 VDDA.t102 25.3822
R1404 VDDA.t47 VDDA.t28 25.3822
R1405 VDDA.n355 VDDA.t118 24.6255
R1406 VDDA.n44 VDDA.t129 24.6255
R1407 VDDA.n50 VDDA.t31 24.6255
R1408 VDDA.n283 VDDA.t122 24.6255
R1409 VDDA.n346 VDDA.t114 24.6255
R1410 VDDA.n51 VDDA.t108 24.6255
R1411 VDDA.n191 VDDA.t99 24.6255
R1412 VDDA.n191 VDDA.t76 24.6255
R1413 VDDA.n188 VDDA.t38 24.6255
R1414 VDDA.n188 VDDA.t8 24.6255
R1415 VDDA.t73 VDDA.n255 24.6255
R1416 VDDA.n255 VDDA.t1 24.6255
R1417 VDDA.n211 VDDA.t101 24.6255
R1418 VDDA.n211 VDDA.t59 24.6255
R1419 VDDA.n214 VDDA.t40 24.6255
R1420 VDDA.n214 VDDA.t3 24.6255
R1421 VDDA.n231 VDDA.t66 24.6255
R1422 VDDA.n231 VDDA.t83 24.6255
R1423 VDDA.t66 VDDA.n230 24.6255
R1424 VDDA.n175 VDDA.t77 24.6255
R1425 VDDA.n256 VDDA.t73 24.6255
R1426 VDDA.n260 VDDA.t60 24.6255
R1427 VDDA.n220 VDDA.n217 24.361
R1428 VDDA.n196 VDDA.n192 22.4005
R1429 VDDA.n247 VDDA.n246 22.4005
R1430 VDDA.n248 VDDA.n180 22.4005
R1431 VDDA.n105 VDDA.n96 22.0449
R1432 VDDA.n116 VDDA.t56 19.7005
R1433 VDDA.n97 VDDA.t53 19.7005
R1434 VDDA.n67 VDDA.t79 19.7005
R1435 VDDA.n67 VDDA.t52 19.7005
R1436 VDDA.n70 VDDA.t85 19.7005
R1437 VDDA.n70 VDDA.t12 19.7005
R1438 VDDA.n73 VDDA.t29 19.7005
R1439 VDDA.n73 VDDA.t33 19.7005
R1440 VDDA.n76 VDDA.t14 19.7005
R1441 VDDA.n76 VDDA.t5 19.7005
R1442 VDDA.t56 VDDA.n81 19.7005
R1443 VDDA.n81 VDDA.t16 19.7005
R1444 VDDA.n32 VDDA.n24 19.2005
R1445 VDDA.t104 VDDA.t13 18.1303
R1446 VDDA.t116 VDDA.t51 18.1303
R1447 VDDA.n273 VDDA.n272 17.6005
R1448 VDDA.n397 VDDA.n396 16.0005
R1449 VDDA.n129 VDDA.n128 16.0005
R1450 VDDA.n91 VDDA.n90 16.0005
R1451 VDDA.n111 VDDA.n110 16.0005
R1452 VDDA.n86 VDDA.n83 16.0005
R1453 VDDA.n192 VDDA.n174 16.0005
R1454 VDDA.n208 VDDA.n180 16.0005
R1455 VDDA.n246 VDDA.n245 16.0005
R1456 VDDA.n233 VDDA.n232 16.0005
R1457 VDDA.n171 VDDA 15.7005
R1458 VDDA.n272 VDDA.n271 15.6449
R1459 VDDA.n229 VDDA.n220 15.6449
R1460 VDDA.n293 VDDA.n281 13.8989
R1461 VDDA.n398 VDDA.n30 12.8005
R1462 VDDA.n415 VDDA.n24 12.8005
R1463 VDDA.n280 VDDA.n171 12.7493
R1464 VDDA.n281 VDDA.n280 12.3383
R1465 VDDA.n280 VDDA.n279 11.579
R1466 VDDA.n343 VDDA.t24 11.4924
R1467 VDDA.t109 VDDA.n335 11.4924
R1468 VDDA.n327 VDDA.t106 11.4924
R1469 VDDA.n405 VDDA.t127 11.4924
R1470 VDDA.n411 VDDA.t119 11.4924
R1471 VDDA.t126 VDDA.t11 10.8784
R1472 VDDA.n96 VDDA.n65 9.613
R1473 VDDA.n274 VDDA.n273 9.6005
R1474 VDDA.n254 VDDA.n186 9.6005
R1475 VDDA.n202 VDDA.n189 9.6005
R1476 VDDA.n170 VDDA.n63 9.3005
R1477 VDDA.n169 VDDA.n168 9.3005
R1478 VDDA.n167 VDDA.n64 9.3005
R1479 VDDA.n166 VDDA.n165 9.3005
R1480 VDDA.n164 VDDA.n163 9.3005
R1481 VDDA.n162 VDDA.n66 9.3005
R1482 VDDA.n160 VDDA.n159 9.3005
R1483 VDDA.n158 VDDA.n68 9.3005
R1484 VDDA.n157 VDDA.n156 9.3005
R1485 VDDA.n155 VDDA.n69 9.3005
R1486 VDDA.n153 VDDA.n152 9.3005
R1487 VDDA.n151 VDDA.n71 9.3005
R1488 VDDA.n150 VDDA.n149 9.3005
R1489 VDDA.n148 VDDA.n72 9.3005
R1490 VDDA.n146 VDDA.n145 9.3005
R1491 VDDA.n144 VDDA.n74 9.3005
R1492 VDDA.n143 VDDA.n142 9.3005
R1493 VDDA.n141 VDDA.n75 9.3005
R1494 VDDA.n139 VDDA.n138 9.3005
R1495 VDDA.n133 VDDA.n80 9.3005
R1496 VDDA.n135 VDDA.n134 9.3005
R1497 VDDA.n136 VDDA.n77 9.3005
R1498 VDDA.n233 VDDA.n216 9.3005
R1499 VDDA.n235 VDDA.n234 9.3005
R1500 VDDA.n236 VDDA.n215 9.3005
R1501 VDDA.n238 VDDA.n237 9.3005
R1502 VDDA.n240 VDDA.n213 9.3005
R1503 VDDA.n242 VDDA.n241 9.3005
R1504 VDDA.n243 VDDA.n212 9.3005
R1505 VDDA.n245 VDDA.n244 9.3005
R1506 VDDA.n246 VDDA.n210 9.3005
R1507 VDDA.n247 VDDA.n209 9.3005
R1508 VDDA.n249 VDDA.n248 9.3005
R1509 VDDA.n250 VDDA.n180 9.3005
R1510 VDDA.n251 VDDA.n208 9.3005
R1511 VDDA.n253 VDDA.n252 9.3005
R1512 VDDA.n254 VDDA.n207 9.3005
R1513 VDDA.n206 VDDA.n186 9.3005
R1514 VDDA.n205 VDDA.n204 9.3005
R1515 VDDA.n203 VDDA.n187 9.3005
R1516 VDDA.n202 VDDA.n201 9.3005
R1517 VDDA.n200 VDDA.n189 9.3005
R1518 VDDA.n199 VDDA.n198 9.3005
R1519 VDDA.n197 VDDA.n190 9.3005
R1520 VDDA.n196 VDDA.n195 9.3005
R1521 VDDA.n194 VDDA.n192 9.3005
R1522 VDDA.n193 VDDA.n174 9.3005
R1523 VDDA.n273 VDDA.n173 9.3005
R1524 VDDA.n275 VDDA.n274 9.3005
R1525 VDDA.n276 VDDA.n172 9.3005
R1526 VDDA.n278 VDDA.n277 9.3005
R1527 VDDA.n517 VDDA.n0 9.3005
R1528 VDDA.n295 VDDA.n294 9.3005
R1529 VDDA.n296 VDDA.n62 9.3005
R1530 VDDA.n298 VDDA.n297 9.3005
R1531 VDDA.n299 VDDA.n61 9.3005
R1532 VDDA.n301 VDDA.n300 9.3005
R1533 VDDA.n302 VDDA.n59 9.3005
R1534 VDDA.n306 VDDA.n305 9.3005
R1535 VDDA.n304 VDDA.n60 9.3005
R1536 VDDA.n303 VDDA.n42 9.3005
R1537 VDDA.n374 VDDA.n373 9.3005
R1538 VDDA.n375 VDDA.n40 9.3005
R1539 VDDA.n377 VDDA.n376 9.3005
R1540 VDDA.n378 VDDA.n39 9.3005
R1541 VDDA.n380 VDDA.n379 9.3005
R1542 VDDA.n382 VDDA.n381 9.3005
R1543 VDDA.n383 VDDA.n37 9.3005
R1544 VDDA.n385 VDDA.n384 9.3005
R1545 VDDA.n386 VDDA.n36 9.3005
R1546 VDDA.n388 VDDA.n387 9.3005
R1547 VDDA.n391 VDDA.n33 9.3005
R1548 VDDA.n393 VDDA.n392 9.3005
R1549 VDDA.n394 VDDA.n30 9.3005
R1550 VDDA.n396 VDDA.n395 9.3005
R1551 VDDA.n32 VDDA.n23 9.3005
R1552 VDDA.n416 VDDA.n415 9.3005
R1553 VDDA.n417 VDDA.n22 9.3005
R1554 VDDA.n419 VDDA.n418 9.3005
R1555 VDDA.n15 VDDA.n14 9.3005
R1556 VDDA.n488 VDDA.n487 9.3005
R1557 VDDA.n489 VDDA.n13 9.3005
R1558 VDDA.n491 VDDA.n490 9.3005
R1559 VDDA.n492 VDDA.n12 9.3005
R1560 VDDA.n494 VDDA.n493 9.3005
R1561 VDDA.n495 VDDA.n11 9.3005
R1562 VDDA.n497 VDDA.n496 9.3005
R1563 VDDA.n498 VDDA.n10 9.3005
R1564 VDDA.n500 VDDA.n499 9.3005
R1565 VDDA.n502 VDDA.n501 9.3005
R1566 VDDA.n504 VDDA.n6 9.3005
R1567 VDDA.n506 VDDA.n505 9.3005
R1568 VDDA.n507 VDDA.n5 9.3005
R1569 VDDA.n509 VDDA.n508 9.3005
R1570 VDDA.n510 VDDA.n4 9.3005
R1571 VDDA.n512 VDDA.n511 9.3005
R1572 VDDA.n513 VDDA.n3 9.3005
R1573 VDDA.n515 VDDA.n514 9.3005
R1574 VDDA.n442 VDDA.n440 9.14336
R1575 VDDA.n479 VDDA.n477 9.14336
R1576 VDDA.n423 VDDA.n21 9.14336
R1577 VDDA.n401 VDDA.n29 9.14336
R1578 VDDA.n331 VDDA.n329 9.14336
R1579 VDDA.n436 VDDA.n435 9.14336
R1580 VDDA.n473 VDDA.n472 9.14336
R1581 VDDA.n408 VDDA.n407 9.14336
R1582 VDDA.n324 VDDA.n323 9.14336
R1583 VDDA.n340 VDDA.n339 9.14336
R1584 VDDA.t86 VDDA.t22 7.66179
R1585 VDDA.n126 VDDA.n125 7.25241
R1586 VDDA.n361 VDDA.n360 7.11161
R1587 VDDA.n358 VDDA.n356 7.11161
R1588 VDDA.n367 VDDA.n366 7.11161
R1589 VDDA.n371 VDDA.n43 7.11161
R1590 VDDA.n312 VDDA.n311 7.11161
R1591 VDDA.n309 VDDA.n307 7.11161
R1592 VDDA.n288 VDDA.n287 7.11161
R1593 VDDA.n292 VDDA.n282 7.11161
R1594 VDDA.n352 VDDA.n351 7.11161
R1595 VDDA.n349 VDDA.n347 7.11161
R1596 VDDA.n58 VDDA.n57 7.11161
R1597 VDDA.n54 VDDA.n53 7.11161
R1598 VDDA.n123 VDDA.n122 7.11161
R1599 VDDA.n120 VDDA.n119 7.11161
R1600 VDDA.n105 VDDA.n104 7.11161
R1601 VDDA.n102 VDDA.n99 7.11161
R1602 VDDA.n271 VDDA.n176 7.11161
R1603 VDDA.n266 VDDA.n264 7.11161
R1604 VDDA.n229 VDDA.n228 7.11161
R1605 VDDA.n222 VDDA.n219 7.11161
R1606 VDDA.n232 VDDA.n217 6.54033
R1607 VDDA.n382 VDDA.n38 6.4005
R1608 VDDA.n414 VDDA.n22 6.4005
R1609 VDDA.n420 VDDA.n419 6.4005
R1610 VDDA.n486 VDDA.n13 6.4005
R1611 VDDA.n499 VDDA.n9 6.4005
R1612 VDDA.n504 VDDA.n503 6.4005
R1613 VDDA.n516 VDDA.n515 6.4005
R1614 VDDA.n138 VDDA.n137 6.4005
R1615 VDDA.n465 VDDA.n461 5.81868
R1616 VDDA.n454 VDDA.n450 5.81868
R1617 VDDA.n336 VDDA.n34 5.33286
R1618 VDDA.n443 VDDA.n1 5.33286
R1619 VDDA.n480 VDDA.n16 5.33286
R1620 VDDA.n424 VDDA.n421 5.33286
R1621 VDDA.n402 VDDA.n399 5.33286
R1622 VDDA.n332 VDDA.n35 5.33286
R1623 VDDA.n433 VDDA.n2 5.33286
R1624 VDDA.n485 VDDA.n17 5.33286
R1625 VDDA.n413 VDDA.n25 5.33286
R1626 VDDA.n321 VDDA.n31 5.33286
R1627 VDDA.n444 VDDA.n440 3.75335
R1628 VDDA.n443 VDDA.n442 3.75335
R1629 VDDA.n481 VDDA.n477 3.75335
R1630 VDDA.n480 VDDA.n479 3.75335
R1631 VDDA.n425 VDDA.n21 3.75335
R1632 VDDA.n424 VDDA.n423 3.75335
R1633 VDDA.n403 VDDA.n29 3.75335
R1634 VDDA.n402 VDDA.n401 3.75335
R1635 VDDA.n333 VDDA.n329 3.75335
R1636 VDDA.n332 VDDA.n331 3.75335
R1637 VDDA.n436 VDDA.n433 3.75335
R1638 VDDA.n435 VDDA.n434 3.75335
R1639 VDDA.n472 VDDA.n17 3.75335
R1640 VDDA.n473 VDDA.n471 3.75335
R1641 VDDA.n407 VDDA.n25 3.75335
R1642 VDDA.n408 VDDA.n406 3.75335
R1643 VDDA.n324 VDDA.n321 3.75335
R1644 VDDA.n323 VDDA.n322 3.75335
R1645 VDDA.n340 VDDA.n336 3.75335
R1646 VDDA.n339 VDDA.n338 3.75335
R1647 VDDA.n360 VDDA.n359 3.53508
R1648 VDDA.n359 VDDA.n358 3.53508
R1649 VDDA.n366 VDDA.n365 3.53508
R1650 VDDA.n365 VDDA.n43 3.53508
R1651 VDDA.n311 VDDA.n310 3.53508
R1652 VDDA.n310 VDDA.n309 3.53508
R1653 VDDA.n287 VDDA.n286 3.53508
R1654 VDDA.n286 VDDA.n282 3.53508
R1655 VDDA.n351 VDDA.n350 3.53508
R1656 VDDA.n350 VDDA.n349 3.53508
R1657 VDDA.n57 VDDA.n52 3.53508
R1658 VDDA.n54 VDDA.n52 3.53508
R1659 VDDA.n122 VDDA.n121 3.53508
R1660 VDDA.n119 VDDA.n117 3.53508
R1661 VDDA.n121 VDDA.n120 3.53508
R1662 VDDA.n104 VDDA.n103 3.53508
R1663 VDDA.n99 VDDA.n98 3.53508
R1664 VDDA.n103 VDDA.n102 3.53508
R1665 VDDA.n265 VDDA.n176 3.53508
R1666 VDDA.n266 VDDA.n265 3.53508
R1667 VDDA.n228 VDDA.n218 3.53508
R1668 VDDA.n222 VDDA.n218 3.53508
R1669 VDDA.n468 VDDA.n467 3.40194
R1670 VDDA.n466 VDDA.n462 3.40194
R1671 VDDA.n457 VDDA.n456 3.40194
R1672 VDDA.n455 VDDA.n451 3.40194
R1673 VDDA.n372 VDDA.n40 3.2005
R1674 VDDA.n389 VDDA.n388 3.2005
R1675 VDDA.n390 VDDA.n389 3.2005
R1676 VDDA.n398 VDDA.n397 3.2005
R1677 VDDA.n240 VDDA.n239 3.2005
R1678 VDDA.n239 VDDA.n238 3.2005
R1679 VDDA.n467 VDDA.n461 2.39444
R1680 VDDA.n466 VDDA.n465 2.39444
R1681 VDDA.n456 VDDA.n450 2.39444
R1682 VDDA.n455 VDDA.n454 2.39444
R1683 VDDA.n462 VDDA.n7 2.32777
R1684 VDDA.n457 VDDA.n8 2.32777
R1685 VDDA.n182 VDDA.n181 2.27782
R1686 VDDA.n183 VDDA.n182 2.27782
R1687 VDDA.n259 VDDA.n257 2.27782
R1688 VDDA.n185 VDDA.n183 2.27782
R1689 VDDA.n261 VDDA.n181 2.27782
R1690 VDDA.n257 VDDA.n185 2.27782
R1691 VDDA.n217 VDDA.n216 0.703395
R1692 VDDA.n295 VDDA.n281 0.193961
R1693 VDDA.n171 VDDA.n63 0.188
R1694 VDDA.n134 VDDA.n133 0.15675
R1695 VDDA.n134 VDDA.n77 0.15675
R1696 VDDA.n139 VDDA.n77 0.15675
R1697 VDDA.n142 VDDA.n141 0.15675
R1698 VDDA.n142 VDDA.n74 0.15675
R1699 VDDA.n146 VDDA.n74 0.15675
R1700 VDDA.n149 VDDA.n148 0.15675
R1701 VDDA.n149 VDDA.n71 0.15675
R1702 VDDA.n153 VDDA.n71 0.15675
R1703 VDDA.n156 VDDA.n155 0.15675
R1704 VDDA.n156 VDDA.n68 0.15675
R1705 VDDA.n160 VDDA.n68 0.15675
R1706 VDDA.n163 VDDA.n162 0.15675
R1707 VDDA.n167 VDDA.n166 0.15675
R1708 VDDA.n168 VDDA.n167 0.15675
R1709 VDDA.n168 VDDA.n63 0.15675
R1710 VDDA.n235 VDDA.n216 0.15675
R1711 VDDA.n236 VDDA.n235 0.15675
R1712 VDDA.n237 VDDA.n236 0.15675
R1713 VDDA.n237 VDDA.n213 0.15675
R1714 VDDA.n242 VDDA.n213 0.15675
R1715 VDDA.n243 VDDA.n242 0.15675
R1716 VDDA.n244 VDDA.n243 0.15675
R1717 VDDA.n244 VDDA.n210 0.15675
R1718 VDDA.n210 VDDA.n209 0.15675
R1719 VDDA.n249 VDDA.n209 0.15675
R1720 VDDA.n250 VDDA.n249 0.15675
R1721 VDDA.n251 VDDA.n250 0.15675
R1722 VDDA.n252 VDDA.n251 0.15675
R1723 VDDA.n252 VDDA.n207 0.15675
R1724 VDDA.n207 VDDA.n206 0.15675
R1725 VDDA.n206 VDDA.n205 0.15675
R1726 VDDA.n205 VDDA.n187 0.15675
R1727 VDDA.n201 VDDA.n187 0.15675
R1728 VDDA.n201 VDDA.n200 0.15675
R1729 VDDA.n200 VDDA.n199 0.15675
R1730 VDDA.n199 VDDA.n190 0.15675
R1731 VDDA.n195 VDDA.n190 0.15675
R1732 VDDA.n195 VDDA.n194 0.15675
R1733 VDDA.n194 VDDA.n193 0.15675
R1734 VDDA.n193 VDDA.n173 0.15675
R1735 VDDA.n275 VDDA.n173 0.15675
R1736 VDDA.n276 VDDA.n275 0.15675
R1737 VDDA.n277 VDDA.n276 0.15675
R1738 VDDA.n296 VDDA.n295 0.15675
R1739 VDDA.n297 VDDA.n296 0.15675
R1740 VDDA.n297 VDDA.n61 0.15675
R1741 VDDA.n301 VDDA.n61 0.15675
R1742 VDDA.n302 VDDA.n301 0.15675
R1743 VDDA.n305 VDDA.n302 0.15675
R1744 VDDA.n305 VDDA.n304 0.15675
R1745 VDDA.n304 VDDA.n303 0.15675
R1746 VDDA.n375 VDDA.n374 0.15675
R1747 VDDA.n376 VDDA.n375 0.15675
R1748 VDDA.n376 VDDA.n39 0.15675
R1749 VDDA.n380 VDDA.n39 0.15675
R1750 VDDA.n381 VDDA.n380 0.15675
R1751 VDDA.n381 VDDA.n37 0.15675
R1752 VDDA.n385 VDDA.n37 0.15675
R1753 VDDA.n386 VDDA.n385 0.15675
R1754 VDDA.n387 VDDA.n386 0.15675
R1755 VDDA.n387 VDDA.n33 0.15675
R1756 VDDA.n393 VDDA.n33 0.15675
R1757 VDDA.n394 VDDA.n393 0.15675
R1758 VDDA.n395 VDDA.n394 0.15675
R1759 VDDA.n395 VDDA.n23 0.15675
R1760 VDDA.n416 VDDA.n23 0.15675
R1761 VDDA.n417 VDDA.n416 0.15675
R1762 VDDA.n418 VDDA.n417 0.15675
R1763 VDDA.n418 VDDA.n14 0.15675
R1764 VDDA.n488 VDDA.n14 0.15675
R1765 VDDA.n489 VDDA.n488 0.15675
R1766 VDDA.n490 VDDA.n489 0.15675
R1767 VDDA.n490 VDDA.n12 0.15675
R1768 VDDA.n494 VDDA.n12 0.15675
R1769 VDDA.n495 VDDA.n494 0.15675
R1770 VDDA.n496 VDDA.n495 0.15675
R1771 VDDA.n496 VDDA.n10 0.15675
R1772 VDDA.n500 VDDA.n10 0.15675
R1773 VDDA.n501 VDDA.n500 0.15675
R1774 VDDA.n501 VDDA.n6 0.15675
R1775 VDDA.n506 VDDA.n6 0.15675
R1776 VDDA.n507 VDDA.n506 0.15675
R1777 VDDA.n508 VDDA.n507 0.15675
R1778 VDDA.n508 VDDA.n4 0.15675
R1779 VDDA.n512 VDDA.n4 0.15675
R1780 VDDA.n513 VDDA.n512 0.15675
R1781 VDDA.n514 VDDA.n513 0.15675
R1782 VDDA.n514 VDDA.n0 0.15675
R1783 VDDA VDDA.n0 0.1255
R1784 VDDA.n277 VDDA 0.122375
R1785 VDDA.n132 VDDA.n131 0.100307
R1786 VDDA.n133 VDDA.n132 0.09425
R1787 VDDA.n141 VDDA.n140 0.09425
R1788 VDDA.n148 VDDA.n147 0.09425
R1789 VDDA.n155 VDDA.n154 0.09425
R1790 VDDA.n162 VDDA.n161 0.09425
R1791 VDDA.n166 VDDA.n65 0.09425
R1792 VDDA.n303 VDDA.n41 0.078625
R1793 VDDA.n374 VDDA.n41 0.078625
R1794 VDDA.n140 VDDA.n139 0.063
R1795 VDDA.n147 VDDA.n146 0.063
R1796 VDDA.n154 VDDA.n153 0.063
R1797 VDDA.n161 VDDA.n160 0.063
R1798 VDDA.n163 VDDA.n65 0.063
R1799 VDDA.n279 VDDA 0.0505
R1800 pfd_8_0.DOWN_PFD_b.t2 pfd_8_0.DOWN_PFD_b.n1 203.528
R1801 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 203.528
R1802 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R1803 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t1 183.935
R1804 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R1805 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R1806 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R1807 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R1808 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R1809 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R1810 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R1811 pfd_8_0.DOWN_b.t1 pfd_8_0.DOWN_b.n2 211.847
R1812 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t0 173.055
R1813 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R1814 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R1815 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R1816 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R1817 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R1818 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R1819 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R1820 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t0 221.411
R1821 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t1 24.0005
R1822 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R1823 a_870_1400.t0 a_870_1400.t1 39.4005
R1824 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t2 605.311
R1825 pfd_8_0.DOWN.t0 pfd_8_0.DOWN.n0 240.327
R1826 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 148.736
R1827 pfd_8_0.UP_input.n14 pfd_8_0.UP_input.n13 424.447
R1828 pfd_8_0.UP_input.n14 pfd_8_0.UP_input.n12 354.048
R1829 pfd_8_0.UP_input.t18 pfd_8_0.UP_input.n11 326.658
R1830 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n1 313
R1831 pfd_8_0.UP_input.n9 pfd_8_0.UP_input.t15 297.233
R1832 pfd_8_0.UP_input.t17 pfd_8_0.UP_input.n10 297.233
R1833 pfd_8_0.UP_input.n17 pfd_8_0.UP_input.t21 297.233
R1834 pfd_8_0.UP_input.n18 pfd_8_0.UP_input.t21 297.233
R1835 pfd_8_0.UP_input.t19 pfd_8_0.UP_input.n19 297.233
R1836 pfd_8_0.UP_input.n21 pfd_8_0.UP_input.t1 281.596
R1837 pfd_8_0.UP_input.n8 pfd_8_0.UP_input.n4 257.067
R1838 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 246.275
R1839 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n0 242.601
R1840 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t0 241.928
R1841 pfd_8_0.UP_input.n8 pfd_8_0.UP_input.n7 226.942
R1842 pfd_8_0.UP_input.n11 pfd_8_0.UP_input.n4 226.942
R1843 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 220.8
R1844 pfd_8_0.UP_input.n15 pfd_8_0.UP_input.n14 220.8
R1845 pfd_8_0.UP_input.n10 pfd_8_0.UP_input.n9 216.9
R1846 pfd_8_0.UP_input.n19 pfd_8_0.UP_input.n18 216.9
R1847 pfd_8_0.UP_input.n17 pfd_8_0.UP_input.n16 216.9
R1848 pfd_8_0.UP_input.n22 pfd_8_0.UP_input.n20 215.107
R1849 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t12 209.928
R1850 pfd_8_0.UP_input.n20 pfd_8_0.UP_input.n16 184.768
R1851 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t2 145.535
R1852 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n5 144
R1853 pfd_8_0.UP_input.n21 pfd_8_0.UP_input.t3 118.666
R1854 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.t15 92.3838
R1855 pfd_8_0.UP_input.n11 pfd_8_0.UP_input.t17 92.3838
R1856 pfd_8_0.UP_input.n9 pfd_8_0.UP_input.t14 80.3338
R1857 pfd_8_0.UP_input.t14 pfd_8_0.UP_input.n8 80.3338
R1858 pfd_8_0.UP_input.n10 pfd_8_0.UP_input.t20 80.3338
R1859 pfd_8_0.UP_input.t20 pfd_8_0.UP_input.n4 80.3338
R1860 pfd_8_0.UP_input.n18 pfd_8_0.UP_input.t22 80.3338
R1861 pfd_8_0.UP_input.t22 pfd_8_0.UP_input.n17 80.3338
R1862 pfd_8_0.UP_input.n19 pfd_8_0.UP_input.t13 80.3338
R1863 pfd_8_0.UP_input.t13 pfd_8_0.UP_input.n16 80.3338
R1864 pfd_8_0.UP_input.n20 pfd_8_0.UP_input.t19 80.3338
R1865 pfd_8_0.UP_input.n23 pfd_8_0.UP_input.n22 78.9255
R1866 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t16 70.0829
R1867 pfd_8_0.UP_input.n15 pfd_8_0.UP_input.t18 63.6829
R1868 opamp_cell_4_0.VOUT pfd_8_0.UP_input.n3 62.4005
R1869 pfd_8_0.UP_input.n23 pfd_8_0.UP_input.n15 60.8005
R1870 pfd_8_0.UP_input.n22 pfd_8_0.UP_input.n21 60.2361
R1871 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t10 60.0005
R1872 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t9 60.0005
R1873 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t8 60.0005
R1874 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t11 60.0005
R1875 pfd_8_0.UP_input.n13 pfd_8_0.UP_input.t4 49.2505
R1876 pfd_8_0.UP_input.n13 pfd_8_0.UP_input.t7 49.2505
R1877 pfd_8_0.UP_input.n12 pfd_8_0.UP_input.t6 49.2505
R1878 pfd_8_0.UP_input.n12 pfd_8_0.UP_input.t5 49.2505
R1879 opamp_cell_4_0.VOUT pfd_8_0.UP_input.n23 1.6005
R1880 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t8 377.567
R1881 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t9 297.233
R1882 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 243.44
R1883 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 224.496
R1884 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t7 216.9
R1885 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 196.262
R1886 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R1887 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R1888 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t6 136.567
R1889 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R1890 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 50.088
R1891 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t3 24.6255
R1892 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R1893 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t5 24.6255
R1894 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t4 24.6255
R1895 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t0 15.0005
R1896 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t1 15.0005
R1897 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.138
R1898 a_6320_5840.n7 a_6320_5840.n5 482.582
R1899 a_6320_5840.n10 a_6320_5840.t7 304.634
R1900 a_6320_5840.n3 a_6320_5840.t5 304.634
R1901 a_6320_5840.t9 a_6320_5840.n10 277.914
R1902 a_6320_5840.n3 a_6320_5840.t6 276.289
R1903 a_6320_5840.n8 a_6320_5840.n1 204.201
R1904 a_6320_5840.n4 a_6320_5840.n2 204.201
R1905 a_6320_5840.n9 a_6320_5840.n0 204.201
R1906 a_6320_5840.n7 a_6320_5840.n6 120.981
R1907 a_6320_5840.n8 a_6320_5840.n4 74.6672
R1908 a_6320_5840.n9 a_6320_5840.n8 74.6672
R1909 a_6320_5840.n1 a_6320_5840.t1 60.0005
R1910 a_6320_5840.n1 a_6320_5840.t11 60.0005
R1911 a_6320_5840.t6 a_6320_5840.n2 60.0005
R1912 a_6320_5840.n2 a_6320_5840.t2 60.0005
R1913 a_6320_5840.n0 a_6320_5840.t10 60.0005
R1914 a_6320_5840.n0 a_6320_5840.t8 60.0005
R1915 a_6320_5840.n8 a_6320_5840.n7 37.763
R1916 a_6320_5840.n5 a_6320_5840.t4 24.0005
R1917 a_6320_5840.n5 a_6320_5840.t3 24.0005
R1918 a_6320_5840.n6 a_6320_5840.t0 24.0005
R1919 a_6320_5840.n6 a_6320_5840.t12 24.0005
R1920 a_6320_5840.n4 a_6320_5840.n3 16.0005
R1921 a_6320_5840.n10 a_6320_5840.n9 16.0005
R1922 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_right.n6 1010.36
R1923 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 416.101
R1924 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 354.048
R1925 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 289.2
R1926 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R1927 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R1928 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R1929 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 284.2
R1930 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R1931 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R1932 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 208.868
R1933 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t0 60.0005
R1934 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R1935 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t2 49.2505
R1936 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R1937 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 401.668
R1938 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R1939 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R1940 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t0 252.248
R1941 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R1942 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R1943 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R1944 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R1945 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t5 60.0005
R1946 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t4 60.0005
R1947 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R1948 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R1949 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t1 49.2505
R1950 a_6490_4630.t2 a_6490_4630.n6 1112.76
R1951 a_6490_4630.n3 a_6490_4630.n2 416.863
R1952 a_6490_4630.n2 a_6490_4630.n1 366.848
R1953 a_6490_4630.n2 a_6490_4630.n0 271.401
R1954 a_6490_4630.n3 a_6490_4630.t5 208.868
R1955 a_6490_4630.n6 a_6490_4630.t6 208.868
R1956 a_6490_4630.n5 a_6490_4630.t7 208.868
R1957 a_6490_4630.n4 a_6490_4630.t8 208.868
R1958 a_6490_4630.n6 a_6490_4630.n5 208.868
R1959 a_6490_4630.n5 a_6490_4630.n4 208.868
R1960 a_6490_4630.n4 a_6490_4630.n3 193.804
R1961 a_6490_4630.n0 a_6490_4630.t4 60.0005
R1962 a_6490_4630.n0 a_6490_4630.t3 60.0005
R1963 a_6490_4630.n1 a_6490_4630.t1 49.2505
R1964 a_6490_4630.n1 a_6490_4630.t0 49.2505
R1965 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R1966 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R1967 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R1968 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R1969 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t0 172.458
R1970 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R1971 pfd_8_0.before_Reset.t1 pfd_8_0.before_Reset.n2 19.7005
R1972 a_2350_1400.t0 a_2350_1400.n2 500.086
R1973 a_2350_1400.n1 a_2350_1400.n0 473.334
R1974 a_2350_1400.n0 a_2350_1400.t3 465.933
R1975 a_2350_1400.t0 a_2350_1400.n2 461.389
R1976 a_2350_1400.n0 a_2350_1400.t2 321.334
R1977 a_2350_1400.n1 a_2350_1400.t1 177.577
R1978 a_2350_1400.n2 a_2350_1400.n1 48.3899
R1979 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t8 918.318
R1980 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R1981 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R1982 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R1983 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R1984 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R1985 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R1986 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R1987 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R1988 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R1989 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R1990 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R1991 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t4 120.501
R1992 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t0 120.501
R1993 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t2 120.501
R1994 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R1995 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t6 120.501
R1996 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R1997 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R1998 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R1999 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R2000 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R2001 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t1 19.7005
R2002 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t5 19.7005
R2003 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t7 19.7005
R2004 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t3 19.7005
R2005 F_REF.n0 F_REF.t0 514.134
R2006 F_REF.n0 F_REF.t1 273.134
R2007 F_REF F_REF.n0 216.9
R2008 a_n30_1400.t0 a_n30_1400.t1 39.4005
R2009 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R2010 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R2011 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R2012 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R2013 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R2014 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R2015 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R2016 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R2017 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R2018 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R2019 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R2020 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R2021 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R2022 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R2023 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R2024 pfd_8_0.I_IN.n4 pfd_8_0.I_IN.n3 1269.42
R2025 pfd_8_0.I_IN.n4 pfd_8_0.I_IN.t0 275.325
R2026 pfd_8_0.I_IN.n6 pfd_8_0.I_IN.n5 248.4
R2027 pfd_8_0.I_IN.n1 pfd_8_0.I_IN.t5 238.892
R2028 charge_pump_cell_6_0.I_IN pfd_8_0.I_IN.n6 214.4
R2029 pfd_8_0.I_IN.n1 pfd_8_0.I_IN.t4 161.371
R2030 pfd_8_0.I_IN.n2 pfd_8_0.I_IN.n1 160.639
R2031 pfd_8_0.I_IN.n3 pfd_8_0.I_IN.t6 151.792
R2032 pfd_8_0.I_IN.n5 pfd_8_0.I_IN.t2 140.583
R2033 pfd_8_0.I_IN.n5 pfd_8_0.I_IN.t0 140.583
R2034 pfd_8_0.I_IN.n2 pfd_8_0.I_IN.n0 95.4614
R2035 pfd_8_0.I_IN.t2 pfd_8_0.I_IN.n4 80.3338
R2036 pfd_8_0.I_IN.n3 pfd_8_0.I_IN.t7 44.2902
R2037 pfd_8_0.I_IN.n0 pfd_8_0.I_IN.t3 15.0005
R2038 pfd_8_0.I_IN.n0 pfd_8_0.I_IN.t1 15.0005
R2039 pfd_8_0.I_IN.n6 pfd_8_0.I_IN.n2 3.2005
R2040 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.t3 377.567
R2041 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t5 326.658
R2042 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t0 229.127
R2043 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 225.601
R2044 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 196.817
R2045 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t2 158.335
R2046 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t1 158.335
R2047 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 121.6
R2048 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN_input.n2 92.3838
R2049 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t4 92.3838
R2050 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 3.2005
R2051 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R2052 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R2053 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R2054 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R2055 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R2056 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R2057 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R2058 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R2059 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R2060 pfd_8_0.QB.n4 pfd_8_0.QB.t2 221.411
R2061 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R2062 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R2063 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R2064 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R2065 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R2066 a_1910_2020.t0 a_1910_2020.t1 48.0005
R2067 a_6220_5810.n4 a_6220_5810.t12 317.317
R2068 a_6220_5810.n2 a_6220_5810.t11 317.317
R2069 a_6220_5810.n5 a_6220_5810.n4 257.067
R2070 a_6220_5810.n3 a_6220_5810.n2 257.067
R2071 a_6220_5810.n10 a_6220_5810.n9 257.067
R2072 a_6220_5810.t8 a_6220_5810.n12 194.478
R2073 a_6220_5810.n8 a_6220_5810.n7 152
R2074 a_6220_5810.n12 a_6220_5810.n11 152
R2075 a_6220_5810.n1 a_6220_5810.n0 120.981
R2076 a_6220_5810.n7 a_6220_5810.n6 117.781
R2077 a_6220_5810.n7 a_6220_5810.n1 108.8
R2078 a_6220_5810.n8 a_6220_5810.n5 85.6894
R2079 a_6220_5810.n11 a_6220_5810.n3 85.6894
R2080 a_6220_5810.n11 a_6220_5810.n10 85.6894
R2081 a_6220_5810.n9 a_6220_5810.n8 85.6894
R2082 a_6220_5810.n4 a_6220_5810.t10 60.2505
R2083 a_6220_5810.n5 a_6220_5810.t0 60.2505
R2084 a_6220_5810.n2 a_6220_5810.t9 60.2505
R2085 a_6220_5810.n3 a_6220_5810.t2 60.2505
R2086 a_6220_5810.n10 a_6220_5810.t6 60.2505
R2087 a_6220_5810.n9 a_6220_5810.t4 60.2505
R2088 a_6220_5810.n6 a_6220_5810.t5 24.0005
R2089 a_6220_5810.n6 a_6220_5810.t1 24.0005
R2090 a_6220_5810.n0 a_6220_5810.t3 24.0005
R2091 a_6220_5810.n0 a_6220_5810.t7 24.0005
R2092 a_6220_5810.n12 a_6220_5810.n1 3.2005
R2093 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R2094 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R2095 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R2096 pfd_8_0.UP_PFD_b.t0 pfd_8_0.UP_PFD_b.n1 219.528
R2097 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t1 167.935
R2098 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R2099 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R2100 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R2101 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R2102 pfd_8_0.UP.t0 pfd_8_0.UP.n3 229.127
R2103 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R2104 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R2105 pfd_8_0.UP.n3 pfd_8_0.UP.t1 158.335
R2106 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R2107 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R2108 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R2109 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R2110 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R2111 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R2112 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R2113 pfd_8_0.E.t0 pfd_8_0.E.n4 221.411
R2114 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R2115 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R2116 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R2117 pfd_8_0.E.n1 pfd_8_0.E.t1 24.0005
R2118 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R2119 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R2120 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R2121 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R2122 pfd_8_0.E_b.t1 pfd_8_0.E_b.n2 221.411
R2123 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R2124 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R2125 a_1390_1400.t0 a_1390_1400.t1 39.4005
R2126 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R2127 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R2128 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R2129 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R2130 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R2131 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R2132 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R2133 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t0 221.411
R2134 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t1 24.0005
R2135 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R2136 a_870_640.t0 a_870_640.t1 39.4005
R2137 loop_filter_2_0.R1_C1.t0 loop_filter_2_0.R1_C1.t1 167.429
R2138 a_2530_190.t0 a_2530_190.n2 500.086
R2139 a_2530_190.n0 a_2530_190.t2 465.933
R2140 a_2530_190.t0 a_2530_190.n2 461.389
R2141 a_2530_190.n1 a_2530_190.n0 392.623
R2142 a_2530_190.n0 a_2530_190.t3 321.334
R2143 a_2530_190.n1 a_2530_190.t1 177.577
R2144 a_2530_190.n2 a_2530_190.n1 48.3899
R2145 a_2200_190.t0 a_2200_190.n2 500.086
R2146 a_2200_190.n1 a_2200_190.n0 473.334
R2147 a_2200_190.n0 a_2200_190.t2 465.933
R2148 a_2200_190.t0 a_2200_190.n2 461.389
R2149 a_2200_190.n0 a_2200_190.t3 321.334
R2150 a_2200_190.n1 a_2200_190.t1 177.577
R2151 a_2200_190.n2 a_2200_190.n1 48.3898
R2152 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R2153 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R2154 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R2155 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R2156 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R2157 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R2158 pfd_8_0.F.t0 pfd_8_0.F.n4 221.411
R2159 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R2160 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R2161 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R2162 pfd_8_0.F.n1 pfd_8_0.F.t1 24.0005
R2163 a_9360_6440.t0 a_9360_6440.t1 245.883
R2164 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 778.601
R2165 pfd_8_0.UP_b.t0 pfd_8_0.UP_b.n0 209.928
R2166 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t1 177.536
R2167 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R2168 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R2169 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R2170 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R2171 pfd_8_0.F_b.t1 pfd_8_0.F_b.n2 221.411
R2172 pfd_8_0.F_b.n1 pfd_8_0.F_b.t0 24.0005
R2173 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R2174 a_1390_640.t0 a_1390_640.t1 39.4005
R2175 a_490_640.t0 a_490_640.t1 39.4005
R2176 charge_pump_cell_6_0.UP_b.n0 charge_pump_cell_6_0.UP_b.t0 0.00505063
R2177 charge_pump_cell_6_0.UP_b charge_pump_cell_6_0.UP_b.n0 12.0576
R2178 charge_pump_cell_6_0.UP_b.n0 charge_pump_cell_6_0.UP_b.t1 323.788
R2179 a_490_1400.t0 a_490_1400.t1 39.4005
R2180 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R2181 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R2182 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R2183 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R2184 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R2185 pfd_8_0.Reset.t0 pfd_8_0.Reset.n3 288.37
R2186 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R2187 pfd_8_0.Reset.n3 pfd_8_0.Reset.t1 177.577
R2188 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R2189 charge_pump_cell_6_0.DOWN charge_pump_cell_6_0.DOWN.t0 12.0533
R2190 a_1870_190.t0 a_1870_190.n2 500.086
R2191 a_1870_190.n1 a_1870_190.n0 473.334
R2192 a_1870_190.n0 a_1870_190.t2 465.933
R2193 a_1870_190.t0 a_1870_190.n2 461.389
R2194 a_1870_190.n0 a_1870_190.t3 321.334
R2195 a_1870_190.n1 a_1870_190.t1 177.577
R2196 a_1870_190.n2 a_1870_190.n1 48.3898
R2197 a_n30_640.t0 a_n30_640.t1 39.4005
R2198 F_VCO.n0 F_VCO.t0 514.134
R2199 F_VCO.n0 F_VCO.t1 273.134
R2200 F_VCO F_VCO.n0 216.9
C0 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN- 0.010861f
C1 pfd_8_0.QB VDDA 2.7499f
C2 VDDA opamp_cell_4_0.VIN+ 0.924492f
C3 charge_pump_cell_6_0.UP_b opamp_cell_4_0.p_bias 0.041967f
C4 pfd_8_0.QB_b VDDA 0.511838f
C5 pfd_8_0.QB pfd_8_0.QB_b 0.388258f
C6 pfd_8_0.QA_b VDDA 0.52066f
C7 VDDA F_REF 0.098433f
C8 VDDA opamp_cell_4_0.VIN- 0.171047f
C9 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN- 0.133176f
C10 charge_pump_cell_6_0.UP_b charge_pump_cell_6_0.DOWN 0.049574f
C11 pfd_8_0.QA_b F_REF 0.027208f
C12 VDDA pfd_8_0.QA 0.550605f
C13 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN_input 0.200808f
C14 pfd_8_0.QB pfd_8_0.QA 0.074487f
C15 opamp_cell_4_0.p_bias VDDA 2.86573f
C16 VDDA F_VCO 0.12889f
C17 pfd_8_0.QB F_VCO 0.058558f
C18 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.098414f
C19 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C20 F_REF pfd_8_0.QA 0.056f
C21 charge_pump_cell_6_0.UP_b VDDA 0.396833f
C22 pfd_8_0.QB_b F_VCO 0.039516f
C23 charge_pump_cell_6_0.UP_b opamp_cell_4_0.VIN+ 0.011697f
C24 VDDA pfd_8_0.DOWN_input 0.221393f
C25 opamp_cell_4_0.VIN+ pfd_8_0.DOWN_input 0.072856f
C26 F_VCO V_OUT 0.389374f
C27 F_REF V_OUT 0.277742f
C28 VDDA V_OUT 45.160034f
C29 charge_pump_cell_6_0.DOWN V_OUT 2.98421f
C30 pfd_8_0.DOWN_input V_OUT 3.49455f
C31 pfd_8_0.QB_b V_OUT 1.05311f
C32 pfd_8_0.QB V_OUT 1.307381f
C33 pfd_8_0.QA V_OUT 3.10102f
C34 pfd_8_0.QA_b V_OUT 1.05138f
C35 charge_pump_cell_6_0.UP_b V_OUT 6.21267f
C36 opamp_cell_4_0.VIN+ V_OUT 3.98071f
C37 opamp_cell_4_0.VIN- V_OUT 1.2483f
C38 opamp_cell_4_0.p_bias V_OUT 3.989291f
C39 pfd_8_0.QB.t7 V_OUT 0.066708f
C40 pfd_8_0.QB.t8 V_OUT 0.031333f
C41 pfd_8_0.QB.n0 V_OUT 0.096363f
C42 pfd_8_0.QB.t3 V_OUT 0.066708f
C43 pfd_8_0.QB.t4 V_OUT 0.100569f
C44 pfd_8_0.QB.n1 V_OUT 1.20598f
C45 pfd_8_0.QB.t5 V_OUT 0.067367f
C46 pfd_8_0.QB.t6 V_OUT 0.029539f
C47 pfd_8_0.QB.n2 V_OUT 0.170164f
C48 pfd_8_0.QB.t2 V_OUT 0.14186f
C49 pfd_8_0.QB.t0 V_OUT 0.026953f
C50 pfd_8_0.QB.t1 V_OUT 0.026953f
C51 pfd_8_0.QB.n3 V_OUT 0.143916f
C52 pfd_8_0.QB.n4 V_OUT 0.255686f
C53 pfd_8_0.QB.n5 V_OUT 0.218372f
C54 opamp_cell_4_0.p_bias.t8 V_OUT 1.66267f
C55 opamp_cell_4_0.p_bias.t1 V_OUT 0.019693f
C56 opamp_cell_4_0.p_bias.t5 V_OUT 0.019693f
C57 opamp_cell_4_0.p_bias.n0 V_OUT 0.054067f
C58 opamp_cell_4_0.p_bias.t7 V_OUT 0.019693f
C59 opamp_cell_4_0.p_bias.t3 V_OUT 0.019693f
C60 opamp_cell_4_0.p_bias.n1 V_OUT 0.054067f
C61 opamp_cell_4_0.p_bias.n2 V_OUT 0.068502f
C62 opamp_cell_4_0.p_bias.t0 V_OUT 0.054353f
C63 opamp_cell_4_0.p_bias.t2 V_OUT 0.054353f
C64 opamp_cell_4_0.p_bias.t6 V_OUT 0.054353f
C65 opamp_cell_4_0.p_bias.t11 V_OUT 0.054353f
C66 opamp_cell_4_0.p_bias.t9 V_OUT 0.074733f
C67 opamp_cell_4_0.p_bias.n3 V_OUT 0.04185f
C68 opamp_cell_4_0.p_bias.n4 V_OUT 0.029697f
C69 opamp_cell_4_0.p_bias.n5 V_OUT 0.012761f
C70 opamp_cell_4_0.p_bias.n6 V_OUT 0.029697f
C71 opamp_cell_4_0.p_bias.n7 V_OUT 0.029697f
C72 opamp_cell_4_0.p_bias.t4 V_OUT 0.054353f
C73 opamp_cell_4_0.p_bias.t12 V_OUT 0.054353f
C74 opamp_cell_4_0.p_bias.t10 V_OUT 0.074733f
C75 opamp_cell_4_0.p_bias.n8 V_OUT 0.04185f
C76 opamp_cell_4_0.p_bias.n9 V_OUT 0.029697f
C77 opamp_cell_4_0.p_bias.n10 V_OUT 0.012761f
C78 opamp_cell_4_0.p_bias.n11 V_OUT 0.120625f
C79 opamp_cell_4_0.VIN+.t8 V_OUT 0.023149f
C80 opamp_cell_4_0.VIN+.t7 V_OUT 0.016337f
C81 opamp_cell_4_0.VIN+.n0 V_OUT 0.042889f
C82 opamp_cell_4_0.VIN+.t9 V_OUT 0.014474f
C83 opamp_cell_4_0.VIN+.n1 V_OUT 0.038113f
C84 opamp_cell_4_0.VIN+.n2 V_OUT 0.297842f
C85 opamp_cell_4_0.VIN+.t3 V_OUT 0.039604f
C86 opamp_cell_4_0.VIN+.t2 V_OUT 0.039604f
C87 opamp_cell_4_0.VIN+.n3 V_OUT 0.097602f
C88 opamp_cell_4_0.VIN+.t0 V_OUT 0.039604f
C89 opamp_cell_4_0.VIN+.t1 V_OUT 0.039604f
C90 opamp_cell_4_0.VIN+.n4 V_OUT 0.265157f
C91 opamp_cell_4_0.VIN+.n5 V_OUT 0.416646f
C92 opamp_cell_4_0.VIN+.t5 V_OUT 0.039604f
C93 opamp_cell_4_0.VIN+.t4 V_OUT 0.039604f
C94 opamp_cell_4_0.VIN+.n6 V_OUT 0.097602f
C95 opamp_cell_4_0.VIN+.n7 V_OUT 0.468809f
C96 pfd_8_0.UP_input.t16 V_OUT 2.22616f
C97 pfd_8_0.UP_input.n2 V_OUT 0.022396f
C98 pfd_8_0.UP_input.n3 V_OUT 0.019378f
C99 pfd_8_0.UP_input.n4 V_OUT 0.011811f
C100 pfd_8_0.UP_input.t20 V_OUT 0.013068f
C101 pfd_8_0.UP_input.t15 V_OUT 0.022473f
C102 pfd_8_0.UP_input.t2 V_OUT 0.010448f
C103 pfd_8_0.UP_input.t0 V_OUT 0.025333f
C104 pfd_8_0.UP_input.n5 V_OUT 0.031065f
C105 pfd_8_0.UP_input.t12 V_OUT 0.023005f
C106 pfd_8_0.UP_input.n6 V_OUT 0.108905f
C107 pfd_8_0.UP_input.n7 V_OUT 0.023305f
C108 pfd_8_0.UP_input.n8 V_OUT 0.011811f
C109 pfd_8_0.UP_input.t14 V_OUT 0.013068f
C110 pfd_8_0.UP_input.n9 V_OUT 0.015753f
C111 pfd_8_0.UP_input.n10 V_OUT 0.015753f
C112 pfd_8_0.UP_input.t17 V_OUT 0.022473f
C113 pfd_8_0.UP_input.n11 V_OUT 0.022906f
C114 pfd_8_0.UP_input.t18 V_OUT 3.24153f
C115 pfd_8_0.UP_input.n14 V_OUT 0.030112f
C116 pfd_8_0.UP_input.n15 V_OUT 0.019856f
C117 pfd_8_0.UP_input.n16 V_OUT 0.012216f
C118 pfd_8_0.UP_input.t13 V_OUT 0.013068f
C119 pfd_8_0.UP_input.t21 V_OUT 0.029916f
C120 pfd_8_0.UP_input.n17 V_OUT 0.015753f
C121 pfd_8_0.UP_input.t22 V_OUT 0.013068f
C122 pfd_8_0.UP_input.n18 V_OUT 0.015753f
C123 pfd_8_0.UP_input.n19 V_OUT 0.015753f
C124 pfd_8_0.UP_input.t19 V_OUT 0.021492f
C125 pfd_8_0.UP_input.n20 V_OUT 0.014914f
C126 pfd_8_0.UP_input.t1 V_OUT 0.027948f
C127 pfd_8_0.UP_input.n21 V_OUT 0.035654f
C128 pfd_8_0.UP_input.n22 V_OUT 0.188444f
C129 pfd_8_0.UP_input.n23 V_OUT 0.110692f
C130 VDDA.n1 V_OUT 0.011281f
C131 VDDA.n2 V_OUT 0.011281f
C132 VDDA.n16 V_OUT 0.011281f
C133 VDDA.t22 V_OUT 0.047758f
C134 VDDA.t120 V_OUT 0.01732f
C135 VDDA.n24 V_OUT 0.018969f
C136 VDDA.t127 V_OUT 0.047758f
C137 VDDA.n31 V_OUT 0.011281f
C138 VDDA.n34 V_OUT 0.010259f
C139 VDDA.n35 V_OUT 0.011281f
C140 VDDA.n41 V_OUT 0.043944f
C141 VDDA.n43 V_OUT 0.010271f
C142 VDDA.n44 V_OUT 0.017118f
C143 VDDA.t30 V_OUT 0.160962f
C144 VDDA.n50 V_OUT 0.017118f
C145 VDDA.n51 V_OUT 0.017118f
C146 VDDA.n53 V_OUT 0.010366f
C147 VDDA.n54 V_OUT 0.010271f
C148 VDDA.n57 V_OUT 0.010271f
C149 VDDA.n58 V_OUT 0.012107f
C150 VDDA.n67 V_OUT 0.014937f
C151 VDDA.n70 V_OUT 0.014937f
C152 VDDA.n73 V_OUT 0.014937f
C153 VDDA.n76 V_OUT 0.014937f
C154 VDDA.n79 V_OUT 0.015944f
C155 VDDA.n81 V_OUT 0.014937f
C156 VDDA.n83 V_OUT 0.012338f
C157 VDDA.t70 V_OUT 0.010226f
C158 VDDA.t63 V_OUT 0.013084f
C159 VDDA.n87 V_OUT 0.078421f
C160 VDDA.t62 V_OUT 0.192072f
C161 VDDA.t92 V_OUT 0.097171f
C162 VDDA.t90 V_OUT 0.097171f
C163 VDDA.t88 V_OUT 0.097171f
C164 VDDA.t94 V_OUT 0.097171f
C165 VDDA.t68 V_OUT 0.110251f
C166 VDDA.n90 V_OUT 0.012338f
C167 VDDA.t49 V_OUT 0.010226f
C168 VDDA.n92 V_OUT 0.021462f
C169 VDDA.t50 V_OUT 0.028263f
C170 VDDA.n97 V_OUT 0.021397f
C171 VDDA.n98 V_OUT 0.010209f
C172 VDDA.n99 V_OUT 0.010271f
C173 VDDA.n102 V_OUT 0.010271f
C174 VDDA.n104 V_OUT 0.010271f
C175 VDDA.n107 V_OUT 0.155099f
C176 VDDA.t34 V_OUT 0.074747f
C177 VDDA.t51 V_OUT 0.048585f
C178 VDDA.t116 V_OUT 0.057929f
C179 VDDA.t117 V_OUT 0.065403f
C180 VDDA.t78 V_OUT 0.048585f
C181 VDDA.t125 V_OUT 0.074747f
C182 VDDA.t11 V_OUT 0.048585f
C183 VDDA.t126 V_OUT 0.054191f
C184 VDDA.t35 V_OUT 0.069141f
C185 VDDA.t84 V_OUT 0.095302f
C186 VDDA.t32 V_OUT 0.100908f
C187 VDDA.n108 V_OUT 0.08054f
C188 VDDA.t28 V_OUT 0.061666f
C189 VDDA.t47 V_OUT 0.061666f
C190 VDDA.t102 V_OUT 0.061666f
C191 VDDA.t4 V_OUT 0.048585f
C192 VDDA.t41 V_OUT 0.074747f
C193 VDDA.t13 V_OUT 0.048585f
C194 VDDA.t104 V_OUT 0.057929f
C195 VDDA.t80 V_OUT 0.065403f
C196 VDDA.t15 V_OUT 0.048585f
C197 VDDA.t44 V_OUT 0.074747f
C198 VDDA.t55 V_OUT 0.061666f
C199 VDDA.t45 V_OUT 0.013084f
C200 VDDA.n110 V_OUT 0.012338f
C201 VDDA.n112 V_OUT 0.025501f
C202 VDDA.n113 V_OUT 0.08055f
C203 VDDA.t54 V_OUT 0.028842f
C204 VDDA.t56 V_OUT 0.014265f
C205 VDDA.n116 V_OUT 0.021397f
C206 VDDA.n117 V_OUT 0.010209f
C207 VDDA.n119 V_OUT 0.010271f
C208 VDDA.n120 V_OUT 0.010271f
C209 VDDA.n122 V_OUT 0.010271f
C210 VDDA.n123 V_OUT 0.020153f
C211 VDDA.n125 V_OUT 0.059797f
C212 VDDA.n126 V_OUT 0.071197f
C213 VDDA.n127 V_OUT 0.021462f
C214 VDDA.n129 V_OUT 0.012338f
C215 VDDA.n130 V_OUT 0.01766f
C216 VDDA.n131 V_OUT 0.051309f
C217 VDDA.n132 V_OUT 0.051555f
C218 VDDA.n140 V_OUT 0.049996f
C219 VDDA.n147 V_OUT 0.049996f
C220 VDDA.n154 V_OUT 0.049996f
C221 VDDA.n161 V_OUT 0.049996f
C222 VDDA.n171 V_OUT 0.033572f
C223 VDDA.n175 V_OUT 0.017118f
C224 VDDA.n176 V_OUT 0.010271f
C225 VDDA.t58 V_OUT 0.071152f
C226 VDDA.n182 V_OUT 0.015976f
C227 VDDA.n185 V_OUT 0.015976f
C228 VDDA.n188 V_OUT 0.016498f
C229 VDDA.n189 V_OUT 0.023215f
C230 VDDA.n191 V_OUT 0.016498f
C231 VDDA.n192 V_OUT 0.023215f
C232 VDDA.n211 V_OUT 0.016498f
C233 VDDA.n214 V_OUT 0.016498f
C234 VDDA.n216 V_OUT 0.014676f
C235 VDDA.t64 V_OUT 0.028441f
C236 VDDA.n220 V_OUT 0.011186f
C237 VDDA.n222 V_OUT 0.010271f
C238 VDDA.t100 V_OUT 0.072807f
C239 VDDA.t2 V_OUT 0.072807f
C240 VDDA.t39 V_OUT 0.072807f
C241 VDDA.t82 V_OUT 0.072807f
C242 VDDA.t65 V_OUT 0.071152f
C243 VDDA.n225 V_OUT 0.064533f
C244 VDDA.n228 V_OUT 0.010271f
C245 VDDA.n229 V_OUT 0.010364f
C246 VDDA.n230 V_OUT 0.017118f
C247 VDDA.t66 V_OUT 0.011412f
C248 VDDA.n231 V_OUT 0.016498f
C249 VDDA.n232 V_OUT 0.023509f
C250 VDDA.n239 V_OUT 0.022074f
C251 VDDA.n246 V_OUT 0.023215f
C252 VDDA.n254 V_OUT 0.023215f
C253 VDDA.n255 V_OUT 0.016498f
C254 VDDA.t73 V_OUT 0.011412f
C255 VDDA.n256 V_OUT 0.017118f
C256 VDDA.t57 V_OUT 0.026837f
C257 VDDA.t71 V_OUT 0.026837f
C258 VDDA.n258 V_OUT 0.01209f
C259 VDDA.n259 V_OUT 0.020603f
C260 VDDA.n260 V_OUT 0.017118f
C261 VDDA.n261 V_OUT 0.01941f
C262 VDDA.n263 V_OUT 0.069497f
C263 VDDA.t72 V_OUT 0.071152f
C264 VDDA.t0 V_OUT 0.072807f
C265 VDDA.t37 V_OUT 0.072807f
C266 VDDA.t7 V_OUT 0.072807f
C267 VDDA.t98 V_OUT 0.072807f
C268 VDDA.t75 V_OUT 0.071152f
C269 VDDA.n264 V_OUT 0.010366f
C270 VDDA.n266 V_OUT 0.010271f
C271 VDDA.n269 V_OUT 0.064533f
C272 VDDA.n271 V_OUT 0.011486f
C273 VDDA.t74 V_OUT 0.028441f
C274 VDDA.n279 V_OUT 0.023362f
C275 VDDA.n280 V_OUT 0.244464f
C276 VDDA.n281 V_OUT 0.04381f
C277 VDDA.n282 V_OUT 0.010271f
C278 VDDA.n283 V_OUT 0.017118f
C279 VDDA.t121 V_OUT 0.168037f
C280 VDDA.t19 V_OUT 0.182188f
C281 VDDA.n287 V_OUT 0.010271f
C282 VDDA.n288 V_OUT 0.010366f
C283 VDDA.n290 V_OUT 0.137968f
C284 VDDA.n292 V_OUT 0.012107f
C285 VDDA.n307 V_OUT 0.012107f
C286 VDDA.n309 V_OUT 0.010271f
C287 VDDA.n311 V_OUT 0.010271f
C288 VDDA.n312 V_OUT 0.010366f
C289 VDDA.n314 V_OUT 0.137968f
C290 VDDA.t115 V_OUT 0.137968f
C291 VDDA.t106 V_OUT 0.047758f
C292 VDDA.t128 V_OUT 0.012035f
C293 VDDA.n322 V_OUT 0.011114f
C294 VDDA.n327 V_OUT 0.068984f
C295 VDDA.t25 V_OUT 0.012035f
C296 VDDA.n333 V_OUT 0.011114f
C297 VDDA.n335 V_OUT 0.068984f
C298 VDDA.t109 V_OUT 0.047758f
C299 VDDA.t24 V_OUT 0.047758f
C300 VDDA.t110 V_OUT 0.012035f
C301 VDDA.n338 V_OUT 0.010062f
C302 VDDA.n343 V_OUT 0.097285f
C303 VDDA.n346 V_OUT 0.017118f
C304 VDDA.n347 V_OUT 0.010366f
C305 VDDA.n349 V_OUT 0.010271f
C306 VDDA.n351 V_OUT 0.010271f
C307 VDDA.n352 V_OUT 0.012107f
C308 VDDA.n355 V_OUT 0.017118f
C309 VDDA.n356 V_OUT 0.012107f
C310 VDDA.n358 V_OUT 0.010271f
C311 VDDA.n360 V_OUT 0.010271f
C312 VDDA.n361 V_OUT 0.010366f
C313 VDDA.n363 V_OUT 0.150349f
C314 VDDA.t113 V_OUT 0.137968f
C315 VDDA.n366 V_OUT 0.010271f
C316 VDDA.n367 V_OUT 0.010366f
C317 VDDA.n369 V_OUT 0.137968f
C318 VDDA.n371 V_OUT 0.012107f
C319 VDDA.n399 V_OUT 0.011281f
C320 VDDA.t107 V_OUT 0.012035f
C321 VDDA.n403 V_OUT 0.011114f
C322 VDDA.n405 V_OUT 0.068984f
C323 VDDA.t23 V_OUT 0.012035f
C324 VDDA.n406 V_OUT 0.011114f
C325 VDDA.t86 V_OUT 0.042452f
C326 VDDA.t119 V_OUT 0.04422f
C327 VDDA.n411 V_OUT 0.068984f
C328 VDDA.n413 V_OUT 0.011281f
C329 VDDA.n421 V_OUT 0.011068f
C330 VDDA.t87 V_OUT 0.011976f
C331 VDDA.n425 V_OUT 0.011114f
C332 VDDA.n427 V_OUT 0.093747f
C333 VDDA.t111 V_OUT 0.012035f
C334 VDDA.n434 V_OUT 0.011114f
C335 VDDA.t97 V_OUT 0.012035f
C336 VDDA.n444 V_OUT 0.011114f
C337 VDDA.n446 V_OUT 0.10436f
C338 VDDA.t96 V_OUT 0.086672f
C339 VDDA.t17 V_OUT 0.183957f
C340 VDDA.t124 V_OUT 0.183957f
C341 VDDA.t26 V_OUT 0.086672f
C342 VDDA.n450 V_OUT 0.012553f
C343 VDDA.n451 V_OUT 0.015024f
C344 VDDA.n454 V_OUT 0.012553f
C345 VDDA.t18 V_OUT 0.012041f
C346 VDDA.n457 V_OUT 0.012514f
C347 VDDA.n461 V_OUT 0.012553f
C348 VDDA.n462 V_OUT 0.012514f
C349 VDDA.n465 V_OUT 0.012553f
C350 VDDA.t10 V_OUT 0.012041f
C351 VDDA.n468 V_OUT 0.015024f
C352 VDDA.n470 V_OUT 0.095516f
C353 VDDA.t9 V_OUT 0.086672f
C354 VDDA.t6 V_OUT 0.183957f
C355 VDDA.t112 V_OUT 0.183957f
C356 VDDA.t20 V_OUT 0.086672f
C357 VDDA.t36 V_OUT 0.012035f
C358 VDDA.n471 V_OUT 0.011114f
C359 VDDA.t21 V_OUT 0.012035f
C360 VDDA.n481 V_OUT 0.011114f
C361 VDDA.n483 V_OUT 0.097285f
C362 VDDA.n485 V_OUT 0.011281f
C363 a_5970_4630.t6 V_OUT 0.030769f
C364 a_5970_4630.n0 V_OUT 0.124795f
C365 a_5970_4630.t12 V_OUT 0.020325f
C366 a_5970_4630.t11 V_OUT 0.020325f
C367 a_5970_4630.t10 V_OUT 0.020325f
C368 a_5970_4630.n1 V_OUT 0.044943f
C369 a_5970_4630.t9 V_OUT 0.020325f
C370 a_5970_4630.t4 V_OUT 0.020325f
C371 a_5970_4630.n2 V_OUT 0.044943f
C372 a_5970_4630.t5 V_OUT 0.077457f
C373 a_5970_4630.t3 V_OUT 0.030769f
C374 a_5970_4630.n3 V_OUT 0.097952f
C375 a_5970_4630.n4 V_OUT 0.087903f
C376 a_5970_4630.n5 V_OUT 0.089425f
C377 a_5970_4630.t2 V_OUT 0.050813f
C378 a_5970_4630.t1 V_OUT 0.050813f
C379 a_5970_4630.n6 V_OUT 0.295522f
C380 a_5970_4630.t0 V_OUT 0.050813f
C381 a_5970_4630.t8 V_OUT 0.050813f
C382 a_5970_4630.n7 V_OUT 0.144587f
C383 a_5970_4630.n8 V_OUT 0.360746f
C384 a_5970_4630.n9 V_OUT 0.13437f
C385 a_5970_4630.n10 V_OUT 0.085474f
C386 a_5970_4630.n11 V_OUT 0.045257f
C387 a_5970_4630.t7 V_OUT 0.100208f
.ends

