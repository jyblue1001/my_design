magic
tech sky130A
timestamp 1748864850
<< pwell >>
rect 2990 2830 5010 2930
rect 2810 2400 5190 2700
rect 2565 1900 2715 2000
rect 2745 1900 3985 2000
rect 4015 1900 5255 2000
rect -45 1685 130 1725
rect 3165 1615 3805 1665
rect 4195 1615 4835 1665
rect 2835 1210 3955 1460
rect 4045 1210 5165 1460
rect 2940 980 5060 1080
rect 2990 785 5010 885
<< nmos >>
rect 3030 2830 3080 2930
rect 3120 2830 3170 2930
rect 3210 2830 3260 2930
rect 3300 2830 3350 2930
rect 3390 2830 3440 2930
rect 3480 2830 3530 2930
rect 3570 2830 3620 2930
rect 3660 2830 3710 2930
rect 3750 2830 3800 2930
rect 3840 2830 3890 2930
rect 3930 2830 3980 2930
rect 4020 2830 4070 2930
rect 4110 2830 4160 2930
rect 4200 2830 4250 2930
rect 4290 2830 4340 2930
rect 4380 2830 4430 2930
rect 4470 2830 4520 2930
rect 4560 2830 4610 2930
rect 4650 2830 4700 2930
rect 4740 2830 4790 2930
rect 4830 2830 4880 2930
rect 4920 2830 4970 2930
rect 2850 2400 2900 2700
rect 2940 2400 2990 2700
rect 3030 2400 3080 2700
rect 3120 2400 3170 2700
rect 3210 2400 3260 2700
rect 3300 2400 3350 2700
rect 3390 2400 3440 2700
rect 3480 2400 3530 2700
rect 3570 2400 3620 2700
rect 3660 2400 3710 2700
rect 3750 2400 3800 2700
rect 3840 2400 3890 2700
rect 3930 2400 3980 2700
rect 4020 2400 4070 2700
rect 4110 2400 4160 2700
rect 4200 2400 4250 2700
rect 4290 2400 4340 2700
rect 4380 2400 4430 2700
rect 4470 2400 4520 2700
rect 4560 2400 4610 2700
rect 4650 2400 4700 2700
rect 4740 2400 4790 2700
rect 4830 2400 4880 2700
rect 4920 2400 4970 2700
rect 5010 2400 5060 2700
rect 5100 2400 5150 2700
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4055 1900 4075 2000
rect 4115 1900 4135 2000
rect 4175 1900 4195 2000
rect 4235 1900 4255 2000
rect 4295 1900 4315 2000
rect 4355 1900 4375 2000
rect 4415 1900 4435 2000
rect 4475 1900 4495 2000
rect 4535 1900 4555 2000
rect 4595 1900 4615 2000
rect 4655 1900 4675 2000
rect 4715 1900 4735 2000
rect 4775 1900 4795 2000
rect 4835 1900 4855 2000
rect 4895 1900 4915 2000
rect 4955 1900 4975 2000
rect 5015 1900 5035 2000
rect 5075 1900 5095 2000
rect 5135 1900 5155 2000
rect 5195 1900 5215 2000
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4235 1615 4255 1665
rect 4295 1615 4315 1665
rect 4355 1615 4375 1665
rect 4415 1615 4435 1665
rect 4475 1615 4495 1665
rect 4535 1615 4555 1665
rect 4595 1615 4615 1665
rect 4655 1615 4675 1665
rect 4715 1615 4735 1665
rect 4775 1615 4795 1665
rect 2875 1210 3375 1460
rect 3415 1210 3915 1460
rect 4085 1210 4585 1460
rect 4625 1210 5125 1460
rect 2980 980 3980 1080
rect 4020 980 5020 1080
rect 3030 785 3080 885
rect 3120 785 3170 885
rect 3210 785 3260 885
rect 3300 785 3350 885
rect 3390 785 3440 885
rect 3480 785 3530 885
rect 3570 785 3620 885
rect 3660 785 3710 885
rect 3750 785 3800 885
rect 3840 785 3890 885
rect 3930 785 3980 885
rect 4020 785 4070 885
rect 4110 785 4160 885
rect 4200 785 4250 885
rect 4290 785 4340 885
rect 4380 785 4430 885
rect 4470 785 4520 885
rect 4560 785 4610 885
rect 4650 785 4700 885
rect 4740 785 4790 885
rect 4830 785 4880 885
rect 4920 785 4970 885
<< ndiff >>
rect 2990 2915 3030 2930
rect 2990 2895 3000 2915
rect 3020 2895 3030 2915
rect 2990 2865 3030 2895
rect 2990 2845 3000 2865
rect 3020 2845 3030 2865
rect 2990 2830 3030 2845
rect 3080 2915 3120 2930
rect 3080 2895 3090 2915
rect 3110 2895 3120 2915
rect 3080 2865 3120 2895
rect 3080 2845 3090 2865
rect 3110 2845 3120 2865
rect 3080 2830 3120 2845
rect 3170 2915 3210 2930
rect 3170 2895 3180 2915
rect 3200 2895 3210 2915
rect 3170 2865 3210 2895
rect 3170 2845 3180 2865
rect 3200 2845 3210 2865
rect 3170 2830 3210 2845
rect 3260 2915 3300 2930
rect 3260 2895 3270 2915
rect 3290 2895 3300 2915
rect 3260 2865 3300 2895
rect 3260 2845 3270 2865
rect 3290 2845 3300 2865
rect 3260 2830 3300 2845
rect 3350 2915 3390 2930
rect 3350 2895 3360 2915
rect 3380 2895 3390 2915
rect 3350 2865 3390 2895
rect 3350 2845 3360 2865
rect 3380 2845 3390 2865
rect 3350 2830 3390 2845
rect 3440 2915 3480 2930
rect 3440 2895 3450 2915
rect 3470 2895 3480 2915
rect 3440 2865 3480 2895
rect 3440 2845 3450 2865
rect 3470 2845 3480 2865
rect 3440 2830 3480 2845
rect 3530 2915 3570 2930
rect 3530 2895 3540 2915
rect 3560 2895 3570 2915
rect 3530 2865 3570 2895
rect 3530 2845 3540 2865
rect 3560 2845 3570 2865
rect 3530 2830 3570 2845
rect 3620 2915 3660 2930
rect 3620 2895 3630 2915
rect 3650 2895 3660 2915
rect 3620 2865 3660 2895
rect 3620 2845 3630 2865
rect 3650 2845 3660 2865
rect 3620 2830 3660 2845
rect 3710 2915 3750 2930
rect 3710 2895 3720 2915
rect 3740 2895 3750 2915
rect 3710 2865 3750 2895
rect 3710 2845 3720 2865
rect 3740 2845 3750 2865
rect 3710 2830 3750 2845
rect 3800 2915 3840 2930
rect 3800 2895 3810 2915
rect 3830 2895 3840 2915
rect 3800 2865 3840 2895
rect 3800 2845 3810 2865
rect 3830 2845 3840 2865
rect 3800 2830 3840 2845
rect 3890 2915 3930 2930
rect 3890 2895 3900 2915
rect 3920 2895 3930 2915
rect 3890 2865 3930 2895
rect 3890 2845 3900 2865
rect 3920 2845 3930 2865
rect 3890 2830 3930 2845
rect 3980 2915 4020 2930
rect 3980 2895 3990 2915
rect 4010 2895 4020 2915
rect 3980 2865 4020 2895
rect 3980 2845 3990 2865
rect 4010 2845 4020 2865
rect 3980 2830 4020 2845
rect 4070 2915 4110 2930
rect 4070 2895 4080 2915
rect 4100 2895 4110 2915
rect 4070 2865 4110 2895
rect 4070 2845 4080 2865
rect 4100 2845 4110 2865
rect 4070 2830 4110 2845
rect 4160 2915 4200 2930
rect 4160 2895 4170 2915
rect 4190 2895 4200 2915
rect 4160 2865 4200 2895
rect 4160 2845 4170 2865
rect 4190 2845 4200 2865
rect 4160 2830 4200 2845
rect 4250 2915 4290 2930
rect 4250 2895 4260 2915
rect 4280 2895 4290 2915
rect 4250 2865 4290 2895
rect 4250 2845 4260 2865
rect 4280 2845 4290 2865
rect 4250 2830 4290 2845
rect 4340 2915 4380 2930
rect 4340 2895 4350 2915
rect 4370 2895 4380 2915
rect 4340 2865 4380 2895
rect 4340 2845 4350 2865
rect 4370 2845 4380 2865
rect 4340 2830 4380 2845
rect 4430 2915 4470 2930
rect 4430 2895 4440 2915
rect 4460 2895 4470 2915
rect 4430 2865 4470 2895
rect 4430 2845 4440 2865
rect 4460 2845 4470 2865
rect 4430 2830 4470 2845
rect 4520 2915 4560 2930
rect 4520 2895 4530 2915
rect 4550 2895 4560 2915
rect 4520 2865 4560 2895
rect 4520 2845 4530 2865
rect 4550 2845 4560 2865
rect 4520 2830 4560 2845
rect 4610 2915 4650 2930
rect 4610 2895 4620 2915
rect 4640 2895 4650 2915
rect 4610 2865 4650 2895
rect 4610 2845 4620 2865
rect 4640 2845 4650 2865
rect 4610 2830 4650 2845
rect 4700 2915 4740 2930
rect 4700 2895 4710 2915
rect 4730 2895 4740 2915
rect 4700 2865 4740 2895
rect 4700 2845 4710 2865
rect 4730 2845 4740 2865
rect 4700 2830 4740 2845
rect 4790 2915 4830 2930
rect 4790 2895 4800 2915
rect 4820 2895 4830 2915
rect 4790 2865 4830 2895
rect 4790 2845 4800 2865
rect 4820 2845 4830 2865
rect 4790 2830 4830 2845
rect 4880 2915 4920 2930
rect 4880 2895 4890 2915
rect 4910 2895 4920 2915
rect 4880 2865 4920 2895
rect 4880 2845 4890 2865
rect 4910 2845 4920 2865
rect 4880 2830 4920 2845
rect 4970 2915 5010 2930
rect 4970 2895 4980 2915
rect 5000 2895 5010 2915
rect 4970 2865 5010 2895
rect 4970 2845 4980 2865
rect 5000 2845 5010 2865
rect 4970 2830 5010 2845
rect 2810 2685 2850 2700
rect 2810 2665 2820 2685
rect 2840 2665 2850 2685
rect 2810 2635 2850 2665
rect 2810 2615 2820 2635
rect 2840 2615 2850 2635
rect 2810 2585 2850 2615
rect 2810 2565 2820 2585
rect 2840 2565 2850 2585
rect 2810 2535 2850 2565
rect 2810 2515 2820 2535
rect 2840 2515 2850 2535
rect 2810 2485 2850 2515
rect 2810 2465 2820 2485
rect 2840 2465 2850 2485
rect 2810 2435 2850 2465
rect 2810 2415 2820 2435
rect 2840 2415 2850 2435
rect 2810 2400 2850 2415
rect 2900 2685 2940 2700
rect 2900 2665 2910 2685
rect 2930 2665 2940 2685
rect 2900 2635 2940 2665
rect 2900 2615 2910 2635
rect 2930 2615 2940 2635
rect 2900 2585 2940 2615
rect 2900 2565 2910 2585
rect 2930 2565 2940 2585
rect 2900 2535 2940 2565
rect 2900 2515 2910 2535
rect 2930 2515 2940 2535
rect 2900 2485 2940 2515
rect 2900 2465 2910 2485
rect 2930 2465 2940 2485
rect 2900 2435 2940 2465
rect 2900 2415 2910 2435
rect 2930 2415 2940 2435
rect 2900 2400 2940 2415
rect 2990 2685 3030 2700
rect 2990 2665 3000 2685
rect 3020 2665 3030 2685
rect 2990 2635 3030 2665
rect 2990 2615 3000 2635
rect 3020 2615 3030 2635
rect 2990 2585 3030 2615
rect 2990 2565 3000 2585
rect 3020 2565 3030 2585
rect 2990 2535 3030 2565
rect 2990 2515 3000 2535
rect 3020 2515 3030 2535
rect 2990 2485 3030 2515
rect 2990 2465 3000 2485
rect 3020 2465 3030 2485
rect 2990 2435 3030 2465
rect 2990 2415 3000 2435
rect 3020 2415 3030 2435
rect 2990 2400 3030 2415
rect 3080 2685 3120 2700
rect 3080 2665 3090 2685
rect 3110 2665 3120 2685
rect 3080 2635 3120 2665
rect 3080 2615 3090 2635
rect 3110 2615 3120 2635
rect 3080 2585 3120 2615
rect 3080 2565 3090 2585
rect 3110 2565 3120 2585
rect 3080 2535 3120 2565
rect 3080 2515 3090 2535
rect 3110 2515 3120 2535
rect 3080 2485 3120 2515
rect 3080 2465 3090 2485
rect 3110 2465 3120 2485
rect 3080 2435 3120 2465
rect 3080 2415 3090 2435
rect 3110 2415 3120 2435
rect 3080 2400 3120 2415
rect 3170 2685 3210 2700
rect 3170 2665 3180 2685
rect 3200 2665 3210 2685
rect 3170 2635 3210 2665
rect 3170 2615 3180 2635
rect 3200 2615 3210 2635
rect 3170 2585 3210 2615
rect 3170 2565 3180 2585
rect 3200 2565 3210 2585
rect 3170 2535 3210 2565
rect 3170 2515 3180 2535
rect 3200 2515 3210 2535
rect 3170 2485 3210 2515
rect 3170 2465 3180 2485
rect 3200 2465 3210 2485
rect 3170 2435 3210 2465
rect 3170 2415 3180 2435
rect 3200 2415 3210 2435
rect 3170 2400 3210 2415
rect 3260 2685 3300 2700
rect 3260 2665 3270 2685
rect 3290 2665 3300 2685
rect 3260 2635 3300 2665
rect 3260 2615 3270 2635
rect 3290 2615 3300 2635
rect 3260 2585 3300 2615
rect 3260 2565 3270 2585
rect 3290 2565 3300 2585
rect 3260 2535 3300 2565
rect 3260 2515 3270 2535
rect 3290 2515 3300 2535
rect 3260 2485 3300 2515
rect 3260 2465 3270 2485
rect 3290 2465 3300 2485
rect 3260 2435 3300 2465
rect 3260 2415 3270 2435
rect 3290 2415 3300 2435
rect 3260 2400 3300 2415
rect 3350 2685 3390 2700
rect 3350 2665 3360 2685
rect 3380 2665 3390 2685
rect 3350 2635 3390 2665
rect 3350 2615 3360 2635
rect 3380 2615 3390 2635
rect 3350 2585 3390 2615
rect 3350 2565 3360 2585
rect 3380 2565 3390 2585
rect 3350 2535 3390 2565
rect 3350 2515 3360 2535
rect 3380 2515 3390 2535
rect 3350 2485 3390 2515
rect 3350 2465 3360 2485
rect 3380 2465 3390 2485
rect 3350 2435 3390 2465
rect 3350 2415 3360 2435
rect 3380 2415 3390 2435
rect 3350 2400 3390 2415
rect 3440 2685 3480 2700
rect 3440 2665 3450 2685
rect 3470 2665 3480 2685
rect 3440 2635 3480 2665
rect 3440 2615 3450 2635
rect 3470 2615 3480 2635
rect 3440 2585 3480 2615
rect 3440 2565 3450 2585
rect 3470 2565 3480 2585
rect 3440 2535 3480 2565
rect 3440 2515 3450 2535
rect 3470 2515 3480 2535
rect 3440 2485 3480 2515
rect 3440 2465 3450 2485
rect 3470 2465 3480 2485
rect 3440 2435 3480 2465
rect 3440 2415 3450 2435
rect 3470 2415 3480 2435
rect 3440 2400 3480 2415
rect 3530 2685 3570 2700
rect 3530 2665 3540 2685
rect 3560 2665 3570 2685
rect 3530 2635 3570 2665
rect 3530 2615 3540 2635
rect 3560 2615 3570 2635
rect 3530 2585 3570 2615
rect 3530 2565 3540 2585
rect 3560 2565 3570 2585
rect 3530 2535 3570 2565
rect 3530 2515 3540 2535
rect 3560 2515 3570 2535
rect 3530 2485 3570 2515
rect 3530 2465 3540 2485
rect 3560 2465 3570 2485
rect 3530 2435 3570 2465
rect 3530 2415 3540 2435
rect 3560 2415 3570 2435
rect 3530 2400 3570 2415
rect 3620 2685 3660 2700
rect 3620 2665 3630 2685
rect 3650 2665 3660 2685
rect 3620 2635 3660 2665
rect 3620 2615 3630 2635
rect 3650 2615 3660 2635
rect 3620 2585 3660 2615
rect 3620 2565 3630 2585
rect 3650 2565 3660 2585
rect 3620 2535 3660 2565
rect 3620 2515 3630 2535
rect 3650 2515 3660 2535
rect 3620 2485 3660 2515
rect 3620 2465 3630 2485
rect 3650 2465 3660 2485
rect 3620 2435 3660 2465
rect 3620 2415 3630 2435
rect 3650 2415 3660 2435
rect 3620 2400 3660 2415
rect 3710 2685 3750 2700
rect 3710 2665 3720 2685
rect 3740 2665 3750 2685
rect 3710 2635 3750 2665
rect 3710 2615 3720 2635
rect 3740 2615 3750 2635
rect 3710 2585 3750 2615
rect 3710 2565 3720 2585
rect 3740 2565 3750 2585
rect 3710 2535 3750 2565
rect 3710 2515 3720 2535
rect 3740 2515 3750 2535
rect 3710 2485 3750 2515
rect 3710 2465 3720 2485
rect 3740 2465 3750 2485
rect 3710 2435 3750 2465
rect 3710 2415 3720 2435
rect 3740 2415 3750 2435
rect 3710 2400 3750 2415
rect 3800 2685 3840 2700
rect 3800 2665 3810 2685
rect 3830 2665 3840 2685
rect 3800 2635 3840 2665
rect 3800 2615 3810 2635
rect 3830 2615 3840 2635
rect 3800 2585 3840 2615
rect 3800 2565 3810 2585
rect 3830 2565 3840 2585
rect 3800 2535 3840 2565
rect 3800 2515 3810 2535
rect 3830 2515 3840 2535
rect 3800 2485 3840 2515
rect 3800 2465 3810 2485
rect 3830 2465 3840 2485
rect 3800 2435 3840 2465
rect 3800 2415 3810 2435
rect 3830 2415 3840 2435
rect 3800 2400 3840 2415
rect 3890 2685 3930 2700
rect 3890 2665 3900 2685
rect 3920 2665 3930 2685
rect 3890 2635 3930 2665
rect 3890 2615 3900 2635
rect 3920 2615 3930 2635
rect 3890 2585 3930 2615
rect 3890 2565 3900 2585
rect 3920 2565 3930 2585
rect 3890 2535 3930 2565
rect 3890 2515 3900 2535
rect 3920 2515 3930 2535
rect 3890 2485 3930 2515
rect 3890 2465 3900 2485
rect 3920 2465 3930 2485
rect 3890 2435 3930 2465
rect 3890 2415 3900 2435
rect 3920 2415 3930 2435
rect 3890 2400 3930 2415
rect 3980 2685 4020 2700
rect 3980 2665 3990 2685
rect 4010 2665 4020 2685
rect 3980 2635 4020 2665
rect 3980 2615 3990 2635
rect 4010 2615 4020 2635
rect 3980 2585 4020 2615
rect 3980 2565 3990 2585
rect 4010 2565 4020 2585
rect 3980 2535 4020 2565
rect 3980 2515 3990 2535
rect 4010 2515 4020 2535
rect 3980 2485 4020 2515
rect 3980 2465 3990 2485
rect 4010 2465 4020 2485
rect 3980 2435 4020 2465
rect 3980 2415 3990 2435
rect 4010 2415 4020 2435
rect 3980 2400 4020 2415
rect 4070 2685 4110 2700
rect 4070 2665 4080 2685
rect 4100 2665 4110 2685
rect 4070 2635 4110 2665
rect 4070 2615 4080 2635
rect 4100 2615 4110 2635
rect 4070 2585 4110 2615
rect 4070 2565 4080 2585
rect 4100 2565 4110 2585
rect 4070 2535 4110 2565
rect 4070 2515 4080 2535
rect 4100 2515 4110 2535
rect 4070 2485 4110 2515
rect 4070 2465 4080 2485
rect 4100 2465 4110 2485
rect 4070 2435 4110 2465
rect 4070 2415 4080 2435
rect 4100 2415 4110 2435
rect 4070 2400 4110 2415
rect 4160 2685 4200 2700
rect 4160 2665 4170 2685
rect 4190 2665 4200 2685
rect 4160 2635 4200 2665
rect 4160 2615 4170 2635
rect 4190 2615 4200 2635
rect 4160 2585 4200 2615
rect 4160 2565 4170 2585
rect 4190 2565 4200 2585
rect 4160 2535 4200 2565
rect 4160 2515 4170 2535
rect 4190 2515 4200 2535
rect 4160 2485 4200 2515
rect 4160 2465 4170 2485
rect 4190 2465 4200 2485
rect 4160 2435 4200 2465
rect 4160 2415 4170 2435
rect 4190 2415 4200 2435
rect 4160 2400 4200 2415
rect 4250 2685 4290 2700
rect 4250 2665 4260 2685
rect 4280 2665 4290 2685
rect 4250 2635 4290 2665
rect 4250 2615 4260 2635
rect 4280 2615 4290 2635
rect 4250 2585 4290 2615
rect 4250 2565 4260 2585
rect 4280 2565 4290 2585
rect 4250 2535 4290 2565
rect 4250 2515 4260 2535
rect 4280 2515 4290 2535
rect 4250 2485 4290 2515
rect 4250 2465 4260 2485
rect 4280 2465 4290 2485
rect 4250 2435 4290 2465
rect 4250 2415 4260 2435
rect 4280 2415 4290 2435
rect 4250 2400 4290 2415
rect 4340 2685 4380 2700
rect 4340 2665 4350 2685
rect 4370 2665 4380 2685
rect 4340 2635 4380 2665
rect 4340 2615 4350 2635
rect 4370 2615 4380 2635
rect 4340 2585 4380 2615
rect 4340 2565 4350 2585
rect 4370 2565 4380 2585
rect 4340 2535 4380 2565
rect 4340 2515 4350 2535
rect 4370 2515 4380 2535
rect 4340 2485 4380 2515
rect 4340 2465 4350 2485
rect 4370 2465 4380 2485
rect 4340 2435 4380 2465
rect 4340 2415 4350 2435
rect 4370 2415 4380 2435
rect 4340 2400 4380 2415
rect 4430 2685 4470 2700
rect 4430 2665 4440 2685
rect 4460 2665 4470 2685
rect 4430 2635 4470 2665
rect 4430 2615 4440 2635
rect 4460 2615 4470 2635
rect 4430 2585 4470 2615
rect 4430 2565 4440 2585
rect 4460 2565 4470 2585
rect 4430 2535 4470 2565
rect 4430 2515 4440 2535
rect 4460 2515 4470 2535
rect 4430 2485 4470 2515
rect 4430 2465 4440 2485
rect 4460 2465 4470 2485
rect 4430 2435 4470 2465
rect 4430 2415 4440 2435
rect 4460 2415 4470 2435
rect 4430 2400 4470 2415
rect 4520 2685 4560 2700
rect 4520 2665 4530 2685
rect 4550 2665 4560 2685
rect 4520 2635 4560 2665
rect 4520 2615 4530 2635
rect 4550 2615 4560 2635
rect 4520 2585 4560 2615
rect 4520 2565 4530 2585
rect 4550 2565 4560 2585
rect 4520 2535 4560 2565
rect 4520 2515 4530 2535
rect 4550 2515 4560 2535
rect 4520 2485 4560 2515
rect 4520 2465 4530 2485
rect 4550 2465 4560 2485
rect 4520 2435 4560 2465
rect 4520 2415 4530 2435
rect 4550 2415 4560 2435
rect 4520 2400 4560 2415
rect 4610 2685 4650 2700
rect 4610 2665 4620 2685
rect 4640 2665 4650 2685
rect 4610 2635 4650 2665
rect 4610 2615 4620 2635
rect 4640 2615 4650 2635
rect 4610 2585 4650 2615
rect 4610 2565 4620 2585
rect 4640 2565 4650 2585
rect 4610 2535 4650 2565
rect 4610 2515 4620 2535
rect 4640 2515 4650 2535
rect 4610 2485 4650 2515
rect 4610 2465 4620 2485
rect 4640 2465 4650 2485
rect 4610 2435 4650 2465
rect 4610 2415 4620 2435
rect 4640 2415 4650 2435
rect 4610 2400 4650 2415
rect 4700 2685 4740 2700
rect 4700 2665 4710 2685
rect 4730 2665 4740 2685
rect 4700 2635 4740 2665
rect 4700 2615 4710 2635
rect 4730 2615 4740 2635
rect 4700 2585 4740 2615
rect 4700 2565 4710 2585
rect 4730 2565 4740 2585
rect 4700 2535 4740 2565
rect 4700 2515 4710 2535
rect 4730 2515 4740 2535
rect 4700 2485 4740 2515
rect 4700 2465 4710 2485
rect 4730 2465 4740 2485
rect 4700 2435 4740 2465
rect 4700 2415 4710 2435
rect 4730 2415 4740 2435
rect 4700 2400 4740 2415
rect 4790 2685 4830 2700
rect 4790 2665 4800 2685
rect 4820 2665 4830 2685
rect 4790 2635 4830 2665
rect 4790 2615 4800 2635
rect 4820 2615 4830 2635
rect 4790 2585 4830 2615
rect 4790 2565 4800 2585
rect 4820 2565 4830 2585
rect 4790 2535 4830 2565
rect 4790 2515 4800 2535
rect 4820 2515 4830 2535
rect 4790 2485 4830 2515
rect 4790 2465 4800 2485
rect 4820 2465 4830 2485
rect 4790 2435 4830 2465
rect 4790 2415 4800 2435
rect 4820 2415 4830 2435
rect 4790 2400 4830 2415
rect 4880 2685 4920 2700
rect 4880 2665 4890 2685
rect 4910 2665 4920 2685
rect 4880 2635 4920 2665
rect 4880 2615 4890 2635
rect 4910 2615 4920 2635
rect 4880 2585 4920 2615
rect 4880 2565 4890 2585
rect 4910 2565 4920 2585
rect 4880 2535 4920 2565
rect 4880 2515 4890 2535
rect 4910 2515 4920 2535
rect 4880 2485 4920 2515
rect 4880 2465 4890 2485
rect 4910 2465 4920 2485
rect 4880 2435 4920 2465
rect 4880 2415 4890 2435
rect 4910 2415 4920 2435
rect 4880 2400 4920 2415
rect 4970 2685 5010 2700
rect 4970 2665 4980 2685
rect 5000 2665 5010 2685
rect 4970 2635 5010 2665
rect 4970 2615 4980 2635
rect 5000 2615 5010 2635
rect 4970 2585 5010 2615
rect 4970 2565 4980 2585
rect 5000 2565 5010 2585
rect 4970 2535 5010 2565
rect 4970 2515 4980 2535
rect 5000 2515 5010 2535
rect 4970 2485 5010 2515
rect 4970 2465 4980 2485
rect 5000 2465 5010 2485
rect 4970 2435 5010 2465
rect 4970 2415 4980 2435
rect 5000 2415 5010 2435
rect 4970 2400 5010 2415
rect 5060 2685 5100 2700
rect 5060 2665 5070 2685
rect 5090 2665 5100 2685
rect 5060 2635 5100 2665
rect 5060 2615 5070 2635
rect 5090 2615 5100 2635
rect 5060 2585 5100 2615
rect 5060 2565 5070 2585
rect 5090 2565 5100 2585
rect 5060 2535 5100 2565
rect 5060 2515 5070 2535
rect 5090 2515 5100 2535
rect 5060 2485 5100 2515
rect 5060 2465 5070 2485
rect 5090 2465 5100 2485
rect 5060 2435 5100 2465
rect 5060 2415 5070 2435
rect 5090 2415 5100 2435
rect 5060 2400 5100 2415
rect 5150 2685 5190 2700
rect 5150 2665 5160 2685
rect 5180 2665 5190 2685
rect 5150 2635 5190 2665
rect 5150 2615 5160 2635
rect 5180 2615 5190 2635
rect 5150 2585 5190 2615
rect 5150 2565 5160 2585
rect 5180 2565 5190 2585
rect 5150 2535 5190 2565
rect 5150 2515 5160 2535
rect 5180 2515 5190 2535
rect 5150 2485 5190 2515
rect 5150 2465 5160 2485
rect 5180 2465 5190 2485
rect 5150 2435 5190 2465
rect 5150 2415 5160 2435
rect 5180 2415 5190 2435
rect 5150 2400 5190 2415
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 3945 1935 3985 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 3945 1900 3985 1915
rect 4015 1985 4055 2000
rect 4015 1965 4025 1985
rect 4045 1965 4055 1985
rect 4015 1935 4055 1965
rect 4015 1915 4025 1935
rect 4045 1915 4055 1935
rect 4015 1900 4055 1915
rect 4075 1985 4115 2000
rect 4075 1965 4085 1985
rect 4105 1965 4115 1985
rect 4075 1935 4115 1965
rect 4075 1915 4085 1935
rect 4105 1915 4115 1935
rect 4075 1900 4115 1915
rect 4135 1985 4175 2000
rect 4135 1965 4145 1985
rect 4165 1965 4175 1985
rect 4135 1935 4175 1965
rect 4135 1915 4145 1935
rect 4165 1915 4175 1935
rect 4135 1900 4175 1915
rect 4195 1985 4235 2000
rect 4195 1965 4205 1985
rect 4225 1965 4235 1985
rect 4195 1935 4235 1965
rect 4195 1915 4205 1935
rect 4225 1915 4235 1935
rect 4195 1900 4235 1915
rect 4255 1985 4295 2000
rect 4255 1965 4265 1985
rect 4285 1965 4295 1985
rect 4255 1935 4295 1965
rect 4255 1915 4265 1935
rect 4285 1915 4295 1935
rect 4255 1900 4295 1915
rect 4315 1985 4355 2000
rect 4315 1965 4325 1985
rect 4345 1965 4355 1985
rect 4315 1935 4355 1965
rect 4315 1915 4325 1935
rect 4345 1915 4355 1935
rect 4315 1900 4355 1915
rect 4375 1985 4415 2000
rect 4375 1965 4385 1985
rect 4405 1965 4415 1985
rect 4375 1935 4415 1965
rect 4375 1915 4385 1935
rect 4405 1915 4415 1935
rect 4375 1900 4415 1915
rect 4435 1985 4475 2000
rect 4435 1965 4445 1985
rect 4465 1965 4475 1985
rect 4435 1935 4475 1965
rect 4435 1915 4445 1935
rect 4465 1915 4475 1935
rect 4435 1900 4475 1915
rect 4495 1985 4535 2000
rect 4495 1965 4505 1985
rect 4525 1965 4535 1985
rect 4495 1935 4535 1965
rect 4495 1915 4505 1935
rect 4525 1915 4535 1935
rect 4495 1900 4535 1915
rect 4555 1985 4595 2000
rect 4555 1965 4565 1985
rect 4585 1965 4595 1985
rect 4555 1935 4595 1965
rect 4555 1915 4565 1935
rect 4585 1915 4595 1935
rect 4555 1900 4595 1915
rect 4615 1985 4655 2000
rect 4615 1965 4625 1985
rect 4645 1965 4655 1985
rect 4615 1935 4655 1965
rect 4615 1915 4625 1935
rect 4645 1915 4655 1935
rect 4615 1900 4655 1915
rect 4675 1985 4715 2000
rect 4675 1965 4685 1985
rect 4705 1965 4715 1985
rect 4675 1935 4715 1965
rect 4675 1915 4685 1935
rect 4705 1915 4715 1935
rect 4675 1900 4715 1915
rect 4735 1985 4775 2000
rect 4735 1965 4745 1985
rect 4765 1965 4775 1985
rect 4735 1935 4775 1965
rect 4735 1915 4745 1935
rect 4765 1915 4775 1935
rect 4735 1900 4775 1915
rect 4795 1985 4835 2000
rect 4795 1965 4805 1985
rect 4825 1965 4835 1985
rect 4795 1935 4835 1965
rect 4795 1915 4805 1935
rect 4825 1915 4835 1935
rect 4795 1900 4835 1915
rect 4855 1985 4895 2000
rect 4855 1965 4865 1985
rect 4885 1965 4895 1985
rect 4855 1935 4895 1965
rect 4855 1915 4865 1935
rect 4885 1915 4895 1935
rect 4855 1900 4895 1915
rect 4915 1985 4955 2000
rect 4915 1965 4925 1985
rect 4945 1965 4955 1985
rect 4915 1935 4955 1965
rect 4915 1915 4925 1935
rect 4945 1915 4955 1935
rect 4915 1900 4955 1915
rect 4975 1985 5015 2000
rect 4975 1965 4985 1985
rect 5005 1965 5015 1985
rect 4975 1935 5015 1965
rect 4975 1915 4985 1935
rect 5005 1915 5015 1935
rect 4975 1900 5015 1915
rect 5035 1985 5075 2000
rect 5035 1965 5045 1985
rect 5065 1965 5075 1985
rect 5035 1935 5075 1965
rect 5035 1915 5045 1935
rect 5065 1915 5075 1935
rect 5035 1900 5075 1915
rect 5095 1985 5135 2000
rect 5095 1965 5105 1985
rect 5125 1965 5135 1985
rect 5095 1935 5135 1965
rect 5095 1915 5105 1935
rect 5125 1915 5135 1935
rect 5095 1900 5135 1915
rect 5155 1985 5195 2000
rect 5155 1965 5165 1985
rect 5185 1965 5195 1985
rect 5155 1935 5195 1965
rect 5155 1915 5165 1935
rect 5185 1915 5195 1935
rect 5155 1900 5195 1915
rect 5215 1985 5255 2000
rect 5215 1965 5225 1985
rect 5245 1965 5255 1985
rect 5215 1935 5255 1965
rect 5215 1915 5225 1935
rect 5245 1915 5255 1935
rect 5215 1900 5255 1915
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4195 1650 4235 1665
rect 4195 1630 4205 1650
rect 4225 1630 4235 1650
rect 4195 1615 4235 1630
rect 4255 1650 4295 1665
rect 4255 1630 4265 1650
rect 4285 1630 4295 1650
rect 4255 1615 4295 1630
rect 4315 1650 4355 1665
rect 4315 1630 4325 1650
rect 4345 1630 4355 1650
rect 4315 1615 4355 1630
rect 4375 1650 4415 1665
rect 4375 1630 4385 1650
rect 4405 1630 4415 1650
rect 4375 1615 4415 1630
rect 4435 1650 4475 1665
rect 4435 1630 4445 1650
rect 4465 1630 4475 1650
rect 4435 1615 4475 1630
rect 4495 1650 4535 1665
rect 4495 1630 4505 1650
rect 4525 1630 4535 1650
rect 4495 1615 4535 1630
rect 4555 1650 4595 1665
rect 4555 1630 4565 1650
rect 4585 1630 4595 1650
rect 4555 1615 4595 1630
rect 4615 1650 4655 1665
rect 4615 1630 4625 1650
rect 4645 1630 4655 1650
rect 4615 1615 4655 1630
rect 4675 1650 4715 1665
rect 4675 1630 4685 1650
rect 4705 1630 4715 1650
rect 4675 1615 4715 1630
rect 4735 1650 4775 1665
rect 4735 1630 4745 1650
rect 4765 1630 4775 1650
rect 4735 1615 4775 1630
rect 4795 1650 4835 1665
rect 4795 1630 4805 1650
rect 4825 1630 4835 1650
rect 4795 1615 4835 1630
rect 2835 1445 2875 1460
rect 2835 1425 2845 1445
rect 2865 1425 2875 1445
rect 2835 1395 2875 1425
rect 2835 1375 2845 1395
rect 2865 1375 2875 1395
rect 2835 1345 2875 1375
rect 2835 1325 2845 1345
rect 2865 1325 2875 1345
rect 2835 1295 2875 1325
rect 2835 1275 2845 1295
rect 2865 1275 2875 1295
rect 2835 1245 2875 1275
rect 2835 1225 2845 1245
rect 2865 1225 2875 1245
rect 2835 1210 2875 1225
rect 3375 1445 3415 1460
rect 3375 1425 3385 1445
rect 3405 1425 3415 1445
rect 3375 1395 3415 1425
rect 3375 1375 3385 1395
rect 3405 1375 3415 1395
rect 3375 1345 3415 1375
rect 3375 1325 3385 1345
rect 3405 1325 3415 1345
rect 3375 1295 3415 1325
rect 3375 1275 3385 1295
rect 3405 1275 3415 1295
rect 3375 1245 3415 1275
rect 3375 1225 3385 1245
rect 3405 1225 3415 1245
rect 3375 1210 3415 1225
rect 3915 1445 3955 1460
rect 3915 1425 3925 1445
rect 3945 1425 3955 1445
rect 3915 1395 3955 1425
rect 3915 1375 3925 1395
rect 3945 1375 3955 1395
rect 3915 1345 3955 1375
rect 3915 1325 3925 1345
rect 3945 1325 3955 1345
rect 3915 1295 3955 1325
rect 3915 1275 3925 1295
rect 3945 1275 3955 1295
rect 3915 1245 3955 1275
rect 3915 1225 3925 1245
rect 3945 1225 3955 1245
rect 3915 1210 3955 1225
rect 4045 1445 4085 1460
rect 4045 1425 4055 1445
rect 4075 1425 4085 1445
rect 4045 1395 4085 1425
rect 4045 1375 4055 1395
rect 4075 1375 4085 1395
rect 4045 1345 4085 1375
rect 4045 1325 4055 1345
rect 4075 1325 4085 1345
rect 4045 1295 4085 1325
rect 4045 1275 4055 1295
rect 4075 1275 4085 1295
rect 4045 1245 4085 1275
rect 4045 1225 4055 1245
rect 4075 1225 4085 1245
rect 4045 1210 4085 1225
rect 4585 1445 4625 1460
rect 4585 1425 4595 1445
rect 4615 1425 4625 1445
rect 4585 1395 4625 1425
rect 4585 1375 4595 1395
rect 4615 1375 4625 1395
rect 4585 1345 4625 1375
rect 4585 1325 4595 1345
rect 4615 1325 4625 1345
rect 4585 1295 4625 1325
rect 4585 1275 4595 1295
rect 4615 1275 4625 1295
rect 4585 1245 4625 1275
rect 4585 1225 4595 1245
rect 4615 1225 4625 1245
rect 4585 1210 4625 1225
rect 5125 1445 5165 1460
rect 5125 1425 5135 1445
rect 5155 1425 5165 1445
rect 5125 1395 5165 1425
rect 5125 1375 5135 1395
rect 5155 1375 5165 1395
rect 5125 1345 5165 1375
rect 5125 1325 5135 1345
rect 5155 1325 5165 1345
rect 5125 1295 5165 1325
rect 5125 1275 5135 1295
rect 5155 1275 5165 1295
rect 5125 1245 5165 1275
rect 5125 1225 5135 1245
rect 5155 1225 5165 1245
rect 5125 1210 5165 1225
rect 2940 1065 2980 1080
rect 2940 1045 2950 1065
rect 2970 1045 2980 1065
rect 2940 1015 2980 1045
rect 2940 995 2950 1015
rect 2970 995 2980 1015
rect 2940 980 2980 995
rect 3980 1065 4020 1080
rect 3980 1045 3990 1065
rect 4010 1045 4020 1065
rect 3980 1015 4020 1045
rect 3980 995 3990 1015
rect 4010 995 4020 1015
rect 3980 980 4020 995
rect 5020 1065 5060 1080
rect 5020 1045 5030 1065
rect 5050 1045 5060 1065
rect 5020 1015 5060 1045
rect 5020 995 5030 1015
rect 5050 995 5060 1015
rect 5020 980 5060 995
rect 2990 870 3030 885
rect 2990 850 3000 870
rect 3020 850 3030 870
rect 2990 820 3030 850
rect 2990 800 3000 820
rect 3020 800 3030 820
rect 2990 785 3030 800
rect 3080 870 3120 885
rect 3080 850 3090 870
rect 3110 850 3120 870
rect 3080 820 3120 850
rect 3080 800 3090 820
rect 3110 800 3120 820
rect 3080 785 3120 800
rect 3170 870 3210 885
rect 3170 850 3180 870
rect 3200 850 3210 870
rect 3170 820 3210 850
rect 3170 800 3180 820
rect 3200 800 3210 820
rect 3170 785 3210 800
rect 3260 870 3300 885
rect 3260 850 3270 870
rect 3290 850 3300 870
rect 3260 820 3300 850
rect 3260 800 3270 820
rect 3290 800 3300 820
rect 3260 785 3300 800
rect 3350 870 3390 885
rect 3350 850 3360 870
rect 3380 850 3390 870
rect 3350 820 3390 850
rect 3350 800 3360 820
rect 3380 800 3390 820
rect 3350 785 3390 800
rect 3440 870 3480 885
rect 3440 850 3450 870
rect 3470 850 3480 870
rect 3440 820 3480 850
rect 3440 800 3450 820
rect 3470 800 3480 820
rect 3440 785 3480 800
rect 3530 870 3570 885
rect 3530 850 3540 870
rect 3560 850 3570 870
rect 3530 820 3570 850
rect 3530 800 3540 820
rect 3560 800 3570 820
rect 3530 785 3570 800
rect 3620 870 3660 885
rect 3620 850 3630 870
rect 3650 850 3660 870
rect 3620 820 3660 850
rect 3620 800 3630 820
rect 3650 800 3660 820
rect 3620 785 3660 800
rect 3710 870 3750 885
rect 3710 850 3720 870
rect 3740 850 3750 870
rect 3710 820 3750 850
rect 3710 800 3720 820
rect 3740 800 3750 820
rect 3710 785 3750 800
rect 3800 870 3840 885
rect 3800 850 3810 870
rect 3830 850 3840 870
rect 3800 820 3840 850
rect 3800 800 3810 820
rect 3830 800 3840 820
rect 3800 785 3840 800
rect 3890 870 3930 885
rect 3890 850 3900 870
rect 3920 850 3930 870
rect 3890 820 3930 850
rect 3890 800 3900 820
rect 3920 800 3930 820
rect 3890 785 3930 800
rect 3980 870 4020 885
rect 3980 850 3990 870
rect 4010 850 4020 870
rect 3980 820 4020 850
rect 3980 800 3990 820
rect 4010 800 4020 820
rect 3980 785 4020 800
rect 4070 870 4110 885
rect 4070 850 4080 870
rect 4100 850 4110 870
rect 4070 820 4110 850
rect 4070 800 4080 820
rect 4100 800 4110 820
rect 4070 785 4110 800
rect 4160 870 4200 885
rect 4160 850 4170 870
rect 4190 850 4200 870
rect 4160 820 4200 850
rect 4160 800 4170 820
rect 4190 800 4200 820
rect 4160 785 4200 800
rect 4250 870 4290 885
rect 4250 850 4260 870
rect 4280 850 4290 870
rect 4250 820 4290 850
rect 4250 800 4260 820
rect 4280 800 4290 820
rect 4250 785 4290 800
rect 4340 870 4380 885
rect 4340 850 4350 870
rect 4370 850 4380 870
rect 4340 820 4380 850
rect 4340 800 4350 820
rect 4370 800 4380 820
rect 4340 785 4380 800
rect 4430 870 4470 885
rect 4430 850 4440 870
rect 4460 850 4470 870
rect 4430 820 4470 850
rect 4430 800 4440 820
rect 4460 800 4470 820
rect 4430 785 4470 800
rect 4520 870 4560 885
rect 4520 850 4530 870
rect 4550 850 4560 870
rect 4520 820 4560 850
rect 4520 800 4530 820
rect 4550 800 4560 820
rect 4520 785 4560 800
rect 4610 870 4650 885
rect 4610 850 4620 870
rect 4640 850 4650 870
rect 4610 820 4650 850
rect 4610 800 4620 820
rect 4640 800 4650 820
rect 4610 785 4650 800
rect 4700 870 4740 885
rect 4700 850 4710 870
rect 4730 850 4740 870
rect 4700 820 4740 850
rect 4700 800 4710 820
rect 4730 800 4740 820
rect 4700 785 4740 800
rect 4790 870 4830 885
rect 4790 850 4800 870
rect 4820 850 4830 870
rect 4790 820 4830 850
rect 4790 800 4800 820
rect 4820 800 4830 820
rect 4790 785 4830 800
rect 4880 870 4920 885
rect 4880 850 4890 870
rect 4910 850 4920 870
rect 4880 820 4920 850
rect 4880 800 4890 820
rect 4910 800 4920 820
rect 4880 785 4920 800
rect 4970 870 5010 885
rect 4970 850 4980 870
rect 5000 850 5010 870
rect 4970 820 5010 850
rect 4970 800 4980 820
rect 5000 800 5010 820
rect 4970 785 5010 800
<< ndiffc >>
rect 3000 2895 3020 2915
rect 3000 2845 3020 2865
rect 3090 2895 3110 2915
rect 3090 2845 3110 2865
rect 3180 2895 3200 2915
rect 3180 2845 3200 2865
rect 3270 2895 3290 2915
rect 3270 2845 3290 2865
rect 3360 2895 3380 2915
rect 3360 2845 3380 2865
rect 3450 2895 3470 2915
rect 3450 2845 3470 2865
rect 3540 2895 3560 2915
rect 3540 2845 3560 2865
rect 3630 2895 3650 2915
rect 3630 2845 3650 2865
rect 3720 2895 3740 2915
rect 3720 2845 3740 2865
rect 3810 2895 3830 2915
rect 3810 2845 3830 2865
rect 3900 2895 3920 2915
rect 3900 2845 3920 2865
rect 3990 2895 4010 2915
rect 3990 2845 4010 2865
rect 4080 2895 4100 2915
rect 4080 2845 4100 2865
rect 4170 2895 4190 2915
rect 4170 2845 4190 2865
rect 4260 2895 4280 2915
rect 4260 2845 4280 2865
rect 4350 2895 4370 2915
rect 4350 2845 4370 2865
rect 4440 2895 4460 2915
rect 4440 2845 4460 2865
rect 4530 2895 4550 2915
rect 4530 2845 4550 2865
rect 4620 2895 4640 2915
rect 4620 2845 4640 2865
rect 4710 2895 4730 2915
rect 4710 2845 4730 2865
rect 4800 2895 4820 2915
rect 4800 2845 4820 2865
rect 4890 2895 4910 2915
rect 4890 2845 4910 2865
rect 4980 2895 5000 2915
rect 4980 2845 5000 2865
rect 2820 2665 2840 2685
rect 2820 2615 2840 2635
rect 2820 2565 2840 2585
rect 2820 2515 2840 2535
rect 2820 2465 2840 2485
rect 2820 2415 2840 2435
rect 2910 2665 2930 2685
rect 2910 2615 2930 2635
rect 2910 2565 2930 2585
rect 2910 2515 2930 2535
rect 2910 2465 2930 2485
rect 2910 2415 2930 2435
rect 3000 2665 3020 2685
rect 3000 2615 3020 2635
rect 3000 2565 3020 2585
rect 3000 2515 3020 2535
rect 3000 2465 3020 2485
rect 3000 2415 3020 2435
rect 3090 2665 3110 2685
rect 3090 2615 3110 2635
rect 3090 2565 3110 2585
rect 3090 2515 3110 2535
rect 3090 2465 3110 2485
rect 3090 2415 3110 2435
rect 3180 2665 3200 2685
rect 3180 2615 3200 2635
rect 3180 2565 3200 2585
rect 3180 2515 3200 2535
rect 3180 2465 3200 2485
rect 3180 2415 3200 2435
rect 3270 2665 3290 2685
rect 3270 2615 3290 2635
rect 3270 2565 3290 2585
rect 3270 2515 3290 2535
rect 3270 2465 3290 2485
rect 3270 2415 3290 2435
rect 3360 2665 3380 2685
rect 3360 2615 3380 2635
rect 3360 2565 3380 2585
rect 3360 2515 3380 2535
rect 3360 2465 3380 2485
rect 3360 2415 3380 2435
rect 3450 2665 3470 2685
rect 3450 2615 3470 2635
rect 3450 2565 3470 2585
rect 3450 2515 3470 2535
rect 3450 2465 3470 2485
rect 3450 2415 3470 2435
rect 3540 2665 3560 2685
rect 3540 2615 3560 2635
rect 3540 2565 3560 2585
rect 3540 2515 3560 2535
rect 3540 2465 3560 2485
rect 3540 2415 3560 2435
rect 3630 2665 3650 2685
rect 3630 2615 3650 2635
rect 3630 2565 3650 2585
rect 3630 2515 3650 2535
rect 3630 2465 3650 2485
rect 3630 2415 3650 2435
rect 3720 2665 3740 2685
rect 3720 2615 3740 2635
rect 3720 2565 3740 2585
rect 3720 2515 3740 2535
rect 3720 2465 3740 2485
rect 3720 2415 3740 2435
rect 3810 2665 3830 2685
rect 3810 2615 3830 2635
rect 3810 2565 3830 2585
rect 3810 2515 3830 2535
rect 3810 2465 3830 2485
rect 3810 2415 3830 2435
rect 3900 2665 3920 2685
rect 3900 2615 3920 2635
rect 3900 2565 3920 2585
rect 3900 2515 3920 2535
rect 3900 2465 3920 2485
rect 3900 2415 3920 2435
rect 3990 2665 4010 2685
rect 3990 2615 4010 2635
rect 3990 2565 4010 2585
rect 3990 2515 4010 2535
rect 3990 2465 4010 2485
rect 3990 2415 4010 2435
rect 4080 2665 4100 2685
rect 4080 2615 4100 2635
rect 4080 2565 4100 2585
rect 4080 2515 4100 2535
rect 4080 2465 4100 2485
rect 4080 2415 4100 2435
rect 4170 2665 4190 2685
rect 4170 2615 4190 2635
rect 4170 2565 4190 2585
rect 4170 2515 4190 2535
rect 4170 2465 4190 2485
rect 4170 2415 4190 2435
rect 4260 2665 4280 2685
rect 4260 2615 4280 2635
rect 4260 2565 4280 2585
rect 4260 2515 4280 2535
rect 4260 2465 4280 2485
rect 4260 2415 4280 2435
rect 4350 2665 4370 2685
rect 4350 2615 4370 2635
rect 4350 2565 4370 2585
rect 4350 2515 4370 2535
rect 4350 2465 4370 2485
rect 4350 2415 4370 2435
rect 4440 2665 4460 2685
rect 4440 2615 4460 2635
rect 4440 2565 4460 2585
rect 4440 2515 4460 2535
rect 4440 2465 4460 2485
rect 4440 2415 4460 2435
rect 4530 2665 4550 2685
rect 4530 2615 4550 2635
rect 4530 2565 4550 2585
rect 4530 2515 4550 2535
rect 4530 2465 4550 2485
rect 4530 2415 4550 2435
rect 4620 2665 4640 2685
rect 4620 2615 4640 2635
rect 4620 2565 4640 2585
rect 4620 2515 4640 2535
rect 4620 2465 4640 2485
rect 4620 2415 4640 2435
rect 4710 2665 4730 2685
rect 4710 2615 4730 2635
rect 4710 2565 4730 2585
rect 4710 2515 4730 2535
rect 4710 2465 4730 2485
rect 4710 2415 4730 2435
rect 4800 2665 4820 2685
rect 4800 2615 4820 2635
rect 4800 2565 4820 2585
rect 4800 2515 4820 2535
rect 4800 2465 4820 2485
rect 4800 2415 4820 2435
rect 4890 2665 4910 2685
rect 4890 2615 4910 2635
rect 4890 2565 4910 2585
rect 4890 2515 4910 2535
rect 4890 2465 4910 2485
rect 4890 2415 4910 2435
rect 4980 2665 5000 2685
rect 4980 2615 5000 2635
rect 4980 2565 5000 2585
rect 4980 2515 5000 2535
rect 4980 2465 5000 2485
rect 4980 2415 5000 2435
rect 5070 2665 5090 2685
rect 5070 2615 5090 2635
rect 5070 2565 5090 2585
rect 5070 2515 5090 2535
rect 5070 2465 5090 2485
rect 5070 2415 5090 2435
rect 5160 2665 5180 2685
rect 5160 2615 5180 2635
rect 5160 2565 5180 2585
rect 5160 2515 5180 2535
rect 5160 2465 5180 2485
rect 5160 2415 5180 2435
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 3955 1915 3975 1935
rect 4025 1965 4045 1985
rect 4025 1915 4045 1935
rect 4085 1965 4105 1985
rect 4085 1915 4105 1935
rect 4145 1965 4165 1985
rect 4145 1915 4165 1935
rect 4205 1965 4225 1985
rect 4205 1915 4225 1935
rect 4265 1965 4285 1985
rect 4265 1915 4285 1935
rect 4325 1965 4345 1985
rect 4325 1915 4345 1935
rect 4385 1965 4405 1985
rect 4385 1915 4405 1935
rect 4445 1965 4465 1985
rect 4445 1915 4465 1935
rect 4505 1965 4525 1985
rect 4505 1915 4525 1935
rect 4565 1965 4585 1985
rect 4565 1915 4585 1935
rect 4625 1965 4645 1985
rect 4625 1915 4645 1935
rect 4685 1965 4705 1985
rect 4685 1915 4705 1935
rect 4745 1965 4765 1985
rect 4745 1915 4765 1935
rect 4805 1965 4825 1985
rect 4805 1915 4825 1935
rect 4865 1965 4885 1985
rect 4865 1915 4885 1935
rect 4925 1965 4945 1985
rect 4925 1915 4945 1935
rect 4985 1965 5005 1985
rect 4985 1915 5005 1935
rect 5045 1965 5065 1985
rect 5045 1915 5065 1935
rect 5105 1965 5125 1985
rect 5105 1915 5125 1935
rect 5165 1965 5185 1985
rect 5165 1915 5185 1935
rect 5225 1965 5245 1985
rect 5225 1915 5245 1935
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4205 1630 4225 1650
rect 4265 1630 4285 1650
rect 4325 1630 4345 1650
rect 4385 1630 4405 1650
rect 4445 1630 4465 1650
rect 4505 1630 4525 1650
rect 4565 1630 4585 1650
rect 4625 1630 4645 1650
rect 4685 1630 4705 1650
rect 4745 1630 4765 1650
rect 4805 1630 4825 1650
rect 2845 1425 2865 1445
rect 2845 1375 2865 1395
rect 2845 1325 2865 1345
rect 2845 1275 2865 1295
rect 2845 1225 2865 1245
rect 3385 1425 3405 1445
rect 3385 1375 3405 1395
rect 3385 1325 3405 1345
rect 3385 1275 3405 1295
rect 3385 1225 3405 1245
rect 3925 1425 3945 1445
rect 3925 1375 3945 1395
rect 3925 1325 3945 1345
rect 3925 1275 3945 1295
rect 3925 1225 3945 1245
rect 4055 1425 4075 1445
rect 4055 1375 4075 1395
rect 4055 1325 4075 1345
rect 4055 1275 4075 1295
rect 4055 1225 4075 1245
rect 4595 1425 4615 1445
rect 4595 1375 4615 1395
rect 4595 1325 4615 1345
rect 4595 1275 4615 1295
rect 4595 1225 4615 1245
rect 5135 1425 5155 1445
rect 5135 1375 5155 1395
rect 5135 1325 5155 1345
rect 5135 1275 5155 1295
rect 5135 1225 5155 1245
rect 2950 1045 2970 1065
rect 2950 995 2970 1015
rect 3990 1045 4010 1065
rect 3990 995 4010 1015
rect 5030 1045 5050 1065
rect 5030 995 5050 1015
rect 3000 850 3020 870
rect 3000 800 3020 820
rect 3090 850 3110 870
rect 3090 800 3110 820
rect 3180 850 3200 870
rect 3180 800 3200 820
rect 3270 850 3290 870
rect 3270 800 3290 820
rect 3360 850 3380 870
rect 3360 800 3380 820
rect 3450 850 3470 870
rect 3450 800 3470 820
rect 3540 850 3560 870
rect 3540 800 3560 820
rect 3630 850 3650 870
rect 3630 800 3650 820
rect 3720 850 3740 870
rect 3720 800 3740 820
rect 3810 850 3830 870
rect 3810 800 3830 820
rect 3900 850 3920 870
rect 3900 800 3920 820
rect 3990 850 4010 870
rect 3990 800 4010 820
rect 4080 850 4100 870
rect 4080 800 4100 820
rect 4170 850 4190 870
rect 4170 800 4190 820
rect 4260 850 4280 870
rect 4260 800 4280 820
rect 4350 850 4370 870
rect 4350 800 4370 820
rect 4440 850 4460 870
rect 4440 800 4460 820
rect 4530 850 4550 870
rect 4530 800 4550 820
rect 4620 850 4640 870
rect 4620 800 4640 820
rect 4710 850 4730 870
rect 4710 800 4730 820
rect 4800 850 4820 870
rect 4800 800 4820 820
rect 4890 850 4910 870
rect 4890 800 4910 820
rect 4980 850 5000 870
rect 4980 800 5000 820
<< psubdiff >>
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
<< psubdiffcont >>
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
<< poly >>
rect 3135 2975 3170 2985
rect 3135 2955 3140 2975
rect 3160 2955 3170 2975
rect 3135 2945 3170 2955
rect 4830 2975 4865 2985
rect 4830 2955 4840 2975
rect 4860 2955 4865 2975
rect 4830 2945 4865 2955
rect 3030 2930 3080 2945
rect 3120 2930 3170 2945
rect 3210 2930 3260 2945
rect 3300 2930 3350 2945
rect 3390 2930 3440 2945
rect 3480 2930 3530 2945
rect 3570 2930 3620 2945
rect 3660 2930 3710 2945
rect 3750 2930 3800 2945
rect 3840 2930 3890 2945
rect 3930 2930 3980 2945
rect 4020 2930 4070 2945
rect 4110 2930 4160 2945
rect 4200 2930 4250 2945
rect 4290 2930 4340 2945
rect 4380 2930 4430 2945
rect 4470 2930 4520 2945
rect 4560 2930 4610 2945
rect 4650 2930 4700 2945
rect 4740 2930 4790 2945
rect 4830 2930 4880 2945
rect 4920 2930 4970 2945
rect 3030 2815 3080 2830
rect 2990 2805 3080 2815
rect 3120 2820 3170 2830
rect 3210 2820 3260 2830
rect 3300 2820 3350 2830
rect 3390 2820 3440 2830
rect 3480 2820 3530 2830
rect 3570 2820 3620 2830
rect 3660 2820 3710 2830
rect 3750 2820 3800 2830
rect 3840 2820 3890 2830
rect 3930 2820 3980 2830
rect 4020 2820 4070 2830
rect 4110 2820 4160 2830
rect 4200 2820 4250 2830
rect 4290 2820 4340 2830
rect 4380 2820 4430 2830
rect 4470 2820 4520 2830
rect 4560 2820 4610 2830
rect 4650 2820 4700 2830
rect 4740 2820 4790 2830
rect 4830 2820 4880 2830
rect 3120 2805 4880 2820
rect 4920 2815 4970 2830
rect 4920 2805 5010 2815
rect 2990 2785 3000 2805
rect 3020 2800 3080 2805
rect 4920 2800 4980 2805
rect 3020 2785 3030 2800
rect 2990 2775 3030 2785
rect 4970 2785 4980 2800
rect 5000 2785 5010 2805
rect 4970 2775 5010 2785
rect 2850 2700 2900 2715
rect 2940 2700 2990 2715
rect 3030 2700 3080 2715
rect 3120 2700 3170 2715
rect 3210 2700 3260 2715
rect 3300 2700 3350 2715
rect 3390 2700 3440 2715
rect 3480 2700 3530 2715
rect 3570 2700 3620 2715
rect 3660 2700 3710 2715
rect 3750 2700 3800 2715
rect 3840 2700 3890 2715
rect 3930 2700 3980 2715
rect 4020 2700 4070 2715
rect 4110 2700 4160 2715
rect 4200 2700 4250 2715
rect 4290 2700 4340 2715
rect 4380 2700 4430 2715
rect 4470 2700 4520 2715
rect 4560 2700 4610 2715
rect 4650 2700 4700 2715
rect 4740 2700 4790 2715
rect 4830 2700 4880 2715
rect 4920 2700 4970 2715
rect 5010 2700 5060 2715
rect 5100 2700 5150 2715
rect 2850 2390 2900 2400
rect 2810 2375 2900 2390
rect 2940 2390 2990 2400
rect 3030 2390 3080 2400
rect 3120 2390 3170 2400
rect 3210 2390 3260 2400
rect 3300 2390 3350 2400
rect 3390 2390 3440 2400
rect 3480 2390 3530 2400
rect 3570 2390 3620 2400
rect 3660 2390 3710 2400
rect 3750 2390 3800 2400
rect 3840 2390 3890 2400
rect 3930 2390 3980 2400
rect 4020 2390 4070 2400
rect 4110 2390 4160 2400
rect 4200 2390 4250 2400
rect 4290 2390 4340 2400
rect 4380 2390 4430 2400
rect 4470 2390 4520 2400
rect 4560 2390 4610 2400
rect 4650 2390 4700 2400
rect 4740 2390 4790 2400
rect 4830 2390 4880 2400
rect 4920 2390 4970 2400
rect 5010 2390 5060 2400
rect 2940 2375 5060 2390
rect 5100 2390 5150 2400
rect 5100 2375 5190 2390
rect 2810 2355 2820 2375
rect 2840 2355 2850 2375
rect 2810 2345 2850 2355
rect 2990 2370 3030 2375
rect 2990 2350 3000 2370
rect 3020 2350 3030 2370
rect 2990 2340 3030 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 5150 2355 5160 2375
rect 5180 2355 5190 2375
rect 5150 2345 5190 2355
rect 2745 2045 2785 2055
rect 2745 2025 2755 2045
rect 2775 2030 2785 2045
rect 3945 2045 3985 2055
rect 3945 2030 3955 2045
rect 2775 2025 2805 2030
rect 2745 2015 2805 2025
rect 3925 2025 3955 2030
rect 3975 2025 3985 2045
rect 3925 2015 3985 2025
rect 4015 2045 4055 2055
rect 4015 2025 4025 2045
rect 4045 2030 4055 2045
rect 5215 2045 5255 2055
rect 5215 2030 5225 2045
rect 4045 2025 4075 2030
rect 4015 2015 4075 2025
rect 5195 2025 5225 2030
rect 5245 2025 5255 2045
rect 5195 2015 5255 2025
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4055 2000 4075 2015
rect 4115 2000 4135 2015
rect 4175 2000 4195 2015
rect 4235 2000 4255 2015
rect 4295 2000 4315 2015
rect 4355 2000 4375 2015
rect 4415 2000 4435 2015
rect 4475 2000 4495 2015
rect 4535 2000 4555 2015
rect 4595 2000 4615 2015
rect 4655 2000 4675 2015
rect 4715 2000 4735 2015
rect 4775 2000 4795 2015
rect 4835 2000 4855 2015
rect 4895 2000 4915 2015
rect 4955 2000 4975 2015
rect 5015 2000 5035 2015
rect 5075 2000 5095 2015
rect 5135 2000 5155 2015
rect 5195 2000 5215 2015
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1885 3945 1900
rect 4055 1885 4075 1900
rect 4115 1885 4135 1900
rect 4175 1890 4195 1900
rect 4235 1890 4255 1900
rect 4295 1890 4315 1900
rect 4355 1890 4375 1900
rect 3855 1875 3895 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 4105 1875 4145 1885
rect 4175 1875 4375 1890
rect 4415 1890 4435 1900
rect 4475 1890 4495 1900
rect 4415 1875 4495 1890
rect 4535 1890 4555 1900
rect 4595 1890 4615 1900
rect 4655 1890 4675 1900
rect 4715 1890 4735 1900
rect 4535 1875 4735 1890
rect 4775 1890 4795 1900
rect 4835 1890 4855 1900
rect 4775 1875 4855 1890
rect 4895 1890 4915 1900
rect 4955 1890 4975 1900
rect 5015 1890 5035 1900
rect 5075 1890 5095 1900
rect 4895 1875 5095 1890
rect 5135 1885 5155 1900
rect 5195 1885 5215 1900
rect 5125 1875 5165 1885
rect 4105 1855 4115 1875
rect 4135 1855 4145 1875
rect 4105 1845 4145 1855
rect 4315 1855 4325 1875
rect 4345 1855 4355 1875
rect 4315 1845 4355 1855
rect 4435 1855 4445 1875
rect 4465 1855 4475 1875
rect 4435 1845 4475 1855
rect 4675 1855 4685 1875
rect 4705 1855 4715 1875
rect 4675 1845 4715 1855
rect 4795 1855 4805 1875
rect 4825 1855 4835 1875
rect 4795 1845 4835 1855
rect 5035 1855 5045 1875
rect 5065 1855 5075 1875
rect 5035 1845 5075 1855
rect 5125 1855 5135 1875
rect 5155 1855 5165 1875
rect 5125 1845 5165 1855
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4735 1755 4775 1765
rect 4735 1735 4745 1755
rect 4765 1735 4775 1755
rect 4735 1720 4775 1735
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4235 1705 4775 1720
rect 4235 1665 4255 1705
rect 4295 1665 4315 1680
rect 4355 1665 4375 1680
rect 4415 1665 4435 1705
rect 4475 1665 4495 1705
rect 4535 1665 4555 1680
rect 4595 1665 4615 1680
rect 4655 1665 4675 1705
rect 4715 1665 4735 1705
rect 4775 1665 4795 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4235 1600 4255 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4295 1575 4315 1615
rect 4355 1575 4375 1615
rect 4415 1600 4435 1615
rect 4475 1600 4495 1615
rect 4535 1575 4555 1615
rect 4595 1575 4615 1615
rect 4655 1600 4675 1615
rect 4715 1600 4735 1615
rect 4775 1600 4795 1615
rect 4775 1590 4835 1600
rect 4775 1575 4805 1590
rect 4295 1570 4805 1575
rect 4825 1570 4835 1590
rect 4295 1560 4835 1570
rect 2875 1460 3375 1475
rect 3415 1460 3915 1475
rect 4085 1460 4585 1475
rect 4625 1460 5125 1475
rect 2875 1195 3375 1210
rect 3415 1195 3915 1210
rect 4085 1195 4585 1210
rect 4625 1195 5125 1210
rect 3020 1125 3060 1135
rect 3020 1105 3030 1125
rect 3050 1105 3060 1125
rect 3020 1095 3060 1105
rect 3100 1125 3140 1135
rect 3100 1105 3110 1125
rect 3130 1105 3140 1125
rect 3100 1095 3140 1105
rect 3180 1125 3220 1135
rect 3180 1105 3190 1125
rect 3210 1105 3220 1125
rect 3180 1095 3220 1105
rect 3260 1125 3300 1135
rect 3260 1105 3270 1125
rect 3290 1105 3300 1125
rect 3260 1095 3300 1105
rect 3340 1125 3380 1135
rect 3340 1105 3350 1125
rect 3370 1105 3380 1125
rect 3340 1095 3380 1105
rect 3420 1125 3460 1135
rect 3420 1105 3430 1125
rect 3450 1105 3460 1125
rect 3420 1095 3460 1105
rect 3500 1125 3540 1135
rect 3500 1105 3510 1125
rect 3530 1105 3540 1125
rect 3500 1095 3540 1105
rect 3580 1125 3620 1135
rect 3580 1105 3590 1125
rect 3610 1105 3620 1125
rect 3580 1095 3620 1105
rect 3660 1125 3700 1135
rect 3660 1105 3670 1125
rect 3690 1105 3700 1125
rect 3660 1095 3700 1105
rect 3740 1125 3780 1135
rect 3740 1105 3750 1125
rect 3770 1105 3780 1125
rect 3740 1095 3780 1105
rect 3820 1125 3860 1135
rect 3820 1105 3830 1125
rect 3850 1105 3860 1125
rect 3820 1095 3860 1105
rect 3900 1125 3940 1135
rect 3900 1105 3910 1125
rect 3930 1105 3940 1125
rect 3900 1095 3940 1105
rect 4060 1125 4100 1135
rect 4060 1105 4070 1125
rect 4090 1105 4100 1125
rect 4060 1095 4100 1105
rect 4140 1125 4180 1135
rect 4140 1105 4150 1125
rect 4170 1105 4180 1125
rect 4140 1095 4180 1105
rect 4220 1125 4260 1135
rect 4220 1105 4230 1125
rect 4250 1105 4260 1125
rect 4220 1095 4260 1105
rect 4300 1125 4340 1135
rect 4300 1105 4310 1125
rect 4330 1105 4340 1125
rect 4300 1095 4340 1105
rect 4380 1125 4420 1135
rect 4380 1105 4390 1125
rect 4410 1105 4420 1125
rect 4380 1095 4420 1105
rect 4460 1125 4500 1135
rect 4460 1105 4470 1125
rect 4490 1105 4500 1125
rect 4460 1095 4500 1105
rect 4540 1125 4580 1135
rect 4540 1105 4550 1125
rect 4570 1105 4580 1125
rect 4540 1095 4580 1105
rect 4620 1125 4660 1135
rect 4620 1105 4630 1125
rect 4650 1105 4660 1125
rect 4620 1095 4660 1105
rect 4700 1125 4740 1135
rect 4700 1105 4710 1125
rect 4730 1105 4740 1125
rect 4700 1095 4740 1105
rect 4780 1125 4820 1135
rect 4780 1105 4790 1125
rect 4810 1105 4820 1125
rect 4780 1095 4820 1105
rect 4860 1125 4900 1135
rect 4860 1105 4870 1125
rect 4890 1105 4900 1125
rect 4860 1095 4900 1105
rect 4940 1125 4980 1135
rect 4940 1105 4950 1125
rect 4970 1105 4980 1125
rect 4940 1095 4980 1105
rect 2980 1080 3980 1095
rect 4020 1080 5020 1095
rect 2980 965 3980 980
rect 4020 965 5020 980
rect 2990 930 3030 940
rect 2990 910 3000 930
rect 3020 910 3030 930
rect 4970 930 5010 940
rect 4970 910 4980 930
rect 5000 910 5010 930
rect 2990 895 3080 910
rect 3030 885 3080 895
rect 3120 895 4880 910
rect 3120 885 3170 895
rect 3210 885 3260 895
rect 3300 885 3350 895
rect 3390 885 3440 895
rect 3480 885 3530 895
rect 3570 885 3620 895
rect 3660 885 3710 895
rect 3750 885 3800 895
rect 3840 885 3890 895
rect 3930 885 3980 895
rect 4020 885 4070 895
rect 4110 885 4160 895
rect 4200 885 4250 895
rect 4290 885 4340 895
rect 4380 885 4430 895
rect 4470 885 4520 895
rect 4560 885 4610 895
rect 4650 885 4700 895
rect 4740 885 4790 895
rect 4830 885 4880 895
rect 4920 895 5010 910
rect 4920 885 4970 895
rect 3030 770 3080 785
rect 3120 770 3170 785
rect 3210 770 3260 785
rect 3300 770 3350 785
rect 3390 770 3440 785
rect 3480 770 3530 785
rect 3570 770 3620 785
rect 3660 770 3710 785
rect 3750 770 3800 785
rect 3840 770 3890 785
rect 3930 770 3980 785
rect 4020 770 4070 785
rect 4110 770 4160 785
rect 4200 770 4250 785
rect 4290 770 4340 785
rect 4380 770 4430 785
rect 4470 770 4520 785
rect 4560 770 4610 785
rect 4650 770 4700 785
rect 4740 770 4790 785
rect 4830 770 4880 785
rect 4920 770 4970 785
<< polycont >>
rect 3140 2955 3160 2975
rect 4840 2955 4860 2975
rect 3000 2785 3020 2805
rect 4980 2785 5000 2805
rect 2820 2355 2840 2375
rect 3000 2350 3020 2370
rect 3895 2355 3915 2375
rect 5160 2355 5180 2375
rect 2755 2025 2775 2045
rect 3955 2025 3975 2045
rect 4025 2025 4045 2045
rect 5225 2025 5245 2045
rect 2630 1855 2650 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 4115 1855 4135 1875
rect 4325 1855 4345 1875
rect 4445 1855 4465 1875
rect 4685 1855 4705 1875
rect 4805 1855 4825 1875
rect 5045 1855 5065 1875
rect 5135 1855 5155 1875
rect 3235 1735 3255 1755
rect 4745 1735 4765 1755
rect 3175 1570 3195 1590
rect 4805 1570 4825 1590
rect 3030 1105 3050 1125
rect 3110 1105 3130 1125
rect 3190 1105 3210 1125
rect 3270 1105 3290 1125
rect 3350 1105 3370 1125
rect 3430 1105 3450 1125
rect 3510 1105 3530 1125
rect 3590 1105 3610 1125
rect 3670 1105 3690 1125
rect 3750 1105 3770 1125
rect 3830 1105 3850 1125
rect 3910 1105 3930 1125
rect 4070 1105 4090 1125
rect 4150 1105 4170 1125
rect 4230 1105 4250 1125
rect 4310 1105 4330 1125
rect 4390 1105 4410 1125
rect 4470 1105 4490 1125
rect 4550 1105 4570 1125
rect 4630 1105 4650 1125
rect 4710 1105 4730 1125
rect 4790 1105 4810 1125
rect 4870 1105 4890 1125
rect 4950 1105 4970 1125
rect 3000 910 3020 930
rect 4980 910 5000 930
<< xpolycontact >>
rect 85 3170 305 3205
rect 910 3170 1130 3205
rect 1290 3165 1510 3200
rect 2110 3165 2330 3200
rect 85 3110 305 3145
rect 910 3110 1130 3145
rect 1290 3105 1510 3140
rect 2110 3105 2330 3140
rect 85 3030 305 3065
rect 905 3030 1125 3065
rect 1290 3045 1510 3080
rect 2110 3045 2330 3080
rect 85 2970 305 3005
rect 905 2970 1125 3005
rect 1290 2985 1510 3020
rect 2110 2985 2330 3020
rect 1290 2925 1510 2960
rect 2110 2925 2330 2960
rect 1290 2865 1510 2900
rect 2110 2865 2330 2900
rect 85 2820 305 2855
rect 355 2820 575 2855
rect 1290 2805 1510 2840
rect 1740 2805 1960 2840
rect 85 2760 305 2795
rect 355 2760 575 2795
<< xpolyres >>
rect 305 3170 910 3205
rect 1510 3165 2110 3200
rect 305 3110 910 3145
rect 1510 3105 2110 3140
rect 305 3030 905 3065
rect 1510 3045 2110 3080
rect 305 2970 905 3005
rect 1510 2985 2110 3020
rect 1510 2925 2110 2960
rect 1510 2865 2110 2900
rect 305 2820 355 2855
rect 1510 2805 1740 2840
rect 305 2760 355 2795
<< locali >>
rect 1250 3495 1280 3525
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1195 3310 1225 3340
rect 3135 3310 3165 3340
rect 3395 3305 3425 3335
rect 5345 3305 5375 3335
rect 1150 3255 1180 3285
rect 4885 3255 4915 3285
rect 5395 3255 5425 3285
rect 2740 3210 2770 3240
rect 40 3200 85 3205
rect 40 3175 50 3200
rect 75 3175 85 3200
rect 40 3170 85 3175
rect 1110 3145 1130 3170
rect 1245 3195 1290 3200
rect 1245 3170 1255 3195
rect 1280 3170 1290 3195
rect 1245 3165 1290 3170
rect 2330 3165 2370 3200
rect 40 3140 85 3145
rect 40 3115 50 3140
rect 75 3115 85 3140
rect 40 3110 85 3115
rect 1245 3135 1290 3140
rect 1245 3110 1255 3135
rect 1280 3110 1290 3135
rect 1245 3105 1290 3110
rect 1150 3070 1180 3100
rect 2295 3080 2330 3105
rect 40 3060 85 3065
rect 40 3035 50 3060
rect 75 3035 85 3060
rect 40 3030 85 3035
rect 1105 3005 1125 3030
rect 40 3000 85 3005
rect 40 2975 50 3000
rect 75 2975 85 3000
rect 40 2970 85 2975
rect 1250 3045 1290 3080
rect 1250 2900 1270 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 3135 3110 3165 3140
rect 4835 3110 4865 3140
rect 5300 3110 5330 3140
rect 3985 3050 4015 3080
rect 2330 2985 2370 3020
rect 3445 3005 3475 3035
rect 3805 3005 3835 3035
rect 4345 3005 4375 3035
rect 4705 3005 4735 3035
rect 1290 2960 1325 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3075 2975 3115 2985
rect 3075 2955 3085 2975
rect 3105 2955 3115 2975
rect 3075 2945 3115 2955
rect 3135 2975 3170 2985
rect 3135 2955 3140 2975
rect 3160 2955 3170 2975
rect 3135 2945 3170 2955
rect 3260 2975 3300 2985
rect 3260 2955 3270 2975
rect 3290 2955 3300 2975
rect 3260 2945 3300 2955
rect 3440 2975 3480 2985
rect 3440 2955 3450 2975
rect 3470 2955 3480 2975
rect 3440 2945 3480 2955
rect 3620 2975 3660 2985
rect 3620 2955 3630 2975
rect 3650 2955 3660 2975
rect 3620 2945 3660 2955
rect 3800 2975 3840 2985
rect 3800 2955 3810 2975
rect 3830 2955 3840 2975
rect 3800 2945 3840 2955
rect 3980 2975 4020 2985
rect 3980 2955 3990 2975
rect 4010 2955 4020 2975
rect 3980 2945 4020 2955
rect 4160 2975 4200 2985
rect 4160 2955 4170 2975
rect 4190 2955 4200 2975
rect 4160 2945 4200 2955
rect 4340 2975 4380 2985
rect 4340 2955 4350 2975
rect 4370 2955 4380 2975
rect 4340 2945 4380 2955
rect 4520 2975 4560 2985
rect 4520 2955 4530 2975
rect 4550 2955 4560 2975
rect 4520 2945 4560 2955
rect 4700 2975 4740 2985
rect 4700 2955 4710 2975
rect 4730 2955 4740 2975
rect 4700 2945 4740 2955
rect 4830 2975 4865 2985
rect 4830 2955 4840 2975
rect 4860 2955 4865 2975
rect 4830 2945 4865 2955
rect 4885 2975 4920 2985
rect 4885 2955 4890 2975
rect 4910 2955 4920 2975
rect 4885 2945 4920 2955
rect 3090 2925 3110 2945
rect 3270 2925 3290 2945
rect 3450 2925 3470 2945
rect 3630 2925 3650 2945
rect 3810 2925 3830 2945
rect 3990 2925 4010 2945
rect 4170 2925 4190 2945
rect 4350 2925 4370 2945
rect 4530 2925 4550 2945
rect 4710 2925 4730 2945
rect 4890 2925 4910 2945
rect 2995 2915 3025 2925
rect 1250 2865 1290 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2995 2895 3000 2915
rect 3020 2895 3025 2915
rect 2995 2865 3025 2895
rect -55 2825 -25 2855
rect 40 2850 85 2855
rect 40 2825 50 2850
rect 75 2825 85 2850
rect 40 2820 85 2825
rect 575 2850 620 2855
rect 575 2825 585 2850
rect 610 2825 620 2850
rect 575 2820 620 2825
rect 1195 2820 1225 2850
rect 2995 2845 3000 2865
rect 3020 2845 3025 2865
rect 1245 2835 1290 2840
rect 1245 2810 1255 2835
rect 1280 2810 1290 2835
rect 1245 2805 1290 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2995 2835 3025 2845
rect 3085 2915 3115 2925
rect 3085 2895 3090 2915
rect 3110 2895 3115 2915
rect 3085 2865 3115 2895
rect 3085 2845 3090 2865
rect 3110 2845 3115 2865
rect 3085 2835 3115 2845
rect 3175 2915 3205 2925
rect 3175 2895 3180 2915
rect 3200 2895 3205 2915
rect 3175 2865 3205 2895
rect 3175 2845 3180 2865
rect 3200 2845 3205 2865
rect 3175 2835 3205 2845
rect 3265 2915 3295 2925
rect 3265 2895 3270 2915
rect 3290 2895 3295 2915
rect 3265 2865 3295 2895
rect 3265 2845 3270 2865
rect 3290 2845 3295 2865
rect 3265 2835 3295 2845
rect 3355 2915 3385 2925
rect 3355 2895 3360 2915
rect 3380 2895 3385 2915
rect 3355 2865 3385 2895
rect 3355 2845 3360 2865
rect 3380 2845 3385 2865
rect 3355 2835 3385 2845
rect 3445 2915 3475 2925
rect 3445 2895 3450 2915
rect 3470 2895 3475 2915
rect 3445 2865 3475 2895
rect 3445 2845 3450 2865
rect 3470 2845 3475 2865
rect 3445 2835 3475 2845
rect 3535 2915 3565 2925
rect 3535 2895 3540 2915
rect 3560 2895 3565 2915
rect 3535 2865 3565 2895
rect 3535 2845 3540 2865
rect 3560 2845 3565 2865
rect 3535 2835 3565 2845
rect 3625 2915 3655 2925
rect 3625 2895 3630 2915
rect 3650 2895 3655 2915
rect 3625 2865 3655 2895
rect 3625 2845 3630 2865
rect 3650 2845 3655 2865
rect 3625 2835 3655 2845
rect 3715 2915 3745 2925
rect 3715 2895 3720 2915
rect 3740 2895 3745 2915
rect 3715 2865 3745 2895
rect 3715 2845 3720 2865
rect 3740 2845 3745 2865
rect 3715 2835 3745 2845
rect 3805 2915 3835 2925
rect 3805 2895 3810 2915
rect 3830 2895 3835 2915
rect 3805 2865 3835 2895
rect 3805 2845 3810 2865
rect 3830 2845 3835 2865
rect 3805 2835 3835 2845
rect 3895 2915 3925 2925
rect 3895 2895 3900 2915
rect 3920 2895 3925 2915
rect 3895 2865 3925 2895
rect 3895 2845 3900 2865
rect 3920 2845 3925 2865
rect 3895 2835 3925 2845
rect 3985 2915 4015 2925
rect 3985 2895 3990 2915
rect 4010 2895 4015 2915
rect 3985 2865 4015 2895
rect 3985 2845 3990 2865
rect 4010 2845 4015 2865
rect 3985 2835 4015 2845
rect 4075 2915 4105 2925
rect 4075 2895 4080 2915
rect 4100 2895 4105 2915
rect 4075 2865 4105 2895
rect 4075 2845 4080 2865
rect 4100 2845 4105 2865
rect 4075 2835 4105 2845
rect 4165 2915 4195 2925
rect 4165 2895 4170 2915
rect 4190 2895 4195 2915
rect 4165 2865 4195 2895
rect 4165 2845 4170 2865
rect 4190 2845 4195 2865
rect 4165 2835 4195 2845
rect 4255 2915 4285 2925
rect 4255 2895 4260 2915
rect 4280 2895 4285 2915
rect 4255 2865 4285 2895
rect 4255 2845 4260 2865
rect 4280 2845 4285 2865
rect 4255 2835 4285 2845
rect 4345 2915 4375 2925
rect 4345 2895 4350 2915
rect 4370 2895 4375 2915
rect 4345 2865 4375 2895
rect 4345 2845 4350 2865
rect 4370 2845 4375 2865
rect 4345 2835 4375 2845
rect 4435 2915 4465 2925
rect 4435 2895 4440 2915
rect 4460 2895 4465 2915
rect 4435 2865 4465 2895
rect 4435 2845 4440 2865
rect 4460 2845 4465 2865
rect 4435 2835 4465 2845
rect 4525 2915 4555 2925
rect 4525 2895 4530 2915
rect 4550 2895 4555 2915
rect 4525 2865 4555 2895
rect 4525 2845 4530 2865
rect 4550 2845 4555 2865
rect 4525 2835 4555 2845
rect 4615 2915 4645 2925
rect 4615 2895 4620 2915
rect 4640 2895 4645 2915
rect 4615 2865 4645 2895
rect 4615 2845 4620 2865
rect 4640 2845 4645 2865
rect 4615 2835 4645 2845
rect 4705 2915 4735 2925
rect 4705 2895 4710 2915
rect 4730 2895 4735 2915
rect 4705 2865 4735 2895
rect 4705 2845 4710 2865
rect 4730 2845 4735 2865
rect 4705 2835 4735 2845
rect 4795 2915 4825 2925
rect 4795 2895 4800 2915
rect 4820 2895 4825 2915
rect 4795 2865 4825 2895
rect 4795 2845 4800 2865
rect 4820 2845 4825 2865
rect 4795 2835 4825 2845
rect 4885 2915 4915 2925
rect 4885 2895 4890 2915
rect 4910 2895 4915 2915
rect 4885 2865 4915 2895
rect 4885 2845 4890 2865
rect 4910 2845 4915 2865
rect 4885 2835 4915 2845
rect 4975 2915 5005 2925
rect 4975 2895 4980 2915
rect 5000 2895 5005 2915
rect 4975 2865 5005 2895
rect 4975 2845 4980 2865
rect 5000 2845 5005 2865
rect 4975 2835 5005 2845
rect 3000 2815 3020 2835
rect 3180 2815 3200 2835
rect 3360 2815 3380 2835
rect 3540 2815 3560 2835
rect 3720 2815 3740 2835
rect 3900 2815 3920 2835
rect 4080 2815 4100 2835
rect 4260 2815 4280 2835
rect 4440 2815 4460 2835
rect 4620 2815 4640 2835
rect 4800 2815 4820 2835
rect 4980 2815 5000 2835
rect 2990 2805 3030 2815
rect -10 2765 20 2795
rect 40 2790 85 2795
rect 40 2765 50 2790
rect 75 2765 85 2790
rect 40 2760 85 2765
rect 575 2790 620 2795
rect 575 2765 585 2790
rect 610 2765 620 2790
rect 575 2760 620 2765
rect 2620 2755 2660 2795
rect 2990 2785 3000 2805
rect 3020 2785 3030 2805
rect 2990 2775 3030 2785
rect 3170 2805 3210 2815
rect 3170 2785 3180 2805
rect 3200 2785 3210 2805
rect 3170 2775 3210 2785
rect 3350 2805 3390 2815
rect 3350 2785 3360 2805
rect 3380 2785 3390 2805
rect 3350 2775 3390 2785
rect 3530 2805 3570 2815
rect 3530 2785 3540 2805
rect 3560 2785 3570 2805
rect 3530 2775 3570 2785
rect 3710 2805 3750 2815
rect 3710 2785 3720 2805
rect 3740 2785 3750 2805
rect 3710 2775 3750 2785
rect 3890 2805 3930 2815
rect 3890 2785 3900 2805
rect 3920 2785 3930 2805
rect 3890 2775 3930 2785
rect 4070 2805 4110 2815
rect 4070 2785 4080 2805
rect 4100 2785 4110 2805
rect 4070 2775 4110 2785
rect 4250 2805 4290 2815
rect 4250 2785 4260 2805
rect 4280 2785 4290 2805
rect 4250 2775 4290 2785
rect 4430 2805 4470 2815
rect 4430 2785 4440 2805
rect 4460 2785 4470 2805
rect 4430 2775 4470 2785
rect 4610 2805 4650 2815
rect 4610 2785 4620 2805
rect 4640 2785 4650 2805
rect 4610 2775 4650 2785
rect 4790 2805 4830 2815
rect 4790 2785 4800 2805
rect 4820 2785 4830 2805
rect 4790 2775 4830 2785
rect 4970 2805 5010 2815
rect 4970 2785 4980 2805
rect 5000 2785 5010 2805
rect 4970 2775 5010 2785
rect 1250 2715 1280 2745
rect 2150 2710 2190 2750
rect 2990 2745 3030 2755
rect 2990 2725 3000 2745
rect 3020 2725 3030 2745
rect 2990 2715 3030 2725
rect 3170 2745 3210 2755
rect 3170 2725 3180 2745
rect 3200 2725 3210 2745
rect 3170 2715 3210 2725
rect 3350 2745 3390 2755
rect 3350 2725 3360 2745
rect 3380 2725 3390 2745
rect 3350 2715 3390 2725
rect 3530 2745 3570 2755
rect 3530 2725 3540 2745
rect 3560 2725 3570 2745
rect 3530 2715 3570 2725
rect 3710 2745 3750 2755
rect 3710 2725 3720 2745
rect 3740 2725 3750 2745
rect 3710 2715 3750 2725
rect 3890 2745 3930 2755
rect 3890 2725 3900 2745
rect 3920 2725 3930 2745
rect 3890 2715 3930 2725
rect 4070 2745 4110 2755
rect 4070 2725 4080 2745
rect 4100 2725 4110 2745
rect 4070 2715 4110 2725
rect 4250 2745 4290 2755
rect 4250 2725 4260 2745
rect 4280 2725 4290 2745
rect 4250 2715 4290 2725
rect 4430 2745 4470 2755
rect 4430 2725 4440 2745
rect 4460 2725 4470 2745
rect 4430 2715 4470 2725
rect 4610 2745 4650 2755
rect 4610 2725 4620 2745
rect 4640 2725 4650 2745
rect 4610 2715 4650 2725
rect 4790 2745 4830 2755
rect 4790 2725 4800 2745
rect 4820 2725 4830 2745
rect 4790 2715 4830 2725
rect 4970 2745 5010 2755
rect 4970 2725 4980 2745
rect 5000 2725 5010 2745
rect 4970 2715 5010 2725
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3000 2695 3020 2715
rect 3180 2695 3200 2715
rect 3360 2695 3380 2715
rect 3540 2695 3560 2715
rect 3720 2695 3740 2715
rect 3900 2695 3920 2715
rect 4080 2695 4100 2715
rect 4260 2695 4280 2715
rect 4440 2695 4460 2715
rect 4620 2695 4640 2715
rect 4800 2695 4820 2715
rect 4980 2695 5000 2715
rect 2815 2685 2845 2695
rect 2815 2665 2820 2685
rect 2840 2665 2845 2685
rect 2815 2635 2845 2665
rect 2815 2615 2820 2635
rect 2840 2615 2845 2635
rect 2815 2585 2845 2615
rect 2815 2565 2820 2585
rect 2840 2565 2845 2585
rect 2815 2535 2845 2565
rect 2815 2515 2820 2535
rect 2840 2515 2845 2535
rect 2815 2485 2845 2515
rect 2815 2465 2820 2485
rect 2840 2465 2845 2485
rect 2815 2435 2845 2465
rect 2815 2415 2820 2435
rect 2840 2415 2845 2435
rect 2815 2405 2845 2415
rect 2905 2685 2935 2695
rect 2905 2665 2910 2685
rect 2930 2665 2935 2685
rect 2905 2635 2935 2665
rect 2905 2615 2910 2635
rect 2930 2615 2935 2635
rect 2905 2585 2935 2615
rect 2905 2565 2910 2585
rect 2930 2565 2935 2585
rect 2905 2535 2935 2565
rect 2905 2515 2910 2535
rect 2930 2515 2935 2535
rect 2905 2485 2935 2515
rect 2905 2465 2910 2485
rect 2930 2465 2935 2485
rect 2905 2435 2935 2465
rect 2905 2415 2910 2435
rect 2930 2415 2935 2435
rect 2905 2405 2935 2415
rect 2995 2685 3025 2695
rect 2995 2665 3000 2685
rect 3020 2665 3025 2685
rect 2995 2635 3025 2665
rect 2995 2615 3000 2635
rect 3020 2615 3025 2635
rect 2995 2585 3025 2615
rect 2995 2565 3000 2585
rect 3020 2565 3025 2585
rect 2995 2535 3025 2565
rect 2995 2515 3000 2535
rect 3020 2515 3025 2535
rect 2995 2485 3025 2515
rect 2995 2465 3000 2485
rect 3020 2465 3025 2485
rect 2995 2435 3025 2465
rect 2995 2415 3000 2435
rect 3020 2415 3025 2435
rect 2995 2405 3025 2415
rect 3085 2685 3115 2695
rect 3085 2665 3090 2685
rect 3110 2665 3115 2685
rect 3085 2635 3115 2665
rect 3085 2615 3090 2635
rect 3110 2615 3115 2635
rect 3085 2585 3115 2615
rect 3085 2565 3090 2585
rect 3110 2565 3115 2585
rect 3085 2535 3115 2565
rect 3085 2515 3090 2535
rect 3110 2515 3115 2535
rect 3085 2485 3115 2515
rect 3085 2465 3090 2485
rect 3110 2465 3115 2485
rect 3085 2435 3115 2465
rect 3085 2415 3090 2435
rect 3110 2415 3115 2435
rect 3085 2405 3115 2415
rect 3175 2685 3205 2695
rect 3175 2665 3180 2685
rect 3200 2665 3205 2685
rect 3175 2635 3205 2665
rect 3175 2615 3180 2635
rect 3200 2615 3205 2635
rect 3175 2585 3205 2615
rect 3175 2565 3180 2585
rect 3200 2565 3205 2585
rect 3175 2535 3205 2565
rect 3175 2515 3180 2535
rect 3200 2515 3205 2535
rect 3175 2485 3205 2515
rect 3175 2465 3180 2485
rect 3200 2465 3205 2485
rect 3175 2435 3205 2465
rect 3175 2415 3180 2435
rect 3200 2415 3205 2435
rect 3175 2405 3205 2415
rect 3265 2685 3295 2695
rect 3265 2665 3270 2685
rect 3290 2665 3295 2685
rect 3265 2635 3295 2665
rect 3265 2615 3270 2635
rect 3290 2615 3295 2635
rect 3265 2585 3295 2615
rect 3265 2565 3270 2585
rect 3290 2565 3295 2585
rect 3265 2535 3295 2565
rect 3265 2515 3270 2535
rect 3290 2515 3295 2535
rect 3265 2485 3295 2515
rect 3265 2465 3270 2485
rect 3290 2465 3295 2485
rect 3265 2435 3295 2465
rect 3265 2415 3270 2435
rect 3290 2415 3295 2435
rect 3265 2405 3295 2415
rect 3355 2685 3385 2695
rect 3355 2665 3360 2685
rect 3380 2665 3385 2685
rect 3355 2635 3385 2665
rect 3355 2615 3360 2635
rect 3380 2615 3385 2635
rect 3355 2585 3385 2615
rect 3355 2565 3360 2585
rect 3380 2565 3385 2585
rect 3355 2535 3385 2565
rect 3355 2515 3360 2535
rect 3380 2515 3385 2535
rect 3355 2485 3385 2515
rect 3355 2465 3360 2485
rect 3380 2465 3385 2485
rect 3355 2435 3385 2465
rect 3355 2415 3360 2435
rect 3380 2415 3385 2435
rect 3355 2405 3385 2415
rect 3445 2685 3475 2695
rect 3445 2665 3450 2685
rect 3470 2665 3475 2685
rect 3445 2635 3475 2665
rect 3445 2615 3450 2635
rect 3470 2615 3475 2635
rect 3445 2585 3475 2615
rect 3445 2565 3450 2585
rect 3470 2565 3475 2585
rect 3445 2535 3475 2565
rect 3445 2515 3450 2535
rect 3470 2515 3475 2535
rect 3445 2485 3475 2515
rect 3445 2465 3450 2485
rect 3470 2465 3475 2485
rect 3445 2435 3475 2465
rect 3445 2415 3450 2435
rect 3470 2415 3475 2435
rect 3445 2405 3475 2415
rect 3535 2685 3565 2695
rect 3535 2665 3540 2685
rect 3560 2665 3565 2685
rect 3535 2635 3565 2665
rect 3535 2615 3540 2635
rect 3560 2615 3565 2635
rect 3535 2585 3565 2615
rect 3535 2565 3540 2585
rect 3560 2565 3565 2585
rect 3535 2535 3565 2565
rect 3535 2515 3540 2535
rect 3560 2515 3565 2535
rect 3535 2485 3565 2515
rect 3535 2465 3540 2485
rect 3560 2465 3565 2485
rect 3535 2435 3565 2465
rect 3535 2415 3540 2435
rect 3560 2415 3565 2435
rect 3535 2405 3565 2415
rect 3625 2685 3655 2695
rect 3625 2665 3630 2685
rect 3650 2665 3655 2685
rect 3625 2635 3655 2665
rect 3625 2615 3630 2635
rect 3650 2615 3655 2635
rect 3625 2585 3655 2615
rect 3625 2565 3630 2585
rect 3650 2565 3655 2585
rect 3625 2535 3655 2565
rect 3625 2515 3630 2535
rect 3650 2515 3655 2535
rect 3625 2485 3655 2515
rect 3625 2465 3630 2485
rect 3650 2465 3655 2485
rect 3625 2435 3655 2465
rect 3625 2415 3630 2435
rect 3650 2415 3655 2435
rect 3625 2405 3655 2415
rect 3715 2685 3745 2695
rect 3715 2665 3720 2685
rect 3740 2665 3745 2685
rect 3715 2635 3745 2665
rect 3715 2615 3720 2635
rect 3740 2615 3745 2635
rect 3715 2585 3745 2615
rect 3715 2565 3720 2585
rect 3740 2565 3745 2585
rect 3715 2535 3745 2565
rect 3715 2515 3720 2535
rect 3740 2515 3745 2535
rect 3715 2485 3745 2515
rect 3715 2465 3720 2485
rect 3740 2465 3745 2485
rect 3715 2435 3745 2465
rect 3715 2415 3720 2435
rect 3740 2415 3745 2435
rect 3715 2405 3745 2415
rect 3805 2685 3835 2695
rect 3805 2665 3810 2685
rect 3830 2665 3835 2685
rect 3805 2635 3835 2665
rect 3805 2615 3810 2635
rect 3830 2615 3835 2635
rect 3805 2585 3835 2615
rect 3805 2565 3810 2585
rect 3830 2565 3835 2585
rect 3805 2535 3835 2565
rect 3805 2515 3810 2535
rect 3830 2515 3835 2535
rect 3805 2485 3835 2515
rect 3805 2465 3810 2485
rect 3830 2465 3835 2485
rect 3805 2435 3835 2465
rect 3805 2415 3810 2435
rect 3830 2415 3835 2435
rect 3805 2405 3835 2415
rect 3895 2685 3925 2695
rect 3895 2665 3900 2685
rect 3920 2665 3925 2685
rect 3895 2635 3925 2665
rect 3895 2615 3900 2635
rect 3920 2615 3925 2635
rect 3895 2585 3925 2615
rect 3895 2565 3900 2585
rect 3920 2565 3925 2585
rect 3895 2535 3925 2565
rect 3895 2515 3900 2535
rect 3920 2515 3925 2535
rect 3895 2485 3925 2515
rect 3895 2465 3900 2485
rect 3920 2465 3925 2485
rect 3895 2435 3925 2465
rect 3895 2415 3900 2435
rect 3920 2415 3925 2435
rect 3895 2405 3925 2415
rect 3985 2685 4015 2695
rect 3985 2665 3990 2685
rect 4010 2665 4015 2685
rect 3985 2635 4015 2665
rect 3985 2615 3990 2635
rect 4010 2615 4015 2635
rect 3985 2585 4015 2615
rect 3985 2565 3990 2585
rect 4010 2565 4015 2585
rect 3985 2535 4015 2565
rect 3985 2515 3990 2535
rect 4010 2515 4015 2535
rect 3985 2485 4015 2515
rect 3985 2465 3990 2485
rect 4010 2465 4015 2485
rect 3985 2435 4015 2465
rect 3985 2415 3990 2435
rect 4010 2415 4015 2435
rect 3985 2405 4015 2415
rect 4075 2685 4105 2695
rect 4075 2665 4080 2685
rect 4100 2665 4105 2685
rect 4075 2635 4105 2665
rect 4075 2615 4080 2635
rect 4100 2615 4105 2635
rect 4075 2585 4105 2615
rect 4075 2565 4080 2585
rect 4100 2565 4105 2585
rect 4075 2535 4105 2565
rect 4075 2515 4080 2535
rect 4100 2515 4105 2535
rect 4075 2485 4105 2515
rect 4075 2465 4080 2485
rect 4100 2465 4105 2485
rect 4075 2435 4105 2465
rect 4075 2415 4080 2435
rect 4100 2415 4105 2435
rect 4075 2405 4105 2415
rect 4165 2685 4195 2695
rect 4165 2665 4170 2685
rect 4190 2665 4195 2685
rect 4165 2635 4195 2665
rect 4165 2615 4170 2635
rect 4190 2615 4195 2635
rect 4165 2585 4195 2615
rect 4165 2565 4170 2585
rect 4190 2565 4195 2585
rect 4165 2535 4195 2565
rect 4165 2515 4170 2535
rect 4190 2515 4195 2535
rect 4165 2485 4195 2515
rect 4165 2465 4170 2485
rect 4190 2465 4195 2485
rect 4165 2435 4195 2465
rect 4165 2415 4170 2435
rect 4190 2415 4195 2435
rect 4165 2405 4195 2415
rect 4255 2685 4285 2695
rect 4255 2665 4260 2685
rect 4280 2665 4285 2685
rect 4255 2635 4285 2665
rect 4255 2615 4260 2635
rect 4280 2615 4285 2635
rect 4255 2585 4285 2615
rect 4255 2565 4260 2585
rect 4280 2565 4285 2585
rect 4255 2535 4285 2565
rect 4255 2515 4260 2535
rect 4280 2515 4285 2535
rect 4255 2485 4285 2515
rect 4255 2465 4260 2485
rect 4280 2465 4285 2485
rect 4255 2435 4285 2465
rect 4255 2415 4260 2435
rect 4280 2415 4285 2435
rect 4255 2405 4285 2415
rect 4345 2685 4375 2695
rect 4345 2665 4350 2685
rect 4370 2665 4375 2685
rect 4345 2635 4375 2665
rect 4345 2615 4350 2635
rect 4370 2615 4375 2635
rect 4345 2585 4375 2615
rect 4345 2565 4350 2585
rect 4370 2565 4375 2585
rect 4345 2535 4375 2565
rect 4345 2515 4350 2535
rect 4370 2515 4375 2535
rect 4345 2485 4375 2515
rect 4345 2465 4350 2485
rect 4370 2465 4375 2485
rect 4345 2435 4375 2465
rect 4345 2415 4350 2435
rect 4370 2415 4375 2435
rect 4345 2405 4375 2415
rect 4435 2685 4465 2695
rect 4435 2665 4440 2685
rect 4460 2665 4465 2685
rect 4435 2635 4465 2665
rect 4435 2615 4440 2635
rect 4460 2615 4465 2635
rect 4435 2585 4465 2615
rect 4435 2565 4440 2585
rect 4460 2565 4465 2585
rect 4435 2535 4465 2565
rect 4435 2515 4440 2535
rect 4460 2515 4465 2535
rect 4435 2485 4465 2515
rect 4435 2465 4440 2485
rect 4460 2465 4465 2485
rect 4435 2435 4465 2465
rect 4435 2415 4440 2435
rect 4460 2415 4465 2435
rect 4435 2405 4465 2415
rect 4525 2685 4555 2695
rect 4525 2665 4530 2685
rect 4550 2665 4555 2685
rect 4525 2635 4555 2665
rect 4525 2615 4530 2635
rect 4550 2615 4555 2635
rect 4525 2585 4555 2615
rect 4525 2565 4530 2585
rect 4550 2565 4555 2585
rect 4525 2535 4555 2565
rect 4525 2515 4530 2535
rect 4550 2515 4555 2535
rect 4525 2485 4555 2515
rect 4525 2465 4530 2485
rect 4550 2465 4555 2485
rect 4525 2435 4555 2465
rect 4525 2415 4530 2435
rect 4550 2415 4555 2435
rect 4525 2405 4555 2415
rect 4615 2685 4645 2695
rect 4615 2665 4620 2685
rect 4640 2665 4645 2685
rect 4615 2635 4645 2665
rect 4615 2615 4620 2635
rect 4640 2615 4645 2635
rect 4615 2585 4645 2615
rect 4615 2565 4620 2585
rect 4640 2565 4645 2585
rect 4615 2535 4645 2565
rect 4615 2515 4620 2535
rect 4640 2515 4645 2535
rect 4615 2485 4645 2515
rect 4615 2465 4620 2485
rect 4640 2465 4645 2485
rect 4615 2435 4645 2465
rect 4615 2415 4620 2435
rect 4640 2415 4645 2435
rect 4615 2405 4645 2415
rect 4705 2685 4735 2695
rect 4705 2665 4710 2685
rect 4730 2665 4735 2685
rect 4705 2635 4735 2665
rect 4705 2615 4710 2635
rect 4730 2615 4735 2635
rect 4705 2585 4735 2615
rect 4705 2565 4710 2585
rect 4730 2565 4735 2585
rect 4705 2535 4735 2565
rect 4705 2515 4710 2535
rect 4730 2515 4735 2535
rect 4705 2485 4735 2515
rect 4705 2465 4710 2485
rect 4730 2465 4735 2485
rect 4705 2435 4735 2465
rect 4705 2415 4710 2435
rect 4730 2415 4735 2435
rect 4705 2405 4735 2415
rect 4795 2685 4825 2695
rect 4795 2665 4800 2685
rect 4820 2665 4825 2685
rect 4795 2635 4825 2665
rect 4795 2615 4800 2635
rect 4820 2615 4825 2635
rect 4795 2585 4825 2615
rect 4795 2565 4800 2585
rect 4820 2565 4825 2585
rect 4795 2535 4825 2565
rect 4795 2515 4800 2535
rect 4820 2515 4825 2535
rect 4795 2485 4825 2515
rect 4795 2465 4800 2485
rect 4820 2465 4825 2485
rect 4795 2435 4825 2465
rect 4795 2415 4800 2435
rect 4820 2415 4825 2435
rect 4795 2405 4825 2415
rect 4885 2685 4915 2695
rect 4885 2665 4890 2685
rect 4910 2665 4915 2685
rect 4885 2635 4915 2665
rect 4885 2615 4890 2635
rect 4910 2615 4915 2635
rect 4885 2585 4915 2615
rect 4885 2565 4890 2585
rect 4910 2565 4915 2585
rect 4885 2535 4915 2565
rect 4885 2515 4890 2535
rect 4910 2515 4915 2535
rect 4885 2485 4915 2515
rect 4885 2465 4890 2485
rect 4910 2465 4915 2485
rect 4885 2435 4915 2465
rect 4885 2415 4890 2435
rect 4910 2415 4915 2435
rect 4885 2405 4915 2415
rect 4975 2685 5005 2695
rect 4975 2665 4980 2685
rect 5000 2665 5005 2685
rect 4975 2635 5005 2665
rect 4975 2615 4980 2635
rect 5000 2615 5005 2635
rect 4975 2585 5005 2615
rect 4975 2565 4980 2585
rect 5000 2565 5005 2585
rect 4975 2535 5005 2565
rect 4975 2515 4980 2535
rect 5000 2515 5005 2535
rect 4975 2485 5005 2515
rect 4975 2465 4980 2485
rect 5000 2465 5005 2485
rect 4975 2435 5005 2465
rect 4975 2415 4980 2435
rect 5000 2415 5005 2435
rect 4975 2405 5005 2415
rect 5065 2685 5095 2695
rect 5065 2665 5070 2685
rect 5090 2665 5095 2685
rect 5065 2635 5095 2665
rect 5065 2615 5070 2635
rect 5090 2615 5095 2635
rect 5065 2585 5095 2615
rect 5065 2565 5070 2585
rect 5090 2565 5095 2585
rect 5065 2535 5095 2565
rect 5065 2515 5070 2535
rect 5090 2515 5095 2535
rect 5065 2485 5095 2515
rect 5065 2465 5070 2485
rect 5090 2465 5095 2485
rect 5065 2435 5095 2465
rect 5065 2415 5070 2435
rect 5090 2415 5095 2435
rect 5065 2405 5095 2415
rect 5155 2685 5185 2695
rect 5155 2665 5160 2685
rect 5180 2665 5185 2685
rect 5155 2635 5185 2665
rect 5155 2615 5160 2635
rect 5180 2615 5185 2635
rect 5155 2585 5185 2615
rect 5155 2565 5160 2585
rect 5180 2565 5185 2585
rect 5155 2535 5185 2565
rect 5155 2515 5160 2535
rect 5180 2515 5185 2535
rect 5155 2485 5185 2515
rect 5155 2465 5160 2485
rect 5180 2465 5185 2485
rect 5155 2435 5185 2465
rect 5155 2415 5160 2435
rect 5180 2415 5185 2435
rect 5155 2405 5185 2415
rect 2820 2385 2840 2405
rect 2910 2385 2930 2405
rect 3090 2385 3110 2405
rect 2810 2375 2850 2385
rect 2810 2355 2820 2375
rect 2840 2355 2850 2375
rect 2810 2345 2850 2355
rect 2900 2375 2940 2385
rect 2900 2355 2910 2375
rect 2930 2355 2940 2375
rect 2900 2345 2940 2355
rect 2990 2370 3030 2380
rect 2990 2350 3000 2370
rect 3020 2350 3030 2370
rect 2625 2315 2655 2345
rect 2990 2340 3030 2350
rect 3080 2375 3120 2385
rect 3080 2355 3090 2375
rect 3110 2355 3120 2375
rect 3080 2345 3120 2355
rect 3270 2340 3290 2405
rect 3450 2385 3470 2405
rect 3440 2375 3480 2385
rect 3440 2355 3450 2375
rect 3470 2355 3480 2375
rect 3440 2345 3480 2355
rect 3630 2340 3650 2405
rect 3810 2385 3830 2405
rect 3990 2385 4010 2405
rect 4170 2385 4190 2405
rect 3800 2375 3840 2385
rect 3800 2355 3810 2375
rect 3830 2355 3840 2375
rect 3800 2345 3840 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3980 2375 4020 2385
rect 3980 2355 3990 2375
rect 4010 2355 4020 2375
rect 3980 2345 4020 2355
rect 4150 2375 4190 2385
rect 4150 2355 4160 2375
rect 4180 2355 4190 2375
rect 4150 2345 4190 2355
rect 4350 2340 4370 2405
rect 4530 2385 4550 2405
rect 4520 2375 4560 2385
rect 4520 2355 4530 2375
rect 4550 2355 4560 2375
rect 4520 2345 4560 2355
rect 4710 2340 4730 2405
rect 4890 2385 4910 2405
rect 5070 2385 5090 2405
rect 5160 2385 5180 2405
rect 4880 2375 4920 2385
rect 4880 2355 4890 2375
rect 4910 2355 4920 2375
rect 4880 2345 4920 2355
rect 5060 2375 5100 2385
rect 5060 2355 5070 2375
rect 5090 2355 5100 2375
rect 5060 2345 5100 2355
rect 5150 2375 5190 2385
rect 5150 2355 5160 2375
rect 5180 2355 5190 2375
rect 5150 2345 5190 2355
rect 3260 2330 3300 2340
rect 3260 2310 3270 2330
rect 3290 2310 3300 2330
rect 3260 2300 3300 2310
rect 3620 2330 3660 2340
rect 3620 2310 3630 2330
rect 3650 2310 3660 2330
rect 3620 2300 3660 2310
rect 4340 2330 4380 2340
rect 4340 2310 4350 2330
rect 4370 2310 4380 2330
rect 4340 2300 4380 2310
rect 4700 2330 4740 2340
rect 4700 2310 4710 2330
rect 4730 2310 4740 2330
rect 4700 2300 4740 2310
rect 2740 2260 2770 2290
rect 3440 2285 3480 2295
rect 3440 2265 3450 2285
rect 3470 2265 3480 2285
rect 3440 2255 3480 2265
rect 4520 2285 4560 2295
rect 4520 2265 4530 2285
rect 4550 2265 4560 2285
rect 4520 2255 4560 2265
rect 5255 2260 5285 2290
rect 2430 2215 2460 2245
rect 3085 2215 3115 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3265 2120 3295 2150
rect 4080 2115 4110 2145
rect 5300 2115 5330 2145
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 4135 2090 4175 2100
rect 4135 2070 4145 2090
rect 4165 2070 4175 2090
rect 4135 2060 4175 2070
rect 4255 2090 4295 2100
rect 4255 2070 4265 2090
rect 4285 2070 4295 2090
rect 4255 2060 4295 2070
rect 4375 2090 4415 2100
rect 4375 2070 4385 2090
rect 4405 2070 4415 2090
rect 4375 2060 4415 2070
rect 4495 2090 4535 2100
rect 4495 2070 4505 2090
rect 4525 2070 4535 2090
rect 4495 2060 4535 2070
rect 4615 2090 4655 2100
rect 4615 2070 4625 2090
rect 4645 2070 4655 2090
rect 4615 2060 4655 2070
rect 4735 2090 4775 2100
rect 4735 2070 4745 2090
rect 4765 2070 4775 2090
rect 4735 2060 4775 2070
rect 4855 2090 4895 2100
rect 4855 2070 4865 2090
rect 4885 2070 4895 2090
rect 4855 2060 4895 2070
rect 4975 2090 5015 2100
rect 4975 2070 4985 2090
rect 5005 2070 5015 2090
rect 4975 2060 5015 2070
rect 5095 2090 5135 2100
rect 5095 2070 5105 2090
rect 5125 2070 5135 2090
rect 5095 2060 5135 2070
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect 2745 2045 2785 2055
rect 2745 2025 2755 2045
rect 2775 2025 2785 2045
rect 2745 2015 2785 2025
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2015
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3945 2045 3985 2055
rect 3945 2025 3955 2045
rect 3975 2025 3985 2045
rect 3945 2015 3985 2025
rect 4015 2045 4055 2055
rect 4015 2025 4025 2045
rect 4045 2025 4055 2045
rect 4015 2015 4055 2025
rect 4075 2045 4115 2055
rect 4075 2025 4085 2045
rect 4105 2025 4115 2045
rect 4075 2015 4115 2025
rect 3895 1995 3915 2015
rect 3955 1995 3975 2015
rect 4025 1995 4045 2015
rect 4085 1995 4105 2015
rect 4145 1995 4165 2060
rect 4265 1995 4285 2060
rect 4385 1995 4405 2060
rect 4435 2045 4475 2055
rect 4435 2025 4445 2045
rect 4465 2025 4475 2045
rect 4435 2015 4475 2025
rect 4445 1995 4465 2015
rect 4505 1995 4525 2060
rect 4625 1995 4645 2060
rect 4745 1995 4765 2060
rect 4795 2045 4835 2055
rect 4795 2025 4805 2045
rect 4825 2025 4835 2045
rect 4795 2015 4835 2025
rect 4805 1995 4825 2015
rect 4865 1995 4885 2060
rect 4985 1995 5005 2060
rect 5105 1995 5125 2060
rect 5155 2045 5195 2055
rect 5155 2025 5165 2045
rect 5185 2025 5195 2045
rect 5155 2015 5195 2025
rect 5215 2045 5255 2055
rect 5215 2025 5225 2045
rect 5245 2025 5255 2045
rect 5215 2015 5255 2025
rect 5165 1995 5185 2015
rect 5225 1995 5245 2015
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 3980 1995
rect 3950 1965 3955 1985
rect 3975 1965 3980 1985
rect 3950 1935 3980 1965
rect 3950 1915 3955 1935
rect 3975 1915 3980 1935
rect 3950 1905 3980 1915
rect 4020 1985 4050 1995
rect 4020 1965 4025 1985
rect 4045 1965 4050 1985
rect 4020 1935 4050 1965
rect 4020 1915 4025 1935
rect 4045 1915 4050 1935
rect 4020 1905 4050 1915
rect 4080 1985 4110 1995
rect 4080 1965 4085 1985
rect 4105 1965 4110 1985
rect 4080 1935 4110 1965
rect 4080 1915 4085 1935
rect 4105 1915 4110 1935
rect 4080 1905 4110 1915
rect 4140 1985 4170 1995
rect 4140 1965 4145 1985
rect 4165 1965 4170 1985
rect 4140 1935 4170 1965
rect 4140 1915 4145 1935
rect 4165 1915 4170 1935
rect 4140 1905 4170 1915
rect 4200 1985 4230 1995
rect 4200 1965 4205 1985
rect 4225 1965 4230 1985
rect 4200 1935 4230 1965
rect 4200 1915 4205 1935
rect 4225 1915 4230 1935
rect 4200 1905 4230 1915
rect 4260 1985 4290 1995
rect 4260 1965 4265 1985
rect 4285 1965 4290 1985
rect 4260 1935 4290 1965
rect 4260 1915 4265 1935
rect 4285 1915 4290 1935
rect 4260 1905 4290 1915
rect 4320 1985 4350 1995
rect 4320 1965 4325 1985
rect 4345 1965 4350 1985
rect 4320 1935 4350 1965
rect 4320 1915 4325 1935
rect 4345 1915 4350 1935
rect 4320 1905 4350 1915
rect 4380 1985 4410 1995
rect 4380 1965 4385 1985
rect 4405 1965 4410 1985
rect 4380 1935 4410 1965
rect 4380 1915 4385 1935
rect 4405 1915 4410 1935
rect 4380 1905 4410 1915
rect 4440 1985 4470 1995
rect 4440 1965 4445 1985
rect 4465 1965 4470 1985
rect 4440 1935 4470 1965
rect 4440 1915 4445 1935
rect 4465 1915 4470 1935
rect 4440 1905 4470 1915
rect 4500 1985 4530 1995
rect 4500 1965 4505 1985
rect 4525 1965 4530 1985
rect 4500 1935 4530 1965
rect 4500 1915 4505 1935
rect 4525 1915 4530 1935
rect 4500 1905 4530 1915
rect 4560 1985 4590 1995
rect 4560 1965 4565 1985
rect 4585 1965 4590 1985
rect 4560 1935 4590 1965
rect 4560 1915 4565 1935
rect 4585 1915 4590 1935
rect 4560 1905 4590 1915
rect 4620 1985 4650 1995
rect 4620 1965 4625 1985
rect 4645 1965 4650 1985
rect 4620 1935 4650 1965
rect 4620 1915 4625 1935
rect 4645 1915 4650 1935
rect 4620 1905 4650 1915
rect 4680 1985 4710 1995
rect 4680 1965 4685 1985
rect 4705 1965 4710 1985
rect 4680 1935 4710 1965
rect 4680 1915 4685 1935
rect 4705 1915 4710 1935
rect 4680 1905 4710 1915
rect 4740 1985 4770 1995
rect 4740 1965 4745 1985
rect 4765 1965 4770 1985
rect 4740 1935 4770 1965
rect 4740 1915 4745 1935
rect 4765 1915 4770 1935
rect 4740 1905 4770 1915
rect 4800 1985 4830 1995
rect 4800 1965 4805 1985
rect 4825 1965 4830 1985
rect 4800 1935 4830 1965
rect 4800 1915 4805 1935
rect 4825 1915 4830 1935
rect 4800 1905 4830 1915
rect 4860 1985 4890 1995
rect 4860 1965 4865 1985
rect 4885 1965 4890 1985
rect 4860 1935 4890 1965
rect 4860 1915 4865 1935
rect 4885 1915 4890 1935
rect 4860 1905 4890 1915
rect 4920 1985 4950 1995
rect 4920 1965 4925 1985
rect 4945 1965 4950 1985
rect 4920 1935 4950 1965
rect 4920 1915 4925 1935
rect 4945 1915 4950 1935
rect 4920 1905 4950 1915
rect 4980 1985 5010 1995
rect 4980 1965 4985 1985
rect 5005 1965 5010 1985
rect 4980 1935 5010 1965
rect 4980 1915 4985 1935
rect 5005 1915 5010 1935
rect 4980 1905 5010 1915
rect 5040 1985 5070 1995
rect 5040 1965 5045 1985
rect 5065 1965 5070 1985
rect 5040 1935 5070 1965
rect 5040 1915 5045 1935
rect 5065 1915 5070 1935
rect 5040 1905 5070 1915
rect 5100 1985 5130 1995
rect 5100 1965 5105 1985
rect 5125 1965 5130 1985
rect 5100 1935 5130 1965
rect 5100 1915 5105 1935
rect 5125 1915 5130 1935
rect 5100 1905 5130 1915
rect 5160 1985 5190 1995
rect 5160 1965 5165 1985
rect 5185 1965 5190 1985
rect 5160 1935 5190 1965
rect 5160 1915 5165 1935
rect 5185 1915 5190 1935
rect 5160 1905 5190 1915
rect 5220 1985 5250 1995
rect 5220 1965 5225 1985
rect 5245 1965 5250 1985
rect 5220 1935 5250 1965
rect 5220 1915 5225 1935
rect 5245 1915 5250 1935
rect 5220 1905 5250 1915
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 4205 1885 4225 1905
rect 4325 1885 4345 1905
rect 4565 1885 4585 1905
rect 4685 1885 4705 1905
rect 4925 1885 4945 1905
rect 5045 1885 5065 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 4105 1875 4145 1885
rect 4105 1855 4115 1875
rect 4135 1855 4145 1875
rect 4105 1845 4145 1855
rect 4195 1875 4235 1885
rect 4195 1855 4205 1875
rect 4225 1855 4235 1875
rect 4195 1845 4235 1855
rect 4315 1875 4355 1885
rect 4315 1855 4325 1875
rect 4345 1855 4355 1875
rect 4315 1845 4355 1855
rect 4435 1875 4475 1885
rect 4435 1855 4445 1875
rect 4465 1855 4475 1875
rect 4435 1845 4475 1855
rect 4555 1875 4595 1885
rect 4555 1855 4565 1875
rect 4585 1855 4595 1875
rect 4555 1845 4595 1855
rect 4675 1875 4715 1885
rect 4675 1855 4685 1875
rect 4705 1855 4715 1875
rect 4675 1845 4715 1855
rect 4795 1875 4835 1885
rect 4795 1855 4805 1875
rect 4825 1855 4835 1875
rect 4795 1845 4835 1855
rect 4915 1875 4955 1885
rect 4915 1855 4925 1875
rect 4945 1855 4955 1875
rect 4915 1845 4955 1855
rect 5035 1875 5075 1885
rect 5035 1855 5045 1875
rect 5065 1855 5075 1875
rect 5035 1845 5075 1855
rect 5125 1875 5165 1885
rect 5125 1855 5135 1875
rect 5155 1855 5165 1875
rect 5125 1845 5165 1855
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4105 1785 4145 1825
rect 4195 1815 4235 1825
rect 4195 1795 4205 1815
rect 4225 1795 4235 1815
rect 4195 1785 4235 1795
rect 4435 1785 4475 1825
rect 4555 1815 4595 1825
rect 4555 1795 4565 1815
rect 4585 1795 4595 1815
rect 4555 1785 4595 1795
rect 4795 1785 4835 1825
rect 4915 1815 4955 1825
rect 4915 1795 4925 1815
rect 4945 1795 4955 1815
rect 4915 1785 4955 1795
rect 5125 1785 5165 1825
rect 5345 1790 5375 1820
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4195 1755 4235 1765
rect 4195 1735 4205 1755
rect 4225 1735 4235 1755
rect 4195 1725 4235 1735
rect 4435 1755 4475 1765
rect 4435 1735 4445 1755
rect 4465 1735 4475 1755
rect 4435 1725 4475 1735
rect 4675 1755 4715 1765
rect 4675 1735 4685 1755
rect 4705 1735 4715 1755
rect 4675 1725 4715 1735
rect 4735 1755 4775 1765
rect 4735 1735 4745 1755
rect 4765 1735 4775 1755
rect 4735 1725 4775 1735
rect 5255 1730 5285 1760
rect 3165 1710 3205 1720
rect 2155 1680 2185 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4205 1660 4225 1725
rect 4315 1710 4355 1720
rect 4315 1690 4325 1710
rect 4345 1690 4355 1710
rect 4315 1680 4355 1690
rect 4325 1660 4345 1680
rect 4445 1660 4465 1725
rect 4555 1710 4595 1720
rect 4555 1690 4565 1710
rect 4585 1690 4595 1710
rect 4555 1680 4595 1690
rect 4565 1660 4585 1680
rect 4685 1660 4705 1725
rect 4795 1710 4835 1720
rect 4795 1690 4805 1710
rect 4825 1690 4835 1710
rect 4795 1680 4835 1690
rect 4805 1660 4825 1680
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 4200 1650 4230 1660
rect 4200 1630 4205 1650
rect 4225 1630 4230 1650
rect 4200 1620 4230 1630
rect 4260 1650 4290 1660
rect 4260 1630 4265 1650
rect 4285 1630 4290 1650
rect 4260 1620 4290 1630
rect 4320 1650 4350 1660
rect 4320 1630 4325 1650
rect 4345 1630 4350 1650
rect 4320 1620 4350 1630
rect 4380 1650 4410 1660
rect 4380 1630 4385 1650
rect 4405 1630 4410 1650
rect 4380 1620 4410 1630
rect 4440 1650 4470 1660
rect 4440 1630 4445 1650
rect 4465 1630 4470 1650
rect 4440 1620 4470 1630
rect 4500 1650 4530 1660
rect 4500 1630 4505 1650
rect 4525 1630 4530 1650
rect 4500 1620 4530 1630
rect 4560 1650 4590 1660
rect 4560 1630 4565 1650
rect 4585 1630 4590 1650
rect 4560 1620 4590 1630
rect 4620 1650 4650 1660
rect 4620 1630 4625 1650
rect 4645 1630 4650 1650
rect 4620 1620 4650 1630
rect 4680 1650 4710 1660
rect 4680 1630 4685 1650
rect 4705 1630 4710 1650
rect 4680 1620 4710 1630
rect 4740 1650 4770 1660
rect 4740 1630 4745 1650
rect 4765 1630 4770 1650
rect 4740 1620 4770 1630
rect 4800 1650 4830 1660
rect 4800 1630 4805 1650
rect 4825 1630 4830 1650
rect 4800 1620 4830 1630
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4265 1550 4285 1620
rect 4385 1550 4405 1620
rect 4505 1550 4525 1620
rect 4625 1550 4645 1620
rect 4745 1550 4765 1620
rect 4795 1590 4835 1600
rect 4795 1570 4805 1590
rect 4825 1570 4835 1590
rect 4795 1560 4835 1570
rect 5395 1565 5425 1595
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4255 1540 4295 1550
rect 4255 1520 4265 1540
rect 4285 1520 4295 1540
rect 4255 1510 4295 1520
rect 4375 1540 4415 1550
rect 4375 1520 4385 1540
rect 4405 1520 4415 1540
rect 4375 1510 4415 1520
rect 4495 1540 4535 1550
rect 4495 1520 4505 1540
rect 4525 1520 4535 1540
rect 4495 1510 4535 1520
rect 4615 1540 4655 1550
rect 4615 1520 4625 1540
rect 4645 1520 4655 1540
rect 4615 1510 4655 1520
rect 4735 1540 4775 1550
rect 4735 1520 4745 1540
rect 4765 1520 4775 1540
rect 4735 1510 4775 1520
rect 2835 1485 2875 1495
rect 2835 1465 2845 1485
rect 2865 1465 2875 1485
rect 2835 1455 2875 1465
rect 3915 1485 3955 1495
rect 3915 1465 3925 1485
rect 3945 1465 3955 1485
rect 3915 1455 3955 1465
rect 4045 1485 4085 1495
rect 4045 1465 4055 1485
rect 4075 1465 4085 1485
rect 4045 1455 4085 1465
rect 5125 1485 5165 1495
rect 5125 1465 5135 1485
rect 5155 1465 5165 1485
rect 5125 1455 5165 1465
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1445 2870 1455
rect 2840 1425 2845 1445
rect 2865 1425 2870 1445
rect 2840 1395 2870 1425
rect 2840 1375 2845 1395
rect 2865 1375 2870 1395
rect 2840 1345 2870 1375
rect 2840 1325 2845 1345
rect 2865 1325 2870 1345
rect 2840 1295 2870 1325
rect 2840 1275 2845 1295
rect 2865 1275 2870 1295
rect 2840 1245 2870 1275
rect 2840 1225 2845 1245
rect 2865 1225 2870 1245
rect 2840 1215 2870 1225
rect 3380 1445 3410 1455
rect 3380 1425 3385 1445
rect 3405 1425 3410 1445
rect 3380 1395 3410 1425
rect 3380 1375 3385 1395
rect 3405 1375 3410 1395
rect 3380 1345 3410 1375
rect 3380 1325 3385 1345
rect 3405 1325 3410 1345
rect 3380 1295 3410 1325
rect 3380 1275 3385 1295
rect 3405 1275 3410 1295
rect 3380 1245 3410 1275
rect 3380 1225 3385 1245
rect 3405 1225 3410 1245
rect 3380 1215 3410 1225
rect 3920 1445 3950 1455
rect 3920 1425 3925 1445
rect 3945 1425 3950 1445
rect 3920 1395 3950 1425
rect 3920 1375 3925 1395
rect 3945 1375 3950 1395
rect 3920 1345 3950 1375
rect 3920 1325 3925 1345
rect 3945 1325 3950 1345
rect 3920 1295 3950 1325
rect 3920 1275 3925 1295
rect 3945 1275 3950 1295
rect 3920 1245 3950 1275
rect 3920 1225 3925 1245
rect 3945 1225 3950 1245
rect 3920 1215 3950 1225
rect 4050 1445 4080 1455
rect 4050 1425 4055 1445
rect 4075 1425 4080 1445
rect 4050 1395 4080 1425
rect 4050 1375 4055 1395
rect 4075 1375 4080 1395
rect 4050 1345 4080 1375
rect 4050 1325 4055 1345
rect 4075 1325 4080 1345
rect 4050 1295 4080 1325
rect 4050 1275 4055 1295
rect 4075 1275 4080 1295
rect 4050 1245 4080 1275
rect 4050 1225 4055 1245
rect 4075 1225 4080 1245
rect 4050 1215 4080 1225
rect 4590 1445 4620 1455
rect 4590 1425 4595 1445
rect 4615 1425 4620 1445
rect 4590 1395 4620 1425
rect 4590 1375 4595 1395
rect 4615 1375 4620 1395
rect 4590 1345 4620 1375
rect 4590 1325 4595 1345
rect 4615 1325 4620 1345
rect 4590 1295 4620 1325
rect 4590 1275 4595 1295
rect 4615 1275 4620 1295
rect 4590 1245 4620 1275
rect 4590 1225 4595 1245
rect 4615 1225 4620 1245
rect 4590 1215 4620 1225
rect 5130 1445 5160 1455
rect 5130 1425 5135 1445
rect 5155 1425 5160 1445
rect 5130 1395 5160 1425
rect 5130 1375 5135 1395
rect 5155 1375 5160 1395
rect 5130 1345 5160 1375
rect 5130 1325 5135 1345
rect 5155 1325 5160 1345
rect 5130 1295 5160 1325
rect 5130 1275 5135 1295
rect 5155 1275 5160 1295
rect 5130 1245 5160 1275
rect 5130 1225 5135 1245
rect 5155 1225 5160 1245
rect 5130 1215 5160 1225
rect 3385 1195 3405 1215
rect 4595 1195 4615 1215
rect 3375 1185 3415 1195
rect 3375 1165 3385 1185
rect 3405 1165 3415 1185
rect 3375 1155 3415 1165
rect 4585 1185 4625 1195
rect 4585 1165 4595 1185
rect 4615 1165 4625 1185
rect 4585 1155 4625 1165
rect 2940 1125 2980 1135
rect 2940 1105 2950 1125
rect 2970 1105 2980 1125
rect 2940 1095 2980 1105
rect 3020 1125 3060 1135
rect 3020 1105 3030 1125
rect 3050 1105 3060 1125
rect 3020 1095 3060 1105
rect 3100 1125 3140 1135
rect 3100 1105 3110 1125
rect 3130 1105 3140 1125
rect 3100 1095 3140 1105
rect 3180 1125 3220 1135
rect 3180 1105 3190 1125
rect 3210 1105 3220 1125
rect 3180 1095 3220 1105
rect 3260 1125 3300 1135
rect 3260 1105 3270 1125
rect 3290 1105 3300 1125
rect 3260 1095 3300 1105
rect 3340 1125 3380 1135
rect 3340 1105 3350 1125
rect 3370 1105 3380 1125
rect 3340 1095 3380 1105
rect 3420 1125 3460 1135
rect 3420 1105 3430 1125
rect 3450 1105 3460 1125
rect 3420 1095 3460 1105
rect 3500 1125 3540 1135
rect 3500 1105 3510 1125
rect 3530 1105 3540 1125
rect 3500 1095 3540 1105
rect 3580 1125 3620 1135
rect 3580 1105 3590 1125
rect 3610 1105 3620 1125
rect 3580 1095 3620 1105
rect 3660 1125 3700 1135
rect 3660 1105 3670 1125
rect 3690 1105 3700 1125
rect 3660 1095 3700 1105
rect 3740 1125 3780 1135
rect 3740 1105 3750 1125
rect 3770 1105 3780 1125
rect 3740 1095 3780 1105
rect 3820 1125 3860 1135
rect 3820 1105 3830 1125
rect 3850 1105 3860 1125
rect 3820 1095 3860 1105
rect 3900 1125 3940 1135
rect 3900 1105 3910 1125
rect 3930 1105 3940 1125
rect 3900 1095 3940 1105
rect 3980 1125 4020 1135
rect 3980 1105 3990 1125
rect 4010 1105 4020 1125
rect 3980 1095 4020 1105
rect 4060 1125 4100 1135
rect 4060 1105 4070 1125
rect 4090 1105 4100 1125
rect 4060 1095 4100 1105
rect 4140 1125 4180 1135
rect 4140 1105 4150 1125
rect 4170 1105 4180 1125
rect 4140 1095 4180 1105
rect 4220 1125 4260 1135
rect 4220 1105 4230 1125
rect 4250 1105 4260 1125
rect 4220 1095 4260 1105
rect 4300 1125 4340 1135
rect 4300 1105 4310 1125
rect 4330 1105 4340 1125
rect 4300 1095 4340 1105
rect 4380 1125 4420 1135
rect 4380 1105 4390 1125
rect 4410 1105 4420 1125
rect 4380 1095 4420 1105
rect 4460 1125 4500 1135
rect 4460 1105 4470 1125
rect 4490 1105 4500 1125
rect 4460 1095 4500 1105
rect 4540 1125 4580 1135
rect 4540 1105 4550 1125
rect 4570 1105 4580 1125
rect 4540 1095 4580 1105
rect 4620 1125 4660 1135
rect 4620 1105 4630 1125
rect 4650 1105 4660 1125
rect 4620 1095 4660 1105
rect 4700 1125 4740 1135
rect 4700 1105 4710 1125
rect 4730 1105 4740 1125
rect 4700 1095 4740 1105
rect 4780 1125 4820 1135
rect 4780 1105 4790 1125
rect 4810 1105 4820 1125
rect 4780 1095 4820 1105
rect 4860 1125 4900 1135
rect 4860 1105 4870 1125
rect 4890 1105 4900 1125
rect 4860 1095 4900 1105
rect 4940 1125 4980 1135
rect 4940 1105 4950 1125
rect 4970 1105 4980 1125
rect 4940 1095 4980 1105
rect 2950 1075 2970 1095
rect 3990 1075 4010 1095
rect 2945 1065 2975 1075
rect 2945 1050 2950 1065
rect 2930 1045 2950 1050
rect 2970 1045 2975 1065
rect 2430 1000 2460 1030
rect 2625 1015 2655 1045
rect 2905 1040 2975 1045
rect 2905 1020 2910 1040
rect 2930 1020 2975 1040
rect 2905 1015 2975 1020
rect 2930 1010 2950 1015
rect 2945 995 2950 1010
rect 2970 995 2975 1015
rect 2945 985 2975 995
rect 3985 1065 4015 1075
rect 3985 1045 3990 1065
rect 4010 1045 4015 1065
rect 3985 1015 4015 1045
rect 3985 995 3990 1015
rect 4010 995 4015 1015
rect 3985 985 4015 995
rect 5025 1065 5055 1075
rect 5025 1045 5030 1065
rect 5050 1050 5055 1065
rect 5050 1045 5095 1050
rect 5025 1040 5095 1045
rect 5025 1020 5065 1040
rect 5085 1020 5095 1040
rect 5025 1015 5095 1020
rect 5025 995 5030 1015
rect 5050 1010 5095 1015
rect 5050 995 5055 1010
rect 5025 985 5055 995
rect 2990 930 3030 940
rect 2990 910 3000 930
rect 3020 910 3030 930
rect 2990 900 3030 910
rect 3170 930 3210 940
rect 3170 910 3180 930
rect 3200 910 3210 930
rect 3170 900 3210 910
rect 3350 930 3390 940
rect 3350 910 3360 930
rect 3380 910 3390 930
rect 3350 900 3390 910
rect 3530 930 3570 940
rect 3530 910 3540 930
rect 3560 910 3570 930
rect 3530 900 3570 910
rect 3710 930 3750 940
rect 3710 910 3720 930
rect 3740 910 3750 930
rect 3710 900 3750 910
rect 3890 930 3930 940
rect 3890 910 3900 930
rect 3920 910 3930 930
rect 3890 900 3930 910
rect 4070 930 4110 940
rect 4070 910 4080 930
rect 4100 910 4110 930
rect 4070 900 4110 910
rect 4250 930 4290 940
rect 4250 910 4260 930
rect 4280 910 4290 930
rect 4250 900 4290 910
rect 4430 930 4470 940
rect 4430 910 4440 930
rect 4460 910 4470 930
rect 4430 900 4470 910
rect 4610 930 4650 940
rect 4610 910 4620 930
rect 4640 910 4650 930
rect 4610 900 4650 910
rect 4790 930 4830 940
rect 4790 910 4800 930
rect 4820 910 4830 930
rect 4790 900 4830 910
rect 4970 930 5010 940
rect 4970 910 4980 930
rect 5000 910 5010 930
rect 4970 900 5010 910
rect 3000 880 3020 900
rect 3180 880 3200 900
rect 3360 880 3380 900
rect 3540 880 3560 900
rect 3720 880 3740 900
rect 3900 880 3920 900
rect 4080 880 4100 900
rect 4260 880 4280 900
rect 4440 880 4460 900
rect 4620 880 4640 900
rect 4800 880 4820 900
rect 4980 880 5000 900
rect 2995 870 3025 880
rect 2995 850 3000 870
rect 3020 850 3025 870
rect 2995 820 3025 850
rect 2995 800 3000 820
rect 3020 800 3025 820
rect 2995 790 3025 800
rect 3085 870 3115 880
rect 3085 850 3090 870
rect 3110 850 3115 870
rect 3085 820 3115 850
rect 3085 800 3090 820
rect 3110 800 3115 820
rect 3085 790 3115 800
rect 3175 870 3205 880
rect 3175 850 3180 870
rect 3200 850 3205 870
rect 3175 820 3205 850
rect 3175 800 3180 820
rect 3200 800 3205 820
rect 3175 790 3205 800
rect 3265 870 3295 880
rect 3265 850 3270 870
rect 3290 850 3295 870
rect 3265 820 3295 850
rect 3265 800 3270 820
rect 3290 800 3295 820
rect 3265 790 3295 800
rect 3355 870 3385 880
rect 3355 850 3360 870
rect 3380 850 3385 870
rect 3355 820 3385 850
rect 3355 800 3360 820
rect 3380 800 3385 820
rect 3355 790 3385 800
rect 3445 870 3475 880
rect 3445 850 3450 870
rect 3470 850 3475 870
rect 3445 820 3475 850
rect 3445 800 3450 820
rect 3470 800 3475 820
rect 3445 790 3475 800
rect 3535 870 3565 880
rect 3535 850 3540 870
rect 3560 850 3565 870
rect 3535 820 3565 850
rect 3535 800 3540 820
rect 3560 800 3565 820
rect 3535 790 3565 800
rect 3625 870 3655 880
rect 3625 850 3630 870
rect 3650 850 3655 870
rect 3625 820 3655 850
rect 3625 800 3630 820
rect 3650 800 3655 820
rect 3625 790 3655 800
rect 3715 870 3745 880
rect 3715 850 3720 870
rect 3740 850 3745 870
rect 3715 820 3745 850
rect 3715 800 3720 820
rect 3740 800 3745 820
rect 3715 790 3745 800
rect 3805 870 3835 880
rect 3805 850 3810 870
rect 3830 850 3835 870
rect 3805 820 3835 850
rect 3805 800 3810 820
rect 3830 800 3835 820
rect 3805 790 3835 800
rect 3895 870 3925 880
rect 3895 850 3900 870
rect 3920 850 3925 870
rect 3895 820 3925 850
rect 3895 800 3900 820
rect 3920 800 3925 820
rect 3895 790 3925 800
rect 3985 870 4015 880
rect 3985 850 3990 870
rect 4010 850 4015 870
rect 3985 820 4015 850
rect 3985 800 3990 820
rect 4010 800 4015 820
rect 3985 790 4015 800
rect 4075 870 4105 880
rect 4075 850 4080 870
rect 4100 850 4105 870
rect 4075 820 4105 850
rect 4075 800 4080 820
rect 4100 800 4105 820
rect 4075 790 4105 800
rect 4165 870 4195 880
rect 4165 850 4170 870
rect 4190 850 4195 870
rect 4165 820 4195 850
rect 4165 800 4170 820
rect 4190 800 4195 820
rect 4165 790 4195 800
rect 4255 870 4285 880
rect 4255 850 4260 870
rect 4280 850 4285 870
rect 4255 820 4285 850
rect 4255 800 4260 820
rect 4280 800 4285 820
rect 4255 790 4285 800
rect 4345 870 4375 880
rect 4345 850 4350 870
rect 4370 850 4375 870
rect 4345 820 4375 850
rect 4345 800 4350 820
rect 4370 800 4375 820
rect 4345 790 4375 800
rect 4435 870 4465 880
rect 4435 850 4440 870
rect 4460 850 4465 870
rect 4435 820 4465 850
rect 4435 800 4440 820
rect 4460 800 4465 820
rect 4435 790 4465 800
rect 4525 870 4555 880
rect 4525 850 4530 870
rect 4550 850 4555 870
rect 4525 820 4555 850
rect 4525 800 4530 820
rect 4550 800 4555 820
rect 4525 790 4555 800
rect 4615 870 4645 880
rect 4615 850 4620 870
rect 4640 850 4645 870
rect 4615 820 4645 850
rect 4615 800 4620 820
rect 4640 800 4645 820
rect 4615 790 4645 800
rect 4705 870 4735 880
rect 4705 850 4710 870
rect 4730 850 4735 870
rect 4705 820 4735 850
rect 4705 800 4710 820
rect 4730 800 4735 820
rect 4705 790 4735 800
rect 4795 870 4825 880
rect 4795 850 4800 870
rect 4820 850 4825 870
rect 4795 820 4825 850
rect 4795 800 4800 820
rect 4820 800 4825 820
rect 4795 790 4825 800
rect 4885 870 4915 880
rect 4885 850 4890 870
rect 4910 850 4915 870
rect 4885 820 4915 850
rect 4885 800 4890 820
rect 4910 800 4915 820
rect 4885 790 4915 800
rect 4975 870 5005 880
rect 4975 850 4980 870
rect 5000 850 5005 870
rect 4975 820 5005 850
rect 4975 800 4980 820
rect 5000 800 5005 820
rect 4975 790 5005 800
rect 3090 755 3110 790
rect 3270 770 3290 790
rect 3450 770 3470 790
rect 3630 770 3650 790
rect 3810 770 3830 790
rect 3990 770 4010 790
rect 4170 770 4190 790
rect 4350 770 4370 790
rect 4530 770 4550 790
rect 4710 770 4730 790
rect 4890 770 4910 790
rect 3260 760 3300 770
rect 2525 720 2555 750
rect 3080 745 3120 755
rect 3080 725 3090 745
rect 3110 725 3120 745
rect 3260 740 3270 760
rect 3290 740 3300 760
rect 3260 730 3300 740
rect 3440 760 3480 770
rect 3440 740 3450 760
rect 3470 740 3480 760
rect 3440 730 3480 740
rect 3620 760 3660 770
rect 3620 740 3630 760
rect 3650 740 3660 760
rect 3620 730 3660 740
rect 3800 760 3840 770
rect 3800 740 3810 760
rect 3830 740 3840 760
rect 3800 730 3840 740
rect 3980 760 4020 770
rect 3980 740 3990 760
rect 4010 740 4020 760
rect 3980 730 4020 740
rect 4160 760 4200 770
rect 4160 740 4170 760
rect 4190 740 4200 760
rect 4160 730 4200 740
rect 4340 760 4380 770
rect 4340 740 4350 760
rect 4370 740 4380 760
rect 4340 730 4380 740
rect 4520 760 4560 770
rect 4520 740 4530 760
rect 4550 740 4560 760
rect 4520 730 4560 740
rect 4700 760 4740 770
rect 4700 740 4710 760
rect 4730 740 4740 760
rect 4700 730 4740 740
rect 4880 760 4920 770
rect 4880 740 4890 760
rect 4910 740 4920 760
rect 4880 730 4920 740
rect 3080 715 3120 725
rect 3445 680 3475 710
rect 3805 680 3835 710
rect 4165 680 4195 710
<< viali >>
rect 50 3175 75 3200
rect 1255 3170 1280 3195
rect 50 3115 75 3140
rect 1255 3110 1280 3135
rect 50 3035 75 3060
rect 50 2975 75 3000
rect 2340 2930 2365 2955
rect 3085 2955 3105 2975
rect 3140 2955 3160 2975
rect 3270 2955 3290 2975
rect 3450 2955 3470 2975
rect 3630 2955 3650 2975
rect 3810 2955 3830 2975
rect 3990 2955 4010 2975
rect 4170 2955 4190 2975
rect 4350 2955 4370 2975
rect 4530 2955 4550 2975
rect 4710 2955 4730 2975
rect 4840 2955 4860 2975
rect 4890 2955 4910 2975
rect 2340 2870 2365 2895
rect 50 2825 75 2850
rect 585 2825 610 2850
rect 1255 2810 1280 2835
rect 1970 2810 1995 2835
rect 50 2765 75 2790
rect 585 2765 610 2790
rect 3000 2785 3020 2805
rect 3180 2785 3200 2805
rect 3360 2785 3380 2805
rect 3540 2785 3560 2805
rect 3720 2785 3740 2805
rect 3900 2785 3920 2805
rect 4080 2785 4100 2805
rect 4260 2785 4280 2805
rect 4440 2785 4460 2805
rect 4620 2785 4640 2805
rect 4800 2785 4820 2805
rect 4980 2785 5000 2805
rect 3000 2725 3020 2745
rect 3180 2725 3200 2745
rect 3360 2725 3380 2745
rect 3540 2725 3560 2745
rect 3720 2725 3740 2745
rect 3900 2725 3920 2745
rect 4080 2725 4100 2745
rect 4260 2725 4280 2745
rect 4440 2725 4460 2745
rect 4620 2725 4640 2745
rect 4800 2725 4820 2745
rect 4980 2725 5000 2745
rect 2910 2355 2930 2375
rect 3000 2350 3020 2370
rect 3090 2355 3110 2375
rect 3450 2355 3470 2375
rect 3810 2355 3830 2375
rect 3895 2355 3915 2375
rect 3990 2355 4010 2375
rect 4160 2355 4180 2375
rect 4530 2355 4550 2375
rect 4890 2355 4910 2375
rect 5070 2355 5090 2375
rect 3270 2310 3290 2330
rect 3630 2310 3650 2330
rect 4350 2310 4370 2330
rect 4710 2310 4730 2330
rect 3450 2265 3470 2285
rect 4530 2265 4550 2285
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 4145 2070 4165 2090
rect 4265 2070 4285 2090
rect 4385 2070 4405 2090
rect 4505 2070 4525 2090
rect 4625 2070 4645 2090
rect 4745 2070 4765 2090
rect 4865 2070 4885 2090
rect 4985 2070 5005 2090
rect 5105 2070 5125 2090
rect 2630 2025 2650 2045
rect 2815 2025 2835 2045
rect -35 1695 -15 1715
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4085 2025 4105 2045
rect 4445 2025 4465 2045
rect 4805 2025 4825 2045
rect 5165 2025 5185 2045
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 3865 1855 3885 1875
rect 4115 1855 4135 1875
rect 4205 1855 4225 1875
rect 4325 1855 4345 1875
rect 4445 1855 4465 1875
rect 4565 1855 4585 1875
rect 4685 1855 4705 1875
rect 4805 1855 4825 1875
rect 4925 1855 4945 1875
rect 5045 1855 5065 1875
rect 5135 1855 5155 1875
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4205 1795 4225 1815
rect 4565 1795 4585 1815
rect 4925 1795 4945 1815
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4205 1735 4225 1755
rect 4445 1735 4465 1755
rect 4685 1735 4705 1755
rect 4745 1735 4765 1755
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4325 1690 4345 1710
rect 4565 1690 4585 1710
rect 4805 1690 4825 1710
rect 3175 1570 3195 1590
rect 4805 1570 4825 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4265 1520 4285 1540
rect 4385 1520 4405 1540
rect 4505 1520 4525 1540
rect 4625 1520 4645 1540
rect 4745 1520 4765 1540
rect 2845 1465 2865 1485
rect 3925 1465 3945 1485
rect 4055 1465 4075 1485
rect 5135 1465 5155 1485
rect 3385 1165 3405 1185
rect 4595 1165 4615 1185
rect 2950 1105 2970 1125
rect 3030 1105 3050 1125
rect 3110 1105 3130 1125
rect 3190 1105 3210 1125
rect 3270 1105 3290 1125
rect 3350 1105 3370 1125
rect 3430 1105 3450 1125
rect 3510 1105 3530 1125
rect 3590 1105 3610 1125
rect 3670 1105 3690 1125
rect 3750 1105 3770 1125
rect 3830 1105 3850 1125
rect 3910 1105 3930 1125
rect 3990 1105 4010 1125
rect 4070 1105 4090 1125
rect 4150 1105 4170 1125
rect 4230 1105 4250 1125
rect 4310 1105 4330 1125
rect 4390 1105 4410 1125
rect 4470 1105 4490 1125
rect 4550 1105 4570 1125
rect 4630 1105 4650 1125
rect 4710 1105 4730 1125
rect 4790 1105 4810 1125
rect 4870 1105 4890 1125
rect 4950 1105 4970 1125
rect 2910 1020 2930 1040
rect 5065 1020 5085 1040
rect 3000 910 3020 930
rect 3180 910 3200 930
rect 3360 910 3380 930
rect 3540 910 3560 930
rect 3720 910 3740 930
rect 3900 910 3920 930
rect 4080 910 4100 930
rect 4260 910 4280 930
rect 4440 910 4460 930
rect 4620 910 4640 930
rect 4800 910 4820 930
rect 4980 910 5000 930
rect 3090 725 3110 745
rect 3270 740 3290 760
rect 3450 740 3470 760
rect 3630 740 3650 760
rect 3810 740 3830 760
rect 3990 740 4010 760
rect 4170 740 4190 760
rect 4350 740 4370 760
rect 4530 740 4550 760
rect 4710 740 4730 760
rect 4890 740 4910 760
<< metal1 >>
rect 1245 3525 1285 3530
rect 1245 3495 1250 3525
rect 1280 3495 1285 3525
rect 1245 3490 1285 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1190 3340 1230 3345
rect 1190 3310 1195 3340
rect 1225 3310 1230 3340
rect 1190 3305 1230 3310
rect 1145 3285 1185 3290
rect 1145 3255 1150 3285
rect 1180 3255 1185 3285
rect 1145 3250 1185 3255
rect 40 3170 45 3205
rect 80 3170 85 3205
rect 40 3110 45 3145
rect 80 3110 85 3145
rect 1155 3105 1175 3250
rect 1145 3100 1185 3105
rect 1145 3070 1150 3100
rect 1180 3070 1185 3100
rect 1145 3065 1185 3070
rect 40 3030 45 3065
rect 80 3030 85 3065
rect 40 2970 45 3005
rect 80 2970 85 3005
rect 1200 2855 1220 3305
rect 1255 3200 1275 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1245 3165 1250 3200
rect 1285 3165 1290 3200
rect 1255 3140 1275 3165
rect 1245 3105 1250 3140
rect 1285 3105 1290 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 40 2820 45 2855
rect 80 2820 85 2855
rect 575 2820 580 2855
rect 615 2820 620 2855
rect 1190 2850 1230 2855
rect 1190 2820 1195 2850
rect 1225 2820 1230 2850
rect 2340 2840 2360 2860
rect 1190 2815 1230 2820
rect 1245 2805 1250 2840
rect 1285 2805 1290 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 40 2760 45 2795
rect 80 2760 85 2795
rect 575 2760 580 2795
rect 615 2760 620 2795
rect 1255 2750 1275 2805
rect 2330 2800 2370 2805
rect 1245 2745 1285 2750
rect 1245 2715 1250 2745
rect 1280 2715 1285 2745
rect 1245 2710 1285 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 955 1710 1305 1870
rect 955 1680 1270 1710
rect 1300 1680 1305 1710
rect 955 1520 1305 1680
rect 1635 1190 1985 2200
rect 2160 1715 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2150 1710 2190 1715
rect 2150 1680 2155 1710
rect 2185 1680 2190 1710
rect 2150 1675 2190 1680
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3130 3340 3170 3345
rect 3130 3310 3135 3340
rect 3165 3310 3170 3340
rect 3130 3305 3170 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 1035 2175 1190
rect 2435 1035 2455 1725
rect 275 1030 2215 1035
rect 275 1000 2180 1030
rect 2210 1000 2215 1030
rect 275 995 2215 1000
rect 2425 1030 2465 1035
rect 2425 1000 2430 1030
rect 2460 1000 2465 1030
rect 2425 995 2465 1000
rect 275 840 2175 995
rect 2530 755 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3140 3145 3160 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5340 3335 5380 3340
rect 5340 3305 5345 3335
rect 5375 3305 5380 3335
rect 5340 3300 5380 3305
rect 4880 3285 4920 3290
rect 4880 3255 4885 3285
rect 4915 3255 4920 3285
rect 4880 3250 4920 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3130 3140 3170 3145
rect 3130 3110 3135 3140
rect 3165 3110 3170 3140
rect 3130 3105 3170 3110
rect 4830 3140 4870 3145
rect 4830 3110 4835 3140
rect 4865 3110 4870 3140
rect 4830 3105 4870 3110
rect 3140 2985 3160 3105
rect 3980 3080 4020 3085
rect 3980 3050 3985 3080
rect 4015 3050 4020 3080
rect 3980 3045 4020 3050
rect 3440 3035 3480 3040
rect 3440 3005 3445 3035
rect 3475 3005 3480 3035
rect 3440 3000 3480 3005
rect 3800 3035 3840 3040
rect 3800 3005 3805 3035
rect 3835 3005 3840 3035
rect 3800 3000 3840 3005
rect 3450 2985 3470 3000
rect 3810 2985 3830 3000
rect 3990 2985 4010 3045
rect 4340 3035 4380 3040
rect 4340 3005 4345 3035
rect 4375 3005 4380 3035
rect 4340 3000 4380 3005
rect 4700 3035 4740 3040
rect 4700 3005 4705 3035
rect 4735 3005 4740 3035
rect 4700 3000 4740 3005
rect 4350 2985 4370 3000
rect 4710 2985 4730 3000
rect 4840 2985 4860 3105
rect 4890 2985 4910 3250
rect 5295 3140 5335 3145
rect 5295 3110 5300 3140
rect 5330 3110 5335 3140
rect 5295 3105 5335 3110
rect 3075 2980 3115 2985
rect 3075 2950 3080 2980
rect 3110 2950 3115 2980
rect 3075 2945 3115 2950
rect 3135 2975 3170 2985
rect 3135 2955 3140 2975
rect 3160 2955 3170 2975
rect 3135 2945 3170 2955
rect 3260 2980 3300 2985
rect 3260 2950 3265 2980
rect 3295 2950 3300 2980
rect 3260 2945 3300 2950
rect 3440 2975 3480 2985
rect 3440 2955 3450 2975
rect 3470 2955 3480 2975
rect 3440 2945 3480 2955
rect 3620 2980 3660 2985
rect 3620 2950 3625 2980
rect 3655 2950 3660 2980
rect 3620 2945 3660 2950
rect 3800 2975 3840 2985
rect 3800 2955 3810 2975
rect 3830 2955 3840 2975
rect 3800 2945 3840 2955
rect 3980 2975 4020 2985
rect 3980 2955 3990 2975
rect 4010 2955 4020 2975
rect 3980 2945 4020 2955
rect 4160 2980 4200 2985
rect 4160 2950 4165 2980
rect 4195 2950 4200 2980
rect 4160 2945 4200 2950
rect 4340 2975 4380 2985
rect 4340 2955 4350 2975
rect 4370 2955 4380 2975
rect 4340 2945 4380 2955
rect 4520 2980 4560 2985
rect 4520 2950 4525 2980
rect 4555 2950 4560 2980
rect 4520 2945 4560 2950
rect 4700 2975 4740 2985
rect 4700 2955 4710 2975
rect 4730 2955 4740 2975
rect 4700 2945 4740 2955
rect 4830 2975 4865 2985
rect 4830 2955 4840 2975
rect 4860 2955 4865 2975
rect 4830 2945 4865 2955
rect 4885 2975 4920 2985
rect 4885 2955 4890 2975
rect 4910 2955 4920 2975
rect 4885 2945 4920 2955
rect 2990 2810 3030 2815
rect 2990 2780 2995 2810
rect 3025 2780 3030 2810
rect 2990 2775 3030 2780
rect 3170 2810 3210 2815
rect 3170 2780 3175 2810
rect 3205 2780 3210 2810
rect 3170 2775 3210 2780
rect 3350 2810 3390 2815
rect 3350 2780 3355 2810
rect 3385 2780 3390 2810
rect 3350 2775 3390 2780
rect 3530 2810 3570 2815
rect 3530 2780 3535 2810
rect 3565 2780 3570 2810
rect 3530 2775 3570 2780
rect 3710 2810 3750 2815
rect 3710 2780 3715 2810
rect 3745 2780 3750 2810
rect 3710 2775 3750 2780
rect 3890 2810 3930 2815
rect 3890 2780 3895 2810
rect 3925 2780 3930 2810
rect 3890 2775 3930 2780
rect 4070 2810 4110 2815
rect 4070 2780 4075 2810
rect 4105 2780 4110 2810
rect 4070 2775 4110 2780
rect 4250 2810 4290 2815
rect 4250 2780 4255 2810
rect 4285 2780 4290 2810
rect 4250 2775 4290 2780
rect 4430 2810 4470 2815
rect 4430 2780 4435 2810
rect 4465 2780 4470 2810
rect 4430 2775 4470 2780
rect 4610 2810 4650 2815
rect 4610 2780 4615 2810
rect 4645 2780 4650 2810
rect 4610 2775 4650 2780
rect 4790 2810 4830 2815
rect 4790 2780 4795 2810
rect 4825 2780 4830 2810
rect 4790 2775 4830 2780
rect 4970 2810 5010 2815
rect 4970 2780 4975 2810
rect 5005 2780 5010 2810
rect 4970 2775 5010 2780
rect 4980 2755 5000 2775
rect 2990 2750 3030 2755
rect 2990 2720 2995 2750
rect 3025 2720 3030 2750
rect 2990 2715 3030 2720
rect 3170 2750 3210 2755
rect 3170 2720 3175 2750
rect 3205 2720 3210 2750
rect 3170 2715 3210 2720
rect 3350 2750 3390 2755
rect 3350 2720 3355 2750
rect 3385 2720 3390 2750
rect 3350 2715 3390 2720
rect 3530 2750 3570 2755
rect 3530 2720 3535 2750
rect 3565 2720 3570 2750
rect 3530 2715 3570 2720
rect 3710 2750 3750 2755
rect 3710 2720 3715 2750
rect 3745 2720 3750 2750
rect 3710 2715 3750 2720
rect 3890 2750 3930 2755
rect 3890 2720 3895 2750
rect 3925 2720 3930 2750
rect 3890 2715 3930 2720
rect 4070 2750 4110 2755
rect 4070 2720 4075 2750
rect 4105 2720 4110 2750
rect 4070 2715 4110 2720
rect 4250 2750 4290 2755
rect 4250 2720 4255 2750
rect 4285 2720 4290 2750
rect 4250 2715 4290 2720
rect 4430 2750 4470 2755
rect 4430 2720 4435 2750
rect 4465 2720 4470 2750
rect 4430 2715 4470 2720
rect 4610 2750 4650 2755
rect 4610 2720 4615 2750
rect 4645 2720 4650 2750
rect 4610 2715 4650 2720
rect 4790 2750 4830 2755
rect 4790 2720 4795 2750
rect 4825 2720 4830 2750
rect 4790 2715 4830 2720
rect 4970 2750 5010 2755
rect 4970 2720 4975 2750
rect 5005 2720 5010 2750
rect 4970 2715 5010 2720
rect 2900 2375 2940 2385
rect 3080 2380 3120 2385
rect 2900 2355 2910 2375
rect 2930 2355 2940 2375
rect 2900 2345 2940 2355
rect 2990 2375 3030 2380
rect 2990 2345 2995 2375
rect 3025 2345 3030 2375
rect 3080 2350 3085 2380
rect 3115 2350 3120 2380
rect 3080 2345 3120 2350
rect 3440 2375 3480 2385
rect 3440 2355 3450 2375
rect 3470 2355 3480 2375
rect 3440 2345 3480 2355
rect 3800 2380 3840 2385
rect 3800 2350 3805 2380
rect 3835 2350 3840 2380
rect 3800 2345 3840 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3980 2375 4020 2385
rect 3980 2355 3990 2375
rect 4010 2355 4020 2375
rect 3980 2345 4020 2355
rect 4150 2380 4190 2385
rect 4150 2350 4155 2380
rect 4185 2350 4190 2380
rect 4150 2345 4190 2350
rect 4520 2375 4560 2385
rect 4520 2355 4530 2375
rect 4550 2355 4560 2375
rect 4520 2345 4560 2355
rect 4880 2380 4920 2385
rect 4880 2350 4885 2380
rect 4915 2350 4920 2380
rect 4880 2345 4920 2350
rect 5060 2375 5100 2385
rect 5060 2355 5070 2375
rect 5090 2355 5100 2375
rect 5060 2345 5100 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 2910 2205 2930 2345
rect 2990 2340 3030 2345
rect 3090 2250 3110 2345
rect 3260 2335 3300 2340
rect 3260 2305 3265 2335
rect 3295 2305 3300 2335
rect 3260 2300 3300 2305
rect 3080 2245 3120 2250
rect 3080 2215 3085 2245
rect 3115 2215 3120 2245
rect 3080 2210 3120 2215
rect 2900 2200 2940 2205
rect 2900 2170 2905 2200
rect 2935 2170 2940 2200
rect 2900 2165 2940 2170
rect 3270 2155 3290 2300
rect 3450 2295 3470 2345
rect 3620 2335 3660 2340
rect 3620 2305 3625 2335
rect 3655 2305 3660 2335
rect 3620 2300 3660 2305
rect 3440 2290 3480 2295
rect 3440 2260 3445 2290
rect 3475 2260 3480 2290
rect 3440 2255 3480 2260
rect 3260 2150 3300 2155
rect 3260 2120 3265 2150
rect 3295 2120 3300 2150
rect 3260 2115 3300 2120
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3990 2205 4010 2345
rect 4340 2335 4380 2340
rect 4340 2305 4345 2335
rect 4375 2305 4380 2335
rect 4340 2300 4380 2305
rect 4530 2295 4550 2345
rect 4700 2335 4740 2340
rect 4700 2305 4705 2335
rect 4735 2305 4740 2335
rect 4700 2300 4740 2305
rect 4520 2290 4560 2295
rect 4520 2260 4525 2290
rect 4555 2260 4560 2290
rect 4520 2255 4560 2260
rect 5070 2205 5090 2345
rect 5250 2290 5290 2295
rect 5250 2260 5255 2290
rect 5285 2260 5290 2290
rect 5250 2255 5290 2260
rect 3980 2200 4020 2205
rect 3980 2170 3985 2200
rect 4015 2170 4020 2200
rect 3980 2165 4020 2170
rect 5060 2200 5100 2205
rect 5060 2170 5065 2200
rect 5095 2170 5100 2200
rect 5060 2165 5100 2170
rect 4075 2145 4115 2150
rect 4075 2115 4080 2145
rect 4110 2115 4115 2145
rect 4075 2110 4115 2115
rect 4085 2055 4105 2110
rect 4135 2095 4175 2100
rect 4135 2065 4140 2095
rect 4170 2065 4175 2095
rect 4135 2060 4175 2065
rect 4255 2095 4295 2100
rect 4255 2065 4260 2095
rect 4290 2065 4295 2095
rect 4255 2060 4295 2065
rect 4375 2095 4415 2100
rect 4375 2065 4380 2095
rect 4410 2065 4415 2095
rect 4375 2060 4415 2065
rect 4495 2095 4535 2100
rect 4495 2065 4500 2095
rect 4530 2065 4535 2095
rect 4495 2060 4535 2065
rect 4615 2095 4655 2100
rect 4615 2065 4620 2095
rect 4650 2065 4655 2095
rect 4615 2060 4655 2065
rect 4735 2095 4775 2100
rect 4735 2065 4740 2095
rect 4770 2065 4775 2095
rect 4735 2060 4775 2065
rect 4855 2095 4895 2100
rect 4855 2065 4860 2095
rect 4890 2065 4895 2095
rect 4855 2060 4895 2065
rect 4975 2095 5015 2100
rect 4975 2065 4980 2095
rect 5010 2065 5015 2095
rect 4975 2060 5015 2065
rect 5095 2095 5135 2100
rect 5095 2065 5100 2095
rect 5130 2065 5135 2095
rect 5095 2060 5135 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3945 2055
rect 3885 2020 3890 2050
rect 3920 2020 3945 2050
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2675 1725 2715 1730
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1050 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1495 2865 1510
rect 3925 1495 3945 2015
rect 4055 2050 4115 2055
rect 4055 2020 4080 2050
rect 4110 2020 4115 2050
rect 4055 2015 4115 2020
rect 4435 2050 4475 2055
rect 4435 2020 4440 2050
rect 4470 2020 4475 2050
rect 4435 2015 4475 2020
rect 4795 2050 4835 2055
rect 4795 2020 4800 2050
rect 4830 2020 4835 2050
rect 4795 2015 4835 2020
rect 5155 2050 5195 2055
rect 5155 2020 5160 2050
rect 5190 2020 5195 2050
rect 5155 2015 5195 2020
rect 4055 1495 4075 2015
rect 4105 1875 4145 1885
rect 4105 1855 4115 1875
rect 4135 1855 4145 1875
rect 4105 1845 4145 1855
rect 4195 1875 4235 1885
rect 4195 1855 4205 1875
rect 4225 1855 4235 1875
rect 4195 1845 4235 1855
rect 4315 1880 4355 1885
rect 4315 1850 4320 1880
rect 4350 1850 4355 1880
rect 4315 1845 4355 1850
rect 4435 1875 4475 1885
rect 4435 1855 4445 1875
rect 4465 1855 4475 1875
rect 4435 1845 4475 1855
rect 4555 1875 4595 1885
rect 4555 1855 4565 1875
rect 4585 1855 4595 1875
rect 4555 1845 4595 1855
rect 4675 1880 4715 1885
rect 4675 1850 4680 1880
rect 4710 1850 4715 1880
rect 4675 1845 4715 1850
rect 4795 1875 4835 1885
rect 4795 1855 4805 1875
rect 4825 1855 4835 1875
rect 4795 1845 4835 1855
rect 4915 1875 4955 1885
rect 4915 1855 4925 1875
rect 4945 1855 4955 1875
rect 4915 1845 4955 1855
rect 5035 1880 5075 1885
rect 5035 1850 5040 1880
rect 5070 1850 5075 1880
rect 5035 1845 5075 1850
rect 5125 1875 5165 1885
rect 5125 1855 5135 1875
rect 5155 1855 5165 1875
rect 5125 1845 5165 1855
rect 4115 1825 4135 1845
rect 4205 1825 4225 1845
rect 4445 1825 4465 1845
rect 4565 1825 4585 1845
rect 4105 1820 4145 1825
rect 4105 1790 4110 1820
rect 4140 1790 4145 1820
rect 4105 1785 4145 1790
rect 4195 1820 4235 1825
rect 4195 1790 4200 1820
rect 4230 1790 4235 1820
rect 4195 1785 4235 1790
rect 4435 1820 4475 1825
rect 4435 1790 4440 1820
rect 4470 1790 4475 1820
rect 4435 1785 4475 1790
rect 4555 1820 4595 1825
rect 4555 1790 4560 1820
rect 4590 1790 4595 1820
rect 4555 1785 4595 1790
rect 4195 1760 4235 1765
rect 4195 1730 4200 1760
rect 4230 1730 4235 1760
rect 4195 1725 4235 1730
rect 4435 1760 4475 1765
rect 4435 1730 4440 1760
rect 4470 1730 4475 1760
rect 4435 1725 4475 1730
rect 4565 1720 4585 1785
rect 4685 1765 4705 1845
rect 4805 1825 4825 1845
rect 4925 1825 4945 1845
rect 5135 1825 5155 1845
rect 4795 1820 4835 1825
rect 4795 1790 4800 1820
rect 4830 1790 4835 1820
rect 4795 1785 4835 1790
rect 4915 1820 4955 1825
rect 4915 1790 4920 1820
rect 4950 1790 4955 1820
rect 4915 1785 4955 1790
rect 5125 1820 5165 1825
rect 5125 1790 5130 1820
rect 5160 1790 5165 1820
rect 5125 1785 5165 1790
rect 5260 1765 5280 2255
rect 5305 2150 5325 3105
rect 5295 2145 5335 2150
rect 5295 2115 5300 2145
rect 5330 2115 5335 2145
rect 5295 2110 5335 2115
rect 5350 1825 5370 3300
rect 5390 3285 5430 3290
rect 5390 3255 5395 3285
rect 5425 3255 5430 3285
rect 5390 3250 5430 3255
rect 5340 1820 5380 1825
rect 5340 1790 5345 1820
rect 5375 1790 5380 1820
rect 5340 1785 5380 1790
rect 4675 1760 4715 1765
rect 4675 1730 4680 1760
rect 4710 1730 4715 1760
rect 4675 1725 4715 1730
rect 4735 1760 4775 1765
rect 4735 1730 4740 1760
rect 4770 1730 4775 1760
rect 4735 1725 4775 1730
rect 5250 1760 5290 1765
rect 5250 1730 5255 1760
rect 5285 1730 5290 1760
rect 5250 1725 5290 1730
rect 4315 1715 4355 1720
rect 4315 1685 4320 1715
rect 4350 1685 4355 1715
rect 4315 1680 4355 1685
rect 4555 1715 4595 1720
rect 4555 1685 4560 1715
rect 4590 1685 4595 1715
rect 4555 1680 4595 1685
rect 4795 1715 4835 1720
rect 4795 1685 4800 1715
rect 4830 1685 4835 1715
rect 4795 1680 4835 1685
rect 5400 1600 5420 3250
rect 4795 1595 4835 1600
rect 4795 1565 4800 1595
rect 4830 1565 4835 1595
rect 4795 1560 4835 1565
rect 5390 1595 5430 1600
rect 5390 1565 5395 1595
rect 5425 1565 5430 1595
rect 5390 1560 5430 1565
rect 4255 1545 4295 1550
rect 4255 1515 4260 1545
rect 4290 1515 4295 1545
rect 4255 1510 4295 1515
rect 4375 1545 4415 1550
rect 4375 1515 4380 1545
rect 4410 1515 4415 1545
rect 4375 1510 4415 1515
rect 4495 1545 4535 1550
rect 4495 1515 4500 1545
rect 4530 1515 4535 1545
rect 4495 1510 4535 1515
rect 4615 1545 4655 1550
rect 4615 1515 4620 1545
rect 4650 1515 4655 1545
rect 4615 1510 4655 1515
rect 4735 1545 4775 1550
rect 4735 1515 4740 1545
rect 4770 1515 4775 1545
rect 4735 1510 4775 1515
rect 5125 1545 5165 1550
rect 5125 1515 5130 1545
rect 5160 1515 5165 1545
rect 5125 1510 5165 1515
rect 5135 1495 5155 1510
rect 2835 1485 2875 1495
rect 2835 1465 2845 1485
rect 2865 1465 2875 1485
rect 2835 1455 2875 1465
rect 3915 1485 3955 1495
rect 3915 1465 3925 1485
rect 3945 1465 3955 1485
rect 3915 1455 3955 1465
rect 4045 1485 4085 1495
rect 4045 1465 4055 1485
rect 4075 1465 4085 1485
rect 4045 1455 4085 1465
rect 5125 1485 5165 1495
rect 5125 1465 5135 1485
rect 5155 1465 5165 1485
rect 5125 1455 5165 1465
rect 3375 1190 3415 1195
rect 3375 1160 3380 1190
rect 3410 1160 3415 1190
rect 3375 1155 3415 1160
rect 4585 1190 4625 1195
rect 4585 1160 4590 1190
rect 4620 1160 4625 1190
rect 4585 1155 4625 1160
rect 2940 1130 2980 1135
rect 2940 1100 2945 1130
rect 2975 1100 2980 1130
rect 2940 1095 2980 1100
rect 3020 1130 3060 1135
rect 3020 1100 3025 1130
rect 3055 1100 3060 1130
rect 3020 1095 3060 1100
rect 3100 1130 3140 1135
rect 3100 1100 3105 1130
rect 3135 1100 3140 1130
rect 3100 1095 3140 1100
rect 3180 1130 3220 1135
rect 3180 1100 3185 1130
rect 3215 1100 3220 1130
rect 3180 1095 3220 1100
rect 3260 1130 3300 1135
rect 3260 1100 3265 1130
rect 3295 1100 3300 1130
rect 3260 1095 3300 1100
rect 3340 1130 3380 1135
rect 3340 1100 3345 1130
rect 3375 1100 3380 1130
rect 3340 1095 3380 1100
rect 3420 1130 3460 1135
rect 3420 1100 3425 1130
rect 3455 1100 3460 1130
rect 3420 1095 3460 1100
rect 3500 1130 3540 1135
rect 3500 1100 3505 1130
rect 3535 1100 3540 1130
rect 3500 1095 3540 1100
rect 3580 1130 3620 1135
rect 3580 1100 3585 1130
rect 3615 1100 3620 1130
rect 3580 1095 3620 1100
rect 3660 1130 3700 1135
rect 3660 1100 3665 1130
rect 3695 1100 3700 1130
rect 3660 1095 3700 1100
rect 3740 1130 3780 1135
rect 3740 1100 3745 1130
rect 3775 1100 3780 1130
rect 3740 1095 3780 1100
rect 3820 1130 3860 1135
rect 3820 1100 3825 1130
rect 3855 1100 3860 1130
rect 3820 1095 3860 1100
rect 3900 1130 3940 1135
rect 3900 1100 3905 1130
rect 3935 1100 3940 1130
rect 3900 1095 3940 1100
rect 3980 1130 4020 1135
rect 3980 1100 3985 1130
rect 4015 1100 4020 1130
rect 3980 1095 4020 1100
rect 4060 1130 4100 1135
rect 4060 1100 4065 1130
rect 4095 1100 4100 1130
rect 4060 1095 4100 1100
rect 4140 1130 4180 1135
rect 4140 1100 4145 1130
rect 4175 1100 4180 1130
rect 4140 1095 4180 1100
rect 4220 1130 4260 1135
rect 4220 1100 4225 1130
rect 4255 1100 4260 1130
rect 4220 1095 4260 1100
rect 4300 1130 4340 1135
rect 4300 1100 4305 1130
rect 4335 1100 4340 1130
rect 4300 1095 4340 1100
rect 4380 1130 4420 1135
rect 4380 1100 4385 1130
rect 4415 1100 4420 1130
rect 4380 1095 4420 1100
rect 4460 1130 4500 1135
rect 4460 1100 4465 1130
rect 4495 1100 4500 1130
rect 4460 1095 4500 1100
rect 4540 1130 4580 1135
rect 4540 1100 4545 1130
rect 4575 1100 4580 1130
rect 4540 1095 4580 1100
rect 4620 1130 4660 1135
rect 4620 1100 4625 1130
rect 4655 1100 4660 1130
rect 4620 1095 4660 1100
rect 4700 1130 4740 1135
rect 4700 1100 4705 1130
rect 4735 1100 4740 1130
rect 4700 1095 4740 1100
rect 4780 1130 4820 1135
rect 4780 1100 4785 1130
rect 4815 1100 4820 1130
rect 4780 1095 4820 1100
rect 4860 1130 4900 1135
rect 4860 1100 4865 1130
rect 4895 1100 4900 1130
rect 4860 1095 4900 1100
rect 4940 1130 4980 1135
rect 4940 1100 4945 1130
rect 4975 1100 4980 1130
rect 4940 1095 4980 1100
rect 2620 1045 2660 1050
rect 2620 1015 2625 1045
rect 2655 1015 2660 1045
rect 2620 1010 2660 1015
rect 2900 1045 2940 1050
rect 2900 1015 2905 1045
rect 2935 1015 2940 1045
rect 2900 1010 2940 1015
rect 5055 1045 5095 1050
rect 5055 1015 5060 1045
rect 5090 1015 5095 1045
rect 5055 1010 5095 1015
rect 2990 935 3030 940
rect 2990 905 2995 935
rect 3025 905 3030 935
rect 2990 900 3030 905
rect 3170 935 3210 940
rect 3170 905 3175 935
rect 3205 905 3210 935
rect 3170 900 3210 905
rect 3350 935 3390 940
rect 3350 905 3355 935
rect 3385 905 3390 935
rect 3350 900 3390 905
rect 3530 935 3570 940
rect 3530 905 3535 935
rect 3565 905 3570 935
rect 3530 900 3570 905
rect 3710 935 3750 940
rect 3710 905 3715 935
rect 3745 905 3750 935
rect 3710 900 3750 905
rect 3890 935 3930 940
rect 3890 905 3895 935
rect 3925 905 3930 935
rect 3890 900 3930 905
rect 4070 935 4110 940
rect 4070 905 4075 935
rect 4105 905 4110 935
rect 4070 900 4110 905
rect 4250 935 4290 940
rect 4250 905 4255 935
rect 4285 905 4290 935
rect 4250 900 4290 905
rect 4430 935 4470 940
rect 4430 905 4435 935
rect 4465 905 4470 935
rect 4430 900 4470 905
rect 4610 935 4650 940
rect 4610 905 4615 935
rect 4645 905 4650 935
rect 4610 900 4650 905
rect 4790 935 4830 940
rect 4790 905 4795 935
rect 4825 905 4830 935
rect 4790 900 4830 905
rect 4970 935 5010 940
rect 4970 905 4975 935
rect 5005 905 5010 935
rect 4970 900 5010 905
rect 3260 760 3300 770
rect 2520 750 2560 755
rect 2520 720 2525 750
rect 2555 720 2560 750
rect 2520 715 2560 720
rect 3080 750 3120 755
rect 3080 720 3085 750
rect 3115 720 3120 750
rect 3260 740 3270 760
rect 3290 740 3300 760
rect 3260 730 3300 740
rect 3440 760 3480 770
rect 3440 740 3450 760
rect 3470 740 3480 760
rect 3440 730 3480 740
rect 3620 765 3660 770
rect 3620 735 3625 765
rect 3655 735 3660 765
rect 3620 730 3660 735
rect 3800 760 3840 770
rect 3800 740 3810 760
rect 3830 740 3840 760
rect 3800 730 3840 740
rect 3980 765 4020 770
rect 3980 735 3985 765
rect 4015 735 4020 765
rect 3980 730 4020 735
rect 4160 760 4200 770
rect 4160 740 4170 760
rect 4190 740 4200 760
rect 4160 730 4200 740
rect 4340 765 4380 770
rect 4340 735 4345 765
rect 4375 735 4380 765
rect 4340 730 4380 735
rect 4520 765 4560 770
rect 4520 735 4525 765
rect 4555 735 4560 765
rect 4520 730 4560 735
rect 4700 765 4740 770
rect 4700 735 4705 765
rect 4735 735 4740 765
rect 4700 730 4740 735
rect 4880 765 4920 770
rect 4880 735 4885 765
rect 4915 735 4920 765
rect 4880 730 4920 735
rect 3080 715 3120 720
rect 3270 295 3290 730
rect 3450 715 3470 730
rect 3810 715 3830 730
rect 3440 710 3480 715
rect 3440 680 3445 710
rect 3475 680 3480 710
rect 3440 675 3480 680
rect 3800 710 3840 715
rect 3800 680 3805 710
rect 3835 680 3840 710
rect 3800 675 3840 680
rect 3810 295 3830 675
rect 3990 295 4010 730
rect 4170 715 4190 730
rect 4160 710 4200 715
rect 4160 680 4165 710
rect 4195 680 4200 710
rect 4160 675 4200 680
rect 4710 295 4730 730
<< via1 >>
rect 1250 3495 1280 3525
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1195 3310 1225 3340
rect 1150 3255 1180 3285
rect 45 3200 80 3205
rect 45 3175 50 3200
rect 50 3175 75 3200
rect 75 3175 80 3200
rect 45 3170 80 3175
rect 45 3140 80 3145
rect 45 3115 50 3140
rect 50 3115 75 3140
rect 75 3115 80 3140
rect 45 3110 80 3115
rect 1150 3070 1180 3100
rect 45 3060 80 3065
rect 45 3035 50 3060
rect 50 3035 75 3060
rect 75 3035 80 3060
rect 45 3030 80 3035
rect 45 3000 80 3005
rect 45 2975 50 3000
rect 50 2975 75 3000
rect 75 2975 80 3000
rect 45 2970 80 2975
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1250 3195 1285 3200
rect 1250 3170 1255 3195
rect 1255 3170 1280 3195
rect 1280 3170 1285 3195
rect 1250 3165 1285 3170
rect 1250 3135 1285 3140
rect 1250 3110 1255 3135
rect 1255 3110 1280 3135
rect 1280 3110 1285 3135
rect 1250 3105 1285 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 45 2850 80 2855
rect 45 2825 50 2850
rect 50 2825 75 2850
rect 75 2825 80 2850
rect 45 2820 80 2825
rect 580 2850 615 2855
rect 580 2825 585 2850
rect 585 2825 610 2850
rect 610 2825 615 2850
rect 580 2820 615 2825
rect 1195 2820 1225 2850
rect 1250 2835 1285 2840
rect 1250 2810 1255 2835
rect 1255 2810 1280 2835
rect 1280 2810 1285 2835
rect 1250 2805 1285 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 45 2790 80 2795
rect 45 2765 50 2790
rect 50 2765 75 2790
rect 75 2765 80 2790
rect 45 2760 80 2765
rect 580 2790 615 2795
rect 580 2765 585 2790
rect 585 2765 610 2790
rect 610 2765 615 2790
rect 580 2760 615 2765
rect 1250 2715 1280 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1300 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2155 1680 2185 1710
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3135 3310 3165 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2180 1000 2210 1030
rect 2430 1000 2460 1030
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5345 3305 5375 3335
rect 4885 3255 4915 3285
rect 4445 3155 4475 3185
rect 3135 3110 3165 3140
rect 4835 3110 4865 3140
rect 3985 3050 4015 3080
rect 3445 3005 3475 3035
rect 3805 3005 3835 3035
rect 4345 3005 4375 3035
rect 4705 3005 4735 3035
rect 5300 3110 5330 3140
rect 3080 2975 3110 2980
rect 3080 2955 3085 2975
rect 3085 2955 3105 2975
rect 3105 2955 3110 2975
rect 3080 2950 3110 2955
rect 3265 2975 3295 2980
rect 3265 2955 3270 2975
rect 3270 2955 3290 2975
rect 3290 2955 3295 2975
rect 3265 2950 3295 2955
rect 3625 2975 3655 2980
rect 3625 2955 3630 2975
rect 3630 2955 3650 2975
rect 3650 2955 3655 2975
rect 3625 2950 3655 2955
rect 4165 2975 4195 2980
rect 4165 2955 4170 2975
rect 4170 2955 4190 2975
rect 4190 2955 4195 2975
rect 4165 2950 4195 2955
rect 4525 2975 4555 2980
rect 4525 2955 4530 2975
rect 4530 2955 4550 2975
rect 4550 2955 4555 2975
rect 4525 2950 4555 2955
rect 2995 2805 3025 2810
rect 2995 2785 3000 2805
rect 3000 2785 3020 2805
rect 3020 2785 3025 2805
rect 2995 2780 3025 2785
rect 3175 2805 3205 2810
rect 3175 2785 3180 2805
rect 3180 2785 3200 2805
rect 3200 2785 3205 2805
rect 3175 2780 3205 2785
rect 3355 2805 3385 2810
rect 3355 2785 3360 2805
rect 3360 2785 3380 2805
rect 3380 2785 3385 2805
rect 3355 2780 3385 2785
rect 3535 2805 3565 2810
rect 3535 2785 3540 2805
rect 3540 2785 3560 2805
rect 3560 2785 3565 2805
rect 3535 2780 3565 2785
rect 3715 2805 3745 2810
rect 3715 2785 3720 2805
rect 3720 2785 3740 2805
rect 3740 2785 3745 2805
rect 3715 2780 3745 2785
rect 3895 2805 3925 2810
rect 3895 2785 3900 2805
rect 3900 2785 3920 2805
rect 3920 2785 3925 2805
rect 3895 2780 3925 2785
rect 4075 2805 4105 2810
rect 4075 2785 4080 2805
rect 4080 2785 4100 2805
rect 4100 2785 4105 2805
rect 4075 2780 4105 2785
rect 4255 2805 4285 2810
rect 4255 2785 4260 2805
rect 4260 2785 4280 2805
rect 4280 2785 4285 2805
rect 4255 2780 4285 2785
rect 4435 2805 4465 2810
rect 4435 2785 4440 2805
rect 4440 2785 4460 2805
rect 4460 2785 4465 2805
rect 4435 2780 4465 2785
rect 4615 2805 4645 2810
rect 4615 2785 4620 2805
rect 4620 2785 4640 2805
rect 4640 2785 4645 2805
rect 4615 2780 4645 2785
rect 4795 2805 4825 2810
rect 4795 2785 4800 2805
rect 4800 2785 4820 2805
rect 4820 2785 4825 2805
rect 4795 2780 4825 2785
rect 4975 2805 5005 2810
rect 4975 2785 4980 2805
rect 4980 2785 5000 2805
rect 5000 2785 5005 2805
rect 4975 2780 5005 2785
rect 2995 2745 3025 2750
rect 2995 2725 3000 2745
rect 3000 2725 3020 2745
rect 3020 2725 3025 2745
rect 2995 2720 3025 2725
rect 3175 2745 3205 2750
rect 3175 2725 3180 2745
rect 3180 2725 3200 2745
rect 3200 2725 3205 2745
rect 3175 2720 3205 2725
rect 3355 2745 3385 2750
rect 3355 2725 3360 2745
rect 3360 2725 3380 2745
rect 3380 2725 3385 2745
rect 3355 2720 3385 2725
rect 3535 2745 3565 2750
rect 3535 2725 3540 2745
rect 3540 2725 3560 2745
rect 3560 2725 3565 2745
rect 3535 2720 3565 2725
rect 3715 2745 3745 2750
rect 3715 2725 3720 2745
rect 3720 2725 3740 2745
rect 3740 2725 3745 2745
rect 3715 2720 3745 2725
rect 3895 2745 3925 2750
rect 3895 2725 3900 2745
rect 3900 2725 3920 2745
rect 3920 2725 3925 2745
rect 3895 2720 3925 2725
rect 4075 2745 4105 2750
rect 4075 2725 4080 2745
rect 4080 2725 4100 2745
rect 4100 2725 4105 2745
rect 4075 2720 4105 2725
rect 4255 2745 4285 2750
rect 4255 2725 4260 2745
rect 4260 2725 4280 2745
rect 4280 2725 4285 2745
rect 4255 2720 4285 2725
rect 4435 2745 4465 2750
rect 4435 2725 4440 2745
rect 4440 2725 4460 2745
rect 4460 2725 4465 2745
rect 4435 2720 4465 2725
rect 4615 2745 4645 2750
rect 4615 2725 4620 2745
rect 4620 2725 4640 2745
rect 4640 2725 4645 2745
rect 4615 2720 4645 2725
rect 4795 2745 4825 2750
rect 4795 2725 4800 2745
rect 4800 2725 4820 2745
rect 4820 2725 4825 2745
rect 4795 2720 4825 2725
rect 4975 2745 5005 2750
rect 4975 2725 4980 2745
rect 4980 2725 5000 2745
rect 5000 2725 5005 2745
rect 4975 2720 5005 2725
rect 2995 2370 3025 2375
rect 2995 2350 3000 2370
rect 3000 2350 3020 2370
rect 3020 2350 3025 2370
rect 2995 2345 3025 2350
rect 3085 2375 3115 2380
rect 3085 2355 3090 2375
rect 3090 2355 3110 2375
rect 3110 2355 3115 2375
rect 3085 2350 3115 2355
rect 3805 2375 3835 2380
rect 3805 2355 3810 2375
rect 3810 2355 3830 2375
rect 3830 2355 3835 2375
rect 3805 2350 3835 2355
rect 4155 2375 4185 2380
rect 4155 2355 4160 2375
rect 4160 2355 4180 2375
rect 4180 2355 4185 2375
rect 4155 2350 4185 2355
rect 4885 2375 4915 2380
rect 4885 2355 4890 2375
rect 4890 2355 4910 2375
rect 4910 2355 4915 2375
rect 4885 2350 4915 2355
rect 2740 2260 2770 2290
rect 3265 2330 3295 2335
rect 3265 2310 3270 2330
rect 3270 2310 3290 2330
rect 3290 2310 3295 2330
rect 3265 2305 3295 2310
rect 3085 2215 3115 2245
rect 2905 2170 2935 2200
rect 3625 2330 3655 2335
rect 3625 2310 3630 2330
rect 3630 2310 3650 2330
rect 3650 2310 3655 2330
rect 3625 2305 3655 2310
rect 3445 2285 3475 2290
rect 3445 2265 3450 2285
rect 3450 2265 3470 2285
rect 3470 2265 3475 2285
rect 3445 2260 3475 2265
rect 3265 2120 3295 2150
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4345 2330 4375 2335
rect 4345 2310 4350 2330
rect 4350 2310 4370 2330
rect 4370 2310 4375 2330
rect 4345 2305 4375 2310
rect 4705 2330 4735 2335
rect 4705 2310 4710 2330
rect 4710 2310 4730 2330
rect 4730 2310 4735 2330
rect 4705 2305 4735 2310
rect 4525 2285 4555 2290
rect 4525 2265 4530 2285
rect 4530 2265 4550 2285
rect 4550 2265 4555 2285
rect 4525 2260 4555 2265
rect 5255 2260 5285 2290
rect 3985 2170 4015 2200
rect 5065 2170 5095 2200
rect 4080 2115 4110 2145
rect 4140 2090 4170 2095
rect 4140 2070 4145 2090
rect 4145 2070 4165 2090
rect 4165 2070 4170 2090
rect 4140 2065 4170 2070
rect 4260 2090 4290 2095
rect 4260 2070 4265 2090
rect 4265 2070 4285 2090
rect 4285 2070 4290 2090
rect 4260 2065 4290 2070
rect 4380 2090 4410 2095
rect 4380 2070 4385 2090
rect 4385 2070 4405 2090
rect 4405 2070 4410 2090
rect 4380 2065 4410 2070
rect 4500 2090 4530 2095
rect 4500 2070 4505 2090
rect 4505 2070 4525 2090
rect 4525 2070 4530 2090
rect 4500 2065 4530 2070
rect 4620 2090 4650 2095
rect 4620 2070 4625 2090
rect 4625 2070 4645 2090
rect 4645 2070 4650 2090
rect 4620 2065 4650 2070
rect 4740 2090 4770 2095
rect 4740 2070 4745 2090
rect 4745 2070 4765 2090
rect 4765 2070 4770 2090
rect 4740 2065 4770 2070
rect 4860 2090 4890 2095
rect 4860 2070 4865 2090
rect 4865 2070 4885 2090
rect 4885 2070 4890 2090
rect 4860 2065 4890 2070
rect 4980 2090 5010 2095
rect 4980 2070 4985 2090
rect 4985 2070 5005 2090
rect 5005 2070 5010 2090
rect 4980 2065 5010 2070
rect 5100 2090 5130 2095
rect 5100 2070 5105 2090
rect 5105 2070 5125 2090
rect 5125 2070 5130 2090
rect 5100 2065 5130 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 4080 2045 4110 2050
rect 4080 2025 4085 2045
rect 4085 2025 4105 2045
rect 4105 2025 4110 2045
rect 4080 2020 4110 2025
rect 4440 2045 4470 2050
rect 4440 2025 4445 2045
rect 4445 2025 4465 2045
rect 4465 2025 4470 2045
rect 4440 2020 4470 2025
rect 4800 2045 4830 2050
rect 4800 2025 4805 2045
rect 4805 2025 4825 2045
rect 4825 2025 4830 2045
rect 4800 2020 4830 2025
rect 5160 2045 5190 2050
rect 5160 2025 5165 2045
rect 5165 2025 5185 2045
rect 5185 2025 5190 2045
rect 5160 2020 5190 2025
rect 4320 1875 4350 1880
rect 4320 1855 4325 1875
rect 4325 1855 4345 1875
rect 4345 1855 4350 1875
rect 4320 1850 4350 1855
rect 4680 1875 4710 1880
rect 4680 1855 4685 1875
rect 4685 1855 4705 1875
rect 4705 1855 4710 1875
rect 4680 1850 4710 1855
rect 5040 1875 5070 1880
rect 5040 1855 5045 1875
rect 5045 1855 5065 1875
rect 5065 1855 5070 1875
rect 5040 1850 5070 1855
rect 4110 1790 4140 1820
rect 4200 1815 4230 1820
rect 4200 1795 4205 1815
rect 4205 1795 4225 1815
rect 4225 1795 4230 1815
rect 4200 1790 4230 1795
rect 4440 1790 4470 1820
rect 4560 1815 4590 1820
rect 4560 1795 4565 1815
rect 4565 1795 4585 1815
rect 4585 1795 4590 1815
rect 4560 1790 4590 1795
rect 4200 1755 4230 1760
rect 4200 1735 4205 1755
rect 4205 1735 4225 1755
rect 4225 1735 4230 1755
rect 4200 1730 4230 1735
rect 4440 1755 4470 1760
rect 4440 1735 4445 1755
rect 4445 1735 4465 1755
rect 4465 1735 4470 1755
rect 4440 1730 4470 1735
rect 4800 1790 4830 1820
rect 4920 1815 4950 1820
rect 4920 1795 4925 1815
rect 4925 1795 4945 1815
rect 4945 1795 4950 1815
rect 4920 1790 4950 1795
rect 5130 1790 5160 1820
rect 5300 2115 5330 2145
rect 5395 3255 5425 3285
rect 5345 1790 5375 1820
rect 4680 1755 4710 1760
rect 4680 1735 4685 1755
rect 4685 1735 4705 1755
rect 4705 1735 4710 1755
rect 4680 1730 4710 1735
rect 4740 1755 4770 1760
rect 4740 1735 4745 1755
rect 4745 1735 4765 1755
rect 4765 1735 4770 1755
rect 4740 1730 4770 1735
rect 5255 1730 5285 1760
rect 4320 1710 4350 1715
rect 4320 1690 4325 1710
rect 4325 1690 4345 1710
rect 4345 1690 4350 1710
rect 4320 1685 4350 1690
rect 4560 1710 4590 1715
rect 4560 1690 4565 1710
rect 4565 1690 4585 1710
rect 4585 1690 4590 1710
rect 4560 1685 4590 1690
rect 4800 1710 4830 1715
rect 4800 1690 4805 1710
rect 4805 1690 4825 1710
rect 4825 1690 4830 1710
rect 4800 1685 4830 1690
rect 4800 1590 4830 1595
rect 4800 1570 4805 1590
rect 4805 1570 4825 1590
rect 4825 1570 4830 1590
rect 4800 1565 4830 1570
rect 5395 1565 5425 1595
rect 4260 1540 4290 1545
rect 4260 1520 4265 1540
rect 4265 1520 4285 1540
rect 4285 1520 4290 1540
rect 4260 1515 4290 1520
rect 4380 1540 4410 1545
rect 4380 1520 4385 1540
rect 4385 1520 4405 1540
rect 4405 1520 4410 1540
rect 4380 1515 4410 1520
rect 4500 1540 4530 1545
rect 4500 1520 4505 1540
rect 4505 1520 4525 1540
rect 4525 1520 4530 1540
rect 4500 1515 4530 1520
rect 4620 1540 4650 1545
rect 4620 1520 4625 1540
rect 4625 1520 4645 1540
rect 4645 1520 4650 1540
rect 4620 1515 4650 1520
rect 4740 1540 4770 1545
rect 4740 1520 4745 1540
rect 4745 1520 4765 1540
rect 4765 1520 4770 1540
rect 4740 1515 4770 1520
rect 5130 1515 5160 1545
rect 3380 1185 3410 1190
rect 3380 1165 3385 1185
rect 3385 1165 3405 1185
rect 3405 1165 3410 1185
rect 3380 1160 3410 1165
rect 4590 1185 4620 1190
rect 4590 1165 4595 1185
rect 4595 1165 4615 1185
rect 4615 1165 4620 1185
rect 4590 1160 4620 1165
rect 2945 1125 2975 1130
rect 2945 1105 2950 1125
rect 2950 1105 2970 1125
rect 2970 1105 2975 1125
rect 2945 1100 2975 1105
rect 3025 1125 3055 1130
rect 3025 1105 3030 1125
rect 3030 1105 3050 1125
rect 3050 1105 3055 1125
rect 3025 1100 3055 1105
rect 3105 1125 3135 1130
rect 3105 1105 3110 1125
rect 3110 1105 3130 1125
rect 3130 1105 3135 1125
rect 3105 1100 3135 1105
rect 3185 1125 3215 1130
rect 3185 1105 3190 1125
rect 3190 1105 3210 1125
rect 3210 1105 3215 1125
rect 3185 1100 3215 1105
rect 3265 1125 3295 1130
rect 3265 1105 3270 1125
rect 3270 1105 3290 1125
rect 3290 1105 3295 1125
rect 3265 1100 3295 1105
rect 3345 1125 3375 1130
rect 3345 1105 3350 1125
rect 3350 1105 3370 1125
rect 3370 1105 3375 1125
rect 3345 1100 3375 1105
rect 3425 1125 3455 1130
rect 3425 1105 3430 1125
rect 3430 1105 3450 1125
rect 3450 1105 3455 1125
rect 3425 1100 3455 1105
rect 3505 1125 3535 1130
rect 3505 1105 3510 1125
rect 3510 1105 3530 1125
rect 3530 1105 3535 1125
rect 3505 1100 3535 1105
rect 3585 1125 3615 1130
rect 3585 1105 3590 1125
rect 3590 1105 3610 1125
rect 3610 1105 3615 1125
rect 3585 1100 3615 1105
rect 3665 1125 3695 1130
rect 3665 1105 3670 1125
rect 3670 1105 3690 1125
rect 3690 1105 3695 1125
rect 3665 1100 3695 1105
rect 3745 1125 3775 1130
rect 3745 1105 3750 1125
rect 3750 1105 3770 1125
rect 3770 1105 3775 1125
rect 3745 1100 3775 1105
rect 3825 1125 3855 1130
rect 3825 1105 3830 1125
rect 3830 1105 3850 1125
rect 3850 1105 3855 1125
rect 3825 1100 3855 1105
rect 3905 1125 3935 1130
rect 3905 1105 3910 1125
rect 3910 1105 3930 1125
rect 3930 1105 3935 1125
rect 3905 1100 3935 1105
rect 3985 1125 4015 1130
rect 3985 1105 3990 1125
rect 3990 1105 4010 1125
rect 4010 1105 4015 1125
rect 3985 1100 4015 1105
rect 4065 1125 4095 1130
rect 4065 1105 4070 1125
rect 4070 1105 4090 1125
rect 4090 1105 4095 1125
rect 4065 1100 4095 1105
rect 4145 1125 4175 1130
rect 4145 1105 4150 1125
rect 4150 1105 4170 1125
rect 4170 1105 4175 1125
rect 4145 1100 4175 1105
rect 4225 1125 4255 1130
rect 4225 1105 4230 1125
rect 4230 1105 4250 1125
rect 4250 1105 4255 1125
rect 4225 1100 4255 1105
rect 4305 1125 4335 1130
rect 4305 1105 4310 1125
rect 4310 1105 4330 1125
rect 4330 1105 4335 1125
rect 4305 1100 4335 1105
rect 4385 1125 4415 1130
rect 4385 1105 4390 1125
rect 4390 1105 4410 1125
rect 4410 1105 4415 1125
rect 4385 1100 4415 1105
rect 4465 1125 4495 1130
rect 4465 1105 4470 1125
rect 4470 1105 4490 1125
rect 4490 1105 4495 1125
rect 4465 1100 4495 1105
rect 4545 1125 4575 1130
rect 4545 1105 4550 1125
rect 4550 1105 4570 1125
rect 4570 1105 4575 1125
rect 4545 1100 4575 1105
rect 4625 1125 4655 1130
rect 4625 1105 4630 1125
rect 4630 1105 4650 1125
rect 4650 1105 4655 1125
rect 4625 1100 4655 1105
rect 4705 1125 4735 1130
rect 4705 1105 4710 1125
rect 4710 1105 4730 1125
rect 4730 1105 4735 1125
rect 4705 1100 4735 1105
rect 4785 1125 4815 1130
rect 4785 1105 4790 1125
rect 4790 1105 4810 1125
rect 4810 1105 4815 1125
rect 4785 1100 4815 1105
rect 4865 1125 4895 1130
rect 4865 1105 4870 1125
rect 4870 1105 4890 1125
rect 4890 1105 4895 1125
rect 4865 1100 4895 1105
rect 4945 1125 4975 1130
rect 4945 1105 4950 1125
rect 4950 1105 4970 1125
rect 4970 1105 4975 1125
rect 4945 1100 4975 1105
rect 2625 1015 2655 1045
rect 2905 1040 2935 1045
rect 2905 1020 2910 1040
rect 2910 1020 2930 1040
rect 2930 1020 2935 1040
rect 2905 1015 2935 1020
rect 5060 1040 5090 1045
rect 5060 1020 5065 1040
rect 5065 1020 5085 1040
rect 5085 1020 5090 1040
rect 5060 1015 5090 1020
rect 2995 930 3025 935
rect 2995 910 3000 930
rect 3000 910 3020 930
rect 3020 910 3025 930
rect 2995 905 3025 910
rect 3175 930 3205 935
rect 3175 910 3180 930
rect 3180 910 3200 930
rect 3200 910 3205 930
rect 3175 905 3205 910
rect 3355 930 3385 935
rect 3355 910 3360 930
rect 3360 910 3380 930
rect 3380 910 3385 930
rect 3355 905 3385 910
rect 3535 930 3565 935
rect 3535 910 3540 930
rect 3540 910 3560 930
rect 3560 910 3565 930
rect 3535 905 3565 910
rect 3715 930 3745 935
rect 3715 910 3720 930
rect 3720 910 3740 930
rect 3740 910 3745 930
rect 3715 905 3745 910
rect 3895 930 3925 935
rect 3895 910 3900 930
rect 3900 910 3920 930
rect 3920 910 3925 930
rect 3895 905 3925 910
rect 4075 930 4105 935
rect 4075 910 4080 930
rect 4080 910 4100 930
rect 4100 910 4105 930
rect 4075 905 4105 910
rect 4255 930 4285 935
rect 4255 910 4260 930
rect 4260 910 4280 930
rect 4280 910 4285 930
rect 4255 905 4285 910
rect 4435 930 4465 935
rect 4435 910 4440 930
rect 4440 910 4460 930
rect 4460 910 4465 930
rect 4435 905 4465 910
rect 4615 930 4645 935
rect 4615 910 4620 930
rect 4620 910 4640 930
rect 4640 910 4645 930
rect 4615 905 4645 910
rect 4795 930 4825 935
rect 4795 910 4800 930
rect 4800 910 4820 930
rect 4820 910 4825 930
rect 4795 905 4825 910
rect 4975 930 5005 935
rect 4975 910 4980 930
rect 4980 910 5000 930
rect 5000 910 5005 930
rect 4975 905 5005 910
rect 2525 720 2555 750
rect 3085 745 3115 750
rect 3085 725 3090 745
rect 3090 725 3110 745
rect 3110 725 3115 745
rect 3085 720 3115 725
rect 3625 760 3655 765
rect 3625 740 3630 760
rect 3630 740 3650 760
rect 3650 740 3655 760
rect 3625 735 3655 740
rect 3985 760 4015 765
rect 3985 740 3990 760
rect 3990 740 4010 760
rect 4010 740 4015 760
rect 3985 735 4015 740
rect 4345 760 4375 765
rect 4345 740 4350 760
rect 4350 740 4370 760
rect 4370 740 4375 760
rect 4345 735 4375 740
rect 4525 760 4555 765
rect 4525 740 4530 760
rect 4530 740 4550 760
rect 4550 740 4555 760
rect 4525 735 4555 740
rect 4705 760 4735 765
rect 4705 740 4710 760
rect 4710 740 4730 760
rect 4730 740 4735 760
rect 4705 735 4735 740
rect 4885 760 4915 765
rect 4885 740 4890 760
rect 4890 740 4910 760
rect 4910 740 4915 760
rect 4885 735 4915 740
rect 3445 680 3475 710
rect 3805 680 3835 710
rect 4165 680 4195 710
<< metal2 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5530 4990 5570 4995
rect 5530 4960 5535 4990
rect 5565 4960 5570 4990
rect 5530 4955 5570 4960
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1245 3525 1285 3530
rect 1245 3520 1250 3525
rect -75 3500 1250 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1245 3495 1250 3500
rect 1280 3495 1285 3525
rect 1245 3490 1285 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5530 3445 5570 3450
rect 5530 3440 5535 3445
rect 5175 3420 5535 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5530 3415 5535 3420
rect 5565 3415 5570 3445
rect 5530 3410 5570 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1190 3340 1230 3345
rect 1190 3310 1195 3340
rect 1225 3335 1230 3340
rect 3130 3340 3170 3345
rect 3130 3335 3135 3340
rect 1225 3315 3135 3335
rect 1225 3310 1230 3315
rect 1190 3305 1230 3310
rect 3130 3310 3135 3315
rect 3165 3310 3170 3340
rect 3130 3305 3170 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5340 3335 5380 3340
rect 5340 3330 5345 3335
rect 3425 3310 5345 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5340 3305 5345 3310
rect 5375 3305 5380 3335
rect 5340 3300 5380 3305
rect 1145 3285 1185 3290
rect 1145 3255 1150 3285
rect 1180 3280 1185 3285
rect 4880 3285 4920 3290
rect 4880 3280 4885 3285
rect 1180 3260 4885 3280
rect 1180 3255 1185 3260
rect 1145 3250 1185 3255
rect 4880 3255 4885 3260
rect 4915 3280 4920 3285
rect 5390 3285 5430 3290
rect 5390 3280 5395 3285
rect 4915 3260 5395 3280
rect 4915 3255 4920 3260
rect 4880 3250 4920 3255
rect 5390 3255 5395 3260
rect 5425 3255 5430 3285
rect 5390 3250 5430 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 40 3215 2740 3235
rect 40 3205 85 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 40 3170 45 3205
rect 80 3170 85 3205
rect 1245 3165 1250 3200
rect 1285 3165 1290 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 40 3135 45 3145
rect -75 3115 45 3135
rect -75 3110 -70 3115
rect 40 3110 45 3115
rect 80 3110 85 3145
rect 3130 3140 3170 3145
rect -110 3105 -70 3110
rect 1245 3105 1250 3140
rect 1285 3105 1290 3140
rect 3130 3110 3135 3140
rect 3165 3135 3170 3140
rect 4830 3140 4870 3145
rect 4830 3135 4835 3140
rect 3165 3115 4835 3135
rect 3165 3110 3170 3115
rect 3130 3105 3170 3110
rect 4830 3110 4835 3115
rect 4865 3135 4870 3140
rect 5295 3140 5335 3145
rect 5295 3135 5300 3140
rect 4865 3115 5300 3135
rect 4865 3110 4870 3115
rect 4830 3105 4870 3110
rect 5295 3110 5300 3115
rect 5330 3110 5335 3140
rect 5295 3105 5335 3110
rect 1145 3100 1185 3105
rect 1145 3095 1150 3100
rect 40 3075 1150 3095
rect 40 3065 85 3075
rect 1145 3070 1150 3075
rect 1180 3070 1185 3100
rect 1145 3065 1185 3070
rect 3980 3080 4020 3085
rect 40 3030 45 3065
rect 80 3030 85 3065
rect 3980 3050 3985 3080
rect 4015 3075 4020 3080
rect 4015 3055 6080 3075
rect 4015 3050 4020 3055
rect 3980 3045 4020 3050
rect 3440 3035 3480 3040
rect 3440 3005 3445 3035
rect 3475 3030 3480 3035
rect 3800 3035 3840 3040
rect 3800 3030 3805 3035
rect 3475 3010 3805 3030
rect 3475 3005 3480 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 40 2995 45 3005
rect -75 2975 45 2995
rect -75 2970 -70 2975
rect 40 2970 45 2975
rect 80 2970 85 3005
rect 3440 3000 3480 3005
rect 3800 3005 3805 3010
rect 3835 3030 3840 3035
rect 4340 3035 4380 3040
rect 4340 3030 4345 3035
rect 3835 3010 4345 3030
rect 3835 3005 3840 3010
rect 3800 3000 3840 3005
rect 4340 3005 4345 3010
rect 4375 3030 4380 3035
rect 4700 3035 4740 3040
rect 4700 3030 4705 3035
rect 4375 3010 4705 3030
rect 4375 3005 4380 3010
rect 4340 3000 4380 3005
rect 4700 3005 4705 3010
rect 4735 3030 4740 3035
rect 4735 3010 6080 3030
rect 4735 3005 4740 3010
rect 4700 3000 4740 3005
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3075 2980 3115 2985
rect 3075 2975 3080 2980
rect 2555 2955 3080 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3075 2950 3080 2955
rect 3110 2950 3115 2980
rect 3075 2945 3115 2950
rect 3260 2980 3300 2985
rect 3260 2950 3265 2980
rect 3295 2975 3300 2980
rect 3620 2980 3660 2985
rect 3620 2975 3625 2980
rect 3295 2955 3625 2975
rect 3295 2950 3300 2955
rect 3260 2945 3300 2950
rect 3620 2950 3625 2955
rect 3655 2975 3660 2980
rect 4160 2980 4200 2985
rect 4160 2975 4165 2980
rect 3655 2955 4165 2975
rect 3655 2950 3660 2955
rect 3620 2945 3660 2950
rect 4160 2950 4165 2955
rect 4195 2975 4200 2980
rect 4520 2980 4560 2985
rect 4520 2975 4525 2980
rect 4195 2955 4525 2975
rect 4195 2950 4200 2955
rect 4160 2945 4200 2950
rect 4520 2950 4525 2955
rect 4555 2975 4560 2980
rect 4555 2955 6080 2975
rect 4555 2950 4560 2955
rect 4520 2945 4560 2950
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 40 2850 45 2855
rect -25 2830 45 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 40 2820 45 2830
rect 80 2820 85 2855
rect 575 2820 580 2855
rect 615 2845 620 2855
rect 1190 2850 1230 2855
rect 1190 2845 1195 2850
rect 615 2825 1195 2845
rect 615 2820 620 2825
rect 1190 2820 1195 2825
rect 1225 2820 1230 2850
rect 1190 2815 1230 2820
rect 1245 2805 1250 2840
rect 1285 2805 1290 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 2330 2800 2370 2805
rect 2990 2810 3030 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 40 2785 45 2795
rect 20 2765 45 2785
rect -15 2760 25 2765
rect 40 2760 45 2765
rect 80 2760 85 2795
rect 575 2760 580 2795
rect 615 2785 620 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 615 2765 2625 2785
rect 615 2760 620 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2990 2780 2995 2810
rect 3025 2805 3030 2810
rect 3170 2810 3210 2815
rect 3170 2805 3175 2810
rect 3025 2785 3175 2805
rect 3025 2780 3030 2785
rect 2990 2775 3030 2780
rect 3170 2780 3175 2785
rect 3205 2805 3210 2810
rect 3350 2810 3390 2815
rect 3350 2805 3355 2810
rect 3205 2785 3355 2805
rect 3205 2780 3210 2785
rect 3170 2775 3210 2780
rect 3350 2780 3355 2785
rect 3385 2805 3390 2810
rect 3530 2810 3570 2815
rect 3530 2805 3535 2810
rect 3385 2785 3535 2805
rect 3385 2780 3390 2785
rect 3350 2775 3390 2780
rect 3530 2780 3535 2785
rect 3565 2805 3570 2810
rect 3710 2810 3750 2815
rect 3710 2805 3715 2810
rect 3565 2785 3715 2805
rect 3565 2780 3570 2785
rect 3530 2775 3570 2780
rect 3710 2780 3715 2785
rect 3745 2805 3750 2810
rect 3890 2810 3930 2815
rect 3890 2805 3895 2810
rect 3745 2785 3895 2805
rect 3745 2780 3750 2785
rect 3710 2775 3750 2780
rect 3890 2780 3895 2785
rect 3925 2805 3930 2810
rect 4070 2810 4110 2815
rect 4070 2805 4075 2810
rect 3925 2785 4075 2805
rect 3925 2780 3930 2785
rect 3890 2775 3930 2780
rect 4070 2780 4075 2785
rect 4105 2805 4110 2810
rect 4250 2810 4290 2815
rect 4250 2805 4255 2810
rect 4105 2785 4255 2805
rect 4105 2780 4110 2785
rect 4070 2775 4110 2780
rect 4250 2780 4255 2785
rect 4285 2805 4290 2810
rect 4430 2810 4470 2815
rect 4430 2805 4435 2810
rect 4285 2785 4435 2805
rect 4285 2780 4290 2785
rect 4250 2775 4290 2780
rect 4430 2780 4435 2785
rect 4465 2805 4470 2810
rect 4610 2810 4650 2815
rect 4610 2805 4615 2810
rect 4465 2785 4615 2805
rect 4465 2780 4470 2785
rect 4430 2775 4470 2780
rect 4610 2780 4615 2785
rect 4645 2805 4650 2810
rect 4790 2810 4830 2815
rect 4790 2805 4795 2810
rect 4645 2785 4795 2805
rect 4645 2780 4650 2785
rect 4610 2775 4650 2780
rect 4790 2780 4795 2785
rect 4825 2805 4830 2810
rect 4970 2810 5010 2815
rect 4970 2805 4975 2810
rect 4825 2785 4975 2805
rect 4825 2780 4830 2785
rect 4790 2775 4830 2780
rect 4970 2780 4975 2785
rect 5005 2805 5010 2810
rect 5530 2810 5570 2815
rect 5530 2805 5535 2810
rect 5005 2785 5535 2805
rect 5005 2780 5010 2785
rect 4970 2775 5010 2780
rect 5530 2780 5535 2785
rect 5565 2780 5570 2810
rect 5530 2775 5570 2780
rect 2620 2755 2660 2760
rect 2990 2750 3030 2755
rect 1245 2745 1285 2750
rect 1245 2715 1250 2745
rect 1280 2740 1285 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1280 2720 2155 2740
rect 1280 2715 1285 2720
rect 1245 2710 1285 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 2990 2720 2995 2750
rect 3025 2745 3030 2750
rect 3170 2750 3210 2755
rect 3170 2745 3175 2750
rect 3025 2725 3175 2745
rect 3025 2720 3030 2725
rect 2990 2715 3030 2720
rect 3170 2720 3175 2725
rect 3205 2745 3210 2750
rect 3350 2750 3390 2755
rect 3350 2745 3355 2750
rect 3205 2725 3355 2745
rect 3205 2720 3210 2725
rect 3170 2715 3210 2720
rect 3350 2720 3355 2725
rect 3385 2745 3390 2750
rect 3530 2750 3570 2755
rect 3530 2745 3535 2750
rect 3385 2725 3535 2745
rect 3385 2720 3390 2725
rect 3350 2715 3390 2720
rect 3530 2720 3535 2725
rect 3565 2745 3570 2750
rect 3710 2750 3750 2755
rect 3710 2745 3715 2750
rect 3565 2725 3715 2745
rect 3565 2720 3570 2725
rect 3530 2715 3570 2720
rect 3710 2720 3715 2725
rect 3745 2745 3750 2750
rect 3890 2750 3930 2755
rect 3890 2745 3895 2750
rect 3745 2725 3895 2745
rect 3745 2720 3750 2725
rect 3710 2715 3750 2720
rect 3890 2720 3895 2725
rect 3925 2745 3930 2750
rect 4070 2750 4110 2755
rect 4070 2745 4075 2750
rect 3925 2725 4075 2745
rect 3925 2720 3930 2725
rect 3890 2715 3930 2720
rect 4070 2720 4075 2725
rect 4105 2745 4110 2750
rect 4250 2750 4290 2755
rect 4250 2745 4255 2750
rect 4105 2725 4255 2745
rect 4105 2720 4110 2725
rect 4070 2715 4110 2720
rect 4250 2720 4255 2725
rect 4285 2745 4290 2750
rect 4430 2750 4470 2755
rect 4430 2745 4435 2750
rect 4285 2725 4435 2745
rect 4285 2720 4290 2725
rect 4250 2715 4290 2720
rect 4430 2720 4435 2725
rect 4465 2745 4470 2750
rect 4610 2750 4650 2755
rect 4610 2745 4615 2750
rect 4465 2725 4615 2745
rect 4465 2720 4470 2725
rect 4430 2715 4470 2720
rect 4610 2720 4615 2725
rect 4645 2745 4650 2750
rect 4790 2750 4830 2755
rect 4790 2745 4795 2750
rect 4645 2725 4795 2745
rect 4645 2720 4650 2725
rect 4610 2715 4650 2720
rect 4790 2720 4795 2725
rect 4825 2745 4830 2750
rect 4970 2750 5010 2755
rect 4970 2745 4975 2750
rect 4825 2725 4975 2745
rect 4825 2720 4830 2725
rect 4790 2715 4830 2720
rect 4970 2720 4975 2725
rect 5005 2720 5010 2750
rect 4970 2715 5010 2720
rect 2150 2710 2190 2715
rect 3080 2380 3120 2385
rect 2990 2375 3030 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 2990 2345 2995 2375
rect 3025 2345 3030 2375
rect 3080 2350 3085 2380
rect 3115 2375 3120 2380
rect 3800 2380 3840 2385
rect 3800 2375 3805 2380
rect 3115 2355 3805 2375
rect 3115 2350 3120 2355
rect 3080 2345 3120 2350
rect 3800 2350 3805 2355
rect 3835 2375 3840 2380
rect 4150 2380 4190 2385
rect 4150 2375 4155 2380
rect 3835 2355 4155 2375
rect 3835 2350 3840 2355
rect 3800 2345 3840 2350
rect 4150 2350 4155 2355
rect 4185 2375 4190 2380
rect 4880 2380 4920 2385
rect 4880 2375 4885 2380
rect 4185 2355 4885 2375
rect 4185 2350 4190 2355
rect 4150 2345 4190 2350
rect 4880 2350 4885 2355
rect 4915 2350 4920 2380
rect 4880 2345 4920 2350
rect 2990 2340 3030 2345
rect 2655 2320 3030 2340
rect 3260 2335 3300 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3260 2305 3265 2335
rect 3295 2330 3300 2335
rect 3620 2335 3660 2340
rect 3620 2330 3625 2335
rect 3295 2310 3625 2330
rect 3295 2305 3300 2310
rect 3260 2300 3300 2305
rect 3620 2305 3625 2310
rect 3655 2330 3660 2335
rect 4340 2335 4380 2340
rect 4340 2330 4345 2335
rect 3655 2310 4345 2330
rect 3655 2305 3660 2310
rect 3620 2300 3660 2305
rect 4340 2305 4345 2310
rect 4375 2330 4380 2335
rect 4700 2335 4740 2340
rect 4700 2330 4705 2335
rect 4375 2310 4705 2330
rect 4375 2305 4380 2310
rect 4340 2300 4380 2305
rect 4700 2305 4705 2310
rect 4735 2305 4740 2335
rect 4700 2300 4740 2305
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3440 2290 3480 2295
rect 3440 2285 3445 2290
rect 2770 2265 3445 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3440 2260 3445 2265
rect 3475 2285 3480 2290
rect 4520 2290 4560 2295
rect 4520 2285 4525 2290
rect 3475 2265 4525 2285
rect 3475 2260 3480 2265
rect 3440 2255 3480 2260
rect 4520 2260 4525 2265
rect 4555 2285 4560 2290
rect 5250 2290 5290 2295
rect 5250 2285 5255 2290
rect 4555 2265 5255 2285
rect 4555 2260 4560 2265
rect 4520 2255 4560 2260
rect 5250 2260 5255 2265
rect 5285 2260 5290 2290
rect 5250 2255 5290 2260
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3080 2245 3120 2250
rect 3080 2240 3085 2245
rect 2460 2220 3085 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3080 2215 3085 2220
rect 3115 2215 3120 2245
rect 3080 2210 3120 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 2900 2200 2940 2205
rect 2900 2195 2905 2200
rect 2365 2175 2905 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 2900 2170 2905 2175
rect 2935 2195 2940 2200
rect 3980 2200 4020 2205
rect 3980 2195 3985 2200
rect 2935 2175 3985 2195
rect 2935 2170 2940 2175
rect 2900 2165 2940 2170
rect 3980 2170 3985 2175
rect 4015 2195 4020 2200
rect 5060 2200 5100 2205
rect 5060 2195 5065 2200
rect 4015 2175 5065 2195
rect 4015 2170 4020 2175
rect 3980 2165 4020 2170
rect 5060 2170 5065 2175
rect 5095 2170 5100 2200
rect 5060 2165 5100 2170
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3260 2150 3300 2155
rect 3260 2145 3265 2150
rect 2415 2125 3265 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3260 2120 3265 2125
rect 3295 2120 3300 2150
rect 3260 2115 3300 2120
rect 4075 2145 4115 2150
rect 4075 2115 4080 2145
rect 4110 2140 4115 2145
rect 5295 2145 5335 2150
rect 5295 2140 5300 2145
rect 4110 2120 5300 2140
rect 4110 2115 4115 2120
rect 4075 2110 4115 2115
rect 5295 2115 5300 2120
rect 5330 2115 5335 2145
rect 5295 2110 5335 2115
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 4135 2095 4175 2100
rect 4135 2065 4140 2095
rect 4170 2090 4175 2095
rect 4255 2095 4295 2100
rect 4255 2090 4260 2095
rect 4170 2070 4260 2090
rect 4170 2065 4175 2070
rect 4135 2060 4175 2065
rect 4255 2065 4260 2070
rect 4290 2090 4295 2095
rect 4375 2095 4415 2100
rect 4375 2090 4380 2095
rect 4290 2070 4380 2090
rect 4290 2065 4295 2070
rect 4255 2060 4295 2065
rect 4375 2065 4380 2070
rect 4410 2090 4415 2095
rect 4495 2095 4535 2100
rect 4495 2090 4500 2095
rect 4410 2070 4500 2090
rect 4410 2065 4415 2070
rect 4375 2060 4415 2065
rect 4495 2065 4500 2070
rect 4530 2090 4535 2095
rect 4615 2095 4655 2100
rect 4615 2090 4620 2095
rect 4530 2070 4620 2090
rect 4530 2065 4535 2070
rect 4495 2060 4535 2065
rect 4615 2065 4620 2070
rect 4650 2090 4655 2095
rect 4735 2095 4775 2100
rect 4735 2090 4740 2095
rect 4650 2070 4740 2090
rect 4650 2065 4655 2070
rect 4615 2060 4655 2065
rect 4735 2065 4740 2070
rect 4770 2090 4775 2095
rect 4855 2095 4895 2100
rect 4855 2090 4860 2095
rect 4770 2070 4860 2090
rect 4770 2065 4775 2070
rect 4735 2060 4775 2065
rect 4855 2065 4860 2070
rect 4890 2090 4895 2095
rect 4975 2095 5015 2100
rect 4975 2090 4980 2095
rect 4890 2070 4980 2090
rect 4890 2065 4895 2070
rect 4855 2060 4895 2065
rect 4975 2065 4980 2070
rect 5010 2090 5015 2095
rect 5095 2095 5135 2100
rect 5095 2090 5100 2095
rect 5010 2070 5100 2090
rect 5010 2065 5015 2070
rect 4975 2060 5015 2065
rect 5095 2065 5100 2070
rect 5130 2065 5135 2095
rect 5095 2060 5135 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4075 2050 4115 2055
rect 4075 2020 4080 2050
rect 4110 2045 4115 2050
rect 4435 2050 4475 2055
rect 4435 2045 4440 2050
rect 4110 2025 4440 2045
rect 4110 2020 4115 2025
rect 4075 2015 4115 2020
rect 4435 2020 4440 2025
rect 4470 2045 4475 2050
rect 4795 2050 4835 2055
rect 4795 2045 4800 2050
rect 4470 2025 4800 2045
rect 4470 2020 4475 2025
rect 4435 2015 4475 2020
rect 4795 2020 4800 2025
rect 4830 2045 4835 2050
rect 5155 2050 5195 2055
rect 5155 2045 5160 2050
rect 4830 2025 5160 2045
rect 4830 2020 4835 2025
rect 4795 2015 4835 2020
rect 5155 2020 5160 2025
rect 5190 2020 5195 2050
rect 5155 2015 5195 2020
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4195 1845 4235 1885
rect 4315 1880 4355 1885
rect 4315 1850 4320 1880
rect 4350 1875 4355 1880
rect 4555 1875 4595 1885
rect 4675 1880 4715 1885
rect 4675 1875 4680 1880
rect 4350 1855 4680 1875
rect 4350 1850 4355 1855
rect 4315 1845 4355 1850
rect 4555 1845 4595 1855
rect 4675 1850 4680 1855
rect 4710 1875 4715 1880
rect 4915 1875 4955 1885
rect 5035 1880 5075 1885
rect 5035 1875 5040 1880
rect 4710 1855 5040 1875
rect 4710 1850 4715 1855
rect 4675 1845 4715 1850
rect 4915 1845 4955 1855
rect 5035 1850 5040 1855
rect 5070 1875 5075 1880
rect 5070 1855 5165 1875
rect 5070 1850 5075 1855
rect 5035 1845 5075 1850
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4105 1820 4145 1825
rect 4105 1790 4110 1820
rect 4140 1815 4145 1820
rect 4195 1820 4235 1825
rect 4195 1815 4200 1820
rect 4140 1795 4200 1815
rect 4140 1790 4145 1795
rect 4105 1785 4145 1790
rect 4195 1790 4200 1795
rect 4230 1815 4235 1820
rect 4435 1820 4475 1825
rect 4435 1815 4440 1820
rect 4230 1795 4440 1815
rect 4230 1790 4235 1795
rect 4195 1785 4235 1790
rect 4435 1790 4440 1795
rect 4470 1815 4475 1820
rect 4555 1820 4595 1825
rect 4555 1815 4560 1820
rect 4470 1795 4560 1815
rect 4470 1790 4475 1795
rect 4435 1785 4475 1790
rect 4555 1790 4560 1795
rect 4590 1815 4595 1820
rect 4795 1820 4835 1825
rect 4795 1815 4800 1820
rect 4590 1795 4800 1815
rect 4590 1790 4595 1795
rect 4555 1785 4595 1790
rect 4795 1790 4800 1795
rect 4830 1815 4835 1820
rect 4915 1820 4955 1825
rect 4915 1815 4920 1820
rect 4830 1795 4920 1815
rect 4830 1790 4835 1795
rect 4795 1785 4835 1790
rect 4915 1790 4920 1795
rect 4950 1815 4955 1820
rect 5125 1820 5165 1825
rect 5125 1815 5130 1820
rect 4950 1795 5130 1815
rect 4950 1790 4955 1795
rect 4915 1785 4955 1790
rect 5125 1790 5130 1795
rect 5160 1815 5165 1820
rect 5340 1820 5380 1825
rect 5340 1815 5345 1820
rect 5160 1795 5345 1815
rect 5160 1790 5165 1795
rect 5125 1785 5165 1790
rect 5340 1790 5345 1795
rect 5375 1790 5380 1820
rect 5340 1785 5380 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2710 1735 3230 1755
rect 2710 1730 2715 1735
rect 2675 1725 2715 1730
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4195 1760 4235 1765
rect 4195 1730 4200 1760
rect 4230 1755 4235 1760
rect 4435 1760 4475 1765
rect 4435 1755 4440 1760
rect 4230 1735 4440 1755
rect 4230 1730 4235 1735
rect 4195 1725 4235 1730
rect 4435 1730 4440 1735
rect 4470 1755 4475 1760
rect 4675 1760 4715 1765
rect 4675 1755 4680 1760
rect 4470 1735 4680 1755
rect 4470 1730 4475 1735
rect 4435 1725 4475 1730
rect 4675 1730 4680 1735
rect 4710 1730 4715 1760
rect 4675 1725 4715 1730
rect 4735 1760 4775 1765
rect 4735 1730 4740 1760
rect 4770 1755 4775 1760
rect 5250 1760 5290 1765
rect 5250 1755 5255 1760
rect 4770 1735 5255 1755
rect 4770 1730 4775 1735
rect 4735 1725 4775 1730
rect 5250 1730 5255 1735
rect 5285 1755 5290 1760
rect 5285 1735 6080 1755
rect 5285 1730 5290 1735
rect 5250 1725 5290 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1265 1710 1305 1715
rect 1265 1680 1270 1710
rect 1300 1705 1305 1710
rect 2150 1710 2190 1715
rect 2150 1705 2155 1710
rect 1300 1685 2155 1705
rect 1300 1680 1305 1685
rect 1265 1675 1305 1680
rect 2150 1680 2155 1685
rect 2185 1680 2190 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4315 1715 4355 1720
rect 4315 1685 4320 1715
rect 4350 1710 4355 1715
rect 4555 1715 4595 1720
rect 4555 1710 4560 1715
rect 4350 1690 4560 1710
rect 4350 1685 4355 1690
rect 4315 1680 4355 1685
rect 4555 1685 4560 1690
rect 4590 1710 4595 1715
rect 4795 1715 4835 1720
rect 4795 1710 4800 1715
rect 4590 1690 4800 1710
rect 4590 1685 4595 1690
rect 4555 1680 4595 1685
rect 4795 1685 4800 1690
rect 4830 1685 4835 1715
rect 4795 1680 4835 1685
rect 2150 1675 2190 1680
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4795 1595 4835 1600
rect 4795 1565 4800 1595
rect 4830 1590 4835 1595
rect 5390 1595 5430 1600
rect 5390 1590 5395 1595
rect 4830 1570 5395 1590
rect 4830 1565 4835 1570
rect 4795 1560 4835 1565
rect 5390 1565 5395 1570
rect 5425 1565 5430 1595
rect 5390 1560 5430 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4255 1545 4295 1550
rect 4255 1515 4260 1545
rect 4290 1540 4295 1545
rect 4375 1545 4415 1550
rect 4375 1540 4380 1545
rect 4290 1520 4380 1540
rect 4290 1515 4295 1520
rect 4255 1510 4295 1515
rect 4375 1515 4380 1520
rect 4410 1540 4415 1545
rect 4495 1545 4535 1550
rect 4495 1540 4500 1545
rect 4410 1520 4500 1540
rect 4410 1515 4415 1520
rect 4375 1510 4415 1515
rect 4495 1515 4500 1520
rect 4530 1540 4535 1545
rect 4615 1545 4655 1550
rect 4615 1540 4620 1545
rect 4530 1520 4620 1540
rect 4530 1515 4535 1520
rect 4495 1510 4535 1515
rect 4615 1515 4620 1520
rect 4650 1540 4655 1545
rect 4735 1545 4775 1550
rect 4735 1540 4740 1545
rect 4650 1520 4740 1540
rect 4650 1515 4655 1520
rect 4615 1510 4655 1515
rect 4735 1515 4740 1520
rect 4770 1540 4775 1545
rect 5125 1545 5165 1550
rect 5125 1540 5130 1545
rect 4770 1520 5130 1540
rect 4770 1515 4775 1520
rect 4735 1510 4775 1515
rect 5125 1515 5130 1520
rect 5160 1515 5165 1545
rect 5125 1510 5165 1515
rect 3375 1190 3415 1195
rect 3375 1160 3380 1190
rect 3410 1185 3415 1190
rect 4585 1190 4625 1195
rect 4585 1185 4590 1190
rect 3410 1165 4590 1185
rect 3410 1160 3415 1165
rect 3375 1155 3415 1160
rect 4585 1160 4590 1165
rect 4620 1185 4625 1190
rect 5445 1190 5485 1195
rect 5445 1185 5450 1190
rect 4620 1165 5450 1185
rect 4620 1160 4625 1165
rect 4585 1155 4625 1160
rect 5445 1160 5450 1165
rect 5480 1160 5485 1190
rect 5445 1155 5485 1160
rect 2940 1130 2980 1135
rect 2940 1100 2945 1130
rect 2975 1125 2980 1130
rect 3020 1130 3060 1135
rect 3020 1125 3025 1130
rect 2975 1105 3025 1125
rect 2975 1100 2980 1105
rect 2940 1095 2980 1100
rect 3020 1100 3025 1105
rect 3055 1125 3060 1130
rect 3100 1130 3140 1135
rect 3100 1125 3105 1130
rect 3055 1105 3105 1125
rect 3055 1100 3060 1105
rect 3020 1095 3060 1100
rect 3100 1100 3105 1105
rect 3135 1125 3140 1130
rect 3180 1130 3220 1135
rect 3180 1125 3185 1130
rect 3135 1105 3185 1125
rect 3135 1100 3140 1105
rect 3100 1095 3140 1100
rect 3180 1100 3185 1105
rect 3215 1125 3220 1130
rect 3260 1130 3300 1135
rect 3260 1125 3265 1130
rect 3215 1105 3265 1125
rect 3215 1100 3220 1105
rect 3180 1095 3220 1100
rect 3260 1100 3265 1105
rect 3295 1125 3300 1130
rect 3340 1130 3380 1135
rect 3340 1125 3345 1130
rect 3295 1105 3345 1125
rect 3295 1100 3300 1105
rect 3260 1095 3300 1100
rect 3340 1100 3345 1105
rect 3375 1125 3380 1130
rect 3420 1130 3460 1135
rect 3420 1125 3425 1130
rect 3375 1105 3425 1125
rect 3375 1100 3380 1105
rect 3340 1095 3380 1100
rect 3420 1100 3425 1105
rect 3455 1125 3460 1130
rect 3500 1130 3540 1135
rect 3500 1125 3505 1130
rect 3455 1105 3505 1125
rect 3455 1100 3460 1105
rect 3420 1095 3460 1100
rect 3500 1100 3505 1105
rect 3535 1125 3540 1130
rect 3580 1130 3620 1135
rect 3580 1125 3585 1130
rect 3535 1105 3585 1125
rect 3535 1100 3540 1105
rect 3500 1095 3540 1100
rect 3580 1100 3585 1105
rect 3615 1125 3620 1130
rect 3660 1130 3700 1135
rect 3660 1125 3665 1130
rect 3615 1105 3665 1125
rect 3615 1100 3620 1105
rect 3580 1095 3620 1100
rect 3660 1100 3665 1105
rect 3695 1125 3700 1130
rect 3740 1130 3780 1135
rect 3740 1125 3745 1130
rect 3695 1105 3745 1125
rect 3695 1100 3700 1105
rect 3660 1095 3700 1100
rect 3740 1100 3745 1105
rect 3775 1125 3780 1130
rect 3820 1130 3860 1135
rect 3820 1125 3825 1130
rect 3775 1105 3825 1125
rect 3775 1100 3780 1105
rect 3740 1095 3780 1100
rect 3820 1100 3825 1105
rect 3855 1125 3860 1130
rect 3900 1130 3940 1135
rect 3900 1125 3905 1130
rect 3855 1105 3905 1125
rect 3855 1100 3860 1105
rect 3820 1095 3860 1100
rect 3900 1100 3905 1105
rect 3935 1100 3940 1130
rect 3900 1095 3940 1100
rect 3980 1130 4020 1135
rect 3980 1100 3985 1130
rect 4015 1125 4020 1130
rect 4060 1130 4100 1135
rect 4060 1125 4065 1130
rect 4015 1105 4065 1125
rect 4015 1100 4020 1105
rect 3980 1095 4020 1100
rect 4060 1100 4065 1105
rect 4095 1125 4100 1130
rect 4140 1130 4180 1135
rect 4140 1125 4145 1130
rect 4095 1105 4145 1125
rect 4095 1100 4100 1105
rect 4060 1095 4100 1100
rect 4140 1100 4145 1105
rect 4175 1125 4180 1130
rect 4220 1130 4260 1135
rect 4220 1125 4225 1130
rect 4175 1105 4225 1125
rect 4175 1100 4180 1105
rect 4140 1095 4180 1100
rect 4220 1100 4225 1105
rect 4255 1125 4260 1130
rect 4300 1130 4340 1135
rect 4300 1125 4305 1130
rect 4255 1105 4305 1125
rect 4255 1100 4260 1105
rect 4220 1095 4260 1100
rect 4300 1100 4305 1105
rect 4335 1125 4340 1130
rect 4380 1130 4420 1135
rect 4380 1125 4385 1130
rect 4335 1105 4385 1125
rect 4335 1100 4340 1105
rect 4300 1095 4340 1100
rect 4380 1100 4385 1105
rect 4415 1125 4420 1130
rect 4460 1130 4500 1135
rect 4460 1125 4465 1130
rect 4415 1105 4465 1125
rect 4415 1100 4420 1105
rect 4380 1095 4420 1100
rect 4460 1100 4465 1105
rect 4495 1125 4500 1130
rect 4540 1130 4580 1135
rect 4540 1125 4545 1130
rect 4495 1105 4545 1125
rect 4495 1100 4500 1105
rect 4460 1095 4500 1100
rect 4540 1100 4545 1105
rect 4575 1125 4580 1130
rect 4620 1130 4660 1135
rect 4620 1125 4625 1130
rect 4575 1105 4625 1125
rect 4575 1100 4580 1105
rect 4540 1095 4580 1100
rect 4620 1100 4625 1105
rect 4655 1125 4660 1130
rect 4700 1130 4740 1135
rect 4700 1125 4705 1130
rect 4655 1105 4705 1125
rect 4655 1100 4660 1105
rect 4620 1095 4660 1100
rect 4700 1100 4705 1105
rect 4735 1125 4740 1130
rect 4780 1130 4820 1135
rect 4780 1125 4785 1130
rect 4735 1105 4785 1125
rect 4735 1100 4740 1105
rect 4700 1095 4740 1100
rect 4780 1100 4785 1105
rect 4815 1125 4820 1130
rect 4860 1130 4900 1135
rect 4860 1125 4865 1130
rect 4815 1105 4865 1125
rect 4815 1100 4820 1105
rect 4780 1095 4820 1100
rect 4860 1100 4865 1105
rect 4895 1125 4900 1130
rect 4940 1130 4980 1135
rect 4940 1125 4945 1130
rect 4895 1105 4945 1125
rect 4895 1100 4900 1105
rect 4860 1095 4900 1100
rect 4940 1100 4945 1105
rect 4975 1100 4980 1130
rect 4940 1095 4980 1100
rect 2620 1045 2660 1050
rect 2175 1030 2215 1035
rect 2175 1000 2180 1030
rect 2210 1025 2215 1030
rect 2425 1030 2465 1035
rect 2425 1025 2430 1030
rect 2210 1005 2430 1025
rect 2210 1000 2215 1005
rect 2175 995 2215 1000
rect 2425 1000 2430 1005
rect 2460 1000 2465 1030
rect 2620 1015 2625 1045
rect 2655 1040 2660 1045
rect 2900 1045 2940 1050
rect 2900 1040 2905 1045
rect 2655 1020 2905 1040
rect 2655 1015 2660 1020
rect 2620 1010 2660 1015
rect 2900 1015 2905 1020
rect 2935 1015 2940 1045
rect 2900 1010 2940 1015
rect 5055 1045 5095 1050
rect 5055 1015 5060 1045
rect 5090 1040 5095 1045
rect 5445 1045 5485 1050
rect 5445 1040 5450 1045
rect 5090 1020 5450 1040
rect 5090 1015 5095 1020
rect 5055 1010 5095 1015
rect 5445 1015 5450 1020
rect 5480 1015 5485 1045
rect 5445 1010 5485 1015
rect 2425 995 2465 1000
rect 2990 935 3030 940
rect 2990 905 2995 935
rect 3025 930 3030 935
rect 3170 935 3210 940
rect 3170 930 3175 935
rect 3025 910 3175 930
rect 3025 905 3030 910
rect 2990 900 3030 905
rect 3170 905 3175 910
rect 3205 930 3210 935
rect 3350 935 3390 940
rect 3350 930 3355 935
rect 3205 910 3355 930
rect 3205 905 3210 910
rect 3170 900 3210 905
rect 3350 905 3355 910
rect 3385 930 3390 935
rect 3530 935 3570 940
rect 3530 930 3535 935
rect 3385 910 3535 930
rect 3385 905 3390 910
rect 3350 900 3390 905
rect 3530 905 3535 910
rect 3565 930 3570 935
rect 3710 935 3750 940
rect 3710 930 3715 935
rect 3565 910 3715 930
rect 3565 905 3570 910
rect 3530 900 3570 905
rect 3710 905 3715 910
rect 3745 930 3750 935
rect 3890 935 3930 940
rect 3890 930 3895 935
rect 3745 910 3895 930
rect 3745 905 3750 910
rect 3710 900 3750 905
rect 3890 905 3895 910
rect 3925 930 3930 935
rect 4070 935 4110 940
rect 4070 930 4075 935
rect 3925 910 4075 930
rect 3925 905 3930 910
rect 3890 900 3930 905
rect 4070 905 4075 910
rect 4105 930 4110 935
rect 4250 935 4290 940
rect 4250 930 4255 935
rect 4105 910 4255 930
rect 4105 905 4110 910
rect 4070 900 4110 905
rect 4250 905 4255 910
rect 4285 930 4290 935
rect 4430 935 4470 940
rect 4430 930 4435 935
rect 4285 910 4435 930
rect 4285 905 4290 910
rect 4250 900 4290 905
rect 4430 905 4435 910
rect 4465 930 4470 935
rect 4610 935 4650 940
rect 4610 930 4615 935
rect 4465 910 4615 930
rect 4465 905 4470 910
rect 4430 900 4470 905
rect 4610 905 4615 910
rect 4645 930 4650 935
rect 4790 935 4830 940
rect 4790 930 4795 935
rect 4645 910 4795 930
rect 4645 905 4650 910
rect 4610 900 4650 905
rect 4790 905 4795 910
rect 4825 930 4830 935
rect 4970 935 5010 940
rect 4970 930 4975 935
rect 4825 910 4975 930
rect 4825 905 4830 910
rect 4790 900 4830 905
rect 4970 905 4975 910
rect 5005 930 5010 935
rect 5445 935 5485 940
rect 5445 930 5450 935
rect 5005 910 5450 930
rect 5005 905 5010 910
rect 4970 900 5010 905
rect 5445 905 5450 910
rect 5480 905 5485 935
rect 5445 900 5485 905
rect 3620 765 3660 770
rect 2520 750 2560 755
rect 2520 720 2525 750
rect 2555 745 2560 750
rect 3080 750 3120 755
rect 3080 745 3085 750
rect 2555 725 3085 745
rect 2555 720 2560 725
rect 2520 715 2560 720
rect 3080 720 3085 725
rect 3115 720 3120 750
rect 3620 735 3625 765
rect 3655 760 3660 765
rect 3980 765 4020 770
rect 3980 760 3985 765
rect 3655 740 3985 760
rect 3655 735 3660 740
rect 3620 730 3660 735
rect 3980 735 3985 740
rect 4015 760 4020 765
rect 4340 765 4380 770
rect 4340 760 4345 765
rect 4015 740 4345 760
rect 4015 735 4020 740
rect 3980 730 4020 735
rect 4340 735 4345 740
rect 4375 735 4380 765
rect 4340 730 4380 735
rect 4520 765 4560 770
rect 4520 735 4525 765
rect 4555 760 4560 765
rect 4700 765 4740 770
rect 4700 760 4705 765
rect 4555 740 4705 760
rect 4555 735 4560 740
rect 4520 730 4560 735
rect 4700 735 4705 740
rect 4735 760 4740 765
rect 4880 765 4920 770
rect 4880 760 4885 765
rect 4735 740 4885 760
rect 4735 735 4740 740
rect 4700 730 4740 735
rect 4880 735 4885 740
rect 4915 735 4920 765
rect 4880 730 4920 735
rect 3080 715 3120 720
rect 3440 710 3480 715
rect 3440 680 3445 710
rect 3475 705 3480 710
rect 3800 710 3840 715
rect 3800 705 3805 710
rect 3475 685 3805 705
rect 3475 680 3480 685
rect 3440 675 3480 680
rect 3800 680 3805 685
rect 3835 705 3840 710
rect 4160 710 4200 715
rect 4160 705 4165 710
rect 3835 685 4165 705
rect 3835 680 3840 685
rect 3800 675 3840 680
rect 4160 680 4165 685
rect 4195 680 4200 710
rect 4160 675 4200 680
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
<< via2 >>
rect -190 4960 -160 4990
rect 5535 4960 5565 4990
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5535 3415 5565 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect 5535 2780 5565 2810
rect -105 1690 -75 1720
rect 5450 1160 5480 1190
rect 5450 1015 5480 1045
rect 5450 905 5480 935
rect -190 545 -160 575
<< metal3 >>
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5525 4995 5575 5000
rect 5525 4955 5530 4995
rect 5570 4955 5575 4995
rect 5525 4950 5575 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5440 4910 5490 4915
rect 5440 4870 5445 4910
rect 5485 4870 5490 4910
rect 5440 4865 5490 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 1720 -70 2970
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5445 1190 5485 4865
rect 5445 1160 5450 1190
rect 5480 1160 5485 1190
rect 5445 1045 5485 1160
rect 5445 1015 5450 1045
rect 5480 1015 5485 1045
rect 5445 935 5485 1015
rect 5445 905 5450 935
rect 5480 905 5485 935
rect 5445 665 5485 905
rect 5530 3445 5570 4950
rect 5530 3415 5535 3445
rect 5565 3415 5570 3445
rect 5530 2810 5570 3415
rect 5530 2780 5535 2810
rect 5565 2780 5570 2810
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5440 660 5490 665
rect 5440 620 5445 660
rect 5485 620 5490 660
rect 5440 615 5490 620
rect 5530 585 5570 2780
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5525 580 5575 585
rect 5525 540 5530 580
rect 5570 540 5575 580
rect 5525 535 5575 540
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5530 4990 5570 4995
rect 5530 4960 5535 4990
rect 5535 4960 5565 4990
rect 5565 4960 5570 4990
rect 5530 4955 5570 4960
rect -110 4870 -70 4910
rect 5445 4870 5485 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect -110 620 -70 660
rect 5445 620 5485 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5530 540 5570 580
<< mimcap >>
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
<< mimcapcontact >>
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 5140 3675 5180 3715
<< metal4 >>
rect -200 4995 5575 5000
rect -200 4955 -195 4995
rect -155 4955 5530 4995
rect 5570 4955 5575 4995
rect -200 4950 5575 4955
rect -115 4910 5490 4915
rect -115 4870 -110 4910
rect -70 4870 5445 4910
rect 5485 4870 5490 4910
rect -115 4865 5490 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -115 660 5490 665
rect -115 620 -110 660
rect -70 620 5445 660
rect 5485 620 5490 660
rect -115 615 5490 620
rect -200 580 5575 585
rect -200 540 -195 580
rect -155 540 5530 580
rect 5570 540 5575 580
rect -200 535 5575 540
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal3 5570 4400 5570 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5485 4175 5485 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 3270 350 3270 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3820 295 3820 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4010 350 4010 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4720 295 4720 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal2 6060 3075 6060 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6080 3020 6080 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6060 2955 6060 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6080 1745 6080 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
<< end >>
