magic
tech sky130A
timestamp 1737793922
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 0 0 1 0
box -19 -24 157 296
<< end >>
