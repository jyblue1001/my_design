* PEX produced on Mon Sep  1 11:23:19 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from pll_bgr_magic.ext - technology: sky130A

.subckt pll_bgr_magic V_OSC VDDA GNDA F_REF
X0 GNDA.t268 GNDA.t266 GNDA.t268 GNDA.t267 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X1 a_5970_4630.t5 V_CONT.t8 a_6200_5250.t1 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 GNDA.t92 a_6200_5250.t4 a_6200_5250.t5 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 GNDA.t282 pfd_8_0.F_b.t3 pfd_8_0.F.t2 GNDA.t281 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X4 a_6330_n1530.t2 VCO_FD_magic_0.div120_2_0.div4.t2 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 bgr_0.V_TOP.t13 bgr_0.1st_Vout_1.t11 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X6 pfd_8_0.QB_b.t2 pfd_8_0.QB.t3 a_n30_630.t1 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X7 VCO_FD_magic_0.vco2_3_0.V9.t1 V_OSC.t2 VCO_FD_magic_0.vco2_3_0.V6.t1 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X8 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 bgr_0.Vin+.t5 bgr_0.V_TOP.t14 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X10 BGR_CURRENT_OUT.t14 bgr_0.V2.t10 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X11 BGR_CURRENT_OUT.t13 bgr_0.V2.t11 VDDA.t413 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X12 bgr_0.V2.t9 VDDA.t335 VDDA.t337 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X13 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 VCO_FD_magic_0.div120_2_0.div24.t3 GNDA.t323 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 GNDA.t34 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 VDDA.t257 pfd_8_0.Reset.t2 a_1390_630.t1 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X17 bgr_0.V_p_2.t9 bgr_0.V1.t7 a_n1450_5080.t14 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X18 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 pfd_8_0.E.t1 pfd_8_0.E_b.t3 a_870_1390.t1 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X20 GNDA.t98 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X21 VDDA.t6 VCO_FD_magic_0.div120_2_0.div2.t2 a_7630_n1530.t2 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 pfd_8_0.UP_b.t2 pfd_8_0.UP.t2 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X23 pfd_8_0.UP_input.t3 pfd_8_0.UP_b.t0 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X24 GNDA.t221 GNDA.t260 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X25 VDDA.t27 VCO_FD_magic_0.vco2_3_0.V1.t3 VCO_FD_magic_0.vco2_3_0.V4.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X26 GNDA.t68 pfd_8_0.QB.t4 pfd_8_0.QB_b.t1 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X27 VDDA.t42 pfd_8_0.opamp_out.t10 opamp_cell_4_0.VIN+.t3 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X28 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.n_left.t6 VDDA.t230 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X29 GNDA.t221 GNDA.t265 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X30 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 pfd_8_0.opamp_out.t7 opamp_cell_4_0.n_right.t5 VDDA.t218 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X32 opamp_cell_4_0.n_right.t3 opamp_cell_4_0.VIN+.t6 a_6320_5840.t9 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X33 GNDA.t190 VCO_FD_magic_0.div120_2_0.div8.t2 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X34 pfd_8_0.opamp_out.t9 a_6490_4630.t5 GNDA.t316 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 bgr_0.1st_Vout_1.t9 bgr_0.V_mir1.t17 VDDA.t359 VDDA.t358 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X36 VDDA.t262 GNDA.t328 VCO_FD_magic_0.vco2_3_0.V4.t2 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X37 GNDA.t302 pfd_8_0.Reset.t3 pfd_8_0.F_b.t2 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X38 a_3280_11518.t1 bgr_0.Vin-.t1 GNDA.t187 sky130_fd_pr__res_xhigh_po_0p35 l=6
X39 bgr_0.V_TOP.t15 VDDA.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VDDA.t54 a_6330_n1530.t3 VCO_FD_magic_0.div120_2_0.div8.t1 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X41 bgr_0.V_TOP.t16 VDDA.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X43 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 GNDA.t145 BGR_CURRENT_OUT.t3 BGR_CURRENT_OUT.t4 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X45 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 VCO_FD_magic_0.div120_2_0.div4.t3 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 VDDA.t18 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t7 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X47 VDDA.t8 a_n1450_5080.t10 a_n1450_5080.t11 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X48 BGR_CURRENT_OUT.t12 bgr_0.V2.t12 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X49 VDDA.t73 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 a_7630_n1530.t3 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X51 VDDA.t200 bgr_0.1st_Vout_2.t13 bgr_0.V2.t6 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X52 bgr_0.1st_Vout_1.t8 bgr_0.V_mir1.t18 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 bgr_0.V_TOP.t17 VDDA.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 bgr_0.cap_res2.t0 bgr_0.V2.t0 GNDA.t76 sky130_fd_pr__res_high_po_0p35 l=2.05
X55 pfd_8_0.E.t0 pfd_8_0.QA_b.t3 GNDA.t194 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X56 bgr_0.Vin-.t7 bgr_0.V_TOP.t18 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X57 bgr_0.V_TOP.t7 VDDA.t332 VDDA.t334 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X58 VDDA.t175 bgr_0.V2.t13 bgr_0.V_CUR_REF_REG.t9 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X59 VDDA.t60 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t12 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X60 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t13 bgr_0.V_p_2.t4 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X61 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VDDA.t374 opamp_cell_4_0.p_bias.t9 a_5970_4630.t11 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X63 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 a_6200_5250.t0 V_CONT.t9 a_5970_4630.t4 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X65 a_6200_5250.t3 a_6200_5250.t2 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X66 VDDA.t108 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X67 VDDA.t372 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X68 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 VDDA.t331 VDDA.t328 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X70 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X71 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 VCO_FD_magic_0.div120_2_0.div8.t3 GNDA.t106 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X72 bgr_0.1st_Vout_2.t5 bgr_0.V_CUR_REF_REG.t14 bgr_0.V_p_2.t2 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X73 a_8930_n1530.t0 V_OSC.t3 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X74 VDDA.t327 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X75 a_n30_630.t0 F_VCO.t2 VDDA.t82 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X76 VDDA.t422 pfd_8_0.UP_input.t4 V_CONT.t7 VDDA.t421 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X77 a_6220_5810.t8 a_6220_5810.t7 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X78 VDDA.t65 bgr_0.1st_Vout_1.t17 bgr_0.V_TOP.t11 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 VDDA.t133 bgr_0.V_TOP.t19 a_n1130_7570.t5 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X80 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 VCO_FD_magic_0.div120_2_0.div24.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X82 GNDA.t87 F_VCO.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X83 GNDA.t290 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X84 VDDA.t386 a_2200_180.t2 a_1870_180.t1 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X85 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 a_6330_n1530.t4 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X86 GNDA.t176 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 VCO_FD_magic_0.div120_2_0.div8.t0 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X87 bgr_0.V_TOP.t20 VDDA.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 a_6320_5840.t2 a_6220_5810.t9 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X89 pfd_8_0.QA_b.t2 F_REF.t0 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X90 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X91 BGR_CURRENT_OUT.t11 bgr_0.V2.t14 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X92 a_n1450_5080.t16 bgr_0.V1.t8 bgr_0.V_p_2.t8 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X93 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X94 pfd_8_0.QB_b.t0 F_VCO.t4 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X95 a_5970_4630.t3 opamp_cell_4_0.p_bias.t10 VDDA.t216 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X96 VDDA.t240 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t6 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X97 GNDA.t182 VDDA.t423 bgr_0.V_p_2.t10 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X98 a_490_630.t1 pfd_8_0.QB_b.t3 pfd_8_0.QB.t2 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X99 VDDA.t365 pfd_8_0.Reset.t4 a_1390_1390.t1 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X100 BGR_CURRENT_OUT.t2 BGR_CURRENT_OUT.t1 GNDA.t157 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X101 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VDDA.t324 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X103 pfd_8_0.opamp_out.t11 a_9360_3514.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X104 V_CONT.t6 loop_filter_2_0.R1_C1.t1 GNDA.t298 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X105 GNDA.t264 GNDA.t261 GNDA.t263 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X106 GNDA.t259 GNDA.t257 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X107 a_2530_180.t1 a_2350_1390.t2 VDDA.t248 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X108 GNDA.t212 a_n1490_9910.t1 GNDA.t211 sky130_fd_pr__res_xhigh_po_0p35 l=6
X109 GNDA.t306 a_2200_180.t3 a_1870_180.t0 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X110 opamp_cell_4_0.p_bias.t5 opamp_cell_4_0.p_bias.t4 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X111 GNDA.t205 a_7630_n1530.t4 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X112 VCO_FD_magic_0.vco2_3_0.V1.t2 V_CONT.t10 GNDA.t147 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X113 VDDA.t104 bgr_0.V_TOP.t21 bgr_0.Vin-.t6 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X114 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.QB.t5 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X115 VDDA.t355 bgr_0.V_mir1.t20 bgr_0.1st_Vout_1.t7 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X116 V_OSC.t1 VCO_FD_magic_0.vco2_3_0.V8.t2 VCO_FD_magic_0.vco2_3_0.V3.t0 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X117 pfd_8_0.QB.t1 pfd_8_0.QB_b.t4 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X118 V_CONT.t1 pfd_8_0.UP_input.t5 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X119 bgr_0.V_TOP.t22 VDDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 GNDA.t46 VCO_FD_magic_0.div120_2_0.div24.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X121 VDDA.t320 VDDA.t318 VDDA.t320 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X122 bgr_0.V_mir1.t0 bgr_0.Vin-.t8 bgr_0.V_p_1.t4 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X123 VDDA.t317 VDDA.t315 bgr_0.V_TOP.t6 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X124 bgr_0.V_CUR_REF_REG.t8 bgr_0.V2.t15 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X125 bgr_0.V2.t7 VDDA.t424 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X126 GNDA.t256 GNDA.t253 GNDA.t255 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X127 GNDA.t252 GNDA.t249 GNDA.t251 GNDA.t250 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X128 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 GNDA.t135 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X129 bgr_0.V1.t2 VDDA.t312 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X130 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 a_8930_n1530.t3 GNDA.t320 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X131 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X132 bgr_0.1st_Vout_2.t9 a_n1450_5080.t17 VDDA.t242 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X133 GNDA.t180 VDDA.t425 VCO_FD_magic_0.vco2_3_0.V3.t2 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X134 a_n2040_11368.t1 a_n1920_10290.t0 GNDA.t210 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X135 GNDA.t325 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X136 bgr_0.V2.t5 bgr_0.1st_Vout_2.t16 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 pfd_8_0.opamp_out.t12 a_9360_6440.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X138 VDDA.t361 bgr_0.V_mir1.t21 bgr_0.1st_Vout_1.t10 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X139 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t6 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X140 GNDA.t137 F_VCO.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X141 BGR_CURRENT_OUT.t16 VDDA.t309 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X142 pfd_8_0.E_b.t1 pfd_8_0.E.t3 GNDA.t276 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X143 GNDA.t248 GNDA.t245 GNDA.t247 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X144 pfd_8_0.UP_input.t1 pfd_8_0.UP.t3 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X145 GNDA.t85 a_6220_5810.t10 a_6320_5840.t1 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X146 bgr_0.1st_Vout_1.t5 bgr_0.V_mir1.t22 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X147 pfd_8_0.DOWN_b.t0 GNDA.t329 pfd_8_0.DOWN_PFD_b.t2 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X148 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 VDDA.t226 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X149 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 GNDA.t314 bgr_0.V_CUR_REF_REG.t12 GNDA.t313 sky130_fd_pr__res_xhigh_po_0p35 l=1
X152 GNDA.t164 a_6220_5810.t5 a_6220_5810.t6 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X153 GNDA.t244 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X154 bgr_0.1st_Vout_1.t3 bgr_0.Vin+.t6 bgr_0.V_p_1.t9 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X155 a_3280_11518.t0 a_3160_9910.t0 GNDA.t59 sky130_fd_pr__res_xhigh_po_0p35 l=6
X156 a_5970_4630.t10 a_5970_4630.t9 a_5970_4630.t10 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X157 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 GNDA.t240 GNDA.t238 GNDA.t240 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X159 VDDA.t246 pfd_8_0.UP_input.t6 V_CONT.t4 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X160 bgr_0.V_CUR_REF_REG.t7 bgr_0.V2.t16 VDDA.t382 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X161 bgr_0.V_CUR_REF_REG.t6 bgr_0.V2.t17 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X162 pfd_8_0.DOWN_b.t1 VDDA.t426 pfd_8_0.DOWN_PFD_b.t3 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X163 bgr_0.V_TOP.t23 VDDA.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 GNDA.t330 loop_filter_2_0.R1_C1.t0 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X165 VDDA.t12 VCO_FD_magic_0.div120_2_0.div4.t4 a_6330_n1530.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X166 GNDA.t27 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1.t1 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X167 VDDA.t308 VDDA.t306 VDDA.t308 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X168 bgr_0.V_TOP.t24 VDDA.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t15 bgr_0.1st_Vout_2.t0 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X170 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t2 VDDA.t416 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X171 GNDA.t237 GNDA.t235 GNDA.t237 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X172 bgr_0.V_mir1.t16 bgr_0.V_mir1.t15 VDDA.t363 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X173 bgr_0.V_p_2.t3 bgr_0.V_CUR_REF_REG.t16 bgr_0.1st_Vout_2.t6 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X174 bgr_0.V_CUR_REF_REG.t11 VDDA.t303 VDDA.t305 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X175 bgr_0.V_TOP.t25 VDDA.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 bgr_0.V_TOP.t26 VDDA.t251 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 GNDA.t8 VCO_FD_magic_0.div120_2_0.div24.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X178 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 GNDA.t56 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X180 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VDDA.t253 bgr_0.V_TOP.t27 bgr_0.Vin+.t4 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X182 VDDA.t16 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X183 GNDA.t148 V_CONT.t11 VCO_FD_magic_0.vco2_3_0.V7.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X184 VDDA.t205 pfd_8_0.QA.t3 pfd_8_0.before_Reset.t1 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X185 a_2350_1390.t1 pfd_8_0.before_Reset.t3 GNDA.t312 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X186 GNDA.t75 VDDA.t427 VCO_FD_magic_0.vco2_3_0.V5.t2 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X187 VDDA.t237 VCO_FD_magic_0.vco2_3_0.V1.t4 VCO_FD_magic_0.vco2_3_0.V2.t1 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X188 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t4 VDDA.t113 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X189 bgr_0.V_mir1.t14 bgr_0.V_mir1.t13 VDDA.t353 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X190 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t3 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X191 bgr_0.1st_Vout_2.t1 a_n1450_5080.t18 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X192 opamp_cell_4_0.VIN+.t2 pfd_8_0.opamp_out.t13 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X193 VDDA.t1 opamp_cell_4_0.n_right.t6 pfd_8_0.opamp_out.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X194 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VDDA.t302 VDDA.t300 BGR_CURRENT_OUT.t15 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X196 GNDA.t66 a_6490_4630.t6 pfd_8_0.opamp_out.t1 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X197 a_n1610_11518.t0 bgr_0.Vin+.t0 GNDA.t114 sky130_fd_pr__res_xhigh_po_0p35 l=6
X198 bgr_0.V_p_1.t3 bgr_0.Vin-.t9 bgr_0.V_mir1.t1 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X199 VDDA.t167 pfd_8_0.E.t4 a_490_1390.t1 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X200 VDDA.t405 bgr_0.1st_Vout_2.t20 bgr_0.V2.t4 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X201 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div8.t4 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X202 V_CONT.t2 pfd_8_0.UP_input.t7 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X203 a_8930_n1530.t2 V_OSC.t4 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X204 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VDDA.t261 GNDA.t331 VCO_FD_magic_0.vco2_3_0.V2.t2 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X206 VDDA.t212 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 F_VCO.t1 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X207 VDDA.t228 a_n1450_5080.t19 bgr_0.1st_Vout_2.t8 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X208 VDDA.t48 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X209 GNDA.t100 pfd_8_0.QA.t5 pfd_8_0.QA_b.t1 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X210 bgr_0.V_mir1.t12 bgr_0.V_mir1.t11 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X211 bgr_0.V_p_1.t2 bgr_0.Vin-.t10 bgr_0.V_mir1.t3 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X212 GNDA.t300 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 VCO_FD_magic_0.div120_2_0.div24.t2 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X213 bgr_0.V_TOP.t28 VDDA.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 bgr_0.V_CUR_REF_REG.t5 bgr_0.V2.t18 VDDA.t407 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X215 VCO_FD_magic_0.vco2_3_0.V9.t0 V_OSC.t5 VCO_FD_magic_0.vco2_3_0.V7.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X216 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 F_VCO.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X217 a_7630_n1530.t0 VCO_FD_magic_0.div120_2_0.div2.t3 GNDA.t278 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X218 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X219 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN_b.t4 BGR_CURRENT_OUT.t0 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X221 bgr_0.V_TOP.t29 VDDA.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VDDA.t36 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X223 a_1910_2010.t1 pfd_8_0.QB.t7 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X224 a_6320_5840.t11 V_CONT.t12 opamp_cell_4_0.n_left.t5 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X225 VCO_FD_magic_0.vco2_3_0.V8.t0 VCO_FD_magic_0.vco2_3_0.V9.t2 VCO_FD_magic_0.vco2_3_0.V4.t1 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X226 bgr_0.V_p_1.t8 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t4 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X227 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 GNDA.t170 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X229 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 a_8930_n1530.t4 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X230 GNDA.t58 VCO_FD_magic_0.div120_2_0.div24.t7 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X231 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 GNDA.t119 VCO_FD_magic_0.div120_2_0.div2.t4 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X233 VDDA.t409 bgr_0.V2.t19 BGR_CURRENT_OUT.t10 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X234 GNDA.t207 VDDA.t428 bgr_0.V_TOP.t3 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X235 VDDA.t80 a_n1450_5080.t20 bgr_0.1st_Vout_2.t2 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X236 VDDA.t142 bgr_0.V_TOP.t30 a_n1130_7570.t4 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X237 pfd_8_0.UP_input.t0 pfd_8_0.UP.t4 pfd_8_0.opamp_out.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X238 bgr_0.V_TOP.t31 VDDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 pfd_8_0.QA.t0 pfd_8_0.QA_b.t4 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X240 bgr_0.Vin-.t5 bgr_0.V_TOP.t32 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X241 bgr_0.V_TOP.t10 bgr_0.1st_Vout_1.t25 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X242 VDDA.t159 a_8930_n1530.t5 VCO_FD_magic_0.div120_2_0.div2.t0 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X243 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN.t3 BGR_CURRENT_OUT.t17 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X244 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN.t2 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X245 a_n1450_5080.t13 bgr_0.V1.t9 bgr_0.V_p_2.t7 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X246 GNDA.t292 a_n1920_10290.t1 GNDA.t291 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X247 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X248 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 VCO_FD_magic_0.div120_2_0.div8.t5 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X249 a_870_630.t0 pfd_8_0.QB_b.t5 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X250 VDDA.t349 bgr_0.V_mir1.t9 bgr_0.V_mir1.t10 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X251 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div24.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X252 VDDA.t163 a_2530_180.t2 a_2200_180.t1 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X253 GNDA.t140 a_6330_n1530.t5 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X254 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 a_6330_n1530.t6 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X255 bgr_0.V_CUR_REF_REG.t4 bgr_0.V2.t20 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X256 a_5970_4630.t8 a_5970_4630.t6 a_5970_4630.t7 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X257 VDDA.t341 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X258 GNDA.t234 GNDA.t231 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X259 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 bgr_0.V1.t6 bgr_0.V_TOP.t33 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X261 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 pfd_8_0.opamp_out.t8 opamp_cell_4_0.n_right.t7 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X263 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 F_VCO.t7 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X264 pfd_8_0.opamp_out.t3 a_6490_4630.t7 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X265 GNDA.t221 GNDA.t230 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X266 VDDA.t394 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X267 VDDA.t351 bgr_0.V_mir1.t7 bgr_0.V_mir1.t8 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 VDDA.t93 a_n1450_5080.t8 a_n1450_5080.t9 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X269 pfd_8_0.F.t0 pfd_8_0.QB_b.t6 GNDA.t133 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X270 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 a_7630_n1530.t5 GNDA.t152 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X271 GNDA.t54 a_2530_180.t3 a_2200_180.t0 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X272 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t5 GNDA.t327 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X273 GNDA.t221 GNDA.t229 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X274 VDDA.t171 bgr_0.V2.t21 BGR_CURRENT_OUT.t9 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X275 bgr_0.V2.t3 bgr_0.1st_Vout_2.t24 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X276 bgr_0.V_TOP.t34 VDDA.t187 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 GNDA.t200 pfd_8_0.E_b.t4 pfd_8_0.E.t2 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X278 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 VCO_FD_magic_0.div120_2_0.div24.t9 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X279 VDDA.t299 VDDA.t296 VDDA.t298 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X280 a_n2040_11368.t0 bgr_0.V1.t0 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X281 a_870_1390.t0 pfd_8_0.QA_b.t5 VDDA.t208 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X282 pfd_8_0.UP_b.t1 pfd_8_0.UP.t5 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X283 bgr_0.Vin-.t2 a_n1130_7570.t6 bgr_0.V_TOP.t2 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X284 bgr_0.V2.t2 bgr_0.1st_Vout_2.t25 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X285 a_1390_630.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t0 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X286 opamp_cell_4_0.p_bias.t3 opamp_cell_4_0.p_bias.t2 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X287 GNDA.t221 GNDA.t228 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X288 bgr_0.1st_Vout_1.t0 bgr_0.Vin+.t8 bgr_0.V_p_1.t7 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X289 VDDA.t345 bgr_0.V_mir1.t5 bgr_0.V_mir1.t6 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X290 opamp_cell_4_0.p_bias.t8 a_6220_5810.t0 GNDA.t111 sky130_fd_pr__res_xhigh_po_5p73 l=1
X291 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 GNDA.t160 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X293 VDDA.t52 VCO_FD_magic_0.vco2_3_0.V1.t5 VCO_FD_magic_0.vco2_3_0.V6.t0 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X294 bgr_0.V_TOP.t35 VDDA.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 GNDA.t318 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 VCO_FD_magic_0.div120_2_0.div2.t1 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X296 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X297 bgr_0.Vin+.t3 bgr_0.V_TOP.t36 VDDA.t418 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X298 GNDA.t332 V_CONT.t5 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X299 opamp_cell_4_0.n_left.t1 opamp_cell_4_0.n_left.t0 VDDA.t259 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X300 GNDA.t150 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 F_VCO.t0 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X301 VDDA.t420 bgr_0.V_TOP.t37 bgr_0.Vin-.t4 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X302 opamp_cell_4_0.n_left.t4 V_CONT.t13 a_6320_5840.t10 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X303 bgr_0.V_TOP.t38 VDDA.t366 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X305 a_5970_4630.t2 opamp_cell_4_0.p_bias.t11 VDDA.t151 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X306 VDDA.t181 bgr_0.1st_Vout_1.t28 bgr_0.V_TOP.t9 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 VDDA.t260 GNDA.t333 VCO_FD_magic_0.vco2_3_0.V6.t2 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X308 VDDA.t145 VCO_FD_magic_0.div120_2_0.div24.t10 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X309 bgr_0.V_mir1.t2 bgr_0.Vin-.t11 bgr_0.V_p_1.t1 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X310 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VDDA.t165 VCO_FD_magic_0.div120_2_0.div24.t11 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X312 pfd_8_0.F_b.t1 pfd_8_0.F.t4 GNDA.t272 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X313 VDDA.t99 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X314 VDDA.t364 pfd_8_0.F.t5 a_490_630.t0 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X315 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 a_n1610_11518.t1 a_n1490_9910.t0 GNDA.t162 sky130_fd_pr__res_xhigh_po_0p35 l=6
X317 VDDA.t295 VDDA.t293 VDDA.t295 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X318 VDDA.t292 VDDA.t290 bgr_0.V1.t1 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X319 GNDA.t221 GNDA.t227 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X320 a_9360_6440.t0 a_6490_4630.t0 GNDA.t153 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X321 a_n30_1390.t1 F_REF.t1 VDDA.t231 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X322 VDDA.t378 bgr_0.V2.t22 BGR_CURRENT_OUT.t8 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X323 bgr_0.V_p_2.t6 bgr_0.V1.t10 a_n1450_5080.t15 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X324 VDDA.t289 VDDA.t287 bgr_0.V_TOP.t5 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X325 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 GNDA.t226 GNDA.t224 GNDA.t226 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X327 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 GNDA.t94 a_6220_5810.t3 a_6220_5810.t4 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X329 VDDA.t286 VDDA.t283 VDDA.t285 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X330 VDDA.t67 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t2 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X331 GNDA.t126 a_6490_4630.t8 pfd_8_0.opamp_out.t4 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X332 GNDA.t270 pfd_8_0.F.t6 pfd_8_0.QB.t0 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X333 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_0.Vin+.t1 GNDA.t161 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X335 GNDA.t221 GNDA.t222 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X336 VCO_FD_magic_0.div120_2_0.div24.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X337 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 VCO_FD_magic_0.div120_2_0.div24.t12 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X338 VDDA.t78 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 VCO_FD_magic_0.div120_2_0.div24.t1 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X339 GNDA.t21 a_6220_5810.t11 a_6320_5840.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X340 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 GNDA.t295 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X341 VDDA.t282 VDDA.t280 bgr_0.V_CUR_REF_REG.t10 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X342 VDDA.t376 opamp_cell_4_0.p_bias.t12 a_5970_4630.t12 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X343 VDDA.t368 bgr_0.V_TOP.t39 bgr_0.Vin+.t2 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X344 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t30 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X345 a_7630_n1530.t1 VCO_FD_magic_0.div120_2_0.div2.t5 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X346 bgr_0.V_TOP.t40 VDDA.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 a_5970_4630.t0 opamp_cell_4_0.VIN+.t7 a_6490_4630.t2 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X348 a_n1450_5080.t7 a_n1450_5080.t6 VDDA.t244 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X349 GNDA.t274 a_6200_5250.t6 a_6490_4630.t4 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X350 bgr_0.V_p_1.t10 VDDA.t429 GNDA.t209 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X351 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X352 a_n1130_7570.t3 bgr_0.V_TOP.t41 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X353 VDDA.t370 a_n1450_5080.t21 bgr_0.1st_Vout_2.t10 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X354 bgr_0.V_TOP.t42 VDDA.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 opamp_cell_4_0.n_right.t4 a_9360_3514.t1 GNDA.t153 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X356 bgr_0.START_UP_NFET1.t1 a_n1130_7570.t0 a_n1130_7570.t1 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X357 VDDA.t380 bgr_0.V2.t23 BGR_CURRENT_OUT.t7 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X358 VDDA.t153 opamp_cell_4_0.p_bias.t0 opamp_cell_4_0.p_bias.t1 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X359 GNDA.t280 pfd_8_0.Reset.t5 pfd_8_0.E_b.t0 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X360 a_1390_1390.t0 pfd_8_0.E.t5 pfd_8_0.E_b.t2 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X361 a_6330_n1530.t0 VCO_FD_magic_0.div120_2_0.div4.t5 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X362 VDDA.t279 VDDA.t276 VDDA.t278 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X363 VDDA.t275 VDDA.t273 bgr_0.V2.t8 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X364 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 VDDA.t202 VCO_FD_magic_0.div120_2_0.div8.t6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X366 a_6320_5840.t7 a_6320_5840.t5 a_6320_5840.t6 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X367 VDDA.t415 V_OSC.t6 a_8930_n1530.t1 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X368 bgr_0.V_p_1.t6 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X369 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 a_2530_180.t0 a_2350_1390.t3 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X371 a_6320_5840.t12 a_6220_5810.t12 GNDA.t304 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X372 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X374 GNDA.t64 VCO_FD_magic_0.div120_2_0.div4.t6 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 GNDA.t184 pfd_8_0.DOWN_input.t4 V_CONT.t3 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X376 GNDA.t221 GNDA.t220 bgr_0.Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X377 a_n1130_7570.t2 bgr_0.V_TOP.t43 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X378 VDDA.t91 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X379 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VDDA.t272 VDDA.t270 VDDA.t272 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X381 bgr_0.V_p_1.t0 bgr_0.Vin-.t12 bgr_0.V_mir1.t4 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X382 VDDA.t396 bgr_0.V2.t24 bgr_0.V_CUR_REF_REG.t3 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X383 bgr_0.V_TOP.t0 a_n1130_7570.t7 bgr_0.Vin-.t0 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X384 a_6320_5840.t4 a_6320_5840.t3 a_6320_5840.t4 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X385 VDDA.t401 a_7630_n1530.t6 VCO_FD_magic_0.div120_2_0.div4.t1 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X386 a_6220_5810.t2 a_6220_5810.t1 GNDA.t83 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X387 VDDA.t97 a_n1450_5080.t4 a_n1450_5080.t5 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X388 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 VCO_FD_magic_0.div120_2_0.div24.t13 VDDA.t210 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X389 GNDA.t307 V_CONT.t14 VCO_FD_magic_0.vco2_3_0.V3.t1 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X390 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 VCO_FD_magic_0.div120_2_0.div2.t6 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X391 GNDA.t166 BGR_CURRENT_OUT.t18 opamp_cell_4_0.VIN+.t5 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X392 a_n1450_5080.t12 bgr_0.V1.t11 bgr_0.V_p_2.t5 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X393 V_OSC.t0 VCO_FD_magic_0.vco2_3_0.V8.t3 VCO_FD_magic_0.vco2_3_0.V2.t0 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X394 GNDA.t96 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X395 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 GNDA.t284 a_8930_n1530.t6 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X397 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X398 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 a_8930_n1530.t7 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X399 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VDDA.t398 bgr_0.V2.t25 BGR_CURRENT_OUT.t6 VDDA.t397 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X401 bgr_0.V1.t5 bgr_0.V_TOP.t44 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X402 GNDA.t221 GNDA.t223 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X403 bgr_0.V_TOP.t45 VDDA.t184 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t155 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X405 VDDA.t161 a_1870_180.t2 pfd_8_0.Reset.t0 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X406 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X407 VDDA.t76 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X408 bgr_0.V_TOP.t46 VDDA.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 GNDA.t29 VDDA.t430 VCO_FD_magic_0.vco2_3_0.V7.t2 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X410 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 a_2350_1390.t0 pfd_8_0.before_Reset.t4 VDDA.t115 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X412 a_6490_4630.t1 opamp_cell_4_0.VIN+.t8 a_5970_4630.t1 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X413 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 a_6330_n1530.t7 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X414 a_6490_4630.t3 a_6200_5250.t7 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X415 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VDDA.t88 bgr_0.1st_Vout_2.t34 bgr_0.V2.t1 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X417 VDDA.t20 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X418 GNDA.t288 a_1870_180.t3 pfd_8_0.Reset.t1 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X419 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X420 bgr_0.1st_Vout_2.t4 a_n1450_5080.t22 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X421 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 a_7630_n1530.t7 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X422 V_CONT.t0 pfd_8_0.DOWN_input.t5 GNDA.t31 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X423 pfd_8_0.QA_b.t0 pfd_8_0.QA.t6 a_n30_1390.t0 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X424 VDDA.t147 bgr_0.V2.t26 bgr_0.V_CUR_REF_REG.t2 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X425 GNDA.t43 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 VCO_FD_magic_0.div120_2_0.div4.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X426 VDDA.t140 bgr_0.V_TOP.t47 bgr_0.V1.t4 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X427 GNDA.t102 a_3160_9910.t1 GNDA.t101 sky130_fd_pr__res_xhigh_po_0p35 l=6
X428 VDDA.t392 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t1 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X429 VCO_FD_magic_0.vco2_3_0.V8.t1 VCO_FD_magic_0.vco2_3_0.V9.t3 VCO_FD_magic_0.vco2_3_0.V5.t0 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X430 VDDA.t149 bgr_0.V2.t27 bgr_0.V_CUR_REF_REG.t1 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X431 VDDA.t24 bgr_0.V_TOP.t48 bgr_0.V1.t3 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X432 a_n1450_5080.t3 a_n1450_5080.t2 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X433 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 VCO_FD_magic_0.div120_2_0.div24.t14 GNDA.t203 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X434 GNDA.t72 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X435 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 opamp_cell_4_0.VIN+.t4 BGR_CURRENT_OUT.t19 GNDA.t168 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X437 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 pfd_8_0.before_Reset.t0 pfd_8_0.QA.t7 a_1910_2010.t0 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X439 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 GNDA.t186 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X440 GNDA.t308 V_CONT.t15 VCO_FD_magic_0.vco2_3_0.V5.t1 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X441 pfd_8_0.before_Reset.t2 pfd_8_0.QB.t8 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X442 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X444 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X445 VDDA.t233 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t0 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X446 a_6320_5840.t8 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t2 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X447 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X448 BGR_CURRENT_OUT.t5 bgr_0.V2.t28 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X449 bgr_0.1st_Vout_1.t2 bgr_0.Vin+.t10 bgr_0.V_p_1.t5 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X450 GNDA.t2 pfd_8_0.E.t6 pfd_8_0.QA.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X451 pfd_8_0.UP_input.t2 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t6 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X452 a_490_1390.t0 pfd_8_0.QA_b.t6 pfd_8_0.QA.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X453 a_n1450_5080.t1 a_n1450_5080.t0 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X454 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 pfd_8_0.F.t1 pfd_8_0.F_b.t4 a_870_630.t1 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X456 bgr_0.cap_res1.t0 bgr_0.V_TOP.t1 GNDA.t62 sky130_fd_pr__res_high_po_0p35 l=2.05
X457 GNDA.t219 GNDA.t217 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X458 VCO_FD_magic_0.vco2_3_0.V1.t1 VCO_FD_magic_0.vco2_3_0.V1.t0 VDDA.t343 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X459 bgr_0.V_TOP.t4 VDDA.t267 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X460 bgr_0.V_p_2.t1 bgr_0.V_CUR_REF_REG.t17 bgr_0.1st_Vout_2.t3 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X461 bgr_0.V_TOP.t49 VDDA.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 opamp_cell_4_0.VIN+.t0 pfd_8_0.opamp_out.t15 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X463 VDDA.t157 bgr_0.V2.t29 bgr_0.V_CUR_REF_REG.t0 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
R0 GNDA.n2402 GNDA.n360 323538
R1 GNDA.n1094 GNDA.n106 215600
R2 GNDA.t149 GNDA.n2764 164510
R3 GNDA.n1095 GNDA.n1086 158481
R4 GNDA.n360 GNDA.t40 132387
R5 GNDA.n1095 GNDA.n1094 103400
R6 GNDA.n2490 GNDA.n106 39732
R7 GNDA.n194 GNDA.n193 36300
R8 GNDA.n2402 GNDA.n2401 29837.5
R9 GNDA.n1086 GNDA.n361 9511.11
R10 GNDA.n2400 GNDA.n361 8900
R11 GNDA.n302 GNDA.n301 8097.04
R12 GNDA.n2765 GNDA.n23 6000.99
R13 GNDA.n2403 GNDA.n2402 4738.46
R14 GNDA.n2400 GNDA.n2399 4458.3
R15 GNDA.n1087 GNDA.n1086 4106.67
R16 GNDA.t221 GNDA.n361 4106.67
R17 GNDA.n2401 GNDA.n2400 3344.05
R18 GNDA.n24 GNDA.t298 2012.26
R19 GNDA.t99 GNDA.t69 1670.37
R20 GNDA.n2765 GNDA.t149 1622.77
R21 GNDA.n2403 GNDA.t275 1568.52
R22 GNDA.n1900 GNDA.n1899 1515.29
R23 GNDA.n1927 GNDA.n1072 1515.29
R24 GNDA.n1901 GNDA.n1900 1482.87
R25 GNDA.n1971 GNDA.n1072 1482.87
R26 GNDA.n1964 GNDA.n1933 1214.72
R27 GNDA.n1964 GNDA.n1963 1214.72
R28 GNDA.n1963 GNDA.n1962 1214.72
R29 GNDA.n1962 GNDA.n1936 1214.72
R30 GNDA.n1936 GNDA.n382 1214.72
R31 GNDA.n1954 GNDA.n381 1214.72
R32 GNDA.n1954 GNDA.n1953 1214.72
R33 GNDA.n1953 GNDA.n1952 1214.72
R34 GNDA.n1952 GNDA.n1948 1214.72
R35 GNDA.n1948 GNDA.n380 1214.72
R36 GNDA.n1864 GNDA.n1824 1214.72
R37 GNDA.n1864 GNDA.n1863 1214.72
R38 GNDA.n1863 GNDA.n1862 1214.72
R39 GNDA.n1862 GNDA.n1832 1214.72
R40 GNDA.n1832 GNDA.n370 1214.72
R41 GNDA.n1854 GNDA.n371 1214.72
R42 GNDA.n1854 GNDA.n1853 1214.72
R43 GNDA.n1853 GNDA.n1852 1214.72
R44 GNDA.n1852 GNDA.n1843 1214.72
R45 GNDA.n1843 GNDA.n372 1214.72
R46 GNDA.n226 GNDA.n69 1204.13
R47 GNDA.n225 GNDA.n58 1204.13
R48 GNDA.n196 GNDA.n47 1204.13
R49 GNDA.n172 GNDA.n171 1186
R50 GNDA.n306 GNDA.n305 1186
R51 GNDA.n130 GNDA.n129 1186
R52 GNDA.n179 GNDA.n178 1186
R53 GNDA.n2527 GNDA.n2526 1182.8
R54 GNDA.n2492 GNDA.n83 1182.8
R55 GNDA.n2401 GNDA.n23 1176.24
R56 GNDA.n185 GNDA.n180 1173.78
R57 GNDA.n192 GNDA.n186 1173.78
R58 GNDA.n2763 GNDA.n25 1173.78
R59 GNDA.n2745 GNDA.n24 1170
R60 GNDA.t221 GNDA.n382 823.313
R61 GNDA.t221 GNDA.n370 823.313
R62 GNDA.n2764 GNDA.n24 798.423
R63 GNDA.n2452 GNDA.t311 794.444
R64 GNDA.n2451 GNDA.t321 794.444
R65 GNDA.t73 GNDA.t154 767.181
R66 GNDA.t86 GNDA.t322 744.615
R67 GNDA.n1877 GNDA.n367 729.283
R68 GNDA.n1877 GNDA.n1875 729.283
R69 GNDA.n1883 GNDA.n1875 729.283
R70 GNDA.n1884 GNDA.n1883 729.283
R71 GNDA.n1885 GNDA.n1884 729.283
R72 GNDA.n1891 GNDA.n1871 729.283
R73 GNDA.n1892 GNDA.n1891 729.283
R74 GNDA.n1893 GNDA.n1892 729.283
R75 GNDA.n1893 GNDA.n1825 729.283
R76 GNDA.n1899 GNDA.n1825 729.283
R77 GNDA.n1901 GNDA.n1820 729.283
R78 GNDA.n1908 GNDA.n1820 729.283
R79 GNDA.n1909 GNDA.n1908 729.283
R80 GNDA.n1910 GNDA.n1909 729.283
R81 GNDA.n1910 GNDA.n1080 729.283
R82 GNDA.n1918 GNDA.n1917 729.283
R83 GNDA.n1918 GNDA.n1076 729.283
R84 GNDA.n1925 GNDA.n1076 729.283
R85 GNDA.n1926 GNDA.n1925 729.283
R86 GNDA.n1927 GNDA.n1926 729.283
R87 GNDA.n1972 GNDA.n1971 729.283
R88 GNDA.n1973 GNDA.n1972 729.283
R89 GNDA.n1973 GNDA.n1068 729.283
R90 GNDA.n1979 GNDA.n1068 729.283
R91 GNDA.n1980 GNDA.n1979 729.283
R92 GNDA.n1981 GNDA.n1064 729.283
R93 GNDA.n1988 GNDA.n1064 729.283
R94 GNDA.n1989 GNDA.n1988 729.283
R95 GNDA.n1990 GNDA.n1989 729.283
R96 GNDA.n1990 GNDA.n373 729.283
R97 GNDA.n180 GNDA.t328 728.524
R98 GNDA.n186 GNDA.t333 728.524
R99 GNDA.n25 GNDA.t331 728.524
R100 GNDA.n191 GNDA.n190 686.717
R101 GNDA.n184 GNDA.n32 686.717
R102 GNDA.n2762 GNDA.n2761 686.717
R103 GNDA.n1788 GNDA.n1787 686.717
R104 GNDA.n1807 GNDA.n1806 686.717
R105 GNDA.n1098 GNDA.n1097 686.717
R106 GNDA.n1097 GNDA.n1085 686.717
R107 GNDA.n1799 GNDA.n1798 686.717
R108 GNDA.n1780 GNDA.n1779 686.717
R109 GNDA.n2762 GNDA.n27 686.717
R110 GNDA.n184 GNDA.n183 686.717
R111 GNDA.n191 GNDA.n188 686.717
R112 GNDA.n251 GNDA.n250 669.307
R113 GNDA.n254 GNDA.n253 669.307
R114 GNDA.n272 GNDA.n271 669.307
R115 GNDA.n275 GNDA.n274 669.307
R116 GNDA.n299 GNDA.n298 669.307
R117 GNDA.n293 GNDA.n195 669.307
R118 GNDA.n1680 GNDA.n1679 669.307
R119 GNDA.n1763 GNDA.n1762 669.307
R120 GNDA.n1813 GNDA.n1081 654.447
R121 GNDA.t143 GNDA.t159 591.035
R122 GNDA.n2768 GNDA.n2767 585.003
R123 GNDA.n2405 GNDA.n2404 585.003
R124 GNDA.n2453 GNDA.n2452 585.001
R125 GNDA.n2407 GNDA.n2406 585.001
R126 GNDA.n359 GNDA.n347 585.001
R127 GNDA.n358 GNDA.n344 585.001
R128 GNDA.n2451 GNDA.n2450 585.001
R129 GNDA.n1093 GNDA.n1092 585.001
R130 GNDA.n1091 GNDA.n1090 585.001
R131 GNDA.n1089 GNDA.n1088 585.001
R132 GNDA.n2494 GNDA.n2493 585.001
R133 GNDA.n2491 GNDA.n101 585.001
R134 GNDA.n2525 GNDA.n2524 585.001
R135 GNDA.n2773 GNDA.n2772 585.001
R136 GNDA.n2771 GNDA.n19 585.001
R137 GNDA.n2770 GNDA.n16 585.001
R138 GNDA.n2769 GNDA.n13 585.001
R139 GNDA.n2766 GNDA.n2 585.001
R140 GNDA.n170 GNDA.n169 585.001
R141 GNDA.n304 GNDA.n303 585.001
R142 GNDA.n1323 GNDA.n1322 585
R143 GNDA.n1325 GNDA.n1324 585
R144 GNDA.n1327 GNDA.n1326 585
R145 GNDA.n1329 GNDA.n1328 585
R146 GNDA.n1331 GNDA.n1330 585
R147 GNDA.n1333 GNDA.n1332 585
R148 GNDA.n1335 GNDA.n1334 585
R149 GNDA.n1337 GNDA.n1336 585
R150 GNDA.n1339 GNDA.n1338 585
R151 GNDA.n1341 GNDA.n1340 585
R152 GNDA.n1342 GNDA.n631 585
R153 GNDA.n2237 GNDA.n631 585
R154 GNDA.n1344 GNDA.n1343 585
R155 GNDA.n1345 GNDA.n1344 585
R156 GNDA.n612 GNDA.n611 585
R157 GNDA.n614 GNDA.n613 585
R158 GNDA.n616 GNDA.n615 585
R159 GNDA.n618 GNDA.n617 585
R160 GNDA.n620 GNDA.n619 585
R161 GNDA.n622 GNDA.n621 585
R162 GNDA.n624 GNDA.n623 585
R163 GNDA.n625 GNDA.n590 585
R164 GNDA.n628 GNDA.n627 585
R165 GNDA.n626 GNDA.n589 585
R166 GNDA.n579 GNDA.n578 585
R167 GNDA.n2237 GNDA.n579 585
R168 GNDA.n2240 GNDA.n2239 585
R169 GNDA.n2240 GNDA.n577 585
R170 GNDA.n2235 GNDA.n2234 585
R171 GNDA.n2233 GNDA.n638 585
R172 GNDA.n2232 GNDA.n637 585
R173 GNDA.n2237 GNDA.n637 585
R174 GNDA.n2231 GNDA.n2230 585
R175 GNDA.n2229 GNDA.n2228 585
R176 GNDA.n2227 GNDA.n2226 585
R177 GNDA.n2225 GNDA.n2224 585
R178 GNDA.n2223 GNDA.n2222 585
R179 GNDA.n2221 GNDA.n2220 585
R180 GNDA.n2219 GNDA.n2218 585
R181 GNDA.n2217 GNDA.n2216 585
R182 GNDA.n2215 GNDA.n2214 585
R183 GNDA.n2214 GNDA.n2213 585
R184 GNDA.n2113 GNDA.n917 585
R185 GNDA.n917 GNDA.n380 585
R186 GNDA.n1947 GNDA.n916 585
R187 GNDA.n1948 GNDA.n1947 585
R188 GNDA.n1950 GNDA.n1946 585
R189 GNDA.n1952 GNDA.n1946 585
R190 GNDA.n1949 GNDA.n1945 585
R191 GNDA.n1953 GNDA.n1945 585
R192 GNDA.n1944 GNDA.n1942 585
R193 GNDA.n1954 GNDA.n1944 585
R194 GNDA.n1943 GNDA.n1940 585
R195 GNDA.n1943 GNDA.n381 585
R196 GNDA.n1958 GNDA.n1939 585
R197 GNDA.n1939 GNDA.n382 585
R198 GNDA.n1959 GNDA.n1938 585
R199 GNDA.n1938 GNDA.n1936 585
R200 GNDA.n1960 GNDA.n1935 585
R201 GNDA.n1962 GNDA.n1935 585
R202 GNDA.n1934 GNDA.n1931 585
R203 GNDA.n1963 GNDA.n1934 585
R204 GNDA.n1966 GNDA.n1930 585
R205 GNDA.n1964 GNDA.n1930 585
R206 GNDA.n1967 GNDA.n1929 585
R207 GNDA.n1933 GNDA.n1929 585
R208 GNDA.n1967 GNDA.n1073 585
R209 GNDA.n1933 GNDA.n1073 585
R210 GNDA.n1966 GNDA.n1965 585
R211 GNDA.n1965 GNDA.n1964 585
R212 GNDA.n1932 GNDA.n1931 585
R213 GNDA.n1963 GNDA.n1932 585
R214 GNDA.n1961 GNDA.n1960 585
R215 GNDA.n1962 GNDA.n1961 585
R216 GNDA.n1959 GNDA.n1937 585
R217 GNDA.n1937 GNDA.n1936 585
R218 GNDA.n1958 GNDA.n1957 585
R219 GNDA.n1957 GNDA.n382 585
R220 GNDA.n1956 GNDA.n1940 585
R221 GNDA.n1956 GNDA.n381 585
R222 GNDA.n1955 GNDA.n1942 585
R223 GNDA.n1955 GNDA.n1954 585
R224 GNDA.n1949 GNDA.n1941 585
R225 GNDA.n1953 GNDA.n1941 585
R226 GNDA.n1951 GNDA.n1950 585
R227 GNDA.n1952 GNDA.n1951 585
R228 GNDA.n916 GNDA.n915 585
R229 GNDA.n1948 GNDA.n915 585
R230 GNDA.n2114 GNDA.n2113 585
R231 GNDA.n2114 GNDA.n380 585
R232 GNDA.n2364 GNDA.n441 585
R233 GNDA.n888 GNDA.n440 585
R234 GNDA.n891 GNDA.n890 585
R235 GNDA.n896 GNDA.n886 585
R236 GNDA.n897 GNDA.n885 585
R237 GNDA.n898 GNDA.n883 585
R238 GNDA.n882 GNDA.n879 585
R239 GNDA.n904 GNDA.n878 585
R240 GNDA.n905 GNDA.n877 585
R241 GNDA.n906 GNDA.n875 585
R242 GNDA.n874 GNDA.n870 585
R243 GNDA.n911 GNDA.n869 585
R244 GNDA.n911 GNDA.n910 585
R245 GNDA.n908 GNDA.n870 585
R246 GNDA.n907 GNDA.n906 585
R247 GNDA.n907 GNDA.n383 585
R248 GNDA.n905 GNDA.n872 585
R249 GNDA.n904 GNDA.n903 585
R250 GNDA.n901 GNDA.n879 585
R251 GNDA.n899 GNDA.n898 585
R252 GNDA.n897 GNDA.n880 585
R253 GNDA.n896 GNDA.n895 585
R254 GNDA.n893 GNDA.n891 585
R255 GNDA.n440 GNDA.n439 585
R256 GNDA.n2365 GNDA.n2364 585
R257 GNDA.n2365 GNDA.n383 585
R258 GNDA.n1668 GNDA.n1148 585
R259 GNDA.n1169 GNDA.n1149 585
R260 GNDA.n1664 GNDA.n1663 585
R261 GNDA.n1168 GNDA.n1167 585
R262 GNDA.n1172 GNDA.n1171 585
R263 GNDA.n1656 GNDA.n1655 585
R264 GNDA.n1654 GNDA.n1653 585
R265 GNDA.n1652 GNDA.n1176 585
R266 GNDA.n1175 GNDA.n1174 585
R267 GNDA.n1646 GNDA.n1645 585
R268 GNDA.n1644 GNDA.n1643 585
R269 GNDA.n1642 GNDA.n1446 585
R270 GNDA.n1642 GNDA.n1641 585
R271 GNDA.n1643 GNDA.n1177 585
R272 GNDA.n1647 GNDA.n1646 585
R273 GNDA.n1649 GNDA.n1174 585
R274 GNDA.n1652 GNDA.n1651 585
R275 GNDA.n1653 GNDA.n1173 585
R276 GNDA.n1657 GNDA.n1656 585
R277 GNDA.n1659 GNDA.n1172 585
R278 GNDA.n1660 GNDA.n1168 585
R279 GNDA.n1663 GNDA.n1662 585
R280 GNDA.n1170 GNDA.n1169 585
R281 GNDA.n1554 GNDA.n1148 585
R282 GNDA.n1399 GNDA.n1211 585
R283 GNDA.n1400 GNDA.n1209 585
R284 GNDA.n1403 GNDA.n1208 585
R285 GNDA.n1404 GNDA.n1206 585
R286 GNDA.n1407 GNDA.n1205 585
R287 GNDA.n1408 GNDA.n1203 585
R288 GNDA.n1411 GNDA.n1202 585
R289 GNDA.n1412 GNDA.n1200 585
R290 GNDA.n1413 GNDA.n1199 585
R291 GNDA.n1197 GNDA.n1190 585
R292 GNDA.n1419 GNDA.n1189 585
R293 GNDA.n1420 GNDA.n1187 585
R294 GNDA.n1420 GNDA.n1185 585
R295 GNDA.n1419 GNDA.n1418 585
R296 GNDA.n1191 GNDA.n1190 585
R297 GNDA.n1414 GNDA.n1413 585
R298 GNDA.n1412 GNDA.n1196 585
R299 GNDA.n1411 GNDA.n1410 585
R300 GNDA.n1409 GNDA.n1408 585
R301 GNDA.n1407 GNDA.n1406 585
R302 GNDA.n1405 GNDA.n1404 585
R303 GNDA.n1403 GNDA.n1402 585
R304 GNDA.n1401 GNDA.n1400 585
R305 GNDA.n1399 GNDA.n1398 585
R306 GNDA.n2370 GNDA.n431 585
R307 GNDA.n2371 GNDA.n422 585
R308 GNDA.n2374 GNDA.n421 585
R309 GNDA.n2375 GNDA.n420 585
R310 GNDA.n2378 GNDA.n419 585
R311 GNDA.n2379 GNDA.n418 585
R312 GNDA.n2382 GNDA.n417 585
R313 GNDA.n2384 GNDA.n416 585
R314 GNDA.n2385 GNDA.n415 585
R315 GNDA.n2386 GNDA.n414 585
R316 GNDA.n423 GNDA.n406 585
R317 GNDA.n2392 GNDA.n402 585
R318 GNDA.n2392 GNDA.n2391 585
R319 GNDA.n408 GNDA.n406 585
R320 GNDA.n2387 GNDA.n2386 585
R321 GNDA.n2385 GNDA.n413 585
R322 GNDA.n2384 GNDA.n2383 585
R323 GNDA.n2382 GNDA.n2381 585
R324 GNDA.n2380 GNDA.n2379 585
R325 GNDA.n2378 GNDA.n2377 585
R326 GNDA.n2376 GNDA.n2375 585
R327 GNDA.n2374 GNDA.n2373 585
R328 GNDA.n2372 GNDA.n2371 585
R329 GNDA.n2370 GNDA.n2369 585
R330 GNDA.n1848 GNDA.n682 585
R331 GNDA.n682 GNDA.n372 585
R332 GNDA.n1849 GNDA.n1846 585
R333 GNDA.n1846 GNDA.n1843 585
R334 GNDA.n1850 GNDA.n1842 585
R335 GNDA.n1852 GNDA.n1842 585
R336 GNDA.n1845 GNDA.n1841 585
R337 GNDA.n1853 GNDA.n1841 585
R338 GNDA.n1840 GNDA.n1838 585
R339 GNDA.n1854 GNDA.n1840 585
R340 GNDA.n1839 GNDA.n1836 585
R341 GNDA.n1839 GNDA.n371 585
R342 GNDA.n1858 GNDA.n1835 585
R343 GNDA.n1835 GNDA.n370 585
R344 GNDA.n1859 GNDA.n1834 585
R345 GNDA.n1834 GNDA.n1832 585
R346 GNDA.n1860 GNDA.n1831 585
R347 GNDA.n1862 GNDA.n1831 585
R348 GNDA.n1830 GNDA.n1828 585
R349 GNDA.n1863 GNDA.n1830 585
R350 GNDA.n1866 GNDA.n1827 585
R351 GNDA.n1864 GNDA.n1827 585
R352 GNDA.n1868 GNDA.n1867 585
R353 GNDA.n1868 GNDA.n1824 585
R354 GNDA.n1867 GNDA.n1823 585
R355 GNDA.n1824 GNDA.n1823 585
R356 GNDA.n1866 GNDA.n1865 585
R357 GNDA.n1865 GNDA.n1864 585
R358 GNDA.n1829 GNDA.n1828 585
R359 GNDA.n1863 GNDA.n1829 585
R360 GNDA.n1861 GNDA.n1860 585
R361 GNDA.n1862 GNDA.n1861 585
R362 GNDA.n1859 GNDA.n1833 585
R363 GNDA.n1833 GNDA.n1832 585
R364 GNDA.n1858 GNDA.n1857 585
R365 GNDA.n1857 GNDA.n370 585
R366 GNDA.n1856 GNDA.n1836 585
R367 GNDA.n1856 GNDA.n371 585
R368 GNDA.n1855 GNDA.n1838 585
R369 GNDA.n1855 GNDA.n1854 585
R370 GNDA.n1845 GNDA.n1837 585
R371 GNDA.n1853 GNDA.n1837 585
R372 GNDA.n1851 GNDA.n1850 585
R373 GNDA.n1852 GNDA.n1851 585
R374 GNDA.n1849 GNDA.n1844 585
R375 GNDA.n1844 GNDA.n1843 585
R376 GNDA.n1848 GNDA.n1847 585
R377 GNDA.n1847 GNDA.n372 585
R378 GNDA.n1898 GNDA.n1897 585
R379 GNDA.n1899 GNDA.n1898 585
R380 GNDA.n1896 GNDA.n1826 585
R381 GNDA.n1826 GNDA.n1825 585
R382 GNDA.n1895 GNDA.n1894 585
R383 GNDA.n1894 GNDA.n1893 585
R384 GNDA.n1870 GNDA.n1869 585
R385 GNDA.n1892 GNDA.n1870 585
R386 GNDA.n1890 GNDA.n1889 585
R387 GNDA.n1891 GNDA.n1890 585
R388 GNDA.n1888 GNDA.n1872 585
R389 GNDA.n1872 GNDA.n1871 585
R390 GNDA.n1887 GNDA.n1886 585
R391 GNDA.n1886 GNDA.n1885 585
R392 GNDA.n1874 GNDA.n1873 585
R393 GNDA.n1884 GNDA.n1874 585
R394 GNDA.n1882 GNDA.n1881 585
R395 GNDA.n1883 GNDA.n1882 585
R396 GNDA.n1880 GNDA.n1876 585
R397 GNDA.n1876 GNDA.n1875 585
R398 GNDA.n1879 GNDA.n1878 585
R399 GNDA.n1878 GNDA.n1877 585
R400 GNDA.n640 GNDA.n639 585
R401 GNDA.n639 GNDA.n367 585
R402 GNDA.n1928 GNDA.n1074 585
R403 GNDA.n1928 GNDA.n1927 585
R404 GNDA.n1922 GNDA.n1075 585
R405 GNDA.n1926 GNDA.n1075 585
R406 GNDA.n1924 GNDA.n1923 585
R407 GNDA.n1925 GNDA.n1924 585
R408 GNDA.n1921 GNDA.n1077 585
R409 GNDA.n1077 GNDA.n1076 585
R410 GNDA.n1920 GNDA.n1919 585
R411 GNDA.n1919 GNDA.n1918 585
R412 GNDA.n1079 GNDA.n1078 585
R413 GNDA.n1917 GNDA.n1079 585
R414 GNDA.n1913 GNDA.n1912 585
R415 GNDA.n1912 GNDA.n1080 585
R416 GNDA.n1911 GNDA.n1818 585
R417 GNDA.n1911 GNDA.n1910 585
R418 GNDA.n1905 GNDA.n1819 585
R419 GNDA.n1909 GNDA.n1819 585
R420 GNDA.n1907 GNDA.n1906 585
R421 GNDA.n1908 GNDA.n1907 585
R422 GNDA.n1904 GNDA.n1821 585
R423 GNDA.n1821 GNDA.n1820 585
R424 GNDA.n1903 GNDA.n1902 585
R425 GNDA.n1902 GNDA.n1901 585
R426 GNDA.n1992 GNDA.n1061 585
R427 GNDA.n1992 GNDA.n373 585
R428 GNDA.n1991 GNDA.n1063 585
R429 GNDA.n1991 GNDA.n1990 585
R430 GNDA.n1985 GNDA.n1062 585
R431 GNDA.n1989 GNDA.n1062 585
R432 GNDA.n1987 GNDA.n1986 585
R433 GNDA.n1988 GNDA.n1987 585
R434 GNDA.n1984 GNDA.n1065 585
R435 GNDA.n1065 GNDA.n1064 585
R436 GNDA.n1983 GNDA.n1982 585
R437 GNDA.n1982 GNDA.n1981 585
R438 GNDA.n1067 GNDA.n1066 585
R439 GNDA.n1980 GNDA.n1067 585
R440 GNDA.n1978 GNDA.n1977 585
R441 GNDA.n1979 GNDA.n1978 585
R442 GNDA.n1976 GNDA.n1069 585
R443 GNDA.n1069 GNDA.n1068 585
R444 GNDA.n1975 GNDA.n1974 585
R445 GNDA.n1974 GNDA.n1973 585
R446 GNDA.n1071 GNDA.n1070 585
R447 GNDA.n1972 GNDA.n1071 585
R448 GNDA.n1970 GNDA.n1969 585
R449 GNDA.n1971 GNDA.n1970 585
R450 GNDA.n1083 GNDA.n1082 585
R451 GNDA.n1916 GNDA.n1915 585
R452 GNDA.t221 GNDA.n1916 585
R453 GNDA.n2395 GNDA.n2394 585
R454 GNDA.n403 GNDA.n401 585
R455 GNDA.n592 GNDA.n591 585
R456 GNDA.n594 GNDA.n593 585
R457 GNDA.n596 GNDA.n595 585
R458 GNDA.n598 GNDA.n597 585
R459 GNDA.n600 GNDA.n599 585
R460 GNDA.n602 GNDA.n601 585
R461 GNDA.n604 GNDA.n603 585
R462 GNDA.n606 GNDA.n605 585
R463 GNDA.n608 GNDA.n607 585
R464 GNDA.n610 GNDA.n609 585
R465 GNDA.n868 GNDA.n867 585
R466 GNDA.n866 GNDA.n865 585
R467 GNDA.n864 GNDA.n863 585
R468 GNDA.n862 GNDA.n861 585
R469 GNDA.n860 GNDA.n859 585
R470 GNDA.n858 GNDA.n857 585
R471 GNDA.n856 GNDA.n855 585
R472 GNDA.n854 GNDA.n853 585
R473 GNDA.n852 GNDA.n851 585
R474 GNDA.n850 GNDA.n849 585
R475 GNDA.n848 GNDA.n847 585
R476 GNDA.n407 GNDA.n404 585
R477 GNDA.n825 GNDA.n824 585
R478 GNDA.n827 GNDA.n826 585
R479 GNDA.n829 GNDA.n828 585
R480 GNDA.n831 GNDA.n830 585
R481 GNDA.n833 GNDA.n832 585
R482 GNDA.n835 GNDA.n834 585
R483 GNDA.n837 GNDA.n836 585
R484 GNDA.n839 GNDA.n838 585
R485 GNDA.n841 GNDA.n840 585
R486 GNDA.n843 GNDA.n842 585
R487 GNDA.n845 GNDA.n844 585
R488 GNDA.n871 GNDA.n846 585
R489 GNDA.n2117 GNDA.n405 585
R490 GNDA.n2117 GNDA.n2116 585
R491 GNDA.n2212 GNDA.n641 585
R492 GNDA.n2199 GNDA.n642 585
R493 GNDA.n2208 GNDA.n2207 585
R494 GNDA.n661 GNDA.n659 585
R495 GNDA.n2124 GNDA.n2123 585
R496 GNDA.n2128 GNDA.n2127 585
R497 GNDA.n2130 GNDA.n2129 585
R498 GNDA.n2137 GNDA.n2136 585
R499 GNDA.n2135 GNDA.n2121 585
R500 GNDA.n2143 GNDA.n2142 585
R501 GNDA.n2145 GNDA.n2144 585
R502 GNDA.n2119 GNDA.n2118 585
R503 GNDA.n913 GNDA.n684 585
R504 GNDA.n2116 GNDA.n684 585
R505 GNDA.n683 GNDA.n405 585
R506 GNDA.n2116 GNDA.n683 585
R507 GNDA.n994 GNDA.n993 585
R508 GNDA.n1018 GNDA.n996 585
R509 GNDA.n1020 GNDA.n1019 585
R510 GNDA.n1016 GNDA.n1015 585
R511 GNDA.n1014 GNDA.n1013 585
R512 GNDA.n1009 GNDA.n1008 585
R513 GNDA.n1007 GNDA.n1006 585
R514 GNDA.n1002 GNDA.n1001 585
R515 GNDA.n1000 GNDA.n920 585
R516 GNDA.n1028 GNDA.n1027 585
R517 GNDA.n1030 GNDA.n1029 585
R518 GNDA.n1033 GNDA.n1032 585
R519 GNDA.n2115 GNDA.n913 585
R520 GNDA.n2116 GNDA.n2115 585
R521 GNDA.n2111 GNDA.n914 585
R522 GNDA.n2109 GNDA.n2108 585
R523 GNDA.n2107 GNDA.n2106 585
R524 GNDA.n2023 GNDA.n1036 585
R525 GNDA.n2025 GNDA.n2024 585
R526 GNDA.n2029 GNDA.n2028 585
R527 GNDA.n2031 GNDA.n2030 585
R528 GNDA.n2038 GNDA.n2037 585
R529 GNDA.n2036 GNDA.n2021 585
R530 GNDA.n2044 GNDA.n2043 585
R531 GNDA.n2046 GNDA.n2045 585
R532 GNDA.n2019 GNDA.n2018 585
R533 GNDA.n1300 GNDA.n1186 585
R534 GNDA.n1303 GNDA.n1302 585
R535 GNDA.n1305 GNDA.n1304 585
R536 GNDA.n1307 GNDA.n1298 585
R537 GNDA.n1309 GNDA.n1308 585
R538 GNDA.n1310 GNDA.n1297 585
R539 GNDA.n1312 GNDA.n1311 585
R540 GNDA.n1314 GNDA.n1295 585
R541 GNDA.n1316 GNDA.n1315 585
R542 GNDA.n1317 GNDA.n1294 585
R543 GNDA.n1319 GNDA.n1318 585
R544 GNDA.n1321 GNDA.n1293 585
R545 GNDA.n1445 GNDA.n1444 585
R546 GNDA.n1443 GNDA.n1442 585
R547 GNDA.n1441 GNDA.n1180 585
R548 GNDA.n1439 GNDA.n1438 585
R549 GNDA.n1437 GNDA.n1181 585
R550 GNDA.n1436 GNDA.n1435 585
R551 GNDA.n1433 GNDA.n1182 585
R552 GNDA.n1431 GNDA.n1430 585
R553 GNDA.n1429 GNDA.n1183 585
R554 GNDA.n1428 GNDA.n1427 585
R555 GNDA.n1425 GNDA.n1184 585
R556 GNDA.n1423 GNDA.n1422 585
R557 GNDA.n1620 GNDA.n1619 585
R558 GNDA.n1621 GNDA.n1454 585
R559 GNDA.n1623 GNDA.n1622 585
R560 GNDA.n1625 GNDA.n1452 585
R561 GNDA.n1627 GNDA.n1626 585
R562 GNDA.n1628 GNDA.n1451 585
R563 GNDA.n1630 GNDA.n1629 585
R564 GNDA.n1632 GNDA.n1449 585
R565 GNDA.n1634 GNDA.n1633 585
R566 GNDA.n1635 GNDA.n1448 585
R567 GNDA.n1637 GNDA.n1636 585
R568 GNDA.n1639 GNDA.n1447 585
R569 GNDA.n435 GNDA.n434 585
R570 GNDA.n2367 GNDA.n435 585
R571 GNDA.n2355 GNDA.n2354 585
R572 GNDA.n2352 GNDA.n576 585
R573 GNDA.n2243 GNDA.n2242 585
R574 GNDA.n2347 GNDA.n2346 585
R575 GNDA.n2345 GNDA.n2344 585
R576 GNDA.n2271 GNDA.n2247 585
R577 GNDA.n2273 GNDA.n2272 585
R578 GNDA.n2278 GNDA.n2277 585
R579 GNDA.n2276 GNDA.n2269 585
R580 GNDA.n2284 GNDA.n2283 585
R581 GNDA.n2286 GNDA.n2285 585
R582 GNDA.n2267 GNDA.n2266 585
R583 GNDA.n437 GNDA.n436 585
R584 GNDA.n2367 GNDA.n436 585
R585 GNDA.n2368 GNDA.n434 585
R586 GNDA.n2368 GNDA.n2367 585
R587 GNDA.n458 GNDA.n433 585
R588 GNDA.n569 GNDA.n568 585
R589 GNDA.n460 GNDA.n457 585
R590 GNDA.n563 GNDA.n562 585
R591 GNDA.n561 GNDA.n560 585
R592 GNDA.n486 GNDA.n464 585
R593 GNDA.n488 GNDA.n487 585
R594 GNDA.n493 GNDA.n492 585
R595 GNDA.n491 GNDA.n484 585
R596 GNDA.n499 GNDA.n498 585
R597 GNDA.n501 GNDA.n500 585
R598 GNDA.n451 GNDA.n442 585
R599 GNDA.n2366 GNDA.n437 585
R600 GNDA.n2367 GNDA.n2366 585
R601 GNDA.n2362 GNDA.n438 585
R602 GNDA.n2360 GNDA.n2359 585
R603 GNDA.n766 GNDA.n445 585
R604 GNDA.n786 GNDA.n785 585
R605 GNDA.n784 GNDA.n783 585
R606 GNDA.n779 GNDA.n778 585
R607 GNDA.n777 GNDA.n776 585
R608 GNDA.n772 GNDA.n771 585
R609 GNDA.n770 GNDA.n695 585
R610 GNDA.n795 GNDA.n794 585
R611 GNDA.n797 GNDA.n796 585
R612 GNDA.n800 GNDA.n799 585
R613 GNDA.n1111 GNDA.n1110 585
R614 GNDA.n1760 GNDA.n1759 585
R615 GNDA.n1761 GNDA.n1760 585
R616 GNDA.n1678 GNDA.n1673 585
R617 GNDA.n1675 GNDA.n1672 585
R618 GNDA.n1681 GNDA.n1672 585
R619 GNDA.n1805 GNDA.n1794 585
R620 GNDA.n1804 GNDA.n1803 585
R621 GNDA.n1804 GNDA.t173 585
R622 GNDA.n1801 GNDA.n1797 585
R623 GNDA.n1786 GNDA.n1785 585
R624 GNDA.n1783 GNDA.n1775 585
R625 GNDA.n1775 GNDA.t107 585
R626 GNDA.n1778 GNDA.n1776 585
R627 GNDA.n1395 GNDA.n1394 585
R628 GNDA.n1394 GNDA.n1393 585
R629 GNDA.n1347 GNDA.n1346 585
R630 GNDA.n1346 GNDA.n369 585
R631 GNDA.n1348 GNDA.n1229 585
R632 GNDA.n1229 GNDA.n1228 585
R633 GNDA.n1358 GNDA.n1357 585
R634 GNDA.n1359 GNDA.n1358 585
R635 GNDA.n1231 GNDA.n1227 585
R636 GNDA.n1360 GNDA.n1227 585
R637 GNDA.n1363 GNDA.n1362 585
R638 GNDA.n1362 GNDA.n1361 585
R639 GNDA.n1364 GNDA.n1222 585
R640 GNDA.n1222 GNDA.n368 585
R641 GNDA.n1373 GNDA.n1372 585
R642 GNDA.n1374 GNDA.n1373 585
R643 GNDA.n1223 GNDA.n1221 585
R644 GNDA.n1375 GNDA.n1221 585
R645 GNDA.n1379 GNDA.n1378 585
R646 GNDA.n1378 GNDA.n1377 585
R647 GNDA.n1380 GNDA.n1215 585
R648 GNDA.n1376 GNDA.n1215 585
R649 GNDA.n1390 GNDA.n1389 585
R650 GNDA.n1391 GNDA.n1390 585
R651 GNDA.n1387 GNDA.n1214 585
R652 GNDA.n1392 GNDA.n1214 585
R653 GNDA.n1669 GNDA.n1147 585
R654 GNDA.n1670 GNDA.n1669 585
R655 GNDA.n1397 GNDA.n1395 585
R656 GNDA.n1397 GNDA.n1396 585
R657 GNDA.n1212 GNDA.n1114 585
R658 GNDA.n1114 GNDA.n1112 585
R659 GNDA.n1757 GNDA.n1756 585
R660 GNDA.n1758 GNDA.n1757 585
R661 GNDA.n1117 GNDA.n1115 585
R662 GNDA.n1115 GNDA.n1113 585
R663 GNDA.n1751 GNDA.n1750 585
R664 GNDA.n1750 GNDA.n1749 585
R665 GNDA.n1123 GNDA.n1121 585
R666 GNDA.n1748 GNDA.n1121 585
R667 GNDA.n1746 GNDA.n1745 585
R668 GNDA.n1747 GNDA.n1746 585
R669 GNDA.n1152 GNDA.n1122 585
R670 GNDA.n1162 GNDA.n1122 585
R671 GNDA.n1160 GNDA.n1159 585
R672 GNDA.n1161 GNDA.n1160 585
R673 GNDA.n1154 GNDA.n1151 585
R674 GNDA.n1151 GNDA.n1150 585
R675 GNDA.n1144 GNDA.n1143 585
R676 GNDA.n1146 GNDA.n1144 585
R677 GNDA.n1684 GNDA.n1683 585
R678 GNDA.n1683 GNDA.n1682 585
R679 GNDA.n1494 GNDA.n1145 585
R680 GNDA.n1671 GNDA.n1145 585
R681 GNDA.n1555 GNDA.n1147 585
R682 GNDA.n1556 GNDA.n1555 585
R683 GNDA.n1552 GNDA.n1551 585
R684 GNDA.n1557 GNDA.n1552 585
R685 GNDA.n1559 GNDA.n1492 585
R686 GNDA.n1559 GNDA.n1558 585
R687 GNDA.n1582 GNDA.n1581 585
R688 GNDA.n1581 GNDA.n1580 585
R689 GNDA.n1563 GNDA.n1560 585
R690 GNDA.n1579 GNDA.n1560 585
R691 GNDA.n1577 GNDA.n1576 585
R692 GNDA.n1578 GNDA.n1577 585
R693 GNDA.n1572 GNDA.n1562 585
R694 GNDA.n1562 GNDA.n1561 585
R695 GNDA.n1566 GNDA.n1565 585
R696 GNDA.n1565 GNDA.n377 585
R697 GNDA.n1567 GNDA.n1468 585
R698 GNDA.n1468 GNDA.n1467 585
R699 GNDA.n1590 GNDA.n1589 585
R700 GNDA.n1591 GNDA.n1590 585
R701 GNDA.n1470 GNDA.n1465 585
R702 GNDA.n1592 GNDA.n1465 585
R703 GNDA.n1594 GNDA.n1466 585
R704 GNDA.n1594 GNDA.n1593 585
R705 GNDA.n1595 GNDA.n1464 585
R706 GNDA.n1595 GNDA.n378 585
R707 GNDA.n1600 GNDA.n1463 585
R708 GNDA.n1602 GNDA.n1601 585
R709 GNDA.n1604 GNDA.n1461 585
R710 GNDA.n1606 GNDA.n1605 585
R711 GNDA.n1607 GNDA.n1460 585
R712 GNDA.n1609 GNDA.n1608 585
R713 GNDA.n1611 GNDA.n1458 585
R714 GNDA.n1613 GNDA.n1612 585
R715 GNDA.n1614 GNDA.n1457 585
R716 GNDA.n1616 GNDA.n1615 585
R717 GNDA.n1618 GNDA.n1455 585
R718 GNDA.n1596 GNDA.n362 585
R719 GNDA.n805 GNDA.n692 585
R720 GNDA.n807 GNDA.n806 585
R721 GNDA.n809 GNDA.n690 585
R722 GNDA.n811 GNDA.n810 585
R723 GNDA.n812 GNDA.n689 585
R724 GNDA.n814 GNDA.n813 585
R725 GNDA.n816 GNDA.n687 585
R726 GNDA.n818 GNDA.n817 585
R727 GNDA.n819 GNDA.n686 585
R728 GNDA.n821 GNDA.n820 585
R729 GNDA.n823 GNDA.n685 585
R730 GNDA.n801 GNDA.n362 585
R731 GNDA.n2014 GNDA.n2013 585
R732 GNDA.n2012 GNDA.n1056 585
R733 GNDA.n2011 GNDA.n2010 585
R734 GNDA.n2008 GNDA.n1057 585
R735 GNDA.n2006 GNDA.n2005 585
R736 GNDA.n2004 GNDA.n1058 585
R737 GNDA.n2003 GNDA.n2002 585
R738 GNDA.n2000 GNDA.n1059 585
R739 GNDA.n1998 GNDA.n1997 585
R740 GNDA.n1996 GNDA.n1060 585
R741 GNDA.n1995 GNDA.n1994 585
R742 GNDA.n2017 GNDA.n362 585
R743 GNDA.n297 GNDA.n197 585
R744 GNDA.n295 GNDA.n294 585
R745 GNDA.n212 GNDA.n208 585
R746 GNDA.n210 GNDA.n207 585
R747 GNDA.n231 GNDA.n227 585
R748 GNDA.n229 GNDA.n224 585
R749 GNDA.n2488 GNDA.n2487 585
R750 GNDA.n2489 GNDA.n2488 585
R751 GNDA.n2486 GNDA.n109 585
R752 GNDA.n2484 GNDA.n2483 585
R753 GNDA.n2482 GNDA.n108 585
R754 GNDA.n2489 GNDA.n108 585
R755 GNDA.n359 GNDA.n358 570.37
R756 GNDA.n2511 GNDA.t329 566.966
R757 GNDA.n2452 GNDA.t40 550
R758 GNDA.t311 GNDA.n2451 550
R759 GNDA.n358 GNDA.t51 550
R760 GNDA.t279 GNDA.n359 550
R761 GNDA.n2405 GNDA.t193 550
R762 GNDA.t1 GNDA.n2405 550
R763 GNDA.n2406 GNDA.t108 550
R764 GNDA.n1093 GNDA.t134 550
R765 GNDA.n1091 GNDA.t120 550
R766 GNDA.t221 GNDA.n380 512.884
R767 GNDA.t221 GNDA.n372 512.884
R768 GNDA.t169 GNDA.n2489 504.512
R769 GNDA.t221 GNDA.t26 501.745
R770 GNDA.t221 GNDA.t81 501.745
R771 GNDA.t287 GNDA.t216 496.411
R772 GNDA.n2491 GNDA.t299 462.565
R773 GNDA.t51 GNDA.t321 448.149
R774 GNDA.t275 GNDA.t279 448.149
R775 GNDA.t193 GNDA.t199 448.149
R776 GNDA.t69 GNDA.t1 448.149
R777 GNDA.t108 GNDA.t99 448.149
R778 GNDA.t53 GNDA.n2771 440
R779 GNDA.n302 GNDA.n106 421.277
R780 GNDA.t221 GNDA.n381 391.411
R781 GNDA.t221 GNDA.n371 391.411
R782 GNDA.n1885 GNDA.t221 380.848
R783 GNDA.t221 GNDA.n1080 380.848
R784 GNDA.t221 GNDA.n1980 380.848
R785 GNDA.n2525 GNDA.t49 372.308
R786 GNDA.t254 GNDA.t30 363.911
R787 GNDA.t134 GNDA.n1091 362.767
R788 GNDA.t120 GNDA.n1089 362.767
R789 GNDA.t115 GNDA.t67 361.026
R790 GNDA.n1087 GNDA.n360 351.065
R791 GNDA.t221 GNDA.n1871 348.435
R792 GNDA.n1917 GNDA.t221 348.435
R793 GNDA.n1981 GNDA.t221 348.435
R794 GNDA.n252 GNDA.t246 347.368
R795 GNDA.n228 GNDA.t266 336.329
R796 GNDA.n228 GNDA.t245 336.329
R797 GNDA.n209 GNDA.t217 336.329
R798 GNDA.n209 GNDA.t253 336.329
R799 GNDA.t221 GNDA.n364 172.876
R800 GNDA.n1666 GNDA.t221 172.876
R801 GNDA.n2406 GNDA.n23 325.926
R802 GNDA.n1416 GNDA.t221 172.615
R803 GNDA.t221 GNDA.n365 172.615
R804 GNDA.n2481 GNDA.t241 320.7
R805 GNDA.n292 GNDA.t224 320.7
R806 GNDA.t18 GNDA.t136 315.897
R807 GNDA.t277 GNDA.t225 306.015
R808 GNDA.t15 GNDA.t165 306.015
R809 GNDA.t156 GNDA.t105 306.015
R810 GNDA.n123 GNDA.t235 304.634
R811 GNDA.n173 GNDA.t261 304.634
R812 GNDA.n307 GNDA.t231 304.634
R813 GNDA.n128 GNDA.t238 304.634
R814 GNDA.n2526 GNDA.t289 304.615
R815 GNDA.n225 GNDA.t218 297.745
R816 GNDA.t144 GNDA.n226 297.745
R817 GNDA.n2559 GNDA.t137 295.933
R818 GNDA.n93 GNDA.t155 295.933
R819 GNDA.n2611 GNDA.t300 295.933
R820 GNDA.t71 GNDA.t287 293.334
R821 GNDA.n168 GNDA.t257 292.584
R822 GNDA.n115 GNDA.t249 292.584
R823 GNDA.n300 GNDA.n196 281.204
R824 GNDA.n2237 GNDA.n630 264.301
R825 GNDA.n2238 GNDA.n2237 264.301
R826 GNDA.n2237 GNDA.n584 264.301
R827 GNDA.n1599 GNDA.n1598 264.301
R828 GNDA.n804 GNDA.n803 264.301
R829 GNDA.n2016 GNDA.n1055 264.301
R830 GNDA.t27 GNDA.n1085 260
R831 GNDA.n1098 GNDA.t27 260
R832 GNDA.n2761 GNDA.t307 260
R833 GNDA.t307 GNDA.n27 260
R834 GNDA.n2492 GNDA.t310 259.488
R835 GNDA.n1619 GNDA.n1618 259.416
R836 GNDA.n1446 GNDA.n1445 259.416
R837 GNDA.n824 GNDA.n823 259.416
R838 GNDA.n869 GNDA.n868 259.416
R839 GNDA.n1994 GNDA.n1992 259.416
R840 GNDA.n1929 GNDA.n1928 259.416
R841 GNDA.n1898 GNDA.n1868 259.416
R842 GNDA.n2395 GNDA.n402 259.416
R843 GNDA.n1300 GNDA.n1187 259.416
R844 GNDA.n1721 GNDA.n1140 258.334
R845 GNDA.n1533 GNDA.n1532 258.334
R846 GNDA.n538 GNDA.n481 258.334
R847 GNDA.n749 GNDA.n748 258.334
R848 GNDA.n976 GNDA.n975 258.334
R849 GNDA.n2184 GNDA.n2183 258.334
R850 GNDA.n2323 GNDA.n2264 258.334
R851 GNDA.n1278 GNDA.n1236 258.334
R852 GNDA.n2085 GNDA.n2084 258.334
R853 GNDA.t221 GNDA.n1081 257.779
R854 GNDA.n1094 GNDA.n1093 257.447
R855 GNDA.n2551 GNDA.n2550 256.207
R856 GNDA.n2237 GNDA.n636 254.34
R857 GNDA.n2237 GNDA.n635 254.34
R858 GNDA.n2237 GNDA.n634 254.34
R859 GNDA.n2237 GNDA.n633 254.34
R860 GNDA.n2237 GNDA.n632 254.34
R861 GNDA.n2237 GNDA.n585 254.34
R862 GNDA.n2237 GNDA.n586 254.34
R863 GNDA.n2237 GNDA.n587 254.34
R864 GNDA.n2237 GNDA.n588 254.34
R865 GNDA.n2237 GNDA.n629 254.34
R866 GNDA.n2237 GNDA.n2236 254.34
R867 GNDA.n2237 GNDA.n580 254.34
R868 GNDA.n2237 GNDA.n581 254.34
R869 GNDA.n2237 GNDA.n582 254.34
R870 GNDA.n2237 GNDA.n583 254.34
R871 GNDA.n887 GNDA.n366 254.34
R872 GNDA.n889 GNDA.n366 254.34
R873 GNDA.n884 GNDA.n366 254.34
R874 GNDA.n881 GNDA.n366 254.34
R875 GNDA.n876 GNDA.n366 254.34
R876 GNDA.n873 GNDA.n366 254.34
R877 GNDA.n909 GNDA.n383 254.34
R878 GNDA.n902 GNDA.n383 254.34
R879 GNDA.n900 GNDA.n383 254.34
R880 GNDA.n894 GNDA.n383 254.34
R881 GNDA.n892 GNDA.n383 254.34
R882 GNDA.n1667 GNDA.n1666 254.34
R883 GNDA.n1666 GNDA.n1665 254.34
R884 GNDA.n1666 GNDA.n1166 254.34
R885 GNDA.n1666 GNDA.n1165 254.34
R886 GNDA.n1666 GNDA.n1164 254.34
R887 GNDA.n1666 GNDA.n1163 254.34
R888 GNDA.n1640 GNDA.n365 254.34
R889 GNDA.n1648 GNDA.n365 254.34
R890 GNDA.n1650 GNDA.n365 254.34
R891 GNDA.n1658 GNDA.n365 254.34
R892 GNDA.n1661 GNDA.n365 254.34
R893 GNDA.n1553 GNDA.n365 254.34
R894 GNDA.n1210 GNDA.n364 254.34
R895 GNDA.n1207 GNDA.n364 254.34
R896 GNDA.n1204 GNDA.n364 254.34
R897 GNDA.n1201 GNDA.n364 254.34
R898 GNDA.n1198 GNDA.n364 254.34
R899 GNDA.n1188 GNDA.n364 254.34
R900 GNDA.n1417 GNDA.n1416 254.34
R901 GNDA.n1416 GNDA.n1415 254.34
R902 GNDA.n1416 GNDA.n1195 254.34
R903 GNDA.n1416 GNDA.n1194 254.34
R904 GNDA.n1416 GNDA.n1193 254.34
R905 GNDA.n1416 GNDA.n1192 254.34
R906 GNDA.n430 GNDA.n429 254.34
R907 GNDA.n429 GNDA.n428 254.34
R908 GNDA.n429 GNDA.n427 254.34
R909 GNDA.n429 GNDA.n426 254.34
R910 GNDA.n429 GNDA.n425 254.34
R911 GNDA.n429 GNDA.n424 254.34
R912 GNDA.n2390 GNDA.n2389 254.34
R913 GNDA.n2389 GNDA.n2388 254.34
R914 GNDA.n2389 GNDA.n412 254.34
R915 GNDA.n2389 GNDA.n411 254.34
R916 GNDA.n2389 GNDA.n410 254.34
R917 GNDA.n2389 GNDA.n409 254.34
R918 GNDA.n2397 GNDA.n2396 254.34
R919 GNDA.n2397 GNDA.n400 254.34
R920 GNDA.n2397 GNDA.n399 254.34
R921 GNDA.n2397 GNDA.n398 254.34
R922 GNDA.n2397 GNDA.n397 254.34
R923 GNDA.n2397 GNDA.n396 254.34
R924 GNDA.n2397 GNDA.n395 254.34
R925 GNDA.n2397 GNDA.n394 254.34
R926 GNDA.n2397 GNDA.n393 254.34
R927 GNDA.n2397 GNDA.n392 254.34
R928 GNDA.n2397 GNDA.n391 254.34
R929 GNDA.n2397 GNDA.n390 254.34
R930 GNDA.n2397 GNDA.n389 254.34
R931 GNDA.n2397 GNDA.n388 254.34
R932 GNDA.n2397 GNDA.n387 254.34
R933 GNDA.n2397 GNDA.n386 254.34
R934 GNDA.n2397 GNDA.n385 254.34
R935 GNDA.n2397 GNDA.n384 254.34
R936 GNDA.n2211 GNDA.n2210 254.34
R937 GNDA.n2210 GNDA.n2209 254.34
R938 GNDA.n2210 GNDA.n658 254.34
R939 GNDA.n2210 GNDA.n657 254.34
R940 GNDA.n2210 GNDA.n656 254.34
R941 GNDA.n2210 GNDA.n655 254.34
R942 GNDA.n2210 GNDA.n654 254.34
R943 GNDA.n2210 GNDA.n653 254.34
R944 GNDA.n2210 GNDA.n652 254.34
R945 GNDA.n2210 GNDA.n651 254.34
R946 GNDA.n2210 GNDA.n650 254.34
R947 GNDA.n2210 GNDA.n649 254.34
R948 GNDA.n2210 GNDA.n648 254.34
R949 GNDA.n2210 GNDA.n647 254.34
R950 GNDA.n2210 GNDA.n646 254.34
R951 GNDA.n2210 GNDA.n645 254.34
R952 GNDA.n2210 GNDA.n644 254.34
R953 GNDA.n2210 GNDA.n643 254.34
R954 GNDA.n1301 GNDA.n376 254.34
R955 GNDA.n1306 GNDA.n376 254.34
R956 GNDA.n1299 GNDA.n376 254.34
R957 GNDA.n1313 GNDA.n376 254.34
R958 GNDA.n1296 GNDA.n376 254.34
R959 GNDA.n1320 GNDA.n376 254.34
R960 GNDA.n1179 GNDA.n376 254.34
R961 GNDA.n1440 GNDA.n376 254.34
R962 GNDA.n1434 GNDA.n376 254.34
R963 GNDA.n1432 GNDA.n376 254.34
R964 GNDA.n1426 GNDA.n376 254.34
R965 GNDA.n1424 GNDA.n376 254.34
R966 GNDA.n1456 GNDA.n376 254.34
R967 GNDA.n1624 GNDA.n376 254.34
R968 GNDA.n1453 GNDA.n376 254.34
R969 GNDA.n1631 GNDA.n376 254.34
R970 GNDA.n1450 GNDA.n376 254.34
R971 GNDA.n1638 GNDA.n376 254.34
R972 GNDA.n2357 GNDA.n2356 254.34
R973 GNDA.n2357 GNDA.n575 254.34
R974 GNDA.n2357 GNDA.n574 254.34
R975 GNDA.n2357 GNDA.n573 254.34
R976 GNDA.n2357 GNDA.n572 254.34
R977 GNDA.n2357 GNDA.n571 254.34
R978 GNDA.n2357 GNDA.n570 254.34
R979 GNDA.n2357 GNDA.n456 254.34
R980 GNDA.n2357 GNDA.n455 254.34
R981 GNDA.n2357 GNDA.n454 254.34
R982 GNDA.n2357 GNDA.n453 254.34
R983 GNDA.n2357 GNDA.n452 254.34
R984 GNDA.n2358 GNDA.n2357 254.34
R985 GNDA.n2357 GNDA.n450 254.34
R986 GNDA.n2357 GNDA.n449 254.34
R987 GNDA.n2357 GNDA.n448 254.34
R988 GNDA.n2357 GNDA.n447 254.34
R989 GNDA.n2357 GNDA.n446 254.34
R990 GNDA.n1597 GNDA.n362 254.34
R991 GNDA.n1603 GNDA.n362 254.34
R992 GNDA.n1462 GNDA.n362 254.34
R993 GNDA.n1610 GNDA.n362 254.34
R994 GNDA.n1459 GNDA.n362 254.34
R995 GNDA.n1617 GNDA.n362 254.34
R996 GNDA.n802 GNDA.n362 254.34
R997 GNDA.n808 GNDA.n362 254.34
R998 GNDA.n691 GNDA.n362 254.34
R999 GNDA.n815 GNDA.n362 254.34
R1000 GNDA.n688 GNDA.n362 254.34
R1001 GNDA.n822 GNDA.n362 254.34
R1002 GNDA.n2015 GNDA.n362 254.34
R1003 GNDA.n2009 GNDA.n362 254.34
R1004 GNDA.n2007 GNDA.n362 254.34
R1005 GNDA.n2001 GNDA.n362 254.34
R1006 GNDA.n1999 GNDA.n362 254.34
R1007 GNDA.n1993 GNDA.n362 254.34
R1008 GNDA.n1762 GNDA.n1761 250.349
R1009 GNDA.n1681 GNDA.n1680 250.349
R1010 GNDA.n300 GNDA.n299 250.349
R1011 GNDA.n300 GNDA.n195 250.349
R1012 GNDA.n273 GNDA.n272 250.349
R1013 GNDA.n274 GNDA.n273 250.349
R1014 GNDA.n252 GNDA.n251 250.349
R1015 GNDA.n253 GNDA.n252 250.349
R1016 GNDA.n2489 GNDA.n107 250.349
R1017 GNDA.n1641 GNDA.n1639 249.663
R1018 GNDA.n1423 GNDA.n1185 249.663
R1019 GNDA.n910 GNDA.n871 249.663
R1020 GNDA.n2391 GNDA.n407 249.663
R1021 GNDA.n1970 GNDA.n1073 249.663
R1022 GNDA.n1902 GNDA.n1823 249.663
R1023 GNDA.n2235 GNDA.n639 249.663
R1024 GNDA.n611 GNDA.n610 249.663
R1025 GNDA.n1322 GNDA.n1321 249.663
R1026 GNDA.t10 GNDA.t309 248.206
R1027 GNDA.n2493 GNDA.n2492 248.206
R1028 GNDA.t185 GNDA.t55 248.206
R1029 GNDA.t294 GNDA.t97 248.206
R1030 GNDA.t202 GNDA.t45 248.206
R1031 GNDA.t269 GNDA.t18 248.206
R1032 GNDA.t136 GNDA.t115 248.206
R1033 GNDA.n2552 GNDA.n2549 247.934
R1034 GNDA.n2566 GNDA.n2544 247.934
R1035 GNDA.n2543 GNDA.n2542 247.934
R1036 GNDA.n2538 GNDA.n2537 247.934
R1037 GNDA.n2534 GNDA.n2533 247.934
R1038 GNDA.n2590 GNDA.n2530 247.934
R1039 GNDA.n2617 GNDA.n88 247.934
R1040 GNDA.n87 GNDA.n86 247.934
R1041 GNDA.n2637 GNDA.n78 247.934
R1042 GNDA.n77 GNDA.n76 247.934
R1043 GNDA.n2650 GNDA.n71 246.714
R1044 GNDA.n1786 GNDA.n1775 246.25
R1045 GNDA.n1778 GNDA.n1775 246.25
R1046 GNDA.n1805 GNDA.n1804 246.25
R1047 GNDA.n1804 GNDA.n1797 246.25
R1048 GNDA.n178 GNDA.t237 245
R1049 GNDA.n172 GNDA.t264 245
R1050 GNDA.n306 GNDA.t234 245
R1051 GNDA.n129 GNDA.t240 245
R1052 GNDA.n1097 GNDA.n1096 241.643
R1053 GNDA.n1806 GNDA.t173 241.643
R1054 GNDA.n1798 GNDA.t173 241.643
R1055 GNDA.n1787 GNDA.t107 241.643
R1056 GNDA.n1779 GNDA.t107 241.643
R1057 GNDA.n2763 GNDA.n2762 241.643
R1058 GNDA.n185 GNDA.n184 241.643
R1059 GNDA.n192 GNDA.n191 241.643
R1060 GNDA.t3 GNDA.n2770 236.923
R1061 GNDA.t62 GNDA.n106 236.078
R1062 GNDA.n2527 GNDA.t290 233
R1063 GNDA.n83 GNDA.t11 233
R1064 GNDA.n182 GNDA.t75 233
R1065 GNDA.n187 GNDA.t29 233
R1066 GNDA.n26 GNDA.t180 233
R1067 GNDA.t55 GNDA.t47 225.642
R1068 GNDA.n2526 GNDA.n2525 225.642
R1069 GNDA.n67 GNDA.n66 219.133
R1070 GNDA.n2662 GNDA.n65 219.133
R1071 GNDA.n61 GNDA.n60 219.133
R1072 GNDA.n56 GNDA.n55 219.133
R1073 GNDA.n2684 GNDA.n54 219.133
R1074 GNDA.n50 GNDA.n49 219.133
R1075 GNDA.n45 GNDA.n44 219.133
R1076 GNDA.n2706 GNDA.n43 219.133
R1077 GNDA.n39 GNDA.n38 219.133
R1078 GNDA.t211 GNDA.t181 218.802
R1079 GNDA.n2764 GNDA.t146 212.904
R1080 GNDA.n175 GNDA.n125 204.201
R1081 GNDA.n309 GNDA.n120 204.201
R1082 GNDA.n308 GNDA.n122 204.201
R1083 GNDA.n127 GNDA.n121 204.201
R1084 GNDA.n174 GNDA.n126 204.201
R1085 GNDA.n177 GNDA.n176 204.201
R1086 GNDA.t305 GNDA.t3 203.077
R1087 GNDA.t33 GNDA.t269 203.077
R1088 GNDA.t67 GNDA.t35 203.077
R1089 GNDA.t22 GNDA.t324 203.077
R1090 GNDA.n3 GNDA.t68 198.058
R1091 GNDA.n2814 GNDA.t19 198.058
R1092 GNDA.n2802 GNDA.t282 198.058
R1093 GNDA.n11 GNDA.t272 198.058
R1094 GNDA.n356 GNDA.t100 198.058
R1095 GNDA.n2416 GNDA.t70 198.058
R1096 GNDA.n2428 GNDA.t200 198.058
R1097 GNDA.n348 GNDA.t276 198.058
R1098 GNDA.n227 GNDA.n224 197
R1099 GNDA.n208 GNDA.n207 197
R1100 GNDA.n294 GNDA.n197 197
R1101 GNDA.n1673 GNDA.n1672 197
R1102 GNDA.n1760 GNDA.n1111 197
R1103 GNDA.n1596 GNDA.n1595 197
R1104 GNDA.n1669 GNDA.n1145 197
R1105 GNDA.n801 GNDA.n800 197
R1106 GNDA.n451 GNDA.n436 197
R1107 GNDA.n2018 GNDA.n2017 197
R1108 GNDA.n1032 GNDA.n684 197
R1109 GNDA.n2118 GNDA.n2117 197
R1110 GNDA.n2266 GNDA.n435 197
R1111 GNDA.n1394 GNDA.n1214 197
R1112 GNDA.n2488 GNDA.n109 197
R1113 GNDA.n2483 GNDA.n108 197
R1114 GNDA.t221 GNDA.n373 194.476
R1115 GNDA.n2772 GNDA.t6 191.796
R1116 GNDA.t313 GNDA.n1095 188.828
R1117 GNDA.n1555 GNDA.n1552 187.249
R1118 GNDA.n1397 GNDA.n1114 187.249
R1119 GNDA.n2366 GNDA.n438 187.249
R1120 GNDA.n2368 GNDA.n433 187.249
R1121 GNDA.n2115 GNDA.n914 187.249
R1122 GNDA.n993 GNDA.n683 187.249
R1123 GNDA.n2213 GNDA.n2212 187.249
R1124 GNDA.n2355 GNDA.n577 187.249
R1125 GNDA.n1346 GNDA.n1345 187.249
R1126 GNDA.n250 GNDA.n223 185
R1127 GNDA.n254 GNDA.n223 185
R1128 GNDA.n271 GNDA.n206 185
R1129 GNDA.n275 GNDA.n206 185
R1130 GNDA.n298 GNDA.n198 185
R1131 GNDA.n293 GNDA.n198 185
R1132 GNDA.n1788 GNDA.n1774 185
R1133 GNDA.n1781 GNDA.n1780 185
R1134 GNDA.n1807 GNDA.n1796 185
R1135 GNDA.n1803 GNDA.n1796 185
R1136 GNDA.n1807 GNDA.n1793 185
R1137 GNDA.n1799 GNDA.n1793 185
R1138 GNDA.n1723 GNDA.n1140 185
R1139 GNDA.n1738 GNDA.n1737 185
R1140 GNDA.n1736 GNDA.n1141 185
R1141 GNDA.n1735 GNDA.n1734 185
R1142 GNDA.n1733 GNDA.n1732 185
R1143 GNDA.n1731 GNDA.n1730 185
R1144 GNDA.n1729 GNDA.n1728 185
R1145 GNDA.n1727 GNDA.n1726 185
R1146 GNDA.n1725 GNDA.n1724 185
R1147 GNDA.n1706 GNDA.n1705 185
R1148 GNDA.n1708 GNDA.n1707 185
R1149 GNDA.n1710 GNDA.n1709 185
R1150 GNDA.n1712 GNDA.n1711 185
R1151 GNDA.n1714 GNDA.n1713 185
R1152 GNDA.n1716 GNDA.n1715 185
R1153 GNDA.n1718 GNDA.n1717 185
R1154 GNDA.n1720 GNDA.n1719 185
R1155 GNDA.n1722 GNDA.n1721 185
R1156 GNDA.n1688 GNDA.n1687 185
R1157 GNDA.n1690 GNDA.n1689 185
R1158 GNDA.n1692 GNDA.n1691 185
R1159 GNDA.n1694 GNDA.n1693 185
R1160 GNDA.n1696 GNDA.n1695 185
R1161 GNDA.n1698 GNDA.n1697 185
R1162 GNDA.n1700 GNDA.n1699 185
R1163 GNDA.n1702 GNDA.n1701 185
R1164 GNDA.n1704 GNDA.n1703 185
R1165 GNDA.n1534 GNDA.n1533 185
R1166 GNDA.n1536 GNDA.n1535 185
R1167 GNDA.n1538 GNDA.n1537 185
R1168 GNDA.n1540 GNDA.n1539 185
R1169 GNDA.n1542 GNDA.n1541 185
R1170 GNDA.n1544 GNDA.n1543 185
R1171 GNDA.n1546 GNDA.n1545 185
R1172 GNDA.n1548 GNDA.n1547 185
R1173 GNDA.n1549 GNDA.n1490 185
R1174 GNDA.n1516 GNDA.n1515 185
R1175 GNDA.n1518 GNDA.n1517 185
R1176 GNDA.n1520 GNDA.n1519 185
R1177 GNDA.n1522 GNDA.n1521 185
R1178 GNDA.n1524 GNDA.n1523 185
R1179 GNDA.n1526 GNDA.n1525 185
R1180 GNDA.n1528 GNDA.n1527 185
R1181 GNDA.n1530 GNDA.n1529 185
R1182 GNDA.n1532 GNDA.n1531 185
R1183 GNDA.n1498 GNDA.n1497 185
R1184 GNDA.n1500 GNDA.n1499 185
R1185 GNDA.n1502 GNDA.n1501 185
R1186 GNDA.n1504 GNDA.n1503 185
R1187 GNDA.n1506 GNDA.n1505 185
R1188 GNDA.n1508 GNDA.n1507 185
R1189 GNDA.n1510 GNDA.n1509 185
R1190 GNDA.n1512 GNDA.n1511 185
R1191 GNDA.n1514 GNDA.n1513 185
R1192 GNDA.n1473 GNDA.n1472 185
R1193 GNDA.n1588 GNDA.n1587 185
R1194 GNDA.n1471 GNDA.n1469 185
R1195 GNDA.n1569 GNDA.n1568 185
R1196 GNDA.n1571 GNDA.n1570 185
R1197 GNDA.n1575 GNDA.n1574 185
R1198 GNDA.n1573 GNDA.n1564 185
R1199 GNDA.n1493 GNDA.n1491 185
R1200 GNDA.n1584 GNDA.n1583 185
R1201 GNDA.n1686 GNDA.n1685 185
R1202 GNDA.n1156 GNDA.n1155 185
R1203 GNDA.n1158 GNDA.n1157 185
R1204 GNDA.n1153 GNDA.n1125 185
R1205 GNDA.n1744 GNDA.n1743 185
R1206 GNDA.n1741 GNDA.n1124 185
R1207 GNDA.n1740 GNDA.n1120 185
R1208 GNDA.n1753 GNDA.n1752 185
R1209 GNDA.n1755 GNDA.n1754 185
R1210 GNDA.n540 GNDA.n481 185
R1211 GNDA.n555 GNDA.n554 185
R1212 GNDA.n553 GNDA.n482 185
R1213 GNDA.n552 GNDA.n551 185
R1214 GNDA.n550 GNDA.n549 185
R1215 GNDA.n548 GNDA.n547 185
R1216 GNDA.n546 GNDA.n545 185
R1217 GNDA.n544 GNDA.n543 185
R1218 GNDA.n542 GNDA.n541 185
R1219 GNDA.n523 GNDA.n522 185
R1220 GNDA.n525 GNDA.n524 185
R1221 GNDA.n527 GNDA.n526 185
R1222 GNDA.n529 GNDA.n528 185
R1223 GNDA.n531 GNDA.n530 185
R1224 GNDA.n533 GNDA.n532 185
R1225 GNDA.n535 GNDA.n534 185
R1226 GNDA.n537 GNDA.n536 185
R1227 GNDA.n539 GNDA.n538 185
R1228 GNDA.n505 GNDA.n504 185
R1229 GNDA.n507 GNDA.n506 185
R1230 GNDA.n509 GNDA.n508 185
R1231 GNDA.n511 GNDA.n510 185
R1232 GNDA.n513 GNDA.n512 185
R1233 GNDA.n515 GNDA.n514 185
R1234 GNDA.n517 GNDA.n516 185
R1235 GNDA.n519 GNDA.n518 185
R1236 GNDA.n521 GNDA.n520 185
R1237 GNDA.n503 GNDA.n502 185
R1238 GNDA.n497 GNDA.n496 185
R1239 GNDA.n495 GNDA.n494 185
R1240 GNDA.n490 GNDA.n489 185
R1241 GNDA.n485 GNDA.n466 185
R1242 GNDA.n559 GNDA.n558 185
R1243 GNDA.n465 GNDA.n463 185
R1244 GNDA.n565 GNDA.n564 185
R1245 GNDA.n567 GNDA.n566 185
R1246 GNDA.n750 GNDA.n749 185
R1247 GNDA.n752 GNDA.n751 185
R1248 GNDA.n754 GNDA.n753 185
R1249 GNDA.n756 GNDA.n755 185
R1250 GNDA.n758 GNDA.n757 185
R1251 GNDA.n760 GNDA.n759 185
R1252 GNDA.n762 GNDA.n761 185
R1253 GNDA.n764 GNDA.n763 185
R1254 GNDA.n765 GNDA.n443 185
R1255 GNDA.n732 GNDA.n731 185
R1256 GNDA.n734 GNDA.n733 185
R1257 GNDA.n736 GNDA.n735 185
R1258 GNDA.n738 GNDA.n737 185
R1259 GNDA.n740 GNDA.n739 185
R1260 GNDA.n742 GNDA.n741 185
R1261 GNDA.n744 GNDA.n743 185
R1262 GNDA.n746 GNDA.n745 185
R1263 GNDA.n748 GNDA.n747 185
R1264 GNDA.n707 GNDA.n693 185
R1265 GNDA.n716 GNDA.n715 185
R1266 GNDA.n718 GNDA.n717 185
R1267 GNDA.n720 GNDA.n719 185
R1268 GNDA.n722 GNDA.n721 185
R1269 GNDA.n724 GNDA.n723 185
R1270 GNDA.n726 GNDA.n725 185
R1271 GNDA.n728 GNDA.n727 185
R1272 GNDA.n730 GNDA.n729 185
R1273 GNDA.n697 GNDA.n694 185
R1274 GNDA.n793 GNDA.n792 185
R1275 GNDA.n769 GNDA.n696 185
R1276 GNDA.n775 GNDA.n774 185
R1277 GNDA.n773 GNDA.n768 185
R1278 GNDA.n782 GNDA.n781 185
R1279 GNDA.n780 GNDA.n767 185
R1280 GNDA.n788 GNDA.n787 185
R1281 GNDA.n789 GNDA.n444 185
R1282 GNDA.n977 GNDA.n976 185
R1283 GNDA.n979 GNDA.n978 185
R1284 GNDA.n981 GNDA.n980 185
R1285 GNDA.n983 GNDA.n982 185
R1286 GNDA.n985 GNDA.n984 185
R1287 GNDA.n987 GNDA.n986 185
R1288 GNDA.n989 GNDA.n988 185
R1289 GNDA.n991 GNDA.n990 185
R1290 GNDA.n992 GNDA.n940 185
R1291 GNDA.n959 GNDA.n958 185
R1292 GNDA.n961 GNDA.n960 185
R1293 GNDA.n963 GNDA.n962 185
R1294 GNDA.n965 GNDA.n964 185
R1295 GNDA.n967 GNDA.n966 185
R1296 GNDA.n969 GNDA.n968 185
R1297 GNDA.n971 GNDA.n970 185
R1298 GNDA.n973 GNDA.n972 185
R1299 GNDA.n975 GNDA.n974 185
R1300 GNDA.n932 GNDA.n918 185
R1301 GNDA.n943 GNDA.n942 185
R1302 GNDA.n945 GNDA.n944 185
R1303 GNDA.n947 GNDA.n946 185
R1304 GNDA.n949 GNDA.n948 185
R1305 GNDA.n951 GNDA.n950 185
R1306 GNDA.n953 GNDA.n952 185
R1307 GNDA.n955 GNDA.n954 185
R1308 GNDA.n957 GNDA.n956 185
R1309 GNDA.n922 GNDA.n919 185
R1310 GNDA.n1026 GNDA.n1025 185
R1311 GNDA.n999 GNDA.n921 185
R1312 GNDA.n1005 GNDA.n1004 185
R1313 GNDA.n1003 GNDA.n998 185
R1314 GNDA.n1012 GNDA.n1011 185
R1315 GNDA.n1010 GNDA.n997 185
R1316 GNDA.n1017 GNDA.n941 185
R1317 GNDA.n1022 GNDA.n1021 185
R1318 GNDA.n2185 GNDA.n2184 185
R1319 GNDA.n2187 GNDA.n2186 185
R1320 GNDA.n2189 GNDA.n2188 185
R1321 GNDA.n2191 GNDA.n2190 185
R1322 GNDA.n2193 GNDA.n2192 185
R1323 GNDA.n2195 GNDA.n2194 185
R1324 GNDA.n2197 GNDA.n2196 185
R1325 GNDA.n2198 GNDA.n680 185
R1326 GNDA.n2202 GNDA.n2201 185
R1327 GNDA.n2167 GNDA.n2166 185
R1328 GNDA.n2169 GNDA.n2168 185
R1329 GNDA.n2171 GNDA.n2170 185
R1330 GNDA.n2173 GNDA.n2172 185
R1331 GNDA.n2175 GNDA.n2174 185
R1332 GNDA.n2177 GNDA.n2176 185
R1333 GNDA.n2179 GNDA.n2178 185
R1334 GNDA.n2181 GNDA.n2180 185
R1335 GNDA.n2183 GNDA.n2182 185
R1336 GNDA.n2149 GNDA.n2148 185
R1337 GNDA.n2151 GNDA.n2150 185
R1338 GNDA.n2153 GNDA.n2152 185
R1339 GNDA.n2155 GNDA.n2154 185
R1340 GNDA.n2157 GNDA.n2156 185
R1341 GNDA.n2159 GNDA.n2158 185
R1342 GNDA.n2161 GNDA.n2160 185
R1343 GNDA.n2163 GNDA.n2162 185
R1344 GNDA.n2165 GNDA.n2164 185
R1345 GNDA.n2147 GNDA.n2146 185
R1346 GNDA.n2141 GNDA.n2140 185
R1347 GNDA.n2139 GNDA.n2138 185
R1348 GNDA.n2134 GNDA.n2133 185
R1349 GNDA.n2132 GNDA.n2131 185
R1350 GNDA.n2126 GNDA.n2125 185
R1351 GNDA.n2122 GNDA.n663 185
R1352 GNDA.n2206 GNDA.n2205 185
R1353 GNDA.n662 GNDA.n660 185
R1354 GNDA.n2325 GNDA.n2264 185
R1355 GNDA.n2339 GNDA.n2338 185
R1356 GNDA.n2337 GNDA.n2265 185
R1357 GNDA.n2336 GNDA.n2335 185
R1358 GNDA.n2334 GNDA.n2333 185
R1359 GNDA.n2332 GNDA.n2331 185
R1360 GNDA.n2330 GNDA.n2329 185
R1361 GNDA.n2328 GNDA.n2327 185
R1362 GNDA.n2326 GNDA.n2241 185
R1363 GNDA.n2308 GNDA.n2307 185
R1364 GNDA.n2310 GNDA.n2309 185
R1365 GNDA.n2312 GNDA.n2311 185
R1366 GNDA.n2314 GNDA.n2313 185
R1367 GNDA.n2316 GNDA.n2315 185
R1368 GNDA.n2318 GNDA.n2317 185
R1369 GNDA.n2320 GNDA.n2319 185
R1370 GNDA.n2322 GNDA.n2321 185
R1371 GNDA.n2324 GNDA.n2323 185
R1372 GNDA.n2290 GNDA.n2289 185
R1373 GNDA.n2292 GNDA.n2291 185
R1374 GNDA.n2294 GNDA.n2293 185
R1375 GNDA.n2296 GNDA.n2295 185
R1376 GNDA.n2298 GNDA.n2297 185
R1377 GNDA.n2300 GNDA.n2299 185
R1378 GNDA.n2302 GNDA.n2301 185
R1379 GNDA.n2304 GNDA.n2303 185
R1380 GNDA.n2306 GNDA.n2305 185
R1381 GNDA.n2288 GNDA.n2287 185
R1382 GNDA.n2282 GNDA.n2281 185
R1383 GNDA.n2280 GNDA.n2279 185
R1384 GNDA.n2275 GNDA.n2274 185
R1385 GNDA.n2270 GNDA.n2249 185
R1386 GNDA.n2343 GNDA.n2342 185
R1387 GNDA.n2248 GNDA.n2246 185
R1388 GNDA.n2349 GNDA.n2348 185
R1389 GNDA.n2351 GNDA.n2350 185
R1390 GNDA.n1278 GNDA.n1277 185
R1391 GNDA.n1280 GNDA.n1235 185
R1392 GNDA.n1283 GNDA.n1282 185
R1393 GNDA.n1284 GNDA.n1234 185
R1394 GNDA.n1286 GNDA.n1285 185
R1395 GNDA.n1288 GNDA.n1233 185
R1396 GNDA.n1291 GNDA.n1290 185
R1397 GNDA.n1292 GNDA.n1232 185
R1398 GNDA.n1351 GNDA.n1350 185
R1399 GNDA.n1260 GNDA.n1240 185
R1400 GNDA.n1262 GNDA.n1261 185
R1401 GNDA.n1264 GNDA.n1239 185
R1402 GNDA.n1267 GNDA.n1266 185
R1403 GNDA.n1268 GNDA.n1238 185
R1404 GNDA.n1270 GNDA.n1269 185
R1405 GNDA.n1272 GNDA.n1237 185
R1406 GNDA.n1275 GNDA.n1274 185
R1407 GNDA.n1276 GNDA.n1236 185
R1408 GNDA.n1386 GNDA.n1385 185
R1409 GNDA.n1245 GNDA.n1217 185
R1410 GNDA.n1247 GNDA.n1246 185
R1411 GNDA.n1249 GNDA.n1243 185
R1412 GNDA.n1251 GNDA.n1250 185
R1413 GNDA.n1252 GNDA.n1242 185
R1414 GNDA.n1254 GNDA.n1253 185
R1415 GNDA.n1256 GNDA.n1241 185
R1416 GNDA.n1259 GNDA.n1258 185
R1417 GNDA.n1384 GNDA.n1216 185
R1418 GNDA.n1382 GNDA.n1381 185
R1419 GNDA.n1220 GNDA.n1219 185
R1420 GNDA.n1371 GNDA.n1370 185
R1421 GNDA.n1368 GNDA.n1224 185
R1422 GNDA.n1366 GNDA.n1365 185
R1423 GNDA.n1226 GNDA.n1225 185
R1424 GNDA.n1356 GNDA.n1355 185
R1425 GNDA.n1353 GNDA.n1230 185
R1426 GNDA.n2086 GNDA.n2085 185
R1427 GNDA.n2088 GNDA.n2087 185
R1428 GNDA.n2090 GNDA.n2089 185
R1429 GNDA.n2092 GNDA.n2091 185
R1430 GNDA.n2094 GNDA.n2093 185
R1431 GNDA.n2096 GNDA.n2095 185
R1432 GNDA.n2098 GNDA.n2097 185
R1433 GNDA.n2100 GNDA.n2099 185
R1434 GNDA.n2101 GNDA.n1034 185
R1435 GNDA.n2068 GNDA.n2067 185
R1436 GNDA.n2070 GNDA.n2069 185
R1437 GNDA.n2072 GNDA.n2071 185
R1438 GNDA.n2074 GNDA.n2073 185
R1439 GNDA.n2076 GNDA.n2075 185
R1440 GNDA.n2078 GNDA.n2077 185
R1441 GNDA.n2080 GNDA.n2079 185
R1442 GNDA.n2082 GNDA.n2081 185
R1443 GNDA.n2084 GNDA.n2083 185
R1444 GNDA.n2050 GNDA.n2049 185
R1445 GNDA.n2052 GNDA.n2051 185
R1446 GNDA.n2054 GNDA.n2053 185
R1447 GNDA.n2056 GNDA.n2055 185
R1448 GNDA.n2058 GNDA.n2057 185
R1449 GNDA.n2060 GNDA.n2059 185
R1450 GNDA.n2062 GNDA.n2061 185
R1451 GNDA.n2064 GNDA.n2063 185
R1452 GNDA.n2066 GNDA.n2065 185
R1453 GNDA.n2048 GNDA.n2047 185
R1454 GNDA.n2042 GNDA.n2041 185
R1455 GNDA.n2040 GNDA.n2039 185
R1456 GNDA.n2035 GNDA.n2034 185
R1457 GNDA.n2033 GNDA.n2032 185
R1458 GNDA.n2027 GNDA.n2026 185
R1459 GNDA.n2022 GNDA.n1038 185
R1460 GNDA.n2105 GNDA.n2104 185
R1461 GNDA.n1037 GNDA.n1035 185
R1462 GNDA.n2487 GNDA.n110 185
R1463 GNDA.n2482 GNDA.n110 185
R1464 GNDA.t44 GNDA.t63 181.956
R1465 GNDA.t204 GNDA.t77 181.956
R1466 GNDA.t42 GNDA.t151 181.956
R1467 GNDA.t131 GNDA.t189 181.956
R1468 GNDA.t112 GNDA.t139 181.956
R1469 GNDA.t285 GNDA.t175 181.956
R1470 GNDA.t57 GNDA.t110 181.956
R1471 GNDA.t197 GNDA.t95 181.956
R1472 GNDA.t159 GNDA.t197 181.956
R1473 GNDA.t326 GNDA.t143 180.513
R1474 GNDA.t310 GNDA.t185 180.513
R1475 GNDA.n1616 GNDA.n1457 175.546
R1476 GNDA.n1612 GNDA.n1611 175.546
R1477 GNDA.n1609 GNDA.n1460 175.546
R1478 GNDA.n1605 GNDA.n1604 175.546
R1479 GNDA.n1602 GNDA.n1463 175.546
R1480 GNDA.n1637 GNDA.n1448 175.546
R1481 GNDA.n1633 GNDA.n1632 175.546
R1482 GNDA.n1630 GNDA.n1451 175.546
R1483 GNDA.n1626 GNDA.n1625 175.546
R1484 GNDA.n1623 GNDA.n1454 175.546
R1485 GNDA.n1559 GNDA.n1552 175.546
R1486 GNDA.n1581 GNDA.n1559 175.546
R1487 GNDA.n1581 GNDA.n1560 175.546
R1488 GNDA.n1577 GNDA.n1560 175.546
R1489 GNDA.n1577 GNDA.n1562 175.546
R1490 GNDA.n1565 GNDA.n1562 175.546
R1491 GNDA.n1565 GNDA.n1468 175.546
R1492 GNDA.n1590 GNDA.n1468 175.546
R1493 GNDA.n1590 GNDA.n1465 175.546
R1494 GNDA.n1594 GNDA.n1465 175.546
R1495 GNDA.n1595 GNDA.n1594 175.546
R1496 GNDA.n1647 GNDA.n1177 175.546
R1497 GNDA.n1651 GNDA.n1649 175.546
R1498 GNDA.n1657 GNDA.n1173 175.546
R1499 GNDA.n1660 GNDA.n1659 175.546
R1500 GNDA.n1662 GNDA.n1170 175.546
R1501 GNDA.n1418 GNDA.n1191 175.546
R1502 GNDA.n1414 GNDA.n1196 175.546
R1503 GNDA.n1410 GNDA.n1409 175.546
R1504 GNDA.n1406 GNDA.n1405 175.546
R1505 GNDA.n1402 GNDA.n1401 175.546
R1506 GNDA.n1427 GNDA.n1425 175.546
R1507 GNDA.n1431 GNDA.n1183 175.546
R1508 GNDA.n1435 GNDA.n1433 175.546
R1509 GNDA.n1439 GNDA.n1181 175.546
R1510 GNDA.n1442 GNDA.n1441 175.546
R1511 GNDA.n1757 GNDA.n1114 175.546
R1512 GNDA.n1757 GNDA.n1115 175.546
R1513 GNDA.n1750 GNDA.n1115 175.546
R1514 GNDA.n1750 GNDA.n1121 175.546
R1515 GNDA.n1746 GNDA.n1121 175.546
R1516 GNDA.n1746 GNDA.n1122 175.546
R1517 GNDA.n1160 GNDA.n1122 175.546
R1518 GNDA.n1160 GNDA.n1151 175.546
R1519 GNDA.n1151 GNDA.n1144 175.546
R1520 GNDA.n1683 GNDA.n1144 175.546
R1521 GNDA.n1683 GNDA.n1145 175.546
R1522 GNDA.n1645 GNDA.n1644 175.546
R1523 GNDA.n1176 GNDA.n1175 175.546
R1524 GNDA.n1655 GNDA.n1654 175.546
R1525 GNDA.n1171 GNDA.n1167 175.546
R1526 GNDA.n1664 GNDA.n1149 175.546
R1527 GNDA.n821 GNDA.n686 175.546
R1528 GNDA.n817 GNDA.n816 175.546
R1529 GNDA.n814 GNDA.n689 175.546
R1530 GNDA.n810 GNDA.n809 175.546
R1531 GNDA.n807 GNDA.n692 175.546
R1532 GNDA.n844 GNDA.n843 175.546
R1533 GNDA.n840 GNDA.n839 175.546
R1534 GNDA.n836 GNDA.n835 175.546
R1535 GNDA.n832 GNDA.n831 175.546
R1536 GNDA.n828 GNDA.n827 175.546
R1537 GNDA.n2359 GNDA.n445 175.546
R1538 GNDA.n785 GNDA.n784 175.546
R1539 GNDA.n778 GNDA.n777 175.546
R1540 GNDA.n771 GNDA.n770 175.546
R1541 GNDA.n796 GNDA.n795 175.546
R1542 GNDA.n908 GNDA.n907 175.546
R1543 GNDA.n907 GNDA.n872 175.546
R1544 GNDA.n903 GNDA.n901 175.546
R1545 GNDA.n899 GNDA.n880 175.546
R1546 GNDA.n895 GNDA.n893 175.546
R1547 GNDA.n2365 GNDA.n439 175.546
R1548 GNDA.n2387 GNDA.n408 175.546
R1549 GNDA.n2383 GNDA.n413 175.546
R1550 GNDA.n2381 GNDA.n2380 175.546
R1551 GNDA.n2377 GNDA.n2376 175.546
R1552 GNDA.n2373 GNDA.n2372 175.546
R1553 GNDA.n849 GNDA.n848 175.546
R1554 GNDA.n853 GNDA.n852 175.546
R1555 GNDA.n857 GNDA.n856 175.546
R1556 GNDA.n861 GNDA.n860 175.546
R1557 GNDA.n865 GNDA.n864 175.546
R1558 GNDA.n569 GNDA.n457 175.546
R1559 GNDA.n562 GNDA.n561 175.546
R1560 GNDA.n487 GNDA.n486 175.546
R1561 GNDA.n492 GNDA.n491 175.546
R1562 GNDA.n500 GNDA.n499 175.546
R1563 GNDA.n875 GNDA.n874 175.546
R1564 GNDA.n878 GNDA.n877 175.546
R1565 GNDA.n883 GNDA.n882 175.546
R1566 GNDA.n886 GNDA.n885 175.546
R1567 GNDA.n890 GNDA.n888 175.546
R1568 GNDA.n1998 GNDA.n1060 175.546
R1569 GNDA.n2002 GNDA.n2000 175.546
R1570 GNDA.n2006 GNDA.n1058 175.546
R1571 GNDA.n2010 GNDA.n2008 175.546
R1572 GNDA.n2014 GNDA.n1056 175.546
R1573 GNDA.n1970 GNDA.n1071 175.546
R1574 GNDA.n1974 GNDA.n1071 175.546
R1575 GNDA.n1974 GNDA.n1069 175.546
R1576 GNDA.n1978 GNDA.n1069 175.546
R1577 GNDA.n1978 GNDA.n1067 175.546
R1578 GNDA.n1982 GNDA.n1067 175.546
R1579 GNDA.n1982 GNDA.n1065 175.546
R1580 GNDA.n1987 GNDA.n1065 175.546
R1581 GNDA.n1987 GNDA.n1062 175.546
R1582 GNDA.n1991 GNDA.n1062 175.546
R1583 GNDA.n1992 GNDA.n1991 175.546
R1584 GNDA.n2108 GNDA.n2107 175.546
R1585 GNDA.n2024 GNDA.n2023 175.546
R1586 GNDA.n2030 GNDA.n2029 175.546
R1587 GNDA.n2037 GNDA.n2036 175.546
R1588 GNDA.n2045 GNDA.n2044 175.546
R1589 GNDA.n1965 GNDA.n1073 175.546
R1590 GNDA.n1965 GNDA.n1932 175.546
R1591 GNDA.n1961 GNDA.n1932 175.546
R1592 GNDA.n1961 GNDA.n1937 175.546
R1593 GNDA.n1957 GNDA.n1937 175.546
R1594 GNDA.n1957 GNDA.n1956 175.546
R1595 GNDA.n1956 GNDA.n1955 175.546
R1596 GNDA.n1955 GNDA.n1941 175.546
R1597 GNDA.n1951 GNDA.n1941 175.546
R1598 GNDA.n1951 GNDA.n915 175.546
R1599 GNDA.n2114 GNDA.n915 175.546
R1600 GNDA.n1865 GNDA.n1823 175.546
R1601 GNDA.n1865 GNDA.n1829 175.546
R1602 GNDA.n1861 GNDA.n1829 175.546
R1603 GNDA.n1861 GNDA.n1833 175.546
R1604 GNDA.n1857 GNDA.n1833 175.546
R1605 GNDA.n1857 GNDA.n1856 175.546
R1606 GNDA.n1856 GNDA.n1855 175.546
R1607 GNDA.n1855 GNDA.n1837 175.546
R1608 GNDA.n1851 GNDA.n1837 175.546
R1609 GNDA.n1851 GNDA.n1844 175.546
R1610 GNDA.n1847 GNDA.n1844 175.546
R1611 GNDA.n1902 GNDA.n1821 175.546
R1612 GNDA.n1907 GNDA.n1821 175.546
R1613 GNDA.n1907 GNDA.n1819 175.546
R1614 GNDA.n1911 GNDA.n1819 175.546
R1615 GNDA.n1912 GNDA.n1911 175.546
R1616 GNDA.n1912 GNDA.n1079 175.546
R1617 GNDA.n1919 GNDA.n1079 175.546
R1618 GNDA.n1919 GNDA.n1077 175.546
R1619 GNDA.n1924 GNDA.n1077 175.546
R1620 GNDA.n1924 GNDA.n1075 175.546
R1621 GNDA.n1928 GNDA.n1075 175.546
R1622 GNDA.n1019 GNDA.n1018 175.546
R1623 GNDA.n1015 GNDA.n1014 175.546
R1624 GNDA.n1008 GNDA.n1007 175.546
R1625 GNDA.n1001 GNDA.n1000 175.546
R1626 GNDA.n1029 GNDA.n1028 175.546
R1627 GNDA.n1930 GNDA.n1929 175.546
R1628 GNDA.n1934 GNDA.n1930 175.546
R1629 GNDA.n1935 GNDA.n1934 175.546
R1630 GNDA.n1938 GNDA.n1935 175.546
R1631 GNDA.n1939 GNDA.n1938 175.546
R1632 GNDA.n1943 GNDA.n1939 175.546
R1633 GNDA.n1944 GNDA.n1943 175.546
R1634 GNDA.n1945 GNDA.n1944 175.546
R1635 GNDA.n1946 GNDA.n1945 175.546
R1636 GNDA.n1947 GNDA.n1946 175.546
R1637 GNDA.n1947 GNDA.n917 175.546
R1638 GNDA.n1868 GNDA.n1827 175.546
R1639 GNDA.n1830 GNDA.n1827 175.546
R1640 GNDA.n1831 GNDA.n1830 175.546
R1641 GNDA.n1834 GNDA.n1831 175.546
R1642 GNDA.n1835 GNDA.n1834 175.546
R1643 GNDA.n1839 GNDA.n1835 175.546
R1644 GNDA.n1840 GNDA.n1839 175.546
R1645 GNDA.n1841 GNDA.n1840 175.546
R1646 GNDA.n1842 GNDA.n1841 175.546
R1647 GNDA.n1846 GNDA.n1842 175.546
R1648 GNDA.n1846 GNDA.n682 175.546
R1649 GNDA.n1878 GNDA.n639 175.546
R1650 GNDA.n1878 GNDA.n1876 175.546
R1651 GNDA.n1882 GNDA.n1876 175.546
R1652 GNDA.n1882 GNDA.n1874 175.546
R1653 GNDA.n1886 GNDA.n1874 175.546
R1654 GNDA.n1886 GNDA.n1872 175.546
R1655 GNDA.n1890 GNDA.n1872 175.546
R1656 GNDA.n1890 GNDA.n1870 175.546
R1657 GNDA.n1894 GNDA.n1870 175.546
R1658 GNDA.n1894 GNDA.n1826 175.546
R1659 GNDA.n1898 GNDA.n1826 175.546
R1660 GNDA.n2208 GNDA.n642 175.546
R1661 GNDA.n2123 GNDA.n659 175.546
R1662 GNDA.n2129 GNDA.n2128 175.546
R1663 GNDA.n2136 GNDA.n2135 175.546
R1664 GNDA.n2144 GNDA.n2143 175.546
R1665 GNDA.n638 GNDA.n637 175.546
R1666 GNDA.n2230 GNDA.n637 175.546
R1667 GNDA.n2228 GNDA.n2227 175.546
R1668 GNDA.n2224 GNDA.n2223 175.546
R1669 GNDA.n2220 GNDA.n2219 175.546
R1670 GNDA.n2216 GNDA.n2215 175.546
R1671 GNDA.n423 GNDA.n414 175.546
R1672 GNDA.n416 GNDA.n415 175.546
R1673 GNDA.n418 GNDA.n417 175.546
R1674 GNDA.n420 GNDA.n419 175.546
R1675 GNDA.n422 GNDA.n421 175.546
R1676 GNDA.n607 GNDA.n606 175.546
R1677 GNDA.n603 GNDA.n602 175.546
R1678 GNDA.n599 GNDA.n598 175.546
R1679 GNDA.n595 GNDA.n594 175.546
R1680 GNDA.n591 GNDA.n401 175.546
R1681 GNDA.n2242 GNDA.n576 175.546
R1682 GNDA.n2346 GNDA.n2345 175.546
R1683 GNDA.n2272 GNDA.n2271 175.546
R1684 GNDA.n2277 GNDA.n2276 175.546
R1685 GNDA.n2285 GNDA.n2284 175.546
R1686 GNDA.n615 GNDA.n614 175.546
R1687 GNDA.n619 GNDA.n618 175.546
R1688 GNDA.n623 GNDA.n622 175.546
R1689 GNDA.n628 GNDA.n590 175.546
R1690 GNDA.n589 GNDA.n579 175.546
R1691 GNDA.n2239 GNDA.n579 175.546
R1692 GNDA.n1197 GNDA.n1189 175.546
R1693 GNDA.n1200 GNDA.n1199 175.546
R1694 GNDA.n1203 GNDA.n1202 175.546
R1695 GNDA.n1206 GNDA.n1205 175.546
R1696 GNDA.n1209 GNDA.n1208 175.546
R1697 GNDA.n1319 GNDA.n1294 175.546
R1698 GNDA.n1315 GNDA.n1314 175.546
R1699 GNDA.n1312 GNDA.n1297 175.546
R1700 GNDA.n1308 GNDA.n1307 175.546
R1701 GNDA.n1305 GNDA.n1302 175.546
R1702 GNDA.n1346 GNDA.n1229 175.546
R1703 GNDA.n1358 GNDA.n1229 175.546
R1704 GNDA.n1358 GNDA.n1227 175.546
R1705 GNDA.n1362 GNDA.n1227 175.546
R1706 GNDA.n1362 GNDA.n1222 175.546
R1707 GNDA.n1373 GNDA.n1222 175.546
R1708 GNDA.n1373 GNDA.n1221 175.546
R1709 GNDA.n1378 GNDA.n1221 175.546
R1710 GNDA.n1378 GNDA.n1215 175.546
R1711 GNDA.n1390 GNDA.n1215 175.546
R1712 GNDA.n1390 GNDA.n1214 175.546
R1713 GNDA.n1326 GNDA.n1325 175.546
R1714 GNDA.n1330 GNDA.n1329 175.546
R1715 GNDA.n1334 GNDA.n1333 175.546
R1716 GNDA.n1338 GNDA.n1337 175.546
R1717 GNDA.n1340 GNDA.n631 175.546
R1718 GNDA.n1343 GNDA.n631 175.546
R1719 GNDA.n429 GNDA.n363 173.881
R1720 GNDA.t221 GNDA.n366 172.876
R1721 GNDA.t221 GNDA.n383 172.615
R1722 GNDA.n2389 GNDA.n363 171.624
R1723 GNDA.n2746 GNDA.n2745 171.494
R1724 GNDA.n250 GNDA.n228 166.63
R1725 GNDA.n271 GNDA.n209 166.63
R1726 GNDA.n1687 GNDA.n1686 163.333
R1727 GNDA.n1497 GNDA.n1473 163.333
R1728 GNDA.n504 GNDA.n503 163.333
R1729 GNDA.n707 GNDA.n697 163.333
R1730 GNDA.n932 GNDA.n922 163.333
R1731 GNDA.n2148 GNDA.n2147 163.333
R1732 GNDA.n2289 GNDA.n2288 163.333
R1733 GNDA.n1385 GNDA.n1384 163.333
R1734 GNDA.n2049 GNDA.n2048 163.333
R1735 GNDA.t221 GNDA.n367 162.064
R1736 GNDA.t37 GNDA.t301 157.95
R1737 GNDA.t141 GNDA.t271 157.95
R1738 GNDA.t281 GNDA.t7 157.95
R1739 GNDA.t132 GNDA.t79 157.95
R1740 GNDA.n1916 GNDA.n1082 157.601
R1741 GNDA.t267 GNDA.t285 157.143
R1742 GNDA.n1719 GNDA.n1718 150
R1743 GNDA.n1715 GNDA.n1714 150
R1744 GNDA.n1711 GNDA.n1710 150
R1745 GNDA.n1707 GNDA.n1706 150
R1746 GNDA.n1703 GNDA.n1702 150
R1747 GNDA.n1699 GNDA.n1698 150
R1748 GNDA.n1695 GNDA.n1694 150
R1749 GNDA.n1691 GNDA.n1690 150
R1750 GNDA.n1754 GNDA.n1753 150
R1751 GNDA.n1741 GNDA.n1740 150
R1752 GNDA.n1743 GNDA.n1125 150
R1753 GNDA.n1157 GNDA.n1156 150
R1754 GNDA.n1738 GNDA.n1141 150
R1755 GNDA.n1734 GNDA.n1733 150
R1756 GNDA.n1730 GNDA.n1729 150
R1757 GNDA.n1726 GNDA.n1725 150
R1758 GNDA.n1529 GNDA.n1528 150
R1759 GNDA.n1525 GNDA.n1524 150
R1760 GNDA.n1521 GNDA.n1520 150
R1761 GNDA.n1517 GNDA.n1516 150
R1762 GNDA.n1513 GNDA.n1512 150
R1763 GNDA.n1509 GNDA.n1508 150
R1764 GNDA.n1505 GNDA.n1504 150
R1765 GNDA.n1501 GNDA.n1500 150
R1766 GNDA.n1584 GNDA.n1491 150
R1767 GNDA.n1574 GNDA.n1573 150
R1768 GNDA.n1570 GNDA.n1569 150
R1769 GNDA.n1587 GNDA.n1471 150
R1770 GNDA.n1537 GNDA.n1536 150
R1771 GNDA.n1541 GNDA.n1540 150
R1772 GNDA.n1545 GNDA.n1544 150
R1773 GNDA.n1547 GNDA.n1490 150
R1774 GNDA.n536 GNDA.n535 150
R1775 GNDA.n532 GNDA.n531 150
R1776 GNDA.n528 GNDA.n527 150
R1777 GNDA.n524 GNDA.n523 150
R1778 GNDA.n520 GNDA.n519 150
R1779 GNDA.n516 GNDA.n515 150
R1780 GNDA.n512 GNDA.n511 150
R1781 GNDA.n508 GNDA.n507 150
R1782 GNDA.n566 GNDA.n565 150
R1783 GNDA.n558 GNDA.n465 150
R1784 GNDA.n489 GNDA.n466 150
R1785 GNDA.n496 GNDA.n495 150
R1786 GNDA.n555 GNDA.n482 150
R1787 GNDA.n551 GNDA.n550 150
R1788 GNDA.n547 GNDA.n546 150
R1789 GNDA.n543 GNDA.n542 150
R1790 GNDA.n745 GNDA.n744 150
R1791 GNDA.n741 GNDA.n740 150
R1792 GNDA.n737 GNDA.n736 150
R1793 GNDA.n733 GNDA.n732 150
R1794 GNDA.n729 GNDA.n728 150
R1795 GNDA.n725 GNDA.n724 150
R1796 GNDA.n721 GNDA.n720 150
R1797 GNDA.n717 GNDA.n716 150
R1798 GNDA.n789 GNDA.n788 150
R1799 GNDA.n781 GNDA.n780 150
R1800 GNDA.n774 GNDA.n773 150
R1801 GNDA.n792 GNDA.n696 150
R1802 GNDA.n753 GNDA.n752 150
R1803 GNDA.n757 GNDA.n756 150
R1804 GNDA.n761 GNDA.n760 150
R1805 GNDA.n765 GNDA.n764 150
R1806 GNDA.n972 GNDA.n971 150
R1807 GNDA.n968 GNDA.n967 150
R1808 GNDA.n964 GNDA.n963 150
R1809 GNDA.n960 GNDA.n959 150
R1810 GNDA.n956 GNDA.n955 150
R1811 GNDA.n952 GNDA.n951 150
R1812 GNDA.n948 GNDA.n947 150
R1813 GNDA.n944 GNDA.n943 150
R1814 GNDA.n1022 GNDA.n941 150
R1815 GNDA.n1011 GNDA.n1010 150
R1816 GNDA.n1004 GNDA.n1003 150
R1817 GNDA.n1025 GNDA.n921 150
R1818 GNDA.n980 GNDA.n979 150
R1819 GNDA.n984 GNDA.n983 150
R1820 GNDA.n988 GNDA.n987 150
R1821 GNDA.n990 GNDA.n940 150
R1822 GNDA.n2180 GNDA.n2179 150
R1823 GNDA.n2176 GNDA.n2175 150
R1824 GNDA.n2172 GNDA.n2171 150
R1825 GNDA.n2168 GNDA.n2167 150
R1826 GNDA.n2164 GNDA.n2163 150
R1827 GNDA.n2160 GNDA.n2159 150
R1828 GNDA.n2156 GNDA.n2155 150
R1829 GNDA.n2152 GNDA.n2151 150
R1830 GNDA.n2205 GNDA.n662 150
R1831 GNDA.n2125 GNDA.n663 150
R1832 GNDA.n2133 GNDA.n2132 150
R1833 GNDA.n2140 GNDA.n2139 150
R1834 GNDA.n2188 GNDA.n2187 150
R1835 GNDA.n2192 GNDA.n2191 150
R1836 GNDA.n2196 GNDA.n2195 150
R1837 GNDA.n2202 GNDA.n680 150
R1838 GNDA.n2321 GNDA.n2320 150
R1839 GNDA.n2317 GNDA.n2316 150
R1840 GNDA.n2313 GNDA.n2312 150
R1841 GNDA.n2309 GNDA.n2308 150
R1842 GNDA.n2305 GNDA.n2304 150
R1843 GNDA.n2301 GNDA.n2300 150
R1844 GNDA.n2297 GNDA.n2296 150
R1845 GNDA.n2293 GNDA.n2292 150
R1846 GNDA.n2350 GNDA.n2349 150
R1847 GNDA.n2342 GNDA.n2248 150
R1848 GNDA.n2274 GNDA.n2249 150
R1849 GNDA.n2281 GNDA.n2280 150
R1850 GNDA.n2339 GNDA.n2265 150
R1851 GNDA.n2335 GNDA.n2334 150
R1852 GNDA.n2331 GNDA.n2330 150
R1853 GNDA.n2327 GNDA.n2326 150
R1854 GNDA.n1274 GNDA.n1272 150
R1855 GNDA.n1270 GNDA.n1238 150
R1856 GNDA.n1266 GNDA.n1264 150
R1857 GNDA.n1262 GNDA.n1240 150
R1858 GNDA.n1258 GNDA.n1256 150
R1859 GNDA.n1254 GNDA.n1242 150
R1860 GNDA.n1250 GNDA.n1249 150
R1861 GNDA.n1247 GNDA.n1245 150
R1862 GNDA.n1355 GNDA.n1353 150
R1863 GNDA.n1366 GNDA.n1225 150
R1864 GNDA.n1370 GNDA.n1368 150
R1865 GNDA.n1382 GNDA.n1219 150
R1866 GNDA.n1282 GNDA.n1280 150
R1867 GNDA.n1286 GNDA.n1234 150
R1868 GNDA.n1290 GNDA.n1288 150
R1869 GNDA.n1351 GNDA.n1232 150
R1870 GNDA.n2081 GNDA.n2080 150
R1871 GNDA.n2077 GNDA.n2076 150
R1872 GNDA.n2073 GNDA.n2072 150
R1873 GNDA.n2069 GNDA.n2068 150
R1874 GNDA.n2065 GNDA.n2064 150
R1875 GNDA.n2061 GNDA.n2060 150
R1876 GNDA.n2057 GNDA.n2056 150
R1877 GNDA.n2053 GNDA.n2052 150
R1878 GNDA.n2104 GNDA.n1037 150
R1879 GNDA.n2026 GNDA.n1038 150
R1880 GNDA.n2034 GNDA.n2033 150
R1881 GNDA.n2041 GNDA.n2040 150
R1882 GNDA.n2089 GNDA.n2088 150
R1883 GNDA.n2093 GNDA.n2092 150
R1884 GNDA.n2097 GNDA.n2096 150
R1885 GNDA.n2101 GNDA.n2100 150
R1886 GNDA.n2769 GNDA.t37 146.667
R1887 GNDA.t79 GNDA.n2768 146.667
R1888 GNDA.n2766 GNDA.t116 146.667
R1889 GNDA.n185 GNDA.t179 146.667
R1890 GNDA.n192 GNDA.t74 146.667
R1891 GNDA.n1671 GNDA.n1670 146.041
R1892 GNDA.t195 GNDA.t28 145.09
R1893 GNDA.n273 GNDA.t151 140.602
R1894 GNDA.n252 GNDA.t112 140.602
R1895 GNDA.n2490 GNDA.t169 140.602
R1896 GNDA.n1396 GNDA.n1112 138.81
R1897 GNDA.n1393 GNDA.t24 135.919
R1898 GNDA.n303 GNDA.t252 134.501
R1899 GNDA.n169 GNDA.t259 134.501
R1900 GNDA.t17 GNDA.n1556 134.474
R1901 GNDA.n1796 GNDA.n1795 134.268
R1902 GNDA.n1795 GNDA.n1793 134.268
R1903 GNDA.n1598 GNDA.n1597 132.721
R1904 GNDA.n803 GNDA.n802 132.721
R1905 GNDA.n2016 GNDA.n2015 132.721
R1906 GNDA.n7 GNDA.t270 130.713
R1907 GNDA.n1360 GNDA.n1359 130.136
R1908 GNDA.n1375 GNDA.n1374 130.136
R1909 GNDA.n1392 GNDA.n1391 130.136
R1910 GNDA.n1758 GNDA.n1113 130.136
R1911 GNDA.n1749 GNDA.n1113 130.136
R1912 GNDA.n1749 GNDA.n1748 130.136
R1913 GNDA.n1748 GNDA.n1747 130.136
R1914 GNDA.n1162 GNDA.n1161 130.136
R1915 GNDA.n1161 GNDA.n1150 130.136
R1916 GNDA.n1150 GNDA.n1146 130.136
R1917 GNDA.n1682 GNDA.n1146 130.136
R1918 GNDA.n1558 GNDA.n1557 130.136
R1919 GNDA.n1578 GNDA.n1561 130.136
R1920 GNDA.n1592 GNDA.n1591 130.136
R1921 GNDA.n2 GNDA.t23 130.001
R1922 GNDA.n13 GNDA.t302 130.001
R1923 GNDA.n16 GNDA.t288 130.001
R1924 GNDA.n19 GNDA.t306 130.001
R1925 GNDA.n2773 GNDA.t54 130.001
R1926 GNDA.n2407 GNDA.t109 130.001
R1927 GNDA.n347 GNDA.t280 130.001
R1928 GNDA.n344 GNDA.t52 130.001
R1929 GNDA.n2450 GNDA.t312 130.001
R1930 GNDA.n2453 GNDA.t41 130.001
R1931 GNDA.n8 GNDA.t133 130.001
R1932 GNDA.n352 GNDA.t194 130.001
R1933 GNDA.n353 GNDA.t2 130.001
R1934 GNDA.n2760 GNDA.t147 128.562
R1935 GNDA.n181 GNDA.t308 127.754
R1936 GNDA.n189 GNDA.t148 127.754
R1937 GNDA.n1396 GNDA.t221 125.797
R1938 GNDA.n1579 GNDA.t201 125.797
R1939 GNDA.n1467 GNDA.t89 125.797
R1940 GNDA.n1555 GNDA.n1554 124.832
R1941 GNDA.n1398 GNDA.n1397 124.832
R1942 GNDA.n1669 GNDA.n1668 124.832
R1943 GNDA.n2366 GNDA.n2365 124.832
R1944 GNDA.n2369 GNDA.n2368 124.832
R1945 GNDA.n441 GNDA.n436 124.832
R1946 GNDA.n2115 GNDA.n2114 124.832
R1947 GNDA.n1847 GNDA.n683 124.832
R1948 GNDA.n917 GNDA.n684 124.832
R1949 GNDA.n2117 GNDA.n682 124.832
R1950 GNDA.n435 GNDA.n431 124.832
R1951 GNDA.n1394 GNDA.n1211 124.832
R1952 GNDA.n1670 GNDA.t221 124.352
R1953 GNDA.t63 GNDA.t183 124.061
R1954 GNDA.t77 GNDA.t254 124.061
R1955 GNDA.t189 GNDA.t167 124.061
R1956 GNDA.t242 GNDA.t57 124.061
R1957 GNDA.n2524 GNDA.t50 122.501
R1958 GNDA.n101 GNDA.t48 122.501
R1959 GNDA.n2494 GNDA.t327 122.501
R1960 GNDA.n1092 GNDA.t61 122.501
R1961 GNDA.n1088 GNDA.t121 122.501
R1962 GNDA.n1090 GNDA.t135 122.501
R1963 GNDA.n1361 GNDA.t38 120.013
R1964 GNDA.n1377 GNDA.t32 120.013
R1965 GNDA.n1096 GNDA.t208 119.891
R1966 GNDA.t60 GNDA.t0 118.04
R1967 GNDA.t291 GNDA.t114 113.897
R1968 GNDA.t154 GNDA.t49 112.822
R1969 GNDA.t6 GNDA.t53 112.822
R1970 GNDA.n1815 GNDA.t292 111.049
R1971 GNDA.n1811 GNDA.t314 110.925
R1972 GNDA.n1812 GNDA.t102 110.659
R1973 GNDA.n1815 GNDA.t212 110.591
R1974 GNDA.n170 GNDA.t158 110.141
R1975 GNDA.n301 GNDA.t317 107.519
R1976 GNDA.t199 GNDA.n2403 101.853
R1977 GNDA.n1779 GNDA.n1778 101.718
R1978 GNDA.n1798 GNDA.n1797 101.718
R1979 GNDA.n1806 GNDA.n1805 101.718
R1980 GNDA.n1787 GNDA.n1786 101.718
R1981 GNDA.t97 GNDA.n2491 101.538
R1982 GNDA.t216 GNDA.n2769 101.538
R1983 GNDA.n2768 GNDA.t33 101.538
R1984 GNDA.t324 GNDA.n2766 101.538
R1985 GNDA.t221 GNDA.n376 47.6748
R1986 GNDA.t283 GNDA.t123 98.1749
R1987 GNDA.t319 GNDA.t283 98.1749
R1988 GNDA.n134 GNDA.n133 97.8707
R1989 GNDA.n138 GNDA.n137 97.8707
R1990 GNDA.n142 GNDA.n141 97.8707
R1991 GNDA.n144 GNDA.n143 97.8707
R1992 GNDA.n315 GNDA.n314 97.8707
R1993 GNDA.n1228 GNDA.t122 96.8786
R1994 GNDA.t127 GNDA.n130 95.7752
R1995 GNDA.n171 GNDA.t262 93.1969
R1996 GNDA.n179 GNDA.t236 92.9582
R1997 GNDA.n282 GNDA.n281 92.2612
R1998 GNDA.n290 GNDA.n289 92.2612
R1999 GNDA.n268 GNDA.n267 92.2612
R2000 GNDA.n261 GNDA.n218 92.2612
R2001 GNDA.n247 GNDA.n246 92.2612
R2002 GNDA.n240 GNDA.n239 92.2612
R2003 GNDA.n230 GNDA.n223 91.3721
R2004 GNDA.n249 GNDA.n248 91.3721
R2005 GNDA.n248 GNDA.n222 91.3721
R2006 GNDA.n211 GNDA.n206 91.3721
R2007 GNDA.n270 GNDA.n269 91.3721
R2008 GNDA.n269 GNDA.n205 91.3721
R2009 GNDA.n1593 GNDA.t138 91.0948
R2010 GNDA.n1784 GNDA.n1774 91.069
R2011 GNDA.n1777 GNDA.n1774 91.069
R2012 GNDA.n1781 GNDA.n1773 91.069
R2013 GNDA.n1782 GNDA.n1781 91.069
R2014 GNDA.n1800 GNDA.n1796 91.069
R2015 GNDA.n1802 GNDA.n1793 91.069
R2016 GNDA.n296 GNDA.n198 90.7567
R2017 GNDA.n2485 GNDA.n110 90.7567
R2018 GNDA.t301 GNDA.t141 90.2569
R2019 GNDA.t271 GNDA.t86 90.2569
R2020 GNDA.t322 GNDA.t281 90.2569
R2021 GNDA.t7 GNDA.t132 90.2569
R2022 GNDA.t215 GNDA.t127 87.3244
R2023 GNDA.t25 GNDA.t26 86.757
R2024 GNDA.t171 GNDA.t81 86.757
R2025 GNDA.n2745 GNDA.t332 86.0829
R2026 GNDA.n305 GNDA.t250 84.5075
R2027 GNDA.n1762 GNDA.n1111 84.306
R2028 GNDA.n1680 GNDA.n1673 84.306
R2029 GNDA.n299 GNDA.n197 84.306
R2030 GNDA.n294 GNDA.n195 84.306
R2031 GNDA.n272 GNDA.n208 84.306
R2032 GNDA.n274 GNDA.n207 84.306
R2033 GNDA.n251 GNDA.n227 84.306
R2034 GNDA.n253 GNDA.n224 84.306
R2035 GNDA.n109 GNDA.n107 84.306
R2036 GNDA.n2483 GNDA.n107 84.306
R2037 GNDA.n309 GNDA.n121 83.2005
R2038 GNDA.n309 GNDA.n308 83.2005
R2039 GNDA.n2745 GNDA.t330 82.8829
R2040 GNDA.n1761 GNDA.n1112 82.4192
R2041 GNDA.n1580 GNDA.t88 82.4192
R2042 GNDA.t192 GNDA.n377 82.4192
R2043 GNDA.n1593 GNDA.t191 82.4192
R2044 GNDA.n1933 GNDA.n1072 80.9821
R2045 GNDA.n1900 GNDA.n1824 80.9821
R2046 GNDA.n1228 GNDA.t172 76.6354
R2047 GNDA.t174 GNDA.n368 76.6354
R2048 GNDA.t9 GNDA.n1376 76.6354
R2049 GNDA.n1681 GNDA.n1671 76.6354
R2050 GNDA.t221 GNDA.n363 76.3879
R2051 GNDA.n1617 GNDA.n1616 76.3222
R2052 GNDA.n1612 GNDA.n1459 76.3222
R2053 GNDA.n1610 GNDA.n1609 76.3222
R2054 GNDA.n1605 GNDA.n1462 76.3222
R2055 GNDA.n1603 GNDA.n1602 76.3222
R2056 GNDA.n1638 GNDA.n1637 76.3222
R2057 GNDA.n1633 GNDA.n1450 76.3222
R2058 GNDA.n1631 GNDA.n1630 76.3222
R2059 GNDA.n1626 GNDA.n1453 76.3222
R2060 GNDA.n1624 GNDA.n1623 76.3222
R2061 GNDA.n1619 GNDA.n1456 76.3222
R2062 GNDA.n1641 GNDA.n1640 76.3222
R2063 GNDA.n1648 GNDA.n1647 76.3222
R2064 GNDA.n1651 GNDA.n1650 76.3222
R2065 GNDA.n1658 GNDA.n1657 76.3222
R2066 GNDA.n1661 GNDA.n1660 76.3222
R2067 GNDA.n1553 GNDA.n1170 76.3222
R2068 GNDA.n1417 GNDA.n1185 76.3222
R2069 GNDA.n1415 GNDA.n1191 76.3222
R2070 GNDA.n1196 GNDA.n1195 76.3222
R2071 GNDA.n1409 GNDA.n1194 76.3222
R2072 GNDA.n1405 GNDA.n1193 76.3222
R2073 GNDA.n1401 GNDA.n1192 76.3222
R2074 GNDA.n1425 GNDA.n1424 76.3222
R2075 GNDA.n1426 GNDA.n1183 76.3222
R2076 GNDA.n1433 GNDA.n1432 76.3222
R2077 GNDA.n1434 GNDA.n1181 76.3222
R2078 GNDA.n1441 GNDA.n1440 76.3222
R2079 GNDA.n1445 GNDA.n1179 76.3222
R2080 GNDA.n1446 GNDA.n1163 76.3222
R2081 GNDA.n1645 GNDA.n1164 76.3222
R2082 GNDA.n1176 GNDA.n1165 76.3222
R2083 GNDA.n1655 GNDA.n1166 76.3222
R2084 GNDA.n1665 GNDA.n1167 76.3222
R2085 GNDA.n1667 GNDA.n1149 76.3222
R2086 GNDA.n822 GNDA.n821 76.3222
R2087 GNDA.n817 GNDA.n688 76.3222
R2088 GNDA.n815 GNDA.n814 76.3222
R2089 GNDA.n810 GNDA.n691 76.3222
R2090 GNDA.n808 GNDA.n807 76.3222
R2091 GNDA.n844 GNDA.n384 76.3222
R2092 GNDA.n840 GNDA.n385 76.3222
R2093 GNDA.n836 GNDA.n386 76.3222
R2094 GNDA.n832 GNDA.n387 76.3222
R2095 GNDA.n828 GNDA.n388 76.3222
R2096 GNDA.n824 GNDA.n389 76.3222
R2097 GNDA.n2358 GNDA.n438 76.3222
R2098 GNDA.n450 GNDA.n445 76.3222
R2099 GNDA.n784 GNDA.n449 76.3222
R2100 GNDA.n777 GNDA.n448 76.3222
R2101 GNDA.n770 GNDA.n447 76.3222
R2102 GNDA.n796 GNDA.n446 76.3222
R2103 GNDA.n910 GNDA.n909 76.3222
R2104 GNDA.n902 GNDA.n872 76.3222
R2105 GNDA.n901 GNDA.n900 76.3222
R2106 GNDA.n894 GNDA.n880 76.3222
R2107 GNDA.n893 GNDA.n892 76.3222
R2108 GNDA.n2391 GNDA.n2390 76.3222
R2109 GNDA.n2388 GNDA.n2387 76.3222
R2110 GNDA.n2383 GNDA.n412 76.3222
R2111 GNDA.n2380 GNDA.n411 76.3222
R2112 GNDA.n2376 GNDA.n410 76.3222
R2113 GNDA.n2372 GNDA.n409 76.3222
R2114 GNDA.n848 GNDA.n390 76.3222
R2115 GNDA.n852 GNDA.n391 76.3222
R2116 GNDA.n856 GNDA.n392 76.3222
R2117 GNDA.n860 GNDA.n393 76.3222
R2118 GNDA.n864 GNDA.n394 76.3222
R2119 GNDA.n868 GNDA.n395 76.3222
R2120 GNDA.n570 GNDA.n433 76.3222
R2121 GNDA.n457 GNDA.n456 76.3222
R2122 GNDA.n561 GNDA.n455 76.3222
R2123 GNDA.n487 GNDA.n454 76.3222
R2124 GNDA.n491 GNDA.n453 76.3222
R2125 GNDA.n500 GNDA.n452 76.3222
R2126 GNDA.n873 GNDA.n869 76.3222
R2127 GNDA.n876 GNDA.n875 76.3222
R2128 GNDA.n881 GNDA.n878 76.3222
R2129 GNDA.n884 GNDA.n883 76.3222
R2130 GNDA.n889 GNDA.n886 76.3222
R2131 GNDA.n888 GNDA.n887 76.3222
R2132 GNDA.n1993 GNDA.n1060 76.3222
R2133 GNDA.n2000 GNDA.n1999 76.3222
R2134 GNDA.n2001 GNDA.n1058 76.3222
R2135 GNDA.n2008 GNDA.n2007 76.3222
R2136 GNDA.n2009 GNDA.n1056 76.3222
R2137 GNDA.n914 GNDA.n648 76.3222
R2138 GNDA.n2107 GNDA.n647 76.3222
R2139 GNDA.n2024 GNDA.n646 76.3222
R2140 GNDA.n2030 GNDA.n645 76.3222
R2141 GNDA.n2036 GNDA.n644 76.3222
R2142 GNDA.n2045 GNDA.n643 76.3222
R2143 GNDA.n993 GNDA.n654 76.3222
R2144 GNDA.n1019 GNDA.n653 76.3222
R2145 GNDA.n1014 GNDA.n652 76.3222
R2146 GNDA.n1007 GNDA.n651 76.3222
R2147 GNDA.n1000 GNDA.n650 76.3222
R2148 GNDA.n1029 GNDA.n649 76.3222
R2149 GNDA.n2212 GNDA.n2211 76.3222
R2150 GNDA.n2209 GNDA.n2208 76.3222
R2151 GNDA.n2123 GNDA.n658 76.3222
R2152 GNDA.n2129 GNDA.n657 76.3222
R2153 GNDA.n2135 GNDA.n656 76.3222
R2154 GNDA.n2144 GNDA.n655 76.3222
R2155 GNDA.n2236 GNDA.n2235 76.3222
R2156 GNDA.n2230 GNDA.n580 76.3222
R2157 GNDA.n2227 GNDA.n581 76.3222
R2158 GNDA.n2223 GNDA.n582 76.3222
R2159 GNDA.n2219 GNDA.n583 76.3222
R2160 GNDA.n424 GNDA.n402 76.3222
R2161 GNDA.n425 GNDA.n414 76.3222
R2162 GNDA.n426 GNDA.n416 76.3222
R2163 GNDA.n427 GNDA.n418 76.3222
R2164 GNDA.n428 GNDA.n420 76.3222
R2165 GNDA.n430 GNDA.n422 76.3222
R2166 GNDA.n607 GNDA.n396 76.3222
R2167 GNDA.n603 GNDA.n397 76.3222
R2168 GNDA.n599 GNDA.n398 76.3222
R2169 GNDA.n595 GNDA.n399 76.3222
R2170 GNDA.n591 GNDA.n400 76.3222
R2171 GNDA.n2396 GNDA.n2395 76.3222
R2172 GNDA.n2356 GNDA.n2355 76.3222
R2173 GNDA.n2242 GNDA.n575 76.3222
R2174 GNDA.n2345 GNDA.n574 76.3222
R2175 GNDA.n2272 GNDA.n573 76.3222
R2176 GNDA.n2276 GNDA.n572 76.3222
R2177 GNDA.n2285 GNDA.n571 76.3222
R2178 GNDA.n611 GNDA.n585 76.3222
R2179 GNDA.n615 GNDA.n586 76.3222
R2180 GNDA.n619 GNDA.n587 76.3222
R2181 GNDA.n623 GNDA.n588 76.3222
R2182 GNDA.n629 GNDA.n628 76.3222
R2183 GNDA.n1188 GNDA.n1187 76.3222
R2184 GNDA.n1198 GNDA.n1197 76.3222
R2185 GNDA.n1201 GNDA.n1200 76.3222
R2186 GNDA.n1204 GNDA.n1203 76.3222
R2187 GNDA.n1207 GNDA.n1206 76.3222
R2188 GNDA.n1210 GNDA.n1209 76.3222
R2189 GNDA.n1320 GNDA.n1319 76.3222
R2190 GNDA.n1315 GNDA.n1296 76.3222
R2191 GNDA.n1313 GNDA.n1312 76.3222
R2192 GNDA.n1308 GNDA.n1299 76.3222
R2193 GNDA.n1306 GNDA.n1305 76.3222
R2194 GNDA.n1301 GNDA.n1300 76.3222
R2195 GNDA.n1322 GNDA.n636 76.3222
R2196 GNDA.n1326 GNDA.n635 76.3222
R2197 GNDA.n1330 GNDA.n634 76.3222
R2198 GNDA.n1334 GNDA.n633 76.3222
R2199 GNDA.n1338 GNDA.n632 76.3222
R2200 GNDA.n1325 GNDA.n636 76.3222
R2201 GNDA.n1329 GNDA.n635 76.3222
R2202 GNDA.n1333 GNDA.n634 76.3222
R2203 GNDA.n1337 GNDA.n633 76.3222
R2204 GNDA.n1340 GNDA.n632 76.3222
R2205 GNDA.n614 GNDA.n585 76.3222
R2206 GNDA.n618 GNDA.n586 76.3222
R2207 GNDA.n622 GNDA.n587 76.3222
R2208 GNDA.n590 GNDA.n588 76.3222
R2209 GNDA.n629 GNDA.n589 76.3222
R2210 GNDA.n2236 GNDA.n638 76.3222
R2211 GNDA.n2228 GNDA.n580 76.3222
R2212 GNDA.n2224 GNDA.n581 76.3222
R2213 GNDA.n2220 GNDA.n582 76.3222
R2214 GNDA.n2216 GNDA.n583 76.3222
R2215 GNDA.n887 GNDA.n441 76.3222
R2216 GNDA.n890 GNDA.n889 76.3222
R2217 GNDA.n885 GNDA.n884 76.3222
R2218 GNDA.n882 GNDA.n881 76.3222
R2219 GNDA.n877 GNDA.n876 76.3222
R2220 GNDA.n874 GNDA.n873 76.3222
R2221 GNDA.n909 GNDA.n908 76.3222
R2222 GNDA.n903 GNDA.n902 76.3222
R2223 GNDA.n900 GNDA.n899 76.3222
R2224 GNDA.n895 GNDA.n894 76.3222
R2225 GNDA.n892 GNDA.n439 76.3222
R2226 GNDA.n1668 GNDA.n1667 76.3222
R2227 GNDA.n1665 GNDA.n1664 76.3222
R2228 GNDA.n1171 GNDA.n1166 76.3222
R2229 GNDA.n1654 GNDA.n1165 76.3222
R2230 GNDA.n1175 GNDA.n1164 76.3222
R2231 GNDA.n1644 GNDA.n1163 76.3222
R2232 GNDA.n1640 GNDA.n1177 76.3222
R2233 GNDA.n1649 GNDA.n1648 76.3222
R2234 GNDA.n1650 GNDA.n1173 76.3222
R2235 GNDA.n1659 GNDA.n1658 76.3222
R2236 GNDA.n1662 GNDA.n1661 76.3222
R2237 GNDA.n1554 GNDA.n1553 76.3222
R2238 GNDA.n1211 GNDA.n1210 76.3222
R2239 GNDA.n1208 GNDA.n1207 76.3222
R2240 GNDA.n1205 GNDA.n1204 76.3222
R2241 GNDA.n1202 GNDA.n1201 76.3222
R2242 GNDA.n1199 GNDA.n1198 76.3222
R2243 GNDA.n1189 GNDA.n1188 76.3222
R2244 GNDA.n1418 GNDA.n1417 76.3222
R2245 GNDA.n1415 GNDA.n1414 76.3222
R2246 GNDA.n1410 GNDA.n1195 76.3222
R2247 GNDA.n1406 GNDA.n1194 76.3222
R2248 GNDA.n1402 GNDA.n1193 76.3222
R2249 GNDA.n1398 GNDA.n1192 76.3222
R2250 GNDA.n431 GNDA.n430 76.3222
R2251 GNDA.n428 GNDA.n421 76.3222
R2252 GNDA.n427 GNDA.n419 76.3222
R2253 GNDA.n426 GNDA.n417 76.3222
R2254 GNDA.n425 GNDA.n415 76.3222
R2255 GNDA.n424 GNDA.n423 76.3222
R2256 GNDA.n2390 GNDA.n408 76.3222
R2257 GNDA.n2388 GNDA.n413 76.3222
R2258 GNDA.n2381 GNDA.n412 76.3222
R2259 GNDA.n2377 GNDA.n411 76.3222
R2260 GNDA.n2373 GNDA.n410 76.3222
R2261 GNDA.n2369 GNDA.n409 76.3222
R2262 GNDA.n2396 GNDA.n401 76.3222
R2263 GNDA.n594 GNDA.n400 76.3222
R2264 GNDA.n598 GNDA.n399 76.3222
R2265 GNDA.n602 GNDA.n398 76.3222
R2266 GNDA.n606 GNDA.n397 76.3222
R2267 GNDA.n610 GNDA.n396 76.3222
R2268 GNDA.n865 GNDA.n395 76.3222
R2269 GNDA.n861 GNDA.n394 76.3222
R2270 GNDA.n857 GNDA.n393 76.3222
R2271 GNDA.n853 GNDA.n392 76.3222
R2272 GNDA.n849 GNDA.n391 76.3222
R2273 GNDA.n407 GNDA.n390 76.3222
R2274 GNDA.n827 GNDA.n389 76.3222
R2275 GNDA.n831 GNDA.n388 76.3222
R2276 GNDA.n835 GNDA.n387 76.3222
R2277 GNDA.n839 GNDA.n386 76.3222
R2278 GNDA.n843 GNDA.n385 76.3222
R2279 GNDA.n871 GNDA.n384 76.3222
R2280 GNDA.n2211 GNDA.n642 76.3222
R2281 GNDA.n2209 GNDA.n659 76.3222
R2282 GNDA.n2128 GNDA.n658 76.3222
R2283 GNDA.n2136 GNDA.n657 76.3222
R2284 GNDA.n2143 GNDA.n656 76.3222
R2285 GNDA.n2118 GNDA.n655 76.3222
R2286 GNDA.n1018 GNDA.n654 76.3222
R2287 GNDA.n1015 GNDA.n653 76.3222
R2288 GNDA.n1008 GNDA.n652 76.3222
R2289 GNDA.n1001 GNDA.n651 76.3222
R2290 GNDA.n1028 GNDA.n650 76.3222
R2291 GNDA.n1032 GNDA.n649 76.3222
R2292 GNDA.n2108 GNDA.n648 76.3222
R2293 GNDA.n2023 GNDA.n647 76.3222
R2294 GNDA.n2029 GNDA.n646 76.3222
R2295 GNDA.n2037 GNDA.n645 76.3222
R2296 GNDA.n2044 GNDA.n644 76.3222
R2297 GNDA.n2018 GNDA.n643 76.3222
R2298 GNDA.n1302 GNDA.n1301 76.3222
R2299 GNDA.n1307 GNDA.n1306 76.3222
R2300 GNDA.n1299 GNDA.n1297 76.3222
R2301 GNDA.n1314 GNDA.n1313 76.3222
R2302 GNDA.n1296 GNDA.n1294 76.3222
R2303 GNDA.n1321 GNDA.n1320 76.3222
R2304 GNDA.n1442 GNDA.n1179 76.3222
R2305 GNDA.n1440 GNDA.n1439 76.3222
R2306 GNDA.n1435 GNDA.n1434 76.3222
R2307 GNDA.n1432 GNDA.n1431 76.3222
R2308 GNDA.n1427 GNDA.n1426 76.3222
R2309 GNDA.n1424 GNDA.n1423 76.3222
R2310 GNDA.n1456 GNDA.n1454 76.3222
R2311 GNDA.n1625 GNDA.n1624 76.3222
R2312 GNDA.n1453 GNDA.n1451 76.3222
R2313 GNDA.n1632 GNDA.n1631 76.3222
R2314 GNDA.n1450 GNDA.n1448 76.3222
R2315 GNDA.n1639 GNDA.n1638 76.3222
R2316 GNDA.n2356 GNDA.n576 76.3222
R2317 GNDA.n2346 GNDA.n575 76.3222
R2318 GNDA.n2271 GNDA.n574 76.3222
R2319 GNDA.n2277 GNDA.n573 76.3222
R2320 GNDA.n2284 GNDA.n572 76.3222
R2321 GNDA.n2266 GNDA.n571 76.3222
R2322 GNDA.n570 GNDA.n569 76.3222
R2323 GNDA.n562 GNDA.n456 76.3222
R2324 GNDA.n486 GNDA.n455 76.3222
R2325 GNDA.n492 GNDA.n454 76.3222
R2326 GNDA.n499 GNDA.n453 76.3222
R2327 GNDA.n452 GNDA.n451 76.3222
R2328 GNDA.n2359 GNDA.n2358 76.3222
R2329 GNDA.n785 GNDA.n450 76.3222
R2330 GNDA.n778 GNDA.n449 76.3222
R2331 GNDA.n771 GNDA.n448 76.3222
R2332 GNDA.n795 GNDA.n447 76.3222
R2333 GNDA.n800 GNDA.n446 76.3222
R2334 GNDA.n1597 GNDA.n1463 76.3222
R2335 GNDA.n1604 GNDA.n1603 76.3222
R2336 GNDA.n1462 GNDA.n1460 76.3222
R2337 GNDA.n1611 GNDA.n1610 76.3222
R2338 GNDA.n1459 GNDA.n1457 76.3222
R2339 GNDA.n1618 GNDA.n1617 76.3222
R2340 GNDA.n802 GNDA.n692 76.3222
R2341 GNDA.n809 GNDA.n808 76.3222
R2342 GNDA.n691 GNDA.n689 76.3222
R2343 GNDA.n816 GNDA.n815 76.3222
R2344 GNDA.n688 GNDA.n686 76.3222
R2345 GNDA.n823 GNDA.n822 76.3222
R2346 GNDA.n2015 GNDA.n2014 76.3222
R2347 GNDA.n2010 GNDA.n2009 76.3222
R2348 GNDA.n2007 GNDA.n2006 76.3222
R2349 GNDA.n2002 GNDA.n2001 76.3222
R2350 GNDA.n1999 GNDA.n1998 76.3222
R2351 GNDA.n1994 GNDA.n1993 76.3222
R2352 GNDA.t163 GNDA.t239 76.0568
R2353 GNDA.n1706 GNDA.n1130 74.5978
R2354 GNDA.n1703 GNDA.n1130 74.5978
R2355 GNDA.n1516 GNDA.n1479 74.5978
R2356 GNDA.n1513 GNDA.n1479 74.5978
R2357 GNDA.n523 GNDA.n471 74.5978
R2358 GNDA.n520 GNDA.n471 74.5978
R2359 GNDA.n732 GNDA.n703 74.5978
R2360 GNDA.n729 GNDA.n703 74.5978
R2361 GNDA.n959 GNDA.n928 74.5978
R2362 GNDA.n956 GNDA.n928 74.5978
R2363 GNDA.n2167 GNDA.n669 74.5978
R2364 GNDA.n2164 GNDA.n669 74.5978
R2365 GNDA.n2308 GNDA.n2254 74.5978
R2366 GNDA.n2305 GNDA.n2254 74.5978
R2367 GNDA.n1257 GNDA.n1240 74.5978
R2368 GNDA.n1258 GNDA.n1257 74.5978
R2369 GNDA.n2068 GNDA.n1044 74.5978
R2370 GNDA.n2065 GNDA.n1044 74.5978
R2371 GNDA.n171 GNDA.n170 73.428
R2372 GNDA.t262 GNDA.t315 73.334
R2373 GNDA.t65 GNDA.t236 73.2399
R2374 GNDA.t103 GNDA.t65 73.2399
R2375 GNDA.t125 GNDA.t103 73.2399
R2376 GNDA.t315 GNDA.t125 73.2399
R2377 GNDA.t188 GNDA.t296 73.2399
R2378 GNDA.t273 GNDA.t213 73.2399
R2379 GNDA.t12 GNDA.t232 73.2399
R2380 GNDA.t187 GNDA.t313 71.9351
R2381 GNDA.t59 GNDA.t187 71.9351
R2382 GNDA.t101 GNDA.t59 71.9351
R2383 GNDA.t162 GNDA.t211 71.9351
R2384 GNDA.t114 GNDA.t162 71.9351
R2385 GNDA.t210 GNDA.t291 71.9351
R2386 GNDA.t90 GNDA.t210 71.9351
R2387 GNDA.t258 GNDA.t293 70.6038
R2388 GNDA.t84 GNDA.t91 70.423
R2389 GNDA.n1089 GNDA.n1087 70.2133
R2390 GNDA.n1082 GNDA.n1081 69.4466
R2391 GNDA.n1754 GNDA.n1118 69.3109
R2392 GNDA.n1725 GNDA.n1118 69.3109
R2393 GNDA.n1585 GNDA.n1584 69.3109
R2394 GNDA.n1585 GNDA.n1490 69.3109
R2395 GNDA.n566 GNDA.n461 69.3109
R2396 GNDA.n542 GNDA.n461 69.3109
R2397 GNDA.n790 GNDA.n789 69.3109
R2398 GNDA.n790 GNDA.n765 69.3109
R2399 GNDA.n1023 GNDA.n1022 69.3109
R2400 GNDA.n1023 GNDA.n940 69.3109
R2401 GNDA.n2203 GNDA.n662 69.3109
R2402 GNDA.n2203 GNDA.n2202 69.3109
R2403 GNDA.n2350 GNDA.n2244 69.3109
R2404 GNDA.n2326 GNDA.n2244 69.3109
R2405 GNDA.n1353 GNDA.n1352 69.3109
R2406 GNDA.n1352 GNDA.n1351 69.3109
R2407 GNDA.n2102 GNDA.n1037 69.3109
R2408 GNDA.n2102 GNDA.n2101 69.3109
R2409 GNDA.t221 GNDA.n368 67.9598
R2410 GNDA.t309 GNDA.t326 67.6928
R2411 GNDA.n176 GNDA.n175 66.5605
R2412 GNDA.n175 GNDA.n174 66.5605
R2413 GNDA.t225 GNDA.n196 66.1659
R2414 GNDA.t165 GNDA.n225 66.1659
R2415 GNDA.n226 GNDA.t156 66.1659
R2416 GNDA.n175 GNDA.n124 65.9634
R2417 GNDA.t223 GNDA.n1739 65.8183
R2418 GNDA.t223 GNDA.n1139 65.8183
R2419 GNDA.t223 GNDA.n1138 65.8183
R2420 GNDA.t223 GNDA.n1137 65.8183
R2421 GNDA.t223 GNDA.n1128 65.8183
R2422 GNDA.t223 GNDA.n1135 65.8183
R2423 GNDA.t223 GNDA.n1126 65.8183
R2424 GNDA.t223 GNDA.n1136 65.8183
R2425 GNDA.t223 GNDA.n1134 65.8183
R2426 GNDA.t223 GNDA.n1133 65.8183
R2427 GNDA.t223 GNDA.n1132 65.8183
R2428 GNDA.t223 GNDA.n1131 65.8183
R2429 GNDA.t222 GNDA.n1489 65.8183
R2430 GNDA.t222 GNDA.n1488 65.8183
R2431 GNDA.t222 GNDA.n1487 65.8183
R2432 GNDA.t222 GNDA.n1486 65.8183
R2433 GNDA.t222 GNDA.n1478 65.8183
R2434 GNDA.t222 GNDA.n1484 65.8183
R2435 GNDA.t222 GNDA.n1475 65.8183
R2436 GNDA.t222 GNDA.n1485 65.8183
R2437 GNDA.t222 GNDA.n1483 65.8183
R2438 GNDA.t222 GNDA.n1482 65.8183
R2439 GNDA.t222 GNDA.n1481 65.8183
R2440 GNDA.t222 GNDA.n1480 65.8183
R2441 GNDA.n1586 GNDA.t222 65.8183
R2442 GNDA.t222 GNDA.n1477 65.8183
R2443 GNDA.t222 GNDA.n1476 65.8183
R2444 GNDA.t222 GNDA.n1474 65.8183
R2445 GNDA.t223 GNDA.n1129 65.8183
R2446 GNDA.t223 GNDA.n1127 65.8183
R2447 GNDA.n1742 GNDA.t223 65.8183
R2448 GNDA.t223 GNDA.n1119 65.8183
R2449 GNDA.t220 GNDA.n556 65.8183
R2450 GNDA.t220 GNDA.n480 65.8183
R2451 GNDA.t220 GNDA.n479 65.8183
R2452 GNDA.t220 GNDA.n478 65.8183
R2453 GNDA.t220 GNDA.n469 65.8183
R2454 GNDA.t220 GNDA.n476 65.8183
R2455 GNDA.t220 GNDA.n467 65.8183
R2456 GNDA.t220 GNDA.n477 65.8183
R2457 GNDA.t220 GNDA.n475 65.8183
R2458 GNDA.t220 GNDA.n474 65.8183
R2459 GNDA.t220 GNDA.n473 65.8183
R2460 GNDA.t220 GNDA.n472 65.8183
R2461 GNDA.t220 GNDA.n470 65.8183
R2462 GNDA.t220 GNDA.n468 65.8183
R2463 GNDA.n557 GNDA.t220 65.8183
R2464 GNDA.t220 GNDA.n462 65.8183
R2465 GNDA.t227 GNDA.n714 65.8183
R2466 GNDA.t227 GNDA.n713 65.8183
R2467 GNDA.t227 GNDA.n712 65.8183
R2468 GNDA.t227 GNDA.n711 65.8183
R2469 GNDA.t227 GNDA.n702 65.8183
R2470 GNDA.t227 GNDA.n709 65.8183
R2471 GNDA.t227 GNDA.n699 65.8183
R2472 GNDA.t227 GNDA.n710 65.8183
R2473 GNDA.t227 GNDA.n708 65.8183
R2474 GNDA.t227 GNDA.n706 65.8183
R2475 GNDA.t227 GNDA.n705 65.8183
R2476 GNDA.t227 GNDA.n704 65.8183
R2477 GNDA.n791 GNDA.t227 65.8183
R2478 GNDA.t227 GNDA.n701 65.8183
R2479 GNDA.t227 GNDA.n700 65.8183
R2480 GNDA.t227 GNDA.n698 65.8183
R2481 GNDA.t229 GNDA.n939 65.8183
R2482 GNDA.t229 GNDA.n938 65.8183
R2483 GNDA.t229 GNDA.n937 65.8183
R2484 GNDA.t229 GNDA.n936 65.8183
R2485 GNDA.t229 GNDA.n927 65.8183
R2486 GNDA.t229 GNDA.n934 65.8183
R2487 GNDA.t229 GNDA.n924 65.8183
R2488 GNDA.t229 GNDA.n935 65.8183
R2489 GNDA.t229 GNDA.n933 65.8183
R2490 GNDA.t229 GNDA.n931 65.8183
R2491 GNDA.t229 GNDA.n930 65.8183
R2492 GNDA.t229 GNDA.n929 65.8183
R2493 GNDA.n1024 GNDA.t229 65.8183
R2494 GNDA.t229 GNDA.n926 65.8183
R2495 GNDA.t229 GNDA.n925 65.8183
R2496 GNDA.t229 GNDA.n923 65.8183
R2497 GNDA.t265 GNDA.n679 65.8183
R2498 GNDA.t265 GNDA.n678 65.8183
R2499 GNDA.t265 GNDA.n677 65.8183
R2500 GNDA.t265 GNDA.n676 65.8183
R2501 GNDA.t265 GNDA.n667 65.8183
R2502 GNDA.t265 GNDA.n674 65.8183
R2503 GNDA.t265 GNDA.n664 65.8183
R2504 GNDA.t265 GNDA.n675 65.8183
R2505 GNDA.t265 GNDA.n673 65.8183
R2506 GNDA.t265 GNDA.n672 65.8183
R2507 GNDA.t265 GNDA.n671 65.8183
R2508 GNDA.t265 GNDA.n670 65.8183
R2509 GNDA.t265 GNDA.n668 65.8183
R2510 GNDA.t265 GNDA.n666 65.8183
R2511 GNDA.t265 GNDA.n665 65.8183
R2512 GNDA.n2204 GNDA.t265 65.8183
R2513 GNDA.t230 GNDA.n2340 65.8183
R2514 GNDA.t230 GNDA.n2263 65.8183
R2515 GNDA.t230 GNDA.n2262 65.8183
R2516 GNDA.t230 GNDA.n2261 65.8183
R2517 GNDA.t230 GNDA.n2252 65.8183
R2518 GNDA.t230 GNDA.n2259 65.8183
R2519 GNDA.t230 GNDA.n2250 65.8183
R2520 GNDA.t230 GNDA.n2260 65.8183
R2521 GNDA.t230 GNDA.n2258 65.8183
R2522 GNDA.t230 GNDA.n2257 65.8183
R2523 GNDA.t230 GNDA.n2256 65.8183
R2524 GNDA.t230 GNDA.n2255 65.8183
R2525 GNDA.t230 GNDA.n2253 65.8183
R2526 GNDA.t230 GNDA.n2251 65.8183
R2527 GNDA.n2341 GNDA.t230 65.8183
R2528 GNDA.t230 GNDA.n2245 65.8183
R2529 GNDA.n1279 GNDA.t228 65.8183
R2530 GNDA.n1281 GNDA.t228 65.8183
R2531 GNDA.n1287 GNDA.t228 65.8183
R2532 GNDA.n1289 GNDA.t228 65.8183
R2533 GNDA.n1263 GNDA.t228 65.8183
R2534 GNDA.n1265 GNDA.t228 65.8183
R2535 GNDA.n1271 GNDA.t228 65.8183
R2536 GNDA.n1273 GNDA.t228 65.8183
R2537 GNDA.t228 GNDA.n1218 65.8183
R2538 GNDA.n1248 GNDA.t228 65.8183
R2539 GNDA.n1244 GNDA.t228 65.8183
R2540 GNDA.n1255 GNDA.t228 65.8183
R2541 GNDA.n1383 GNDA.t228 65.8183
R2542 GNDA.n1369 GNDA.t228 65.8183
R2543 GNDA.n1367 GNDA.t228 65.8183
R2544 GNDA.n1354 GNDA.t228 65.8183
R2545 GNDA.t260 GNDA.n1054 65.8183
R2546 GNDA.t260 GNDA.n1053 65.8183
R2547 GNDA.t260 GNDA.n1052 65.8183
R2548 GNDA.t260 GNDA.n1051 65.8183
R2549 GNDA.t260 GNDA.n1042 65.8183
R2550 GNDA.t260 GNDA.n1049 65.8183
R2551 GNDA.t260 GNDA.n1039 65.8183
R2552 GNDA.t260 GNDA.n1050 65.8183
R2553 GNDA.t260 GNDA.n1048 65.8183
R2554 GNDA.t260 GNDA.n1047 65.8183
R2555 GNDA.t260 GNDA.n1046 65.8183
R2556 GNDA.t260 GNDA.n1045 65.8183
R2557 GNDA.t260 GNDA.n1043 65.8183
R2558 GNDA.t260 GNDA.n1041 65.8183
R2559 GNDA.t260 GNDA.n1040 65.8183
R2560 GNDA.n2103 GNDA.t260 65.8183
R2561 GNDA.t129 GNDA.t297 64.7892
R2562 GNDA.t221 GNDA.n1162 62.176
R2563 GNDA.t221 GNDA.n377 62.176
R2564 GNDA.n2774 GNDA.n2773 60.29
R2565 GNDA.n2781 GNDA.n19 60.29
R2566 GNDA.n2787 GNDA.n16 60.29
R2567 GNDA.n2794 GNDA.n13 60.29
R2568 GNDA.n2822 GNDA.n2 60.29
R2569 GNDA.n2408 GNDA.n2407 60.29
R2570 GNDA.n2436 GNDA.n347 60.29
R2571 GNDA.n2442 GNDA.n344 60.29
R2572 GNDA.n2450 GNDA.n2449 60.29
R2573 GNDA.n2454 GNDA.n2453 60.29
R2574 GNDA.n125 GNDA.t104 60.0005
R2575 GNDA.n125 GNDA.t126 60.0005
R2576 GNDA.n120 GNDA.t214 60.0005
R2577 GNDA.n120 GNDA.t92 60.0005
R2578 GNDA.n122 GNDA.t13 60.0005
R2579 GNDA.n122 GNDA.t233 60.0005
R2580 GNDA.t240 GNDA.n127 60.0005
R2581 GNDA.n127 GNDA.t274 60.0005
R2582 GNDA.n126 GNDA.t316 60.0005
R2583 GNDA.n126 GNDA.t263 60.0005
R2584 GNDA.t237 GNDA.n177 60.0005
R2585 GNDA.n177 GNDA.t66 60.0005
R2586 GNDA.n1092 GNDA.n328 59.5478
R2587 GNDA.n1088 GNDA.n334 59.5478
R2588 GNDA.n1090 GNDA.n330 59.5478
R2589 GNDA.n1747 GNDA.t161 59.2841
R2590 GNDA.n2506 GNDA.n101 58.9809
R2591 GNDA.n2524 GNDA.n2523 58.9809
R2592 GNDA.n2495 GNDA.n2494 58.9809
R2593 GNDA.t123 GNDA.n194 58.0127
R2594 GNDA.t183 GNDA.t277 57.8952
R2595 GNDA.t30 GNDA.t44 57.8952
R2596 GNDA.t167 GNDA.t15 57.8952
R2597 GNDA.t246 GNDA.t131 57.8952
R2598 GNDA.t105 GNDA.t242 57.8952
R2599 GNDA.t222 GNDA.n1585 57.8461
R2600 GNDA.t223 GNDA.n1118 57.8461
R2601 GNDA.t220 GNDA.n461 57.8461
R2602 GNDA.t227 GNDA.n790 57.8461
R2603 GNDA.t229 GNDA.n1023 57.8461
R2604 GNDA.t265 GNDA.n2203 57.8461
R2605 GNDA.t230 GNDA.n2244 57.8461
R2606 GNDA.n1352 GNDA.t228 57.8461
R2607 GNDA.t260 GNDA.n2102 57.8461
R2608 GNDA.t206 GNDA.t221 57.8382
R2609 GNDA.t177 GNDA.t221 57.8382
R2610 GNDA.n2493 GNDA.t10 56.4108
R2611 GNDA.n2772 GNDA.t289 56.4108
R2612 GNDA.n2215 GNDA.n584 56.3995
R2613 GNDA.n2239 GNDA.n2238 56.3995
R2614 GNDA.n1343 GNDA.n630 56.3995
R2615 GNDA.n1345 GNDA.n630 56.3995
R2616 GNDA.n2238 GNDA.n577 56.3995
R2617 GNDA.n2213 GNDA.n584 56.3995
R2618 GNDA.n1598 GNDA.n1596 56.3995
R2619 GNDA.n803 GNDA.n801 56.3995
R2620 GNDA.n2017 GNDA.n2016 56.3995
R2621 GNDA.t223 GNDA.n1130 55.2026
R2622 GNDA.t222 GNDA.n1479 55.2026
R2623 GNDA.t220 GNDA.n471 55.2026
R2624 GNDA.t227 GNDA.n703 55.2026
R2625 GNDA.t229 GNDA.n928 55.2026
R2626 GNDA.t265 GNDA.n669 55.2026
R2627 GNDA.t230 GNDA.n2254 55.2026
R2628 GNDA.n1257 GNDA.t228 55.2026
R2629 GNDA.t260 GNDA.n1044 55.2026
R2630 GNDA.n2807 GNDA.n8 54.4005
R2631 GNDA.n2809 GNDA.n7 54.4005
R2632 GNDA.n2598 GNDA.n2527 54.4005
R2633 GNDA.n2421 GNDA.n353 54.4005
R2634 GNDA.n2423 GNDA.n352 54.4005
R2635 GNDA.n2625 GNDA.n83 54.4005
R2636 GNDA.t172 GNDA.n369 53.5003
R2637 GNDA.n1361 GNDA.t174 53.5003
R2638 GNDA.n1377 GNDA.t9 53.5003
R2639 GNDA.n1682 GNDA.n1681 53.5003
R2640 GNDA.n1721 GNDA.n1136 53.3664
R2641 GNDA.n1718 GNDA.n1126 53.3664
R2642 GNDA.n1714 GNDA.n1135 53.3664
R2643 GNDA.n1710 GNDA.n1128 53.3664
R2644 GNDA.n1699 GNDA.n1131 53.3664
R2645 GNDA.n1695 GNDA.n1132 53.3664
R2646 GNDA.n1691 GNDA.n1133 53.3664
R2647 GNDA.n1687 GNDA.n1134 53.3664
R2648 GNDA.n1753 GNDA.n1119 53.3664
R2649 GNDA.n1742 GNDA.n1741 53.3664
R2650 GNDA.n1127 GNDA.n1125 53.3664
R2651 GNDA.n1156 GNDA.n1129 53.3664
R2652 GNDA.n1739 GNDA.n1738 53.3664
R2653 GNDA.n1141 GNDA.n1139 53.3664
R2654 GNDA.n1733 GNDA.n1138 53.3664
R2655 GNDA.n1729 GNDA.n1137 53.3664
R2656 GNDA.n1739 GNDA.n1140 53.3664
R2657 GNDA.n1734 GNDA.n1139 53.3664
R2658 GNDA.n1730 GNDA.n1138 53.3664
R2659 GNDA.n1726 GNDA.n1137 53.3664
R2660 GNDA.n1707 GNDA.n1128 53.3664
R2661 GNDA.n1711 GNDA.n1135 53.3664
R2662 GNDA.n1715 GNDA.n1126 53.3664
R2663 GNDA.n1719 GNDA.n1136 53.3664
R2664 GNDA.n1690 GNDA.n1134 53.3664
R2665 GNDA.n1694 GNDA.n1133 53.3664
R2666 GNDA.n1698 GNDA.n1132 53.3664
R2667 GNDA.n1702 GNDA.n1131 53.3664
R2668 GNDA.n1532 GNDA.n1485 53.3664
R2669 GNDA.n1528 GNDA.n1475 53.3664
R2670 GNDA.n1524 GNDA.n1484 53.3664
R2671 GNDA.n1520 GNDA.n1478 53.3664
R2672 GNDA.n1509 GNDA.n1480 53.3664
R2673 GNDA.n1505 GNDA.n1481 53.3664
R2674 GNDA.n1501 GNDA.n1482 53.3664
R2675 GNDA.n1497 GNDA.n1483 53.3664
R2676 GNDA.n1491 GNDA.n1474 53.3664
R2677 GNDA.n1574 GNDA.n1476 53.3664
R2678 GNDA.n1569 GNDA.n1477 53.3664
R2679 GNDA.n1587 GNDA.n1586 53.3664
R2680 GNDA.n1536 GNDA.n1489 53.3664
R2681 GNDA.n1537 GNDA.n1488 53.3664
R2682 GNDA.n1541 GNDA.n1487 53.3664
R2683 GNDA.n1545 GNDA.n1486 53.3664
R2684 GNDA.n1533 GNDA.n1489 53.3664
R2685 GNDA.n1540 GNDA.n1488 53.3664
R2686 GNDA.n1544 GNDA.n1487 53.3664
R2687 GNDA.n1547 GNDA.n1486 53.3664
R2688 GNDA.n1517 GNDA.n1478 53.3664
R2689 GNDA.n1521 GNDA.n1484 53.3664
R2690 GNDA.n1525 GNDA.n1475 53.3664
R2691 GNDA.n1529 GNDA.n1485 53.3664
R2692 GNDA.n1500 GNDA.n1483 53.3664
R2693 GNDA.n1504 GNDA.n1482 53.3664
R2694 GNDA.n1508 GNDA.n1481 53.3664
R2695 GNDA.n1512 GNDA.n1480 53.3664
R2696 GNDA.n1586 GNDA.n1473 53.3664
R2697 GNDA.n1477 GNDA.n1471 53.3664
R2698 GNDA.n1570 GNDA.n1476 53.3664
R2699 GNDA.n1573 GNDA.n1474 53.3664
R2700 GNDA.n1686 GNDA.n1129 53.3664
R2701 GNDA.n1157 GNDA.n1127 53.3664
R2702 GNDA.n1743 GNDA.n1742 53.3664
R2703 GNDA.n1740 GNDA.n1119 53.3664
R2704 GNDA.n538 GNDA.n477 53.3664
R2705 GNDA.n535 GNDA.n467 53.3664
R2706 GNDA.n531 GNDA.n476 53.3664
R2707 GNDA.n527 GNDA.n469 53.3664
R2708 GNDA.n516 GNDA.n472 53.3664
R2709 GNDA.n512 GNDA.n473 53.3664
R2710 GNDA.n508 GNDA.n474 53.3664
R2711 GNDA.n504 GNDA.n475 53.3664
R2712 GNDA.n565 GNDA.n462 53.3664
R2713 GNDA.n558 GNDA.n557 53.3664
R2714 GNDA.n489 GNDA.n468 53.3664
R2715 GNDA.n496 GNDA.n470 53.3664
R2716 GNDA.n556 GNDA.n555 53.3664
R2717 GNDA.n482 GNDA.n480 53.3664
R2718 GNDA.n550 GNDA.n479 53.3664
R2719 GNDA.n546 GNDA.n478 53.3664
R2720 GNDA.n556 GNDA.n481 53.3664
R2721 GNDA.n551 GNDA.n480 53.3664
R2722 GNDA.n547 GNDA.n479 53.3664
R2723 GNDA.n543 GNDA.n478 53.3664
R2724 GNDA.n524 GNDA.n469 53.3664
R2725 GNDA.n528 GNDA.n476 53.3664
R2726 GNDA.n532 GNDA.n467 53.3664
R2727 GNDA.n536 GNDA.n477 53.3664
R2728 GNDA.n507 GNDA.n475 53.3664
R2729 GNDA.n511 GNDA.n474 53.3664
R2730 GNDA.n515 GNDA.n473 53.3664
R2731 GNDA.n519 GNDA.n472 53.3664
R2732 GNDA.n503 GNDA.n470 53.3664
R2733 GNDA.n495 GNDA.n468 53.3664
R2734 GNDA.n557 GNDA.n466 53.3664
R2735 GNDA.n465 GNDA.n462 53.3664
R2736 GNDA.n748 GNDA.n710 53.3664
R2737 GNDA.n744 GNDA.n699 53.3664
R2738 GNDA.n740 GNDA.n709 53.3664
R2739 GNDA.n736 GNDA.n702 53.3664
R2740 GNDA.n725 GNDA.n704 53.3664
R2741 GNDA.n721 GNDA.n705 53.3664
R2742 GNDA.n717 GNDA.n706 53.3664
R2743 GNDA.n708 GNDA.n707 53.3664
R2744 GNDA.n788 GNDA.n698 53.3664
R2745 GNDA.n781 GNDA.n700 53.3664
R2746 GNDA.n774 GNDA.n701 53.3664
R2747 GNDA.n792 GNDA.n791 53.3664
R2748 GNDA.n752 GNDA.n714 53.3664
R2749 GNDA.n753 GNDA.n713 53.3664
R2750 GNDA.n757 GNDA.n712 53.3664
R2751 GNDA.n761 GNDA.n711 53.3664
R2752 GNDA.n749 GNDA.n714 53.3664
R2753 GNDA.n756 GNDA.n713 53.3664
R2754 GNDA.n760 GNDA.n712 53.3664
R2755 GNDA.n764 GNDA.n711 53.3664
R2756 GNDA.n733 GNDA.n702 53.3664
R2757 GNDA.n737 GNDA.n709 53.3664
R2758 GNDA.n741 GNDA.n699 53.3664
R2759 GNDA.n745 GNDA.n710 53.3664
R2760 GNDA.n716 GNDA.n708 53.3664
R2761 GNDA.n720 GNDA.n706 53.3664
R2762 GNDA.n724 GNDA.n705 53.3664
R2763 GNDA.n728 GNDA.n704 53.3664
R2764 GNDA.n791 GNDA.n697 53.3664
R2765 GNDA.n701 GNDA.n696 53.3664
R2766 GNDA.n773 GNDA.n700 53.3664
R2767 GNDA.n780 GNDA.n698 53.3664
R2768 GNDA.n975 GNDA.n935 53.3664
R2769 GNDA.n971 GNDA.n924 53.3664
R2770 GNDA.n967 GNDA.n934 53.3664
R2771 GNDA.n963 GNDA.n927 53.3664
R2772 GNDA.n952 GNDA.n929 53.3664
R2773 GNDA.n948 GNDA.n930 53.3664
R2774 GNDA.n944 GNDA.n931 53.3664
R2775 GNDA.n933 GNDA.n932 53.3664
R2776 GNDA.n941 GNDA.n923 53.3664
R2777 GNDA.n1011 GNDA.n925 53.3664
R2778 GNDA.n1004 GNDA.n926 53.3664
R2779 GNDA.n1025 GNDA.n1024 53.3664
R2780 GNDA.n979 GNDA.n939 53.3664
R2781 GNDA.n980 GNDA.n938 53.3664
R2782 GNDA.n984 GNDA.n937 53.3664
R2783 GNDA.n988 GNDA.n936 53.3664
R2784 GNDA.n976 GNDA.n939 53.3664
R2785 GNDA.n983 GNDA.n938 53.3664
R2786 GNDA.n987 GNDA.n937 53.3664
R2787 GNDA.n990 GNDA.n936 53.3664
R2788 GNDA.n960 GNDA.n927 53.3664
R2789 GNDA.n964 GNDA.n934 53.3664
R2790 GNDA.n968 GNDA.n924 53.3664
R2791 GNDA.n972 GNDA.n935 53.3664
R2792 GNDA.n943 GNDA.n933 53.3664
R2793 GNDA.n947 GNDA.n931 53.3664
R2794 GNDA.n951 GNDA.n930 53.3664
R2795 GNDA.n955 GNDA.n929 53.3664
R2796 GNDA.n1024 GNDA.n922 53.3664
R2797 GNDA.n926 GNDA.n921 53.3664
R2798 GNDA.n1003 GNDA.n925 53.3664
R2799 GNDA.n1010 GNDA.n923 53.3664
R2800 GNDA.n2183 GNDA.n675 53.3664
R2801 GNDA.n2179 GNDA.n664 53.3664
R2802 GNDA.n2175 GNDA.n674 53.3664
R2803 GNDA.n2171 GNDA.n667 53.3664
R2804 GNDA.n2160 GNDA.n670 53.3664
R2805 GNDA.n2156 GNDA.n671 53.3664
R2806 GNDA.n2152 GNDA.n672 53.3664
R2807 GNDA.n2148 GNDA.n673 53.3664
R2808 GNDA.n2205 GNDA.n2204 53.3664
R2809 GNDA.n2125 GNDA.n665 53.3664
R2810 GNDA.n2133 GNDA.n666 53.3664
R2811 GNDA.n2140 GNDA.n668 53.3664
R2812 GNDA.n2187 GNDA.n679 53.3664
R2813 GNDA.n2188 GNDA.n678 53.3664
R2814 GNDA.n2192 GNDA.n677 53.3664
R2815 GNDA.n2196 GNDA.n676 53.3664
R2816 GNDA.n2184 GNDA.n679 53.3664
R2817 GNDA.n2191 GNDA.n678 53.3664
R2818 GNDA.n2195 GNDA.n677 53.3664
R2819 GNDA.n680 GNDA.n676 53.3664
R2820 GNDA.n2168 GNDA.n667 53.3664
R2821 GNDA.n2172 GNDA.n674 53.3664
R2822 GNDA.n2176 GNDA.n664 53.3664
R2823 GNDA.n2180 GNDA.n675 53.3664
R2824 GNDA.n2151 GNDA.n673 53.3664
R2825 GNDA.n2155 GNDA.n672 53.3664
R2826 GNDA.n2159 GNDA.n671 53.3664
R2827 GNDA.n2163 GNDA.n670 53.3664
R2828 GNDA.n2147 GNDA.n668 53.3664
R2829 GNDA.n2139 GNDA.n666 53.3664
R2830 GNDA.n2132 GNDA.n665 53.3664
R2831 GNDA.n2204 GNDA.n663 53.3664
R2832 GNDA.n2323 GNDA.n2260 53.3664
R2833 GNDA.n2320 GNDA.n2250 53.3664
R2834 GNDA.n2316 GNDA.n2259 53.3664
R2835 GNDA.n2312 GNDA.n2252 53.3664
R2836 GNDA.n2301 GNDA.n2255 53.3664
R2837 GNDA.n2297 GNDA.n2256 53.3664
R2838 GNDA.n2293 GNDA.n2257 53.3664
R2839 GNDA.n2289 GNDA.n2258 53.3664
R2840 GNDA.n2349 GNDA.n2245 53.3664
R2841 GNDA.n2342 GNDA.n2341 53.3664
R2842 GNDA.n2274 GNDA.n2251 53.3664
R2843 GNDA.n2281 GNDA.n2253 53.3664
R2844 GNDA.n2340 GNDA.n2339 53.3664
R2845 GNDA.n2265 GNDA.n2263 53.3664
R2846 GNDA.n2334 GNDA.n2262 53.3664
R2847 GNDA.n2330 GNDA.n2261 53.3664
R2848 GNDA.n2340 GNDA.n2264 53.3664
R2849 GNDA.n2335 GNDA.n2263 53.3664
R2850 GNDA.n2331 GNDA.n2262 53.3664
R2851 GNDA.n2327 GNDA.n2261 53.3664
R2852 GNDA.n2309 GNDA.n2252 53.3664
R2853 GNDA.n2313 GNDA.n2259 53.3664
R2854 GNDA.n2317 GNDA.n2250 53.3664
R2855 GNDA.n2321 GNDA.n2260 53.3664
R2856 GNDA.n2292 GNDA.n2258 53.3664
R2857 GNDA.n2296 GNDA.n2257 53.3664
R2858 GNDA.n2300 GNDA.n2256 53.3664
R2859 GNDA.n2304 GNDA.n2255 53.3664
R2860 GNDA.n2288 GNDA.n2253 53.3664
R2861 GNDA.n2280 GNDA.n2251 53.3664
R2862 GNDA.n2341 GNDA.n2249 53.3664
R2863 GNDA.n2248 GNDA.n2245 53.3664
R2864 GNDA.n1273 GNDA.n1236 53.3664
R2865 GNDA.n1272 GNDA.n1271 53.3664
R2866 GNDA.n1265 GNDA.n1238 53.3664
R2867 GNDA.n1264 GNDA.n1263 53.3664
R2868 GNDA.n1255 GNDA.n1254 53.3664
R2869 GNDA.n1250 GNDA.n1244 53.3664
R2870 GNDA.n1248 GNDA.n1247 53.3664
R2871 GNDA.n1385 GNDA.n1218 53.3664
R2872 GNDA.n1355 GNDA.n1354 53.3664
R2873 GNDA.n1367 GNDA.n1366 53.3664
R2874 GNDA.n1370 GNDA.n1369 53.3664
R2875 GNDA.n1383 GNDA.n1382 53.3664
R2876 GNDA.n1280 GNDA.n1279 53.3664
R2877 GNDA.n1282 GNDA.n1281 53.3664
R2878 GNDA.n1287 GNDA.n1286 53.3664
R2879 GNDA.n1290 GNDA.n1289 53.3664
R2880 GNDA.n1279 GNDA.n1278 53.3664
R2881 GNDA.n1281 GNDA.n1234 53.3664
R2882 GNDA.n1288 GNDA.n1287 53.3664
R2883 GNDA.n1289 GNDA.n1232 53.3664
R2884 GNDA.n1263 GNDA.n1262 53.3664
R2885 GNDA.n1266 GNDA.n1265 53.3664
R2886 GNDA.n1271 GNDA.n1270 53.3664
R2887 GNDA.n1274 GNDA.n1273 53.3664
R2888 GNDA.n1245 GNDA.n1218 53.3664
R2889 GNDA.n1249 GNDA.n1248 53.3664
R2890 GNDA.n1244 GNDA.n1242 53.3664
R2891 GNDA.n1256 GNDA.n1255 53.3664
R2892 GNDA.n1384 GNDA.n1383 53.3664
R2893 GNDA.n1369 GNDA.n1219 53.3664
R2894 GNDA.n1368 GNDA.n1367 53.3664
R2895 GNDA.n1354 GNDA.n1225 53.3664
R2896 GNDA.n2084 GNDA.n1050 53.3664
R2897 GNDA.n2080 GNDA.n1039 53.3664
R2898 GNDA.n2076 GNDA.n1049 53.3664
R2899 GNDA.n2072 GNDA.n1042 53.3664
R2900 GNDA.n2061 GNDA.n1045 53.3664
R2901 GNDA.n2057 GNDA.n1046 53.3664
R2902 GNDA.n2053 GNDA.n1047 53.3664
R2903 GNDA.n2049 GNDA.n1048 53.3664
R2904 GNDA.n2104 GNDA.n2103 53.3664
R2905 GNDA.n2026 GNDA.n1040 53.3664
R2906 GNDA.n2034 GNDA.n1041 53.3664
R2907 GNDA.n2041 GNDA.n1043 53.3664
R2908 GNDA.n2088 GNDA.n1054 53.3664
R2909 GNDA.n2089 GNDA.n1053 53.3664
R2910 GNDA.n2093 GNDA.n1052 53.3664
R2911 GNDA.n2097 GNDA.n1051 53.3664
R2912 GNDA.n2085 GNDA.n1054 53.3664
R2913 GNDA.n2092 GNDA.n1053 53.3664
R2914 GNDA.n2096 GNDA.n1052 53.3664
R2915 GNDA.n2100 GNDA.n1051 53.3664
R2916 GNDA.n2069 GNDA.n1042 53.3664
R2917 GNDA.n2073 GNDA.n1049 53.3664
R2918 GNDA.n2077 GNDA.n1039 53.3664
R2919 GNDA.n2081 GNDA.n1050 53.3664
R2920 GNDA.n2052 GNDA.n1048 53.3664
R2921 GNDA.n2056 GNDA.n1047 53.3664
R2922 GNDA.n2060 GNDA.n1046 53.3664
R2923 GNDA.n2064 GNDA.n1045 53.3664
R2924 GNDA.n2048 GNDA.n1043 53.3664
R2925 GNDA.n2040 GNDA.n1041 53.3664
R2926 GNDA.n2033 GNDA.n1040 53.3664
R2927 GNDA.n2103 GNDA.n1038 53.3664
R2928 GNDA.n194 GNDA.n179 50.7047
R2929 GNDA.n2550 GNDA.t117 48.0005
R2930 GNDA.n2550 GNDA.t150 48.0005
R2931 GNDA.n2549 GNDA.t36 48.0005
R2932 GNDA.n2549 GNDA.t325 48.0005
R2933 GNDA.n2544 GNDA.t80 48.0005
R2934 GNDA.n2544 GNDA.t34 48.0005
R2935 GNDA.n2542 GNDA.t323 48.0005
R2936 GNDA.n2542 GNDA.t8 48.0005
R2937 GNDA.n2537 GNDA.t142 48.0005
R2938 GNDA.n2537 GNDA.t87 48.0005
R2939 GNDA.n2533 GNDA.t4 48.0005
R2940 GNDA.n2533 GNDA.t72 48.0005
R2941 GNDA.n2530 GNDA.t203 48.0005
R2942 GNDA.n2530 GNDA.t46 48.0005
R2943 GNDA.n88 GNDA.t295 48.0005
R2944 GNDA.n88 GNDA.t98 48.0005
R2945 GNDA.n86 GNDA.t186 48.0005
R2946 GNDA.n86 GNDA.t56 48.0005
R2947 GNDA.n78 GNDA.t198 48.0005
R2948 GNDA.n78 GNDA.t160 48.0005
R2949 GNDA.n76 GNDA.t170 48.0005
R2950 GNDA.n76 GNDA.t96 48.0005
R2951 GNDA.n71 GNDA.t106 48.0005
R2952 GNDA.n71 GNDA.t58 48.0005
R2953 GNDA.n66 GNDA.t286 48.0005
R2954 GNDA.n66 GNDA.t176 48.0005
R2955 GNDA.n65 GNDA.t113 48.0005
R2956 GNDA.n65 GNDA.t140 48.0005
R2957 GNDA.n60 GNDA.t16 48.0005
R2958 GNDA.n60 GNDA.t190 48.0005
R2959 GNDA.n55 GNDA.t152 48.0005
R2960 GNDA.n55 GNDA.t43 48.0005
R2961 GNDA.n54 GNDA.t78 48.0005
R2962 GNDA.n54 GNDA.t205 48.0005
R2963 GNDA.n49 GNDA.t278 48.0005
R2964 GNDA.n49 GNDA.t64 48.0005
R2965 GNDA.n44 GNDA.t320 48.0005
R2966 GNDA.n44 GNDA.t318 48.0005
R2967 GNDA.n43 GNDA.t124 48.0005
R2968 GNDA.n43 GNDA.t284 48.0005
R2969 GNDA.n38 GNDA.t196 48.0005
R2970 GNDA.n38 GNDA.t119 48.0005
R2971 GNDA.n2399 GNDA.t90 47.9569
R2972 GNDA.t297 GNDA.t93 47.8878
R2973 GNDA.n1761 GNDA.n1758 47.7166
R2974 GNDA.t88 GNDA.n1579 47.7166
R2975 GNDA.n1467 GNDA.t192 47.7166
R2976 GNDA.t191 GNDA.n378 47.7166
R2977 GNDA.t221 GNDA.n2397 47.6748
R2978 GNDA.t299 GNDA.t73 45.1287
R2979 GNDA.t45 GNDA.t305 45.1287
R2980 GNDA.t35 GNDA.t22 45.1287
R2981 GNDA.t14 GNDA.t153 44.1582
R2982 GNDA.t146 GNDA.n2763 42.5811
R2983 GNDA.n2763 GNDA.t179 42.5811
R2984 GNDA.t74 GNDA.n185 42.5811
R2985 GNDA.t28 GNDA.n192 42.5811
R2986 GNDA.t91 GNDA.t303 42.254
R2987 GNDA.n310 GNDA.n309 41.6005
R2988 GNDA.t317 GNDA.n300 41.3539
R2989 GNDA.n273 GNDA.t204 41.3539
R2990 GNDA.n2489 GNDA.t110 41.3539
R2991 GNDA.t95 GNDA.n2490 41.3539
R2992 GNDA.n2479 GNDA.n2477 41.3005
R2993 GNDA.n301 GNDA.t319 40.1628
R2994 GNDA.t293 GNDA.t20 39.5347
R2995 GNDA.n2747 GNDA.n2746 39.4989
R2996 GNDA.n165 GNDA.n124 39.4985
R2997 GNDA.n194 GNDA.t153 39.427
R2998 GNDA.n1556 GNDA.t5 39.0409
R2999 GNDA.n1558 GNDA.t171 39.0409
R3000 GNDA.n1561 GNDA.t107 39.0409
R3001 GNDA.t138 GNDA.n1592 39.0409
R3002 GNDA.n1393 GNDA.t39 37.595
R3003 GNDA.t239 GNDA.t82 36.6202
R3004 GNDA.t82 GNDA.t273 36.6202
R3005 GNDA.n183 GNDA.n182 35.6576
R3006 GNDA.n2730 GNDA.n32 35.6576
R3007 GNDA.n188 GNDA.n187 35.6576
R3008 GNDA.n190 GNDA.n35 35.6576
R3009 GNDA.t221 GNDA.n378 34.7031
R3010 GNDA.t118 GNDA.t14 34.6958
R3011 GNDA.n27 GNDA.n26 34.3278
R3012 GNDA.n2761 GNDA.n2759 34.3278
R3013 GNDA.t116 GNDA.n2765 33.8467
R3014 GNDA.n1359 GNDA.t122 33.2572
R3015 GNDA.n1374 GNDA.t173 33.2572
R3016 GNDA.n1391 GNDA.t25 33.2572
R3017 GNDA.n2823 GNDA.n2822 33.0991
R3018 GNDA.n2408 GNDA.n0 33.0991
R3019 GNDA.n1789 GNDA.n1788 33.0531
R3020 GNDA.t221 GNDA.n374 32.9056
R3021 GNDA.t221 GNDA.n375 32.9056
R3022 GNDA.n2398 GNDA.t221 32.6313
R3023 GNDA.n1808 GNDA.n1807 32.3969
R3024 GNDA.t221 GNDA.n379 32.2075
R3025 GNDA.n282 GNDA.n280 32.0005
R3026 GNDA.n280 GNDA.n202 32.0005
R3027 GNDA.n288 GNDA.n287 32.0005
R3028 GNDA.n287 GNDA.n200 32.0005
R3029 GNDA.n283 GNDA.n200 32.0005
R3030 GNDA.n213 GNDA.n204 32.0005
R3031 GNDA.n266 GNDA.n216 32.0005
R3032 GNDA.n262 GNDA.n216 32.0005
R3033 GNDA.n262 GNDA.n261 32.0005
R3034 GNDA.n260 GNDA.n219 32.0005
R3035 GNDA.n256 GNDA.n219 32.0005
R3036 GNDA.n255 GNDA.n221 32.0005
R3037 GNDA.n232 GNDA.n221 32.0005
R3038 GNDA.n245 GNDA.n236 32.0005
R3039 GNDA.n241 GNDA.n236 32.0005
R3040 GNDA.n2480 GNDA.n111 32.0005
R3041 GNDA.n165 GNDA.n164 32.0005
R3042 GNDA.n164 GNDA.n163 32.0005
R3043 GNDA.n163 GNDA.n132 32.0005
R3044 GNDA.n159 GNDA.n132 32.0005
R3045 GNDA.n159 GNDA.n158 32.0005
R3046 GNDA.n158 GNDA.n157 32.0005
R3047 GNDA.n157 GNDA.n136 32.0005
R3048 GNDA.n153 GNDA.n136 32.0005
R3049 GNDA.n153 GNDA.n152 32.0005
R3050 GNDA.n152 GNDA.n151 32.0005
R3051 GNDA.n151 GNDA.n140 32.0005
R3052 GNDA.n147 GNDA.n140 32.0005
R3053 GNDA.n147 GNDA.n146 32.0005
R3054 GNDA.n146 GNDA.n119 32.0005
R3055 GNDA.n311 GNDA.n119 32.0005
R3056 GNDA.n317 GNDA.n117 32.0005
R3057 GNDA.n318 GNDA.n317 32.0005
R3058 GNDA.n319 GNDA.n318 32.0005
R3059 GNDA.n319 GNDA.n114 32.0005
R3060 GNDA.n324 GNDA.n114 32.0005
R3061 GNDA.n325 GNDA.n324 32.0005
R3062 GNDA.n2496 GNDA.n104 32.0005
R3063 GNDA.n2500 GNDA.n104 32.0005
R3064 GNDA.n2501 GNDA.n2500 32.0005
R3065 GNDA.n2502 GNDA.n2501 32.0005
R3066 GNDA.n2502 GNDA.n102 32.0005
R3067 GNDA.n2506 GNDA.n102 32.0005
R3068 GNDA.n2507 GNDA.n2506 32.0005
R3069 GNDA.n2508 GNDA.n2507 32.0005
R3070 GNDA.n2508 GNDA.n99 32.0005
R3071 GNDA.n2513 GNDA.n99 32.0005
R3072 GNDA.n2514 GNDA.n2513 32.0005
R3073 GNDA.n2515 GNDA.n2514 32.0005
R3074 GNDA.n2515 GNDA.n96 32.0005
R3075 GNDA.n2522 GNDA.n97 32.0005
R3076 GNDA.n2518 GNDA.n97 32.0005
R3077 GNDA.n2518 GNDA.n22 32.0005
R3078 GNDA.n2775 GNDA.n22 32.0005
R3079 GNDA.n2779 GNDA.n20 32.0005
R3080 GNDA.n2780 GNDA.n2779 32.0005
R3081 GNDA.n2782 GNDA.n17 32.0005
R3082 GNDA.n2786 GNDA.n17 32.0005
R3083 GNDA.n2789 GNDA.n2788 32.0005
R3084 GNDA.n2789 GNDA.n14 32.0005
R3085 GNDA.n2793 GNDA.n14 32.0005
R3086 GNDA.n2796 GNDA.n2795 32.0005
R3087 GNDA.n2796 GNDA.n11 32.0005
R3088 GNDA.n2800 GNDA.n11 32.0005
R3089 GNDA.n2801 GNDA.n2800 32.0005
R3090 GNDA.n2802 GNDA.n2801 32.0005
R3091 GNDA.n2802 GNDA.n9 32.0005
R3092 GNDA.n2806 GNDA.n9 32.0005
R3093 GNDA.n2810 GNDA.n5 32.0005
R3094 GNDA.n2814 GNDA.n5 32.0005
R3095 GNDA.n2815 GNDA.n2814 32.0005
R3096 GNDA.n2816 GNDA.n2815 32.0005
R3097 GNDA.n2816 GNDA.n3 32.0005
R3098 GNDA.n2820 GNDA.n3 32.0005
R3099 GNDA.n2821 GNDA.n2820 32.0005
R3100 GNDA.n2472 GNDA.n328 32.0005
R3101 GNDA.n2472 GNDA.n2471 32.0005
R3102 GNDA.n2471 GNDA.n2470 32.0005
R3103 GNDA.n2467 GNDA.n2466 32.0005
R3104 GNDA.n2466 GNDA.n2465 32.0005
R3105 GNDA.n2465 GNDA.n332 32.0005
R3106 GNDA.n2461 GNDA.n2460 32.0005
R3107 GNDA.n2460 GNDA.n2459 32.0005
R3108 GNDA.n2459 GNDA.n335 32.0005
R3109 GNDA.n2455 GNDA.n335 32.0005
R3110 GNDA.n340 GNDA.n337 32.0005
R3111 GNDA.n340 GNDA.n338 32.0005
R3112 GNDA.n2448 GNDA.n339 32.0005
R3113 GNDA.n2444 GNDA.n339 32.0005
R3114 GNDA.n2444 GNDA.n2443 32.0005
R3115 GNDA.n2441 GNDA.n345 32.0005
R3116 GNDA.n2437 GNDA.n345 32.0005
R3117 GNDA.n2435 GNDA.n2434 32.0005
R3118 GNDA.n2434 GNDA.n348 32.0005
R3119 GNDA.n2430 GNDA.n348 32.0005
R3120 GNDA.n2430 GNDA.n2429 32.0005
R3121 GNDA.n2429 GNDA.n2428 32.0005
R3122 GNDA.n2428 GNDA.n350 32.0005
R3123 GNDA.n2424 GNDA.n350 32.0005
R3124 GNDA.n2420 GNDA.n354 32.0005
R3125 GNDA.n2416 GNDA.n354 32.0005
R3126 GNDA.n2416 GNDA.n2415 32.0005
R3127 GNDA.n2415 GNDA.n2414 32.0005
R3128 GNDA.n2414 GNDA.n356 32.0005
R3129 GNDA.n2410 GNDA.n356 32.0005
R3130 GNDA.n2410 GNDA.n2409 32.0005
R3131 GNDA.n2713 GNDA.n2712 32.0005
R3132 GNDA.n2712 GNDA.n2711 32.0005
R3133 GNDA.n2711 GNDA.n41 32.0005
R3134 GNDA.n2707 GNDA.n41 32.0005
R3135 GNDA.n2705 GNDA.n2704 32.0005
R3136 GNDA.n2701 GNDA.n2700 32.0005
R3137 GNDA.n2700 GNDA.n2699 32.0005
R3138 GNDA.n2696 GNDA.n2695 32.0005
R3139 GNDA.n2695 GNDA.n2694 32.0005
R3140 GNDA.n2691 GNDA.n2690 32.0005
R3141 GNDA.n2690 GNDA.n2689 32.0005
R3142 GNDA.n2689 GNDA.n52 32.0005
R3143 GNDA.n2685 GNDA.n52 32.0005
R3144 GNDA.n2683 GNDA.n2682 32.0005
R3145 GNDA.n2679 GNDA.n2678 32.0005
R3146 GNDA.n2678 GNDA.n2677 32.0005
R3147 GNDA.n2674 GNDA.n2673 32.0005
R3148 GNDA.n2673 GNDA.n2672 32.0005
R3149 GNDA.n2669 GNDA.n2668 32.0005
R3150 GNDA.n2668 GNDA.n2667 32.0005
R3151 GNDA.n2667 GNDA.n63 32.0005
R3152 GNDA.n2663 GNDA.n63 32.0005
R3153 GNDA.n2661 GNDA.n2660 32.0005
R3154 GNDA.n2657 GNDA.n2656 32.0005
R3155 GNDA.n2656 GNDA.n2655 32.0005
R3156 GNDA.n2652 GNDA.n2651 32.0005
R3157 GNDA.n2649 GNDA.n72 32.0005
R3158 GNDA.n2645 GNDA.n72 32.0005
R3159 GNDA.n2645 GNDA.n2644 32.0005
R3160 GNDA.n2644 GNDA.n2643 32.0005
R3161 GNDA.n2643 GNDA.n74 32.0005
R3162 GNDA.n2639 GNDA.n2638 32.0005
R3163 GNDA.n2636 GNDA.n79 32.0005
R3164 GNDA.n2632 GNDA.n79 32.0005
R3165 GNDA.n2632 GNDA.n2631 32.0005
R3166 GNDA.n2631 GNDA.n2630 32.0005
R3167 GNDA.n2630 GNDA.n81 32.0005
R3168 GNDA.n2626 GNDA.n81 32.0005
R3169 GNDA.n2624 GNDA.n2623 32.0005
R3170 GNDA.n2623 GNDA.n84 32.0005
R3171 GNDA.n2619 GNDA.n2618 32.0005
R3172 GNDA.n2616 GNDA.n89 32.0005
R3173 GNDA.n2612 GNDA.n89 32.0005
R3174 GNDA.n2610 GNDA.n2609 32.0005
R3175 GNDA.n2609 GNDA.n91 32.0005
R3176 GNDA.n2605 GNDA.n2604 32.0005
R3177 GNDA.n2604 GNDA.n2603 32.0005
R3178 GNDA.n2603 GNDA.n94 32.0005
R3179 GNDA.n2599 GNDA.n94 32.0005
R3180 GNDA.n2597 GNDA.n2596 32.0005
R3181 GNDA.n2596 GNDA.n2528 32.0005
R3182 GNDA.n2592 GNDA.n2528 32.0005
R3183 GNDA.n2592 GNDA.n2591 32.0005
R3184 GNDA.n2589 GNDA.n2531 32.0005
R3185 GNDA.n2585 GNDA.n2584 32.0005
R3186 GNDA.n2584 GNDA.n2583 32.0005
R3187 GNDA.n2583 GNDA.n2535 32.0005
R3188 GNDA.n2579 GNDA.n2535 32.0005
R3189 GNDA.n2579 GNDA.n2578 32.0005
R3190 GNDA.n2578 GNDA.n2577 32.0005
R3191 GNDA.n2574 GNDA.n2573 32.0005
R3192 GNDA.n2573 GNDA.n2572 32.0005
R3193 GNDA.n2572 GNDA.n2540 32.0005
R3194 GNDA.n2568 GNDA.n2567 32.0005
R3195 GNDA.n2565 GNDA.n2545 32.0005
R3196 GNDA.n2561 GNDA.n2545 32.0005
R3197 GNDA.n2561 GNDA.n2560 32.0005
R3198 GNDA.n2558 GNDA.n2547 32.0005
R3199 GNDA.n2554 GNDA.n2547 32.0005
R3200 GNDA.n2554 GNDA.n2553 32.0005
R3201 GNDA.n2737 GNDA.n28 32.0005
R3202 GNDA.n2737 GNDA.n2736 32.0005
R3203 GNDA.n2736 GNDA.n2735 32.0005
R3204 GNDA.n2735 GNDA.n30 32.0005
R3205 GNDA.n2731 GNDA.n30 32.0005
R3206 GNDA.n2730 GNDA.n2729 32.0005
R3207 GNDA.n2729 GNDA.n33 32.0005
R3208 GNDA.n2725 GNDA.n33 32.0005
R3209 GNDA.n2725 GNDA.n2724 32.0005
R3210 GNDA.n2724 GNDA.n2723 32.0005
R3211 GNDA.n2719 GNDA.n35 32.0005
R3212 GNDA.n2719 GNDA.n2718 32.0005
R3213 GNDA.n2748 GNDA.n2747 32.0005
R3214 GNDA.n2748 GNDA.n2743 32.0005
R3215 GNDA.n2752 GNDA.n2743 32.0005
R3216 GNDA.n2753 GNDA.n2752 32.0005
R3217 GNDA.n2754 GNDA.n2753 32.0005
R3218 GNDA.n2754 GNDA.n2741 32.0005
R3219 GNDA.n2758 GNDA.n2741 32.0005
R3220 GNDA.t20 GNDA.t188 30.9864
R3221 GNDA.n2718 GNDA.n2717 29.4625
R3222 GNDA.n255 GNDA.n254 29.0291
R3223 GNDA.n276 GNDA.n275 29.0291
R3224 GNDA.t221 GNDA.n369 28.9193
R3225 GNDA.t221 GNDA.t173 28.9193
R3226 GNDA.t39 GNDA.t206 28.9193
R3227 GNDA.t5 GNDA.t177 28.9193
R3228 GNDA.t221 GNDA.t107 28.9193
R3229 GNDA.n2470 GNDA.n330 28.8005
R3230 GNDA.n2454 GNDA.n337 28.8005
R3231 GNDA.n2713 GNDA.n39 28.8005
R3232 GNDA.n2691 GNDA.n50 28.8005
R3233 GNDA.n2669 GNDA.n61 28.8005
R3234 GNDA.n2651 GNDA.n2650 28.8005
R3235 GNDA.n2618 GNDA.n2617 28.8005
R3236 GNDA.n93 GNDA.n91 28.8005
R3237 GNDA.n2553 GNDA.n2552 28.8005
R3238 GNDA.n305 GNDA.n304 28.1695
R3239 GNDA.n1723 GNDA.n1722 27.5561
R3240 GNDA.n1534 GNDA.n1531 27.5561
R3241 GNDA.n540 GNDA.n539 27.5561
R3242 GNDA.n750 GNDA.n747 27.5561
R3243 GNDA.n977 GNDA.n974 27.5561
R3244 GNDA.n2185 GNDA.n2182 27.5561
R3245 GNDA.n2325 GNDA.n2324 27.5561
R3246 GNDA.n1277 GNDA.n1276 27.5561
R3247 GNDA.n2086 GNDA.n2083 27.5561
R3248 GNDA.n173 GNDA.n172 27.2005
R3249 GNDA.n178 GNDA.n123 27.2005
R3250 GNDA.n1096 GNDA.t101 26.976
R3251 GNDA.n1705 GNDA.n1704 26.6672
R3252 GNDA.n1515 GNDA.n1514 26.6672
R3253 GNDA.n522 GNDA.n521 26.6672
R3254 GNDA.n731 GNDA.n730 26.6672
R3255 GNDA.n958 GNDA.n957 26.6672
R3256 GNDA.n2166 GNDA.n2165 26.6672
R3257 GNDA.n2307 GNDA.n2306 26.6672
R3258 GNDA.n1260 GNDA.n1259 26.6672
R3259 GNDA.n2067 GNDA.n2066 26.6672
R3260 GNDA.n276 GNDA.n204 25.6005
R3261 GNDA.n246 GNDA.n245 25.6005
R3262 GNDA.n241 GNDA.n240 25.6005
R3263 GNDA.n307 GNDA.n306 25.6005
R3264 GNDA.n129 GNDA.n128 25.6005
R3265 GNDA.n310 GNDA.n117 25.6005
R3266 GNDA GNDA.n325 25.6005
R3267 GNDA.n2496 GNDA.n2495 25.6005
R3268 GNDA.n2523 GNDA.n96 25.6005
R3269 GNDA.n2774 GNDA.n20 25.6005
R3270 GNDA.n2787 GNDA.n2786 25.6005
R3271 GNDA.n2794 GNDA.n2793 25.6005
R3272 GNDA.n2808 GNDA.n2807 25.6005
R3273 GNDA.n334 GNDA.n332 25.6005
R3274 GNDA.n2443 GNDA.n2442 25.6005
R3275 GNDA.n2437 GNDA.n2436 25.6005
R3276 GNDA.n2423 GNDA.n2422 25.6005
R3277 GNDA.n2422 GNDA.n2421 25.6005
R3278 GNDA.n2704 GNDA.n45 25.6005
R3279 GNDA.n2682 GNDA.n56 25.6005
R3280 GNDA.n2660 GNDA.n67 25.6005
R3281 GNDA.n2638 GNDA.n2637 25.6005
R3282 GNDA.n2590 GNDA.n2589 25.6005
R3283 GNDA.n2574 GNDA.n2538 25.6005
R3284 GNDA.n2567 GNDA.n2566 25.6005
R3285 GNDA.n2559 GNDA.n2558 25.6005
R3286 GNDA.n2759 GNDA.n28 25.6005
R3287 GNDA.n1795 GNDA.n1794 25.3679
R3288 GNDA.t93 GNDA.t215 25.3526
R3289 GNDA.n193 GNDA.t195 25.2335
R3290 GNDA.n169 GNDA.n168 24.8279
R3291 GNDA.n303 GNDA.n115 24.8279
R3292 GNDA.t218 GNDA.t42 24.8125
R3293 GNDA.t139 GNDA.t267 24.8125
R3294 GNDA.t175 GNDA.t144 24.8125
R3295 GNDA.n133 GNDA.t259 24.0005
R3296 GNDA.n133 GNDA.t21 24.0005
R3297 GNDA.n137 GNDA.t130 24.0005
R3298 GNDA.n137 GNDA.t94 24.0005
R3299 GNDA.n141 GNDA.t128 24.0005
R3300 GNDA.n141 GNDA.t164 24.0005
R3301 GNDA.n143 GNDA.t83 24.0005
R3302 GNDA.n143 GNDA.t85 24.0005
R3303 GNDA.n314 GNDA.t304 24.0005
R3304 GNDA.n314 GNDA.t251 24.0005
R3305 GNDA.n2399 GNDA.t76 23.9787
R3306 GNDA.n2716 GNDA.n2715 23.1831
R3307 GNDA.t47 GNDA.t294 22.5646
R3308 GNDA.n304 GNDA.n302 22.5357
R3309 GNDA.n2809 GNDA.n2808 22.4005
R3310 GNDA.n2696 GNDA.n47 22.4005
R3311 GNDA.n2674 GNDA.n58 22.4005
R3312 GNDA.n2652 GNDA.n69 22.4005
R3313 GNDA.n87 GNDA.n84 22.4005
R3314 GNDA.n292 GNDA.n291 20.9665
R3315 GNDA.n2717 GNDA.n37 19.4625
R3316 GNDA.n267 GNDA.n213 19.2005
R3317 GNDA.n267 GNDA.n266 19.2005
R3318 GNDA.n2449 GNDA.n2448 19.2005
R3319 GNDA.n2707 GNDA.n2706 19.2005
R3320 GNDA.n2685 GNDA.n2684 19.2005
R3321 GNDA.n2663 GNDA.n2662 19.2005
R3322 GNDA.n77 GNDA.n74 19.2005
R3323 GNDA.n2625 GNDA.n2624 19.2005
R3324 GNDA.n2611 GNDA.n2610 19.2005
R3325 GNDA.n2585 GNDA.n2534 19.2005
R3326 GNDA.n2543 GNDA.n2540 19.2005
R3327 GNDA.n2759 GNDA.n2758 19.2005
R3328 GNDA.n1620 GNDA.n1455 17.5843
R3329 GNDA.n825 GNDA.n685 17.5843
R3330 GNDA.n1995 GNDA.n1061 17.5843
R3331 GNDA.t111 GNDA.t12 17.4653
R3332 GNDA.n1915 GNDA.n1914 16.9605
R3333 GNDA.n2234 GNDA.n640 16.9379
R3334 GNDA.n612 GNDA.n609 16.9379
R3335 GNDA.n1323 GNDA.n1293 16.9379
R3336 GNDA.n130 GNDA.t163 16.9019
R3337 GNDA.n913 GNDA.n912 16.7709
R3338 GNDA.n1178 GNDA.n437 16.7709
R3339 GNDA.n1421 GNDA.n434 16.7709
R3340 GNDA.n2393 GNDA.n405 16.7709
R3341 GNDA.t0 GNDA.t62 16.2817
R3342 GNDA.n2781 GNDA.n2780 16.0005
R3343 GNDA.n2782 GNDA.n2781 16.0005
R3344 GNDA.n1737 GNDA.n1723 16.0005
R3345 GNDA.n1737 GNDA.n1736 16.0005
R3346 GNDA.n1736 GNDA.n1735 16.0005
R3347 GNDA.n1735 GNDA.n1732 16.0005
R3348 GNDA.n1732 GNDA.n1731 16.0005
R3349 GNDA.n1731 GNDA.n1728 16.0005
R3350 GNDA.n1728 GNDA.n1727 16.0005
R3351 GNDA.n1727 GNDA.n1724 16.0005
R3352 GNDA.n1722 GNDA.n1720 16.0005
R3353 GNDA.n1720 GNDA.n1717 16.0005
R3354 GNDA.n1717 GNDA.n1716 16.0005
R3355 GNDA.n1716 GNDA.n1713 16.0005
R3356 GNDA.n1713 GNDA.n1712 16.0005
R3357 GNDA.n1712 GNDA.n1709 16.0005
R3358 GNDA.n1709 GNDA.n1708 16.0005
R3359 GNDA.n1708 GNDA.n1705 16.0005
R3360 GNDA.n1704 GNDA.n1701 16.0005
R3361 GNDA.n1701 GNDA.n1700 16.0005
R3362 GNDA.n1700 GNDA.n1697 16.0005
R3363 GNDA.n1697 GNDA.n1696 16.0005
R3364 GNDA.n1696 GNDA.n1693 16.0005
R3365 GNDA.n1693 GNDA.n1692 16.0005
R3366 GNDA.n1692 GNDA.n1689 16.0005
R3367 GNDA.n1689 GNDA.n1688 16.0005
R3368 GNDA.n1535 GNDA.n1534 16.0005
R3369 GNDA.n1538 GNDA.n1535 16.0005
R3370 GNDA.n1539 GNDA.n1538 16.0005
R3371 GNDA.n1542 GNDA.n1539 16.0005
R3372 GNDA.n1543 GNDA.n1542 16.0005
R3373 GNDA.n1546 GNDA.n1543 16.0005
R3374 GNDA.n1548 GNDA.n1546 16.0005
R3375 GNDA.n1549 GNDA.n1548 16.0005
R3376 GNDA.n1531 GNDA.n1530 16.0005
R3377 GNDA.n1530 GNDA.n1527 16.0005
R3378 GNDA.n1527 GNDA.n1526 16.0005
R3379 GNDA.n1526 GNDA.n1523 16.0005
R3380 GNDA.n1523 GNDA.n1522 16.0005
R3381 GNDA.n1522 GNDA.n1519 16.0005
R3382 GNDA.n1519 GNDA.n1518 16.0005
R3383 GNDA.n1518 GNDA.n1515 16.0005
R3384 GNDA.n1514 GNDA.n1511 16.0005
R3385 GNDA.n1511 GNDA.n1510 16.0005
R3386 GNDA.n1510 GNDA.n1507 16.0005
R3387 GNDA.n1507 GNDA.n1506 16.0005
R3388 GNDA.n1506 GNDA.n1503 16.0005
R3389 GNDA.n1503 GNDA.n1502 16.0005
R3390 GNDA.n1502 GNDA.n1499 16.0005
R3391 GNDA.n1499 GNDA.n1498 16.0005
R3392 GNDA.n554 GNDA.n540 16.0005
R3393 GNDA.n554 GNDA.n553 16.0005
R3394 GNDA.n553 GNDA.n552 16.0005
R3395 GNDA.n552 GNDA.n549 16.0005
R3396 GNDA.n549 GNDA.n548 16.0005
R3397 GNDA.n548 GNDA.n545 16.0005
R3398 GNDA.n545 GNDA.n544 16.0005
R3399 GNDA.n544 GNDA.n541 16.0005
R3400 GNDA.n539 GNDA.n537 16.0005
R3401 GNDA.n537 GNDA.n534 16.0005
R3402 GNDA.n534 GNDA.n533 16.0005
R3403 GNDA.n533 GNDA.n530 16.0005
R3404 GNDA.n530 GNDA.n529 16.0005
R3405 GNDA.n529 GNDA.n526 16.0005
R3406 GNDA.n526 GNDA.n525 16.0005
R3407 GNDA.n525 GNDA.n522 16.0005
R3408 GNDA.n521 GNDA.n518 16.0005
R3409 GNDA.n518 GNDA.n517 16.0005
R3410 GNDA.n517 GNDA.n514 16.0005
R3411 GNDA.n514 GNDA.n513 16.0005
R3412 GNDA.n513 GNDA.n510 16.0005
R3413 GNDA.n510 GNDA.n509 16.0005
R3414 GNDA.n509 GNDA.n506 16.0005
R3415 GNDA.n506 GNDA.n505 16.0005
R3416 GNDA.n751 GNDA.n750 16.0005
R3417 GNDA.n754 GNDA.n751 16.0005
R3418 GNDA.n755 GNDA.n754 16.0005
R3419 GNDA.n758 GNDA.n755 16.0005
R3420 GNDA.n759 GNDA.n758 16.0005
R3421 GNDA.n762 GNDA.n759 16.0005
R3422 GNDA.n763 GNDA.n762 16.0005
R3423 GNDA.n763 GNDA.n443 16.0005
R3424 GNDA.n747 GNDA.n746 16.0005
R3425 GNDA.n746 GNDA.n743 16.0005
R3426 GNDA.n743 GNDA.n742 16.0005
R3427 GNDA.n742 GNDA.n739 16.0005
R3428 GNDA.n739 GNDA.n738 16.0005
R3429 GNDA.n738 GNDA.n735 16.0005
R3430 GNDA.n735 GNDA.n734 16.0005
R3431 GNDA.n734 GNDA.n731 16.0005
R3432 GNDA.n730 GNDA.n727 16.0005
R3433 GNDA.n727 GNDA.n726 16.0005
R3434 GNDA.n726 GNDA.n723 16.0005
R3435 GNDA.n723 GNDA.n722 16.0005
R3436 GNDA.n722 GNDA.n719 16.0005
R3437 GNDA.n719 GNDA.n718 16.0005
R3438 GNDA.n718 GNDA.n715 16.0005
R3439 GNDA.n715 GNDA.n693 16.0005
R3440 GNDA.n978 GNDA.n977 16.0005
R3441 GNDA.n981 GNDA.n978 16.0005
R3442 GNDA.n982 GNDA.n981 16.0005
R3443 GNDA.n985 GNDA.n982 16.0005
R3444 GNDA.n986 GNDA.n985 16.0005
R3445 GNDA.n989 GNDA.n986 16.0005
R3446 GNDA.n991 GNDA.n989 16.0005
R3447 GNDA.n992 GNDA.n991 16.0005
R3448 GNDA.n974 GNDA.n973 16.0005
R3449 GNDA.n973 GNDA.n970 16.0005
R3450 GNDA.n970 GNDA.n969 16.0005
R3451 GNDA.n969 GNDA.n966 16.0005
R3452 GNDA.n966 GNDA.n965 16.0005
R3453 GNDA.n965 GNDA.n962 16.0005
R3454 GNDA.n962 GNDA.n961 16.0005
R3455 GNDA.n961 GNDA.n958 16.0005
R3456 GNDA.n957 GNDA.n954 16.0005
R3457 GNDA.n954 GNDA.n953 16.0005
R3458 GNDA.n953 GNDA.n950 16.0005
R3459 GNDA.n950 GNDA.n949 16.0005
R3460 GNDA.n949 GNDA.n946 16.0005
R3461 GNDA.n946 GNDA.n945 16.0005
R3462 GNDA.n945 GNDA.n942 16.0005
R3463 GNDA.n942 GNDA.n918 16.0005
R3464 GNDA.n2186 GNDA.n2185 16.0005
R3465 GNDA.n2189 GNDA.n2186 16.0005
R3466 GNDA.n2190 GNDA.n2189 16.0005
R3467 GNDA.n2193 GNDA.n2190 16.0005
R3468 GNDA.n2194 GNDA.n2193 16.0005
R3469 GNDA.n2197 GNDA.n2194 16.0005
R3470 GNDA.n2198 GNDA.n2197 16.0005
R3471 GNDA.n2201 GNDA.n2198 16.0005
R3472 GNDA.n2182 GNDA.n2181 16.0005
R3473 GNDA.n2181 GNDA.n2178 16.0005
R3474 GNDA.n2178 GNDA.n2177 16.0005
R3475 GNDA.n2177 GNDA.n2174 16.0005
R3476 GNDA.n2174 GNDA.n2173 16.0005
R3477 GNDA.n2173 GNDA.n2170 16.0005
R3478 GNDA.n2170 GNDA.n2169 16.0005
R3479 GNDA.n2169 GNDA.n2166 16.0005
R3480 GNDA.n2165 GNDA.n2162 16.0005
R3481 GNDA.n2162 GNDA.n2161 16.0005
R3482 GNDA.n2161 GNDA.n2158 16.0005
R3483 GNDA.n2158 GNDA.n2157 16.0005
R3484 GNDA.n2157 GNDA.n2154 16.0005
R3485 GNDA.n2154 GNDA.n2153 16.0005
R3486 GNDA.n2153 GNDA.n2150 16.0005
R3487 GNDA.n2150 GNDA.n2149 16.0005
R3488 GNDA.n2338 GNDA.n2325 16.0005
R3489 GNDA.n2338 GNDA.n2337 16.0005
R3490 GNDA.n2337 GNDA.n2336 16.0005
R3491 GNDA.n2336 GNDA.n2333 16.0005
R3492 GNDA.n2333 GNDA.n2332 16.0005
R3493 GNDA.n2332 GNDA.n2329 16.0005
R3494 GNDA.n2329 GNDA.n2328 16.0005
R3495 GNDA.n2328 GNDA.n2241 16.0005
R3496 GNDA.n2324 GNDA.n2322 16.0005
R3497 GNDA.n2322 GNDA.n2319 16.0005
R3498 GNDA.n2319 GNDA.n2318 16.0005
R3499 GNDA.n2318 GNDA.n2315 16.0005
R3500 GNDA.n2315 GNDA.n2314 16.0005
R3501 GNDA.n2314 GNDA.n2311 16.0005
R3502 GNDA.n2311 GNDA.n2310 16.0005
R3503 GNDA.n2310 GNDA.n2307 16.0005
R3504 GNDA.n2306 GNDA.n2303 16.0005
R3505 GNDA.n2303 GNDA.n2302 16.0005
R3506 GNDA.n2302 GNDA.n2299 16.0005
R3507 GNDA.n2299 GNDA.n2298 16.0005
R3508 GNDA.n2298 GNDA.n2295 16.0005
R3509 GNDA.n2295 GNDA.n2294 16.0005
R3510 GNDA.n2294 GNDA.n2291 16.0005
R3511 GNDA.n2291 GNDA.n2290 16.0005
R3512 GNDA.n1277 GNDA.n1235 16.0005
R3513 GNDA.n1283 GNDA.n1235 16.0005
R3514 GNDA.n1284 GNDA.n1283 16.0005
R3515 GNDA.n1285 GNDA.n1284 16.0005
R3516 GNDA.n1285 GNDA.n1233 16.0005
R3517 GNDA.n1291 GNDA.n1233 16.0005
R3518 GNDA.n1292 GNDA.n1291 16.0005
R3519 GNDA.n1350 GNDA.n1292 16.0005
R3520 GNDA.n1276 GNDA.n1275 16.0005
R3521 GNDA.n1275 GNDA.n1237 16.0005
R3522 GNDA.n1269 GNDA.n1237 16.0005
R3523 GNDA.n1269 GNDA.n1268 16.0005
R3524 GNDA.n1268 GNDA.n1267 16.0005
R3525 GNDA.n1267 GNDA.n1239 16.0005
R3526 GNDA.n1261 GNDA.n1239 16.0005
R3527 GNDA.n1261 GNDA.n1260 16.0005
R3528 GNDA.n1259 GNDA.n1241 16.0005
R3529 GNDA.n1253 GNDA.n1241 16.0005
R3530 GNDA.n1253 GNDA.n1252 16.0005
R3531 GNDA.n1252 GNDA.n1251 16.0005
R3532 GNDA.n1251 GNDA.n1243 16.0005
R3533 GNDA.n1246 GNDA.n1243 16.0005
R3534 GNDA.n1246 GNDA.n1217 16.0005
R3535 GNDA.n1386 GNDA.n1217 16.0005
R3536 GNDA.n2087 GNDA.n2086 16.0005
R3537 GNDA.n2090 GNDA.n2087 16.0005
R3538 GNDA.n2091 GNDA.n2090 16.0005
R3539 GNDA.n2094 GNDA.n2091 16.0005
R3540 GNDA.n2095 GNDA.n2094 16.0005
R3541 GNDA.n2098 GNDA.n2095 16.0005
R3542 GNDA.n2099 GNDA.n2098 16.0005
R3543 GNDA.n2099 GNDA.n1034 16.0005
R3544 GNDA.n2083 GNDA.n2082 16.0005
R3545 GNDA.n2082 GNDA.n2079 16.0005
R3546 GNDA.n2079 GNDA.n2078 16.0005
R3547 GNDA.n2078 GNDA.n2075 16.0005
R3548 GNDA.n2075 GNDA.n2074 16.0005
R3549 GNDA.n2074 GNDA.n2071 16.0005
R3550 GNDA.n2071 GNDA.n2070 16.0005
R3551 GNDA.n2070 GNDA.n2067 16.0005
R3552 GNDA.n2066 GNDA.n2063 16.0005
R3553 GNDA.n2063 GNDA.n2062 16.0005
R3554 GNDA.n2062 GNDA.n2059 16.0005
R3555 GNDA.n2059 GNDA.n2058 16.0005
R3556 GNDA.n2058 GNDA.n2055 16.0005
R3557 GNDA.n2055 GNDA.n2054 16.0005
R3558 GNDA.n2054 GNDA.n2051 16.0005
R3559 GNDA.n2051 GNDA.n2050 16.0005
R3560 GNDA.n2599 GNDA.n2598 16.0005
R3561 GNDA.n2598 GNDA.n2597 16.0005
R3562 GNDA.n326 GNDA 15.7005
R3563 GNDA.n293 GNDA.n292 15.6449
R3564 GNDA.n2482 GNDA.n2481 15.6449
R3565 GNDA.n281 GNDA.t31 15.0005
R3566 GNDA.n281 GNDA.t255 15.0005
R3567 GNDA.n289 GNDA.t226 15.0005
R3568 GNDA.n289 GNDA.t184 15.0005
R3569 GNDA.t219 GNDA.n268 15.0005
R3570 GNDA.n268 GNDA.t166 15.0005
R3571 GNDA.n218 GNDA.t168 15.0005
R3572 GNDA.n218 GNDA.t247 15.0005
R3573 GNDA.t268 GNDA.n247 15.0005
R3574 GNDA.n247 GNDA.t145 15.0005
R3575 GNDA.n239 GNDA.t157 15.0005
R3576 GNDA.n239 GNDA.t243 15.0005
R3577 GNDA.n248 GNDA.t268 15.0005
R3578 GNDA.n223 GNDA.t248 15.0005
R3579 GNDA.n269 GNDA.t219 15.0005
R3580 GNDA.n206 GNDA.t256 15.0005
R3581 GNDA.t226 GNDA.n198 15.0005
R3582 GNDA.n110 GNDA.t244 15.0005
R3583 GNDA.n2210 GNDA.n374 14.555
R3584 GNDA.n2357 GNDA.n375 14.555
R3585 GNDA.n2481 GNDA.n2480 14.4005
R3586 GNDA.n174 GNDA.n173 14.0805
R3587 GNDA.n176 GNDA.n123 14.0805
R3588 GNDA.n2495 GNDA.n105 13.9181
R3589 GNDA.t303 GNDA.t111 13.5216
R3590 GNDA.n2475 GNDA.n2474 12.8163
R3591 GNDA.n276 GNDA.n202 12.8005
R3592 GNDA.n290 GNDA.n288 12.8005
R3593 GNDA.n246 GNDA.n232 12.8005
R3594 GNDA.n240 GNDA.n111 12.8005
R3595 GNDA.n308 GNDA.n307 12.8005
R3596 GNDA.n128 GNDA.n121 12.8005
R3597 GNDA.n1679 GNDA.n1678 12.8005
R3598 GNDA.n1678 GNDA.n1675 12.8005
R3599 GNDA.n1763 GNDA.n1110 12.8005
R3600 GNDA.n1759 GNDA.n1110 12.8005
R3601 GNDA.n2449 GNDA.n338 12.8005
R3602 GNDA.n1813 GNDA.n1083 12.8005
R3603 GNDA.n1915 GNDA.n1083 12.8005
R3604 GNDA.n2706 GNDA.n2705 12.8005
R3605 GNDA.n2684 GNDA.n2683 12.8005
R3606 GNDA.n2662 GNDA.n2661 12.8005
R3607 GNDA.n2639 GNDA.n77 12.8005
R3608 GNDA.n2626 GNDA.n2625 12.8005
R3609 GNDA.n2612 GNDA.n2611 12.8005
R3610 GNDA.n2534 GNDA.n2531 12.8005
R3611 GNDA.n2568 GNDA.n2543 12.8005
R3612 GNDA.n2731 GNDA.n2730 12.8005
R3613 GNDA.n2723 GNDA.n35 12.8005
R3614 GNDA GNDA.n0 12.7806
R3615 GNDA GNDA.n2823 11.8829
R3616 GNDA.n105 GNDA.n37 11.7212
R3617 GNDA.n327 GNDA.n326 11.6918
R3618 GNDA.n2477 GNDA.n2476 11.6542
R3619 GNDA.n1636 GNDA.n1447 11.6369
R3620 GNDA.n1636 GNDA.n1635 11.6369
R3621 GNDA.n1635 GNDA.n1634 11.6369
R3622 GNDA.n1634 GNDA.n1449 11.6369
R3623 GNDA.n1629 GNDA.n1449 11.6369
R3624 GNDA.n1629 GNDA.n1628 11.6369
R3625 GNDA.n1628 GNDA.n1627 11.6369
R3626 GNDA.n1627 GNDA.n1452 11.6369
R3627 GNDA.n1622 GNDA.n1452 11.6369
R3628 GNDA.n1622 GNDA.n1621 11.6369
R3629 GNDA.n1621 GNDA.n1620 11.6369
R3630 GNDA.n1615 GNDA.n1455 11.6369
R3631 GNDA.n1615 GNDA.n1614 11.6369
R3632 GNDA.n1614 GNDA.n1613 11.6369
R3633 GNDA.n1613 GNDA.n1458 11.6369
R3634 GNDA.n1608 GNDA.n1458 11.6369
R3635 GNDA.n1608 GNDA.n1607 11.6369
R3636 GNDA.n1607 GNDA.n1606 11.6369
R3637 GNDA.n1606 GNDA.n1461 11.6369
R3638 GNDA.n1601 GNDA.n1461 11.6369
R3639 GNDA.n1601 GNDA.n1600 11.6369
R3640 GNDA.n820 GNDA.n685 11.6369
R3641 GNDA.n820 GNDA.n819 11.6369
R3642 GNDA.n819 GNDA.n818 11.6369
R3643 GNDA.n818 GNDA.n687 11.6369
R3644 GNDA.n813 GNDA.n687 11.6369
R3645 GNDA.n813 GNDA.n812 11.6369
R3646 GNDA.n812 GNDA.n811 11.6369
R3647 GNDA.n811 GNDA.n690 11.6369
R3648 GNDA.n806 GNDA.n690 11.6369
R3649 GNDA.n806 GNDA.n805 11.6369
R3650 GNDA.n846 GNDA.n845 11.6369
R3651 GNDA.n845 GNDA.n842 11.6369
R3652 GNDA.n842 GNDA.n841 11.6369
R3653 GNDA.n841 GNDA.n838 11.6369
R3654 GNDA.n838 GNDA.n837 11.6369
R3655 GNDA.n837 GNDA.n834 11.6369
R3656 GNDA.n834 GNDA.n833 11.6369
R3657 GNDA.n833 GNDA.n830 11.6369
R3658 GNDA.n830 GNDA.n829 11.6369
R3659 GNDA.n829 GNDA.n826 11.6369
R3660 GNDA.n826 GNDA.n825 11.6369
R3661 GNDA.n847 GNDA.n404 11.6369
R3662 GNDA.n850 GNDA.n847 11.6369
R3663 GNDA.n851 GNDA.n850 11.6369
R3664 GNDA.n854 GNDA.n851 11.6369
R3665 GNDA.n855 GNDA.n854 11.6369
R3666 GNDA.n858 GNDA.n855 11.6369
R3667 GNDA.n859 GNDA.n858 11.6369
R3668 GNDA.n862 GNDA.n859 11.6369
R3669 GNDA.n863 GNDA.n862 11.6369
R3670 GNDA.n866 GNDA.n863 11.6369
R3671 GNDA.n867 GNDA.n866 11.6369
R3672 GNDA.n1879 GNDA.n640 11.6369
R3673 GNDA.n1880 GNDA.n1879 11.6369
R3674 GNDA.n1881 GNDA.n1880 11.6369
R3675 GNDA.n1881 GNDA.n1873 11.6369
R3676 GNDA.n1887 GNDA.n1873 11.6369
R3677 GNDA.n1888 GNDA.n1887 11.6369
R3678 GNDA.n1889 GNDA.n1888 11.6369
R3679 GNDA.n1889 GNDA.n1869 11.6369
R3680 GNDA.n1895 GNDA.n1869 11.6369
R3681 GNDA.n1896 GNDA.n1895 11.6369
R3682 GNDA.n1897 GNDA.n1896 11.6369
R3683 GNDA.n2234 GNDA.n2233 11.6369
R3684 GNDA.n2233 GNDA.n2232 11.6369
R3685 GNDA.n2232 GNDA.n2231 11.6369
R3686 GNDA.n2231 GNDA.n2229 11.6369
R3687 GNDA.n2229 GNDA.n2226 11.6369
R3688 GNDA.n2226 GNDA.n2225 11.6369
R3689 GNDA.n2225 GNDA.n2222 11.6369
R3690 GNDA.n2222 GNDA.n2221 11.6369
R3691 GNDA.n2221 GNDA.n2218 11.6369
R3692 GNDA.n2218 GNDA.n2217 11.6369
R3693 GNDA.n609 GNDA.n608 11.6369
R3694 GNDA.n608 GNDA.n605 11.6369
R3695 GNDA.n605 GNDA.n604 11.6369
R3696 GNDA.n604 GNDA.n601 11.6369
R3697 GNDA.n601 GNDA.n600 11.6369
R3698 GNDA.n600 GNDA.n597 11.6369
R3699 GNDA.n597 GNDA.n596 11.6369
R3700 GNDA.n596 GNDA.n593 11.6369
R3701 GNDA.n593 GNDA.n592 11.6369
R3702 GNDA.n592 GNDA.n403 11.6369
R3703 GNDA.n2394 GNDA.n403 11.6369
R3704 GNDA.n613 GNDA.n612 11.6369
R3705 GNDA.n616 GNDA.n613 11.6369
R3706 GNDA.n617 GNDA.n616 11.6369
R3707 GNDA.n620 GNDA.n617 11.6369
R3708 GNDA.n621 GNDA.n620 11.6369
R3709 GNDA.n624 GNDA.n621 11.6369
R3710 GNDA.n625 GNDA.n624 11.6369
R3711 GNDA.n627 GNDA.n625 11.6369
R3712 GNDA.n627 GNDA.n626 11.6369
R3713 GNDA.n626 GNDA.n578 11.6369
R3714 GNDA.n1324 GNDA.n1323 11.6369
R3715 GNDA.n1327 GNDA.n1324 11.6369
R3716 GNDA.n1328 GNDA.n1327 11.6369
R3717 GNDA.n1331 GNDA.n1328 11.6369
R3718 GNDA.n1332 GNDA.n1331 11.6369
R3719 GNDA.n1335 GNDA.n1332 11.6369
R3720 GNDA.n1336 GNDA.n1335 11.6369
R3721 GNDA.n1339 GNDA.n1336 11.6369
R3722 GNDA.n1341 GNDA.n1339 11.6369
R3723 GNDA.n1342 GNDA.n1341 11.6369
R3724 GNDA.n1996 GNDA.n1995 11.6369
R3725 GNDA.n1997 GNDA.n1996 11.6369
R3726 GNDA.n1997 GNDA.n1059 11.6369
R3727 GNDA.n2003 GNDA.n1059 11.6369
R3728 GNDA.n2004 GNDA.n2003 11.6369
R3729 GNDA.n2005 GNDA.n2004 11.6369
R3730 GNDA.n2005 GNDA.n1057 11.6369
R3731 GNDA.n2011 GNDA.n1057 11.6369
R3732 GNDA.n2012 GNDA.n2011 11.6369
R3733 GNDA.n2013 GNDA.n2012 11.6369
R3734 GNDA.n1969 GNDA.n1070 11.6369
R3735 GNDA.n1975 GNDA.n1070 11.6369
R3736 GNDA.n1976 GNDA.n1975 11.6369
R3737 GNDA.n1977 GNDA.n1976 11.6369
R3738 GNDA.n1977 GNDA.n1066 11.6369
R3739 GNDA.n1983 GNDA.n1066 11.6369
R3740 GNDA.n1984 GNDA.n1983 11.6369
R3741 GNDA.n1986 GNDA.n1984 11.6369
R3742 GNDA.n1986 GNDA.n1985 11.6369
R3743 GNDA.n1985 GNDA.n1063 11.6369
R3744 GNDA.n1063 GNDA.n1061 11.6369
R3745 GNDA.n1904 GNDA.n1903 11.6369
R3746 GNDA.n1906 GNDA.n1904 11.6369
R3747 GNDA.n1906 GNDA.n1905 11.6369
R3748 GNDA.n1905 GNDA.n1818 11.6369
R3749 GNDA.n1913 GNDA.n1818 11.6369
R3750 GNDA.n1920 GNDA.n1078 11.6369
R3751 GNDA.n1921 GNDA.n1920 11.6369
R3752 GNDA.n1923 GNDA.n1921 11.6369
R3753 GNDA.n1923 GNDA.n1922 11.6369
R3754 GNDA.n1922 GNDA.n1074 11.6369
R3755 GNDA.n1422 GNDA.n1184 11.6369
R3756 GNDA.n1428 GNDA.n1184 11.6369
R3757 GNDA.n1429 GNDA.n1428 11.6369
R3758 GNDA.n1430 GNDA.n1429 11.6369
R3759 GNDA.n1430 GNDA.n1182 11.6369
R3760 GNDA.n1436 GNDA.n1182 11.6369
R3761 GNDA.n1437 GNDA.n1436 11.6369
R3762 GNDA.n1438 GNDA.n1437 11.6369
R3763 GNDA.n1438 GNDA.n1180 11.6369
R3764 GNDA.n1443 GNDA.n1180 11.6369
R3765 GNDA.n1444 GNDA.n1443 11.6369
R3766 GNDA.n1318 GNDA.n1293 11.6369
R3767 GNDA.n1318 GNDA.n1317 11.6369
R3768 GNDA.n1317 GNDA.n1316 11.6369
R3769 GNDA.n1316 GNDA.n1295 11.6369
R3770 GNDA.n1311 GNDA.n1295 11.6369
R3771 GNDA.n1311 GNDA.n1310 11.6369
R3772 GNDA.n1310 GNDA.n1309 11.6369
R3773 GNDA.n1309 GNDA.n1298 11.6369
R3774 GNDA.n1304 GNDA.n1298 11.6369
R3775 GNDA.n1304 GNDA.n1303 11.6369
R3776 GNDA.n1303 GNDA.n1186 11.6369
R3777 GNDA.n2771 GNDA.t202 11.2826
R3778 GNDA.n2770 GNDA.t71 11.2826
R3779 GNDA.n2715 GNDA.n39 10.7016
R3780 GNDA.n2552 GNDA.n2551 10.4505
R3781 GNDA.t38 GNDA.n1360 10.1221
R3782 GNDA.t32 GNDA.n1375 10.1221
R3783 GNDA.n1376 GNDA.t26 10.1221
R3784 GNDA.t24 GNDA.n1392 10.1221
R3785 GNDA.n2810 GNDA.n2809 9.6005
R3786 GNDA.n1781 GNDA.t182 9.6005
R3787 GNDA.n1774 GNDA.t178 9.6005
R3788 GNDA.n1793 GNDA.t209 9.6005
R3789 GNDA.n1796 GNDA.t207 9.6005
R3790 GNDA.n2699 GNDA.n47 9.6005
R3791 GNDA.n2677 GNDA.n58 9.6005
R3792 GNDA.n2655 GNDA.n69 9.6005
R3793 GNDA.n2619 GNDA.n87 9.6005
R3794 GNDA.n168 GNDA.n167 9.58175
R3795 GNDA.n321 GNDA.n115 9.58175
R3796 GNDA.n193 GNDA.t118 9.46287
R3797 GNDA.n1679 GNDA.n1674 9.36264
R3798 GNDA.n1759 GNDA.n1108 9.36264
R3799 GNDA.n1814 GNDA.n1813 9.36264
R3800 GNDA.n166 GNDA.n165 9.3005
R3801 GNDA.n164 GNDA.n131 9.3005
R3802 GNDA.n163 GNDA.n162 9.3005
R3803 GNDA.n161 GNDA.n132 9.3005
R3804 GNDA.n160 GNDA.n159 9.3005
R3805 GNDA.n158 GNDA.n135 9.3005
R3806 GNDA.n157 GNDA.n156 9.3005
R3807 GNDA.n155 GNDA.n136 9.3005
R3808 GNDA.n154 GNDA.n153 9.3005
R3809 GNDA.n152 GNDA.n139 9.3005
R3810 GNDA.n151 GNDA.n150 9.3005
R3811 GNDA.n149 GNDA.n140 9.3005
R3812 GNDA.n148 GNDA.n147 9.3005
R3813 GNDA.n146 GNDA.n145 9.3005
R3814 GNDA.n119 GNDA.n118 9.3005
R3815 GNDA.n312 GNDA.n311 9.3005
R3816 GNDA.n313 GNDA.n117 9.3005
R3817 GNDA.n317 GNDA.n316 9.3005
R3818 GNDA.n318 GNDA.n116 9.3005
R3819 GNDA.n320 GNDA.n319 9.3005
R3820 GNDA.n322 GNDA.n114 9.3005
R3821 GNDA.n324 GNDA.n323 9.3005
R3822 GNDA.n325 GNDA.n113 9.3005
R3823 GNDA.n1678 GNDA.n1677 9.3005
R3824 GNDA.n1676 GNDA.n1675 9.3005
R3825 GNDA.n1110 GNDA.n1109 9.3005
R3826 GNDA.n1764 GNDA.n1763 9.3005
R3827 GNDA.n2473 GNDA.n2472 9.3005
R3828 GNDA.n2471 GNDA.n329 9.3005
R3829 GNDA.n2470 GNDA.n2469 9.3005
R3830 GNDA.n2468 GNDA.n2467 9.3005
R3831 GNDA.n2466 GNDA.n331 9.3005
R3832 GNDA.n2465 GNDA.n2464 9.3005
R3833 GNDA.n2463 GNDA.n332 9.3005
R3834 GNDA.n2462 GNDA.n2461 9.3005
R3835 GNDA.n2460 GNDA.n333 9.3005
R3836 GNDA.n2459 GNDA.n2458 9.3005
R3837 GNDA.n2457 GNDA.n335 9.3005
R3838 GNDA.n2456 GNDA.n2455 9.3005
R3839 GNDA.n337 GNDA.n336 9.3005
R3840 GNDA.n341 GNDA.n340 9.3005
R3841 GNDA.n342 GNDA.n338 9.3005
R3842 GNDA.n2448 GNDA.n2447 9.3005
R3843 GNDA.n2446 GNDA.n339 9.3005
R3844 GNDA.n2445 GNDA.n2444 9.3005
R3845 GNDA.n2443 GNDA.n343 9.3005
R3846 GNDA.n2441 GNDA.n2440 9.3005
R3847 GNDA.n2439 GNDA.n345 9.3005
R3848 GNDA.n2438 GNDA.n2437 9.3005
R3849 GNDA.n2435 GNDA.n346 9.3005
R3850 GNDA.n2434 GNDA.n2433 9.3005
R3851 GNDA.n2432 GNDA.n348 9.3005
R3852 GNDA.n2431 GNDA.n2430 9.3005
R3853 GNDA.n2429 GNDA.n349 9.3005
R3854 GNDA.n2428 GNDA.n2427 9.3005
R3855 GNDA.n2426 GNDA.n350 9.3005
R3856 GNDA.n2425 GNDA.n2424 9.3005
R3857 GNDA.n2422 GNDA.n351 9.3005
R3858 GNDA.n2420 GNDA.n2419 9.3005
R3859 GNDA.n2418 GNDA.n354 9.3005
R3860 GNDA.n2417 GNDA.n2416 9.3005
R3861 GNDA.n2415 GNDA.n355 9.3005
R3862 GNDA.n2414 GNDA.n2413 9.3005
R3863 GNDA.n2412 GNDA.n356 9.3005
R3864 GNDA.n2411 GNDA.n2410 9.3005
R3865 GNDA.n2409 GNDA.n357 9.3005
R3866 GNDA.n1084 GNDA.n1083 9.3005
R3867 GNDA.n1915 GNDA.n1817 9.3005
R3868 GNDA.n2553 GNDA.n2548 9.3005
R3869 GNDA.n2555 GNDA.n2554 9.3005
R3870 GNDA.n2556 GNDA.n2547 9.3005
R3871 GNDA.n2558 GNDA.n2557 9.3005
R3872 GNDA.n2560 GNDA.n2546 9.3005
R3873 GNDA.n2562 GNDA.n2561 9.3005
R3874 GNDA.n2563 GNDA.n2545 9.3005
R3875 GNDA.n2565 GNDA.n2564 9.3005
R3876 GNDA.n2567 GNDA.n2541 9.3005
R3877 GNDA.n2569 GNDA.n2568 9.3005
R3878 GNDA.n2570 GNDA.n2540 9.3005
R3879 GNDA.n2572 GNDA.n2571 9.3005
R3880 GNDA.n2573 GNDA.n2539 9.3005
R3881 GNDA.n2575 GNDA.n2574 9.3005
R3882 GNDA.n2577 GNDA.n2576 9.3005
R3883 GNDA.n2578 GNDA.n2536 9.3005
R3884 GNDA.n2580 GNDA.n2579 9.3005
R3885 GNDA.n2581 GNDA.n2535 9.3005
R3886 GNDA.n2583 GNDA.n2582 9.3005
R3887 GNDA.n2584 GNDA.n2532 9.3005
R3888 GNDA.n2586 GNDA.n2585 9.3005
R3889 GNDA.n2587 GNDA.n2531 9.3005
R3890 GNDA.n2589 GNDA.n2588 9.3005
R3891 GNDA.n2591 GNDA.n2529 9.3005
R3892 GNDA.n2593 GNDA.n2592 9.3005
R3893 GNDA.n2594 GNDA.n2528 9.3005
R3894 GNDA.n2596 GNDA.n2595 9.3005
R3895 GNDA.n2597 GNDA.n95 9.3005
R3896 GNDA.n2600 GNDA.n2599 9.3005
R3897 GNDA.n2601 GNDA.n94 9.3005
R3898 GNDA.n2603 GNDA.n2602 9.3005
R3899 GNDA.n2604 GNDA.n92 9.3005
R3900 GNDA.n2606 GNDA.n2605 9.3005
R3901 GNDA.n2607 GNDA.n91 9.3005
R3902 GNDA.n2609 GNDA.n2608 9.3005
R3903 GNDA.n2610 GNDA.n90 9.3005
R3904 GNDA.n2613 GNDA.n2612 9.3005
R3905 GNDA.n2614 GNDA.n89 9.3005
R3906 GNDA.n2616 GNDA.n2615 9.3005
R3907 GNDA.n2618 GNDA.n85 9.3005
R3908 GNDA.n2620 GNDA.n2619 9.3005
R3909 GNDA.n2621 GNDA.n84 9.3005
R3910 GNDA.n2623 GNDA.n2622 9.3005
R3911 GNDA.n2624 GNDA.n82 9.3005
R3912 GNDA.n2627 GNDA.n2626 9.3005
R3913 GNDA.n2628 GNDA.n81 9.3005
R3914 GNDA.n2630 GNDA.n2629 9.3005
R3915 GNDA.n2631 GNDA.n80 9.3005
R3916 GNDA.n2633 GNDA.n2632 9.3005
R3917 GNDA.n2634 GNDA.n79 9.3005
R3918 GNDA.n2636 GNDA.n2635 9.3005
R3919 GNDA.n2638 GNDA.n75 9.3005
R3920 GNDA.n2640 GNDA.n2639 9.3005
R3921 GNDA.n2641 GNDA.n74 9.3005
R3922 GNDA.n2643 GNDA.n2642 9.3005
R3923 GNDA.n2644 GNDA.n73 9.3005
R3924 GNDA.n2646 GNDA.n2645 9.3005
R3925 GNDA.n2647 GNDA.n72 9.3005
R3926 GNDA.n2649 GNDA.n2648 9.3005
R3927 GNDA.n2651 GNDA.n70 9.3005
R3928 GNDA.n2653 GNDA.n2652 9.3005
R3929 GNDA.n2655 GNDA.n2654 9.3005
R3930 GNDA.n2656 GNDA.n68 9.3005
R3931 GNDA.n2658 GNDA.n2657 9.3005
R3932 GNDA.n2660 GNDA.n2659 9.3005
R3933 GNDA.n2661 GNDA.n64 9.3005
R3934 GNDA.n2664 GNDA.n2663 9.3005
R3935 GNDA.n2665 GNDA.n63 9.3005
R3936 GNDA.n2667 GNDA.n2666 9.3005
R3937 GNDA.n2668 GNDA.n62 9.3005
R3938 GNDA.n2670 GNDA.n2669 9.3005
R3939 GNDA.n2672 GNDA.n2671 9.3005
R3940 GNDA.n2673 GNDA.n59 9.3005
R3941 GNDA.n2675 GNDA.n2674 9.3005
R3942 GNDA.n2677 GNDA.n2676 9.3005
R3943 GNDA.n2678 GNDA.n57 9.3005
R3944 GNDA.n2680 GNDA.n2679 9.3005
R3945 GNDA.n2682 GNDA.n2681 9.3005
R3946 GNDA.n2683 GNDA.n53 9.3005
R3947 GNDA.n2686 GNDA.n2685 9.3005
R3948 GNDA.n2687 GNDA.n52 9.3005
R3949 GNDA.n2689 GNDA.n2688 9.3005
R3950 GNDA.n2690 GNDA.n51 9.3005
R3951 GNDA.n2692 GNDA.n2691 9.3005
R3952 GNDA.n2694 GNDA.n2693 9.3005
R3953 GNDA.n2695 GNDA.n48 9.3005
R3954 GNDA.n2697 GNDA.n2696 9.3005
R3955 GNDA.n2699 GNDA.n2698 9.3005
R3956 GNDA.n2700 GNDA.n46 9.3005
R3957 GNDA.n2702 GNDA.n2701 9.3005
R3958 GNDA.n2704 GNDA.n2703 9.3005
R3959 GNDA.n2705 GNDA.n42 9.3005
R3960 GNDA.n2708 GNDA.n2707 9.3005
R3961 GNDA.n2709 GNDA.n41 9.3005
R3962 GNDA.n2711 GNDA.n2710 9.3005
R3963 GNDA.n2712 GNDA.n40 9.3005
R3964 GNDA.n2714 GNDA.n2713 9.3005
R3965 GNDA.n2739 GNDA.n28 9.3005
R3966 GNDA.n2738 GNDA.n2737 9.3005
R3967 GNDA.n2736 GNDA.n29 9.3005
R3968 GNDA.n2735 GNDA.n2734 9.3005
R3969 GNDA.n2733 GNDA.n30 9.3005
R3970 GNDA.n2732 GNDA.n2731 9.3005
R3971 GNDA.n2730 GNDA.n31 9.3005
R3972 GNDA.n2729 GNDA.n2728 9.3005
R3973 GNDA.n2727 GNDA.n33 9.3005
R3974 GNDA.n2726 GNDA.n2725 9.3005
R3975 GNDA.n2724 GNDA.n34 9.3005
R3976 GNDA.n2723 GNDA.n2722 9.3005
R3977 GNDA.n2718 GNDA.n36 9.3005
R3978 GNDA.n2720 GNDA.n2719 9.3005
R3979 GNDA.n2721 GNDA.n35 9.3005
R3980 GNDA.n2759 GNDA.n2740 9.3005
R3981 GNDA.n2747 GNDA.n2744 9.3005
R3982 GNDA.n2749 GNDA.n2748 9.3005
R3983 GNDA.n2750 GNDA.n2743 9.3005
R3984 GNDA.n2752 GNDA.n2751 9.3005
R3985 GNDA.n2753 GNDA.n2742 9.3005
R3986 GNDA.n2755 GNDA.n2754 9.3005
R3987 GNDA.n2756 GNDA.n2741 9.3005
R3988 GNDA.n2758 GNDA.n2757 9.3005
R3989 GNDA.n2479 GNDA.n2478 9.3005
R3990 GNDA.n2480 GNDA.n112 9.3005
R3991 GNDA.n237 GNDA.n111 9.3005
R3992 GNDA.n240 GNDA.n238 9.3005
R3993 GNDA.n242 GNDA.n241 9.3005
R3994 GNDA.n243 GNDA.n236 9.3005
R3995 GNDA.n245 GNDA.n244 9.3005
R3996 GNDA.n246 GNDA.n235 9.3005
R3997 GNDA.n234 GNDA.n232 9.3005
R3998 GNDA.n233 GNDA.n221 9.3005
R3999 GNDA.n255 GNDA.n220 9.3005
R4000 GNDA.n288 GNDA.n199 9.3005
R4001 GNDA.n287 GNDA.n286 9.3005
R4002 GNDA.n285 GNDA.n200 9.3005
R4003 GNDA.n284 GNDA.n283 9.3005
R4004 GNDA.n282 GNDA.n201 9.3005
R4005 GNDA.n280 GNDA.n279 9.3005
R4006 GNDA.n278 GNDA.n202 9.3005
R4007 GNDA.n277 GNDA.n276 9.3005
R4008 GNDA.n204 GNDA.n203 9.3005
R4009 GNDA.n214 GNDA.n213 9.3005
R4010 GNDA.n267 GNDA.n215 9.3005
R4011 GNDA.n266 GNDA.n265 9.3005
R4012 GNDA.n264 GNDA.n216 9.3005
R4013 GNDA.n263 GNDA.n262 9.3005
R4014 GNDA.n261 GNDA.n217 9.3005
R4015 GNDA.n260 GNDA.n259 9.3005
R4016 GNDA.n258 GNDA.n219 9.3005
R4017 GNDA.n257 GNDA.n256 9.3005
R4018 GNDA.n2497 GNDA.n2496 9.3005
R4019 GNDA.n2498 GNDA.n104 9.3005
R4020 GNDA.n2500 GNDA.n2499 9.3005
R4021 GNDA.n2501 GNDA.n103 9.3005
R4022 GNDA.n2503 GNDA.n2502 9.3005
R4023 GNDA.n2504 GNDA.n102 9.3005
R4024 GNDA.n2506 GNDA.n2505 9.3005
R4025 GNDA.n2507 GNDA.n100 9.3005
R4026 GNDA.n2509 GNDA.n2508 9.3005
R4027 GNDA.n2510 GNDA.n99 9.3005
R4028 GNDA.n2513 GNDA.n2512 9.3005
R4029 GNDA.n2514 GNDA.n98 9.3005
R4030 GNDA.n2516 GNDA.n2515 9.3005
R4031 GNDA.n2517 GNDA.n96 9.3005
R4032 GNDA.n2522 GNDA.n2521 9.3005
R4033 GNDA.n2520 GNDA.n97 9.3005
R4034 GNDA.n2519 GNDA.n2518 9.3005
R4035 GNDA.n22 GNDA.n21 9.3005
R4036 GNDA.n2776 GNDA.n2775 9.3005
R4037 GNDA.n2777 GNDA.n20 9.3005
R4038 GNDA.n2779 GNDA.n2778 9.3005
R4039 GNDA.n2780 GNDA.n18 9.3005
R4040 GNDA.n2783 GNDA.n2782 9.3005
R4041 GNDA.n2784 GNDA.n17 9.3005
R4042 GNDA.n2786 GNDA.n2785 9.3005
R4043 GNDA.n2788 GNDA.n15 9.3005
R4044 GNDA.n2790 GNDA.n2789 9.3005
R4045 GNDA.n2791 GNDA.n14 9.3005
R4046 GNDA.n2793 GNDA.n2792 9.3005
R4047 GNDA.n2795 GNDA.n12 9.3005
R4048 GNDA.n2797 GNDA.n2796 9.3005
R4049 GNDA.n2798 GNDA.n11 9.3005
R4050 GNDA.n2800 GNDA.n2799 9.3005
R4051 GNDA.n2801 GNDA.n10 9.3005
R4052 GNDA.n2803 GNDA.n2802 9.3005
R4053 GNDA.n2804 GNDA.n9 9.3005
R4054 GNDA.n2806 GNDA.n2805 9.3005
R4055 GNDA.n2808 GNDA.n6 9.3005
R4056 GNDA.n2811 GNDA.n2810 9.3005
R4057 GNDA.n2812 GNDA.n5 9.3005
R4058 GNDA.n2814 GNDA.n2813 9.3005
R4059 GNDA.n2815 GNDA.n4 9.3005
R4060 GNDA.n2817 GNDA.n2816 9.3005
R4061 GNDA.n2818 GNDA.n3 9.3005
R4062 GNDA.n2820 GNDA.n2819 9.3005
R4063 GNDA.n2821 GNDA.n1 9.3005
R4064 GNDA.t221 GNDA.t161 8.67615
R4065 GNDA.n2116 GNDA.n374 8.60107
R4066 GNDA.n2367 GNDA.n375 8.60107
R4067 GNDA.t296 GNDA.t129 8.4512
R4068 GNDA.t232 GNDA.t250 8.4512
R4069 GNDA.n1810 GNDA.n1809 7.83472
R4070 GNDA.n2474 GNDA.n328 7.49888
R4071 GNDA.n298 GNDA.n297 7.11161
R4072 GNDA.n295 GNDA.n293 7.11161
R4073 GNDA.n2487 GNDA.n2486 7.11161
R4074 GNDA.n2484 GNDA.n2482 7.11161
R4075 GNDA.n912 GNDA.n867 6.72373
R4076 GNDA.n1897 GNDA.n1822 6.72373
R4077 GNDA.n2394 GNDA.n2393 6.72373
R4078 GNDA.n1968 GNDA.n1074 6.72373
R4079 GNDA.n1444 GNDA.n1178 6.72373
R4080 GNDA.n1421 GNDA.n1186 6.72373
R4081 GNDA.n291 GNDA.n290 6.69883
R4082 GNDA.n283 GNDA.n282 6.4005
R4083 GNDA.n261 GNDA.n260 6.4005
R4084 GNDA.n256 GNDA.n255 6.4005
R4085 GNDA.n311 GNDA.n310 6.4005
R4086 GNDA.n2523 GNDA.n2522 6.4005
R4087 GNDA.n2775 GNDA.n2774 6.4005
R4088 GNDA.n2788 GNDA.n2787 6.4005
R4089 GNDA.n2795 GNDA.n2794 6.4005
R4090 GNDA.n2807 GNDA.n2806 6.4005
R4091 GNDA.n2822 GNDA.n2821 6.4005
R4092 GNDA.n2461 GNDA.n334 6.4005
R4093 GNDA.n2442 GNDA.n2441 6.4005
R4094 GNDA.n2436 GNDA.n2435 6.4005
R4095 GNDA.n2424 GNDA.n2423 6.4005
R4096 GNDA.n2421 GNDA.n2420 6.4005
R4097 GNDA.n2409 GNDA.n2408 6.4005
R4098 GNDA.n2701 GNDA.n45 6.4005
R4099 GNDA.n2679 GNDA.n56 6.4005
R4100 GNDA.n2657 GNDA.n67 6.4005
R4101 GNDA.n2637 GNDA.n2636 6.4005
R4102 GNDA.n2591 GNDA.n2590 6.4005
R4103 GNDA.n2577 GNDA.n2538 6.4005
R4104 GNDA.n2566 GNDA.n2565 6.4005
R4105 GNDA.n2560 GNDA.n2559 6.4005
R4106 GNDA.n2480 GNDA.n2479 6.4005
R4107 GNDA.n1810 GNDA.n1099 6.36941
R4108 GNDA.n1447 GNDA.n1178 6.20656
R4109 GNDA.n912 GNDA.n846 6.20656
R4110 GNDA.n2393 GNDA.n404 6.20656
R4111 GNDA.n1969 GNDA.n1968 6.20656
R4112 GNDA.n1903 GNDA.n1822 6.20656
R4113 GNDA.n1422 GNDA.n1421 6.20656
R4114 GNDA.n1095 GNDA.t60 6.10596
R4115 GNDA.n1914 GNDA.n1913 6.07727
R4116 GNDA.n1807 GNDA.n1794 5.81868
R4117 GNDA.n1803 GNDA.n1794 5.81868
R4118 GNDA.n2767 GNDA.n8 5.68939
R4119 GNDA.n2404 GNDA.n352 5.68939
R4120 GNDA.n2404 GNDA.n353 5.68939
R4121 GNDA.n1811 GNDA.n1810 5.64455
R4122 GNDA.n1914 GNDA.n1078 5.5601
R4123 GNDA.n1688 GNDA.n1142 5.51161
R4124 GNDA.n1498 GNDA.n1496 5.51161
R4125 GNDA.n505 GNDA.n483 5.51161
R4126 GNDA.n798 GNDA.n693 5.51161
R4127 GNDA.n1031 GNDA.n918 5.51161
R4128 GNDA.n2149 GNDA.n2120 5.51161
R4129 GNDA.n2290 GNDA.n2268 5.51161
R4130 GNDA.n1388 GNDA.n1386 5.51161
R4131 GNDA.n2050 GNDA.n2020 5.51161
R4132 GNDA.n1599 GNDA.n1464 5.1717
R4133 GNDA.n804 GNDA.n799 5.1717
R4134 GNDA.n2019 GNDA.n1055 5.1717
R4135 GNDA.n2767 GNDA.n7 4.97828
R4136 GNDA.n2214 GNDA.n641 4.9157
R4137 GNDA.n2354 GNDA.n2240 4.9157
R4138 GNDA.n1347 GNDA.n1344 4.9157
R4139 GNDA.n1809 GNDA.n1808 4.69175
R4140 GNDA.n1102 GNDA.n1101 4.5005
R4141 GNDA.n1766 GNDA.n1104 4.5005
R4142 GNDA.n1768 GNDA.n1767 4.5005
R4143 GNDA.n1767 GNDA.n1766 4.5005
R4144 GNDA.n1676 GNDA.n1106 4.5005
R4145 GNDA.n1765 GNDA.n1764 4.5005
R4146 GNDA.n1817 GNDA.n1816 4.5005
R4147 GNDA.n183 GNDA.n181 4.49344
R4148 GNDA.n181 GNDA.n32 4.49344
R4149 GNDA.n189 GNDA.n188 4.49344
R4150 GNDA.n190 GNDA.n189 4.49344
R4151 GNDA.n1557 GNDA.t17 4.33832
R4152 GNDA.n1580 GNDA.t81 4.33832
R4153 GNDA.t201 GNDA.n1578 4.33832
R4154 GNDA.n1591 GNDA.t89 4.33832
R4155 GNDA.n1967 GNDA.n1966 4.26717
R4156 GNDA.n1966 GNDA.n1931 4.26717
R4157 GNDA.n1960 GNDA.n1931 4.26717
R4158 GNDA.n1960 GNDA.n1959 4.26717
R4159 GNDA.n1959 GNDA.n1958 4.26717
R4160 GNDA.n1958 GNDA.n1940 4.26717
R4161 GNDA.n1942 GNDA.n1940 4.26717
R4162 GNDA.n1949 GNDA.n1942 4.26717
R4163 GNDA.n1950 GNDA.n1949 4.26717
R4164 GNDA.n1950 GNDA.n916 4.26717
R4165 GNDA.n2113 GNDA.n916 4.26717
R4166 GNDA.n911 GNDA.n870 4.26717
R4167 GNDA.n906 GNDA.n870 4.26717
R4168 GNDA.n906 GNDA.n905 4.26717
R4169 GNDA.n905 GNDA.n904 4.26717
R4170 GNDA.n904 GNDA.n879 4.26717
R4171 GNDA.n898 GNDA.n879 4.26717
R4172 GNDA.n898 GNDA.n897 4.26717
R4173 GNDA.n897 GNDA.n896 4.26717
R4174 GNDA.n896 GNDA.n891 4.26717
R4175 GNDA.n891 GNDA.n440 4.26717
R4176 GNDA.n2364 GNDA.n440 4.26717
R4177 GNDA.n1643 GNDA.n1642 4.26717
R4178 GNDA.n1646 GNDA.n1643 4.26717
R4179 GNDA.n1646 GNDA.n1174 4.26717
R4180 GNDA.n1652 GNDA.n1174 4.26717
R4181 GNDA.n1653 GNDA.n1652 4.26717
R4182 GNDA.n1656 GNDA.n1653 4.26717
R4183 GNDA.n1656 GNDA.n1172 4.26717
R4184 GNDA.n1172 GNDA.n1168 4.26717
R4185 GNDA.n1663 GNDA.n1168 4.26717
R4186 GNDA.n1663 GNDA.n1169 4.26717
R4187 GNDA.n1169 GNDA.n1148 4.26717
R4188 GNDA.n1420 GNDA.n1419 4.26717
R4189 GNDA.n1419 GNDA.n1190 4.26717
R4190 GNDA.n1413 GNDA.n1190 4.26717
R4191 GNDA.n1413 GNDA.n1412 4.26717
R4192 GNDA.n1412 GNDA.n1411 4.26717
R4193 GNDA.n1411 GNDA.n1408 4.26717
R4194 GNDA.n1408 GNDA.n1407 4.26717
R4195 GNDA.n1407 GNDA.n1404 4.26717
R4196 GNDA.n1404 GNDA.n1403 4.26717
R4197 GNDA.n1403 GNDA.n1400 4.26717
R4198 GNDA.n1400 GNDA.n1399 4.26717
R4199 GNDA.n2392 GNDA.n406 4.26717
R4200 GNDA.n2386 GNDA.n406 4.26717
R4201 GNDA.n2386 GNDA.n2385 4.26717
R4202 GNDA.n2385 GNDA.n2384 4.26717
R4203 GNDA.n2384 GNDA.n2382 4.26717
R4204 GNDA.n2382 GNDA.n2379 4.26717
R4205 GNDA.n2379 GNDA.n2378 4.26717
R4206 GNDA.n2378 GNDA.n2375 4.26717
R4207 GNDA.n2375 GNDA.n2374 4.26717
R4208 GNDA.n2374 GNDA.n2371 4.26717
R4209 GNDA.n2371 GNDA.n2370 4.26717
R4210 GNDA.n1867 GNDA.n1866 4.26717
R4211 GNDA.n1866 GNDA.n1828 4.26717
R4212 GNDA.n1860 GNDA.n1828 4.26717
R4213 GNDA.n1860 GNDA.n1859 4.26717
R4214 GNDA.n1859 GNDA.n1858 4.26717
R4215 GNDA.n1858 GNDA.n1836 4.26717
R4216 GNDA.n1838 GNDA.n1836 4.26717
R4217 GNDA.n1845 GNDA.n1838 4.26717
R4218 GNDA.n1850 GNDA.n1845 4.26717
R4219 GNDA.n1850 GNDA.n1849 4.26717
R4220 GNDA.n1849 GNDA.n1848 4.26717
R4221 GNDA.n1968 GNDA.n1967 3.93531
R4222 GNDA.n912 GNDA.n911 3.93531
R4223 GNDA.n1642 GNDA.n1178 3.93531
R4224 GNDA.n1421 GNDA.n1420 3.93531
R4225 GNDA.n2393 GNDA.n2392 3.93531
R4226 GNDA.n1867 GNDA.n1822 3.93531
R4227 GNDA.n182 GNDA.n180 3.8278
R4228 GNDA.n187 GNDA.n186 3.8278
R4229 GNDA.n26 GNDA.n25 3.8278
R4230 GNDA.n1583 GNDA.n1492 3.7893
R4231 GNDA.n1582 GNDA.n1493 3.7893
R4232 GNDA.n1564 GNDA.n1563 3.7893
R4233 GNDA.n1576 GNDA.n1575 3.7893
R4234 GNDA.n1572 GNDA.n1571 3.7893
R4235 GNDA.n1567 GNDA.n1469 3.7893
R4236 GNDA.n1589 GNDA.n1588 3.7893
R4237 GNDA.n1472 GNDA.n1470 3.7893
R4238 GNDA.n1756 GNDA.n1755 3.7893
R4239 GNDA.n1752 GNDA.n1117 3.7893
R4240 GNDA.n1751 GNDA.n1120 3.7893
R4241 GNDA.n1124 GNDA.n1123 3.7893
R4242 GNDA.n1745 GNDA.n1744 3.7893
R4243 GNDA.n1159 GNDA.n1158 3.7893
R4244 GNDA.n1155 GNDA.n1154 3.7893
R4245 GNDA.n1685 GNDA.n1143 3.7893
R4246 GNDA.n568 GNDA.n567 3.7893
R4247 GNDA.n564 GNDA.n460 3.7893
R4248 GNDA.n563 GNDA.n463 3.7893
R4249 GNDA.n560 GNDA.n559 3.7893
R4250 GNDA.n485 GNDA.n464 3.7893
R4251 GNDA.n494 GNDA.n493 3.7893
R4252 GNDA.n497 GNDA.n484 3.7893
R4253 GNDA.n502 GNDA.n498 3.7893
R4254 GNDA.n2360 GNDA.n444 3.7893
R4255 GNDA.n787 GNDA.n766 3.7893
R4256 GNDA.n786 GNDA.n767 3.7893
R4257 GNDA.n783 GNDA.n782 3.7893
R4258 GNDA.n779 GNDA.n768 3.7893
R4259 GNDA.n772 GNDA.n769 3.7893
R4260 GNDA.n793 GNDA.n695 3.7893
R4261 GNDA.n794 GNDA.n694 3.7893
R4262 GNDA.n1021 GNDA.n996 3.7893
R4263 GNDA.n1020 GNDA.n1017 3.7893
R4264 GNDA.n1016 GNDA.n997 3.7893
R4265 GNDA.n1013 GNDA.n1012 3.7893
R4266 GNDA.n1009 GNDA.n998 3.7893
R4267 GNDA.n1002 GNDA.n999 3.7893
R4268 GNDA.n1026 GNDA.n920 3.7893
R4269 GNDA.n1027 GNDA.n919 3.7893
R4270 GNDA.n2199 GNDA.n660 3.7893
R4271 GNDA.n2207 GNDA.n2206 3.7893
R4272 GNDA.n2122 GNDA.n661 3.7893
R4273 GNDA.n2126 GNDA.n2124 3.7893
R4274 GNDA.n2131 GNDA.n2127 3.7893
R4275 GNDA.n2138 GNDA.n2137 3.7893
R4276 GNDA.n2141 GNDA.n2121 3.7893
R4277 GNDA.n2146 GNDA.n2142 3.7893
R4278 GNDA.n2352 GNDA.n2351 3.7893
R4279 GNDA.n2348 GNDA.n2243 3.7893
R4280 GNDA.n2347 GNDA.n2246 3.7893
R4281 GNDA.n2344 GNDA.n2343 3.7893
R4282 GNDA.n2270 GNDA.n2247 3.7893
R4283 GNDA.n2279 GNDA.n2278 3.7893
R4284 GNDA.n2282 GNDA.n2269 3.7893
R4285 GNDA.n2287 GNDA.n2283 3.7893
R4286 GNDA.n1348 GNDA.n1230 3.7893
R4287 GNDA.n1357 GNDA.n1356 3.7893
R4288 GNDA.n1231 GNDA.n1226 3.7893
R4289 GNDA.n1365 GNDA.n1363 3.7893
R4290 GNDA.n1364 GNDA.n1224 3.7893
R4291 GNDA.n1223 GNDA.n1220 3.7893
R4292 GNDA.n1381 GNDA.n1379 3.7893
R4293 GNDA.n1380 GNDA.n1216 3.7893
R4294 GNDA.n2109 GNDA.n1035 3.7893
R4295 GNDA.n2106 GNDA.n2105 3.7893
R4296 GNDA.n2022 GNDA.n1036 3.7893
R4297 GNDA.n2027 GNDA.n2025 3.7893
R4298 GNDA.n2032 GNDA.n2028 3.7893
R4299 GNDA.n2039 GNDA.n2038 3.7893
R4300 GNDA.n2042 GNDA.n2021 3.7893
R4301 GNDA.n2047 GNDA.n2043 3.7893
R4302 GNDA.n1568 GNDA 3.7381
R4303 GNDA.n1153 GNDA 3.7381
R4304 GNDA.n490 GNDA 3.7381
R4305 GNDA GNDA.n775 3.7381
R4306 GNDA GNDA.n1005 3.7381
R4307 GNDA.n2134 GNDA 3.7381
R4308 GNDA.n2275 GNDA 3.7381
R4309 GNDA GNDA.n1371 3.7381
R4310 GNDA.n2035 GNDA 3.7381
R4311 GNDA.n297 GNDA.n296 3.48951
R4312 GNDA.n296 GNDA.n295 3.48951
R4313 GNDA.n2486 GNDA.n2485 3.48951
R4314 GNDA.n2485 GNDA.n2484 3.48951
R4315 GNDA.n2467 GNDA.n330 3.2005
R4316 GNDA.n2455 GNDA.n2454 3.2005
R4317 GNDA.n2694 GNDA.n50 3.2005
R4318 GNDA.n2672 GNDA.n61 3.2005
R4319 GNDA.n2650 GNDA.n2649 3.2005
R4320 GNDA.n2617 GNDA.n2616 3.2005
R4321 GNDA.n2605 GNDA.n93 3.2005
R4322 GNDA.t208 GNDA.n379 2.96739
R4323 GNDA.n2760 GNDA.n27 2.8779
R4324 GNDA.n2761 GNDA.n2760 2.8779
R4325 GNDA.n1785 GNDA.n1773 2.86505
R4326 GNDA.n1785 GNDA.n1784 2.86505
R4327 GNDA.n1782 GNDA.n1776 2.86505
R4328 GNDA.n1777 GNDA.n1776 2.86505
R4329 GNDA.n1784 GNDA.n1783 2.86505
R4330 GNDA.n1780 GNDA.n1777 2.86505
R4331 GNDA.n1788 GNDA.n1773 2.86505
R4332 GNDA.n1783 GNDA.n1782 2.86505
R4333 GNDA.n1802 GNDA.n1801 2.86505
R4334 GNDA.n1801 GNDA.n1800 2.86505
R4335 GNDA.n1800 GNDA.n1799 2.86505
R4336 GNDA.n1803 GNDA.n1802 2.86505
R4337 GNDA.t158 GNDA.t258 2.82463
R4338 GNDA.t213 GNDA.t84 2.8174
R4339 GNDA.n1551 GNDA.n1550 2.6629
R4340 GNDA.n1212 GNDA.n1116 2.6629
R4341 GNDA.n1495 GNDA.n1494 2.6629
R4342 GNDA.n459 GNDA.n458 2.6629
R4343 GNDA.n2363 GNDA.n442 2.6629
R4344 GNDA.n2362 GNDA.n2361 2.6629
R4345 GNDA.n995 GNDA.n994 2.6629
R4346 GNDA.n2112 GNDA.n1033 2.6629
R4347 GNDA.n2200 GNDA.n641 2.6629
R4348 GNDA.n2119 GNDA.n681 2.6629
R4349 GNDA.n2354 GNDA.n2353 2.6629
R4350 GNDA.n2267 GNDA.n432 2.6629
R4351 GNDA.n1349 GNDA.n1347 2.6629
R4352 GNDA.n1387 GNDA.n1213 2.6629
R4353 GNDA.n2111 GNDA.n2110 2.6629
R4354 GNDA.t181 GNDA.n2398 2.54362
R4355 GNDA.n1551 GNDA.n1495 2.4581
R4356 GNDA.n1496 GNDA.n1464 2.4581
R4357 GNDA.n1213 GNDA.n1212 2.4581
R4358 GNDA.n1494 GNDA.n1142 2.4581
R4359 GNDA.n458 GNDA.n432 2.4581
R4360 GNDA.n483 GNDA.n442 2.4581
R4361 GNDA.n2363 GNDA.n2362 2.4581
R4362 GNDA.n799 GNDA.n798 2.4581
R4363 GNDA.n994 GNDA.n681 2.4581
R4364 GNDA.n1033 GNDA.n1031 2.4581
R4365 GNDA.n2120 GNDA.n2119 2.4581
R4366 GNDA.n2268 GNDA.n2267 2.4581
R4367 GNDA.n1388 GNDA.n1387 2.4581
R4368 GNDA.n2112 GNDA.n2111 2.4581
R4369 GNDA.n2020 GNDA.n2019 2.4581
R4370 GNDA.n1099 GNDA.n1085 2.44675
R4371 GNDA.n1099 GNDA.n1098 2.44675
R4372 GNDA.n1791 GNDA.n1790 2.26187
R4373 GNDA.n249 GNDA.n231 2.25882
R4374 GNDA.n231 GNDA.n230 2.25882
R4375 GNDA.n254 GNDA.n222 2.25882
R4376 GNDA.n230 GNDA.n229 2.25882
R4377 GNDA.n250 GNDA.n249 2.25882
R4378 GNDA.n229 GNDA.n222 2.25882
R4379 GNDA.n270 GNDA.n212 2.25882
R4380 GNDA.n212 GNDA.n211 2.25882
R4381 GNDA.n275 GNDA.n205 2.25882
R4382 GNDA.n211 GNDA.n210 2.25882
R4383 GNDA.n271 GNDA.n270 2.25882
R4384 GNDA.n210 GNDA.n205 2.25882
R4385 GNDA.n1792 GNDA.n1100 2.24063
R4386 GNDA.n1772 GNDA.n1771 2.24063
R4387 GNDA.n1769 GNDA.n1768 2.24063
R4388 GNDA.n1107 GNDA.n1105 2.24063
R4389 GNDA.n1790 GNDA.n1789 2.24063
R4390 GNDA.n1770 GNDA.n1103 2.24063
R4391 GNDA.n1674 GNDA.n1106 2.22018
R4392 GNDA.n1765 GNDA.n1108 2.22018
R4393 GNDA.n1816 GNDA.n1814 2.22018
R4394 GNDA.n2113 GNDA.n2112 2.18124
R4395 GNDA.n2364 GNDA.n2363 2.18124
R4396 GNDA.n1495 GNDA.n1148 2.18124
R4397 GNDA.n1399 GNDA.n1213 2.18124
R4398 GNDA.n2370 GNDA.n432 2.18124
R4399 GNDA.n1848 GNDA.n681 2.18124
R4400 GNDA.n1496 GNDA.n1466 2.1509
R4401 GNDA.n1684 GNDA.n1142 2.1509
R4402 GNDA.n501 GNDA.n483 2.1509
R4403 GNDA.n798 GNDA.n797 2.1509
R4404 GNDA.n1031 GNDA.n1030 2.1509
R4405 GNDA.n2145 GNDA.n2120 2.1509
R4406 GNDA.n2286 GNDA.n2268 2.1509
R4407 GNDA.n1389 GNDA.n1388 2.1509
R4408 GNDA.n2046 GNDA.n2020 2.1509
R4409 GNDA.n1724 GNDA.n1116 2.13383
R4410 GNDA.n1550 GNDA.n1549 2.13383
R4411 GNDA.n541 GNDA.n459 2.13383
R4412 GNDA.n2361 GNDA.n443 2.13383
R4413 GNDA.n995 GNDA.n992 2.13383
R4414 GNDA.n2201 GNDA.n2200 2.13383
R4415 GNDA.n2353 GNDA.n2241 2.13383
R4416 GNDA.n1350 GNDA.n1349 2.13383
R4417 GNDA.n2110 GNDA.n1034 2.13383
R4418 GNDA.n2112 GNDA.n913 2.08643
R4419 GNDA.n2363 GNDA.n437 2.08643
R4420 GNDA.n1495 GNDA.n1147 2.08643
R4421 GNDA.n1395 GNDA.n1213 2.08643
R4422 GNDA.n434 GNDA.n432 2.08643
R4423 GNDA.n681 GNDA.n405 2.08643
R4424 GNDA.n1550 GNDA.n1492 1.9461
R4425 GNDA.n1756 GNDA.n1116 1.9461
R4426 GNDA.n568 GNDA.n459 1.9461
R4427 GNDA.n2361 GNDA.n2360 1.9461
R4428 GNDA.n996 GNDA.n995 1.9461
R4429 GNDA.n2200 GNDA.n2199 1.9461
R4430 GNDA.n2353 GNDA.n2352 1.9461
R4431 GNDA.n1349 GNDA.n1348 1.9461
R4432 GNDA.n2110 GNDA.n2109 1.9461
R4433 GNDA.n2475 GNDA.n327 1.5139
R4434 GNDA.n1600 GNDA.n1599 1.47392
R4435 GNDA.n805 GNDA.n804 1.47392
R4436 GNDA.n2217 GNDA.n2214 1.47392
R4437 GNDA.n2240 GNDA.n578 1.47392
R4438 GNDA.n1344 GNDA.n1342 1.47392
R4439 GNDA.n2013 GNDA.n1055 1.47392
R4440 GNDA.n1816 GNDA.n1815 1.20883
R4441 GNDA.n1816 GNDA.n1812 1.14633
R4442 GNDA.n2237 GNDA.n379 1.12708
R4443 GNDA.n2398 GNDA.n362 0.978912
R4444 GNDA.n2476 GNDA.n2475 0.9781
R4445 GNDA.n1583 GNDA.n1582 0.8197
R4446 GNDA.n1563 GNDA.n1493 0.8197
R4447 GNDA.n1576 GNDA.n1564 0.8197
R4448 GNDA.n1575 GNDA.n1572 0.8197
R4449 GNDA.n1568 GNDA.n1567 0.8197
R4450 GNDA.n1589 GNDA.n1469 0.8197
R4451 GNDA.n1588 GNDA.n1470 0.8197
R4452 GNDA.n1472 GNDA.n1466 0.8197
R4453 GNDA.n1755 GNDA.n1117 0.8197
R4454 GNDA.n1752 GNDA.n1751 0.8197
R4455 GNDA.n1123 GNDA.n1120 0.8197
R4456 GNDA.n1745 GNDA.n1124 0.8197
R4457 GNDA.n1159 GNDA.n1153 0.8197
R4458 GNDA.n1158 GNDA.n1154 0.8197
R4459 GNDA.n1155 GNDA.n1143 0.8197
R4460 GNDA.n1685 GNDA.n1684 0.8197
R4461 GNDA.n567 GNDA.n460 0.8197
R4462 GNDA.n564 GNDA.n563 0.8197
R4463 GNDA.n560 GNDA.n463 0.8197
R4464 GNDA.n559 GNDA.n464 0.8197
R4465 GNDA.n493 GNDA.n490 0.8197
R4466 GNDA.n494 GNDA.n484 0.8197
R4467 GNDA.n498 GNDA.n497 0.8197
R4468 GNDA.n502 GNDA.n501 0.8197
R4469 GNDA.n766 GNDA.n444 0.8197
R4470 GNDA.n787 GNDA.n786 0.8197
R4471 GNDA.n783 GNDA.n767 0.8197
R4472 GNDA.n782 GNDA.n779 0.8197
R4473 GNDA.n775 GNDA.n772 0.8197
R4474 GNDA.n769 GNDA.n695 0.8197
R4475 GNDA.n794 GNDA.n793 0.8197
R4476 GNDA.n797 GNDA.n694 0.8197
R4477 GNDA.n1021 GNDA.n1020 0.8197
R4478 GNDA.n1017 GNDA.n1016 0.8197
R4479 GNDA.n1013 GNDA.n997 0.8197
R4480 GNDA.n1012 GNDA.n1009 0.8197
R4481 GNDA.n1005 GNDA.n1002 0.8197
R4482 GNDA.n999 GNDA.n920 0.8197
R4483 GNDA.n1027 GNDA.n1026 0.8197
R4484 GNDA.n1030 GNDA.n919 0.8197
R4485 GNDA.n2207 GNDA.n660 0.8197
R4486 GNDA.n2206 GNDA.n661 0.8197
R4487 GNDA.n2124 GNDA.n2122 0.8197
R4488 GNDA.n2127 GNDA.n2126 0.8197
R4489 GNDA.n2137 GNDA.n2134 0.8197
R4490 GNDA.n2138 GNDA.n2121 0.8197
R4491 GNDA.n2142 GNDA.n2141 0.8197
R4492 GNDA.n2146 GNDA.n2145 0.8197
R4493 GNDA.n2351 GNDA.n2243 0.8197
R4494 GNDA.n2348 GNDA.n2347 0.8197
R4495 GNDA.n2344 GNDA.n2246 0.8197
R4496 GNDA.n2343 GNDA.n2247 0.8197
R4497 GNDA.n2278 GNDA.n2275 0.8197
R4498 GNDA.n2279 GNDA.n2269 0.8197
R4499 GNDA.n2283 GNDA.n2282 0.8197
R4500 GNDA.n2287 GNDA.n2286 0.8197
R4501 GNDA.n1357 GNDA.n1230 0.8197
R4502 GNDA.n1356 GNDA.n1231 0.8197
R4503 GNDA.n1363 GNDA.n1226 0.8197
R4504 GNDA.n1365 GNDA.n1364 0.8197
R4505 GNDA.n1371 GNDA.n1223 0.8197
R4506 GNDA.n1379 GNDA.n1220 0.8197
R4507 GNDA.n1381 GNDA.n1380 0.8197
R4508 GNDA.n1389 GNDA.n1216 0.8197
R4509 GNDA.n2106 GNDA.n1035 0.8197
R4510 GNDA.n2105 GNDA.n1036 0.8197
R4511 GNDA.n2025 GNDA.n2022 0.8197
R4512 GNDA.n2028 GNDA.n2027 0.8197
R4513 GNDA.n2038 GNDA.n2035 0.8197
R4514 GNDA.n2039 GNDA.n2021 0.8197
R4515 GNDA.n2043 GNDA.n2042 0.8197
R4516 GNDA.n2047 GNDA.n2046 0.8197
R4517 GNDA.n1809 GNDA.n327 0.79984
R4518 GNDA.n291 GNDA.n199 0.703977
R4519 GNDA.n1808 GNDA.n1792 0.65675
R4520 GNDA.n1571 GNDA 0.5637
R4521 GNDA.n1744 GNDA 0.5637
R4522 GNDA GNDA.n485 0.5637
R4523 GNDA GNDA.n768 0.5637
R4524 GNDA GNDA.n998 0.5637
R4525 GNDA.n2131 GNDA 0.5637
R4526 GNDA GNDA.n2270 0.5637
R4527 GNDA.n1224 GNDA 0.5637
R4528 GNDA.n2032 GNDA 0.5637
R4529 GNDA.n1771 GNDA.n1770 0.542167
R4530 GNDA.n2551 GNDA.n2548 0.442364
R4531 GNDA.n1566 GNDA 0.2565
R4532 GNDA.n1152 GNDA 0.2565
R4533 GNDA.n488 GNDA 0.2565
R4534 GNDA.n776 GNDA 0.2565
R4535 GNDA.n1006 GNDA 0.2565
R4536 GNDA GNDA.n2130 0.2565
R4537 GNDA.n2273 GNDA 0.2565
R4538 GNDA.n1372 GNDA 0.2565
R4539 GNDA GNDA.n2031 0.2565
R4540 GNDA.n2474 GNDA.n2473 0.193977
R4541 GNDA.n357 GNDA.n0 0.193881
R4542 GNDA.n2823 GNDA.n1 0.193881
R4543 GNDA.n2497 GNDA.n105 0.193695
R4544 GNDA.n2715 GNDA.n2714 0.193477
R4545 GNDA.n326 GNDA.n113 0.188
R4546 GNDA.n1766 GNDA.n1765 0.188
R4547 GNDA.n1768 GNDA.n1106 0.188
R4548 GNDA.n1812 GNDA.n1811 0.188
R4549 GNDA.n2746 GNDA 0.162727
R4550 GNDA.n166 GNDA.n131 0.15675
R4551 GNDA.n162 GNDA.n161 0.15675
R4552 GNDA.n161 GNDA.n160 0.15675
R4553 GNDA.n160 GNDA.n135 0.15675
R4554 GNDA.n156 GNDA.n155 0.15675
R4555 GNDA.n155 GNDA.n154 0.15675
R4556 GNDA.n154 GNDA.n139 0.15675
R4557 GNDA.n150 GNDA.n149 0.15675
R4558 GNDA.n149 GNDA.n148 0.15675
R4559 GNDA.n148 GNDA.n145 0.15675
R4560 GNDA.n312 GNDA.n118 0.15675
R4561 GNDA.n313 GNDA.n312 0.15675
R4562 GNDA.n316 GNDA.n313 0.15675
R4563 GNDA.n320 GNDA.n116 0.15675
R4564 GNDA.n323 GNDA.n322 0.15675
R4565 GNDA.n323 GNDA.n113 0.15675
R4566 GNDA.n2473 GNDA.n329 0.15675
R4567 GNDA.n2469 GNDA.n329 0.15675
R4568 GNDA.n2469 GNDA.n2468 0.15675
R4569 GNDA.n2468 GNDA.n331 0.15675
R4570 GNDA.n2464 GNDA.n331 0.15675
R4571 GNDA.n2464 GNDA.n2463 0.15675
R4572 GNDA.n2463 GNDA.n2462 0.15675
R4573 GNDA.n2462 GNDA.n333 0.15675
R4574 GNDA.n2458 GNDA.n333 0.15675
R4575 GNDA.n2458 GNDA.n2457 0.15675
R4576 GNDA.n2457 GNDA.n2456 0.15675
R4577 GNDA.n2456 GNDA.n336 0.15675
R4578 GNDA.n341 GNDA.n336 0.15675
R4579 GNDA.n342 GNDA.n341 0.15675
R4580 GNDA.n2447 GNDA.n342 0.15675
R4581 GNDA.n2447 GNDA.n2446 0.15675
R4582 GNDA.n2446 GNDA.n2445 0.15675
R4583 GNDA.n2445 GNDA.n343 0.15675
R4584 GNDA.n2440 GNDA.n343 0.15675
R4585 GNDA.n2440 GNDA.n2439 0.15675
R4586 GNDA.n2439 GNDA.n2438 0.15675
R4587 GNDA.n2438 GNDA.n346 0.15675
R4588 GNDA.n2433 GNDA.n346 0.15675
R4589 GNDA.n2433 GNDA.n2432 0.15675
R4590 GNDA.n2432 GNDA.n2431 0.15675
R4591 GNDA.n2431 GNDA.n349 0.15675
R4592 GNDA.n2427 GNDA.n349 0.15675
R4593 GNDA.n2427 GNDA.n2426 0.15675
R4594 GNDA.n2426 GNDA.n2425 0.15675
R4595 GNDA.n2425 GNDA.n351 0.15675
R4596 GNDA.n2419 GNDA.n351 0.15675
R4597 GNDA.n2419 GNDA.n2418 0.15675
R4598 GNDA.n2418 GNDA.n2417 0.15675
R4599 GNDA.n2417 GNDA.n355 0.15675
R4600 GNDA.n2413 GNDA.n355 0.15675
R4601 GNDA.n2413 GNDA.n2412 0.15675
R4602 GNDA.n2412 GNDA.n2411 0.15675
R4603 GNDA.n2411 GNDA.n357 0.15675
R4604 GNDA.n2714 GNDA.n40 0.15675
R4605 GNDA.n2710 GNDA.n40 0.15675
R4606 GNDA.n2710 GNDA.n2709 0.15675
R4607 GNDA.n2709 GNDA.n2708 0.15675
R4608 GNDA.n2708 GNDA.n42 0.15675
R4609 GNDA.n2703 GNDA.n42 0.15675
R4610 GNDA.n2703 GNDA.n2702 0.15675
R4611 GNDA.n2702 GNDA.n46 0.15675
R4612 GNDA.n2698 GNDA.n46 0.15675
R4613 GNDA.n2698 GNDA.n2697 0.15675
R4614 GNDA.n2697 GNDA.n48 0.15675
R4615 GNDA.n2693 GNDA.n48 0.15675
R4616 GNDA.n2693 GNDA.n2692 0.15675
R4617 GNDA.n2692 GNDA.n51 0.15675
R4618 GNDA.n2688 GNDA.n51 0.15675
R4619 GNDA.n2688 GNDA.n2687 0.15675
R4620 GNDA.n2687 GNDA.n2686 0.15675
R4621 GNDA.n2686 GNDA.n53 0.15675
R4622 GNDA.n2681 GNDA.n53 0.15675
R4623 GNDA.n2681 GNDA.n2680 0.15675
R4624 GNDA.n2680 GNDA.n57 0.15675
R4625 GNDA.n2676 GNDA.n57 0.15675
R4626 GNDA.n2676 GNDA.n2675 0.15675
R4627 GNDA.n2675 GNDA.n59 0.15675
R4628 GNDA.n2671 GNDA.n59 0.15675
R4629 GNDA.n2671 GNDA.n2670 0.15675
R4630 GNDA.n2670 GNDA.n62 0.15675
R4631 GNDA.n2666 GNDA.n62 0.15675
R4632 GNDA.n2666 GNDA.n2665 0.15675
R4633 GNDA.n2665 GNDA.n2664 0.15675
R4634 GNDA.n2664 GNDA.n64 0.15675
R4635 GNDA.n2659 GNDA.n64 0.15675
R4636 GNDA.n2659 GNDA.n2658 0.15675
R4637 GNDA.n2658 GNDA.n68 0.15675
R4638 GNDA.n2654 GNDA.n68 0.15675
R4639 GNDA.n2654 GNDA.n2653 0.15675
R4640 GNDA.n2653 GNDA.n70 0.15675
R4641 GNDA.n2648 GNDA.n70 0.15675
R4642 GNDA.n2648 GNDA.n2647 0.15675
R4643 GNDA.n2647 GNDA.n2646 0.15675
R4644 GNDA.n2646 GNDA.n73 0.15675
R4645 GNDA.n2642 GNDA.n73 0.15675
R4646 GNDA.n2642 GNDA.n2641 0.15675
R4647 GNDA.n2641 GNDA.n2640 0.15675
R4648 GNDA.n2640 GNDA.n75 0.15675
R4649 GNDA.n2635 GNDA.n75 0.15675
R4650 GNDA.n2635 GNDA.n2634 0.15675
R4651 GNDA.n2634 GNDA.n2633 0.15675
R4652 GNDA.n2633 GNDA.n80 0.15675
R4653 GNDA.n2629 GNDA.n80 0.15675
R4654 GNDA.n2629 GNDA.n2628 0.15675
R4655 GNDA.n2628 GNDA.n2627 0.15675
R4656 GNDA.n2627 GNDA.n82 0.15675
R4657 GNDA.n2622 GNDA.n82 0.15675
R4658 GNDA.n2622 GNDA.n2621 0.15675
R4659 GNDA.n2621 GNDA.n2620 0.15675
R4660 GNDA.n2620 GNDA.n85 0.15675
R4661 GNDA.n2615 GNDA.n85 0.15675
R4662 GNDA.n2615 GNDA.n2614 0.15675
R4663 GNDA.n2614 GNDA.n2613 0.15675
R4664 GNDA.n2613 GNDA.n90 0.15675
R4665 GNDA.n2608 GNDA.n90 0.15675
R4666 GNDA.n2608 GNDA.n2607 0.15675
R4667 GNDA.n2607 GNDA.n2606 0.15675
R4668 GNDA.n2606 GNDA.n92 0.15675
R4669 GNDA.n2602 GNDA.n92 0.15675
R4670 GNDA.n2602 GNDA.n2601 0.15675
R4671 GNDA.n2601 GNDA.n2600 0.15675
R4672 GNDA.n2600 GNDA.n95 0.15675
R4673 GNDA.n2595 GNDA.n95 0.15675
R4674 GNDA.n2595 GNDA.n2594 0.15675
R4675 GNDA.n2594 GNDA.n2593 0.15675
R4676 GNDA.n2593 GNDA.n2529 0.15675
R4677 GNDA.n2588 GNDA.n2529 0.15675
R4678 GNDA.n2588 GNDA.n2587 0.15675
R4679 GNDA.n2587 GNDA.n2586 0.15675
R4680 GNDA.n2586 GNDA.n2532 0.15675
R4681 GNDA.n2582 GNDA.n2532 0.15675
R4682 GNDA.n2582 GNDA.n2581 0.15675
R4683 GNDA.n2581 GNDA.n2580 0.15675
R4684 GNDA.n2580 GNDA.n2536 0.15675
R4685 GNDA.n2576 GNDA.n2536 0.15675
R4686 GNDA.n2576 GNDA.n2575 0.15675
R4687 GNDA.n2575 GNDA.n2539 0.15675
R4688 GNDA.n2571 GNDA.n2539 0.15675
R4689 GNDA.n2571 GNDA.n2570 0.15675
R4690 GNDA.n2570 GNDA.n2569 0.15675
R4691 GNDA.n2569 GNDA.n2541 0.15675
R4692 GNDA.n2564 GNDA.n2541 0.15675
R4693 GNDA.n2564 GNDA.n2563 0.15675
R4694 GNDA.n2563 GNDA.n2562 0.15675
R4695 GNDA.n2562 GNDA.n2546 0.15675
R4696 GNDA.n2557 GNDA.n2546 0.15675
R4697 GNDA.n2557 GNDA.n2556 0.15675
R4698 GNDA.n2556 GNDA.n2555 0.15675
R4699 GNDA.n2555 GNDA.n2548 0.15675
R4700 GNDA.n2749 GNDA.n2744 0.15675
R4701 GNDA.n2750 GNDA.n2749 0.15675
R4702 GNDA.n2751 GNDA.n2750 0.15675
R4703 GNDA.n2751 GNDA.n2742 0.15675
R4704 GNDA.n2755 GNDA.n2742 0.15675
R4705 GNDA.n2756 GNDA.n2755 0.15675
R4706 GNDA.n2757 GNDA.n2756 0.15675
R4707 GNDA.n2757 GNDA.n2740 0.15675
R4708 GNDA.n2740 GNDA.n2739 0.15675
R4709 GNDA.n2739 GNDA.n2738 0.15675
R4710 GNDA.n2738 GNDA.n29 0.15675
R4711 GNDA.n2734 GNDA.n29 0.15675
R4712 GNDA.n2734 GNDA.n2733 0.15675
R4713 GNDA.n2733 GNDA.n2732 0.15675
R4714 GNDA.n2732 GNDA.n31 0.15675
R4715 GNDA.n2728 GNDA.n31 0.15675
R4716 GNDA.n2728 GNDA.n2727 0.15675
R4717 GNDA.n2727 GNDA.n2726 0.15675
R4718 GNDA.n2726 GNDA.n34 0.15675
R4719 GNDA.n2722 GNDA.n34 0.15675
R4720 GNDA.n2722 GNDA.n2721 0.15675
R4721 GNDA.n2721 GNDA.n2720 0.15675
R4722 GNDA.n2720 GNDA.n36 0.15675
R4723 GNDA.n286 GNDA.n199 0.15675
R4724 GNDA.n286 GNDA.n285 0.15675
R4725 GNDA.n285 GNDA.n284 0.15675
R4726 GNDA.n284 GNDA.n201 0.15675
R4727 GNDA.n279 GNDA.n201 0.15675
R4728 GNDA.n279 GNDA.n278 0.15675
R4729 GNDA.n278 GNDA.n277 0.15675
R4730 GNDA.n277 GNDA.n203 0.15675
R4731 GNDA.n214 GNDA.n203 0.15675
R4732 GNDA.n215 GNDA.n214 0.15675
R4733 GNDA.n265 GNDA.n215 0.15675
R4734 GNDA.n265 GNDA.n264 0.15675
R4735 GNDA.n264 GNDA.n263 0.15675
R4736 GNDA.n263 GNDA.n217 0.15675
R4737 GNDA.n259 GNDA.n217 0.15675
R4738 GNDA.n259 GNDA.n258 0.15675
R4739 GNDA.n258 GNDA.n257 0.15675
R4740 GNDA.n257 GNDA.n220 0.15675
R4741 GNDA.n233 GNDA.n220 0.15675
R4742 GNDA.n234 GNDA.n233 0.15675
R4743 GNDA.n235 GNDA.n234 0.15675
R4744 GNDA.n244 GNDA.n235 0.15675
R4745 GNDA.n244 GNDA.n243 0.15675
R4746 GNDA.n243 GNDA.n242 0.15675
R4747 GNDA.n242 GNDA.n238 0.15675
R4748 GNDA.n238 GNDA.n237 0.15675
R4749 GNDA.n237 GNDA.n112 0.15675
R4750 GNDA.n2478 GNDA.n112 0.15675
R4751 GNDA.n2498 GNDA.n2497 0.15675
R4752 GNDA.n2499 GNDA.n2498 0.15675
R4753 GNDA.n2499 GNDA.n103 0.15675
R4754 GNDA.n2503 GNDA.n103 0.15675
R4755 GNDA.n2504 GNDA.n2503 0.15675
R4756 GNDA.n2505 GNDA.n2504 0.15675
R4757 GNDA.n2505 GNDA.n100 0.15675
R4758 GNDA.n2509 GNDA.n100 0.15675
R4759 GNDA.n2510 GNDA.n2509 0.15675
R4760 GNDA.n2512 GNDA.n98 0.15675
R4761 GNDA.n2516 GNDA.n98 0.15675
R4762 GNDA.n2517 GNDA.n2516 0.15675
R4763 GNDA.n2521 GNDA.n2517 0.15675
R4764 GNDA.n2521 GNDA.n2520 0.15675
R4765 GNDA.n2520 GNDA.n2519 0.15675
R4766 GNDA.n2519 GNDA.n21 0.15675
R4767 GNDA.n2776 GNDA.n21 0.15675
R4768 GNDA.n2777 GNDA.n2776 0.15675
R4769 GNDA.n2778 GNDA.n2777 0.15675
R4770 GNDA.n2778 GNDA.n18 0.15675
R4771 GNDA.n2783 GNDA.n18 0.15675
R4772 GNDA.n2784 GNDA.n2783 0.15675
R4773 GNDA.n2785 GNDA.n2784 0.15675
R4774 GNDA.n2785 GNDA.n15 0.15675
R4775 GNDA.n2790 GNDA.n15 0.15675
R4776 GNDA.n2791 GNDA.n2790 0.15675
R4777 GNDA.n2792 GNDA.n2791 0.15675
R4778 GNDA.n2792 GNDA.n12 0.15675
R4779 GNDA.n2797 GNDA.n12 0.15675
R4780 GNDA.n2798 GNDA.n2797 0.15675
R4781 GNDA.n2799 GNDA.n2798 0.15675
R4782 GNDA.n2799 GNDA.n10 0.15675
R4783 GNDA.n2803 GNDA.n10 0.15675
R4784 GNDA.n2804 GNDA.n2803 0.15675
R4785 GNDA.n2805 GNDA.n2804 0.15675
R4786 GNDA.n2805 GNDA.n6 0.15675
R4787 GNDA.n2811 GNDA.n6 0.15675
R4788 GNDA.n2812 GNDA.n2811 0.15675
R4789 GNDA.n2813 GNDA.n2812 0.15675
R4790 GNDA.n2813 GNDA.n4 0.15675
R4791 GNDA.n2817 GNDA.n4 0.15675
R4792 GNDA.n2818 GNDA.n2817 0.15675
R4793 GNDA.n2819 GNDA.n2818 0.15675
R4794 GNDA.n2819 GNDA.n1 0.15675
R4795 GNDA.n2716 GNDA.n36 0.141125
R4796 GNDA.n2476 GNDA.n37 0.1321
R4797 GNDA.n167 GNDA.n124 0.131895
R4798 GNDA.n1677 GNDA.n1676 0.1255
R4799 GNDA.n1764 GNDA.n1109 0.1255
R4800 GNDA.n1817 GNDA.n1084 0.1255
R4801 GNDA.n2478 GNDA 0.1255
R4802 GNDA.n2511 GNDA.n2510 0.109875
R4803 GNDA.n134 GNDA.n131 0.09425
R4804 GNDA.n138 GNDA.n135 0.09425
R4805 GNDA.n142 GNDA.n139 0.09425
R4806 GNDA.n145 GNDA.n144 0.09425
R4807 GNDA.n316 GNDA.n315 0.09425
R4808 GNDA.n321 GNDA.n320 0.09425
R4809 GNDA.n167 GNDA.n166 0.063
R4810 GNDA.n162 GNDA.n134 0.063
R4811 GNDA.n156 GNDA.n138 0.063
R4812 GNDA.n150 GNDA.n142 0.063
R4813 GNDA.n144 GNDA.n118 0.063
R4814 GNDA.n315 GNDA.n116 0.063
R4815 GNDA.n322 GNDA.n321 0.063
R4816 GNDA GNDA.n2477 0.063
R4817 GNDA.n1677 GNDA.n1674 0.0626438
R4818 GNDA.n1109 GNDA.n1108 0.0626438
R4819 GNDA.n1814 GNDA.n1084 0.0626438
R4820 GNDA GNDA.n1566 0.0517
R4821 GNDA GNDA.n1152 0.0517
R4822 GNDA GNDA.n488 0.0517
R4823 GNDA.n776 GNDA 0.0517
R4824 GNDA.n1006 GNDA 0.0517
R4825 GNDA.n2130 GNDA 0.0517
R4826 GNDA GNDA.n2273 0.0517
R4827 GNDA.n1372 GNDA 0.0517
R4828 GNDA.n2031 GNDA 0.0517
R4829 GNDA.n2512 GNDA.n2511 0.047375
R4830 GNDA.n2717 GNDA.n2716 0.0430057
R4831 GNDA.n1768 GNDA.n1105 0.0421667
R4832 GNDA GNDA.n2744 0.03175
R4833 GNDA.n1789 GNDA.n1772 0.0217373
R4834 GNDA.n1102 GNDA.n1100 0.0217373
R4835 GNDA.n1770 GNDA.n1769 0.0217373
R4836 GNDA.n1767 GNDA.n1107 0.0217373
R4837 GNDA.n1772 GNDA.n1101 0.0217373
R4838 GNDA.n1771 GNDA.n1100 0.0217373
R4839 GNDA.n1769 GNDA.n1104 0.0217373
R4840 GNDA.n1107 GNDA.n1104 0.0217373
R4841 GNDA.n1791 GNDA.n1101 0.0217373
R4842 GNDA.n1790 GNDA.n1102 0.0217373
R4843 GNDA.n1792 GNDA.n1791 0.0217373
R4844 GNDA.n1766 GNDA.n1103 0.0217373
R4845 GNDA.n1105 GNDA.n1103 0.0217373
R4846 V_CONT.n0 V_CONT.t11 1156.8
R4847 V_CONT.n1 V_CONT.n0 964
R4848 VCO_FD_magic_0.V_CONT V_CONT.n2 562.333
R4849 V_CONT.n2 V_CONT.n1 433.8
R4850 V_CONT.n5 V_CONT.t8 377.567
R4851 V_CONT.n4 V_CONT.t12 297.233
R4852 V_CONT.n9 V_CONT.n8 242.903
R4853 V_CONT.n6 V_CONT.n4 237.851
R4854 V_CONT.n6 V_CONT.n5 232.809
R4855 V_CONT.n5 V_CONT.t9 216.9
R4856 V_CONT.n2 V_CONT.t10 192.8
R4857 V_CONT.n1 V_CONT.t14 192.8
R4858 V_CONT.n0 V_CONT.t15 192.8
R4859 V_CONT.n9 V_CONT.n7 172.502
R4860 VCO_FD_magic_0.V_CONT V_CONT.n13 168.405
R4861 V_CONT.n3 V_CONT.t6 166.368
R4862 V_CONT.n4 V_CONT.t13 136.567
R4863 V_CONT.n12 V_CONT.n11 125.225
R4864 V_CONT.n11 V_CONT.n10 106.662
R4865 V_CONT.n12 opamp_cell_4_0.VIN- 49.9172
R4866 V_CONT.n7 V_CONT.t4 24.6255
R4867 V_CONT.n7 V_CONT.t2 24.6255
R4868 V_CONT.n8 V_CONT.t7 24.6255
R4869 V_CONT.n8 V_CONT.t1 24.6255
R4870 V_CONT.n11 V_CONT.n9 22.4005
R4871 V_CONT.n10 V_CONT.t3 15.0005
R4872 V_CONT.n10 V_CONT.t0 15.0005
R4873 V_CONT.n13 V_CONT.n12 11.5239
R4874 V_CONT.n3 V_CONT.t5 3.82928
R4875 opamp_cell_4_0.VIN- V_CONT.n6 1.29217
R4876 V_CONT.n13 V_CONT.n3 0.09475
R4877 a_6200_5250.n4 a_6200_5250.n0 427.647
R4878 a_6200_5250.n1 a_6200_5250.t6 321.334
R4879 a_6200_5250.n5 a_6200_5250.n4 210.601
R4880 a_6200_5250.n2 a_6200_5250.n1 208.868
R4881 a_6200_5250.n3 a_6200_5250.t2 174.056
R4882 a_6200_5250.n4 a_6200_5250.n3 152
R4883 a_6200_5250.n1 a_6200_5250.t7 112.468
R4884 a_6200_5250.n2 a_6200_5250.t4 112.468
R4885 a_6200_5250.n3 a_6200_5250.n2 61.5894
R4886 a_6200_5250.n5 a_6200_5250.t5 60.0005
R4887 a_6200_5250.t3 a_6200_5250.n5 60.0005
R4888 a_6200_5250.n0 a_6200_5250.t1 49.2505
R4889 a_6200_5250.n0 a_6200_5250.t0 49.2505
R4890 a_5970_4630.n8 a_5970_4630.n6 522.322
R4891 a_5970_4630.n3 a_5970_4630.t6 384.967
R4892 a_5970_4630.n0 a_5970_4630.t9 384.967
R4893 a_5970_4630.n3 a_5970_4630.t8 379.166
R4894 a_5970_4630.t10 a_5970_4630.n0 376.56
R4895 a_5970_4630.n5 a_5970_4630.n1 315.647
R4896 a_5970_4630.n4 a_5970_4630.n2 315.647
R4897 a_5970_4630.n11 a_5970_4630.n10 314.502
R4898 a_5970_4630.n8 a_5970_4630.n7 160.721
R4899 a_5970_4630.n5 a_5970_4630.n4 83.2005
R4900 a_5970_4630.n1 a_5970_4630.t1 49.2505
R4901 a_5970_4630.n1 a_5970_4630.t5 49.2505
R4902 a_5970_4630.n2 a_5970_4630.t4 49.2505
R4903 a_5970_4630.n2 a_5970_4630.t7 49.2505
R4904 a_5970_4630.t10 a_5970_4630.n11 49.2505
R4905 a_5970_4630.n11 a_5970_4630.t0 49.2505
R4906 a_5970_4630.n10 a_5970_4630.n9 42.6672
R4907 a_5970_4630.n9 a_5970_4630.n8 37.763
R4908 a_5970_4630.n9 a_5970_4630.n5 23.4672
R4909 a_5970_4630.n6 a_5970_4630.t11 19.7005
R4910 a_5970_4630.n6 a_5970_4630.t2 19.7005
R4911 a_5970_4630.n7 a_5970_4630.t12 19.7005
R4912 a_5970_4630.n7 a_5970_4630.t3 19.7005
R4913 a_5970_4630.n4 a_5970_4630.n3 16.0005
R4914 a_5970_4630.n10 a_5970_4630.n0 16.0005
R4915 VDDA.t164 VDDA.t220 2804.76
R4916 VDDA.t144 VDDA.t111 2533.33
R4917 VDDA.t15 VDDA.t389 2307.14
R4918 VDDA.t158 VDDA.t185 2216.67
R4919 VDDA.t400 VDDA.t55 2216.67
R4920 VDDA.t53 VDDA.t206 2216.67
R4921 VDDA.t98 VDDA.t77 2126.19
R4922 VDDA.t47 VDDA.t190 1538.1
R4923 VDDA.t340 VDDA.t176 1492.86
R4924 VDDA.t399 VDDA.t225 1492.86
R4925 VDDA.t219 VDDA.t387 1317.78
R4926 VDDA.t90 VDDA.n91 1289.29
R4927 VDDA.t19 VDDA.n90 1289.29
R4928 VDDA.t414 VDDA.t234 1130.95
R4929 VDDA.t5 VDDA.t57 1130.95
R4930 VDDA.t11 VDDA.t116 1130.95
R4931 VDDA.t201 VDDA.t209 1130.95
R4932 VDDA.t37 VDDA.t43 1130.95
R4933 VDDA.t371 VDDA.n97 927.381
R4934 VDDA.t393 VDDA.n95 927.381
R4935 VDDA.t75 VDDA.n94 927.381
R4936 VDDA.t107 VDDA.n92 927.381
R4937 VDDA.n86 VDDA.n75 831.25
R4938 VDDA.n80 VDDA.n78 831.25
R4939 VDDA.n957 VDDA.n949 831.25
R4940 VDDA.n952 VDDA.n951 831.25
R4941 VDDA.n946 VDDA.n938 831.25
R4942 VDDA.n941 VDDA.n940 831.25
R4943 VDDA.n236 VDDA.t78 726.734
R4944 VDDA.n238 VDDA.t38 726.734
R4945 VDDA.t275 VDDA.n390 708.125
R4946 VDDA.n413 VDDA.t275 708.125
R4947 VDDA.n410 VDDA.t337 708.125
R4948 VDDA.t337 VDDA.n391 708.125
R4949 VDDA.t289 VDDA.n370 708.125
R4950 VDDA.n423 VDDA.t289 708.125
R4951 VDDA.n420 VDDA.t269 708.125
R4952 VDDA.t269 VDDA.n371 708.125
R4953 VDDA.t317 VDDA.n603 708.125
R4954 VDDA.n610 VDDA.t317 708.125
R4955 VDDA.t282 VDDA.n630 708.125
R4956 VDDA.n646 VDDA.t282 708.125
R4957 VDDA.t302 VDDA.n617 708.125
R4958 VDDA.n656 VDDA.t302 708.125
R4959 VDDA.n607 VDDA.t334 694.444
R4960 VDDA.t334 VDDA.n604 694.444
R4961 VDDA.n96 VDDA.t159 663.801
R4962 VDDA.n53 VDDA.t401 663.801
R4963 VDDA.n93 VDDA.t54 663.801
R4964 VDDA.n35 VDDA.t16 663.801
R4965 VDDA.n17 VDDA.t165 663.801
R4966 VDDA.n89 VDDA.t212 663.801
R4967 VDDA.n412 VDDA.t274 657.76
R4968 VDDA.n422 VDDA.t288 657.76
R4969 VDDA.n67 VDDA.n66 647.933
R4970 VDDA.n134 VDDA.n133 647.933
R4971 VDDA.n152 VDDA.n59 647.933
R4972 VDDA.n158 VDDA.n56 647.933
R4973 VDDA.n49 VDDA.n48 647.933
R4974 VDDA.n179 VDDA.n178 647.933
R4975 VDDA.n197 VDDA.n41 647.933
R4976 VDDA.n203 VDDA.n38 647.933
R4977 VDDA.n219 VDDA.n218 647.933
R4978 VDDA.n29 VDDA.n28 647.933
R4979 VDDA.n245 VDDA.n23 647.933
R4980 VDDA.n252 VDDA.n20 647.933
R4981 VDDA.n8 VDDA.n7 647.933
R4982 VDDA.n291 VDDA.n290 647.933
R4983 VDDA.n271 VDDA.n12 646.715
R4984 VDDA.n609 VDDA.t316 640.794
R4985 VDDA.n645 VDDA.t281 640.794
R4986 VDDA.n655 VDDA.t301 640.794
R4987 VDDA.n97 VDDA.t158 610.715
R4988 VDDA.n95 VDDA.t400 610.715
R4989 VDDA.n94 VDDA.t53 610.715
R4990 VDDA.n92 VDDA.t15 610.715
R4991 VDDA.n91 VDDA.t164 610.715
R4992 VDDA.n90 VDDA.t211 610.715
R4993 VDDA.n556 VDDA.n554 587.407
R4994 VDDA.n560 VDDA.n557 587.407
R4995 VDDA.n586 VDDA.n585 587.407
R4996 VDDA.n581 VDDA.n547 587.407
R4997 VDDA.n83 VDDA.n75 585
R4998 VDDA.n82 VDDA.n78 585
R4999 VDDA.n950 VDDA.n949 585
R5000 VDDA.n954 VDDA.n952 585
R5001 VDDA.n850 VDDA.n844 585
R5002 VDDA.n845 VDDA.n844 585
R5003 VDDA.n856 VDDA.n344 585
R5004 VDDA.n860 VDDA.n344 585
R5005 VDDA.n801 VDDA.n350 585
R5006 VDDA.n796 VDDA.n350 585
R5007 VDDA.n777 VDDA.n772 585
R5008 VDDA.n781 VDDA.n772 585
R5009 VDDA.n939 VDDA.n938 585
R5010 VDDA.n943 VDDA.n941 585
R5011 VDDA.n841 VDDA.n835 585
R5012 VDDA.n836 VDDA.n835 585
R5013 VDDA.n358 VDDA.n351 585
R5014 VDDA.n353 VDDA.n351 585
R5015 VDDA.n585 VDDA.n584 585
R5016 VDDA.n583 VDDA.n581 585
R5017 VDDA.n567 VDDA.n556 585
R5018 VDDA.n564 VDDA.n557 585
R5019 VDDA.n488 VDDA.n481 585
R5020 VDDA.n466 VDDA.n458 585
R5021 VDDA.n760 VDDA.n664 585
R5022 VDDA.n753 VDDA.n664 585
R5023 VDDA.n750 VDDA.n749 585
R5024 VDDA.n749 VDDA.n748 585
R5025 VDDA.n719 VDDA.n718 585
R5026 VDDA.n719 VDDA.n708 585
R5027 VDDA.t333 VDDA.n608 557.783
R5028 VDDA.t336 VDDA.n411 540.818
R5029 VDDA.t268 VDDA.n421 540.818
R5030 VDDA.n99 VDDA.t430 537.492
R5031 VDDA.n110 VDDA.t427 537.491
R5032 VDDA.n87 VDDA.t425 537.491
R5033 VDDA.t304 VDDA.n644 523.855
R5034 VDDA.t310 VDDA.n654 523.855
R5035 VDDA.t387 VDDA.t414 497.62
R5036 VDDA.t234 VDDA.t371 497.62
R5037 VDDA.t185 VDDA.t5 497.62
R5038 VDDA.t57 VDDA.t393 497.62
R5039 VDDA.t55 VDDA.t11 497.62
R5040 VDDA.t116 VDDA.t75 497.62
R5041 VDDA.t206 VDDA.t201 497.62
R5042 VDDA.t209 VDDA.t107 497.62
R5043 VDDA.t389 VDDA.t340 497.62
R5044 VDDA.t176 VDDA.t98 497.62
R5045 VDDA.t77 VDDA.t37 497.62
R5046 VDDA.t43 VDDA.t47 497.62
R5047 VDDA.t190 VDDA.t90 497.62
R5048 VDDA.t220 VDDA.t72 497.62
R5049 VDDA.t72 VDDA.t399 497.62
R5050 VDDA.t225 VDDA.t144 497.62
R5051 VDDA.t111 VDDA.t19 497.62
R5052 VDDA.t343 VDDA.n76 465.079
R5053 VDDA.n81 VDDA.t343 465.079
R5054 VDDA.n956 VDDA.t208 465.079
R5055 VDDA.t208 VDDA.n955 465.079
R5056 VDDA.n945 VDDA.t14 465.079
R5057 VDDA.t14 VDDA.n944 465.079
R5058 VDDA.n105 VDDA.t52 464.281
R5059 VDDA.n102 VDDA.t52 464.281
R5060 VDDA.n113 VDDA.t27 464.281
R5061 VDDA.t27 VDDA.n72 464.281
R5062 VDDA.t163 VDDA.n825 464.281
R5063 VDDA.n827 VDDA.t163 464.281
R5064 VDDA.n933 VDDA.t231 464.281
R5065 VDDA.t231 VDDA.n932 464.281
R5066 VDDA.n970 VDDA.t365 464.281
R5067 VDDA.t365 VDDA.n969 464.281
R5068 VDDA.n914 VDDA.t110 464.281
R5069 VDDA.t110 VDDA.n913 464.281
R5070 VDDA.n892 VDDA.t115 464.281
R5071 VDDA.t115 VDDA.n891 464.281
R5072 VDDA.n822 VDDA.t248 464.281
R5073 VDDA.t248 VDDA.n821 464.281
R5074 VDDA.t82 VDDA.n922 464.281
R5075 VDDA.n923 VDDA.t82 464.281
R5076 VDDA.t257 VDDA.n317 464.281
R5077 VDDA.n960 VDDA.t257 464.281
R5078 VDDA.t161 VDDA.n325 464.281
R5079 VDDA.n895 VDDA.t161 464.281
R5080 VDDA.t386 VDDA.n810 464.281
R5081 VDDA.n811 VDDA.t386 464.281
R5082 VDDA.n612 VDDA.t315 422.384
R5083 VDDA.n605 VDDA.t332 422.384
R5084 VDDA.n648 VDDA.t280 418.368
R5085 VDDA.n641 VDDA.t303 418.368
R5086 VDDA.n658 VDDA.t300 418.368
R5087 VDDA.n651 VDDA.t309 418.368
R5088 VDDA.n341 VDDA.t426 415.336
R5089 VDDA.t274 VDDA.t120 407.144
R5090 VDDA.t120 VDDA.t227 407.144
R5091 VDDA.t227 VDDA.t241 407.144
R5092 VDDA.t241 VDDA.t7 407.144
R5093 VDDA.t7 VDDA.t9 407.144
R5094 VDDA.t9 VDDA.t404 407.144
R5095 VDDA.t404 VDDA.t118 407.144
R5096 VDDA.t118 VDDA.t369 407.144
R5097 VDDA.t369 VDDA.t178 407.144
R5098 VDDA.t178 VDDA.t96 407.144
R5099 VDDA.t96 VDDA.t338 407.144
R5100 VDDA.t338 VDDA.t199 407.144
R5101 VDDA.t199 VDDA.t197 407.144
R5102 VDDA.t197 VDDA.t79 407.144
R5103 VDDA.t79 VDDA.t39 407.144
R5104 VDDA.t39 VDDA.t92 407.144
R5105 VDDA.t92 VDDA.t243 407.144
R5106 VDDA.t243 VDDA.t87 407.144
R5107 VDDA.t87 VDDA.t336 407.144
R5108 VDDA.t288 VDDA.t49 407.144
R5109 VDDA.t49 VDDA.t344 407.144
R5110 VDDA.t344 VDDA.t346 407.144
R5111 VDDA.t346 VDDA.t360 407.144
R5112 VDDA.t360 VDDA.t356 407.144
R5113 VDDA.t356 VDDA.t180 407.144
R5114 VDDA.t180 VDDA.t249 407.144
R5115 VDDA.t249 VDDA.t350 407.144
R5116 VDDA.t350 VDDA.t352 407.144
R5117 VDDA.t352 VDDA.t354 407.144
R5118 VDDA.t354 VDDA.t358 407.144
R5119 VDDA.t358 VDDA.t64 407.144
R5120 VDDA.t64 VDDA.t402 407.144
R5121 VDDA.t402 VDDA.t348 407.144
R5122 VDDA.t348 VDDA.t362 407.144
R5123 VDDA.t362 VDDA.t239 407.144
R5124 VDDA.t239 VDDA.t213 407.144
R5125 VDDA.t213 VDDA.t59 407.144
R5126 VDDA.t59 VDDA.t268 407.144
R5127 VDDA.n451 VDDA.t306 384.967
R5128 VDDA.n493 VDDA.t321 384.967
R5129 VDDA.n471 VDDA.t276 384.967
R5130 VDDA.n476 VDDA.t270 384.967
R5131 VDDA.n95 VDDA.n53 382.8
R5132 VDDA.n94 VDDA.n93 382.8
R5133 VDDA.n92 VDDA.n35 382.8
R5134 VDDA.n91 VDDA.n17 382.8
R5135 VDDA.n90 VDDA.n89 382.8
R5136 VDDA.n97 VDDA.n96 382.8
R5137 VDDA.n488 VDDA.t293 374.878
R5138 VDDA.t316 VDDA.t63 373.214
R5139 VDDA.t63 VDDA.t222 373.214
R5140 VDDA.t222 VDDA.t333 373.214
R5141 VDDA.t281 VDDA.t194 373.214
R5142 VDDA.t194 VDDA.t395 373.214
R5143 VDDA.t395 VDDA.t383 373.214
R5144 VDDA.t383 VDDA.t174 373.214
R5145 VDDA.t174 VDDA.t381 373.214
R5146 VDDA.t381 VDDA.t146 373.214
R5147 VDDA.t146 VDDA.t168 373.214
R5148 VDDA.t168 VDDA.t156 373.214
R5149 VDDA.t156 VDDA.t406 373.214
R5150 VDDA.t406 VDDA.t148 373.214
R5151 VDDA.t148 VDDA.t304 373.214
R5152 VDDA.t301 VDDA.t154 373.214
R5153 VDDA.t154 VDDA.t408 373.214
R5154 VDDA.t408 VDDA.t412 373.214
R5155 VDDA.t412 VDDA.t397 373.214
R5156 VDDA.t397 VDDA.t410 373.214
R5157 VDDA.t410 VDDA.t170 373.214
R5158 VDDA.t170 VDDA.t172 373.214
R5159 VDDA.t172 VDDA.t377 373.214
R5160 VDDA.t377 VDDA.t192 373.214
R5161 VDDA.t192 VDDA.t379 373.214
R5162 VDDA.t379 VDDA.t310 373.214
R5163 VDDA.n415 VDDA.t273 370.168
R5164 VDDA.n408 VDDA.t335 370.168
R5165 VDDA.n425 VDDA.t287 370.168
R5166 VDDA.n418 VDDA.t267 370.168
R5167 VDDA.n538 VDDA.t290 360.868
R5168 VDDA.n592 VDDA.t312 360.868
R5169 VDDA.t319 VDDA.t245 360.346
R5170 VDDA.t245 VDDA.t29 360.346
R5171 VDDA.t29 VDDA.t421 360.346
R5172 VDDA.t421 VDDA.t21 360.346
R5173 VDDA.t21 VDDA.t297 360.346
R5174 VDDA.t391 VDDA.t326 360.346
R5175 VDDA.t100 VDDA.t391 360.346
R5176 VDDA.t41 VDDA.t100 360.346
R5177 VDDA.t83 VDDA.t41 360.346
R5178 VDDA.t329 VDDA.t83 360.346
R5179 VDDA.n110 VDDA.t262 359.752
R5180 VDDA.n87 VDDA.t261 359.752
R5181 VDDA.n99 VDDA.t260 359.752
R5182 VDDA.n457 VDDA.t283 352.834
R5183 VDDA.n632 VDDA.t305 351.793
R5184 VDDA.n619 VDDA.t311 351.793
R5185 VDDA.n714 VDDA.t319 343.966
R5186 VDDA.n752 VDDA.t297 343.966
R5187 VDDA.t326 VDDA.n752 343.966
R5188 VDDA.n758 VDDA.t329 343.966
R5189 VDDA.n472 VDDA.t279 341.752
R5190 VDDA.n477 VDDA.t272 341.752
R5191 VDDA.n492 VDDA.t324 341.752
R5192 VDDA.n452 VDDA.t308 341.752
R5193 VDDA.n747 VDDA.t325 336.329
R5194 VDDA.n747 VDDA.t296 336.329
R5195 VDDA.n709 VDDA.t318 320.7
R5196 VDDA.n761 VDDA.t328 320.7
R5197 VDDA.n450 VDDA.n448 315.647
R5198 VDDA.n444 VDDA.n443 315.647
R5199 VDDA.n475 VDDA.n474 315.647
R5200 VDDA.n470 VDDA.n469 315.647
R5201 VDDA.n495 VDDA.n447 315.647
R5202 VDDA.n494 VDDA.n449 315.647
R5203 VDDA.n324 VDDA.t205 315.25
R5204 VDDA.t189 VDDA.t238 314.113
R5205 VDDA.t2 VDDA.t89 314.113
R5206 VDDA.t307 VDDA.n452 304.659
R5207 VDDA.n640 VDDA.n639 301.933
R5208 VDDA.n638 VDDA.n637 301.933
R5209 VDDA.n636 VDDA.n635 301.933
R5210 VDDA.n634 VDDA.n633 301.933
R5211 VDDA.n629 VDDA.n628 301.933
R5212 VDDA.n627 VDDA.n626 301.933
R5213 VDDA.n625 VDDA.n624 301.933
R5214 VDDA.n623 VDDA.n622 301.933
R5215 VDDA.n621 VDDA.n620 301.933
R5216 VDDA.n616 VDDA.n615 301.933
R5217 VDDA.n407 VDDA.n406 299.231
R5218 VDDA.n405 VDDA.n404 299.231
R5219 VDDA.n403 VDDA.n402 299.231
R5220 VDDA.n401 VDDA.n400 299.231
R5221 VDDA.n399 VDDA.n398 299.231
R5222 VDDA.n397 VDDA.n396 299.231
R5223 VDDA.n395 VDDA.n394 299.231
R5224 VDDA.n393 VDDA.n392 299.231
R5225 VDDA.n389 VDDA.n388 299.231
R5226 VDDA.n387 VDDA.n386 299.231
R5227 VDDA.n385 VDDA.n384 299.231
R5228 VDDA.n383 VDDA.n382 299.231
R5229 VDDA.n381 VDDA.n380 299.231
R5230 VDDA.n379 VDDA.n378 299.231
R5231 VDDA.n377 VDDA.n376 299.231
R5232 VDDA.n375 VDDA.n374 299.231
R5233 VDDA.n373 VDDA.n372 299.231
R5234 VDDA.n369 VDDA.n368 299.231
R5235 VDDA.n749 VDDA.n672 291.363
R5236 VDDA.n745 VDDA.n670 291.363
R5237 VDDA.n746 VDDA.n745 291.363
R5238 VDDA.n848 VDDA.n844 290.733
R5239 VDDA.n854 VDDA.n344 290.733
R5240 VDDA.n799 VDDA.n350 290.733
R5241 VDDA.n775 VDDA.n772 290.733
R5242 VDDA.n839 VDDA.n835 290.733
R5243 VDDA.n352 VDDA.n351 290.733
R5244 VDDA.n486 VDDA.n481 290.733
R5245 VDDA.n482 VDDA.n481 290.733
R5246 VDDA.n464 VDDA.n458 290.733
R5247 VDDA.n459 VDDA.n458 290.733
R5248 VDDA.n754 VDDA.n664 290.733
R5249 VDDA.n719 VDDA.n707 290.733
R5250 VDDA.t33 VDDA.t291 251.471
R5251 VDDA.t132 VDDA.t33 251.471
R5252 VDDA.t136 VDDA.t132 251.471
R5253 VDDA.t419 VDDA.t136 251.471
R5254 VDDA.t31 VDDA.t419 251.471
R5255 VDDA.t252 VDDA.t31 251.471
R5256 VDDA.t125 VDDA.t252 251.471
R5257 VDDA.t23 VDDA.t125 251.471
R5258 VDDA.t182 VDDA.t23 251.471
R5259 VDDA.t367 VDDA.t182 251.471
R5260 VDDA.t417 VDDA.t367 251.471
R5261 VDDA.t103 VDDA.t417 251.471
R5262 VDDA.t130 VDDA.t103 251.471
R5263 VDDA.t141 VDDA.t130 251.471
R5264 VDDA.t123 VDDA.t141 251.471
R5265 VDDA.t139 VDDA.t123 251.471
R5266 VDDA.t313 VDDA.t139 251.471
R5267 VDDA.n934 VDDA.n933 243.698
R5268 VDDA.n971 VDDA.n970 243.698
R5269 VDDA.n915 VDDA.n914 243.698
R5270 VDDA.n893 VDDA.n892 243.698
R5271 VDDA.n823 VDDA.n822 243.698
R5272 VDDA.n923 VDDA.n920 243.698
R5273 VDDA.n964 VDDA.n960 243.698
R5274 VDDA.n899 VDDA.n895 243.698
R5275 VDDA.n811 VDDA.n808 243.698
R5276 VDDA.n107 VDDA.n106 238.367
R5277 VDDA.n101 VDDA.n88 238.367
R5278 VDDA.n115 VDDA.n114 238.367
R5279 VDDA.n118 VDDA.n117 238.367
R5280 VDDA.n86 VDDA.n85 238.367
R5281 VDDA.n80 VDDA.n79 238.367
R5282 VDDA.n919 VDDA.n301 238.367
R5283 VDDA.n958 VDDA.n957 238.367
R5284 VDDA.n951 VDDA.n918 238.367
R5285 VDDA.n917 VDDA.n316 238.367
R5286 VDDA.n910 VDDA.n319 238.367
R5287 VDDA.n888 VDDA.n327 238.367
R5288 VDDA.n807 VDDA.n335 238.367
R5289 VDDA.n927 VDDA.n302 238.367
R5290 VDDA.n947 VDDA.n946 238.367
R5291 VDDA.n974 VDDA.n973 238.367
R5292 VDDA.n902 VDDA.n901 238.367
R5293 VDDA.n815 VDDA.n331 238.367
R5294 VDDA.n940 VDDA.n936 238.367
R5295 VDDA.n411 VDDA.n410 238.367
R5296 VDDA.n411 VDDA.n391 238.367
R5297 VDDA.n421 VDDA.n420 238.367
R5298 VDDA.n421 VDDA.n371 238.367
R5299 VDDA.n588 VDDA.n587 238.367
R5300 VDDA.n608 VDDA.n607 238.367
R5301 VDDA.n608 VDDA.n604 238.367
R5302 VDDA.n644 VDDA.n643 238.367
R5303 VDDA.n644 VDDA.n631 238.367
R5304 VDDA.n654 VDDA.n653 238.367
R5305 VDDA.n654 VDDA.n618 238.367
R5306 VDDA.t291 VDDA.n572 237.5
R5307 VDDA.n589 VDDA.t313 237.5
R5308 VDDA.n482 VDDA.n453 233.841
R5309 VDDA.n459 VDDA.n455 233.841
R5310 VDDA.n851 VDDA.n850 230.308
R5311 VDDA.n845 VDDA.n804 230.308
R5312 VDDA.n857 VDDA.n856 230.308
R5313 VDDA.n860 VDDA.n859 230.308
R5314 VDDA.n802 VDDA.n801 230.308
R5315 VDDA.n796 VDDA.n346 230.308
R5316 VDDA.n778 VDDA.n777 230.308
R5317 VDDA.n781 VDDA.n780 230.308
R5318 VDDA.n842 VDDA.n841 230.308
R5319 VDDA.n358 VDDA.n348 230.308
R5320 VDDA.n353 VDDA.n347 230.308
R5321 VDDA.n836 VDDA.n833 230.308
R5322 VDDA.n489 VDDA.n488 230.308
R5323 VDDA.n760 VDDA.n759 230.308
R5324 VDDA.n757 VDDA.n753 230.308
R5325 VDDA.n751 VDDA.n750 230.308
R5326 VDDA.n748 VDDA.n667 230.308
R5327 VDDA.t203 VDDA.t3 222.178
R5328 VDDA.n74 VDDA.t342 219.232
R5329 VDDA.t236 VDDA.n74 219.232
R5330 VDDA.n116 VDDA.t26 219.232
R5331 VDDA.n108 VDDA.t51 219.232
R5332 VDDA.n852 VDDA.n832 199.195
R5333 VDDA.n681 VDDA.n680 196.502
R5334 VDDA.n678 VDDA.n677 196.502
R5335 VDDA.n744 VDDA.n743 196.502
R5336 VDDA.n735 VDDA.n700 196.502
R5337 VDDA.n728 VDDA.n703 196.502
R5338 VDDA.n721 VDDA.n720 196.502
R5339 VDDA.n827 VDDA.n806 190.333
R5340 VDDA.n110 VDDA.t26 185.002
R5341 VDDA.t236 VDDA.n87 185.002
R5342 VDDA.n99 VDDA.t51 185.002
R5343 VDDA.n492 VDDA.n491 185.001
R5344 VDDA.n478 VDDA.n477 185.001
R5345 VDDA.n473 VDDA.n472 185.001
R5346 VDDA.n84 VDDA.n83 185
R5347 VDDA.n82 VDDA.n77 185
R5348 VDDA.n112 VDDA.n109 185
R5349 VDDA.n111 VDDA.n73 185
R5350 VDDA.n104 VDDA.n98 185
R5351 VDDA.n103 VDDA.n100 185
R5352 VDDA.n357 VDDA.n356 185
R5353 VDDA.n355 VDDA.n354 185
R5354 VDDA.n840 VDDA.n834 185
R5355 VDDA.n838 VDDA.n837 185
R5356 VDDA.n814 VDDA.n813 185
R5357 VDDA.n812 VDDA.n809 185
R5358 VDDA.n896 VDDA.n326 185
R5359 VDDA.n898 VDDA.n897 185
R5360 VDDA.n961 VDDA.n318 185
R5361 VDDA.n963 VDDA.n962 185
R5362 VDDA.n939 VDDA.n937 185
R5363 VDDA.n943 VDDA.n942 185
R5364 VDDA.n926 VDDA.n925 185
R5365 VDDA.n924 VDDA.n921 185
R5366 VDDA.n776 VDDA.n774 185
R5367 VDDA.n773 VDDA.n771 185
R5368 VDDA.n800 VDDA.n349 185
R5369 VDDA.n798 VDDA.n797 185
R5370 VDDA.n855 VDDA.n853 185
R5371 VDDA.n345 VDDA.n343 185
R5372 VDDA.n849 VDDA.n843 185
R5373 VDDA.n847 VDDA.n846 185
R5374 VDDA.n818 VDDA.n817 185
R5375 VDDA.n820 VDDA.n819 185
R5376 VDDA.n329 VDDA.n328 185
R5377 VDDA.n890 VDDA.n889 185
R5378 VDDA.n321 VDDA.n320 185
R5379 VDDA.n912 VDDA.n911 185
R5380 VDDA.n966 VDDA.n965 185
R5381 VDDA.n968 VDDA.n967 185
R5382 VDDA.n950 VDDA.n948 185
R5383 VDDA.n954 VDDA.n953 185
R5384 VDDA.n929 VDDA.n928 185
R5385 VDDA.n931 VDDA.n930 185
R5386 VDDA.n831 VDDA.n334 185
R5387 VDDA.n832 VDDA.n831 185
R5388 VDDA.n830 VDDA.n829 185
R5389 VDDA.n828 VDDA.n826 185
R5390 VDDA.n832 VDDA.n806 185
R5391 VDDA.n577 VDDA.n575 185
R5392 VDDA.n584 VDDA.n574 185
R5393 VDDA.n589 VDDA.n574 185
R5394 VDDA.n583 VDDA.n582 185
R5395 VDDA.n580 VDDA.n549 185
R5396 VDDA.n591 VDDA.n590 185
R5397 VDDA.n590 VDDA.n589 185
R5398 VDDA.n571 VDDA.n570 185
R5399 VDDA.n572 VDDA.n571 185
R5400 VDDA.n568 VDDA.n553 185
R5401 VDDA.n567 VDDA.n566 185
R5402 VDDA.n565 VDDA.n564 185
R5403 VDDA.n559 VDDA.n558 185
R5404 VDDA.n561 VDDA.n552 185
R5405 VDDA.n572 VDDA.n552 185
R5406 VDDA.n487 VDDA.n480 185
R5407 VDDA.n485 VDDA.n479 185
R5408 VDDA.n490 VDDA.n479 185
R5409 VDDA.n484 VDDA.n483 185
R5410 VDDA.n467 VDDA.n466 185
R5411 VDDA.n468 VDDA.n467 185
R5412 VDDA.n465 VDDA.n456 185
R5413 VDDA.n463 VDDA.n462 185
R5414 VDDA.n461 VDDA.n460 185
R5415 VDDA.n671 VDDA.n668 185
R5416 VDDA.n674 VDDA.n673 185
R5417 VDDA.n666 VDDA.n665 185
R5418 VDDA.n756 VDDA.n755 185
R5419 VDDA.n718 VDDA.n710 185
R5420 VDDA.n714 VDDA.n710 185
R5421 VDDA.n717 VDDA.n716 185
R5422 VDDA.n712 VDDA.n711 185
R5423 VDDA.n713 VDDA.n708 185
R5424 VDDA.n714 VDDA.n713 185
R5425 VDDA.n779 VDDA.t203 172.38
R5426 VDDA.t105 VDDA.n803 172.38
R5427 VDDA.n858 VDDA.t68 172.38
R5428 VDDA.n748 VDDA.n747 166.63
R5429 VDDA.n116 VDDA.t74 158.333
R5430 VDDA.t196 VDDA.n108 158.333
R5431 VDDA.n100 VDDA.n98 150
R5432 VDDA.n109 VDDA.n73 150
R5433 VDDA.n84 VDDA.n77 150
R5434 VDDA.n930 VDDA.n928 150
R5435 VDDA.n953 VDDA.n948 150
R5436 VDDA.n967 VDDA.n965 150
R5437 VDDA.n911 VDDA.n320 150
R5438 VDDA.n889 VDDA.n328 150
R5439 VDDA.n819 VDDA.n817 150
R5440 VDDA.n926 VDDA.n921 150
R5441 VDDA.n942 VDDA.n937 150
R5442 VDDA.n963 VDDA.n318 150
R5443 VDDA.n898 VDDA.n326 150
R5444 VDDA.n814 VDDA.n809 150
R5445 VDDA.n831 VDDA.n830 150
R5446 VDDA.n826 VDDA.n806 150
R5447 VDDA.n575 VDDA.n574 150
R5448 VDDA.n582 VDDA.n574 150
R5449 VDDA.n590 VDDA.n549 150
R5450 VDDA.n571 VDDA.n553 150
R5451 VDDA.n566 VDDA.n565 150
R5452 VDDA.n558 VDDA.n552 150
R5453 VDDA.t152 VDDA.t223 145.038
R5454 VDDA.n593 VDDA.n546 141.712
R5455 VDDA.n594 VDDA.n545 141.712
R5456 VDDA.n595 VDDA.n544 141.712
R5457 VDDA.n596 VDDA.n543 141.712
R5458 VDDA.n597 VDDA.n542 141.712
R5459 VDDA.n598 VDDA.n541 141.712
R5460 VDDA.n599 VDDA.n540 141.712
R5461 VDDA.n600 VDDA.n539 141.712
R5462 VDDA.n824 VDDA.n816 137.904
R5463 VDDA.n900 VDDA.n894 137.904
R5464 VDDA.n779 VDDA.t45 126.412
R5465 VDDA.n803 VDDA.t3 126.412
R5466 VDDA.n858 VDDA.t105 126.412
R5467 VDDA.t68 VDDA.n852 126.412
R5468 VDDA.t237 VDDA.n75 123.126
R5469 VDDA.n78 VDDA.t237 123.126
R5470 VDDA.t167 VDDA.n949 123.126
R5471 VDDA.n952 VDDA.t167 123.126
R5472 VDDA.t364 VDDA.n938 123.126
R5473 VDDA.n941 VDDA.t364 123.126
R5474 VDDA.t292 VDDA.n556 123.126
R5475 VDDA.n557 VDDA.t292 123.126
R5476 VDDA.n585 VDDA.t314 123.126
R5477 VDDA.n581 VDDA.t314 123.126
R5478 VDDA.n846 VDDA.n843 120.001
R5479 VDDA.n853 VDDA.n345 120.001
R5480 VDDA.n797 VDDA.n349 120.001
R5481 VDDA.n774 VDDA.n773 120.001
R5482 VDDA.n837 VDDA.n834 120.001
R5483 VDDA.n356 VDDA.n355 120.001
R5484 VDDA.n480 VDDA.n479 120.001
R5485 VDDA.n483 VDDA.n479 120.001
R5486 VDDA.n467 VDDA.n456 120.001
R5487 VDDA.n462 VDDA.n461 120.001
R5488 VDDA.n756 VDDA.n666 120.001
R5489 VDDA.n673 VDDA.n668 120.001
R5490 VDDA.n716 VDDA.n710 120.001
R5491 VDDA.n713 VDDA.n712 120.001
R5492 VDDA.n526 VDDA.n432 119.737
R5493 VDDA.n519 VDDA.n435 119.737
R5494 VDDA.n512 VDDA.n438 119.737
R5495 VDDA.n505 VDDA.n441 119.737
R5496 VDDA.n497 VDDA.n446 119.737
R5497 VDDA.n491 VDDA.t322 119.656
R5498 VDDA.t74 VDDA.t236 109.615
R5499 VDDA.t26 VDDA.t196 109.615
R5500 VDDA.t51 VDDA.t219 109.615
R5501 VDDA.n490 VDDA.n478 108.779
R5502 VDDA.n972 VDDA.n916 107.258
R5503 VDDA.n972 VDDA.t256 103.427
R5504 VDDA.t13 VDDA.n959 103.427
R5505 VDDA.n959 VDDA.t166 103.427
R5506 VDDA.t81 VDDA.n935 103.427
R5507 VDDA.n916 VDDA.t160 95.7666
R5508 VDDA.t0 VDDA.t307 94.2753
R5509 VDDA.t254 VDDA.t0 94.2753
R5510 VDDA.t66 VDDA.t254 94.2753
R5511 VDDA.t217 VDDA.t66 94.2753
R5512 VDDA.t322 VDDA.t217 94.2753
R5513 VDDA.t232 VDDA.t229 94.2753
R5514 VDDA.t258 VDDA.t277 94.2753
R5515 VDDA.t70 VDDA.n473 94.2753
R5516 VDDA.t266 VDDA.t28 94.2753
R5517 VDDA.t264 VDDA.t263 94.2753
R5518 VDDA.t247 VDDA.t162 91.936
R5519 VDDA.t114 VDDA.t385 91.936
R5520 VDDA.n87 VDDA.n86 90.5056
R5521 VDDA.t204 VDDA.t109 84.2747
R5522 VDDA.t256 VDDA.t189 84.2747
R5523 VDDA.t238 VDDA.t13 84.2747
R5524 VDDA.t166 VDDA.t2 84.2747
R5525 VDDA.t89 VDDA.t81 84.2747
R5526 VDDA.t294 VDDA.t271 83.3974
R5527 VDDA.t375 VDDA.t134 83.3974
R5528 VDDA.n475 VDDA.n444 83.2005
R5529 VDDA.n470 VDDA.n444 83.2005
R5530 VDDA.n495 VDDA.n448 83.2005
R5531 VDDA.n495 VDDA.n494 83.2005
R5532 VDDA.n66 VDDA.t388 78.8005
R5533 VDDA.n66 VDDA.t415 78.8005
R5534 VDDA.n133 VDDA.t235 78.8005
R5535 VDDA.n133 VDDA.t372 78.8005
R5536 VDDA.n59 VDDA.t186 78.8005
R5537 VDDA.n59 VDDA.t6 78.8005
R5538 VDDA.n56 VDDA.t58 78.8005
R5539 VDDA.n56 VDDA.t394 78.8005
R5540 VDDA.n48 VDDA.t56 78.8005
R5541 VDDA.n48 VDDA.t12 78.8005
R5542 VDDA.n178 VDDA.t117 78.8005
R5543 VDDA.n178 VDDA.t76 78.8005
R5544 VDDA.n41 VDDA.t207 78.8005
R5545 VDDA.n41 VDDA.t202 78.8005
R5546 VDDA.n38 VDDA.t210 78.8005
R5547 VDDA.n38 VDDA.t108 78.8005
R5548 VDDA.n218 VDDA.t390 78.8005
R5549 VDDA.n218 VDDA.t341 78.8005
R5550 VDDA.n28 VDDA.t177 78.8005
R5551 VDDA.n28 VDDA.t99 78.8005
R5552 VDDA.n23 VDDA.t44 78.8005
R5553 VDDA.n23 VDDA.t48 78.8005
R5554 VDDA.n20 VDDA.t191 78.8005
R5555 VDDA.n20 VDDA.t91 78.8005
R5556 VDDA.n12 VDDA.t221 78.8005
R5557 VDDA.n12 VDDA.t73 78.8005
R5558 VDDA.n7 VDDA.t226 78.8005
R5559 VDDA.n7 VDDA.t145 78.8005
R5560 VDDA.n290 VDDA.t112 78.8005
R5561 VDDA.n290 VDDA.t20 78.8005
R5562 VDDA.t150 VDDA.t35 76.1455
R5563 VDDA.t284 VDDA.t265 76.1455
R5564 VDDA.n114 VDDA.n110 74.7688
R5565 VDDA.n106 VDDA.n99 74.7688
R5566 VDDA.n803 VDDA.n348 69.8479
R5567 VDDA.n803 VDDA.n347 69.8479
R5568 VDDA.n852 VDDA.n842 69.8479
R5569 VDDA.n852 VDDA.n833 69.8479
R5570 VDDA.n779 VDDA.n778 69.8479
R5571 VDDA.n780 VDDA.n779 69.8479
R5572 VDDA.n803 VDDA.n802 69.8479
R5573 VDDA.n803 VDDA.n346 69.8479
R5574 VDDA.n858 VDDA.n857 69.8479
R5575 VDDA.n859 VDDA.n858 69.8479
R5576 VDDA.n852 VDDA.n851 69.8479
R5577 VDDA.n852 VDDA.n804 69.8479
R5578 VDDA.n490 VDDA.n489 69.8479
R5579 VDDA.n490 VDDA.n453 69.8479
R5580 VDDA.n468 VDDA.n454 69.8479
R5581 VDDA.n468 VDDA.n455 69.8479
R5582 VDDA.n752 VDDA.n751 69.8479
R5583 VDDA.n752 VDDA.n667 69.8479
R5584 VDDA.n759 VDDA.n758 69.8479
R5585 VDDA.n758 VDDA.n757 69.8479
R5586 VDDA.n715 VDDA.n714 69.8479
R5587 VDDA.n496 VDDA.n495 69.3203
R5588 VDDA.t35 VDDA.t17 68.8936
R5589 VDDA.t265 VDDA.n468 68.8936
R5590 VDDA.n85 VDDA.n74 65.8183
R5591 VDDA.n79 VDDA.n74 65.8183
R5592 VDDA.n116 VDDA.n115 65.8183
R5593 VDDA.n117 VDDA.n116 65.8183
R5594 VDDA.n108 VDDA.n107 65.8183
R5595 VDDA.n108 VDDA.n88 65.8183
R5596 VDDA.n816 VDDA.n815 65.8183
R5597 VDDA.n816 VDDA.n808 65.8183
R5598 VDDA.n901 VDDA.n900 65.8183
R5599 VDDA.n900 VDDA.n899 65.8183
R5600 VDDA.n973 VDDA.n972 65.8183
R5601 VDDA.n972 VDDA.n964 65.8183
R5602 VDDA.n959 VDDA.n947 65.8183
R5603 VDDA.n959 VDDA.n936 65.8183
R5604 VDDA.n935 VDDA.n927 65.8183
R5605 VDDA.n935 VDDA.n920 65.8183
R5606 VDDA.n824 VDDA.n823 65.8183
R5607 VDDA.n824 VDDA.n807 65.8183
R5608 VDDA.n894 VDDA.n893 65.8183
R5609 VDDA.n894 VDDA.n327 65.8183
R5610 VDDA.n916 VDDA.n915 65.8183
R5611 VDDA.n916 VDDA.n319 65.8183
R5612 VDDA.n972 VDDA.n971 65.8183
R5613 VDDA.n972 VDDA.n917 65.8183
R5614 VDDA.n959 VDDA.n958 65.8183
R5615 VDDA.n959 VDDA.n918 65.8183
R5616 VDDA.n935 VDDA.n934 65.8183
R5617 VDDA.n935 VDDA.n919 65.8183
R5618 VDDA.n832 VDDA.n805 65.8183
R5619 VDDA.n589 VDDA.n588 65.8183
R5620 VDDA.n589 VDDA.n573 65.8183
R5621 VDDA.n572 VDDA.n550 65.8183
R5622 VDDA.n572 VDDA.n551 65.8183
R5623 VDDA.t271 VDDA.t373 61.6417
R5624 VDDA.t134 VDDA.t215 61.6417
R5625 VDDA.n364 VDDA.t428 58.8005
R5626 VDDA.n363 VDDA.t424 58.8005
R5627 VDDA.n1005 VDDA.n301 58.0576
R5628 VDDA.n975 VDDA.n316 58.0576
R5629 VDDA.n910 VDDA.n909 58.0576
R5630 VDDA.n888 VDDA.n887 58.0576
R5631 VDDA.n878 VDDA.n335 58.0576
R5632 VDDA.n1005 VDDA.n302 58.0576
R5633 VDDA.n975 VDDA.n974 58.0576
R5634 VDDA.n903 VDDA.n902 58.0576
R5635 VDDA.n886 VDDA.n331 58.0576
R5636 VDDA.n879 VDDA.n334 58.0576
R5637 VDDA.n845 VDDA.n338 57.2449
R5638 VDDA.n861 VDDA.n860 57.2449
R5639 VDDA.n796 VDDA.n795 57.2449
R5640 VDDA.n782 VDDA.n781 57.2449
R5641 VDDA.n841 VDDA.n338 57.2449
R5642 VDDA.n795 VDDA.n358 57.2449
R5643 VDDA.n165 VDDA.n53 54.4005
R5644 VDDA.n93 VDDA.n44 54.4005
R5645 VDDA.n210 VDDA.n35 54.4005
R5646 VDDA.n259 VDDA.n17 54.4005
R5647 VDDA.n89 VDDA.n1 54.4005
R5648 VDDA.n96 VDDA.n62 54.4005
R5649 VDDA.n992 VDDA.n307 54.4005
R5650 VDDA.n309 VDDA.n307 54.4005
R5651 VDDA.n309 VDDA.n308 54.4005
R5652 VDDA.n992 VDDA.n308 54.4005
R5653 VDDA.n85 VDDA.n84 53.3664
R5654 VDDA.n79 VDDA.n77 53.3664
R5655 VDDA.n115 VDDA.n109 53.3664
R5656 VDDA.n117 VDDA.n73 53.3664
R5657 VDDA.n107 VDDA.n98 53.3664
R5658 VDDA.n100 VDDA.n88 53.3664
R5659 VDDA.n921 VDDA.n920 53.3664
R5660 VDDA.n942 VDDA.n936 53.3664
R5661 VDDA.n964 VDDA.n963 53.3664
R5662 VDDA.n815 VDDA.n814 53.3664
R5663 VDDA.n809 VDDA.n808 53.3664
R5664 VDDA.n901 VDDA.n326 53.3664
R5665 VDDA.n899 VDDA.n898 53.3664
R5666 VDDA.n973 VDDA.n318 53.3664
R5667 VDDA.n947 VDDA.n937 53.3664
R5668 VDDA.n927 VDDA.n926 53.3664
R5669 VDDA.n823 VDDA.n817 53.3664
R5670 VDDA.n819 VDDA.n807 53.3664
R5671 VDDA.n893 VDDA.n328 53.3664
R5672 VDDA.n889 VDDA.n327 53.3664
R5673 VDDA.n915 VDDA.n320 53.3664
R5674 VDDA.n911 VDDA.n319 53.3664
R5675 VDDA.n971 VDDA.n965 53.3664
R5676 VDDA.n967 VDDA.n917 53.3664
R5677 VDDA.n958 VDDA.n948 53.3664
R5678 VDDA.n953 VDDA.n918 53.3664
R5679 VDDA.n934 VDDA.n928 53.3664
R5680 VDDA.n930 VDDA.n919 53.3664
R5681 VDDA.n830 VDDA.n805 53.3664
R5682 VDDA.n826 VDDA.n805 53.3664
R5683 VDDA.n582 VDDA.n573 53.3664
R5684 VDDA.n588 VDDA.n575 53.3664
R5685 VDDA.n573 VDDA.n549 53.3664
R5686 VDDA.n553 VDDA.n550 53.3664
R5687 VDDA.n565 VDDA.n551 53.3664
R5688 VDDA.n566 VDDA.n550 53.3664
R5689 VDDA.n558 VDDA.n551 53.3664
R5690 VDDA.n473 VDDA.t152 50.7639
R5691 VDDA.t308 VDDA.n450 49.2505
R5692 VDDA.n450 VDDA.t1 49.2505
R5693 VDDA.n443 VDDA.t230 49.2505
R5694 VDDA.n443 VDDA.t36 49.2505
R5695 VDDA.n474 VDDA.t272 49.2505
R5696 VDDA.n474 VDDA.t233 49.2505
R5697 VDDA.n469 VDDA.t259 49.2505
R5698 VDDA.n469 VDDA.t278 49.2505
R5699 VDDA.n447 VDDA.t255 49.2505
R5700 VDDA.n447 VDDA.t67 49.2505
R5701 VDDA.n449 VDDA.t218 49.2505
R5702 VDDA.n449 VDDA.t323 49.2505
R5703 VDDA.n363 VDDA.t423 49.1638
R5704 VDDA.n365 VDDA.t429 48.5162
R5705 VDDA.n1007 VDDA.n1006 47.7005
R5706 VDDA.n837 VDDA.n833 45.3071
R5707 VDDA.n355 VDDA.n347 45.3071
R5708 VDDA.n356 VDDA.n348 45.3071
R5709 VDDA.n842 VDDA.n834 45.3071
R5710 VDDA.n778 VDDA.n774 45.3071
R5711 VDDA.n780 VDDA.n773 45.3071
R5712 VDDA.n802 VDDA.n349 45.3071
R5713 VDDA.n797 VDDA.n346 45.3071
R5714 VDDA.n857 VDDA.n853 45.3071
R5715 VDDA.n859 VDDA.n345 45.3071
R5716 VDDA.n851 VDDA.n843 45.3071
R5717 VDDA.n846 VDDA.n804 45.3071
R5718 VDDA.n483 VDDA.n453 45.3071
R5719 VDDA.n489 VDDA.n480 45.3071
R5720 VDDA.n456 VDDA.n454 45.3071
R5721 VDDA.n461 VDDA.n455 45.3071
R5722 VDDA.n462 VDDA.n454 45.3071
R5723 VDDA.n751 VDDA.n668 45.3071
R5724 VDDA.n673 VDDA.n667 45.3071
R5725 VDDA.n759 VDDA.n666 45.3071
R5726 VDDA.n757 VDDA.n756 45.3071
R5727 VDDA.n716 VDDA.n715 45.3071
R5728 VDDA.n715 VDDA.n712 45.3071
R5729 VDDA.n502 VDDA.n444 41.6005
R5730 VDDA.t223 VDDA.t266 39.886
R5731 VDDA.n496 VDDA.n445 39.4988
R5732 VDDA.n406 VDDA.t244 39.4005
R5733 VDDA.n406 VDDA.t88 39.4005
R5734 VDDA.n404 VDDA.t40 39.4005
R5735 VDDA.n404 VDDA.t93 39.4005
R5736 VDDA.n402 VDDA.t198 39.4005
R5737 VDDA.n402 VDDA.t80 39.4005
R5738 VDDA.n400 VDDA.t339 39.4005
R5739 VDDA.n400 VDDA.t200 39.4005
R5740 VDDA.n398 VDDA.t179 39.4005
R5741 VDDA.n398 VDDA.t97 39.4005
R5742 VDDA.n396 VDDA.t119 39.4005
R5743 VDDA.n396 VDDA.t370 39.4005
R5744 VDDA.n394 VDDA.t10 39.4005
R5745 VDDA.n394 VDDA.t405 39.4005
R5746 VDDA.n392 VDDA.t242 39.4005
R5747 VDDA.n392 VDDA.t8 39.4005
R5748 VDDA.n388 VDDA.t121 39.4005
R5749 VDDA.n388 VDDA.t228 39.4005
R5750 VDDA.n386 VDDA.t214 39.4005
R5751 VDDA.n386 VDDA.t60 39.4005
R5752 VDDA.n384 VDDA.t363 39.4005
R5753 VDDA.n384 VDDA.t240 39.4005
R5754 VDDA.n382 VDDA.t403 39.4005
R5755 VDDA.n382 VDDA.t349 39.4005
R5756 VDDA.n380 VDDA.t359 39.4005
R5757 VDDA.n380 VDDA.t65 39.4005
R5758 VDDA.n378 VDDA.t353 39.4005
R5759 VDDA.n378 VDDA.t355 39.4005
R5760 VDDA.n376 VDDA.t250 39.4005
R5761 VDDA.n376 VDDA.t351 39.4005
R5762 VDDA.n374 VDDA.t357 39.4005
R5763 VDDA.n374 VDDA.t181 39.4005
R5764 VDDA.n372 VDDA.t347 39.4005
R5765 VDDA.n372 VDDA.t361 39.4005
R5766 VDDA.n368 VDDA.t50 39.4005
R5767 VDDA.n368 VDDA.t345 39.4005
R5768 VDDA.n639 VDDA.t407 39.4005
R5769 VDDA.n639 VDDA.t149 39.4005
R5770 VDDA.n637 VDDA.t169 39.4005
R5771 VDDA.n637 VDDA.t157 39.4005
R5772 VDDA.n635 VDDA.t382 39.4005
R5773 VDDA.n635 VDDA.t147 39.4005
R5774 VDDA.n633 VDDA.t384 39.4005
R5775 VDDA.n633 VDDA.t175 39.4005
R5776 VDDA.n628 VDDA.t195 39.4005
R5777 VDDA.n628 VDDA.t396 39.4005
R5778 VDDA.n626 VDDA.t193 39.4005
R5779 VDDA.n626 VDDA.t380 39.4005
R5780 VDDA.n624 VDDA.t173 39.4005
R5781 VDDA.n624 VDDA.t378 39.4005
R5782 VDDA.n622 VDDA.t411 39.4005
R5783 VDDA.n622 VDDA.t171 39.4005
R5784 VDDA.n620 VDDA.t413 39.4005
R5785 VDDA.n620 VDDA.t398 39.4005
R5786 VDDA.n615 VDDA.t155 39.4005
R5787 VDDA.n615 VDDA.t409 39.4005
R5788 VDDA.n768 VDDA.n767 38.1005
R5789 VDDA.n478 VDDA.t294 36.26
R5790 VDDA.t373 VDDA.t232 32.6341
R5791 VDDA.t215 VDDA.t264 32.6341
R5792 VDDA.n750 VDDA.n669 32.2291
R5793 VDDA.n120 VDDA.n70 32.0005
R5794 VDDA.n124 VDDA.n70 32.0005
R5795 VDDA.n125 VDDA.n124 32.0005
R5796 VDDA.n126 VDDA.n125 32.0005
R5797 VDDA.n132 VDDA.n131 32.0005
R5798 VDDA.n135 VDDA.n132 32.0005
R5799 VDDA.n139 VDDA.n64 32.0005
R5800 VDDA.n140 VDDA.n139 32.0005
R5801 VDDA.n141 VDDA.n140 32.0005
R5802 VDDA.n145 VDDA.n144 32.0005
R5803 VDDA.n146 VDDA.n145 32.0005
R5804 VDDA.n146 VDDA.n60 32.0005
R5805 VDDA.n150 VDDA.n60 32.0005
R5806 VDDA.n151 VDDA.n150 32.0005
R5807 VDDA.n153 VDDA.n57 32.0005
R5808 VDDA.n157 VDDA.n57 32.0005
R5809 VDDA.n160 VDDA.n159 32.0005
R5810 VDDA.n160 VDDA.n54 32.0005
R5811 VDDA.n164 VDDA.n54 32.0005
R5812 VDDA.n167 VDDA.n166 32.0005
R5813 VDDA.n167 VDDA.n51 32.0005
R5814 VDDA.n171 VDDA.n51 32.0005
R5815 VDDA.n172 VDDA.n171 32.0005
R5816 VDDA.n173 VDDA.n172 32.0005
R5817 VDDA.n177 VDDA.n176 32.0005
R5818 VDDA.n180 VDDA.n177 32.0005
R5819 VDDA.n184 VDDA.n46 32.0005
R5820 VDDA.n185 VDDA.n184 32.0005
R5821 VDDA.n186 VDDA.n185 32.0005
R5822 VDDA.n190 VDDA.n189 32.0005
R5823 VDDA.n191 VDDA.n190 32.0005
R5824 VDDA.n191 VDDA.n42 32.0005
R5825 VDDA.n195 VDDA.n42 32.0005
R5826 VDDA.n196 VDDA.n195 32.0005
R5827 VDDA.n198 VDDA.n39 32.0005
R5828 VDDA.n202 VDDA.n39 32.0005
R5829 VDDA.n205 VDDA.n204 32.0005
R5830 VDDA.n205 VDDA.n36 32.0005
R5831 VDDA.n209 VDDA.n36 32.0005
R5832 VDDA.n212 VDDA.n211 32.0005
R5833 VDDA.n212 VDDA.n33 32.0005
R5834 VDDA.n216 VDDA.n33 32.0005
R5835 VDDA.n217 VDDA.n216 32.0005
R5836 VDDA.n220 VDDA.n217 32.0005
R5837 VDDA.n224 VDDA.n31 32.0005
R5838 VDDA.n225 VDDA.n224 32.0005
R5839 VDDA.n226 VDDA.n225 32.0005
R5840 VDDA.n230 VDDA.n229 32.0005
R5841 VDDA.n231 VDDA.n230 32.0005
R5842 VDDA.n231 VDDA.n26 32.0005
R5843 VDDA.n235 VDDA.n26 32.0005
R5844 VDDA.n239 VDDA.n237 32.0005
R5845 VDDA.n243 VDDA.n24 32.0005
R5846 VDDA.n244 VDDA.n243 32.0005
R5847 VDDA.n246 VDDA.n21 32.0005
R5848 VDDA.n250 VDDA.n21 32.0005
R5849 VDDA.n251 VDDA.n250 32.0005
R5850 VDDA.n253 VDDA.n18 32.0005
R5851 VDDA.n257 VDDA.n18 32.0005
R5852 VDDA.n258 VDDA.n257 32.0005
R5853 VDDA.n260 VDDA.n15 32.0005
R5854 VDDA.n264 VDDA.n15 32.0005
R5855 VDDA.n265 VDDA.n264 32.0005
R5856 VDDA.n266 VDDA.n265 32.0005
R5857 VDDA.n266 VDDA.n13 32.0005
R5858 VDDA.n270 VDDA.n13 32.0005
R5859 VDDA.n273 VDDA.n272 32.0005
R5860 VDDA.n273 VDDA.n10 32.0005
R5861 VDDA.n277 VDDA.n10 32.0005
R5862 VDDA.n278 VDDA.n277 32.0005
R5863 VDDA.n279 VDDA.n278 32.0005
R5864 VDDA.n283 VDDA.n282 32.0005
R5865 VDDA.n284 VDDA.n283 32.0005
R5866 VDDA.n284 VDDA.n5 32.0005
R5867 VDDA.n288 VDDA.n5 32.0005
R5868 VDDA.n289 VDDA.n288 32.0005
R5869 VDDA.n292 VDDA.n289 32.0005
R5870 VDDA.n296 VDDA.n3 32.0005
R5871 VDDA.n297 VDDA.n296 32.0005
R5872 VDDA.n298 VDDA.n297 32.0005
R5873 VDDA.n783 VDDA.n362 32.0005
R5874 VDDA.n787 VDDA.n362 32.0005
R5875 VDDA.n788 VDDA.n787 32.0005
R5876 VDDA.n789 VDDA.n788 32.0005
R5877 VDDA.n789 VDDA.n359 32.0005
R5878 VDDA.n795 VDDA.n359 32.0005
R5879 VDDA.n795 VDDA.n360 32.0005
R5880 VDDA.n360 VDDA.n342 32.0005
R5881 VDDA.n862 VDDA.n342 32.0005
R5882 VDDA.n866 VDDA.n340 32.0005
R5883 VDDA.n867 VDDA.n866 32.0005
R5884 VDDA.n868 VDDA.n867 32.0005
R5885 VDDA.n872 VDDA.n871 32.0005
R5886 VDDA.n873 VDDA.n872 32.0005
R5887 VDDA.n873 VDDA.n336 32.0005
R5888 VDDA.n877 VDDA.n336 32.0005
R5889 VDDA.n881 VDDA.n880 32.0005
R5890 VDDA.n881 VDDA.n330 32.0005
R5891 VDDA.n885 VDDA.n332 32.0005
R5892 VDDA.n908 VDDA.n322 32.0005
R5893 VDDA.n976 VDDA.n315 32.0005
R5894 VDDA.n980 VDDA.n313 32.0005
R5895 VDDA.n981 VDDA.n980 32.0005
R5896 VDDA.n982 VDDA.n981 32.0005
R5897 VDDA.n982 VDDA.n311 32.0005
R5898 VDDA.n986 VDDA.n311 32.0005
R5899 VDDA.n987 VDDA.n986 32.0005
R5900 VDDA.n988 VDDA.n987 32.0005
R5901 VDDA.n994 VDDA.n993 32.0005
R5902 VDDA.n994 VDDA.n305 32.0005
R5903 VDDA.n998 VDDA.n305 32.0005
R5904 VDDA.n999 VDDA.n998 32.0005
R5905 VDDA.n1000 VDDA.n999 32.0005
R5906 VDDA.n1000 VDDA.n303 32.0005
R5907 VDDA.n1004 VDDA.n303 32.0005
R5908 VDDA.n500 VDDA.n445 32.0005
R5909 VDDA.n501 VDDA.n500 32.0005
R5910 VDDA.n503 VDDA.n440 32.0005
R5911 VDDA.n508 VDDA.n440 32.0005
R5912 VDDA.n509 VDDA.n508 32.0005
R5913 VDDA.n510 VDDA.n509 32.0005
R5914 VDDA.n510 VDDA.n437 32.0005
R5915 VDDA.n515 VDDA.n437 32.0005
R5916 VDDA.n516 VDDA.n515 32.0005
R5917 VDDA.n517 VDDA.n516 32.0005
R5918 VDDA.n517 VDDA.n434 32.0005
R5919 VDDA.n522 VDDA.n434 32.0005
R5920 VDDA.n523 VDDA.n522 32.0005
R5921 VDDA.n524 VDDA.n523 32.0005
R5922 VDDA.n524 VDDA.n431 32.0005
R5923 VDDA.n529 VDDA.n431 32.0005
R5924 VDDA.n530 VDDA.n529 32.0005
R5925 VDDA.n530 VDDA.n429 32.0005
R5926 VDDA.n534 VDDA.n429 32.0005
R5927 VDDA.n535 VDDA.n534 32.0005
R5928 VDDA.n763 VDDA.n661 32.0005
R5929 VDDA.n767 VDDA.n661 32.0005
R5930 VDDA.n687 VDDA.n686 32.0005
R5931 VDDA.n686 VDDA.n685 32.0005
R5932 VDDA.n693 VDDA.n675 32.0005
R5933 VDDA.n693 VDDA.n692 32.0005
R5934 VDDA.n692 VDDA.n691 32.0005
R5935 VDDA.n742 VDDA.n697 32.0005
R5936 VDDA.n737 VDDA.n736 32.0005
R5937 VDDA.n730 VDDA.n729 32.0005
R5938 VDDA.n730 VDDA.n701 32.0005
R5939 VDDA.n734 VDDA.n701 32.0005
R5940 VDDA.n723 VDDA.n722 32.0005
R5941 VDDA.n723 VDDA.n704 32.0005
R5942 VDDA.n727 VDDA.n704 32.0005
R5943 VDDA.n493 VDDA.n492 30.754
R5944 VDDA.n472 VDDA.n471 30.754
R5945 VDDA.n80 VDDA.n71 30.2632
R5946 VDDA.n477 VDDA.n476 30.186
R5947 VDDA.n452 VDDA.n451 30.186
R5948 VDDA.n131 VDDA.n67 28.8005
R5949 VDDA.n144 VDDA.n62 28.8005
R5950 VDDA.n153 VDDA.n152 28.8005
R5951 VDDA.n166 VDDA.n165 28.8005
R5952 VDDA.n176 VDDA.n49 28.8005
R5953 VDDA.n189 VDDA.n44 28.8005
R5954 VDDA.n198 VDDA.n197 28.8005
R5955 VDDA.n211 VDDA.n210 28.8005
R5956 VDDA.n246 VDDA.n245 28.8005
R5957 VDDA.n271 VDDA.n270 28.8005
R5958 VDDA.n862 VDDA.n861 28.8005
R5959 VDDA.n762 VDDA.n663 28.8005
R5960 VDDA.n687 VDDA.n678 28.8005
R5961 VDDA.n743 VDDA.n742 28.8005
R5962 VDDA.n259 VDDA.n258 25.6005
R5963 VDDA.n783 VDDA.n782 25.6005
R5964 VDDA.n868 VDDA.n338 25.6005
R5965 VDDA.n880 VDDA.n879 25.6005
R5966 VDDA.n904 VDDA.n903 25.6005
R5967 VDDA.n909 VDDA.n315 25.6005
R5968 VDDA.n976 VDDA.n975 25.6005
R5969 VDDA.n991 VDDA.n309 25.6005
R5970 VDDA.n992 VDDA.n991 25.6005
R5971 VDDA.n1006 VDDA.n1005 25.6005
R5972 VDDA.n502 VDDA.n501 25.6005
R5973 VDDA VDDA.n535 25.6005
R5974 VDDA.t17 VDDA.t258 25.3822
R5975 VDDA.t277 VDDA.t70 25.3822
R5976 VDDA.n119 VDDA.n118 24.991
R5977 VDDA.n101 VDDA.n68 24.991
R5978 VDDA.n1007 VDDA.n300 24.9182
R5979 VDDA.n844 VDDA.t113 24.6255
R5980 VDDA.n344 VDDA.t106 24.6255
R5981 VDDA.n350 VDDA.t4 24.6255
R5982 VDDA.n772 VDDA.t46 24.6255
R5983 VDDA.n835 VDDA.t69 24.6255
R5984 VDDA.n351 VDDA.t416 24.6255
R5985 VDDA.n680 VDDA.t84 24.6255
R5986 VDDA.n680 VDDA.t330 24.6255
R5987 VDDA.n677 VDDA.t101 24.6255
R5988 VDDA.n677 VDDA.t42 24.6255
R5989 VDDA.t327 VDDA.n744 24.6255
R5990 VDDA.n744 VDDA.t392 24.6255
R5991 VDDA.n700 VDDA.t22 24.6255
R5992 VDDA.n700 VDDA.t298 24.6255
R5993 VDDA.n703 VDDA.t30 24.6255
R5994 VDDA.n703 VDDA.t422 24.6255
R5995 VDDA.n720 VDDA.t320 24.6255
R5996 VDDA.n720 VDDA.t246 24.6255
R5997 VDDA.t320 VDDA.n719 24.6255
R5998 VDDA.n664 VDDA.t331 24.6255
R5999 VDDA.n745 VDDA.t327 24.6255
R6000 VDDA.n749 VDDA.t299 24.6255
R6001 VDDA.n709 VDDA.n706 24.361
R6002 VDDA.n129 VDDA.n128 24.1919
R6003 VDDA.n300 VDDA.n1 23.4989
R6004 VDDA.n592 VDDA.n591 22.8576
R6005 VDDA.n561 VDDA.n538 22.8576
R6006 VDDA.n120 VDDA.n119 22.4005
R6007 VDDA.n126 VDDA.n68 22.4005
R6008 VDDA.n135 VDDA.n134 22.4005
R6009 VDDA.n158 VDDA.n157 22.4005
R6010 VDDA.n180 VDDA.n179 22.4005
R6011 VDDA.n203 VDDA.n202 22.4005
R6012 VDDA.n219 VDDA.n31 22.4005
R6013 VDDA.n226 VDDA.n29 22.4005
R6014 VDDA.n291 VDDA.n3 22.4005
R6015 VDDA.n685 VDDA.n681 22.4005
R6016 VDDA.n736 VDDA.n735 22.4005
R6017 VDDA.n737 VDDA.n669 22.4005
R6018 VDDA.n466 VDDA.n457 22.0449
R6019 VDDA.n481 VDDA.t295 19.7005
R6020 VDDA.n458 VDDA.t286 19.7005
R6021 VDDA.n432 VDDA.t216 19.7005
R6022 VDDA.n432 VDDA.t285 19.7005
R6023 VDDA.n435 VDDA.t224 19.7005
R6024 VDDA.n435 VDDA.t376 19.7005
R6025 VDDA.n438 VDDA.t71 19.7005
R6026 VDDA.n438 VDDA.t153 19.7005
R6027 VDDA.n441 VDDA.t151 19.7005
R6028 VDDA.n441 VDDA.t18 19.7005
R6029 VDDA.t295 VDDA.n446 19.7005
R6030 VDDA.n446 VDDA.t374 19.7005
R6031 VDDA.n237 VDDA.n236 19.2005
R6032 VDDA.n239 VDDA.n238 19.2005
R6033 VDDA.n279 VDDA.n8 19.2005
R6034 VDDA.n332 VDDA.n324 19.2005
R6035 VDDA.t229 VDDA.t150 18.1303
R6036 VDDA.t263 VDDA.t284 18.1303
R6037 VDDA.n762 VDDA.n761 17.6005
R6038 VDDA.n367 VDDA.t85 17.0848
R6039 VDDA.n252 VDDA.n251 16.0005
R6040 VDDA.n253 VDDA.n252 16.0005
R6041 VDDA.n298 VDDA.n1 16.0005
R6042 VDDA.n886 VDDA.n885 16.0005
R6043 VDDA.n494 VDDA.n493 16.0005
R6044 VDDA.n471 VDDA.n470 16.0005
R6045 VDDA.n476 VDDA.n475 16.0005
R6046 VDDA.n451 VDDA.n448 16.0005
R6047 VDDA.n681 VDDA.n663 16.0005
R6048 VDDA.n697 VDDA.n669 16.0005
R6049 VDDA.n735 VDDA.n734 16.0005
R6050 VDDA.n722 VDDA.n721 16.0005
R6051 VDDA.n536 VDDA 15.7005
R6052 VDDA.n761 VDDA.n760 15.6449
R6053 VDDA.n718 VDDA.n709 15.6449
R6054 VDDA.n782 VDDA.n770 13.8989
R6055 VDDA.n546 VDDA.t124 13.1338
R6056 VDDA.n546 VDDA.t140 13.1338
R6057 VDDA.n545 VDDA.t131 13.1338
R6058 VDDA.n545 VDDA.t142 13.1338
R6059 VDDA.n544 VDDA.t418 13.1338
R6060 VDDA.n544 VDDA.t104 13.1338
R6061 VDDA.n543 VDDA.t183 13.1338
R6062 VDDA.n543 VDDA.t368 13.1338
R6063 VDDA.n542 VDDA.t126 13.1338
R6064 VDDA.n542 VDDA.t24 13.1338
R6065 VDDA.n541 VDDA.t32 13.1338
R6066 VDDA.n541 VDDA.t253 13.1338
R6067 VDDA.n540 VDDA.t137 13.1338
R6068 VDDA.n540 VDDA.t420 13.1338
R6069 VDDA.n539 VDDA.t34 13.1338
R6070 VDDA.n539 VDDA.t133 13.1338
R6071 VDDA.n236 VDDA.n235 12.8005
R6072 VDDA.n238 VDDA.n24 12.8005
R6073 VDDA.n282 VDDA.n8 12.8005
R6074 VDDA.n887 VDDA.n330 12.8005
R6075 VDDA.n904 VDDA.n324 12.8005
R6076 VDDA.n770 VDDA.n769 12.343
R6077 VDDA.n537 VDDA.n536 11.6166
R6078 VDDA.n769 VDDA.n768 11.579
R6079 VDDA.n832 VDDA.t247 11.4924
R6080 VDDA.t162 VDDA.n824 11.4924
R6081 VDDA.n816 VDDA.t114 11.4924
R6082 VDDA.n894 VDDA.t385 11.4924
R6083 VDDA.n900 VDDA.t204 11.4924
R6084 VDDA.n593 VDDA.n592 11.0575
R6085 VDDA.t28 VDDA.t375 10.8784
R6086 VDDA.n601 VDDA.n538 10.87
R6087 VDDA.n129 VDDA.n67 10.7016
R6088 VDDA.n660 VDDA.n659 10.508
R6089 VDDA.n457 VDDA.n430 9.613
R6090 VDDA.n134 VDDA.n64 9.6005
R6091 VDDA.n159 VDDA.n158 9.6005
R6092 VDDA.n179 VDDA.n46 9.6005
R6093 VDDA.n204 VDDA.n203 9.6005
R6094 VDDA.n220 VDDA.n219 9.6005
R6095 VDDA.n229 VDDA.n29 9.6005
R6096 VDDA.n292 VDDA.n291 9.6005
R6097 VDDA.n763 VDDA.n762 9.6005
R6098 VDDA.n743 VDDA.n675 9.6005
R6099 VDDA.n691 VDDA.n678 9.6005
R6100 VDDA.n414 VDDA.n390 9.50883
R6101 VDDA.n424 VDDA.n370 9.50883
R6102 VDDA.n570 VDDA.n569 9.50883
R6103 VDDA.n562 VDDA.n561 9.50883
R6104 VDDA.n587 VDDA.n576 9.50883
R6105 VDDA.n591 VDDA.n548 9.50883
R6106 VDDA.n611 VDDA.n603 9.50883
R6107 VDDA.n121 VDDA.n120 9.3005
R6108 VDDA.n122 VDDA.n70 9.3005
R6109 VDDA.n124 VDDA.n123 9.3005
R6110 VDDA.n125 VDDA.n69 9.3005
R6111 VDDA.n127 VDDA.n126 9.3005
R6112 VDDA.n131 VDDA.n130 9.3005
R6113 VDDA.n132 VDDA.n65 9.3005
R6114 VDDA.n136 VDDA.n135 9.3005
R6115 VDDA.n137 VDDA.n64 9.3005
R6116 VDDA.n139 VDDA.n138 9.3005
R6117 VDDA.n140 VDDA.n63 9.3005
R6118 VDDA.n142 VDDA.n141 9.3005
R6119 VDDA.n144 VDDA.n143 9.3005
R6120 VDDA.n145 VDDA.n61 9.3005
R6121 VDDA.n147 VDDA.n146 9.3005
R6122 VDDA.n148 VDDA.n60 9.3005
R6123 VDDA.n150 VDDA.n149 9.3005
R6124 VDDA.n151 VDDA.n58 9.3005
R6125 VDDA.n154 VDDA.n153 9.3005
R6126 VDDA.n155 VDDA.n57 9.3005
R6127 VDDA.n157 VDDA.n156 9.3005
R6128 VDDA.n159 VDDA.n55 9.3005
R6129 VDDA.n161 VDDA.n160 9.3005
R6130 VDDA.n162 VDDA.n54 9.3005
R6131 VDDA.n164 VDDA.n163 9.3005
R6132 VDDA.n166 VDDA.n52 9.3005
R6133 VDDA.n168 VDDA.n167 9.3005
R6134 VDDA.n169 VDDA.n51 9.3005
R6135 VDDA.n171 VDDA.n170 9.3005
R6136 VDDA.n172 VDDA.n50 9.3005
R6137 VDDA.n174 VDDA.n173 9.3005
R6138 VDDA.n176 VDDA.n175 9.3005
R6139 VDDA.n177 VDDA.n47 9.3005
R6140 VDDA.n181 VDDA.n180 9.3005
R6141 VDDA.n182 VDDA.n46 9.3005
R6142 VDDA.n184 VDDA.n183 9.3005
R6143 VDDA.n185 VDDA.n45 9.3005
R6144 VDDA.n187 VDDA.n186 9.3005
R6145 VDDA.n189 VDDA.n188 9.3005
R6146 VDDA.n190 VDDA.n43 9.3005
R6147 VDDA.n192 VDDA.n191 9.3005
R6148 VDDA.n193 VDDA.n42 9.3005
R6149 VDDA.n195 VDDA.n194 9.3005
R6150 VDDA.n196 VDDA.n40 9.3005
R6151 VDDA.n199 VDDA.n198 9.3005
R6152 VDDA.n200 VDDA.n39 9.3005
R6153 VDDA.n202 VDDA.n201 9.3005
R6154 VDDA.n204 VDDA.n37 9.3005
R6155 VDDA.n206 VDDA.n205 9.3005
R6156 VDDA.n207 VDDA.n36 9.3005
R6157 VDDA.n209 VDDA.n208 9.3005
R6158 VDDA.n211 VDDA.n34 9.3005
R6159 VDDA.n213 VDDA.n212 9.3005
R6160 VDDA.n214 VDDA.n33 9.3005
R6161 VDDA.n216 VDDA.n215 9.3005
R6162 VDDA.n217 VDDA.n32 9.3005
R6163 VDDA.n221 VDDA.n220 9.3005
R6164 VDDA.n222 VDDA.n31 9.3005
R6165 VDDA.n224 VDDA.n223 9.3005
R6166 VDDA.n225 VDDA.n30 9.3005
R6167 VDDA.n227 VDDA.n226 9.3005
R6168 VDDA.n229 VDDA.n228 9.3005
R6169 VDDA.n230 VDDA.n27 9.3005
R6170 VDDA.n232 VDDA.n231 9.3005
R6171 VDDA.n233 VDDA.n26 9.3005
R6172 VDDA.n235 VDDA.n234 9.3005
R6173 VDDA.n237 VDDA.n25 9.3005
R6174 VDDA.n240 VDDA.n239 9.3005
R6175 VDDA.n241 VDDA.n24 9.3005
R6176 VDDA.n243 VDDA.n242 9.3005
R6177 VDDA.n244 VDDA.n22 9.3005
R6178 VDDA.n247 VDDA.n246 9.3005
R6179 VDDA.n248 VDDA.n21 9.3005
R6180 VDDA.n250 VDDA.n249 9.3005
R6181 VDDA.n251 VDDA.n19 9.3005
R6182 VDDA.n254 VDDA.n253 9.3005
R6183 VDDA.n255 VDDA.n18 9.3005
R6184 VDDA.n257 VDDA.n256 9.3005
R6185 VDDA.n258 VDDA.n16 9.3005
R6186 VDDA.n261 VDDA.n260 9.3005
R6187 VDDA.n262 VDDA.n15 9.3005
R6188 VDDA.n264 VDDA.n263 9.3005
R6189 VDDA.n265 VDDA.n14 9.3005
R6190 VDDA.n267 VDDA.n266 9.3005
R6191 VDDA.n268 VDDA.n13 9.3005
R6192 VDDA.n270 VDDA.n269 9.3005
R6193 VDDA.n272 VDDA.n11 9.3005
R6194 VDDA.n274 VDDA.n273 9.3005
R6195 VDDA.n275 VDDA.n10 9.3005
R6196 VDDA.n277 VDDA.n276 9.3005
R6197 VDDA.n278 VDDA.n9 9.3005
R6198 VDDA.n280 VDDA.n279 9.3005
R6199 VDDA.n282 VDDA.n281 9.3005
R6200 VDDA.n283 VDDA.n6 9.3005
R6201 VDDA.n285 VDDA.n284 9.3005
R6202 VDDA.n286 VDDA.n5 9.3005
R6203 VDDA.n288 VDDA.n287 9.3005
R6204 VDDA.n289 VDDA.n4 9.3005
R6205 VDDA.n293 VDDA.n292 9.3005
R6206 VDDA.n294 VDDA.n3 9.3005
R6207 VDDA.n296 VDDA.n295 9.3005
R6208 VDDA.n297 VDDA.n2 9.3005
R6209 VDDA.n299 VDDA.n298 9.3005
R6210 VDDA.n414 VDDA.n413 9.3005
R6211 VDDA.n424 VDDA.n423 9.3005
R6212 VDDA.n580 VDDA.n548 9.3005
R6213 VDDA.n583 VDDA.n579 9.3005
R6214 VDDA.n584 VDDA.n578 9.3005
R6215 VDDA.n577 VDDA.n576 9.3005
R6216 VDDA.n562 VDDA.n559 9.3005
R6217 VDDA.n564 VDDA.n563 9.3005
R6218 VDDA.n567 VDDA.n555 9.3005
R6219 VDDA.n569 VDDA.n568 9.3005
R6220 VDDA.n611 VDDA.n610 9.3005
R6221 VDDA.n535 VDDA.n428 9.3005
R6222 VDDA.n534 VDDA.n533 9.3005
R6223 VDDA.n532 VDDA.n429 9.3005
R6224 VDDA.n531 VDDA.n530 9.3005
R6225 VDDA.n529 VDDA.n528 9.3005
R6226 VDDA.n527 VDDA.n431 9.3005
R6227 VDDA.n525 VDDA.n524 9.3005
R6228 VDDA.n523 VDDA.n433 9.3005
R6229 VDDA.n522 VDDA.n521 9.3005
R6230 VDDA.n520 VDDA.n434 9.3005
R6231 VDDA.n518 VDDA.n517 9.3005
R6232 VDDA.n516 VDDA.n436 9.3005
R6233 VDDA.n515 VDDA.n514 9.3005
R6234 VDDA.n513 VDDA.n437 9.3005
R6235 VDDA.n511 VDDA.n510 9.3005
R6236 VDDA.n509 VDDA.n439 9.3005
R6237 VDDA.n508 VDDA.n507 9.3005
R6238 VDDA.n506 VDDA.n440 9.3005
R6239 VDDA.n504 VDDA.n503 9.3005
R6240 VDDA.n498 VDDA.n445 9.3005
R6241 VDDA.n500 VDDA.n499 9.3005
R6242 VDDA.n501 VDDA.n442 9.3005
R6243 VDDA.n722 VDDA.n705 9.3005
R6244 VDDA.n724 VDDA.n723 9.3005
R6245 VDDA.n725 VDDA.n704 9.3005
R6246 VDDA.n727 VDDA.n726 9.3005
R6247 VDDA.n729 VDDA.n702 9.3005
R6248 VDDA.n731 VDDA.n730 9.3005
R6249 VDDA.n732 VDDA.n701 9.3005
R6250 VDDA.n734 VDDA.n733 9.3005
R6251 VDDA.n735 VDDA.n699 9.3005
R6252 VDDA.n736 VDDA.n698 9.3005
R6253 VDDA.n738 VDDA.n737 9.3005
R6254 VDDA.n739 VDDA.n669 9.3005
R6255 VDDA.n740 VDDA.n697 9.3005
R6256 VDDA.n742 VDDA.n741 9.3005
R6257 VDDA.n743 VDDA.n696 9.3005
R6258 VDDA.n695 VDDA.n675 9.3005
R6259 VDDA.n694 VDDA.n693 9.3005
R6260 VDDA.n692 VDDA.n676 9.3005
R6261 VDDA.n691 VDDA.n690 9.3005
R6262 VDDA.n689 VDDA.n678 9.3005
R6263 VDDA.n688 VDDA.n687 9.3005
R6264 VDDA.n686 VDDA.n679 9.3005
R6265 VDDA.n685 VDDA.n684 9.3005
R6266 VDDA.n683 VDDA.n681 9.3005
R6267 VDDA.n682 VDDA.n663 9.3005
R6268 VDDA.n762 VDDA.n662 9.3005
R6269 VDDA.n764 VDDA.n763 9.3005
R6270 VDDA.n765 VDDA.n661 9.3005
R6271 VDDA.n767 VDDA.n766 9.3005
R6272 VDDA.n1006 VDDA.n0 9.3005
R6273 VDDA.n784 VDDA.n783 9.3005
R6274 VDDA.n785 VDDA.n362 9.3005
R6275 VDDA.n787 VDDA.n786 9.3005
R6276 VDDA.n788 VDDA.n361 9.3005
R6277 VDDA.n790 VDDA.n789 9.3005
R6278 VDDA.n791 VDDA.n359 9.3005
R6279 VDDA.n795 VDDA.n794 9.3005
R6280 VDDA.n793 VDDA.n360 9.3005
R6281 VDDA.n792 VDDA.n342 9.3005
R6282 VDDA.n863 VDDA.n862 9.3005
R6283 VDDA.n864 VDDA.n340 9.3005
R6284 VDDA.n866 VDDA.n865 9.3005
R6285 VDDA.n867 VDDA.n339 9.3005
R6286 VDDA.n869 VDDA.n868 9.3005
R6287 VDDA.n871 VDDA.n870 9.3005
R6288 VDDA.n872 VDDA.n337 9.3005
R6289 VDDA.n874 VDDA.n873 9.3005
R6290 VDDA.n875 VDDA.n336 9.3005
R6291 VDDA.n877 VDDA.n876 9.3005
R6292 VDDA.n880 VDDA.n333 9.3005
R6293 VDDA.n882 VDDA.n881 9.3005
R6294 VDDA.n883 VDDA.n330 9.3005
R6295 VDDA.n885 VDDA.n884 9.3005
R6296 VDDA.n332 VDDA.n323 9.3005
R6297 VDDA.n905 VDDA.n904 9.3005
R6298 VDDA.n906 VDDA.n322 9.3005
R6299 VDDA.n908 VDDA.n907 9.3005
R6300 VDDA.n315 VDDA.n314 9.3005
R6301 VDDA.n977 VDDA.n976 9.3005
R6302 VDDA.n978 VDDA.n313 9.3005
R6303 VDDA.n980 VDDA.n979 9.3005
R6304 VDDA.n981 VDDA.n312 9.3005
R6305 VDDA.n983 VDDA.n982 9.3005
R6306 VDDA.n984 VDDA.n311 9.3005
R6307 VDDA.n986 VDDA.n985 9.3005
R6308 VDDA.n987 VDDA.n310 9.3005
R6309 VDDA.n989 VDDA.n988 9.3005
R6310 VDDA.n991 VDDA.n990 9.3005
R6311 VDDA.n993 VDDA.n306 9.3005
R6312 VDDA.n995 VDDA.n994 9.3005
R6313 VDDA.n996 VDDA.n305 9.3005
R6314 VDDA.n998 VDDA.n997 9.3005
R6315 VDDA.n999 VDDA.n304 9.3005
R6316 VDDA.n1001 VDDA.n1000 9.3005
R6317 VDDA.n1002 VDDA.n303 9.3005
R6318 VDDA.n1004 VDDA.n1003 9.3005
R6319 VDDA.n112 VDDA.n111 9.14336
R6320 VDDA.n104 VDDA.n103 9.14336
R6321 VDDA.n931 VDDA.n929 9.14336
R6322 VDDA.n968 VDDA.n966 9.14336
R6323 VDDA.n912 VDDA.n321 9.14336
R6324 VDDA.n890 VDDA.n329 9.14336
R6325 VDDA.n820 VDDA.n818 9.14336
R6326 VDDA.n925 VDDA.n924 9.14336
R6327 VDDA.n962 VDDA.n961 9.14336
R6328 VDDA.n897 VDDA.n896 9.14336
R6329 VDDA.n813 VDDA.n812 9.14336
R6330 VDDA.n829 VDDA.n828 9.14336
R6331 VDDA.n584 VDDA.n577 9.14336
R6332 VDDA.n584 VDDA.n583 9.14336
R6333 VDDA.n583 VDDA.n580 9.14336
R6334 VDDA.n568 VDDA.n567 9.14336
R6335 VDDA.n567 VDDA.n564 9.14336
R6336 VDDA.n564 VDDA.n559 9.14336
R6337 VDDA.t109 VDDA.t160 7.66179
R6338 VDDA.n491 VDDA.n490 7.25241
R6339 VDDA.n850 VDDA.n849 7.11161
R6340 VDDA.n847 VDDA.n845 7.11161
R6341 VDDA.n856 VDDA.n855 7.11161
R6342 VDDA.n860 VDDA.n343 7.11161
R6343 VDDA.n801 VDDA.n800 7.11161
R6344 VDDA.n798 VDDA.n796 7.11161
R6345 VDDA.n777 VDDA.n776 7.11161
R6346 VDDA.n781 VDDA.n771 7.11161
R6347 VDDA.n841 VDDA.n840 7.11161
R6348 VDDA.n838 VDDA.n836 7.11161
R6349 VDDA.n358 VDDA.n357 7.11161
R6350 VDDA.n354 VDDA.n353 7.11161
R6351 VDDA.n488 VDDA.n487 7.11161
R6352 VDDA.n485 VDDA.n484 7.11161
R6353 VDDA.n466 VDDA.n465 7.11161
R6354 VDDA.n463 VDDA.n460 7.11161
R6355 VDDA.n760 VDDA.n665 7.11161
R6356 VDDA.n755 VDDA.n753 7.11161
R6357 VDDA.n718 VDDA.n717 7.11161
R6358 VDDA.n711 VDDA.n708 7.11161
R6359 VDDA.n128 VDDA.n68 7.05969
R6360 VDDA.n119 VDDA.n71 7.05957
R6361 VDDA.n721 VDDA.n706 6.54033
R6362 VDDA.n260 VDDA.n259 6.4005
R6363 VDDA.n871 VDDA.n338 6.4005
R6364 VDDA.n903 VDDA.n322 6.4005
R6365 VDDA.n909 VDDA.n908 6.4005
R6366 VDDA.n975 VDDA.n313 6.4005
R6367 VDDA.n988 VDDA.n309 6.4005
R6368 VDDA.n993 VDDA.n992 6.4005
R6369 VDDA.n1005 VDDA.n1004 6.4005
R6370 VDDA.n503 VDDA.n502 6.4005
R6371 VDDA.n83 VDDA.n82 5.81868
R6372 VDDA.n954 VDDA.n950 5.81868
R6373 VDDA.n943 VDDA.n939 5.81868
R6374 VDDA.n106 VDDA.n105 5.33286
R6375 VDDA.n114 VDDA.n113 5.33286
R6376 VDDA.n118 VDDA.n72 5.33286
R6377 VDDA.n102 VDDA.n101 5.33286
R6378 VDDA.n825 VDDA.n334 5.33286
R6379 VDDA.n932 VDDA.n301 5.33286
R6380 VDDA.n969 VDDA.n316 5.33286
R6381 VDDA.n913 VDDA.n910 5.33286
R6382 VDDA.n891 VDDA.n888 5.33286
R6383 VDDA.n821 VDDA.n335 5.33286
R6384 VDDA.n922 VDDA.n302 5.33286
R6385 VDDA.n974 VDDA.n317 5.33286
R6386 VDDA.n902 VDDA.n325 5.33286
R6387 VDDA.n810 VDDA.n331 5.33286
R6388 VDDA.n587 VDDA.n586 5.33286
R6389 VDDA.n591 VDDA.n547 5.33286
R6390 VDDA.n570 VDDA.n554 5.33286
R6391 VDDA.n561 VDDA.n560 5.33286
R6392 VDDA.n641 VDDA.n640 4.84425
R6393 VDDA.n643 VDDA.n642 4.73979
R6394 VDDA.n647 VDDA.n630 4.73979
R6395 VDDA.n653 VDDA.n652 4.73979
R6396 VDDA.n657 VDDA.n617 4.73979
R6397 VDDA.n642 VDDA.n631 4.6505
R6398 VDDA.n647 VDDA.n646 4.6505
R6399 VDDA.n652 VDDA.n618 4.6505
R6400 VDDA.n657 VDDA.n656 4.6505
R6401 VDDA.n632 VDDA.n631 4.54311
R6402 VDDA.n643 VDDA.n632 4.54311
R6403 VDDA.n619 VDDA.n618 4.54311
R6404 VDDA.n653 VDDA.n619 4.54311
R6405 VDDA.n659 VDDA.n658 4.5005
R6406 VDDA.n651 VDDA.n650 4.5005
R6407 VDDA.n649 VDDA.n648 4.5005
R6408 VDDA.n413 VDDA.n412 4.48641
R6409 VDDA.n412 VDDA.n390 4.48641
R6410 VDDA.n423 VDDA.n422 4.48641
R6411 VDDA.n422 VDDA.n370 4.48641
R6412 VDDA.n610 VDDA.n609 4.48641
R6413 VDDA.n609 VDDA.n603 4.48641
R6414 VDDA.n646 VDDA.n645 4.48641
R6415 VDDA.n645 VDDA.n630 4.48641
R6416 VDDA.n656 VDDA.n655 4.48641
R6417 VDDA.n655 VDDA.n617 4.48641
R6418 VDDA.n427 VDDA.n367 4.18096
R6419 VDDA.n614 VDDA.n613 4.07196
R6420 VDDA.n427 VDDA.n426 4.05633
R6421 VDDA.n113 VDDA.n112 3.75335
R6422 VDDA.n111 VDDA.n72 3.75335
R6423 VDDA.n105 VDDA.n104 3.75335
R6424 VDDA.n103 VDDA.n102 3.75335
R6425 VDDA.n933 VDDA.n929 3.75335
R6426 VDDA.n932 VDDA.n931 3.75335
R6427 VDDA.n970 VDDA.n966 3.75335
R6428 VDDA.n969 VDDA.n968 3.75335
R6429 VDDA.n914 VDDA.n321 3.75335
R6430 VDDA.n913 VDDA.n912 3.75335
R6431 VDDA.n892 VDDA.n329 3.75335
R6432 VDDA.n891 VDDA.n890 3.75335
R6433 VDDA.n822 VDDA.n818 3.75335
R6434 VDDA.n821 VDDA.n820 3.75335
R6435 VDDA.n925 VDDA.n922 3.75335
R6436 VDDA.n924 VDDA.n923 3.75335
R6437 VDDA.n961 VDDA.n317 3.75335
R6438 VDDA.n962 VDDA.n960 3.75335
R6439 VDDA.n896 VDDA.n325 3.75335
R6440 VDDA.n897 VDDA.n895 3.75335
R6441 VDDA.n813 VDDA.n810 3.75335
R6442 VDDA.n812 VDDA.n811 3.75335
R6443 VDDA.n829 VDDA.n825 3.75335
R6444 VDDA.n828 VDDA.n827 3.75335
R6445 VDDA.n586 VDDA.n577 3.75335
R6446 VDDA.n580 VDDA.n547 3.75335
R6447 VDDA.n568 VDDA.n554 3.75335
R6448 VDDA.n560 VDDA.n559 3.75335
R6449 VDDA.n849 VDDA.n848 3.53508
R6450 VDDA.n848 VDDA.n847 3.53508
R6451 VDDA.n855 VDDA.n854 3.53508
R6452 VDDA.n854 VDDA.n343 3.53508
R6453 VDDA.n800 VDDA.n799 3.53508
R6454 VDDA.n799 VDDA.n798 3.53508
R6455 VDDA.n776 VDDA.n775 3.53508
R6456 VDDA.n775 VDDA.n771 3.53508
R6457 VDDA.n840 VDDA.n839 3.53508
R6458 VDDA.n839 VDDA.n838 3.53508
R6459 VDDA.n357 VDDA.n352 3.53508
R6460 VDDA.n354 VDDA.n352 3.53508
R6461 VDDA.n487 VDDA.n486 3.53508
R6462 VDDA.n484 VDDA.n482 3.53508
R6463 VDDA.n486 VDDA.n485 3.53508
R6464 VDDA.n465 VDDA.n464 3.53508
R6465 VDDA.n460 VDDA.n459 3.53508
R6466 VDDA.n464 VDDA.n463 3.53508
R6467 VDDA.n754 VDDA.n665 3.53508
R6468 VDDA.n755 VDDA.n754 3.53508
R6469 VDDA.n717 VDDA.n707 3.53508
R6470 VDDA.n711 VDDA.n707 3.53508
R6471 VDDA.n606 VDDA.n605 3.46433
R6472 VDDA.n409 VDDA.n408 3.41464
R6473 VDDA.n419 VDDA.n418 3.41464
R6474 VDDA.n86 VDDA.n76 3.40194
R6475 VDDA.n81 VDDA.n80 3.40194
R6476 VDDA.n957 VDDA.n956 3.40194
R6477 VDDA.n955 VDDA.n951 3.40194
R6478 VDDA.n946 VDDA.n945 3.40194
R6479 VDDA.n944 VDDA.n940 3.40194
R6480 VDDA.n141 VDDA.n62 3.2005
R6481 VDDA.n152 VDDA.n151 3.2005
R6482 VDDA.n165 VDDA.n164 3.2005
R6483 VDDA.n173 VDDA.n49 3.2005
R6484 VDDA.n186 VDDA.n44 3.2005
R6485 VDDA.n197 VDDA.n196 3.2005
R6486 VDDA.n210 VDDA.n209 3.2005
R6487 VDDA.n245 VDDA.n244 3.2005
R6488 VDDA.n272 VDDA.n271 3.2005
R6489 VDDA.n861 VDDA.n340 3.2005
R6490 VDDA.n878 VDDA.n877 3.2005
R6491 VDDA.n879 VDDA.n878 3.2005
R6492 VDDA.n887 VDDA.n886 3.2005
R6493 VDDA.n729 VDDA.n728 3.2005
R6494 VDDA.n728 VDDA.n727 3.2005
R6495 VDDA.n410 VDDA.n409 3.11118
R6496 VDDA.n420 VDDA.n419 3.11118
R6497 VDDA.n409 VDDA.n391 3.04304
R6498 VDDA.n419 VDDA.n371 3.04304
R6499 VDDA.n607 VDDA.n606 2.96855
R6500 VDDA.n606 VDDA.n604 2.90353
R6501 VDDA.n83 VDDA.n76 2.39444
R6502 VDDA.n82 VDDA.n81 2.39444
R6503 VDDA.n956 VDDA.n950 2.39444
R6504 VDDA.n955 VDDA.n954 2.39444
R6505 VDDA.n945 VDDA.n939 2.39444
R6506 VDDA.n944 VDDA.n943 2.39444
R6507 VDDA.n951 VDDA.n307 2.32777
R6508 VDDA.n946 VDDA.n308 2.32777
R6509 VDDA.n671 VDDA.n670 2.27782
R6510 VDDA.n672 VDDA.n671 2.27782
R6511 VDDA.n748 VDDA.n746 2.27782
R6512 VDDA.n674 VDDA.n672 2.27782
R6513 VDDA.n750 VDDA.n670 2.27782
R6514 VDDA.n746 VDDA.n674 2.27782
R6515 VDDA.n605 VDDA.n602 1.94497
R6516 VDDA.n613 VDDA.n612 1.94497
R6517 VDDA.n408 VDDA.n407 1.90331
R6518 VDDA.n416 VDDA.n415 1.77831
R6519 VDDA.n418 VDDA.n417 1.77831
R6520 VDDA.n426 VDDA.n425 1.77831
R6521 VDDA.n367 VDDA.n365 1.05389
R6522 VDDA.n650 VDDA.n649 0.90675
R6523 VDDA.n364 VDDA.n363 0.75233
R6524 VDDA.n706 VDDA.n705 0.703395
R6525 VDDA.n365 VDDA.n364 0.648711
R6526 VDDA.n614 VDDA.n537 0.48024
R6527 VDDA.n769 VDDA.n660 0.4094
R6528 VDDA.n659 VDDA.n616 0.34425
R6529 VDDA.n621 VDDA.n616 0.34425
R6530 VDDA.n623 VDDA.n621 0.34425
R6531 VDDA.n625 VDDA.n623 0.34425
R6532 VDDA.n627 VDDA.n625 0.34425
R6533 VDDA.n650 VDDA.n627 0.34425
R6534 VDDA.n649 VDDA.n629 0.34425
R6535 VDDA.n634 VDDA.n629 0.34425
R6536 VDDA.n636 VDDA.n634 0.34425
R6537 VDDA.n638 VDDA.n636 0.34425
R6538 VDDA.n640 VDDA.n638 0.34425
R6539 VDDA.n417 VDDA.n416 0.333833
R6540 VDDA.n602 VDDA.n601 0.328625
R6541 VDDA.n415 VDDA.n414 0.2505
R6542 VDDA.n425 VDDA.n424 0.2505
R6543 VDDA.n660 VDDA.n614 0.24524
R6544 VDDA.n612 VDDA.n611 0.229667
R6545 VDDA.n613 VDDA.n602 0.229667
R6546 VDDA.n569 VDDA.n555 0.208833
R6547 VDDA.n563 VDDA.n555 0.208833
R6548 VDDA.n563 VDDA.n562 0.208833
R6549 VDDA.n578 VDDA.n576 0.208833
R6550 VDDA.n579 VDDA.n578 0.208833
R6551 VDDA.n579 VDDA.n548 0.208833
R6552 VDDA.n121 VDDA.n71 0.203053
R6553 VDDA.n537 VDDA.n427 0.20294
R6554 VDDA.n128 VDDA.n127 0.202927
R6555 VDDA.n784 VDDA.n770 0.193961
R6556 VDDA.n300 VDDA.n299 0.193958
R6557 VDDA.n130 VDDA.n129 0.193477
R6558 VDDA.n601 VDDA.n600 0.188
R6559 VDDA.n600 VDDA.n599 0.188
R6560 VDDA.n599 VDDA.n598 0.188
R6561 VDDA.n598 VDDA.n597 0.188
R6562 VDDA.n597 VDDA.n596 0.188
R6563 VDDA.n596 VDDA.n595 0.188
R6564 VDDA.n595 VDDA.n594 0.188
R6565 VDDA.n594 VDDA.n593 0.188
R6566 VDDA.n536 VDDA.n428 0.188
R6567 VDDA.n648 VDDA.n647 0.182048
R6568 VDDA.n658 VDDA.n657 0.182048
R6569 VDDA.n642 VDDA.n641 0.182048
R6570 VDDA.n652 VDDA.n651 0.182048
R6571 VDDA.t61 VDDA.t188 0.1603
R6572 VDDA.t135 VDDA.t61 0.1603
R6573 VDDA.t25 VDDA.t135 0.1603
R6574 VDDA.t184 VDDA.t25 0.1603
R6575 VDDA.t94 VDDA.t184 0.1603
R6576 VDDA.t251 VDDA.t94 0.1603
R6577 VDDA.t143 VDDA.t251 0.1603
R6578 VDDA.t129 VDDA.t143 0.1603
R6579 VDDA.t128 VDDA.t127 0.1603
R6580 VDDA.t95 VDDA.t128 0.1603
R6581 VDDA.t138 VDDA.t95 0.1603
R6582 VDDA.t187 VDDA.t138 0.1603
R6583 VDDA.t122 VDDA.t187 0.1603
R6584 VDDA.t62 VDDA.t122 0.1603
R6585 VDDA.t102 VDDA.t62 0.1603
R6586 VDDA.t85 VDDA.t102 0.1603
R6587 VDDA.t86 VDDA.n366 0.159278
R6588 VDDA.n122 VDDA.n121 0.15675
R6589 VDDA.n123 VDDA.n122 0.15675
R6590 VDDA.n123 VDDA.n69 0.15675
R6591 VDDA.n127 VDDA.n69 0.15675
R6592 VDDA.n130 VDDA.n65 0.15675
R6593 VDDA.n136 VDDA.n65 0.15675
R6594 VDDA.n137 VDDA.n136 0.15675
R6595 VDDA.n138 VDDA.n137 0.15675
R6596 VDDA.n138 VDDA.n63 0.15675
R6597 VDDA.n142 VDDA.n63 0.15675
R6598 VDDA.n143 VDDA.n142 0.15675
R6599 VDDA.n143 VDDA.n61 0.15675
R6600 VDDA.n147 VDDA.n61 0.15675
R6601 VDDA.n148 VDDA.n147 0.15675
R6602 VDDA.n149 VDDA.n148 0.15675
R6603 VDDA.n149 VDDA.n58 0.15675
R6604 VDDA.n154 VDDA.n58 0.15675
R6605 VDDA.n155 VDDA.n154 0.15675
R6606 VDDA.n156 VDDA.n155 0.15675
R6607 VDDA.n156 VDDA.n55 0.15675
R6608 VDDA.n161 VDDA.n55 0.15675
R6609 VDDA.n162 VDDA.n161 0.15675
R6610 VDDA.n163 VDDA.n162 0.15675
R6611 VDDA.n163 VDDA.n52 0.15675
R6612 VDDA.n168 VDDA.n52 0.15675
R6613 VDDA.n169 VDDA.n168 0.15675
R6614 VDDA.n170 VDDA.n169 0.15675
R6615 VDDA.n170 VDDA.n50 0.15675
R6616 VDDA.n174 VDDA.n50 0.15675
R6617 VDDA.n175 VDDA.n174 0.15675
R6618 VDDA.n175 VDDA.n47 0.15675
R6619 VDDA.n181 VDDA.n47 0.15675
R6620 VDDA.n182 VDDA.n181 0.15675
R6621 VDDA.n183 VDDA.n182 0.15675
R6622 VDDA.n183 VDDA.n45 0.15675
R6623 VDDA.n187 VDDA.n45 0.15675
R6624 VDDA.n188 VDDA.n187 0.15675
R6625 VDDA.n188 VDDA.n43 0.15675
R6626 VDDA.n192 VDDA.n43 0.15675
R6627 VDDA.n193 VDDA.n192 0.15675
R6628 VDDA.n194 VDDA.n193 0.15675
R6629 VDDA.n194 VDDA.n40 0.15675
R6630 VDDA.n199 VDDA.n40 0.15675
R6631 VDDA.n200 VDDA.n199 0.15675
R6632 VDDA.n201 VDDA.n200 0.15675
R6633 VDDA.n201 VDDA.n37 0.15675
R6634 VDDA.n206 VDDA.n37 0.15675
R6635 VDDA.n207 VDDA.n206 0.15675
R6636 VDDA.n208 VDDA.n207 0.15675
R6637 VDDA.n208 VDDA.n34 0.15675
R6638 VDDA.n213 VDDA.n34 0.15675
R6639 VDDA.n214 VDDA.n213 0.15675
R6640 VDDA.n215 VDDA.n214 0.15675
R6641 VDDA.n215 VDDA.n32 0.15675
R6642 VDDA.n221 VDDA.n32 0.15675
R6643 VDDA.n222 VDDA.n221 0.15675
R6644 VDDA.n223 VDDA.n222 0.15675
R6645 VDDA.n223 VDDA.n30 0.15675
R6646 VDDA.n227 VDDA.n30 0.15675
R6647 VDDA.n228 VDDA.n227 0.15675
R6648 VDDA.n228 VDDA.n27 0.15675
R6649 VDDA.n232 VDDA.n27 0.15675
R6650 VDDA.n233 VDDA.n232 0.15675
R6651 VDDA.n234 VDDA.n233 0.15675
R6652 VDDA.n234 VDDA.n25 0.15675
R6653 VDDA.n240 VDDA.n25 0.15675
R6654 VDDA.n241 VDDA.n240 0.15675
R6655 VDDA.n242 VDDA.n241 0.15675
R6656 VDDA.n242 VDDA.n22 0.15675
R6657 VDDA.n247 VDDA.n22 0.15675
R6658 VDDA.n248 VDDA.n247 0.15675
R6659 VDDA.n249 VDDA.n248 0.15675
R6660 VDDA.n249 VDDA.n19 0.15675
R6661 VDDA.n254 VDDA.n19 0.15675
R6662 VDDA.n255 VDDA.n254 0.15675
R6663 VDDA.n256 VDDA.n255 0.15675
R6664 VDDA.n256 VDDA.n16 0.15675
R6665 VDDA.n261 VDDA.n16 0.15675
R6666 VDDA.n262 VDDA.n261 0.15675
R6667 VDDA.n263 VDDA.n262 0.15675
R6668 VDDA.n263 VDDA.n14 0.15675
R6669 VDDA.n267 VDDA.n14 0.15675
R6670 VDDA.n268 VDDA.n267 0.15675
R6671 VDDA.n269 VDDA.n268 0.15675
R6672 VDDA.n269 VDDA.n11 0.15675
R6673 VDDA.n274 VDDA.n11 0.15675
R6674 VDDA.n275 VDDA.n274 0.15675
R6675 VDDA.n276 VDDA.n275 0.15675
R6676 VDDA.n276 VDDA.n9 0.15675
R6677 VDDA.n280 VDDA.n9 0.15675
R6678 VDDA.n281 VDDA.n280 0.15675
R6679 VDDA.n281 VDDA.n6 0.15675
R6680 VDDA.n285 VDDA.n6 0.15675
R6681 VDDA.n286 VDDA.n285 0.15675
R6682 VDDA.n287 VDDA.n286 0.15675
R6683 VDDA.n287 VDDA.n4 0.15675
R6684 VDDA.n293 VDDA.n4 0.15675
R6685 VDDA.n294 VDDA.n293 0.15675
R6686 VDDA.n295 VDDA.n294 0.15675
R6687 VDDA.n295 VDDA.n2 0.15675
R6688 VDDA.n299 VDDA.n2 0.15675
R6689 VDDA.n499 VDDA.n498 0.15675
R6690 VDDA.n499 VDDA.n442 0.15675
R6691 VDDA.n504 VDDA.n442 0.15675
R6692 VDDA.n507 VDDA.n506 0.15675
R6693 VDDA.n507 VDDA.n439 0.15675
R6694 VDDA.n511 VDDA.n439 0.15675
R6695 VDDA.n514 VDDA.n513 0.15675
R6696 VDDA.n514 VDDA.n436 0.15675
R6697 VDDA.n518 VDDA.n436 0.15675
R6698 VDDA.n521 VDDA.n520 0.15675
R6699 VDDA.n521 VDDA.n433 0.15675
R6700 VDDA.n525 VDDA.n433 0.15675
R6701 VDDA.n528 VDDA.n527 0.15675
R6702 VDDA.n532 VDDA.n531 0.15675
R6703 VDDA.n533 VDDA.n532 0.15675
R6704 VDDA.n533 VDDA.n428 0.15675
R6705 VDDA.n724 VDDA.n705 0.15675
R6706 VDDA.n725 VDDA.n724 0.15675
R6707 VDDA.n726 VDDA.n725 0.15675
R6708 VDDA.n726 VDDA.n702 0.15675
R6709 VDDA.n731 VDDA.n702 0.15675
R6710 VDDA.n732 VDDA.n731 0.15675
R6711 VDDA.n733 VDDA.n732 0.15675
R6712 VDDA.n733 VDDA.n699 0.15675
R6713 VDDA.n699 VDDA.n698 0.15675
R6714 VDDA.n738 VDDA.n698 0.15675
R6715 VDDA.n739 VDDA.n738 0.15675
R6716 VDDA.n740 VDDA.n739 0.15675
R6717 VDDA.n741 VDDA.n740 0.15675
R6718 VDDA.n741 VDDA.n696 0.15675
R6719 VDDA.n696 VDDA.n695 0.15675
R6720 VDDA.n695 VDDA.n694 0.15675
R6721 VDDA.n694 VDDA.n676 0.15675
R6722 VDDA.n690 VDDA.n676 0.15675
R6723 VDDA.n690 VDDA.n689 0.15675
R6724 VDDA.n689 VDDA.n688 0.15675
R6725 VDDA.n688 VDDA.n679 0.15675
R6726 VDDA.n684 VDDA.n679 0.15675
R6727 VDDA.n684 VDDA.n683 0.15675
R6728 VDDA.n683 VDDA.n682 0.15675
R6729 VDDA.n682 VDDA.n662 0.15675
R6730 VDDA.n764 VDDA.n662 0.15675
R6731 VDDA.n765 VDDA.n764 0.15675
R6732 VDDA.n766 VDDA.n765 0.15675
R6733 VDDA.n785 VDDA.n784 0.15675
R6734 VDDA.n786 VDDA.n785 0.15675
R6735 VDDA.n786 VDDA.n361 0.15675
R6736 VDDA.n790 VDDA.n361 0.15675
R6737 VDDA.n791 VDDA.n790 0.15675
R6738 VDDA.n794 VDDA.n791 0.15675
R6739 VDDA.n794 VDDA.n793 0.15675
R6740 VDDA.n793 VDDA.n792 0.15675
R6741 VDDA.n864 VDDA.n863 0.15675
R6742 VDDA.n865 VDDA.n864 0.15675
R6743 VDDA.n865 VDDA.n339 0.15675
R6744 VDDA.n869 VDDA.n339 0.15675
R6745 VDDA.n870 VDDA.n869 0.15675
R6746 VDDA.n870 VDDA.n337 0.15675
R6747 VDDA.n874 VDDA.n337 0.15675
R6748 VDDA.n875 VDDA.n874 0.15675
R6749 VDDA.n876 VDDA.n875 0.15675
R6750 VDDA.n876 VDDA.n333 0.15675
R6751 VDDA.n882 VDDA.n333 0.15675
R6752 VDDA.n883 VDDA.n882 0.15675
R6753 VDDA.n884 VDDA.n883 0.15675
R6754 VDDA.n884 VDDA.n323 0.15675
R6755 VDDA.n905 VDDA.n323 0.15675
R6756 VDDA.n906 VDDA.n905 0.15675
R6757 VDDA.n907 VDDA.n906 0.15675
R6758 VDDA.n907 VDDA.n314 0.15675
R6759 VDDA.n977 VDDA.n314 0.15675
R6760 VDDA.n978 VDDA.n977 0.15675
R6761 VDDA.n979 VDDA.n978 0.15675
R6762 VDDA.n979 VDDA.n312 0.15675
R6763 VDDA.n983 VDDA.n312 0.15675
R6764 VDDA.n984 VDDA.n983 0.15675
R6765 VDDA.n985 VDDA.n984 0.15675
R6766 VDDA.n985 VDDA.n310 0.15675
R6767 VDDA.n989 VDDA.n310 0.15675
R6768 VDDA.n990 VDDA.n989 0.15675
R6769 VDDA.n990 VDDA.n306 0.15675
R6770 VDDA.n995 VDDA.n306 0.15675
R6771 VDDA.n996 VDDA.n995 0.15675
R6772 VDDA.n997 VDDA.n996 0.15675
R6773 VDDA.n997 VDDA.n304 0.15675
R6774 VDDA.n1001 VDDA.n304 0.15675
R6775 VDDA.n1002 VDDA.n1001 0.15675
R6776 VDDA.n1003 VDDA.n1002 0.15675
R6777 VDDA.n1003 VDDA.n0 0.15675
R6778 VDDA.t127 VDDA.t86 0.137822
R6779 VDDA.n366 VDDA.t129 0.1368
R6780 VDDA.n426 VDDA.n369 0.1255
R6781 VDDA.n373 VDDA.n369 0.1255
R6782 VDDA.n375 VDDA.n373 0.1255
R6783 VDDA.n377 VDDA.n375 0.1255
R6784 VDDA.n379 VDDA.n377 0.1255
R6785 VDDA.n381 VDDA.n379 0.1255
R6786 VDDA.n383 VDDA.n381 0.1255
R6787 VDDA.n385 VDDA.n383 0.1255
R6788 VDDA.n387 VDDA.n385 0.1255
R6789 VDDA.n417 VDDA.n387 0.1255
R6790 VDDA.n416 VDDA.n389 0.1255
R6791 VDDA.n393 VDDA.n389 0.1255
R6792 VDDA.n395 VDDA.n393 0.1255
R6793 VDDA.n397 VDDA.n395 0.1255
R6794 VDDA.n399 VDDA.n397 0.1255
R6795 VDDA.n401 VDDA.n399 0.1255
R6796 VDDA.n403 VDDA.n401 0.1255
R6797 VDDA.n405 VDDA.n403 0.1255
R6798 VDDA.n407 VDDA.n405 0.1255
R6799 VDDA VDDA.n0 0.1255
R6800 VDDA.n766 VDDA 0.122375
R6801 VDDA.n497 VDDA.n496 0.100307
R6802 VDDA.n498 VDDA.n497 0.09425
R6803 VDDA.n506 VDDA.n505 0.09425
R6804 VDDA.n513 VDDA.n512 0.09425
R6805 VDDA.n520 VDDA.n519 0.09425
R6806 VDDA.n527 VDDA.n526 0.09425
R6807 VDDA.n531 VDDA.n430 0.09425
R6808 VDDA.n792 VDDA.n341 0.078625
R6809 VDDA.n863 VDDA.n341 0.078625
R6810 VDDA VDDA.n1007 0.063
R6811 VDDA.n505 VDDA.n504 0.063
R6812 VDDA.n512 VDDA.n511 0.063
R6813 VDDA.n519 VDDA.n518 0.063
R6814 VDDA.n526 VDDA.n525 0.063
R6815 VDDA.n528 VDDA.n430 0.063
R6816 VDDA.n768 VDDA 0.0505
R6817 VDDA.n366 VDDA.t366 0.00152174
R6818 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 517.347
R6819 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R6820 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R6821 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 228.148
R6822 pfd_8_0.F_b.t0 pfd_8_0.F_b.n2 221.411
R6823 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R6824 pfd_8_0.F_b.n1 pfd_8_0.F_b.t1 24.0005
R6825 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R6826 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R6827 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R6828 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R6829 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R6830 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R6831 pfd_8_0.F.t1 pfd_8_0.F.n4 221.411
R6832 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R6833 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R6834 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R6835 pfd_8_0.F.n1 pfd_8_0.F.t0 24.0005
R6836 VCO_FD_magic_0.div120_2_0.div4.t3 VCO_FD_magic_0.div120_2_0.div4.t6 1012.2
R6837 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t1 663.801
R6838 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n1 431.401
R6839 VCO_FD_magic_0.div120_2_0.div4.t2 VCO_FD_magic_0.div120_2_0.div4.t4 401.668
R6840 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t3 361.692
R6841 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t5 353.467
R6842 VCO_FD_magic_0.div120_2_0.div4.t0 VCO_FD_magic_0.div120_2_0.div4.n2 298.921
R6843 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t2 257.067
R6844 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n0 67.2005
R6845 a_6330_n1530.n4 a_6330_n1530.t1 752.333
R6846 a_6330_n1530.t2 a_6330_n1530.n5 752.333
R6847 a_6330_n1530.n0 a_6330_n1530.t3 514.134
R6848 a_6330_n1530.n3 a_6330_n1530.n2 366.856
R6849 a_6330_n1530.n5 a_6330_n1530.t0 254.333
R6850 a_6330_n1530.n3 a_6330_n1530.t6 190.123
R6851 a_6330_n1530.n4 a_6330_n1530.n3 187.201
R6852 a_6330_n1530.n2 a_6330_n1530.n1 176.733
R6853 a_6330_n1530.n1 a_6330_n1530.n0 176.733
R6854 a_6330_n1530.n2 a_6330_n1530.t4 112.468
R6855 a_6330_n1530.n1 a_6330_n1530.t5 112.468
R6856 a_6330_n1530.n0 a_6330_n1530.t7 112.468
R6857 a_6330_n1530.n5 a_6330_n1530.n4 70.4005
R6858 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t25 363.909
R6859 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 351.88
R6860 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 299.252
R6861 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n9 299.25
R6862 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n4 299.25
R6863 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t2 242.968
R6864 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 200.477
R6865 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 199.727
R6866 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t30 194.809
R6867 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t28 194.809
R6868 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t11 194.809
R6869 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t17 194.809
R6870 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 163.097
R6871 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 161.653
R6872 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t1 48.0005
R6873 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t0 48.0005
R6874 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t4 48.0005
R6875 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 48.0005
R6876 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t7 39.4005
R6877 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t9 39.4005
R6878 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t10 39.4005
R6879 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t8 39.4005
R6880 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t6 39.4005
R6881 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t5 39.4005
R6882 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n2 11.6665
R6883 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 5.2505
R6884 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t27 4.8248
R6885 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t22 4.5005
R6886 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R6887 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t31 4.5005
R6888 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t21 4.5005
R6889 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t13 4.5005
R6890 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t33 4.5005
R6891 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t23 4.5005
R6892 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t19 4.5005
R6893 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t36 4.5005
R6894 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t14 4.5005
R6895 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R6896 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R6897 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t12 4.5005
R6898 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t32 4.5005
R6899 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R6900 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R6901 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t35 4.5005
R6902 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t29 4.5005
R6903 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t20 4.5005
R6904 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.2388
R6905 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 2.80435
R6906 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.n0 2.6325
R6907 bgr_0.V_TOP.n1 bgr_0.V_TOP.t33 312.798
R6908 bgr_0.V_TOP bgr_0.V_TOP.t47 312.639
R6909 bgr_0.V_TOP.n44 bgr_0.V_TOP.t44 312.5
R6910 bgr_0.V_TOP.n50 bgr_0.V_TOP.t43 310.401
R6911 bgr_0.V_TOP.n49 bgr_0.V_TOP.t30 310.401
R6912 bgr_0.V_TOP.n48 bgr_0.V_TOP.t18 310.401
R6913 bgr_0.V_TOP.n47 bgr_0.V_TOP.t21 310.401
R6914 bgr_0.V_TOP.n46 bgr_0.V_TOP.t36 310.401
R6915 bgr_0.V_TOP.n45 bgr_0.V_TOP.t39 310.401
R6916 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 310.401
R6917 bgr_0.V_TOP.n4 bgr_0.V_TOP.t32 310.401
R6918 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 310.401
R6919 bgr_0.V_TOP.n2 bgr_0.V_TOP.t41 310.401
R6920 bgr_0.V_TOP.n1 bgr_0.V_TOP.t19 310.401
R6921 bgr_0.V_TOP.n42 bgr_0.V_TOP.t48 308
R6922 bgr_0.V_TOP.n31 bgr_0.V_TOP.n29 306.808
R6923 bgr_0.V_TOP.n7 bgr_0.V_TOP.t14 305.901
R6924 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 301.933
R6925 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 301.933
R6926 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 301.933
R6927 bgr_0.V_TOP.n32 bgr_0.V_TOP.n28 297.433
R6928 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 297.433
R6929 bgr_0.V_TOP.n27 bgr_0.V_TOP.t1 108.898
R6930 bgr_0.V_TOP.n40 bgr_0.V_TOP.t3 98.9217
R6931 bgr_0.V_TOP.n28 bgr_0.V_TOP.t5 39.4005
R6932 bgr_0.V_TOP.n28 bgr_0.V_TOP.t10 39.4005
R6933 bgr_0.V_TOP.n29 bgr_0.V_TOP.t2 39.4005
R6934 bgr_0.V_TOP.n29 bgr_0.V_TOP.t7 39.4005
R6935 bgr_0.V_TOP.n30 bgr_0.V_TOP.t6 39.4005
R6936 bgr_0.V_TOP.n30 bgr_0.V_TOP.t0 39.4005
R6937 bgr_0.V_TOP.n38 bgr_0.V_TOP.t12 39.4005
R6938 bgr_0.V_TOP.n38 bgr_0.V_TOP.t4 39.4005
R6939 bgr_0.V_TOP.n36 bgr_0.V_TOP.t11 39.4005
R6940 bgr_0.V_TOP.n36 bgr_0.V_TOP.t13 39.4005
R6941 bgr_0.V_TOP.n34 bgr_0.V_TOP.t9 39.4005
R6942 bgr_0.V_TOP.n34 bgr_0.V_TOP.t8 39.4005
R6943 bgr_0.V_TOP.n33 bgr_0.V_TOP.n27 13.563
R6944 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 12.3446
R6945 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 4.90675
R6946 bgr_0.V_TOP.n8 bgr_0.V_TOP.t24 4.8248
R6947 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 4.5005
R6948 bgr_0.V_TOP.n41 bgr_0.V_TOP.n0 4.5005
R6949 bgr_0.V_TOP.n43 bgr_0.V_TOP.n42 4.5005
R6950 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 4.5005
R6951 bgr_0.V_TOP.n16 bgr_0.V_TOP.t25 4.5005
R6952 bgr_0.V_TOP.n15 bgr_0.V_TOP.t15 4.5005
R6953 bgr_0.V_TOP.n14 bgr_0.V_TOP.t22 4.5005
R6954 bgr_0.V_TOP.n13 bgr_0.V_TOP.t17 4.5005
R6955 bgr_0.V_TOP.n12 bgr_0.V_TOP.t46 4.5005
R6956 bgr_0.V_TOP.n11 bgr_0.V_TOP.t34 4.5005
R6957 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.5005
R6958 bgr_0.V_TOP.n9 bgr_0.V_TOP.t29 4.5005
R6959 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.5005
R6960 bgr_0.V_TOP.n17 bgr_0.V_TOP.t38 4.5005
R6961 bgr_0.V_TOP.n18 bgr_0.V_TOP.t23 4.5005
R6962 bgr_0.V_TOP.n19 bgr_0.V_TOP.t31 4.5005
R6963 bgr_0.V_TOP.n20 bgr_0.V_TOP.t26 4.5005
R6964 bgr_0.V_TOP.n21 bgr_0.V_TOP.t16 4.5005
R6965 bgr_0.V_TOP.n22 bgr_0.V_TOP.t45 4.5005
R6966 bgr_0.V_TOP.n23 bgr_0.V_TOP.t49 4.5005
R6967 bgr_0.V_TOP.n24 bgr_0.V_TOP.t40 4.5005
R6968 bgr_0.V_TOP.n25 bgr_0.V_TOP.t28 4.5005
R6969 bgr_0.V_TOP.n26 bgr_0.V_TOP.t35 4.5005
R6970 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 1.59425
R6971 bgr_0.V_TOP.n41 bgr_0.V_TOP.n40 1.21925
R6972 bgr_0.V_TOP.n35 bgr_0.V_TOP.n33 1.1255
R6973 bgr_0.V_TOP.n37 bgr_0.V_TOP.n35 1.1255
R6974 bgr_0.V_TOP.n39 bgr_0.V_TOP.n37 1.1255
R6975 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R6976 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R6977 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.3295
R6978 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R6979 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 0.3295
R6980 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R6981 bgr_0.V_TOP.n10 bgr_0.V_TOP.n9 0.3295
R6982 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R6983 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 0.3295
R6984 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 0.3295
R6985 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 0.3295
R6986 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 0.3295
R6987 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 0.3295
R6988 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 0.3295
R6989 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 0.3295
R6990 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 0.3295
R6991 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 0.3248
R6992 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 0.2825
R6993 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 0.28175
R6994 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 0.28175
R6995 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 0.28175
R6996 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 0.28175
R6997 bgr_0.V_TOP.n6 bgr_0.V_TOP.n5 0.28175
R6998 bgr_0.V_TOP.n44 bgr_0.V_TOP.n43 0.28175
R6999 bgr_0.V_TOP.n45 bgr_0.V_TOP.n44 0.28175
R7000 bgr_0.V_TOP.n46 bgr_0.V_TOP.n45 0.28175
R7001 bgr_0.V_TOP.n47 bgr_0.V_TOP.n46 0.28175
R7002 bgr_0.V_TOP.n48 bgr_0.V_TOP.n47 0.28175
R7003 bgr_0.V_TOP.n49 bgr_0.V_TOP.n48 0.28175
R7004 bgr_0.V_TOP.n50 bgr_0.V_TOP.n49 0.28175
R7005 bgr_0.V_TOP.n6 bgr_0.V_TOP.n0 0.141125
R7006 bgr_0.V_TOP.n43 bgr_0.V_TOP.n0 0.141125
R7007 bgr_0.V_TOP bgr_0.V_TOP.n50 0.141125
R7008 bgr_0.V_TOP.n41 bgr_0.V_TOP.n7 0.141125
R7009 bgr_0.V_TOP.n42 bgr_0.V_TOP.n41 0.141125
R7010 pfd_8_0.QB.t8 pfd_8_0.QB.t7 835.467
R7011 pfd_8_0.QB.n1 pfd_8_0.QB.t8 564.496
R7012 pfd_8_0.QB.n2 pfd_8_0.QB.t3 517.347
R7013 pfd_8_0.QB.n0 pfd_8_0.QB.t5 514.134
R7014 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R7015 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R7016 pfd_8_0.QB.n0 pfd_8_0.QB.t6 273.134
R7017 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R7018 pfd_8_0.QB.n2 pfd_8_0.QB.t4 228.148
R7019 pfd_8_0.QB.n4 pfd_8_0.QB.t2 221.411
R7020 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R7021 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R7022 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R7023 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R7024 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R7025 a_n30_630.t0 a_n30_630.t1 39.4005
R7026 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t6 1188.93
R7027 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R7028 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t5 835.467
R7029 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t3 562.333
R7030 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R7031 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R7032 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t4 224.934
R7033 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t2 221.411
R7034 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t1 24.0005
R7035 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t0 24.0005
R7036 V_OSC.t4 V_OSC.t6 401.668
R7037 V_OSC.n1 V_OSC.t0 372.118
R7038 V_OSC.n3 V_OSC.t3 353.467
R7039 V_OSC V_OSC.n3 313.3
R7040 V_OSC.n3 V_OSC.t4 257.067
R7041 V_OSC.n1 V_OSC.t1 247.934
R7042 V_OSC.n2 V_OSC.n1 236.756
R7043 V_OSC.n0 V_OSC.t2 224.934
R7044 V_OSC.n2 V_OSC.n0 224.934
R7045 V_OSC.n0 V_OSC.t5 144.601
R7046 V_OSC V_OSC.n2 120.501
R7047 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t1 421.027
R7048 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t2 348.81
R7049 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.t0 280.05
R7050 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.n0 36.1094
R7051 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.n0 437.733
R7052 VCO_FD_magic_0.vco2_3_0.V9.t1 VCO_FD_magic_0.vco2_3_0.V9.n1 372.118
R7053 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.t0 247.934
R7054 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t2 224.934
R7055 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t3 144.601
R7056 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t34 362.341
R7057 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t25 355.094
R7058 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n8 302.183
R7059 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n6 302.183
R7060 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.n5 302.183
R7061 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t6 242.968
R7062 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n9 200.477
R7063 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 199.727
R7064 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t16 194.809
R7065 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t13 194.809
R7066 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t24 194.809
R7067 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t20 194.809
R7068 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n7 166.03
R7069 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n12 161.53
R7070 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t3 48.0005
R7071 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t7 48.0005
R7072 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t0 48.0005
R7073 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t5 48.0005
R7074 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n2 40.0796
R7075 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t10 39.4005
R7076 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t4 39.4005
R7077 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t8 39.4005
R7078 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t9 39.4005
R7079 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t2 39.4005
R7080 bgr_0.1st_Vout_2.t1 bgr_0.1st_Vout_2.n14 39.4005
R7081 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n11 5.2505
R7082 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n4 4.92238
R7083 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t35 4.8248
R7084 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t36 4.5005
R7085 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t28 4.5005
R7086 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t32 4.5005
R7087 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t29 4.5005
R7088 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R7089 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R7090 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.5005
R7091 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t12 4.5005
R7092 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t31 4.5005
R7093 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t27 4.5005
R7094 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t18 4.5005
R7095 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R7096 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.5005
R7097 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t14 4.5005
R7098 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R7099 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.5005
R7100 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.5005
R7101 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R7102 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.5005
R7103 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n1 3.2388
R7104 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n13 2.90725
R7105 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 2.6325
R7106 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n3 2.2505
R7107 bgr_0.cap_res2.t0 bgr_0.cap_res2.t2 138.543
R7108 bgr_0.cap_res2.t12 bgr_0.cap_res2.t10 0.1603
R7109 bgr_0.cap_res2.t6 bgr_0.cap_res2.t12 0.1603
R7110 bgr_0.cap_res2.t20 bgr_0.cap_res2.t6 0.1603
R7111 bgr_0.cap_res2.t3 bgr_0.cap_res2.t20 0.1603
R7112 bgr_0.cap_res2.t18 bgr_0.cap_res2.t3 0.1603
R7113 bgr_0.cap_res2.t14 bgr_0.cap_res2.t18 0.1603
R7114 bgr_0.cap_res2.t11 bgr_0.cap_res2.t14 0.1603
R7115 bgr_0.cap_res2.t15 bgr_0.cap_res2.t11 0.1603
R7116 bgr_0.cap_res2.t4 bgr_0.cap_res2.t8 0.1603
R7117 bgr_0.cap_res2.t7 bgr_0.cap_res2.t4 0.1603
R7118 bgr_0.cap_res2.t13 bgr_0.cap_res2.t7 0.1603
R7119 bgr_0.cap_res2.t17 bgr_0.cap_res2.t13 0.1603
R7120 bgr_0.cap_res2.t16 bgr_0.cap_res2.t17 0.1603
R7121 bgr_0.cap_res2.t19 bgr_0.cap_res2.t16 0.1603
R7122 bgr_0.cap_res2.t5 bgr_0.cap_res2.t19 0.1603
R7123 bgr_0.cap_res2.t2 bgr_0.cap_res2.t5 0.1603
R7124 bgr_0.cap_res2.t1 bgr_0.cap_res2.n0 0.159278
R7125 bgr_0.cap_res2.t8 bgr_0.cap_res2.t1 0.137822
R7126 bgr_0.cap_res2.n0 bgr_0.cap_res2.t15 0.1368
R7127 bgr_0.cap_res2.n0 bgr_0.cap_res2.t9 0.00152174
R7128 bgr_0.Vin+.n5 bgr_0.Vin+.t8 291.502
R7129 bgr_0.Vin+.n5 bgr_0.Vin+.t9 291.288
R7130 bgr_0.Vin+.n6 bgr_0.Vin+.t6 291.288
R7131 bgr_0.Vin+.n7 bgr_0.Vin+.t7 291.288
R7132 bgr_0.Vin+.n8 bgr_0.Vin+.t10 291.288
R7133 bgr_0.Vin+.n0 bgr_0.Vin+.t1 148.653
R7134 bgr_0.Vin+.n0 bgr_0.Vin+.t0 125.371
R7135 bgr_0.Vin+.n3 bgr_0.Vin+.n1 105.609
R7136 bgr_0.Vin+.n3 bgr_0.Vin+.n2 104.484
R7137 bgr_0.Vin+.n4 bgr_0.Vin+.n0 21.4246
R7138 bgr_0.Vin+.n4 bgr_0.Vin+.n3 14.2349
R7139 bgr_0.Vin+.n1 bgr_0.Vin+.t2 13.1338
R7140 bgr_0.Vin+.n1 bgr_0.Vin+.t3 13.1338
R7141 bgr_0.Vin+.n2 bgr_0.Vin+.t4 13.1338
R7142 bgr_0.Vin+.n2 bgr_0.Vin+.t5 13.1338
R7143 bgr_0.Vin+ bgr_0.Vin+.n4 4.67014
R7144 bgr_0.Vin+ bgr_0.Vin+.n8 1.76657
R7145 bgr_0.Vin+.n8 bgr_0.Vin+.n7 0.643357
R7146 bgr_0.Vin+.n6 bgr_0.Vin+.n5 0.643357
R7147 bgr_0.Vin+.n7 bgr_0.Vin+.n6 0.214786
R7148 bgr_0.V2.n0 bgr_0.V2.t28 403.952
R7149 bgr_0.V2.n18 bgr_0.V2.t27 403.755
R7150 bgr_0.V2.n17 bgr_0.V2.t18 403.755
R7151 bgr_0.V2.n16 bgr_0.V2.t29 403.755
R7152 bgr_0.V2.n15 bgr_0.V2.t20 403.755
R7153 bgr_0.V2.n14 bgr_0.V2.t26 403.755
R7154 bgr_0.V2.n13 bgr_0.V2.t16 403.755
R7155 bgr_0.V2.n12 bgr_0.V2.t13 403.755
R7156 bgr_0.V2.n11 bgr_0.V2.t17 403.755
R7157 bgr_0.V2.n10 bgr_0.V2.t24 403.755
R7158 bgr_0.V2.n9 bgr_0.V2.t15 403.755
R7159 bgr_0.V2.n8 bgr_0.V2.t23 403.755
R7160 bgr_0.V2.n7 bgr_0.V2.t14 403.755
R7161 bgr_0.V2.n6 bgr_0.V2.t22 403.755
R7162 bgr_0.V2.n5 bgr_0.V2.t12 403.755
R7163 bgr_0.V2.n4 bgr_0.V2.t21 403.755
R7164 bgr_0.V2.n3 bgr_0.V2.t10 403.755
R7165 bgr_0.V2.n2 bgr_0.V2.t25 403.755
R7166 bgr_0.V2.n1 bgr_0.V2.t11 403.755
R7167 bgr_0.V2.n0 bgr_0.V2.t19 403.755
R7168 bgr_0.V2.n26 bgr_0.V2.n25 301.933
R7169 bgr_0.V2.n24 bgr_0.V2.n23 301.933
R7170 bgr_0.V2.n22 bgr_0.V2.n21 301.933
R7171 bgr_0.V2.n20 bgr_0.V2.n19 301.933
R7172 bgr_0.V2 bgr_0.V2.t0 116.322
R7173 bgr_0.V2.n20 bgr_0.V2.t7 103.828
R7174 bgr_0.V2.n25 bgr_0.V2.t1 39.4005
R7175 bgr_0.V2.n25 bgr_0.V2.t9 39.4005
R7176 bgr_0.V2.n23 bgr_0.V2.t6 39.4005
R7177 bgr_0.V2.n23 bgr_0.V2.t5 39.4005
R7178 bgr_0.V2.n21 bgr_0.V2.t4 39.4005
R7179 bgr_0.V2.n21 bgr_0.V2.t3 39.4005
R7180 bgr_0.V2.n19 bgr_0.V2.t8 39.4005
R7181 bgr_0.V2.n19 bgr_0.V2.t2 39.4005
R7182 bgr_0.V2.n27 bgr_0.V2.n18 10.3335
R7183 bgr_0.V2.n27 bgr_0.V2.n26 5.313
R7184 bgr_0.V2.n9 bgr_0.V2.n8 1.6255
R7185 bgr_0.V2.n22 bgr_0.V2.n20 1.1255
R7186 bgr_0.V2.n24 bgr_0.V2.n22 1.1255
R7187 bgr_0.V2.n26 bgr_0.V2.n24 1.1255
R7188 bgr_0.V2 bgr_0.V2.n27 0.688
R7189 bgr_0.V2.n1 bgr_0.V2.n0 0.196929
R7190 bgr_0.V2.n2 bgr_0.V2.n1 0.196929
R7191 bgr_0.V2.n3 bgr_0.V2.n2 0.196929
R7192 bgr_0.V2.n4 bgr_0.V2.n3 0.196929
R7193 bgr_0.V2.n5 bgr_0.V2.n4 0.196929
R7194 bgr_0.V2.n6 bgr_0.V2.n5 0.196929
R7195 bgr_0.V2.n7 bgr_0.V2.n6 0.196929
R7196 bgr_0.V2.n8 bgr_0.V2.n7 0.196929
R7197 bgr_0.V2.n10 bgr_0.V2.n9 0.196929
R7198 bgr_0.V2.n11 bgr_0.V2.n10 0.196929
R7199 bgr_0.V2.n12 bgr_0.V2.n11 0.196929
R7200 bgr_0.V2.n13 bgr_0.V2.n12 0.196929
R7201 bgr_0.V2.n14 bgr_0.V2.n13 0.196929
R7202 bgr_0.V2.n15 bgr_0.V2.n14 0.196929
R7203 bgr_0.V2.n16 bgr_0.V2.n15 0.196929
R7204 bgr_0.V2.n17 bgr_0.V2.n16 0.196929
R7205 bgr_0.V2.n18 bgr_0.V2.n17 0.196929
R7206 BGR_CURRENT_OUT.n5 BGR_CURRENT_OUT.n4 1269.42
R7207 BGR_CURRENT_OUT.n23 BGR_CURRENT_OUT.n9 297.663
R7208 BGR_CURRENT_OUT.n21 BGR_CURRENT_OUT.n20 297.663
R7209 bgr_0.CURRENT_OUTPUT BGR_CURRENT_OUT.n11 297.663
R7210 BGR_CURRENT_OUT.n16 BGR_CURRENT_OUT.n14 297.663
R7211 BGR_CURRENT_OUT.n13 BGR_CURRENT_OUT.n12 297.663
R7212 BGR_CURRENT_OUT.n18 BGR_CURRENT_OUT.n17 297.663
R7213 BGR_CURRENT_OUT.n5 BGR_CURRENT_OUT.t1 275.325
R7214 BGR_CURRENT_OUT.n7 BGR_CURRENT_OUT.n6 248.4
R7215 BGR_CURRENT_OUT.n8 BGR_CURRENT_OUT.t17 238.892
R7216 BGR_CURRENT_OUT.n24 BGR_CURRENT_OUT.n8 165.863
R7217 BGR_CURRENT_OUT.n8 BGR_CURRENT_OUT.t0 161.371
R7218 BGR_CURRENT_OUT.n4 BGR_CURRENT_OUT.t18 151.792
R7219 BGR_CURRENT_OUT.n6 BGR_CURRENT_OUT.t3 140.583
R7220 BGR_CURRENT_OUT.n6 BGR_CURRENT_OUT.t1 140.583
R7221 BGR_CURRENT_OUT.n7 BGR_CURRENT_OUT.n3 98.6614
R7222 BGR_CURRENT_OUT.t3 BGR_CURRENT_OUT.n5 80.3338
R7223 BGR_CURRENT_OUT.n4 BGR_CURRENT_OUT.t19 44.2902
R7224 BGR_CURRENT_OUT.n9 BGR_CURRENT_OUT.t7 39.4005
R7225 BGR_CURRENT_OUT.n9 BGR_CURRENT_OUT.t16 39.4005
R7226 BGR_CURRENT_OUT.n20 BGR_CURRENT_OUT.t8 39.4005
R7227 BGR_CURRENT_OUT.n20 BGR_CURRENT_OUT.t11 39.4005
R7228 BGR_CURRENT_OUT.n11 BGR_CURRENT_OUT.t9 39.4005
R7229 BGR_CURRENT_OUT.n11 BGR_CURRENT_OUT.t12 39.4005
R7230 BGR_CURRENT_OUT.n14 BGR_CURRENT_OUT.t10 39.4005
R7231 BGR_CURRENT_OUT.n14 BGR_CURRENT_OUT.t13 39.4005
R7232 BGR_CURRENT_OUT.n12 BGR_CURRENT_OUT.t15 39.4005
R7233 BGR_CURRENT_OUT.n12 BGR_CURRENT_OUT.t5 39.4005
R7234 BGR_CURRENT_OUT.n17 BGR_CURRENT_OUT.t6 39.4005
R7235 BGR_CURRENT_OUT.n17 BGR_CURRENT_OUT.t14 39.4005
R7236 BGR_CURRENT_OUT.n25 BGR_CURRENT_OUT.n24 15.4229
R7237 BGR_CURRENT_OUT.n3 BGR_CURRENT_OUT.t4 15.0005
R7238 BGR_CURRENT_OUT.n3 BGR_CURRENT_OUT.t2 15.0005
R7239 BGR_CURRENT_OUT.n15 BGR_CURRENT_OUT.n13 4.84425
R7240 BGR_CURRENT_OUT.n23 BGR_CURRENT_OUT.n22 4.84425
R7241 BGR_CURRENT_OUT.n16 BGR_CURRENT_OUT.n15 4.5005
R7242 BGR_CURRENT_OUT.n19 bgr_0.CURRENT_OUTPUT 4.5005
R7243 BGR_CURRENT_OUT.n22 BGR_CURRENT_OUT.n21 4.5005
R7244 BGR_CURRENT_OUT.n18 BGR_CURRENT_OUT.n10 4.5005
R7245 BGR_CURRENT_OUT.n0 BGR_CURRENT_OUT.n24 9.36731
R7246 BGR_CURRENT_OUT.n1 BGR_CURRENT_OUT.n13 1.85607
R7247 BGR_CURRENT_OUT.n0 BGR_CURRENT_OUT.n23 1.74185
R7248 BGR_CURRENT_OUT.n21 BGR_CURRENT_OUT.n0 1.74185
R7249 BGR_CURRENT_OUT.n1 BGR_CURRENT_OUT.n16 1.74185
R7250 BGR_CURRENT_OUT.n2 BGR_CURRENT_OUT.n18 1.74185
R7251 bgr_0.CURRENT_OUTPUT BGR_CURRENT_OUT.n2 1.74185
R7252 charge_pump_cell_6_0.I_IN BGR_CURRENT_OUT.n25 1.6005
R7253 BGR_CURRENT_OUT.n25 BGR_CURRENT_OUT.n7 1.6005
R7254 BGR_CURRENT_OUT.n15 BGR_CURRENT_OUT.n10 0.34425
R7255 BGR_CURRENT_OUT.n19 BGR_CURRENT_OUT.n10 0.34425
R7256 BGR_CURRENT_OUT.n22 BGR_CURRENT_OUT.n19 0.34425
R7257 BGR_CURRENT_OUT.n2 BGR_CURRENT_OUT.n0 0.229667
R7258 BGR_CURRENT_OUT.n2 BGR_CURRENT_OUT.n1 0.229667
R7259 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.n2 919.244
R7260 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n7 912.303
R7261 VCO_FD_magic_0.div120_2_0.div24.t7 VCO_FD_magic_0.div120_2_0.div24.t13 819.4
R7262 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.n8 628.734
R7263 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.n1 520.361
R7264 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.n6 364.178
R7265 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t10 337.401
R7266 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.t7 336.25
R7267 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t12 305.267
R7268 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.t2 257.534
R7269 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.t9 192.8
R7270 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.n0 176.733
R7271 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.n5 176.733
R7272 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.n3 160.667
R7273 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.t11 144.601
R7274 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.t4 131.976
R7275 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.t3 128.534
R7276 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t6 128.534
R7277 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.t14 112.468
R7278 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.t5 112.468
R7279 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.t8 112.468
R7280 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.n4 96.4005
R7281 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t1 78.8005
R7282 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t0 78.8005
R7283 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.n9 11.2005
R7284 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n10 6.4005
R7285 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 710.734
R7286 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 553.534
R7287 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 254.333
R7288 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 206.333
R7289 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 70.4005
R7290 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 48.0005
R7291 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 48.0005
R7292 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 12.8005
R7293 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 777.4
R7294 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 514.134
R7295 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 364.178
R7296 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 353.467
R7297 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 353.467
R7298 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 318.702
R7299 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 307.909
R7300 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 289.2
R7301 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 257.079
R7302 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 233
R7303 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 192.8
R7304 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 176.733
R7305 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 112.468
R7306 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 112.468
R7307 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 112.468
R7308 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 112.468
R7309 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 96.4005
R7310 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 38.2642
R7311 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 21.3338
R7312 pfd_8_0.Reset.n1 pfd_8_0.Reset.t4 562.333
R7313 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R7314 pfd_8_0.Reset.n0 pfd_8_0.Reset.t2 417.733
R7315 pfd_8_0.Reset.n0 pfd_8_0.Reset.t3 369.534
R7316 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R7317 pfd_8_0.Reset.t0 pfd_8_0.Reset.n3 288.37
R7318 pfd_8_0.Reset.n1 pfd_8_0.Reset.t5 224.934
R7319 pfd_8_0.Reset.n3 pfd_8_0.Reset.t1 177.577
R7320 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R7321 a_1390_630.t0 a_1390_630.t1 39.4005
R7322 bgr_0.V1.n6 bgr_0.V1.t11 287.762
R7323 bgr_0.V1.n5 bgr_0.V1.t10 287.762
R7324 bgr_0.V1.n5 bgr_0.V1.t9 287.589
R7325 bgr_0.V1.n8 bgr_0.V1.t8 287.012
R7326 bgr_0.V1.n7 bgr_0.V1.t7 287.012
R7327 bgr_0.V1.t0 bgr_0.V1.n9 115.097
R7328 bgr_0.V1.n2 bgr_0.V1.n0 107.266
R7329 bgr_0.V1.n4 bgr_0.V1.n3 105.016
R7330 bgr_0.V1.n2 bgr_0.V1.n1 105.016
R7331 bgr_0.V1.n3 bgr_0.V1.t4 13.1338
R7332 bgr_0.V1.n3 bgr_0.V1.t2 13.1338
R7333 bgr_0.V1.n1 bgr_0.V1.t3 13.1338
R7334 bgr_0.V1.n1 bgr_0.V1.t5 13.1338
R7335 bgr_0.V1.n0 bgr_0.V1.t1 13.1338
R7336 bgr_0.V1.n0 bgr_0.V1.t6 13.1338
R7337 bgr_0.V1.n9 bgr_0.V1.n4 9.0005
R7338 bgr_0.V1.n9 bgr_0.V1.n8 6.78086
R7339 bgr_0.V1.n4 bgr_0.V1.n2 2.2505
R7340 bgr_0.V1.n7 bgr_0.V1.n6 0.579071
R7341 bgr_0.V1.n8 bgr_0.V1.n7 0.282643
R7342 bgr_0.V1.n6 bgr_0.V1.n5 0.2755
R7343 a_n1450_5080.n15 a_n1450_5080.t19 310.488
R7344 a_n1450_5080.n9 a_n1450_5080.t21 310.488
R7345 a_n1450_5080.n0 a_n1450_5080.t20 310.488
R7346 a_n1450_5080.n13 a_n1450_5080.n12 297.433
R7347 a_n1450_5080.n4 a_n1450_5080.n3 297.433
R7348 a_n1450_5080.n19 a_n1450_5080.n18 297.433
R7349 a_n1450_5080.n7 a_n1450_5080.t13 248.133
R7350 a_n1450_5080.n7 a_n1450_5080.n6 199.383
R7351 a_n1450_5080.n8 a_n1450_5080.n5 194.883
R7352 a_n1450_5080.n17 a_n1450_5080.t2 184.097
R7353 a_n1450_5080.n11 a_n1450_5080.t0 184.097
R7354 a_n1450_5080.n2 a_n1450_5080.t6 184.097
R7355 a_n1450_5080.n16 a_n1450_5080.n15 167.094
R7356 a_n1450_5080.n10 a_n1450_5080.n9 167.094
R7357 a_n1450_5080.n1 a_n1450_5080.n0 167.094
R7358 a_n1450_5080.n18 a_n1450_5080.n17 161.3
R7359 a_n1450_5080.n13 a_n1450_5080.n11 161.3
R7360 a_n1450_5080.n4 a_n1450_5080.n2 161.3
R7361 a_n1450_5080.n15 a_n1450_5080.t17 120.501
R7362 a_n1450_5080.n16 a_n1450_5080.t10 120.501
R7363 a_n1450_5080.n9 a_n1450_5080.t22 120.501
R7364 a_n1450_5080.n10 a_n1450_5080.t4 120.501
R7365 a_n1450_5080.n0 a_n1450_5080.t18 120.501
R7366 a_n1450_5080.n1 a_n1450_5080.t8 120.501
R7367 a_n1450_5080.n6 a_n1450_5080.t15 48.0005
R7368 a_n1450_5080.n6 a_n1450_5080.t12 48.0005
R7369 a_n1450_5080.n5 a_n1450_5080.t14 48.0005
R7370 a_n1450_5080.n5 a_n1450_5080.t16 48.0005
R7371 a_n1450_5080.n17 a_n1450_5080.n16 40.7027
R7372 a_n1450_5080.n11 a_n1450_5080.n10 40.7027
R7373 a_n1450_5080.n2 a_n1450_5080.n1 40.7027
R7374 a_n1450_5080.n12 a_n1450_5080.t5 39.4005
R7375 a_n1450_5080.n12 a_n1450_5080.t1 39.4005
R7376 a_n1450_5080.n3 a_n1450_5080.t9 39.4005
R7377 a_n1450_5080.n3 a_n1450_5080.t7 39.4005
R7378 a_n1450_5080.t11 a_n1450_5080.n19 39.4005
R7379 a_n1450_5080.n19 a_n1450_5080.t3 39.4005
R7380 a_n1450_5080.n14 a_n1450_5080.n4 6.6255
R7381 a_n1450_5080.n18 a_n1450_5080.n14 6.6255
R7382 a_n1450_5080.n8 a_n1450_5080.n7 5.2505
R7383 a_n1450_5080.n14 a_n1450_5080.n13 4.5005
R7384 a_n1450_5080.n13 a_n1450_5080.n8 0.78175
R7385 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 199.935
R7386 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 199.53
R7387 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 199.53
R7388 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 199.53
R7389 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 199.53
R7390 bgr_0.V_p_2.n1 bgr_0.V_p_2.t10 97.8998
R7391 bgr_0.V_p_2.n5 bgr_0.V_p_2.t8 48.0005
R7392 bgr_0.V_p_2.n5 bgr_0.V_p_2.t3 48.0005
R7393 bgr_0.V_p_2.n4 bgr_0.V_p_2.t5 48.0005
R7394 bgr_0.V_p_2.n4 bgr_0.V_p_2.t1 48.0005
R7395 bgr_0.V_p_2.n3 bgr_0.V_p_2.t2 48.0005
R7396 bgr_0.V_p_2.n3 bgr_0.V_p_2.t6 48.0005
R7397 bgr_0.V_p_2.n2 bgr_0.V_p_2.t7 48.0005
R7398 bgr_0.V_p_2.n2 bgr_0.V_p_2.t0 48.0005
R7399 bgr_0.V_p_2.n6 bgr_0.V_p_2.t4 48.0005
R7400 bgr_0.V_p_2.t9 bgr_0.V_p_2.n6 48.0005
R7401 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.09425
R7402 bgr_0.cap_res1.t0 bgr_0.cap_res1.t8 130.1
R7403 bgr_0.cap_res1.t7 bgr_0.cap_res1.t14 0.1603
R7404 bgr_0.cap_res1.t2 bgr_0.cap_res1.t7 0.1603
R7405 bgr_0.cap_res1.t16 bgr_0.cap_res1.t2 0.1603
R7406 bgr_0.cap_res1.t9 bgr_0.cap_res1.t16 0.1603
R7407 bgr_0.cap_res1.t5 bgr_0.cap_res1.t9 0.1603
R7408 bgr_0.cap_res1.t20 bgr_0.cap_res1.t5 0.1603
R7409 bgr_0.cap_res1.t10 bgr_0.cap_res1.t20 0.1603
R7410 bgr_0.cap_res1.t3 bgr_0.cap_res1.t10 0.1603
R7411 bgr_0.cap_res1.t6 bgr_0.cap_res1.t17 0.1603
R7412 bgr_0.cap_res1.t13 bgr_0.cap_res1.t6 0.1603
R7413 bgr_0.cap_res1.t19 bgr_0.cap_res1.t13 0.1603
R7414 bgr_0.cap_res1.t4 bgr_0.cap_res1.t19 0.1603
R7415 bgr_0.cap_res1.t11 bgr_0.cap_res1.t4 0.1603
R7416 bgr_0.cap_res1.t15 bgr_0.cap_res1.t11 0.1603
R7417 bgr_0.cap_res1.t1 bgr_0.cap_res1.t15 0.1603
R7418 bgr_0.cap_res1.t8 bgr_0.cap_res1.t1 0.1603
R7419 bgr_0.cap_res1.t12 bgr_0.cap_res1.n0 0.159278
R7420 bgr_0.cap_res1.t17 bgr_0.cap_res1.t12 0.137822
R7421 bgr_0.cap_res1.n0 bgr_0.cap_res1.t3 0.1368
R7422 bgr_0.cap_res1.n0 bgr_0.cap_res1.t18 0.00152174
R7423 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 517.347
R7424 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R7425 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R7426 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 228.148
R7427 pfd_8_0.E_b.t2 pfd_8_0.E_b.n2 221.411
R7428 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R7429 pfd_8_0.E_b.n1 pfd_8_0.E_b.t1 24.0005
R7430 a_870_1390.t0 a_870_1390.t1 39.4005
R7431 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R7432 pfd_8_0.E.n0 pfd_8_0.E.t5 562.333
R7433 pfd_8_0.E.n2 pfd_8_0.E.t4 388.813
R7434 pfd_8_0.E.n2 pfd_8_0.E.t6 356.68
R7435 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R7436 pfd_8_0.E.n0 pfd_8_0.E.t3 224.934
R7437 pfd_8_0.E.t1 pfd_8_0.E.n4 221.411
R7438 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R7439 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R7440 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R7441 pfd_8_0.E.n1 pfd_8_0.E.t0 24.0005
R7442 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 710.734
R7443 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 553.534
R7444 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 254.333
R7445 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 206.333
R7446 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 70.4005
R7447 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 48.0005
R7448 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 48.0005
R7449 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 12.8005
R7450 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 663.801
R7451 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 514.134
R7452 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 479.284
R7453 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 344.8
R7454 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 289.2
R7455 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 275.454
R7456 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 241
R7457 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 112.468
R7458 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 97.9205
R7459 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 64.2672
R7460 VCO_FD_magic_0.div120_2_0.div2.t6 VCO_FD_magic_0.div120_2_0.div2.t4 1012.2
R7461 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t0 663.801
R7462 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n1 431.401
R7463 VCO_FD_magic_0.div120_2_0.div2.t5 VCO_FD_magic_0.div120_2_0.div2.t2 401.668
R7464 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t6 361.692
R7465 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t3 353.467
R7466 VCO_FD_magic_0.div120_2_0.div2.t1 VCO_FD_magic_0.div120_2_0.div2.n2 298.921
R7467 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t5 257.067
R7468 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n0 67.2005
R7469 a_7630_n1530.n0 a_7630_n1530.t1 752.333
R7470 a_7630_n1530.t2 a_7630_n1530.n5 752.333
R7471 a_7630_n1530.n1 a_7630_n1530.t6 514.134
R7472 a_7630_n1530.n4 a_7630_n1530.n3 366.856
R7473 a_7630_n1530.n0 a_7630_n1530.t0 254.333
R7474 a_7630_n1530.n4 a_7630_n1530.t3 190.123
R7475 a_7630_n1530.n5 a_7630_n1530.n4 187.201
R7476 a_7630_n1530.n3 a_7630_n1530.n2 176.733
R7477 a_7630_n1530.n2 a_7630_n1530.n1 176.733
R7478 a_7630_n1530.n3 a_7630_n1530.t7 112.468
R7479 a_7630_n1530.n2 a_7630_n1530.t4 112.468
R7480 a_7630_n1530.n1 a_7630_n1530.t5 112.468
R7481 a_7630_n1530.n5 a_7630_n1530.n0 70.4005
R7482 pfd_8_0.UP.n0 pfd_8_0.UP.t3 1205
R7483 pfd_8_0.UP.n2 pfd_8_0.UP.t2 522.168
R7484 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R7485 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R7486 pfd_8_0.UP.t0 pfd_8_0.UP.n3 229.127
R7487 pfd_8_0.UP.n1 pfd_8_0.UP.t5 217.905
R7488 pfd_8_0.UP.n0 pfd_8_0.UP.t4 208.868
R7489 pfd_8_0.UP.n3 pfd_8_0.UP.t1 158.335
R7490 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R7491 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 501.467
R7492 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R7493 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R7494 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 209.928
R7495 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t1 177.536
R7496 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t0 19.5223
R7497 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t3 326.658
R7498 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t6 297.233
R7499 pfd_8_0.UP_input.t5 pfd_8_0.UP_input.n5 297.233
R7500 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n1 257.067
R7501 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 242.494
R7502 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t2 241.928
R7503 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n1 226.942
R7504 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 226.942
R7505 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n4 216.9
R7506 pfd_8_0.UP_input.t1 pfd_8_0.UP_input.n7 209.928
R7507 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t0 145.536
R7508 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n0 144
R7509 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t6 92.3838
R7510 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t5 92.3838
R7511 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t7 80.3338
R7512 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n3 80.3338
R7513 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t4 80.3338
R7514 pfd_8_0.UP_input.t4 pfd_8_0.UP_input.n1 80.3338
R7515 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R7516 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R7517 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R7518 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R7519 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R7520 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R7521 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R7522 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R7523 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R7524 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R7525 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R7526 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R7527 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R7528 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R7529 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R7530 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R7531 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R7532 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R7533 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R7534 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R7535 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R7536 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R7537 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R7538 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R7539 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R7540 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R7541 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R7542 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R7543 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R7544 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R7545 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R7546 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R7547 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R7548 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R7549 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R7550 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R7551 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R7552 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 65.0299
R7553 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R7554 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R7555 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R7556 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R7557 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R7558 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R7559 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R7560 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R7561 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R7562 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R7563 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R7564 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R7565 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R7566 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 25.7843
R7567 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R7568 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7569 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7570 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7571 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7572 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7573 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7574 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7575 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R7576 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7577 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7578 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7579 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7580 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R7581 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R7582 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7583 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7584 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7585 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7586 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7587 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7588 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7589 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7590 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7591 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7592 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7593 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R7594 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R7595 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R7596 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7597 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7598 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7599 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R7600 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7601 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7602 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7603 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R7604 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7605 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7606 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7607 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7608 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7609 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7610 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7611 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7612 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7613 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7614 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7615 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7616 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R7617 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R7618 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7619 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7620 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7621 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7622 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R7623 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R7624 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R7625 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R7626 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R7627 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R7628 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R7629 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R7630 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R7631 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R7632 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R7633 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R7634 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R7635 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R7636 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R7637 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R7638 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R7639 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R7640 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R7641 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R7642 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R7643 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R7644 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R7645 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R7646 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R7647 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R7648 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R7649 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R7650 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R7651 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R7652 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R7653 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R7654 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R7655 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R7656 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R7657 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R7658 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R7659 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R7660 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R7661 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R7662 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R7663 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R7664 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R7665 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R7666 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R7667 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R7668 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R7669 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R7670 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R7671 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R7672 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R7673 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R7674 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R7675 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R7676 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R7677 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R7678 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R7679 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R7680 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R7681 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R7682 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R7683 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R7684 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R7685 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R7686 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R7687 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R7688 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R7689 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R7690 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R7691 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R7692 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R7693 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R7694 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R7695 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R7696 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R7697 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R7698 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R7699 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R7700 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R7701 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R7702 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7703 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R7704 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R7705 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7706 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R7707 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7708 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R7709 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R7710 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R7711 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R7712 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R7713 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R7714 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R7715 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R7716 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R7717 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R7718 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R7719 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R7720 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R7721 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R7722 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R7723 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 0.290206
R7724 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R7725 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R7726 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R7727 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R7728 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R7729 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R7730 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R7731 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7732 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7733 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7734 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R7735 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7736 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R7737 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R7738 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R7739 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R7740 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R7741 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R7742 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R7743 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R7744 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R7745 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R7746 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R7747 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R7748 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R7749 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R7750 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R7751 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R7752 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R7753 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R7754 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R7755 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R7756 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R7757 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R7758 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R7759 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R7760 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R7761 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R7762 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R7763 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R7764 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R7765 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R7766 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R7767 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R7768 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R7769 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R7770 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R7771 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R7772 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R7773 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R7774 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R7775 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R7776 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R7777 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R7778 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R7779 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R7780 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R7781 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R7782 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R7783 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R7784 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R7785 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R7786 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R7787 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R7788 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R7789 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t5 600.206
R7790 VCO_FD_magic_0.vco2_3_0.V1.t2 VCO_FD_magic_0.vco2_3_0.V1.n5 576.192
R7791 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.n1 568.072
R7792 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n2 392.486
R7793 VCO_FD_magic_0.vco2_3_0.V1.n0 VCO_FD_magic_0.vco2_3_0.V1.t1 289.791
R7794 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n4 168.067
R7795 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.n0 97.9242
R7796 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n3 37.7572
R7797 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t3 32.1338
R7798 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.t4 32.1338
R7799 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.t0 32.1338
R7800 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n0 28.3357
R7801 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t1 421.027
R7802 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t2 348.81
R7803 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.t0 280.05
R7804 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.n0 36.1094
R7805 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 424.447
R7806 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 354.048
R7807 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 313
R7808 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.t14 297.233
R7809 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t14 297.233
R7810 pfd_8_0.opamp_out.t13 pfd_8_0.opamp_out.n11 297.233
R7811 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t6 281.596
R7812 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n0 242.601
R7813 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n2 220.8
R7814 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.n6 220.8
R7815 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n12 218.857
R7816 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.n10 216.9
R7817 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 216.9
R7818 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.n8 184.768
R7819 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t5 118.666
R7820 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 80.3338
R7821 pfd_8_0.opamp_out.t15 pfd_8_0.opamp_out.n9 80.3338
R7822 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t10 80.3338
R7823 pfd_8_0.opamp_out.t10 pfd_8_0.opamp_out.n8 80.3338
R7824 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t13 80.3338
R7825 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 73.0531
R7826 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 70.0829
R7827 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t11 63.6829
R7828 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 62.7569
R7829 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n3 62.4005
R7830 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n7 60.8005
R7831 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t1 60.0005
R7832 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t3 60.0005
R7833 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t4 60.0005
R7834 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t9 60.0005
R7835 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t2 49.2505
R7836 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t7 49.2505
R7837 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t0 49.2505
R7838 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t8 49.2505
R7839 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 1.6005
R7840 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t8 377.567
R7841 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t6 321.334
R7842 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 233.476
R7843 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t7 216.9
R7844 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 199.462
R7845 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 189.898
R7846 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R7847 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R7848 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t9 112.468
R7849 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R7850 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 57.2776
R7851 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R7852 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t0 24.6255
R7853 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t3 24.6255
R7854 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t2 24.6255
R7855 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R7856 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t4 15.0005
R7857 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.20883
R7858 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 359.894
R7859 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R7860 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R7861 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t0 252.248
R7862 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R7863 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R7864 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R7865 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R7866 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t5 60.0005
R7867 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t4 60.0005
R7868 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R7869 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R7870 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t1 49.2505
R7871 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_right.n6 1010.36
R7872 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 404.8
R7873 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 322.048
R7874 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 316.2
R7875 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R7876 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R7877 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R7878 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 232.968
R7879 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R7880 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R7881 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 199.829
R7882 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t2 60.0005
R7883 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t3 60.0005
R7884 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t0 49.2505
R7885 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t1 49.2505
R7886 a_6320_5840.n7 a_6320_5840.n5 482.582
R7887 a_6320_5840.n10 a_6320_5840.t5 304.634
R7888 a_6320_5840.n3 a_6320_5840.t3 304.634
R7889 a_6320_5840.t7 a_6320_5840.n10 277.914
R7890 a_6320_5840.n3 a_6320_5840.t4 276.289
R7891 a_6320_5840.n8 a_6320_5840.n1 204.201
R7892 a_6320_5840.n4 a_6320_5840.n2 204.201
R7893 a_6320_5840.n9 a_6320_5840.n0 204.201
R7894 a_6320_5840.n7 a_6320_5840.n6 120.981
R7895 a_6320_5840.n8 a_6320_5840.n4 74.6672
R7896 a_6320_5840.n9 a_6320_5840.n8 74.6672
R7897 a_6320_5840.n1 a_6320_5840.t9 60.0005
R7898 a_6320_5840.n1 a_6320_5840.t11 60.0005
R7899 a_6320_5840.t4 a_6320_5840.n2 60.0005
R7900 a_6320_5840.n2 a_6320_5840.t8 60.0005
R7901 a_6320_5840.n0 a_6320_5840.t10 60.0005
R7902 a_6320_5840.n0 a_6320_5840.t6 60.0005
R7903 a_6320_5840.n8 a_6320_5840.n7 37.763
R7904 a_6320_5840.n5 a_6320_5840.t1 24.0005
R7905 a_6320_5840.n5 a_6320_5840.t12 24.0005
R7906 a_6320_5840.n6 a_6320_5840.t0 24.0005
R7907 a_6320_5840.n6 a_6320_5840.t2 24.0005
R7908 a_6320_5840.n4 a_6320_5840.n3 16.0005
R7909 a_6320_5840.n10 a_6320_5840.n9 16.0005
R7910 VCO_FD_magic_0.div120_2_0.div8.t5 VCO_FD_magic_0.div120_2_0.div8.t2 1012.2
R7911 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t1 663.801
R7912 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n1 431.401
R7913 VCO_FD_magic_0.div120_2_0.div8.t4 VCO_FD_magic_0.div120_2_0.div8.t6 401.668
R7914 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t5 361.692
R7915 VCO_FD_magic_0.div120_2_0.div8.t0 VCO_FD_magic_0.div120_2_0.div8.n2 298.921
R7916 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t4 257.067
R7917 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t3 208.868
R7918 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n0 67.2005
R7919 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 96.0005
R7920 a_6490_4630.t0 a_6490_4630.n6 1112.76
R7921 a_6490_4630.n3 a_6490_4630.n2 441.433
R7922 a_6490_4630.n2 a_6490_4630.n1 379.647
R7923 a_6490_4630.n2 a_6490_4630.n0 258.601
R7924 a_6490_4630.n6 a_6490_4630.t6 208.868
R7925 a_6490_4630.n5 a_6490_4630.t7 208.868
R7926 a_6490_4630.n4 a_6490_4630.t8 208.868
R7927 a_6490_4630.n3 a_6490_4630.t5 208.868
R7928 a_6490_4630.n6 a_6490_4630.n5 208.868
R7929 a_6490_4630.n5 a_6490_4630.n4 208.868
R7930 a_6490_4630.n4 a_6490_4630.n3 208.868
R7931 a_6490_4630.n0 a_6490_4630.t4 60.0005
R7932 a_6490_4630.n0 a_6490_4630.t3 60.0005
R7933 a_6490_4630.n1 a_6490_4630.t2 49.2505
R7934 a_6490_4630.n1 a_6490_4630.t1 49.2505
R7935 bgr_0.V_mir1.n15 bgr_0.V_mir1.t22 310.488
R7936 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 310.488
R7937 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 310.488
R7938 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 297.433
R7939 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 297.433
R7940 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 297.433
R7941 bgr_0.V_mir1.n7 bgr_0.V_mir1.t3 248.133
R7942 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 199.383
R7943 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 194.883
R7944 bgr_0.V_mir1.n17 bgr_0.V_mir1.t9 184.097
R7945 bgr_0.V_mir1.n11 bgr_0.V_mir1.t7 184.097
R7946 bgr_0.V_mir1.n2 bgr_0.V_mir1.t5 184.097
R7947 bgr_0.V_mir1.n16 bgr_0.V_mir1.n15 167.094
R7948 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7949 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7950 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 161.3
R7951 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 161.3
R7952 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 161.3
R7953 bgr_0.V_mir1.n15 bgr_0.V_mir1.t19 120.501
R7954 bgr_0.V_mir1.n16 bgr_0.V_mir1.t15 120.501
R7955 bgr_0.V_mir1.n9 bgr_0.V_mir1.t20 120.501
R7956 bgr_0.V_mir1.n10 bgr_0.V_mir1.t13 120.501
R7957 bgr_0.V_mir1.n0 bgr_0.V_mir1.t21 120.501
R7958 bgr_0.V_mir1.n1 bgr_0.V_mir1.t11 120.501
R7959 bgr_0.V_mir1.n6 bgr_0.V_mir1.t1 48.0005
R7960 bgr_0.V_mir1.n6 bgr_0.V_mir1.t0 48.0005
R7961 bgr_0.V_mir1.n5 bgr_0.V_mir1.t4 48.0005
R7962 bgr_0.V_mir1.n5 bgr_0.V_mir1.t2 48.0005
R7963 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 40.7027
R7964 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7965 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7966 bgr_0.V_mir1.n12 bgr_0.V_mir1.t8 39.4005
R7967 bgr_0.V_mir1.n12 bgr_0.V_mir1.t14 39.4005
R7968 bgr_0.V_mir1.n3 bgr_0.V_mir1.t6 39.4005
R7969 bgr_0.V_mir1.n3 bgr_0.V_mir1.t12 39.4005
R7970 bgr_0.V_mir1.n19 bgr_0.V_mir1.t10 39.4005
R7971 bgr_0.V_mir1.t16 bgr_0.V_mir1.n19 39.4005
R7972 bgr_0.V_mir1.n14 bgr_0.V_mir1.n4 6.6255
R7973 bgr_0.V_mir1.n18 bgr_0.V_mir1.n14 6.6255
R7974 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.2505
R7975 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 4.5005
R7976 bgr_0.V_mir1.n13 bgr_0.V_mir1.n8 0.78175
R7977 a_3280_11518.t0 a_3280_11518.t1 178.133
R7978 bgr_0.Vin-.n14 bgr_0.Vin-.n13 314.526
R7979 bgr_0.Vin-.n16 bgr_0.Vin-.t8 287.762
R7980 bgr_0.Vin-.n17 bgr_0.Vin-.t9 287.762
R7981 bgr_0.Vin-.n16 bgr_0.Vin-.t10 287.589
R7982 bgr_0.Vin-.n18 bgr_0.Vin-.t11 287.012
R7983 bgr_0.Vin-.n19 bgr_0.Vin-.t12 287.012
R7984 bgr_0.Vin-.n9 bgr_0.Vin-.t1 117.817
R7985 bgr_0.Vin-.n12 bgr_0.Vin-.n10 107.079
R7986 bgr_0.Vin-.n12 bgr_0.Vin-.n11 104.829
R7987 bgr_0.Vin-.n3 bgr_0.Vin-.n2 83.5719
R7988 bgr_0.Vin-.n5 bgr_0.Vin-.n4 83.5719
R7989 bgr_0.Vin-.n4 bgr_0.Vin-.n1 73.8495
R7990 bgr_0.Vin-.t3 bgr_0.Vin-.n0 65.0341
R7991 bgr_0.Vin-.n13 bgr_0.Vin-.t0 39.4005
R7992 bgr_0.Vin-.n13 bgr_0.Vin-.t2 39.4005
R7993 bgr_0.Vin-.n4 bgr_0.Vin-.n3 26.074
R7994 bgr_0.Vin-.n9 bgr_0.Vin-.n8 23.9067
R7995 bgr_0.Vin-.n10 bgr_0.Vin-.t6 13.1338
R7996 bgr_0.Vin-.n10 bgr_0.Vin-.t7 13.1338
R7997 bgr_0.Vin-.n11 bgr_0.Vin-.t4 13.1338
R7998 bgr_0.Vin-.n11 bgr_0.Vin-.t5 13.1338
R7999 bgr_0.Vin-.n15 bgr_0.Vin-.n9 13.0943
R8000 bgr_0.Vin-.n15 bgr_0.Vin-.n14 10.7505
R8001 bgr_0.Vin- bgr_0.Vin-.n15 4.813
R8002 bgr_0.Vin-.n14 bgr_0.Vin-.n12 2.0005
R8003 bgr_0.Vin- bgr_0.Vin-.n19 1.96836
R8004 bgr_0.Vin-.n2 bgr_0.Vin-.n0 1.56483
R8005 bgr_0.Vin-.n7 bgr_0.Vin-.n6 1.5505
R8006 bgr_0.Vin-.n6 bgr_0.Vin-.n5 0.885803
R8007 bgr_0.Vin-.n6 bgr_0.Vin-.n2 0.77514
R8008 bgr_0.Vin-.n5 bgr_0.Vin- 0.756696
R8009 bgr_0.Vin-.n7 bgr_0.Vin-.n1 0.711459
R8010 bgr_0.Vin-.n18 bgr_0.Vin-.n17 0.579071
R8011 bgr_0.Vin- bgr_0.Vin-.n1 0.576566
R8012 bgr_0.Vin-.n8 bgr_0.Vin-.n0 0.531499
R8013 bgr_0.Vin-.n3 bgr_0.Vin-.t3 0.290206
R8014 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.282643
R8015 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.2755
R8016 bgr_0.Vin-.n8 bgr_0.Vin-.n7 0.00817857
R8017 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 755.534
R8018 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 685.134
R8019 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 389.733
R8020 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 340.2
R8021 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 321.334
R8022 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 144.601
R8023 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 19.2005
R8024 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 713.933
R8025 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 327.401
R8026 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 314.233
R8027 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 9.6005
R8028 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t8 918.318
R8029 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R8030 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R8031 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R8032 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R8033 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R8034 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R8035 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R8036 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R8037 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R8038 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R8039 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R8040 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t4 120.501
R8041 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t0 120.501
R8042 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t2 120.501
R8043 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R8044 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t6 120.501
R8045 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R8046 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R8047 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R8048 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R8049 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R8050 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t1 19.7005
R8051 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t5 19.7005
R8052 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t7 19.7005
R8053 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t3 19.7005
R8054 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 723
R8055 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 514.134
R8056 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 332.783
R8057 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 314.921
R8058 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 6.4005
R8059 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 3.2005
R8060 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 157.601
R8061 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 96.0005
R8062 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t3 1188.93
R8063 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R8064 pfd_8_0.QA_b.t3 pfd_8_0.QA_b.t5 835.467
R8065 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t6 562.333
R8066 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R8067 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R8068 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R8069 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t0 221.411
R8070 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t1 24.0005
R8071 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R8072 bgr_0.V_CUR_REF_REG.n6 bgr_0.V_CUR_REF_REG.n4 302.507
R8073 bgr_0.V_CUR_REF_REG.n14 bgr_0.V_CUR_REF_REG.n13 302.163
R8074 bgr_0.V_CUR_REF_REG.n12 bgr_0.V_CUR_REF_REG.n11 302.163
R8075 bgr_0.V_CUR_REF_REG.n10 bgr_0.V_CUR_REF_REG.n9 302.163
R8076 bgr_0.V_CUR_REF_REG.n8 bgr_0.V_CUR_REF_REG.n7 302.163
R8077 bgr_0.V_CUR_REF_REG.n6 bgr_0.V_CUR_REF_REG.n5 302.163
R8078 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t15 291.502
R8079 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t16 291.288
R8080 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t13 291.288
R8081 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t17 291.288
R8082 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t14 291.288
R8083 bgr_0.V_CUR_REF_REG.n15 bgr_0.V_CUR_REF_REG.t12 133.005
R8084 bgr_0.V_CUR_REF_REG.n13 bgr_0.V_CUR_REF_REG.t1 39.4005
R8085 bgr_0.V_CUR_REF_REG.n13 bgr_0.V_CUR_REF_REG.t11 39.4005
R8086 bgr_0.V_CUR_REF_REG.n11 bgr_0.V_CUR_REF_REG.t0 39.4005
R8087 bgr_0.V_CUR_REF_REG.n11 bgr_0.V_CUR_REF_REG.t5 39.4005
R8088 bgr_0.V_CUR_REF_REG.n9 bgr_0.V_CUR_REF_REG.t2 39.4005
R8089 bgr_0.V_CUR_REF_REG.n9 bgr_0.V_CUR_REF_REG.t4 39.4005
R8090 bgr_0.V_CUR_REF_REG.n7 bgr_0.V_CUR_REF_REG.t9 39.4005
R8091 bgr_0.V_CUR_REF_REG.n7 bgr_0.V_CUR_REF_REG.t7 39.4005
R8092 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.t3 39.4005
R8093 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.t6 39.4005
R8094 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t10 39.4005
R8095 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t8 39.4005
R8096 bgr_0.V_CUR_REF_REG.n15 bgr_0.V_CUR_REF_REG.n14 12.0474
R8097 bgr_0.V_CUR_REF_REG bgr_0.V_CUR_REF_REG.n15 4.72371
R8098 bgr_0.V_CUR_REF_REG bgr_0.V_CUR_REF_REG.n3 1.67729
R8099 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 0.643357
R8100 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 0.643357
R8101 bgr_0.V_CUR_REF_REG.n8 bgr_0.V_CUR_REF_REG.n6 0.34425
R8102 bgr_0.V_CUR_REF_REG.n10 bgr_0.V_CUR_REF_REG.n8 0.34425
R8103 bgr_0.V_CUR_REF_REG.n12 bgr_0.V_CUR_REF_REG.n10 0.34425
R8104 bgr_0.V_CUR_REF_REG.n14 bgr_0.V_CUR_REF_REG.n12 0.34425
R8105 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 0.214786
R8106 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 713.933
R8107 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 314.233
R8108 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 308.2
R8109 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 702.201
R8110 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 350.349
R8111 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 276.733
R8112 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 206.333
R8113 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 48.0005
R8114 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 48.0005
R8115 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 48.0005
R8116 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 19.2005
R8117 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 713.933
R8118 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 327.401
R8119 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 314.233
R8120 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 9.6005
R8121 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 702.201
R8122 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 349.433
R8123 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 276.733
R8124 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 206.333
R8125 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 48.0005
R8126 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 48.0005
R8127 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 48.0005
R8128 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 48.0005
R8129 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 742.51
R8130 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 723.534
R8131 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 723.534
R8132 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 684.806
R8133 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 366.856
R8134 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 337.401
R8135 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 305.267
R8136 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 254.333
R8137 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 224.934
R8138 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 190.123
R8139 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 187.201
R8140 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 176.733
R8141 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 176.733
R8142 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 176.733
R8143 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 144.601
R8144 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 131.976
R8145 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 128.534
R8146 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 128.534
R8147 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 112.468
R8148 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 112.468
R8149 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 112.468
R8150 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 70.4005
R8151 a_8930_n1530.n4 a_8930_n1530.t1 752.333
R8152 a_8930_n1530.t2 a_8930_n1530.n5 752.333
R8153 a_8930_n1530.n0 a_8930_n1530.t5 514.134
R8154 a_8930_n1530.n3 a_8930_n1530.n2 366.856
R8155 a_8930_n1530.n5 a_8930_n1530.t0 254.333
R8156 a_8930_n1530.n3 a_8930_n1530.t7 190.123
R8157 a_8930_n1530.n4 a_8930_n1530.n3 187.201
R8158 a_8930_n1530.n2 a_8930_n1530.n1 176.733
R8159 a_8930_n1530.n1 a_8930_n1530.n0 176.733
R8160 a_8930_n1530.n2 a_8930_n1530.t4 112.468
R8161 a_8930_n1530.n1 a_8930_n1530.t6 112.468
R8162 a_8930_n1530.n0 a_8930_n1530.t3 112.468
R8163 a_8930_n1530.n5 a_8930_n1530.n4 70.4005
R8164 F_VCO.n1 F_VCO.t6 772.196
R8165 F_VCO.n3 F_VCO.t1 751.801
R8166 F_VCO.n2 F_VCO.n1 607.465
R8167 F_VCO.t6 F_VCO.t3 514.134
R8168 F_VCO.n4 F_VCO.t2 514.134
R8169 F_VCO.n0 F_VCO.t5 289.2
R8170 F_VCO.n4 F_VCO.t4 273.134
R8171 F_VCO.n2 F_VCO.t0 233
R8172 F_VCO F_VCO.n4 216.9
R8173 F_VCO.n1 F_VCO.n0 208.868
R8174 F_VCO F_VCO.n5 187.053
R8175 F_VCO.n0 F_VCO.t7 176.733
R8176 F_VCO.n3 F_VCO.n2 40.3205
R8177 F_VCO F_VCO.n3 38.4005
R8178 F_VCO.n5 F_VCO 24.1005
R8179 F_VCO.n5 F_VCO 24.1005
R8180 a_6220_5810.n4 a_6220_5810.t12 317.317
R8181 a_6220_5810.n2 a_6220_5810.t11 317.317
R8182 a_6220_5810.n5 a_6220_5810.n4 257.067
R8183 a_6220_5810.n3 a_6220_5810.n2 257.067
R8184 a_6220_5810.n10 a_6220_5810.n9 257.067
R8185 a_6220_5810.t0 a_6220_5810.n12 194.478
R8186 a_6220_5810.n8 a_6220_5810.n7 152
R8187 a_6220_5810.n12 a_6220_5810.n11 152
R8188 a_6220_5810.n1 a_6220_5810.n0 120.981
R8189 a_6220_5810.n7 a_6220_5810.n6 117.781
R8190 a_6220_5810.n7 a_6220_5810.n1 108.8
R8191 a_6220_5810.n8 a_6220_5810.n5 85.6894
R8192 a_6220_5810.n11 a_6220_5810.n3 85.6894
R8193 a_6220_5810.n11 a_6220_5810.n10 85.6894
R8194 a_6220_5810.n9 a_6220_5810.n8 85.6894
R8195 a_6220_5810.n4 a_6220_5810.t10 60.2505
R8196 a_6220_5810.n5 a_6220_5810.t1 60.2505
R8197 a_6220_5810.n2 a_6220_5810.t9 60.2505
R8198 a_6220_5810.n3 a_6220_5810.t3 60.2505
R8199 a_6220_5810.n10 a_6220_5810.t7 60.2505
R8200 a_6220_5810.n9 a_6220_5810.t5 60.2505
R8201 a_6220_5810.n6 a_6220_5810.t6 24.0005
R8202 a_6220_5810.n6 a_6220_5810.t2 24.0005
R8203 a_6220_5810.n0 a_6220_5810.t4 24.0005
R8204 a_6220_5810.n0 a_6220_5810.t8 24.0005
R8205 a_6220_5810.n12 a_6220_5810.n1 3.2005
R8206 a_n1130_7570.n0 a_n1130_7570.t6 238.322
R8207 a_n1130_7570.n0 a_n1130_7570.t7 238.322
R8208 a_n1130_7570.n4 a_n1130_7570.n0 168.8
R8209 a_n1130_7570.n1 a_n1130_7570.t1 130.001
R8210 a_n1130_7570.n3 a_n1130_7570.n2 105.171
R8211 a_n1130_7570.n5 a_n1130_7570.n4 105.171
R8212 a_n1130_7570.n1 a_n1130_7570.t0 81.7085
R8213 a_n1130_7570.n3 a_n1130_7570.n1 46.5739
R8214 a_n1130_7570.n2 a_n1130_7570.t4 13.1338
R8215 a_n1130_7570.n2 a_n1130_7570.t2 13.1338
R8216 a_n1130_7570.t5 a_n1130_7570.n5 13.1338
R8217 a_n1130_7570.n5 a_n1130_7570.t3 13.1338
R8218 a_n1130_7570.n4 a_n1130_7570.n3 3.3755
R8219 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 96.0005
R8220 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 685.134
R8221 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 663.801
R8222 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 534.268
R8223 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 340.521
R8224 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 105.6
R8225 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 21.3338
R8226 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 279.933
R8227 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 251.133
R8228 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 48.0005
R8229 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 48.0005
R8230 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 96.0005
R8231 a_2200_180.t1 a_2200_180.n2 500.086
R8232 a_2200_180.n1 a_2200_180.n0 473.334
R8233 a_2200_180.n0 a_2200_180.t2 465.933
R8234 a_2200_180.t1 a_2200_180.n2 461.389
R8235 a_2200_180.n0 a_2200_180.t3 321.334
R8236 a_2200_180.n1 a_2200_180.t0 177.577
R8237 a_2200_180.n2 a_2200_180.n1 48.3898
R8238 a_1870_180.t1 a_1870_180.n2 500.086
R8239 a_1870_180.n1 a_1870_180.n0 473.334
R8240 a_1870_180.n0 a_1870_180.t2 465.933
R8241 a_1870_180.t1 a_1870_180.n2 461.389
R8242 a_1870_180.n0 a_1870_180.t3 321.334
R8243 a_1870_180.n1 a_1870_180.t0 177.577
R8244 a_1870_180.n2 a_1870_180.n1 48.3898
R8245 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 702.201
R8246 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 349.433
R8247 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 276.733
R8248 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 206.333
R8249 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 48.0005
R8250 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 48.0005
R8251 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 48.0005
R8252 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 48.0005
R8253 F_REF.n0 F_REF.t1 514.134
R8254 F_REF.n0 F_REF.t0 273.134
R8255 F_REF F_REF.n0 216.9
R8256 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 685.134
R8257 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 663.801
R8258 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 534.268
R8259 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 362.921
R8260 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 91.7338
R8261 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 701.467
R8262 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 694.201
R8263 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 321.334
R8264 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 260.521
R8265 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 144.601
R8266 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 54.4005
R8267 a_490_630.t0 a_490_630.t1 39.4005
R8268 a_1390_1390.t0 a_1390_1390.t1 39.4005
R8269 a_9360_3514.t1 a_9360_3514.t0 323.964
R8270 loop_filter_2_0.R1_C1.t1 loop_filter_2_0.R1_C1.t0 167.429
R8271 a_2350_1390.t0 a_2350_1390.n2 500.086
R8272 a_2350_1390.n1 a_2350_1390.n0 473.334
R8273 a_2350_1390.n0 a_2350_1390.t2 465.933
R8274 a_2350_1390.t0 a_2350_1390.n2 461.389
R8275 a_2350_1390.n0 a_2350_1390.t3 321.334
R8276 a_2350_1390.n1 a_2350_1390.t1 177.577
R8277 a_2350_1390.n2 a_2350_1390.n1 48.3899
R8278 a_2530_180.t1 a_2530_180.n2 500.086
R8279 a_2530_180.n0 a_2530_180.t2 465.933
R8280 a_2530_180.t1 a_2530_180.n2 461.389
R8281 a_2530_180.n1 a_2530_180.n0 392.623
R8282 a_2530_180.n0 a_2530_180.t3 321.334
R8283 a_2530_180.n1 a_2530_180.t0 177.577
R8284 a_2530_180.n2 a_2530_180.n1 48.3899
R8285 a_n1490_9910.t0 a_n1490_9910.t1 178.133
R8286 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 702.201
R8287 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 349.433
R8288 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 276.733
R8289 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 206.333
R8290 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 48.0005
R8291 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 48.0005
R8292 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 48.0005
R8293 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 48.0005
R8294 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R8295 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t2 203.528
R8296 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R8297 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 183.935
R8298 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R8299 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.n0 437.733
R8300 VCO_FD_magic_0.vco2_3_0.V8.t0 VCO_FD_magic_0.vco2_3_0.V8.n1 372.118
R8301 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.t1 247.934
R8302 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t3 224.934
R8303 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t2 144.601
R8304 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t0 284.2
R8305 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t2 233
R8306 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.t1 162.857
R8307 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.n0 21.3338
R8308 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 742.201
R8309 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 350.349
R8310 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 254.333
R8311 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 206.333
R8312 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 70.4005
R8313 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 48.0005
R8314 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 48.0005
R8315 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 19.2005
R8316 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 199.935
R8317 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 199.53
R8318 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 199.53
R8319 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 199.53
R8320 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 199.53
R8321 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 55.1744
R8322 bgr_0.V_p_1.n5 bgr_0.V_p_1.t7 48.0005
R8323 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R8324 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8325 bgr_0.V_p_1.n4 bgr_0.V_p_1.t3 48.0005
R8326 bgr_0.V_p_1.n3 bgr_0.V_p_1.t1 48.0005
R8327 bgr_0.V_p_1.n3 bgr_0.V_p_1.t8 48.0005
R8328 bgr_0.V_p_1.n2 bgr_0.V_p_1.t5 48.0005
R8329 bgr_0.V_p_1.n2 bgr_0.V_p_1.t0 48.0005
R8330 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8331 bgr_0.V_p_1.n6 bgr_0.V_p_1.t6 48.0005
R8332 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.09425
R8333 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 441.834
R8334 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 313.3
R8335 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R8336 pfd_8_0.UP_PFD_b.t0 pfd_8_0.UP_PFD_b.n1 219.528
R8337 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t1 167.935
R8338 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 96.0005
R8339 a_n2040_11368.t0 a_n2040_11368.t1 178.133
R8340 a_n1920_10290.t0 a_n1920_10290.t1 178.133
R8341 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 739
R8342 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 349.433
R8343 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 254.333
R8344 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 206.333
R8345 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 70.4005
R8346 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 48.0005
R8347 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 48.0005
R8348 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 22.4005
R8349 a_9360_6440.t0 a_9360_6440.t1 245.883
R8350 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 96.0005
R8351 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R8352 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R8353 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R8354 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R8355 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R8356 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R8357 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R8358 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R8359 a_3160_9910.t0 a_3160_9910.t1 178.133
R8360 bgr_0.START_UP_NFET1.t1 bgr_0.START_UP_NFET1.t0 178.194
R8361 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R8362 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 403.997
R8363 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 240.327
R8364 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 148.736
R8365 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t2 19.987
R8366 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t0 284.2
R8367 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t2 233
R8368 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.t1 162.857
R8369 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.n0 21.3338
R8370 pfd_8_0.QA.t7 pfd_8_0.QA.t3 835.467
R8371 pfd_8_0.QA.n2 pfd_8_0.QA.t6 517.347
R8372 pfd_8_0.QA.n0 pfd_8_0.QA.t4 465.933
R8373 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R8374 pfd_8_0.QA.n1 pfd_8_0.QA.t7 394.267
R8375 pfd_8_0.QA.n0 pfd_8_0.QA.t8 321.334
R8376 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R8377 pfd_8_0.QA.n2 pfd_8_0.QA.t5 228.148
R8378 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R8379 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R8380 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R8381 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R8382 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R8383 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R8384 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R8385 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R8386 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R8387 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R8388 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R8389 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t0 172.458
R8390 pfd_8_0.before_Reset.t1 pfd_8_0.before_Reset.n2 19.7005
R8391 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R8392 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t0 284.2
R8393 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t2 233
R8394 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.t1 162.857
R8395 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.n0 21.3338
R8396 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t0 421.027
R8397 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t2 348.81
R8398 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.t1 284.317
R8399 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.n0 31.8427
R8400 a_n1610_11518.t0 a_n1610_11518.t1 178.133
R8401 a_490_1390.t0 a_490_1390.t1 39.4005
R8402 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 663.801
R8403 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 397.053
R8404 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 348.851
R8405 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN_input.t4 377.567
R8406 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t3 326.658
R8407 pfd_8_0.DOWN_input.n4 pfd_8_0.DOWN_input.n1 242.744
R8408 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t0 229.127
R8409 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 196.817
R8410 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t1 164.736
R8411 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t2 158.335
R8412 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 118.4
R8413 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n0 92.3838
R8414 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t5 92.3838
R8415 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n4 9.6005
R8416 pfd_8_0.DOWN_input.n4 pfd_8_0.DOWN_input.n3 9.6005
R8417 a_1910_2010.t0 a_1910_2010.t1 48.0005
R8418 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 96.0005
R8419 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 96.0005
R8420 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 713.933
R8421 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 327.401
R8422 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 314.233
R8423 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 9.6005
R8424 a_870_630.t0 a_870_630.t1 39.4005
R8425 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 663.801
R8426 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 355.378
R8427 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 276.521
R8428 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 120.534
R8429 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 96.0005
R8430 a_n30_1390.t0 a_n30_1390.t1 39.4005
C0 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div24 0.240642f
C1 pfd_8_0.QA_b F_REF 0.037629f
C2 VCO_FD_magic_0.vco2_3_0.V6 V_OSC 0.019495f
C3 bgr_0.V_TOP VDDA 16.1936f
C4 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div24 0.076865f
C5 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.D 0.163145f
C6 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div24 0.03648f
C7 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.108607f
C8 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div24 0.024014f
C9 VCO_FD_magic_0.div120_2_0.div2_4_1.A VDDA 0.126015f
C10 VCO_FD_magic_0.vco2_3_0.V6 VDDA 0.281338f
C11 VCO_FD_magic_0.vco2_3_0.V2 V_OSC 0.063469f
C12 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.176046f
C13 bgr_0.Vin- bgr_0.V_CUR_REF_REG 0.83728f
C14 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.Vin- 1.05523f
C15 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.169071f
C16 bgr_0.V2 F_REF 0.011728f
C17 VCO_FD_magic_0.div120_2_0.div2_4_2.A VDDA 0.125335f
C18 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div24 0.038583f
C19 F_VCO VDDA 1.24152f
C20 bgr_0.V_TOP bgr_0.Vin+ 2.13503f
C21 VCO_FD_magic_0.vco2_3_0.V2 VDDA 0.410554f
C22 bgr_0.Vin- bgr_0.1st_Vout_1 0.677227f
C23 VCO_FD_magic_0.div120_2_0.div2_4_0.A VDDA 0.125335f
C24 pfd_8_0.QB VDDA 2.75031f
C25 opamp_cell_4_0.VIN+ pfd_8_0.DOWN_input 0.044605f
C26 bgr_0.V_TOP bgr_0.V2 0.351781f
C27 VDDA pfd_8_0.DOWN_input 0.191914f
C28 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.G 0.081976f
C29 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V7 0.010316f
C30 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.021863f
C31 bgr_0.V_CUR_REF_REG VDDA 3.97245f
C32 V_OSC VCO_FD_magic_0.vco2_3_0.V5 0.017652f
C33 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.139506f
C34 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V5 0.010316f
C35 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.03582f
C36 pfd_8_0.QB_b VDDA 0.512644f
C37 bgr_0.1st_Vout_1 VDDA 2.07565f
C38 VDDA VCO_FD_magic_0.vco2_3_0.V5 0.040599f
C39 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.174311f
C40 bgr_0.V_CUR_REF_REG bgr_0.Vin+ 1.39412f
C41 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.Vin+ 1.06306f
C42 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.122602f
C43 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.M 0.117842f
C44 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V3 0.010316f
C45 pfd_8_0.QA VDDA 0.555755f
C46 F_VCO VCO_FD_magic_0.div120_2_0.div24 0.067402f
C47 VDDA VCO_FD_magic_0.div120_2_0.div2_4_1.C 0.111409f
C48 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.C 0.122602f
C49 bgr_0.Vin+ bgr_0.1st_Vout_1 0.298162f
C50 bgr_0.V_CUR_REF_REG bgr_0.V2 0.953674f
C51 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C52 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.18507f
C53 opamp_cell_4_0.p_bias VDDA 2.92833f
C54 bgr_0.Vin- VDDA 2.07276f
C55 bgr_0.V_CUR_REF_REG F_REF 0.050429f
C56 VDDA V_OSC 0.627267f
C57 bgr_0.Vin- bgr_0.Vin+ 4.62486f
C58 bgr_0.V_TOP bgr_0.V_CUR_REF_REG 0.04372f
C59 VCO_FD_magic_0.vco2_3_0.V4 VDDA 0.413959f
C60 pfd_8_0.QB F_VCO 0.060505f
C61 opamp_cell_4_0.VIN+ VDDA 0.834169f
C62 pfd_8_0.QA F_REF 0.060235f
C63 bgr_0.V_TOP bgr_0.1st_Vout_1 3.49786f
C64 bgr_0.Vin- bgr_0.V2 0.013034f
C65 pfd_8_0.QA_b VDDA 0.529765f
C66 V_OSC VCO_FD_magic_0.vco2_3_0.V7 0.108092f
C67 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.G 0.25905f
C68 bgr_0.Vin+ VDDA 1.85713f
C69 F_VCO pfd_8_0.QB_b 0.043478f
C70 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.D 0.144695f
C71 V_OSC VCO_FD_magic_0.vco2_3_0.V3 0.046941f
C72 VDDA VCO_FD_magic_0.vco2_3_0.V7 0.033517f
C73 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.C 0.122602f
C74 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.C 0.125686f
C75 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.533412f
C76 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.D 0.311052f
C77 pfd_8_0.QB pfd_8_0.QB_b 0.388258f
C78 bgr_0.V2 VDDA 8.46559f
C79 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.104998f
C80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.V_CUR_REF_REG 0.802977f
C81 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.G 0.069172f
C82 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.H 0.106696f
C83 VDDA VCO_FD_magic_0.vco2_3_0.V3 0.040599f
C84 bgr_0.V_TOP bgr_0.Vin- 2.07707f
C85 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.482256f
C86 pfd_8_0.QA pfd_8_0.QB 0.074487f
C87 VDDA VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.111144f
C88 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.112235f
C89 VDDA VCO_FD_magic_0.div120_2_0.div2_4_0.C 0.111144f
C90 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.M 0.157966f
C91 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.061186f
C92 VDDA VCO_FD_magic_0.div120_2_0.div24 0.65395f
C93 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.021344f
C94 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.D 0.070599f
C95 VDDA F_REF 0.123677f
C96 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.016448f
C97 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.C 0.060684f
C98 V_OSC GNDA 2.90637f
C99 F_REF GNDA 1.1128f
C100 VDDA GNDA 0.110713p
C101 VCO_FD_magic_0.vco2_3_0.V2 GNDA 0.045471f
C102 VCO_FD_magic_0.vco2_3_0.V4 GNDA 0.045471f
C103 VCO_FD_magic_0.vco2_3_0.V6 GNDA 0.157087f
C104 VCO_FD_magic_0.div120_2_0.div2_4_1.A GNDA 0.200071f
C105 VCO_FD_magic_0.div120_2_0.div2_4_2.A GNDA 0.200074f
C106 VCO_FD_magic_0.div120_2_0.div2_4_0.A GNDA 0.200071f
C107 VCO_FD_magic_0.div120_2_0.div5_2_0.G GNDA 0.195151f
C108 VCO_FD_magic_0.div120_2_0.div5_2_0.I GNDA 0.152847f
C109 VCO_FD_magic_0.div120_2_0.div3_3_0.C GNDA 0.361544f
C110 VCO_FD_magic_0.div120_2_0.div3_3_0.D GNDA 0.302098f
C111 VCO_FD_magic_0.div120_2_0.div3_3_0.H GNDA 0.42371f
C112 VCO_FD_magic_0.div120_2_0.div5_2_0.D GNDA 0.366931f
C113 VCO_FD_magic_0.div120_2_0.div5_2_0.E GNDA 0.297113f
C114 VCO_FD_magic_0.div120_2_0.div5_2_0.J GNDA 0.398143f
C115 VCO_FD_magic_0.div120_2_0.div5_2_0.K GNDA 0.180033f
C116 VCO_FD_magic_0.div120_2_0.div5_2_0.M GNDA 0.397028f
C117 VCO_FD_magic_0.div120_2_0.div2_4_1.C GNDA 0.457612f
C118 VCO_FD_magic_0.div120_2_0.div2_4_2.C GNDA 0.45762f
C119 VCO_FD_magic_0.div120_2_0.div2_4_0.C GNDA 0.461519f
C120 VCO_FD_magic_0.div120_2_0.div24 GNDA 3.78549f
C121 VCO_FD_magic_0.vco2_3_0.V3 GNDA 0.300759f
C122 VCO_FD_magic_0.vco2_3_0.V5 GNDA 0.302737f
C123 VCO_FD_magic_0.vco2_3_0.V7 GNDA 0.314921f
C124 pfd_8_0.DOWN_input GNDA 2.83935f
C125 pfd_8_0.QB_b GNDA 1.04836f
C126 F_VCO GNDA 3.20723f
C127 pfd_8_0.QB GNDA 1.293329f
C128 pfd_8_0.QA GNDA 3.08755f
C129 pfd_8_0.QA_b GNDA 1.03024f
C130 opamp_cell_4_0.VIN+ GNDA 2.53252f
C131 bgr_0.1st_Vout_1 GNDA 9.9405f
C132 opamp_cell_4_0.p_bias GNDA 3.957291f
C133 bgr_0.V_TOP GNDA 8.259795f
C134 bgr_0.V_CUR_REF_REG GNDA 5.420881f
C135 bgr_0.Vin- GNDA 5.523823f
C136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 16.8112f
C137 bgr_0.Vin+ GNDA 4.971383f
C138 bgr_0.V2 GNDA 8.204531f
C139 loop_filter_2_0.R1_C1.t0 GNDA 2.39887f
C140 a_n1130_7570.t7 GNDA 0.016248f
C141 a_n1130_7570.t6 GNDA 0.016248f
C142 a_n1130_7570.n0 GNDA 0.053414f
C143 a_n1130_7570.t0 GNDA 1.72364f
C144 a_n1130_7570.t1 GNDA 0.04531f
C145 a_n1130_7570.n1 GNDA 1.47476f
C146 a_n1130_7570.t4 GNDA 0.04324f
C147 a_n1130_7570.t2 GNDA 0.04324f
C148 a_n1130_7570.n2 GNDA 0.106515f
C149 a_n1130_7570.n3 GNDA 2.1672f
C150 a_n1130_7570.n4 GNDA 1.2172f
C151 a_n1130_7570.t3 GNDA 0.04324f
C152 a_n1130_7570.n5 GNDA 0.106515f
C153 a_n1130_7570.t5 GNDA 0.04324f
C154 bgr_0.V_CUR_REF_REG.t15 GNDA 0.033253f
C155 bgr_0.V_CUR_REF_REG.t14 GNDA 0.033188f
C156 bgr_0.V_CUR_REF_REG.n0 GNDA 0.233433f
C157 bgr_0.V_CUR_REF_REG.t17 GNDA 0.033188f
C158 bgr_0.V_CUR_REF_REG.n1 GNDA 0.145136f
C159 bgr_0.V_CUR_REF_REG.t13 GNDA 0.033188f
C160 bgr_0.V_CUR_REF_REG.n2 GNDA 0.145136f
C161 bgr_0.V_CUR_REF_REG.t16 GNDA 0.033188f
C162 bgr_0.V_CUR_REF_REG.n3 GNDA 0.300128f
C163 bgr_0.V_CUR_REF_REG.t12 GNDA 0.681769f
C164 bgr_0.V_CUR_REF_REG.t10 GNDA 0.021628f
C165 bgr_0.V_CUR_REF_REG.t8 GNDA 0.021628f
C166 bgr_0.V_CUR_REF_REG.n4 GNDA 0.047663f
C167 bgr_0.V_CUR_REF_REG.t3 GNDA 0.021628f
C168 bgr_0.V_CUR_REF_REG.t6 GNDA 0.021628f
C169 bgr_0.V_CUR_REF_REG.n5 GNDA 0.047367f
C170 bgr_0.V_CUR_REF_REG.n6 GNDA 0.55165f
C171 bgr_0.V_CUR_REF_REG.t9 GNDA 0.021628f
C172 bgr_0.V_CUR_REF_REG.t7 GNDA 0.021628f
C173 bgr_0.V_CUR_REF_REG.n7 GNDA 0.047367f
C174 bgr_0.V_CUR_REF_REG.n8 GNDA 0.291113f
C175 bgr_0.V_CUR_REF_REG.t2 GNDA 0.021628f
C176 bgr_0.V_CUR_REF_REG.t4 GNDA 0.021628f
C177 bgr_0.V_CUR_REF_REG.n9 GNDA 0.047367f
C178 bgr_0.V_CUR_REF_REG.n10 GNDA 0.291113f
C179 bgr_0.V_CUR_REF_REG.t0 GNDA 0.021628f
C180 bgr_0.V_CUR_REF_REG.t5 GNDA 0.021628f
C181 bgr_0.V_CUR_REF_REG.n11 GNDA 0.047367f
C182 bgr_0.V_CUR_REF_REG.n12 GNDA 0.291113f
C183 bgr_0.V_CUR_REF_REG.t1 GNDA 0.021628f
C184 bgr_0.V_CUR_REF_REG.t11 GNDA 0.021628f
C185 bgr_0.V_CUR_REF_REG.n13 GNDA 0.047367f
C186 bgr_0.V_CUR_REF_REG.n14 GNDA 1.14445f
C187 bgr_0.V_CUR_REF_REG.n15 GNDA 5.27065f
C188 opamp_cell_4_0.p_bias.t8 GNDA 1.66267f
C189 opamp_cell_4_0.p_bias.t1 GNDA 0.019693f
C190 opamp_cell_4_0.p_bias.t5 GNDA 0.019693f
C191 opamp_cell_4_0.p_bias.n0 GNDA 0.054067f
C192 opamp_cell_4_0.p_bias.t7 GNDA 0.019693f
C193 opamp_cell_4_0.p_bias.t3 GNDA 0.019693f
C194 opamp_cell_4_0.p_bias.n1 GNDA 0.054067f
C195 opamp_cell_4_0.p_bias.n2 GNDA 0.068502f
C196 opamp_cell_4_0.p_bias.t0 GNDA 0.054353f
C197 opamp_cell_4_0.p_bias.t2 GNDA 0.054353f
C198 opamp_cell_4_0.p_bias.t6 GNDA 0.054353f
C199 opamp_cell_4_0.p_bias.t11 GNDA 0.054353f
C200 opamp_cell_4_0.p_bias.t9 GNDA 0.074733f
C201 opamp_cell_4_0.p_bias.n3 GNDA 0.04185f
C202 opamp_cell_4_0.p_bias.n4 GNDA 0.029697f
C203 opamp_cell_4_0.p_bias.n5 GNDA 0.012761f
C204 opamp_cell_4_0.p_bias.n6 GNDA 0.029697f
C205 opamp_cell_4_0.p_bias.n7 GNDA 0.029697f
C206 opamp_cell_4_0.p_bias.t4 GNDA 0.054353f
C207 opamp_cell_4_0.p_bias.t12 GNDA 0.054353f
C208 opamp_cell_4_0.p_bias.t10 GNDA 0.074733f
C209 opamp_cell_4_0.p_bias.n8 GNDA 0.04185f
C210 opamp_cell_4_0.p_bias.n9 GNDA 0.029697f
C211 opamp_cell_4_0.p_bias.n10 GNDA 0.012761f
C212 opamp_cell_4_0.p_bias.n11 GNDA 0.120625f
C213 bgr_0.Vin-.n0 GNDA 0.771457f
C214 bgr_0.Vin-.n1 GNDA 0.586324f
C215 bgr_0.Vin-.n2 GNDA 0.195749f
C216 bgr_0.Vin-.t3 GNDA 0.428234f
C217 bgr_0.Vin-.n3 GNDA 0.114371f
C218 bgr_0.Vin-.n4 GNDA 0.517468f
C219 bgr_0.Vin-.n5 GNDA 0.11416f
C220 bgr_0.Vin-.n6 GNDA 0.115443f
C221 bgr_0.Vin-.n7 GNDA 0.947747f
C222 bgr_0.Vin-.n8 GNDA 1.96817f
C223 bgr_0.Vin-.t1 GNDA 0.187264f
C224 bgr_0.Vin-.n9 GNDA 0.962593f
C225 bgr_0.Vin-.t6 GNDA 0.044358f
C226 bgr_0.Vin-.t7 GNDA 0.044358f
C227 bgr_0.Vin-.n10 GNDA 0.11867f
C228 bgr_0.Vin-.t4 GNDA 0.044358f
C229 bgr_0.Vin-.t5 GNDA 0.044358f
C230 bgr_0.Vin-.n11 GNDA 0.107634f
C231 bgr_0.Vin-.n12 GNDA 1.21683f
C232 bgr_0.Vin-.t0 GNDA 0.014786f
C233 bgr_0.Vin-.t2 GNDA 0.014786f
C234 bgr_0.Vin-.n13 GNDA 0.041682f
C235 bgr_0.Vin-.n14 GNDA 0.860437f
C236 bgr_0.Vin-.n15 GNDA 0.487885f
C237 bgr_0.Vin-.t10 GNDA 0.024477f
C238 bgr_0.Vin-.t8 GNDA 0.023979f
C239 bgr_0.Vin-.n16 GNDA 0.186829f
C240 bgr_0.Vin-.t9 GNDA 0.023979f
C241 bgr_0.Vin-.n17 GNDA 0.099745f
C242 bgr_0.Vin-.t11 GNDA 0.024302f
C243 bgr_0.Vin-.n18 GNDA 0.100457f
C244 bgr_0.Vin-.t12 GNDA 0.024302f
C245 bgr_0.Vin-.n19 GNDA 0.201113f
C246 bgr_0.V_mir1.t10 GNDA 0.018056f
C247 bgr_0.V_mir1.t5 GNDA 0.027505f
C248 bgr_0.V_mir1.t11 GNDA 0.021667f
C249 bgr_0.V_mir1.t21 GNDA 0.021667f
C250 bgr_0.V_mir1.t18 GNDA 0.034973f
C251 bgr_0.V_mir1.n0 GNDA 0.039055f
C252 bgr_0.V_mir1.n1 GNDA 0.02668f
C253 bgr_0.V_mir1.n2 GNDA 0.043175f
C254 bgr_0.V_mir1.t6 GNDA 0.018056f
C255 bgr_0.V_mir1.t12 GNDA 0.018056f
C256 bgr_0.V_mir1.n3 GNDA 0.036969f
C257 bgr_0.V_mir1.n4 GNDA 0.191386f
C258 bgr_0.V_mir1.n5 GNDA 0.019256f
C259 bgr_0.V_mir1.t3 GNDA 0.034183f
C260 bgr_0.V_mir1.n6 GNDA 0.021429f
C261 bgr_0.V_mir1.n7 GNDA 0.554666f
C262 bgr_0.V_mir1.n8 GNDA 0.186578f
C263 bgr_0.V_mir1.t7 GNDA 0.027505f
C264 bgr_0.V_mir1.t13 GNDA 0.021667f
C265 bgr_0.V_mir1.t20 GNDA 0.021667f
C266 bgr_0.V_mir1.t17 GNDA 0.034973f
C267 bgr_0.V_mir1.n9 GNDA 0.039055f
C268 bgr_0.V_mir1.n10 GNDA 0.02668f
C269 bgr_0.V_mir1.n11 GNDA 0.043175f
C270 bgr_0.V_mir1.t8 GNDA 0.018056f
C271 bgr_0.V_mir1.t14 GNDA 0.018056f
C272 bgr_0.V_mir1.n12 GNDA 0.036969f
C273 bgr_0.V_mir1.n13 GNDA 0.239421f
C274 bgr_0.V_mir1.n14 GNDA 0.26218f
C275 bgr_0.V_mir1.t9 GNDA 0.027505f
C276 bgr_0.V_mir1.t15 GNDA 0.021667f
C277 bgr_0.V_mir1.t19 GNDA 0.021667f
C278 bgr_0.V_mir1.t22 GNDA 0.034973f
C279 bgr_0.V_mir1.n15 GNDA 0.039055f
C280 bgr_0.V_mir1.n16 GNDA 0.02668f
C281 bgr_0.V_mir1.n17 GNDA 0.043175f
C282 bgr_0.V_mir1.n18 GNDA 0.191386f
C283 bgr_0.V_mir1.n19 GNDA 0.036969f
C284 bgr_0.V_mir1.t16 GNDA 0.018056f
C285 pfd_8_0.opamp_out.t12 GNDA 1.08371f
C286 pfd_8_0.opamp_out.n2 GNDA 0.010903f
C287 pfd_8_0.opamp_out.t11 GNDA 1.08325f
C288 pfd_8_0.opamp_out.n6 GNDA 0.014659f
C289 pfd_8_0.opamp_out.t14 GNDA 0.014564f
C290 pfd_8_0.opamp_out.t13 GNDA 0.010463f
C291 pfd_8_0.opamp_out.t6 GNDA 0.013605f
C292 pfd_8_0.opamp_out.n13 GNDA 0.018307f
C293 pfd_8_0.opamp_out.n14 GNDA 0.103761f
C294 pfd_8_0.opamp_out.n15 GNDA 0.052015f
C295 VCO_FD_magic_0.vco2_3_0.V1.t1 GNDA 0.104706f
C296 VCO_FD_magic_0.vco2_3_0.V1.n0 GNDA 0.184398f
C297 VCO_FD_magic_0.vco2_3_0.V1.t4 GNDA 0.298444f
C298 VCO_FD_magic_0.vco2_3_0.V1.t3 GNDA 0.298444f
C299 VCO_FD_magic_0.vco2_3_0.V1.t5 GNDA 0.497217f
C300 VCO_FD_magic_0.vco2_3_0.V1.n1 GNDA 0.243367f
C301 VCO_FD_magic_0.vco2_3_0.V1.n2 GNDA 0.217957f
C302 VCO_FD_magic_0.vco2_3_0.V1.t0 GNDA 0.298444f
C303 VCO_FD_magic_0.vco2_3_0.V1.n3 GNDA 0.169192f
C304 VCO_FD_magic_0.vco2_3_0.V1.n4 GNDA 0.045341f
C305 VCO_FD_magic_0.vco2_3_0.V1.n5 GNDA 0.177452f
C306 VCO_FD_magic_0.vco2_3_0.V1.t2 GNDA 0.165036f
C307 pfd_8_0.UP_b.t0 GNDA 1.81459f
C308 pfd_8_0.UP_b.t3 GNDA 0.010202f
C309 pfd_8_0.UP_b.t1 GNDA 0.026993f
C310 pfd_8_0.UP_b.t2 GNDA 0.050413f
C311 pfd_8_0.UP_b.n0 GNDA 0.069085f
C312 pfd_8_0.UP_b.n1 GNDA 0.020893f
C313 charge_pump_cell_6_0.UP_b GNDA 0.207826f
C314 bgr_0.cap_res1.t14 GNDA 0.31433f
C315 bgr_0.cap_res1.t7 GNDA 0.331199f
C316 bgr_0.cap_res1.t2 GNDA 0.331199f
C317 bgr_0.cap_res1.t16 GNDA 0.331199f
C318 bgr_0.cap_res1.t9 GNDA 0.331199f
C319 bgr_0.cap_res1.t5 GNDA 0.331199f
C320 bgr_0.cap_res1.t20 GNDA 0.331199f
C321 bgr_0.cap_res1.t10 GNDA 0.331199f
C322 bgr_0.cap_res1.t3 GNDA 0.315469f
C323 bgr_0.cap_res1.t18 GNDA 0.151964f
C324 bgr_0.cap_res1.n0 GNDA 0.19601f
C325 bgr_0.cap_res1.t12 GNDA 0.344559f
C326 bgr_0.cap_res1.t17 GNDA 0.316794f
C327 bgr_0.cap_res1.t6 GNDA 0.331199f
C328 bgr_0.cap_res1.t13 GNDA 0.331199f
C329 bgr_0.cap_res1.t19 GNDA 0.331199f
C330 bgr_0.cap_res1.t4 GNDA 0.331199f
C331 bgr_0.cap_res1.t11 GNDA 0.331199f
C332 bgr_0.cap_res1.t15 GNDA 0.331199f
C333 bgr_0.cap_res1.t1 GNDA 0.331199f
C334 bgr_0.cap_res1.t8 GNDA 0.722653f
C335 bgr_0.cap_res1.t0 GNDA 0.101437f
C336 a_n1450_5080.t8 GNDA 0.02f
C337 a_n1450_5080.t18 GNDA 0.02f
C338 a_n1450_5080.t20 GNDA 0.032283f
C339 a_n1450_5080.n0 GNDA 0.036051f
C340 a_n1450_5080.n1 GNDA 0.024627f
C341 a_n1450_5080.t6 GNDA 0.025389f
C342 a_n1450_5080.n2 GNDA 0.039854f
C343 a_n1450_5080.t9 GNDA 0.016667f
C344 a_n1450_5080.t7 GNDA 0.016667f
C345 a_n1450_5080.n3 GNDA 0.034125f
C346 a_n1450_5080.n4 GNDA 0.176664f
C347 a_n1450_5080.n5 GNDA 0.017774f
C348 a_n1450_5080.t13 GNDA 0.031554f
C349 a_n1450_5080.n6 GNDA 0.019781f
C350 a_n1450_5080.n7 GNDA 0.511999f
C351 a_n1450_5080.n8 GNDA 0.172226f
C352 a_n1450_5080.t4 GNDA 0.02f
C353 a_n1450_5080.t22 GNDA 0.02f
C354 a_n1450_5080.t21 GNDA 0.032283f
C355 a_n1450_5080.n9 GNDA 0.036051f
C356 a_n1450_5080.n10 GNDA 0.024627f
C357 a_n1450_5080.t0 GNDA 0.025389f
C358 a_n1450_5080.n11 GNDA 0.039854f
C359 a_n1450_5080.t5 GNDA 0.016667f
C360 a_n1450_5080.t1 GNDA 0.016667f
C361 a_n1450_5080.n12 GNDA 0.034125f
C362 a_n1450_5080.n13 GNDA 0.221004f
C363 a_n1450_5080.n14 GNDA 0.242013f
C364 a_n1450_5080.t10 GNDA 0.02f
C365 a_n1450_5080.t17 GNDA 0.02f
C366 a_n1450_5080.t19 GNDA 0.032283f
C367 a_n1450_5080.n15 GNDA 0.036051f
C368 a_n1450_5080.n16 GNDA 0.024627f
C369 a_n1450_5080.t2 GNDA 0.025389f
C370 a_n1450_5080.n17 GNDA 0.039854f
C371 a_n1450_5080.n18 GNDA 0.176664f
C372 a_n1450_5080.t3 GNDA 0.016667f
C373 a_n1450_5080.n19 GNDA 0.034125f
C374 a_n1450_5080.t11 GNDA 0.016667f
C375 bgr_0.V1.t1 GNDA 0.10095f
C376 bgr_0.V1.t6 GNDA 0.10095f
C377 bgr_0.V1.n0 GNDA 0.281599f
C378 bgr_0.V1.t3 GNDA 0.10095f
C379 bgr_0.V1.t5 GNDA 0.10095f
C380 bgr_0.V1.n1 GNDA 0.253459f
C381 bgr_0.V1.n2 GNDA 3.1126f
C382 bgr_0.V1.t4 GNDA 0.10095f
C383 bgr_0.V1.t2 GNDA 0.10095f
C384 bgr_0.V1.n3 GNDA 0.253459f
C385 bgr_0.V1.n4 GNDA 2.34993f
C386 bgr_0.V1.t9 GNDA 0.055705f
C387 bgr_0.V1.t10 GNDA 0.05457f
C388 bgr_0.V1.n5 GNDA 0.425181f
C389 bgr_0.V1.t11 GNDA 0.05457f
C390 bgr_0.V1.n6 GNDA 0.226997f
C391 bgr_0.V1.t7 GNDA 0.055305f
C392 bgr_0.V1.n7 GNDA 0.228617f
C393 bgr_0.V1.t8 GNDA 0.055305f
C394 bgr_0.V1.n8 GNDA 0.780841f
C395 bgr_0.V1.n9 GNDA 4.03498f
C396 bgr_0.V1.t0 GNDA 0.471183f
C397 BGR_CURRENT_OUT.n0 GNDA 2.0431f
C398 BGR_CURRENT_OUT.n1 GNDA 0.097815f
C399 BGR_CURRENT_OUT.n2 GNDA 0.117429f
C400 bgr_0.CURRENT_OUTPUT GNDA 0.059985f
C401 BGR_CURRENT_OUT.t4 GNDA 0.010639f
C402 BGR_CURRENT_OUT.t2 GNDA 0.010639f
C403 BGR_CURRENT_OUT.n3 GNDA 0.041426f
C404 BGR_CURRENT_OUT.t1 GNDA 0.049455f
C405 BGR_CURRENT_OUT.t19 GNDA 0.04628f
C406 BGR_CURRENT_OUT.t18 GNDA 0.062085f
C407 BGR_CURRENT_OUT.n4 GNDA 0.046455f
C408 BGR_CURRENT_OUT.n5 GNDA 0.048543f
C409 BGR_CURRENT_OUT.t3 GNDA 0.03365f
C410 BGR_CURRENT_OUT.n6 GNDA 0.040235f
C411 BGR_CURRENT_OUT.n7 GNDA 0.034459f
C412 BGR_CURRENT_OUT.t0 GNDA 0.037686f
C413 BGR_CURRENT_OUT.t17 GNDA 0.030908f
C414 BGR_CURRENT_OUT.n8 GNDA 0.060622f
C415 BGR_CURRENT_OUT.n10 GNDA 0.018725f
C416 BGR_CURRENT_OUT.n13 GNDA 0.062631f
C417 BGR_CURRENT_OUT.n15 GNDA 0.030586f
C418 BGR_CURRENT_OUT.n16 GNDA 0.059176f
C419 BGR_CURRENT_OUT.n18 GNDA 0.059176f
C420 BGR_CURRENT_OUT.n19 GNDA 0.018725f
C421 BGR_CURRENT_OUT.n21 GNDA 0.059176f
C422 BGR_CURRENT_OUT.n22 GNDA 0.030586f
C423 BGR_CURRENT_OUT.n23 GNDA 0.060082f
C424 BGR_CURRENT_OUT.n24 GNDA 1.61553f
C425 bgr_0.V2.t0 GNDA 0.422109f
C426 bgr_0.V2.t28 GNDA 0.049701f
C427 bgr_0.V2.t19 GNDA 0.049641f
C428 bgr_0.V2.n0 GNDA 0.259633f
C429 bgr_0.V2.t11 GNDA 0.049641f
C430 bgr_0.V2.n1 GNDA 0.136128f
C431 bgr_0.V2.t25 GNDA 0.049641f
C432 bgr_0.V2.n2 GNDA 0.136128f
C433 bgr_0.V2.t10 GNDA 0.049641f
C434 bgr_0.V2.n3 GNDA 0.136128f
C435 bgr_0.V2.t21 GNDA 0.049641f
C436 bgr_0.V2.n4 GNDA 0.136128f
C437 bgr_0.V2.t12 GNDA 0.049641f
C438 bgr_0.V2.n5 GNDA 0.136128f
C439 bgr_0.V2.t22 GNDA 0.049641f
C440 bgr_0.V2.n6 GNDA 0.136128f
C441 bgr_0.V2.t14 GNDA 0.049641f
C442 bgr_0.V2.n7 GNDA 0.136128f
C443 bgr_0.V2.t23 GNDA 0.049641f
C444 bgr_0.V2.n8 GNDA 0.337114f
C445 bgr_0.V2.t15 GNDA 0.049641f
C446 bgr_0.V2.n9 GNDA 0.337114f
C447 bgr_0.V2.t24 GNDA 0.049641f
C448 bgr_0.V2.n10 GNDA 0.136128f
C449 bgr_0.V2.t17 GNDA 0.049641f
C450 bgr_0.V2.n11 GNDA 0.136128f
C451 bgr_0.V2.t13 GNDA 0.049641f
C452 bgr_0.V2.n12 GNDA 0.136128f
C453 bgr_0.V2.t16 GNDA 0.049641f
C454 bgr_0.V2.n13 GNDA 0.136128f
C455 bgr_0.V2.t26 GNDA 0.049641f
C456 bgr_0.V2.n14 GNDA 0.136128f
C457 bgr_0.V2.t20 GNDA 0.049641f
C458 bgr_0.V2.n15 GNDA 0.136128f
C459 bgr_0.V2.t29 GNDA 0.049641f
C460 bgr_0.V2.n16 GNDA 0.136128f
C461 bgr_0.V2.t18 GNDA 0.049641f
C462 bgr_0.V2.n17 GNDA 0.136128f
C463 bgr_0.V2.t27 GNDA 0.049641f
C464 bgr_0.V2.n18 GNDA 0.992373f
C465 bgr_0.V2.t7 GNDA 0.43431f
C466 bgr_0.V2.t8 GNDA 0.028712f
C467 bgr_0.V2.t2 GNDA 0.028712f
C468 bgr_0.V2.n19 GNDA 0.062021f
C469 bgr_0.V2.n20 GNDA 1.41734f
C470 bgr_0.V2.t4 GNDA 0.028712f
C471 bgr_0.V2.t3 GNDA 0.028712f
C472 bgr_0.V2.n21 GNDA 0.062021f
C473 bgr_0.V2.n22 GNDA 0.627074f
C474 bgr_0.V2.t6 GNDA 0.028712f
C475 bgr_0.V2.t5 GNDA 0.028712f
C476 bgr_0.V2.n23 GNDA 0.062021f
C477 bgr_0.V2.n24 GNDA 0.614154f
C478 bgr_0.V2.t1 GNDA 0.028712f
C479 bgr_0.V2.t9 GNDA 0.028712f
C480 bgr_0.V2.n25 GNDA 0.062021f
C481 bgr_0.V2.n26 GNDA 0.715576f
C482 bgr_0.V2.n27 GNDA 1.19812f
C483 bgr_0.Vin+.t0 GNDA 0.342532f
C484 bgr_0.Vin+.t1 GNDA 0.148895f
C485 bgr_0.Vin+.n0 GNDA 2.17873f
C486 bgr_0.Vin+.t2 GNDA 0.051177f
C487 bgr_0.Vin+.t3 GNDA 0.051177f
C488 bgr_0.Vin+.n1 GNDA 0.127304f
C489 bgr_0.Vin+.t4 GNDA 0.051177f
C490 bgr_0.Vin+.t5 GNDA 0.051177f
C491 bgr_0.Vin+.n2 GNDA 0.122338f
C492 bgr_0.Vin+.n3 GNDA 1.74488f
C493 bgr_0.Vin+.n4 GNDA 0.850702f
C494 bgr_0.Vin+.t8 GNDA 0.026228f
C495 bgr_0.Vin+.t9 GNDA 0.026176f
C496 bgr_0.Vin+.n5 GNDA 0.184117f
C497 bgr_0.Vin+.t6 GNDA 0.026176f
C498 bgr_0.Vin+.n6 GNDA 0.114474f
C499 bgr_0.Vin+.t7 GNDA 0.026176f
C500 bgr_0.Vin+.n7 GNDA 0.114474f
C501 bgr_0.Vin+.t10 GNDA 0.026176f
C502 bgr_0.Vin+.n8 GNDA 0.244185f
C503 bgr_0.cap_res2.t10 GNDA 0.293845f
C504 bgr_0.cap_res2.t12 GNDA 0.309615f
C505 bgr_0.cap_res2.t6 GNDA 0.309615f
C506 bgr_0.cap_res2.t20 GNDA 0.309615f
C507 bgr_0.cap_res2.t3 GNDA 0.309615f
C508 bgr_0.cap_res2.t18 GNDA 0.309615f
C509 bgr_0.cap_res2.t14 GNDA 0.309615f
C510 bgr_0.cap_res2.t11 GNDA 0.309615f
C511 bgr_0.cap_res2.t15 GNDA 0.29491f
C512 bgr_0.cap_res2.t9 GNDA 0.14206f
C513 bgr_0.cap_res2.n0 GNDA 0.183237f
C514 bgr_0.cap_res2.t1 GNDA 0.322105f
C515 bgr_0.cap_res2.t8 GNDA 0.296149f
C516 bgr_0.cap_res2.t4 GNDA 0.309615f
C517 bgr_0.cap_res2.t7 GNDA 0.309615f
C518 bgr_0.cap_res2.t13 GNDA 0.309615f
C519 bgr_0.cap_res2.t17 GNDA 0.309615f
C520 bgr_0.cap_res2.t16 GNDA 0.309615f
C521 bgr_0.cap_res2.t19 GNDA 0.309615f
C522 bgr_0.cap_res2.t5 GNDA 0.309615f
C523 bgr_0.cap_res2.t2 GNDA 1.13635f
C524 bgr_0.cap_res2.t0 GNDA 0.196735f
C525 bgr_0.1st_Vout_2.n0 GNDA 1.17563f
C526 bgr_0.1st_Vout_2.n1 GNDA 0.901667f
C527 bgr_0.1st_Vout_2.n2 GNDA 2.31979f
C528 bgr_0.1st_Vout_2.n3 GNDA 0.533984f
C529 bgr_0.1st_Vout_2.n4 GNDA 0.176376f
C530 bgr_0.1st_Vout_2.n5 GNDA 0.289395f
C531 bgr_0.1st_Vout_2.t2 GNDA 0.010305f
C532 bgr_0.1st_Vout_2.t25 GNDA 0.024727f
C533 bgr_0.1st_Vout_2.t8 GNDA 0.010305f
C534 bgr_0.1st_Vout_2.t9 GNDA 0.010305f
C535 bgr_0.1st_Vout_2.n6 GNDA 0.022597f
C536 bgr_0.1st_Vout_2.t20 GNDA 0.015954f
C537 bgr_0.1st_Vout_2.t24 GNDA 0.015954f
C538 bgr_0.1st_Vout_2.n7 GNDA 0.030906f
C539 bgr_0.1st_Vout_2.t10 GNDA 0.010305f
C540 bgr_0.1st_Vout_2.t4 GNDA 0.010305f
C541 bgr_0.1st_Vout_2.n8 GNDA 0.022597f
C542 bgr_0.1st_Vout_2.t6 GNDA 0.018148f
C543 bgr_0.1st_Vout_2.n9 GNDA 0.013021f
C544 bgr_0.1st_Vout_2.n10 GNDA 0.012563f
C545 bgr_0.1st_Vout_2.n11 GNDA 0.335083f
C546 bgr_0.1st_Vout_2.t13 GNDA 0.015954f
C547 bgr_0.1st_Vout_2.t16 GNDA 0.015954f
C548 bgr_0.1st_Vout_2.n12 GNDA 0.029642f
C549 bgr_0.1st_Vout_2.t34 GNDA 0.024402f
C550 bgr_0.1st_Vout_2.t36 GNDA 0.41219f
C551 bgr_0.1st_Vout_2.t35 GNDA 0.419031f
C552 bgr_0.1st_Vout_2.t31 GNDA 0.41219f
C553 bgr_0.1st_Vout_2.t12 GNDA 0.41219f
C554 bgr_0.1st_Vout_2.t17 GNDA 0.41219f
C555 bgr_0.1st_Vout_2.t15 GNDA 0.41219f
C556 bgr_0.1st_Vout_2.t21 GNDA 0.41219f
C557 bgr_0.1st_Vout_2.t29 GNDA 0.41219f
C558 bgr_0.1st_Vout_2.t32 GNDA 0.41219f
C559 bgr_0.1st_Vout_2.t28 GNDA 0.41219f
C560 bgr_0.1st_Vout_2.t27 GNDA 0.41219f
C561 bgr_0.1st_Vout_2.t18 GNDA 0.41219f
C562 bgr_0.1st_Vout_2.t23 GNDA 0.41219f
C563 bgr_0.1st_Vout_2.t19 GNDA 0.41219f
C564 bgr_0.1st_Vout_2.t14 GNDA 0.41219f
C565 bgr_0.1st_Vout_2.t33 GNDA 0.41219f
C566 bgr_0.1st_Vout_2.t11 GNDA 0.41219f
C567 bgr_0.1st_Vout_2.t30 GNDA 0.41219f
C568 bgr_0.1st_Vout_2.t22 GNDA 0.41219f
C569 bgr_0.1st_Vout_2.t26 GNDA 0.41219f
C570 bgr_0.1st_Vout_2.n13 GNDA 0.949966f
C571 bgr_0.1st_Vout_2.n14 GNDA 0.022597f
C572 bgr_0.1st_Vout_2.t1 GNDA 0.010305f
C573 pfd_8_0.QB.t5 GNDA 0.069179f
C574 pfd_8_0.QB.t6 GNDA 0.032493f
C575 pfd_8_0.QB.n0 GNDA 0.099932f
C576 pfd_8_0.QB.t7 GNDA 0.069179f
C577 pfd_8_0.QB.t8 GNDA 0.104293f
C578 pfd_8_0.QB.n1 GNDA 1.25065f
C579 pfd_8_0.QB.t3 GNDA 0.069862f
C580 pfd_8_0.QB.t4 GNDA 0.030633f
C581 pfd_8_0.QB.n2 GNDA 0.176466f
C582 pfd_8_0.QB.t2 GNDA 0.147114f
C583 pfd_8_0.QB.t0 GNDA 0.027951f
C584 pfd_8_0.QB.t1 GNDA 0.027951f
C585 pfd_8_0.QB.n3 GNDA 0.149246f
C586 pfd_8_0.QB.n4 GNDA 0.265156f
C587 pfd_8_0.QB.n5 GNDA 0.226459f
C588 bgr_0.V_TOP.n0 GNDA 0.022936f
C589 bgr_0.V_TOP.t14 GNDA 0.1754f
C590 bgr_0.V_TOP.t33 GNDA 0.175758f
C591 bgr_0.V_TOP.t19 GNDA 0.176515f
C592 bgr_0.V_TOP.n1 GNDA 0.222088f
C593 bgr_0.V_TOP.t41 GNDA 0.176515f
C594 bgr_0.V_TOP.n2 GNDA 0.121656f
C595 bgr_0.V_TOP.t37 GNDA 0.176515f
C596 bgr_0.V_TOP.n3 GNDA 0.121656f
C597 bgr_0.V_TOP.t32 GNDA 0.176515f
C598 bgr_0.V_TOP.n4 GNDA 0.121656f
C599 bgr_0.V_TOP.t27 GNDA 0.176515f
C600 bgr_0.V_TOP.n5 GNDA 0.121656f
C601 bgr_0.V_TOP.n6 GNDA 0.034404f
C602 bgr_0.V_TOP.n7 GNDA 0.078172f
C603 bgr_0.V_TOP.t3 GNDA 0.174413f
C604 bgr_0.V_TOP.t1 GNDA 0.143852f
C605 bgr_0.V_TOP.t25 GNDA 0.509694f
C606 bgr_0.V_TOP.t24 GNDA 0.518153f
C607 bgr_0.V_TOP.t20 GNDA 0.509694f
C608 bgr_0.V_TOP.n8 GNDA 0.338771f
C609 bgr_0.V_TOP.t29 GNDA 0.509694f
C610 bgr_0.V_TOP.n9 GNDA 0.222991f
C611 bgr_0.V_TOP.t42 GNDA 0.509694f
C612 bgr_0.V_TOP.n10 GNDA 0.222991f
C613 bgr_0.V_TOP.t34 GNDA 0.509694f
C614 bgr_0.V_TOP.n11 GNDA 0.222991f
C615 bgr_0.V_TOP.t46 GNDA 0.509694f
C616 bgr_0.V_TOP.n12 GNDA 0.222991f
C617 bgr_0.V_TOP.t17 GNDA 0.509694f
C618 bgr_0.V_TOP.n13 GNDA 0.222991f
C619 bgr_0.V_TOP.t22 GNDA 0.509694f
C620 bgr_0.V_TOP.n14 GNDA 0.222991f
C621 bgr_0.V_TOP.t15 GNDA 0.509694f
C622 bgr_0.V_TOP.n15 GNDA 0.222991f
C623 bgr_0.V_TOP.n16 GNDA 0.222991f
C624 bgr_0.V_TOP.t38 GNDA 0.509694f
C625 bgr_0.V_TOP.n17 GNDA 0.222991f
C626 bgr_0.V_TOP.t23 GNDA 0.509694f
C627 bgr_0.V_TOP.n18 GNDA 0.222991f
C628 bgr_0.V_TOP.t31 GNDA 0.509694f
C629 bgr_0.V_TOP.n19 GNDA 0.222991f
C630 bgr_0.V_TOP.t26 GNDA 0.509694f
C631 bgr_0.V_TOP.n20 GNDA 0.222991f
C632 bgr_0.V_TOP.t16 GNDA 0.509694f
C633 bgr_0.V_TOP.n21 GNDA 0.222991f
C634 bgr_0.V_TOP.t45 GNDA 0.509694f
C635 bgr_0.V_TOP.n22 GNDA 0.222991f
C636 bgr_0.V_TOP.t49 GNDA 0.509694f
C637 bgr_0.V_TOP.n23 GNDA 0.222991f
C638 bgr_0.V_TOP.t40 GNDA 0.509694f
C639 bgr_0.V_TOP.n24 GNDA 0.222991f
C640 bgr_0.V_TOP.t28 GNDA 0.509694f
C641 bgr_0.V_TOP.n25 GNDA 0.221398f
C642 bgr_0.V_TOP.t35 GNDA 0.509694f
C643 bgr_0.V_TOP.n26 GNDA 0.391094f
C644 bgr_0.V_TOP.n27 GNDA 1.20222f
C645 bgr_0.V_TOP.t5 GNDA 0.012742f
C646 bgr_0.V_TOP.t10 GNDA 0.012742f
C647 bgr_0.V_TOP.n28 GNDA 0.02609f
C648 bgr_0.V_TOP.t2 GNDA 0.012742f
C649 bgr_0.V_TOP.t7 GNDA 0.012742f
C650 bgr_0.V_TOP.n29 GNDA 0.029654f
C651 bgr_0.V_TOP.t6 GNDA 0.012742f
C652 bgr_0.V_TOP.t0 GNDA 0.012742f
C653 bgr_0.V_TOP.n30 GNDA 0.02609f
C654 bgr_0.V_TOP.n31 GNDA 0.349463f
C655 bgr_0.V_TOP.n32 GNDA 0.216014f
C656 bgr_0.V_TOP.n33 GNDA 0.654381f
C657 bgr_0.V_TOP.t9 GNDA 0.012742f
C658 bgr_0.V_TOP.t8 GNDA 0.012742f
C659 bgr_0.V_TOP.n34 GNDA 0.027525f
C660 bgr_0.V_TOP.n35 GNDA 0.270646f
C661 bgr_0.V_TOP.t11 GNDA 0.012742f
C662 bgr_0.V_TOP.t13 GNDA 0.012742f
C663 bgr_0.V_TOP.n36 GNDA 0.027525f
C664 bgr_0.V_TOP.n37 GNDA 0.278292f
C665 bgr_0.V_TOP.t12 GNDA 0.012742f
C666 bgr_0.V_TOP.t4 GNDA 0.012742f
C667 bgr_0.V_TOP.n38 GNDA 0.027525f
C668 bgr_0.V_TOP.n39 GNDA 0.259414f
C669 bgr_0.V_TOP.n40 GNDA 0.477123f
C670 bgr_0.V_TOP.n41 GNDA 0.122327f
C671 bgr_0.V_TOP.t48 GNDA 0.174142f
C672 bgr_0.V_TOP.n42 GNDA 0.071785f
C673 bgr_0.V_TOP.n43 GNDA 0.034404f
C674 bgr_0.V_TOP.t44 GNDA 0.175158f
C675 bgr_0.V_TOP.n44 GNDA 0.115368f
C676 bgr_0.V_TOP.t39 GNDA 0.176515f
C677 bgr_0.V_TOP.n45 GNDA 0.121656f
C678 bgr_0.V_TOP.t36 GNDA 0.176515f
C679 bgr_0.V_TOP.n46 GNDA 0.121656f
C680 bgr_0.V_TOP.t21 GNDA 0.176515f
C681 bgr_0.V_TOP.n47 GNDA 0.121656f
C682 bgr_0.V_TOP.t18 GNDA 0.176515f
C683 bgr_0.V_TOP.n48 GNDA 0.121656f
C684 bgr_0.V_TOP.t30 GNDA 0.176515f
C685 bgr_0.V_TOP.n49 GNDA 0.121656f
C686 bgr_0.V_TOP.t43 GNDA 0.176515f
C687 bgr_0.V_TOP.n50 GNDA 0.110188f
C688 bgr_0.V_TOP.t47 GNDA 0.175198f
C689 bgr_0.1st_Vout_1.n0 GNDA 1.02458f
C690 bgr_0.1st_Vout_1.n1 GNDA 0.785813f
C691 bgr_0.1st_Vout_1.n2 GNDA 1.6475f
C692 bgr_0.1st_Vout_1.n3 GNDA 0.153679f
C693 bgr_0.1st_Vout_1.t22 GNDA 0.359229f
C694 bgr_0.1st_Vout_1.t27 GNDA 0.36519f
C695 bgr_0.1st_Vout_1.t36 GNDA 0.359229f
C696 bgr_0.1st_Vout_1.t19 GNDA 0.359229f
C697 bgr_0.1st_Vout_1.t23 GNDA 0.359229f
C698 bgr_0.1st_Vout_1.t33 GNDA 0.359229f
C699 bgr_0.1st_Vout_1.t13 GNDA 0.359229f
C700 bgr_0.1st_Vout_1.t21 GNDA 0.359229f
C701 bgr_0.1st_Vout_1.t31 GNDA 0.359229f
C702 bgr_0.1st_Vout_1.t16 GNDA 0.359229f
C703 bgr_0.1st_Vout_1.t14 GNDA 0.359229f
C704 bgr_0.1st_Vout_1.t34 GNDA 0.359229f
C705 bgr_0.1st_Vout_1.t24 GNDA 0.359229f
C706 bgr_0.1st_Vout_1.t12 GNDA 0.359229f
C707 bgr_0.1st_Vout_1.t32 GNDA 0.359229f
C708 bgr_0.1st_Vout_1.t26 GNDA 0.359229f
C709 bgr_0.1st_Vout_1.t18 GNDA 0.359229f
C710 bgr_0.1st_Vout_1.t35 GNDA 0.359229f
C711 bgr_0.1st_Vout_1.t29 GNDA 0.359229f
C712 bgr_0.1st_Vout_1.t20 GNDA 0.359229f
C713 bgr_0.1st_Vout_1.t25 GNDA 0.021589f
C714 bgr_0.1st_Vout_1.n4 GNDA 0.019024f
C715 bgr_0.1st_Vout_1.t2 GNDA 0.015816f
C716 bgr_0.1st_Vout_1.n5 GNDA 0.011348f
C717 bgr_0.1st_Vout_1.n6 GNDA 0.010949f
C718 bgr_0.1st_Vout_1.n7 GNDA 0.292028f
C719 bgr_0.1st_Vout_1.t28 GNDA 0.013904f
C720 bgr_0.1st_Vout_1.t30 GNDA 0.013904f
C721 bgr_0.1st_Vout_1.n8 GNDA 0.025867f
C722 bgr_0.1st_Vout_1.n9 GNDA 0.019024f
C723 bgr_0.1st_Vout_1.t17 GNDA 0.013904f
C724 bgr_0.1st_Vout_1.t11 GNDA 0.013904f
C725 bgr_0.1st_Vout_1.n10 GNDA 0.026482f
C726 bgr_0.1st_Vout_1.n11 GNDA 0.019024f
C727 bgr_0.1st_Vout_1.t15 GNDA 0.021208f
C728 VDDA.n8 GNDA 0.013807f
C729 VDDA.n17 GNDA 0.012084f
C730 VDDA.n29 GNDA 0.013807f
C731 VDDA.n35 GNDA 0.012084f
C732 VDDA.n49 GNDA 0.013807f
C733 VDDA.n53 GNDA 0.012084f
C734 VDDA.n67 GNDA 0.016447f
C735 VDDA.n71 GNDA 0.151836f
C736 VDDA.t342 GNDA 0.508569f
C737 VDDA.n74 GNDA 0.339046f
C738 VDDA.n75 GNDA 0.012482f
C739 VDDA.n78 GNDA 0.012482f
C740 VDDA.n80 GNDA 0.036533f
C741 VDDA.t343 GNDA 0.022648f
C742 VDDA.n82 GNDA 0.023612f
C743 VDDA.n83 GNDA 0.023612f
C744 VDDA.n86 GNDA 0.042321f
C745 VDDA.t261 GNDA 0.015182f
C746 VDDA.n87 GNDA 0.114002f
C747 VDDA.t236 GNDA 0.262871f
C748 VDDA.t74 GNDA 0.207195f
C749 VDDA.t211 GNDA 0.09748f
C750 VDDA.n89 GNDA 0.012084f
C751 VDDA.n90 GNDA 0.043095f
C752 VDDA.t19 GNDA 0.044514f
C753 VDDA.t111 GNDA 0.075505f
C754 VDDA.t144 GNDA 0.075505f
C755 VDDA.t225 GNDA 0.049585f
C756 VDDA.t399 GNDA 0.049585f
C757 VDDA.t72 GNDA 0.024792f
C758 VDDA.t220 GNDA 0.082266f
C759 VDDA.t164 GNDA 0.085084f
C760 VDDA.n91 GNDA 0.043095f
C761 VDDA.t90 GNDA 0.044514f
C762 VDDA.t190 GNDA 0.050712f
C763 VDDA.t47 GNDA 0.050712f
C764 VDDA.t43 GNDA 0.04057f
C765 VDDA.t37 GNDA 0.04057f
C766 VDDA.t77 GNDA 0.065362f
C767 VDDA.t98 GNDA 0.065362f
C768 VDDA.t176 GNDA 0.049585f
C769 VDDA.t340 GNDA 0.049585f
C770 VDDA.t389 GNDA 0.06987f
C771 VDDA.t15 GNDA 0.072687f
C772 VDDA.n92 GNDA 0.03408f
C773 VDDA.t107 GNDA 0.035498f
C774 VDDA.t209 GNDA 0.04057f
C775 VDDA.t201 GNDA 0.04057f
C776 VDDA.t206 GNDA 0.067616f
C777 VDDA.t53 GNDA 0.070433f
C778 VDDA.n93 GNDA 0.012084f
C779 VDDA.n94 GNDA 0.03408f
C780 VDDA.t75 GNDA 0.035498f
C781 VDDA.t116 GNDA 0.04057f
C782 VDDA.t11 GNDA 0.04057f
C783 VDDA.t55 GNDA 0.067616f
C784 VDDA.t400 GNDA 0.070433f
C785 VDDA.n95 GNDA 0.03408f
C786 VDDA.t393 GNDA 0.035498f
C787 VDDA.t57 GNDA 0.04057f
C788 VDDA.t5 GNDA 0.04057f
C789 VDDA.t185 GNDA 0.067616f
C790 VDDA.t158 GNDA 0.070433f
C791 VDDA.n96 GNDA 0.012084f
C792 VDDA.n97 GNDA 0.03408f
C793 VDDA.t371 GNDA 0.035498f
C794 VDDA.t234 GNDA 0.04057f
C795 VDDA.t414 GNDA 0.04057f
C796 VDDA.t387 GNDA 0.062748f
C797 VDDA.t219 GNDA 0.295215f
C798 VDDA.t51 GNDA 0.262871f
C799 VDDA.t260 GNDA 0.015182f
C800 VDDA.n99 GNDA 0.111819f
C801 VDDA.t52 GNDA 0.022637f
C802 VDDA.n101 GNDA 0.020298f
C803 VDDA.n103 GNDA 0.015026f
C804 VDDA.n104 GNDA 0.015026f
C805 VDDA.n106 GNDA 0.029081f
C806 VDDA.n108 GNDA 0.291956f
C807 VDDA.t196 GNDA 0.207195f
C808 VDDA.t26 GNDA 0.262871f
C809 VDDA.t262 GNDA 0.015182f
C810 VDDA.n110 GNDA 0.111819f
C811 VDDA.n111 GNDA 0.015026f
C812 VDDA.n112 GNDA 0.015026f
C813 VDDA.t27 GNDA 0.022637f
C814 VDDA.n114 GNDA 0.029081f
C815 VDDA.n116 GNDA 0.291956f
C816 VDDA.n118 GNDA 0.020298f
C817 VDDA.n121 GNDA 0.011092f
C818 VDDA.n127 GNDA 0.011011f
C819 VDDA.n128 GNDA 0.155753f
C820 VDDA.n129 GNDA 0.116379f
C821 VDDA.n130 GNDA 0.010559f
C822 VDDA.n134 GNDA 0.013807f
C823 VDDA.n152 GNDA 0.013807f
C824 VDDA.n158 GNDA 0.013807f
C825 VDDA.n179 GNDA 0.013807f
C826 VDDA.n197 GNDA 0.013807f
C827 VDDA.n203 GNDA 0.013807f
C828 VDDA.n219 GNDA 0.013807f
C829 VDDA.n236 GNDA 0.014591f
C830 VDDA.n238 GNDA 0.014591f
C831 VDDA.n245 GNDA 0.013807f
C832 VDDA.n252 GNDA 0.013807f
C833 VDDA.n271 GNDA 0.014592f
C834 VDDA.n291 GNDA 0.013807f
C835 VDDA.n299 GNDA 0.010627f
C836 VDDA.n300 GNDA 0.278635f
C837 VDDA.n301 GNDA 0.021219f
C838 VDDA.n302 GNDA 0.021219f
C839 VDDA.n307 GNDA 0.012021f
C840 VDDA.n308 GNDA 0.012021f
C841 VDDA.n316 GNDA 0.021219f
C842 VDDA.t160 GNDA 0.089833f
C843 VDDA.n321 GNDA 0.015026f
C844 VDDA.t205 GNDA 0.032579f
C845 VDDA.n324 GNDA 0.035681f
C846 VDDA.t385 GNDA 0.089833f
C847 VDDA.n329 GNDA 0.015026f
C848 VDDA.n331 GNDA 0.021219f
C849 VDDA.n334 GNDA 0.019297f
C850 VDDA.n335 GNDA 0.021219f
C851 VDDA.n338 GNDA 0.010191f
C852 VDDA.t426 GNDA 0.01093f
C853 VDDA.n341 GNDA 0.082659f
C854 VDDA.n343 GNDA 0.019319f
C855 VDDA.t106 GNDA 0.010733f
C856 VDDA.n344 GNDA 0.032198f
C857 VDDA.n345 GNDA 0.010733f
C858 VDDA.t3 GNDA 0.302769f
C859 VDDA.n349 GNDA 0.010733f
C860 VDDA.t4 GNDA 0.010733f
C861 VDDA.n350 GNDA 0.032198f
C862 VDDA.t416 GNDA 0.010733f
C863 VDDA.n351 GNDA 0.032198f
C864 VDDA.n353 GNDA 0.019498f
C865 VDDA.n354 GNDA 0.019319f
C866 VDDA.n355 GNDA 0.010733f
C867 VDDA.n356 GNDA 0.010733f
C868 VDDA.n357 GNDA 0.019319f
C869 VDDA.n358 GNDA 0.022774f
C870 VDDA.t428 GNDA 0.507152f
C871 VDDA.t424 GNDA 0.507152f
C872 VDDA.t423 GNDA 0.481819f
C873 VDDA.n363 GNDA 0.932542f
C874 VDDA.n364 GNDA 0.492381f
C875 VDDA.t429 GNDA 0.475945f
C876 VDDA.n365 GNDA 0.584333f
C877 VDDA.t188 GNDA 0.239983f
C878 VDDA.t61 GNDA 0.252862f
C879 VDDA.t135 GNDA 0.252862f
C880 VDDA.t25 GNDA 0.252862f
C881 VDDA.t184 GNDA 0.252862f
C882 VDDA.t94 GNDA 0.252862f
C883 VDDA.t251 GNDA 0.252862f
C884 VDDA.t143 GNDA 0.252862f
C885 VDDA.t129 GNDA 0.240853f
C886 VDDA.t366 GNDA 0.11602f
C887 VDDA.n366 GNDA 0.149649f
C888 VDDA.t86 GNDA 0.263063f
C889 VDDA.t127 GNDA 0.241865f
C890 VDDA.t128 GNDA 0.252862f
C891 VDDA.t95 GNDA 0.252862f
C892 VDDA.t138 GNDA 0.252862f
C893 VDDA.t187 GNDA 0.252862f
C894 VDDA.t122 GNDA 0.252862f
C895 VDDA.t62 GNDA 0.252862f
C896 VDDA.t102 GNDA 0.252862f
C897 VDDA.t85 GNDA 0.390571f
C898 VDDA.n367 GNDA 0.593893f
C899 VDDA.n369 GNDA 0.114767f
C900 VDDA.n370 GNDA 0.016692f
C901 VDDA.n371 GNDA 0.016565f
C902 VDDA.n373 GNDA 0.114767f
C903 VDDA.n375 GNDA 0.114767f
C904 VDDA.n377 GNDA 0.114767f
C905 VDDA.n379 GNDA 0.114767f
C906 VDDA.n381 GNDA 0.114767f
C907 VDDA.n383 GNDA 0.114767f
C908 VDDA.n385 GNDA 0.114767f
C909 VDDA.n387 GNDA 0.114767f
C910 VDDA.n389 GNDA 0.114767f
C911 VDDA.n390 GNDA 0.016692f
C912 VDDA.n391 GNDA 0.016565f
C913 VDDA.n393 GNDA 0.114767f
C914 VDDA.n395 GNDA 0.114767f
C915 VDDA.n397 GNDA 0.114767f
C916 VDDA.n399 GNDA 0.114767f
C917 VDDA.n401 GNDA 0.114767f
C918 VDDA.n403 GNDA 0.114767f
C919 VDDA.n405 GNDA 0.114767f
C920 VDDA.n407 GNDA 0.156386f
C921 VDDA.t335 GNDA 0.010701f
C922 VDDA.n408 GNDA 0.05019f
C923 VDDA.t337 GNDA 0.014933f
C924 VDDA.n410 GNDA 0.016692f
C925 VDDA.n411 GNDA 0.052919f
C926 VDDA.t336 GNDA 0.044553f
C927 VDDA.t87 GNDA 0.036062f
C928 VDDA.t243 GNDA 0.036062f
C929 VDDA.t92 GNDA 0.036062f
C930 VDDA.t39 GNDA 0.036062f
C931 VDDA.t79 GNDA 0.036062f
C932 VDDA.t197 GNDA 0.036062f
C933 VDDA.t199 GNDA 0.036062f
C934 VDDA.t338 GNDA 0.036062f
C935 VDDA.t96 GNDA 0.036062f
C936 VDDA.t178 GNDA 0.036062f
C937 VDDA.t369 GNDA 0.036062f
C938 VDDA.t118 GNDA 0.036062f
C939 VDDA.t404 GNDA 0.036062f
C940 VDDA.t9 GNDA 0.036062f
C941 VDDA.t7 GNDA 0.036062f
C942 VDDA.t241 GNDA 0.036062f
C943 VDDA.t227 GNDA 0.036062f
C944 VDDA.t120 GNDA 0.036062f
C945 VDDA.t274 GNDA 0.054796f
C946 VDDA.n412 GNDA 0.045681f
C947 VDDA.t275 GNDA 0.014933f
C948 VDDA.n413 GNDA 0.016565f
C949 VDDA.n414 GNDA 0.012752f
C950 VDDA.t273 GNDA 0.010701f
C951 VDDA.n415 GNDA 0.035445f
C952 VDDA.n416 GNDA 0.116669f
C953 VDDA.n417 GNDA 0.116669f
C954 VDDA.t267 GNDA 0.010701f
C955 VDDA.n418 GNDA 0.047263f
C956 VDDA.t269 GNDA 0.014933f
C957 VDDA.n420 GNDA 0.016692f
C958 VDDA.n421 GNDA 0.055559f
C959 VDDA.t268 GNDA 0.044919f
C960 VDDA.t59 GNDA 0.036062f
C961 VDDA.t213 GNDA 0.036062f
C962 VDDA.t239 GNDA 0.036062f
C963 VDDA.t362 GNDA 0.036062f
C964 VDDA.t348 GNDA 0.036062f
C965 VDDA.t402 GNDA 0.036062f
C966 VDDA.t64 GNDA 0.036062f
C967 VDDA.t358 GNDA 0.036062f
C968 VDDA.t354 GNDA 0.036062f
C969 VDDA.t352 GNDA 0.036062f
C970 VDDA.t350 GNDA 0.036062f
C971 VDDA.t249 GNDA 0.036062f
C972 VDDA.t180 GNDA 0.036062f
C973 VDDA.t356 GNDA 0.036062f
C974 VDDA.t360 GNDA 0.036062f
C975 VDDA.t346 GNDA 0.036062f
C976 VDDA.t344 GNDA 0.036062f
C977 VDDA.t49 GNDA 0.036062f
C978 VDDA.t288 GNDA 0.053961f
C979 VDDA.n422 GNDA 0.043511f
C980 VDDA.t289 GNDA 0.014933f
C981 VDDA.n423 GNDA 0.016565f
C982 VDDA.n424 GNDA 0.012752f
C983 VDDA.t287 GNDA 0.010701f
C984 VDDA.n425 GNDA 0.035445f
C985 VDDA.n426 GNDA 0.352302f
C986 VDDA.n427 GNDA 0.244315f
C987 VDDA.n430 GNDA 0.01434f
C988 VDDA.t216 GNDA 0.013416f
C989 VDDA.t285 GNDA 0.013416f
C990 VDDA.n432 GNDA 0.028096f
C991 VDDA.t224 GNDA 0.013416f
C992 VDDA.t376 GNDA 0.013416f
C993 VDDA.n435 GNDA 0.028096f
C994 VDDA.t71 GNDA 0.013416f
C995 VDDA.t153 GNDA 0.013416f
C996 VDDA.n438 GNDA 0.028096f
C997 VDDA.t151 GNDA 0.013416f
C998 VDDA.t18 GNDA 0.013416f
C999 VDDA.n441 GNDA 0.028096f
C1000 VDDA.n443 GNDA 0.011866f
C1001 VDDA.n444 GNDA 0.029992f
C1002 VDDA.t374 GNDA 0.013416f
C1003 VDDA.n446 GNDA 0.028096f
C1004 VDDA.n447 GNDA 0.011866f
C1005 VDDA.n448 GNDA 0.023208f
C1006 VDDA.n449 GNDA 0.011866f
C1007 VDDA.t324 GNDA 0.019235f
C1008 VDDA.n450 GNDA 0.011866f
C1009 VDDA.t308 GNDA 0.024611f
C1010 VDDA.n451 GNDA 0.014765f
C1011 VDDA.n452 GNDA 0.14751f
C1012 VDDA.t307 GNDA 0.361287f
C1013 VDDA.t0 GNDA 0.182778f
C1014 VDDA.t254 GNDA 0.182778f
C1015 VDDA.t66 GNDA 0.182778f
C1016 VDDA.t217 GNDA 0.182778f
C1017 VDDA.t322 GNDA 0.207383f
C1018 VDDA.n456 GNDA 0.010733f
C1019 VDDA.t283 GNDA 0.053163f
C1020 VDDA.n457 GNDA 0.018757f
C1021 VDDA.t286 GNDA 0.013416f
C1022 VDDA.n458 GNDA 0.040248f
C1023 VDDA.n459 GNDA 0.019204f
C1024 VDDA.n460 GNDA 0.019319f
C1025 VDDA.n461 GNDA 0.010733f
C1026 VDDA.n462 GNDA 0.010733f
C1027 VDDA.n463 GNDA 0.019319f
C1028 VDDA.n465 GNDA 0.019319f
C1029 VDDA.n466 GNDA 0.018384f
C1030 VDDA.n467 GNDA 0.010733f
C1031 VDDA.n468 GNDA 0.291742f
C1032 VDDA.t265 GNDA 0.140598f
C1033 VDDA.t284 GNDA 0.091389f
C1034 VDDA.t263 GNDA 0.108964f
C1035 VDDA.t264 GNDA 0.123024f
C1036 VDDA.t215 GNDA 0.091389f
C1037 VDDA.t134 GNDA 0.140598f
C1038 VDDA.t375 GNDA 0.091389f
C1039 VDDA.t28 GNDA 0.101934f
C1040 VDDA.t266 GNDA 0.130053f
C1041 VDDA.t223 GNDA 0.179263f
C1042 VDDA.t152 GNDA 0.189808f
C1043 VDDA.t279 GNDA 0.019235f
C1044 VDDA.n469 GNDA 0.011866f
C1045 VDDA.n470 GNDA 0.023208f
C1046 VDDA.n471 GNDA 0.014662f
C1047 VDDA.n472 GNDA 0.040371f
C1048 VDDA.n473 GNDA 0.151496f
C1049 VDDA.t70 GNDA 0.115994f
C1050 VDDA.t277 GNDA 0.115994f
C1051 VDDA.t258 GNDA 0.115994f
C1052 VDDA.t17 GNDA 0.091389f
C1053 VDDA.t35 GNDA 0.140598f
C1054 VDDA.t150 GNDA 0.091389f
C1055 VDDA.t229 GNDA 0.108964f
C1056 VDDA.t232 GNDA 0.123024f
C1057 VDDA.t373 GNDA 0.091389f
C1058 VDDA.t271 GNDA 0.140598f
C1059 VDDA.t294 GNDA 0.115994f
C1060 VDDA.t272 GNDA 0.024611f
C1061 VDDA.n474 GNDA 0.011866f
C1062 VDDA.n475 GNDA 0.023208f
C1063 VDDA.n476 GNDA 0.014765f
C1064 VDDA.n477 GNDA 0.047967f
C1065 VDDA.n478 GNDA 0.137025f
C1066 VDDA.n479 GNDA 0.010733f
C1067 VDDA.n480 GNDA 0.010733f
C1068 VDDA.t293 GNDA 0.054251f
C1069 VDDA.t295 GNDA 0.026832f
C1070 VDDA.n481 GNDA 0.040248f
C1071 VDDA.n482 GNDA 0.019204f
C1072 VDDA.n483 GNDA 0.010733f
C1073 VDDA.n484 GNDA 0.019319f
C1074 VDDA.n485 GNDA 0.019319f
C1075 VDDA.n487 GNDA 0.019319f
C1076 VDDA.n488 GNDA 0.037907f
C1077 VDDA.n490 GNDA 0.110869f
C1078 VDDA.n491 GNDA 0.133921f
C1079 VDDA.n492 GNDA 0.040371f
C1080 VDDA.n493 GNDA 0.014662f
C1081 VDDA.n494 GNDA 0.023208f
C1082 VDDA.n495 GNDA 0.033219f
C1083 VDDA.n496 GNDA 0.096513f
C1084 VDDA.n497 GNDA 0.096974f
C1085 VDDA.n505 GNDA 0.094042f
C1086 VDDA.n512 GNDA 0.094042f
C1087 VDDA.n519 GNDA 0.094042f
C1088 VDDA.n526 GNDA 0.094042f
C1089 VDDA.n536 GNDA 0.045983f
C1090 VDDA.n537 GNDA 0.136853f
C1091 VDDA.t290 GNDA 0.061414f
C1092 VDDA.n538 GNDA 0.023542f
C1093 VDDA.t34 GNDA 0.012879f
C1094 VDDA.t133 GNDA 0.012879f
C1095 VDDA.n539 GNDA 0.050112f
C1096 VDDA.t137 GNDA 0.012879f
C1097 VDDA.t420 GNDA 0.012879f
C1098 VDDA.n540 GNDA 0.050112f
C1099 VDDA.t32 GNDA 0.012879f
C1100 VDDA.t253 GNDA 0.012879f
C1101 VDDA.n541 GNDA 0.050112f
C1102 VDDA.t126 GNDA 0.012879f
C1103 VDDA.t24 GNDA 0.012879f
C1104 VDDA.n542 GNDA 0.050112f
C1105 VDDA.t183 GNDA 0.012879f
C1106 VDDA.t368 GNDA 0.012879f
C1107 VDDA.n543 GNDA 0.050112f
C1108 VDDA.t418 GNDA 0.012879f
C1109 VDDA.t104 GNDA 0.012879f
C1110 VDDA.n544 GNDA 0.050112f
C1111 VDDA.t131 GNDA 0.012879f
C1112 VDDA.t142 GNDA 0.012879f
C1113 VDDA.n545 GNDA 0.050112f
C1114 VDDA.t124 GNDA 0.012879f
C1115 VDDA.t140 GNDA 0.012879f
C1116 VDDA.n546 GNDA 0.050112f
C1117 VDDA.n548 GNDA 0.012108f
C1118 VDDA.n556 GNDA 0.014936f
C1119 VDDA.n557 GNDA 0.014936f
C1120 VDDA.n559 GNDA 0.015026f
C1121 VDDA.n561 GNDA 0.017155f
C1122 VDDA.n562 GNDA 0.012108f
C1123 VDDA.n564 GNDA 0.015026f
C1124 VDDA.n567 GNDA 0.015026f
C1125 VDDA.n568 GNDA 0.015026f
C1126 VDDA.n569 GNDA 0.012108f
C1127 VDDA.n570 GNDA 0.016194f
C1128 VDDA.n572 GNDA 0.120421f
C1129 VDDA.t291 GNDA 0.127719f
C1130 VDDA.t33 GNDA 0.131368f
C1131 VDDA.t132 GNDA 0.131368f
C1132 VDDA.t136 GNDA 0.131368f
C1133 VDDA.t419 GNDA 0.131368f
C1134 VDDA.t31 GNDA 0.131368f
C1135 VDDA.t252 GNDA 0.131368f
C1136 VDDA.t125 GNDA 0.131368f
C1137 VDDA.t23 GNDA 0.131368f
C1138 VDDA.t182 GNDA 0.131368f
C1139 VDDA.t367 GNDA 0.131368f
C1140 VDDA.t417 GNDA 0.131368f
C1141 VDDA.t103 GNDA 0.131368f
C1142 VDDA.t130 GNDA 0.131368f
C1143 VDDA.t141 GNDA 0.131368f
C1144 VDDA.t123 GNDA 0.131368f
C1145 VDDA.t139 GNDA 0.131368f
C1146 VDDA.t313 GNDA 0.127719f
C1147 VDDA.n576 GNDA 0.012108f
C1148 VDDA.n577 GNDA 0.015026f
C1149 VDDA.n580 GNDA 0.015026f
C1150 VDDA.n581 GNDA 0.014936f
C1151 VDDA.n583 GNDA 0.015026f
C1152 VDDA.n584 GNDA 0.015026f
C1153 VDDA.n585 GNDA 0.014936f
C1154 VDDA.n587 GNDA 0.018116f
C1155 VDDA.n589 GNDA 0.120421f
C1156 VDDA.n591 GNDA 0.017155f
C1157 VDDA.t312 GNDA 0.061414f
C1158 VDDA.n592 GNDA 0.024804f
C1159 VDDA.n593 GNDA 0.245437f
C1160 VDDA.n594 GNDA 0.172269f
C1161 VDDA.n595 GNDA 0.172269f
C1162 VDDA.n596 GNDA 0.172269f
C1163 VDDA.n597 GNDA 0.172269f
C1164 VDDA.n598 GNDA 0.172269f
C1165 VDDA.n599 GNDA 0.172269f
C1166 VDDA.n600 GNDA 0.172269f
C1167 VDDA.n601 GNDA 0.145265f
C1168 VDDA.n602 GNDA 0.143252f
C1169 VDDA.n603 GNDA 0.016692f
C1170 VDDA.n604 GNDA 0.017553f
C1171 VDDA.n605 GNDA 0.054633f
C1172 VDDA.t334 GNDA 0.017035f
C1173 VDDA.n607 GNDA 0.01768f
C1174 VDDA.n608 GNDA 0.053749f
C1175 VDDA.t333 GNDA 0.043724f
C1176 VDDA.t222 GNDA 0.033057f
C1177 VDDA.t63 GNDA 0.033057f
C1178 VDDA.t316 GNDA 0.051888f
C1179 VDDA.n609 GNDA 0.042579f
C1180 VDDA.t317 GNDA 0.014933f
C1181 VDDA.n610 GNDA 0.016565f
C1182 VDDA.n611 GNDA 0.012635f
C1183 VDDA.n612 GNDA 0.041154f
C1184 VDDA.n613 GNDA 0.386664f
C1185 VDDA.n614 GNDA 0.124241f
C1186 VDDA.n616 GNDA 0.05083f
C1187 VDDA.n617 GNDA 0.01682f
C1188 VDDA.n618 GNDA 0.016565f
C1189 VDDA.t311 GNDA 0.014933f
C1190 VDDA.n621 GNDA 0.05083f
C1191 VDDA.n623 GNDA 0.05083f
C1192 VDDA.n625 GNDA 0.05083f
C1193 VDDA.n627 GNDA 0.05083f
C1194 VDDA.n629 GNDA 0.05083f
C1195 VDDA.n630 GNDA 0.01682f
C1196 VDDA.n631 GNDA 0.016565f
C1197 VDDA.t305 GNDA 0.014933f
C1198 VDDA.n634 GNDA 0.05083f
C1199 VDDA.n636 GNDA 0.05083f
C1200 VDDA.n638 GNDA 0.05083f
C1201 VDDA.n640 GNDA 0.062795f
C1202 VDDA.n641 GNDA 0.021288f
C1203 VDDA.n642 GNDA 0.02827f
C1204 VDDA.n643 GNDA 0.01682f
C1205 VDDA.n644 GNDA 0.052085f
C1206 VDDA.t304 GNDA 0.042382f
C1207 VDDA.t148 GNDA 0.033057f
C1208 VDDA.t406 GNDA 0.033057f
C1209 VDDA.t156 GNDA 0.033057f
C1210 VDDA.t168 GNDA 0.033057f
C1211 VDDA.t146 GNDA 0.033057f
C1212 VDDA.t381 GNDA 0.033057f
C1213 VDDA.t174 GNDA 0.033057f
C1214 VDDA.t383 GNDA 0.033057f
C1215 VDDA.t395 GNDA 0.033057f
C1216 VDDA.t194 GNDA 0.033057f
C1217 VDDA.t281 GNDA 0.051888f
C1218 VDDA.n645 GNDA 0.042579f
C1219 VDDA.t282 GNDA 0.014933f
C1220 VDDA.n646 GNDA 0.016565f
C1221 VDDA.n647 GNDA 0.02827f
C1222 VDDA.n648 GNDA 0.020374f
C1223 VDDA.n649 GNDA 0.034345f
C1224 VDDA.n650 GNDA 0.034345f
C1225 VDDA.n651 GNDA 0.020374f
C1226 VDDA.n652 GNDA 0.02827f
C1227 VDDA.n653 GNDA 0.01682f
C1228 VDDA.n654 GNDA 0.052085f
C1229 VDDA.t310 GNDA 0.042382f
C1230 VDDA.t379 GNDA 0.033057f
C1231 VDDA.t192 GNDA 0.033057f
C1232 VDDA.t377 GNDA 0.033057f
C1233 VDDA.t172 GNDA 0.033057f
C1234 VDDA.t170 GNDA 0.033057f
C1235 VDDA.t410 GNDA 0.033057f
C1236 VDDA.t397 GNDA 0.033057f
C1237 VDDA.t412 GNDA 0.033057f
C1238 VDDA.t408 GNDA 0.033057f
C1239 VDDA.t154 GNDA 0.033057f
C1240 VDDA.t301 GNDA 0.051888f
C1241 VDDA.n655 GNDA 0.042579f
C1242 VDDA.t302 GNDA 0.014933f
C1243 VDDA.n656 GNDA 0.016565f
C1244 VDDA.n657 GNDA 0.02827f
C1245 VDDA.n658 GNDA 0.020374f
C1246 VDDA.n659 GNDA 0.184748f
C1247 VDDA.n660 GNDA 0.120257f
C1248 VDDA.t331 GNDA 0.010733f
C1249 VDDA.n664 GNDA 0.032198f
C1250 VDDA.n665 GNDA 0.019319f
C1251 VDDA.n666 GNDA 0.010733f
C1252 VDDA.t297 GNDA 0.133837f
C1253 VDDA.n668 GNDA 0.010733f
C1254 VDDA.n669 GNDA 0.013254f
C1255 VDDA.t299 GNDA 0.010733f
C1256 VDDA.n671 GNDA 0.030052f
C1257 VDDA.n673 GNDA 0.010733f
C1258 VDDA.n674 GNDA 0.030052f
C1259 VDDA.t101 GNDA 0.010733f
C1260 VDDA.t42 GNDA 0.010733f
C1261 VDDA.n677 GNDA 0.031032f
C1262 VDDA.n678 GNDA 0.043667f
C1263 VDDA.t84 GNDA 0.010733f
C1264 VDDA.t330 GNDA 0.010733f
C1265 VDDA.n680 GNDA 0.031032f
C1266 VDDA.n681 GNDA 0.043667f
C1267 VDDA.t22 GNDA 0.010733f
C1268 VDDA.t298 GNDA 0.010733f
C1269 VDDA.n700 GNDA 0.031032f
C1270 VDDA.t30 GNDA 0.010733f
C1271 VDDA.t422 GNDA 0.010733f
C1272 VDDA.n703 GNDA 0.031032f
C1273 VDDA.n705 GNDA 0.027606f
C1274 VDDA.n706 GNDA 0.014649f
C1275 VDDA.n708 GNDA 0.017387f
C1276 VDDA.t318 GNDA 0.053498f
C1277 VDDA.n709 GNDA 0.02104f
C1278 VDDA.n710 GNDA 0.010733f
C1279 VDDA.n711 GNDA 0.019319f
C1280 VDDA.n712 GNDA 0.010733f
C1281 VDDA.n713 GNDA 0.010733f
C1282 VDDA.t21 GNDA 0.136949f
C1283 VDDA.t421 GNDA 0.136949f
C1284 VDDA.t29 GNDA 0.136949f
C1285 VDDA.t245 GNDA 0.136949f
C1286 VDDA.t319 GNDA 0.133837f
C1287 VDDA.n714 GNDA 0.121387f
C1288 VDDA.n716 GNDA 0.010733f
C1289 VDDA.n717 GNDA 0.019319f
C1290 VDDA.n718 GNDA 0.019495f
C1291 VDDA.n719 GNDA 0.032198f
C1292 VDDA.t320 GNDA 0.021465f
C1293 VDDA.t246 GNDA 0.010733f
C1294 VDDA.n720 GNDA 0.031032f
C1295 VDDA.n721 GNDA 0.044221f
C1296 VDDA.n728 GNDA 0.041521f
C1297 VDDA.n735 GNDA 0.043667f
C1298 VDDA.n743 GNDA 0.043667f
C1299 VDDA.t392 GNDA 0.010733f
C1300 VDDA.n744 GNDA 0.031032f
C1301 VDDA.t327 GNDA 0.021465f
C1302 VDDA.n745 GNDA 0.032198f
C1303 VDDA.t296 GNDA 0.050481f
C1304 VDDA.t325 GNDA 0.050481f
C1305 VDDA.n747 GNDA 0.022742f
C1306 VDDA.n748 GNDA 0.038755f
C1307 VDDA.n749 GNDA 0.032198f
C1308 VDDA.n750 GNDA 0.036511f
C1309 VDDA.n752 GNDA 0.130724f
C1310 VDDA.t326 GNDA 0.133837f
C1311 VDDA.t391 GNDA 0.136949f
C1312 VDDA.t100 GNDA 0.136949f
C1313 VDDA.t41 GNDA 0.136949f
C1314 VDDA.t83 GNDA 0.136949f
C1315 VDDA.t329 GNDA 0.133837f
C1316 VDDA.n753 GNDA 0.019498f
C1317 VDDA.n755 GNDA 0.019319f
C1318 VDDA.n756 GNDA 0.010733f
C1319 VDDA.n758 GNDA 0.121387f
C1320 VDDA.n760 GNDA 0.021606f
C1321 VDDA.t328 GNDA 0.053498f
C1322 VDDA.n761 GNDA 0.018557f
C1323 VDDA.n768 GNDA 0.043945f
C1324 VDDA.n769 GNDA 0.202191f
C1325 VDDA.n770 GNDA 0.082446f
C1326 VDDA.n771 GNDA 0.019319f
C1327 VDDA.t46 GNDA 0.010733f
C1328 VDDA.n772 GNDA 0.032198f
C1329 VDDA.n773 GNDA 0.010733f
C1330 VDDA.t45 GNDA 0.316078f
C1331 VDDA.t203 GNDA 0.342695f
C1332 VDDA.n774 GNDA 0.010733f
C1333 VDDA.n776 GNDA 0.019319f
C1334 VDDA.n777 GNDA 0.019498f
C1335 VDDA.n779 GNDA 0.259517f
C1336 VDDA.n781 GNDA 0.022774f
C1337 VDDA.n784 GNDA 0.010629f
C1338 VDDA.n795 GNDA 0.012338f
C1339 VDDA.n796 GNDA 0.022774f
C1340 VDDA.n797 GNDA 0.010733f
C1341 VDDA.n798 GNDA 0.019319f
C1342 VDDA.n800 GNDA 0.019319f
C1343 VDDA.n801 GNDA 0.019498f
C1344 VDDA.n803 GNDA 0.259517f
C1345 VDDA.t105 GNDA 0.259517f
C1346 VDDA.t114 GNDA 0.089833f
C1347 VDDA.t386 GNDA 0.022637f
C1348 VDDA.n811 GNDA 0.020906f
C1349 VDDA.n812 GNDA 0.015026f
C1350 VDDA.n813 GNDA 0.015026f
C1351 VDDA.n816 GNDA 0.129758f
C1352 VDDA.n818 GNDA 0.015026f
C1353 VDDA.n820 GNDA 0.015026f
C1354 VDDA.t248 GNDA 0.022637f
C1355 VDDA.n822 GNDA 0.020906f
C1356 VDDA.n824 GNDA 0.129758f
C1357 VDDA.t162 GNDA 0.089833f
C1358 VDDA.t247 GNDA 0.089833f
C1359 VDDA.t163 GNDA 0.022637f
C1360 VDDA.n827 GNDA 0.018927f
C1361 VDDA.n828 GNDA 0.015026f
C1362 VDDA.n829 GNDA 0.015026f
C1363 VDDA.n832 GNDA 0.182993f
C1364 VDDA.n834 GNDA 0.010733f
C1365 VDDA.t69 GNDA 0.010733f
C1366 VDDA.n835 GNDA 0.032198f
C1367 VDDA.n836 GNDA 0.019498f
C1368 VDDA.n837 GNDA 0.010733f
C1369 VDDA.n838 GNDA 0.019319f
C1370 VDDA.n840 GNDA 0.019319f
C1371 VDDA.n841 GNDA 0.022774f
C1372 VDDA.n843 GNDA 0.010733f
C1373 VDDA.t113 GNDA 0.010733f
C1374 VDDA.n844 GNDA 0.032198f
C1375 VDDA.n845 GNDA 0.022774f
C1376 VDDA.n846 GNDA 0.010733f
C1377 VDDA.n847 GNDA 0.019319f
C1378 VDDA.n849 GNDA 0.019319f
C1379 VDDA.n850 GNDA 0.019498f
C1380 VDDA.n852 GNDA 0.282807f
C1381 VDDA.t68 GNDA 0.259517f
C1382 VDDA.n853 GNDA 0.010733f
C1383 VDDA.n855 GNDA 0.019319f
C1384 VDDA.n856 GNDA 0.019498f
C1385 VDDA.n858 GNDA 0.259517f
C1386 VDDA.n860 GNDA 0.022774f
C1387 VDDA.n888 GNDA 0.021219f
C1388 VDDA.n890 GNDA 0.015026f
C1389 VDDA.t115 GNDA 0.022637f
C1390 VDDA.n892 GNDA 0.020906f
C1391 VDDA.n894 GNDA 0.129758f
C1392 VDDA.t161 GNDA 0.022637f
C1393 VDDA.n895 GNDA 0.020906f
C1394 VDDA.n896 GNDA 0.015026f
C1395 VDDA.n897 GNDA 0.015026f
C1396 VDDA.t109 GNDA 0.079851f
C1397 VDDA.t204 GNDA 0.083178f
C1398 VDDA.n900 GNDA 0.129758f
C1399 VDDA.n902 GNDA 0.021219f
C1400 VDDA.n910 GNDA 0.020819f
C1401 VDDA.n912 GNDA 0.015026f
C1402 VDDA.t110 GNDA 0.022526f
C1403 VDDA.n914 GNDA 0.020906f
C1404 VDDA.n916 GNDA 0.176338f
C1405 VDDA.t82 GNDA 0.022637f
C1406 VDDA.n923 GNDA 0.020906f
C1407 VDDA.n924 GNDA 0.015026f
C1408 VDDA.n925 GNDA 0.015026f
C1409 VDDA.n929 GNDA 0.015026f
C1410 VDDA.n931 GNDA 0.015026f
C1411 VDDA.t231 GNDA 0.022637f
C1412 VDDA.n933 GNDA 0.020906f
C1413 VDDA.n935 GNDA 0.196301f
C1414 VDDA.t81 GNDA 0.16303f
C1415 VDDA.t89 GNDA 0.346022f
C1416 VDDA.t2 GNDA 0.346022f
C1417 VDDA.t166 GNDA 0.16303f
C1418 VDDA.n938 GNDA 0.012482f
C1419 VDDA.n939 GNDA 0.023612f
C1420 VDDA.n940 GNDA 0.02826f
C1421 VDDA.n941 GNDA 0.012482f
C1422 VDDA.n943 GNDA 0.023612f
C1423 VDDA.t14 GNDA 0.022648f
C1424 VDDA.n946 GNDA 0.023538f
C1425 VDDA.n949 GNDA 0.012482f
C1426 VDDA.n950 GNDA 0.023612f
C1427 VDDA.n951 GNDA 0.023538f
C1428 VDDA.n952 GNDA 0.012482f
C1429 VDDA.n954 GNDA 0.023612f
C1430 VDDA.t208 GNDA 0.022648f
C1431 VDDA.n957 GNDA 0.02826f
C1432 VDDA.n959 GNDA 0.179665f
C1433 VDDA.t13 GNDA 0.16303f
C1434 VDDA.t238 GNDA 0.346022f
C1435 VDDA.t189 GNDA 0.346022f
C1436 VDDA.t256 GNDA 0.16303f
C1437 VDDA.t257 GNDA 0.022637f
C1438 VDDA.n960 GNDA 0.020906f
C1439 VDDA.n961 GNDA 0.015026f
C1440 VDDA.n962 GNDA 0.015026f
C1441 VDDA.n966 GNDA 0.015026f
C1442 VDDA.n968 GNDA 0.015026f
C1443 VDDA.t365 GNDA 0.022637f
C1444 VDDA.n970 GNDA 0.020906f
C1445 VDDA.n972 GNDA 0.182993f
C1446 VDDA.n974 GNDA 0.021219f
C1447 VDDA.n975 GNDA 0.010283f
C1448 VDDA.n1005 GNDA 0.010283f
C1449 VDDA.n1007 GNDA 0.245974f
C1450 a_5970_4630.t9 GNDA 0.030769f
C1451 a_5970_4630.n0 GNDA 0.124795f
C1452 a_5970_4630.t0 GNDA 0.020325f
C1453 a_5970_4630.t1 GNDA 0.020325f
C1454 a_5970_4630.t5 GNDA 0.020325f
C1455 a_5970_4630.n1 GNDA 0.044943f
C1456 a_5970_4630.t4 GNDA 0.020325f
C1457 a_5970_4630.t7 GNDA 0.020325f
C1458 a_5970_4630.n2 GNDA 0.044943f
C1459 a_5970_4630.t8 GNDA 0.077457f
C1460 a_5970_4630.t6 GNDA 0.030769f
C1461 a_5970_4630.n3 GNDA 0.097952f
C1462 a_5970_4630.n4 GNDA 0.087903f
C1463 a_5970_4630.n5 GNDA 0.089425f
C1464 a_5970_4630.t11 GNDA 0.050813f
C1465 a_5970_4630.t2 GNDA 0.050813f
C1466 a_5970_4630.n6 GNDA 0.295522f
C1467 a_5970_4630.t12 GNDA 0.050813f
C1468 a_5970_4630.t3 GNDA 0.050813f
C1469 a_5970_4630.n7 GNDA 0.144587f
C1470 a_5970_4630.n8 GNDA 0.360746f
C1471 a_5970_4630.n9 GNDA 0.13437f
C1472 a_5970_4630.n10 GNDA 0.085474f
C1473 a_5970_4630.n11 GNDA 0.045257f
C1474 a_5970_4630.t10 GNDA 0.100208f
C1475 V_CONT.t6 GNDA 0.014802f
C1476 V_CONT.t5 GNDA 6.66921f
C1477 V_CONT.n3 GNDA 0.166549f
C1478 V_CONT.n6 GNDA 0.020725f
C1479 opamp_cell_4_0.VIN- GNDA 0.038962f
C1480 V_CONT.n9 GNDA 0.017874f
C1481 V_CONT.n11 GNDA 0.014862f
C1482 V_CONT.n12 GNDA 0.08182f
C1483 V_CONT.n13 GNDA 0.018414f
.ends

