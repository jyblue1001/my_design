magic
tech sky130A
timestamp 1725008253
<< nwell >>
rect -65 695 2225 1385
<< nmos >>
rect 55 190 105 490
rect 155 190 205 490
rect 255 190 305 490
rect 355 190 405 490
rect 455 190 505 490
rect 555 190 605 490
rect 655 190 705 490
rect 755 190 805 490
rect 855 190 905 490
rect 955 190 1005 490
rect 1155 190 1205 490
rect 1255 190 1305 490
rect 1355 190 1405 490
rect 1455 190 1505 490
rect 1555 190 1605 490
rect 1655 190 1705 490
rect 1755 190 1805 490
rect 1855 190 1905 490
rect 1955 190 2005 490
rect 2055 190 2105 490
<< pmos >>
rect 55 1215 105 1365
rect 155 1215 205 1365
rect 255 1215 305 1365
rect 355 1215 405 1365
rect 455 1215 505 1365
rect 555 1215 605 1365
rect 655 1215 705 1365
rect 755 1215 805 1365
rect 855 1215 905 1365
rect 955 1215 1005 1365
rect 1155 1215 1205 1365
rect 1255 1215 1305 1365
rect 1355 1215 1405 1365
rect 1455 1215 1505 1365
rect 1555 1215 1605 1365
rect 1655 1215 1705 1365
rect 1755 1215 1805 1365
rect 1855 1215 1905 1365
rect 1955 1215 2005 1365
rect 2055 1215 2105 1365
rect 55 715 105 1015
rect 155 715 205 1015
rect 255 715 305 1015
rect 355 715 405 1015
rect 455 715 505 1015
rect 555 715 605 1015
rect 655 715 705 1015
rect 755 715 805 1015
rect 855 715 905 1015
rect 955 715 1005 1015
rect 1155 715 1205 1015
rect 1255 715 1305 1015
rect 1355 715 1405 1015
rect 1455 715 1505 1015
rect 1555 715 1605 1015
rect 1655 715 1705 1015
rect 1755 715 1805 1015
rect 1855 715 1905 1015
rect 1955 715 2005 1015
rect 2055 715 2105 1015
<< ndiff >>
rect 5 475 55 490
rect 5 205 20 475
rect 40 205 55 475
rect 5 190 55 205
rect 105 475 155 490
rect 105 205 120 475
rect 140 205 155 475
rect 105 190 155 205
rect 205 475 255 490
rect 205 205 220 475
rect 240 205 255 475
rect 205 190 255 205
rect 305 475 355 490
rect 305 205 320 475
rect 340 205 355 475
rect 305 190 355 205
rect 405 475 455 490
rect 405 205 420 475
rect 440 205 455 475
rect 405 190 455 205
rect 505 475 555 490
rect 505 205 520 475
rect 540 205 555 475
rect 505 190 555 205
rect 605 475 655 490
rect 605 205 620 475
rect 640 205 655 475
rect 605 190 655 205
rect 705 475 755 490
rect 705 205 720 475
rect 740 205 755 475
rect 705 190 755 205
rect 805 475 855 490
rect 805 205 820 475
rect 840 205 855 475
rect 805 190 855 205
rect 905 475 955 490
rect 905 205 920 475
rect 940 205 955 475
rect 905 190 955 205
rect 1005 475 1055 490
rect 1105 475 1155 490
rect 1005 205 1020 475
rect 1040 205 1055 475
rect 1105 205 1120 475
rect 1140 205 1155 475
rect 1005 190 1055 205
rect 1105 190 1155 205
rect 1205 475 1255 490
rect 1205 205 1220 475
rect 1240 205 1255 475
rect 1205 190 1255 205
rect 1305 475 1355 490
rect 1305 205 1320 475
rect 1340 205 1355 475
rect 1305 190 1355 205
rect 1405 475 1455 490
rect 1405 205 1420 475
rect 1440 205 1455 475
rect 1405 190 1455 205
rect 1505 475 1555 490
rect 1505 205 1520 475
rect 1540 205 1555 475
rect 1505 190 1555 205
rect 1605 475 1655 490
rect 1605 205 1620 475
rect 1640 205 1655 475
rect 1605 190 1655 205
rect 1705 475 1755 490
rect 1705 205 1720 475
rect 1740 205 1755 475
rect 1705 190 1755 205
rect 1805 475 1855 490
rect 1805 205 1820 475
rect 1840 205 1855 475
rect 1805 190 1855 205
rect 1905 475 1955 490
rect 1905 205 1920 475
rect 1940 205 1955 475
rect 1905 190 1955 205
rect 2005 475 2055 490
rect 2005 205 2020 475
rect 2040 205 2055 475
rect 2005 190 2055 205
rect 2105 475 2155 490
rect 2105 205 2120 475
rect 2140 205 2155 475
rect 2105 190 2155 205
<< pdiff >>
rect 5 1350 55 1365
rect 5 1230 20 1350
rect 40 1230 55 1350
rect 5 1215 55 1230
rect 105 1350 155 1365
rect 105 1230 120 1350
rect 140 1230 155 1350
rect 105 1215 155 1230
rect 205 1350 255 1365
rect 205 1230 220 1350
rect 240 1230 255 1350
rect 205 1215 255 1230
rect 305 1350 355 1365
rect 305 1230 320 1350
rect 340 1230 355 1350
rect 305 1215 355 1230
rect 405 1350 455 1365
rect 405 1230 420 1350
rect 440 1230 455 1350
rect 405 1215 455 1230
rect 505 1350 555 1365
rect 505 1230 520 1350
rect 540 1230 555 1350
rect 505 1215 555 1230
rect 605 1350 655 1365
rect 605 1230 620 1350
rect 640 1230 655 1350
rect 605 1215 655 1230
rect 705 1350 755 1365
rect 705 1230 720 1350
rect 740 1230 755 1350
rect 705 1215 755 1230
rect 805 1350 855 1365
rect 805 1230 820 1350
rect 840 1230 855 1350
rect 805 1215 855 1230
rect 905 1350 955 1365
rect 905 1230 920 1350
rect 940 1230 955 1350
rect 905 1215 955 1230
rect 1005 1350 1055 1365
rect 1105 1350 1155 1365
rect 1005 1230 1020 1350
rect 1040 1230 1055 1350
rect 1105 1230 1120 1350
rect 1140 1230 1155 1350
rect 1005 1215 1055 1230
rect 1105 1215 1155 1230
rect 1205 1350 1255 1365
rect 1205 1230 1220 1350
rect 1240 1230 1255 1350
rect 1205 1215 1255 1230
rect 1305 1350 1355 1365
rect 1305 1230 1320 1350
rect 1340 1230 1355 1350
rect 1305 1215 1355 1230
rect 1405 1350 1455 1365
rect 1405 1230 1420 1350
rect 1440 1230 1455 1350
rect 1405 1215 1455 1230
rect 1505 1350 1555 1365
rect 1505 1230 1520 1350
rect 1540 1230 1555 1350
rect 1505 1215 1555 1230
rect 1605 1350 1655 1365
rect 1605 1230 1620 1350
rect 1640 1230 1655 1350
rect 1605 1215 1655 1230
rect 1705 1350 1755 1365
rect 1705 1230 1720 1350
rect 1740 1230 1755 1350
rect 1705 1215 1755 1230
rect 1805 1350 1855 1365
rect 1805 1230 1820 1350
rect 1840 1230 1855 1350
rect 1805 1215 1855 1230
rect 1905 1350 1955 1365
rect 1905 1230 1920 1350
rect 1940 1230 1955 1350
rect 1905 1215 1955 1230
rect 2005 1350 2055 1365
rect 2005 1230 2020 1350
rect 2040 1230 2055 1350
rect 2005 1215 2055 1230
rect 2105 1350 2155 1365
rect 2105 1230 2120 1350
rect 2140 1230 2155 1350
rect 2105 1215 2155 1230
rect 5 1000 55 1015
rect 5 730 20 1000
rect 40 730 55 1000
rect 5 715 55 730
rect 105 1000 155 1015
rect 105 730 120 1000
rect 140 730 155 1000
rect 105 715 155 730
rect 205 1000 255 1015
rect 205 730 220 1000
rect 240 730 255 1000
rect 205 715 255 730
rect 305 1000 355 1015
rect 305 730 320 1000
rect 340 730 355 1000
rect 305 715 355 730
rect 405 1000 455 1015
rect 405 730 420 1000
rect 440 730 455 1000
rect 405 715 455 730
rect 505 1000 555 1015
rect 505 730 520 1000
rect 540 730 555 1000
rect 505 715 555 730
rect 605 1000 655 1015
rect 605 730 620 1000
rect 640 730 655 1000
rect 605 715 655 730
rect 705 1000 755 1015
rect 705 730 720 1000
rect 740 730 755 1000
rect 705 715 755 730
rect 805 1000 855 1015
rect 805 730 820 1000
rect 840 730 855 1000
rect 805 715 855 730
rect 905 1000 955 1015
rect 905 730 920 1000
rect 940 730 955 1000
rect 905 715 955 730
rect 1005 1000 1055 1015
rect 1105 1000 1155 1015
rect 1005 730 1020 1000
rect 1040 730 1055 1000
rect 1105 730 1120 1000
rect 1140 730 1155 1000
rect 1005 715 1055 730
rect 1105 715 1155 730
rect 1205 1000 1255 1015
rect 1205 730 1220 1000
rect 1240 730 1255 1000
rect 1205 715 1255 730
rect 1305 1000 1355 1015
rect 1305 730 1320 1000
rect 1340 730 1355 1000
rect 1305 715 1355 730
rect 1405 1000 1455 1015
rect 1405 730 1420 1000
rect 1440 730 1455 1000
rect 1405 715 1455 730
rect 1505 1000 1555 1015
rect 1505 730 1520 1000
rect 1540 730 1555 1000
rect 1505 715 1555 730
rect 1605 1000 1655 1015
rect 1605 730 1620 1000
rect 1640 730 1655 1000
rect 1605 715 1655 730
rect 1705 1000 1755 1015
rect 1705 730 1720 1000
rect 1740 730 1755 1000
rect 1705 715 1755 730
rect 1805 1000 1855 1015
rect 1805 730 1820 1000
rect 1840 730 1855 1000
rect 1805 715 1855 730
rect 1905 1000 1955 1015
rect 1905 730 1920 1000
rect 1940 730 1955 1000
rect 1905 715 1955 730
rect 2005 1000 2055 1015
rect 2005 730 2020 1000
rect 2040 730 2055 1000
rect 2005 715 2055 730
rect 2105 1000 2155 1015
rect 2105 730 2120 1000
rect 2140 730 2155 1000
rect 2105 715 2155 730
<< ndiffc >>
rect 20 205 40 475
rect 120 205 140 475
rect 220 205 240 475
rect 320 205 340 475
rect 420 205 440 475
rect 520 205 540 475
rect 620 205 640 475
rect 720 205 740 475
rect 820 205 840 475
rect 920 205 940 475
rect 1020 205 1040 475
rect 1120 205 1140 475
rect 1220 205 1240 475
rect 1320 205 1340 475
rect 1420 205 1440 475
rect 1520 205 1540 475
rect 1620 205 1640 475
rect 1720 205 1740 475
rect 1820 205 1840 475
rect 1920 205 1940 475
rect 2020 205 2040 475
rect 2120 205 2140 475
<< pdiffc >>
rect 20 1230 40 1350
rect 120 1230 140 1350
rect 220 1230 240 1350
rect 320 1230 340 1350
rect 420 1230 440 1350
rect 520 1230 540 1350
rect 620 1230 640 1350
rect 720 1230 740 1350
rect 820 1230 840 1350
rect 920 1230 940 1350
rect 1020 1230 1040 1350
rect 1120 1230 1140 1350
rect 1220 1230 1240 1350
rect 1320 1230 1340 1350
rect 1420 1230 1440 1350
rect 1520 1230 1540 1350
rect 1620 1230 1640 1350
rect 1720 1230 1740 1350
rect 1820 1230 1840 1350
rect 1920 1230 1940 1350
rect 2020 1230 2040 1350
rect 2120 1230 2140 1350
rect 20 730 40 1000
rect 120 730 140 1000
rect 220 730 240 1000
rect 320 730 340 1000
rect 420 730 440 1000
rect 520 730 540 1000
rect 620 730 640 1000
rect 720 730 740 1000
rect 820 730 840 1000
rect 920 730 940 1000
rect 1020 730 1040 1000
rect 1120 730 1140 1000
rect 1220 730 1240 1000
rect 1320 730 1340 1000
rect 1420 730 1440 1000
rect 1520 730 1540 1000
rect 1620 730 1640 1000
rect 1720 730 1740 1000
rect 1820 730 1840 1000
rect 1920 730 1940 1000
rect 2020 730 2040 1000
rect 2120 730 2140 1000
<< psubdiff >>
rect -45 475 5 490
rect -45 205 -30 475
rect -10 205 5 475
rect -45 190 5 205
rect 1055 475 1105 490
rect 1055 205 1070 475
rect 1090 205 1105 475
rect 1055 190 1105 205
rect 2155 475 2205 490
rect 2155 205 2170 475
rect 2190 205 2205 475
rect 2155 190 2205 205
<< nsubdiff >>
rect -45 1350 5 1365
rect -45 1230 -30 1350
rect -10 1230 5 1350
rect -45 1215 5 1230
rect 1055 1350 1105 1365
rect 1055 1230 1070 1350
rect 1090 1230 1105 1350
rect 1055 1215 1105 1230
rect 2155 1350 2205 1365
rect 2155 1230 2170 1350
rect 2190 1230 2205 1350
rect 2155 1215 2205 1230
rect -45 1000 5 1015
rect -45 730 -30 1000
rect -10 730 5 1000
rect -45 715 5 730
rect 1055 1000 1105 1015
rect 1055 730 1070 1000
rect 1090 730 1105 1000
rect 1055 715 1105 730
rect 2155 1000 2205 1015
rect 2155 730 2170 1000
rect 2190 730 2205 1000
rect 2155 715 2205 730
<< psubdiffcont >>
rect -30 205 -10 475
rect 1070 205 1090 475
rect 2170 205 2190 475
<< nsubdiffcont >>
rect -30 1230 -10 1350
rect 1070 1230 1090 1350
rect 2170 1230 2190 1350
rect -30 730 -10 1000
rect 1070 730 1090 1000
rect 2170 730 2190 1000
<< poly >>
rect 155 1410 205 1425
rect 155 1390 170 1410
rect 190 1390 205 1410
rect 55 1365 105 1380
rect 155 1365 205 1390
rect 255 1410 305 1425
rect 255 1390 270 1410
rect 290 1390 305 1410
rect 255 1365 305 1390
rect 355 1410 405 1425
rect 355 1390 370 1410
rect 390 1390 405 1410
rect 355 1365 405 1390
rect 455 1410 505 1425
rect 455 1390 470 1410
rect 490 1390 505 1410
rect 455 1365 505 1390
rect 555 1410 605 1425
rect 555 1390 570 1410
rect 590 1390 605 1410
rect 555 1365 605 1390
rect 655 1410 705 1425
rect 655 1390 670 1410
rect 690 1390 705 1410
rect 655 1365 705 1390
rect 755 1410 805 1425
rect 755 1390 770 1410
rect 790 1390 805 1410
rect 755 1365 805 1390
rect 855 1410 905 1425
rect 855 1390 870 1410
rect 890 1390 905 1410
rect 855 1365 905 1390
rect 1255 1410 1305 1425
rect 1255 1390 1270 1410
rect 1290 1390 1305 1410
rect 955 1365 1005 1380
rect 1155 1365 1205 1380
rect 1255 1365 1305 1390
rect 1355 1410 1405 1425
rect 1355 1390 1370 1410
rect 1390 1390 1405 1410
rect 1355 1365 1405 1390
rect 1455 1410 1505 1425
rect 1455 1390 1470 1410
rect 1490 1390 1505 1410
rect 1455 1365 1505 1390
rect 1555 1410 1605 1425
rect 1555 1390 1570 1410
rect 1590 1390 1605 1410
rect 1555 1365 1605 1390
rect 1655 1410 1705 1425
rect 1655 1390 1670 1410
rect 1690 1390 1705 1410
rect 1655 1365 1705 1390
rect 1755 1410 1805 1425
rect 1755 1390 1770 1410
rect 1790 1390 1805 1410
rect 1755 1365 1805 1390
rect 1855 1410 1905 1425
rect 1855 1390 1870 1410
rect 1890 1390 1905 1410
rect 1855 1365 1905 1390
rect 1955 1410 2005 1425
rect 1955 1390 1970 1410
rect 1990 1390 2005 1410
rect 1955 1365 2005 1390
rect 2055 1365 2105 1380
rect 55 1205 105 1215
rect 10 1190 105 1205
rect 155 1200 205 1215
rect 255 1200 305 1215
rect 355 1200 405 1215
rect 455 1200 505 1215
rect 555 1200 605 1215
rect 655 1200 705 1215
rect 755 1200 805 1215
rect 855 1200 905 1215
rect 955 1205 1005 1215
rect 1155 1205 1205 1215
rect 955 1190 1205 1205
rect 1255 1200 1305 1215
rect 1355 1200 1405 1215
rect 1455 1200 1505 1215
rect 1555 1200 1605 1215
rect 1655 1200 1705 1215
rect 1755 1200 1805 1215
rect 1855 1200 1905 1215
rect 1955 1200 2005 1215
rect 2055 1205 2105 1215
rect 2055 1190 2150 1205
rect 10 1170 20 1190
rect 40 1170 50 1190
rect 10 1160 50 1170
rect 1060 1170 1070 1190
rect 1090 1170 1100 1190
rect 1060 1160 1100 1170
rect 2110 1170 2120 1190
rect 2140 1170 2150 1190
rect 2110 1160 2150 1170
rect -65 1100 170 1110
rect -65 1080 -55 1100
rect -35 1095 170 1100
rect -35 1080 -25 1095
rect -65 1070 -25 1080
rect 155 1070 170 1095
rect 10 1060 50 1070
rect 10 1040 20 1060
rect 40 1040 50 1060
rect 155 1055 905 1070
rect 10 1025 105 1040
rect 55 1015 105 1025
rect 155 1015 205 1055
rect 255 1015 305 1030
rect 355 1015 405 1030
rect 455 1015 505 1055
rect 555 1015 605 1055
rect 655 1015 705 1030
rect 755 1015 805 1030
rect 855 1015 905 1055
rect 1060 1060 1100 1070
rect 1060 1040 1070 1060
rect 1090 1040 1100 1060
rect 1255 1060 1305 1075
rect 1255 1040 1270 1060
rect 1290 1040 1305 1060
rect 955 1025 1205 1040
rect 955 1015 1005 1025
rect 1155 1015 1205 1025
rect 1255 1015 1305 1040
rect 1355 1060 1405 1075
rect 1355 1040 1370 1060
rect 1390 1040 1405 1060
rect 1355 1015 1405 1040
rect 1455 1060 1505 1075
rect 1455 1040 1470 1060
rect 1490 1040 1505 1060
rect 1455 1015 1505 1040
rect 1555 1060 1605 1075
rect 1555 1040 1570 1060
rect 1590 1040 1605 1060
rect 1555 1015 1605 1040
rect 1655 1060 1705 1075
rect 1655 1040 1670 1060
rect 1690 1040 1705 1060
rect 1655 1015 1705 1040
rect 1755 1060 1805 1075
rect 1755 1040 1770 1060
rect 1790 1040 1805 1060
rect 1755 1015 1805 1040
rect 1855 1060 1905 1075
rect 1855 1040 1870 1060
rect 1890 1040 1905 1060
rect 1855 1015 1905 1040
rect 1955 1060 2005 1075
rect 1955 1040 1970 1060
rect 1990 1040 2005 1060
rect 2110 1060 2150 1070
rect 2110 1040 2120 1060
rect 2140 1040 2150 1060
rect 1955 1015 2005 1040
rect 2055 1025 2150 1040
rect 2055 1015 2105 1025
rect 55 700 105 715
rect 155 700 205 715
rect 255 675 305 715
rect 355 675 405 715
rect 455 700 505 715
rect 555 700 605 715
rect 655 675 705 715
rect 755 675 805 715
rect 855 700 905 715
rect 955 700 1005 715
rect 1155 700 1205 715
rect 1255 700 1305 715
rect 1355 700 1405 715
rect 1455 700 1505 715
rect 1555 700 1605 715
rect 1655 700 1705 715
rect 1755 700 1805 715
rect 1855 700 1905 715
rect 1955 700 2005 715
rect 2055 700 2105 715
rect -65 665 805 675
rect -65 645 -55 665
rect -35 660 805 665
rect -35 645 -25 660
rect -65 635 -25 645
rect 55 490 105 505
rect 155 490 205 505
rect 255 490 305 505
rect 355 490 405 505
rect 455 490 505 505
rect 555 490 605 505
rect 655 490 705 505
rect 755 490 805 505
rect 855 490 905 505
rect 955 490 1005 505
rect 1155 490 1205 505
rect 1255 490 1305 505
rect 1355 490 1405 505
rect 1455 490 1505 505
rect 1555 490 1605 505
rect 1655 490 1705 505
rect 1755 490 1805 505
rect 1855 490 1905 505
rect 1955 490 2005 505
rect 2055 490 2105 505
rect 55 180 105 190
rect 10 165 105 180
rect 155 165 205 190
rect 10 145 20 165
rect 40 145 50 165
rect 10 135 50 145
rect 155 145 170 165
rect 190 145 205 165
rect 155 130 205 145
rect 255 165 305 190
rect 255 145 270 165
rect 290 145 305 165
rect 255 130 305 145
rect 355 165 405 190
rect 355 145 370 165
rect 390 145 405 165
rect 355 130 405 145
rect 455 165 505 190
rect 455 145 470 165
rect 490 145 505 165
rect 455 130 505 145
rect 555 165 605 190
rect 555 145 570 165
rect 590 145 605 165
rect 555 130 605 145
rect 655 165 705 190
rect 655 145 670 165
rect 690 145 705 165
rect 655 130 705 145
rect 755 165 805 190
rect 755 145 770 165
rect 790 145 805 165
rect 755 130 805 145
rect 855 165 905 190
rect 955 180 1005 190
rect 1155 180 1205 190
rect 955 165 1205 180
rect 1255 165 1305 190
rect 855 145 870 165
rect 890 145 905 165
rect 855 130 905 145
rect 1060 145 1070 165
rect 1090 145 1100 165
rect 1060 135 1100 145
rect 1255 145 1270 165
rect 1290 145 1305 165
rect 1255 130 1305 145
rect 1355 165 1405 190
rect 1355 145 1370 165
rect 1390 145 1405 165
rect 1355 130 1405 145
rect 1455 165 1505 190
rect 1455 145 1470 165
rect 1490 145 1505 165
rect 1455 130 1505 145
rect 1555 165 1605 190
rect 1555 145 1570 165
rect 1590 145 1605 165
rect 1555 130 1605 145
rect 1655 165 1705 190
rect 1655 145 1670 165
rect 1690 145 1705 165
rect 1655 130 1705 145
rect 1755 165 1805 190
rect 1755 145 1770 165
rect 1790 145 1805 165
rect 1755 130 1805 145
rect 1855 165 1905 190
rect 1855 145 1870 165
rect 1890 145 1905 165
rect 1855 130 1905 145
rect 1955 165 2005 190
rect 2055 180 2105 190
rect 2055 165 2150 180
rect 1955 145 1970 165
rect 1990 145 2005 165
rect 1955 130 2005 145
rect 2110 145 2120 165
rect 2140 145 2150 165
rect 2110 135 2150 145
<< polycont >>
rect 170 1390 190 1410
rect 270 1390 290 1410
rect 370 1390 390 1410
rect 470 1390 490 1410
rect 570 1390 590 1410
rect 670 1390 690 1410
rect 770 1390 790 1410
rect 870 1390 890 1410
rect 1270 1390 1290 1410
rect 1370 1390 1390 1410
rect 1470 1390 1490 1410
rect 1570 1390 1590 1410
rect 1670 1390 1690 1410
rect 1770 1390 1790 1410
rect 1870 1390 1890 1410
rect 1970 1390 1990 1410
rect 20 1170 40 1190
rect 1070 1170 1090 1190
rect 2120 1170 2140 1190
rect -55 1080 -35 1100
rect 20 1040 40 1060
rect 1070 1040 1090 1060
rect 1270 1040 1290 1060
rect 1370 1040 1390 1060
rect 1470 1040 1490 1060
rect 1570 1040 1590 1060
rect 1670 1040 1690 1060
rect 1770 1040 1790 1060
rect 1870 1040 1890 1060
rect 1970 1040 1990 1060
rect 2120 1040 2140 1060
rect -55 645 -35 665
rect 20 145 40 165
rect 170 145 190 165
rect 270 145 290 165
rect 370 145 390 165
rect 470 145 490 165
rect 570 145 590 165
rect 670 145 690 165
rect 770 145 790 165
rect 870 145 890 165
rect 1070 145 1090 165
rect 1270 145 1290 165
rect 1370 145 1390 165
rect 1470 145 1490 165
rect 1570 145 1590 165
rect 1670 145 1690 165
rect 1770 145 1790 165
rect 1870 145 1890 165
rect 1970 145 1990 165
rect 2120 145 2140 165
<< locali >>
rect -65 1410 2050 1420
rect -65 1390 170 1410
rect 190 1390 270 1410
rect 290 1390 370 1410
rect 390 1390 470 1410
rect 490 1390 570 1410
rect 590 1390 670 1410
rect 690 1390 770 1410
rect 790 1390 870 1410
rect 890 1390 1270 1410
rect 1290 1390 1370 1410
rect 1390 1390 1470 1410
rect 1490 1390 1570 1410
rect 1590 1390 1670 1410
rect 1690 1390 1770 1410
rect 1790 1390 1870 1410
rect 1890 1390 1970 1410
rect 1990 1390 2050 1410
rect -65 1380 2050 1390
rect -40 1350 50 1360
rect -40 1230 -30 1350
rect -10 1230 20 1350
rect 40 1230 50 1350
rect -40 1220 50 1230
rect 110 1350 150 1380
rect 110 1230 120 1350
rect 140 1230 150 1350
rect 110 1220 150 1230
rect 210 1350 250 1360
rect 210 1230 220 1350
rect 240 1230 250 1350
rect 210 1220 250 1230
rect 310 1350 350 1360
rect 310 1230 320 1350
rect 340 1230 350 1350
rect 10 1190 50 1220
rect 10 1170 20 1190
rect 40 1170 50 1190
rect 10 1160 50 1170
rect 310 1135 350 1230
rect 410 1350 450 1360
rect 410 1230 420 1350
rect 440 1230 450 1350
rect 410 1220 450 1230
rect 510 1350 550 1380
rect 510 1230 520 1350
rect 540 1230 550 1350
rect 510 1220 550 1230
rect 610 1350 650 1360
rect 610 1230 620 1350
rect 640 1230 650 1350
rect 610 1220 650 1230
rect 710 1350 750 1360
rect 710 1230 720 1350
rect 740 1230 750 1350
rect 710 1135 750 1230
rect 810 1350 850 1360
rect 810 1230 820 1350
rect 840 1230 850 1350
rect 810 1220 850 1230
rect 910 1350 950 1380
rect 910 1230 920 1350
rect 940 1230 950 1350
rect 910 1220 950 1230
rect 1010 1350 1150 1360
rect 1010 1230 1020 1350
rect 1040 1230 1070 1350
rect 1090 1230 1120 1350
rect 1140 1230 1150 1350
rect 1010 1220 1150 1230
rect 1210 1350 1250 1380
rect 1210 1230 1220 1350
rect 1240 1230 1250 1350
rect 1210 1220 1250 1230
rect 1310 1350 1350 1360
rect 1310 1230 1320 1350
rect 1340 1230 1350 1350
rect 1310 1220 1350 1230
rect 1410 1350 1450 1360
rect 1410 1230 1420 1350
rect 1440 1230 1450 1350
rect 1060 1190 1100 1220
rect 1060 1170 1070 1190
rect 1090 1170 1100 1190
rect 1060 1160 1100 1170
rect 1410 1135 1450 1230
rect 1510 1350 1550 1360
rect 1510 1230 1520 1350
rect 1540 1230 1550 1350
rect 1510 1220 1550 1230
rect 1610 1350 1650 1380
rect 1610 1230 1620 1350
rect 1640 1230 1650 1350
rect 1610 1220 1650 1230
rect 1710 1350 1750 1360
rect 1710 1230 1720 1350
rect 1740 1230 1750 1350
rect 1710 1220 1750 1230
rect 1810 1350 1850 1360
rect 1810 1230 1820 1350
rect 1840 1230 1850 1350
rect 1810 1135 1850 1230
rect 1910 1350 1950 1360
rect 1910 1230 1920 1350
rect 1940 1230 1950 1350
rect 1910 1220 1950 1230
rect 2010 1350 2050 1380
rect 2010 1230 2020 1350
rect 2040 1230 2050 1350
rect 2010 1220 2050 1230
rect 2110 1350 2200 1360
rect 2110 1230 2120 1350
rect 2140 1230 2170 1350
rect 2190 1230 2200 1350
rect 2110 1220 2200 1230
rect 2110 1190 2150 1220
rect 2110 1170 2120 1190
rect 2140 1170 2150 1190
rect 2110 1160 2150 1170
rect -65 1100 -25 1110
rect -65 1080 -55 1100
rect -35 1080 -25 1100
rect -65 1070 -25 1080
rect 210 1095 1850 1135
rect 10 1060 50 1070
rect 10 1040 20 1060
rect 40 1040 50 1060
rect 10 1010 50 1040
rect -40 1000 50 1010
rect -40 730 -30 1000
rect -10 730 20 1000
rect 40 730 50 1000
rect -40 720 50 730
rect 110 1000 150 1010
rect 110 730 120 1000
rect 140 730 150 1000
rect -65 665 -25 675
rect -65 645 -55 665
rect -35 645 -25 665
rect -65 635 -25 645
rect 110 620 150 730
rect 210 1000 250 1095
rect 210 730 220 1000
rect 240 730 250 1000
rect 210 720 250 730
rect 310 1000 350 1010
rect 310 730 320 1000
rect 340 730 350 1000
rect 310 690 350 730
rect 410 1000 450 1095
rect 410 730 420 1000
rect 440 730 450 1000
rect 410 720 450 730
rect 510 1000 550 1010
rect 510 730 520 1000
rect 540 730 550 1000
rect 310 680 390 690
rect 310 660 320 680
rect 380 660 390 680
rect 310 650 390 660
rect 510 620 550 730
rect 610 1000 650 1095
rect 610 730 620 1000
rect 640 730 650 1000
rect 610 720 650 730
rect 710 1000 750 1010
rect 710 730 720 1000
rect 740 730 750 1000
rect 710 690 750 730
rect 810 1000 850 1095
rect 1060 1060 1100 1070
rect 1060 1040 1070 1060
rect 1090 1040 1100 1060
rect 1060 1010 1100 1040
rect 1210 1060 2050 1070
rect 1210 1040 1270 1060
rect 1290 1040 1370 1060
rect 1390 1040 1470 1060
rect 1490 1040 1570 1060
rect 1590 1040 1670 1060
rect 1690 1040 1770 1060
rect 1790 1040 1870 1060
rect 1890 1040 1970 1060
rect 1990 1040 2050 1060
rect 1210 1030 2050 1040
rect 810 730 820 1000
rect 840 730 850 1000
rect 810 720 850 730
rect 910 1000 950 1010
rect 910 730 920 1000
rect 940 730 950 1000
rect 670 680 750 690
rect 670 660 680 680
rect 740 660 750 680
rect 670 650 750 660
rect 910 620 950 730
rect 1010 1000 1150 1010
rect 1010 730 1020 1000
rect 1040 730 1070 1000
rect 1090 730 1120 1000
rect 1140 730 1150 1000
rect 1010 720 1150 730
rect 1210 1000 1250 1030
rect 1210 730 1220 1000
rect 1240 730 1250 1000
rect 1210 690 1250 730
rect 1310 1000 1350 1010
rect 1310 730 1320 1000
rect 1340 730 1350 1000
rect 1310 720 1350 730
rect 1410 1000 1450 1010
rect 1410 730 1420 1000
rect 1440 730 1450 1000
rect 1170 680 1250 690
rect 1170 660 1180 680
rect 1240 660 1250 680
rect 1170 650 1250 660
rect 1410 620 1450 730
rect 1510 1000 1550 1010
rect 1510 730 1520 1000
rect 1540 730 1550 1000
rect 1510 720 1550 730
rect 1610 1000 1650 1030
rect 1610 730 1620 1000
rect 1640 730 1650 1000
rect 1610 720 1650 730
rect 1710 1000 1750 1010
rect 1710 730 1720 1000
rect 1740 730 1750 1000
rect 1710 720 1750 730
rect 1810 1000 1850 1010
rect 1810 730 1820 1000
rect 1840 730 1850 1000
rect 1810 620 1850 730
rect 1910 1000 1950 1010
rect 1910 730 1920 1000
rect 1940 730 1950 1000
rect 1910 720 1950 730
rect 2010 1000 2050 1030
rect 2010 730 2020 1000
rect 2040 730 2050 1000
rect 2010 720 2050 730
rect 2110 1060 2150 1070
rect 2110 1040 2120 1060
rect 2140 1040 2150 1060
rect 2110 1010 2150 1040
rect 2110 1000 2200 1010
rect 2110 730 2120 1000
rect 2140 730 2170 1000
rect 2190 730 2200 1000
rect 2110 720 2200 730
rect 110 580 1250 620
rect 110 550 190 560
rect 110 530 120 550
rect 180 530 190 550
rect 110 520 190 530
rect 310 550 390 560
rect 310 530 320 550
rect 380 530 390 550
rect 310 520 390 530
rect 670 550 750 560
rect 670 530 680 550
rect 740 530 750 550
rect 670 520 750 530
rect -40 475 50 485
rect -40 205 -30 475
rect -10 205 20 475
rect 40 205 50 475
rect -40 195 50 205
rect 10 165 50 195
rect 10 145 20 165
rect 40 145 50 165
rect 10 135 50 145
rect 110 475 150 520
rect 110 205 120 475
rect 140 205 150 475
rect 110 175 150 205
rect 210 475 250 485
rect 210 205 220 475
rect 240 205 250 475
rect 210 195 250 205
rect 310 475 350 520
rect 310 205 320 475
rect 340 205 350 475
rect 310 195 350 205
rect 410 475 450 485
rect 410 205 420 475
rect 440 205 450 475
rect 410 195 450 205
rect 510 475 550 485
rect 510 205 520 475
rect 540 205 550 475
rect 510 175 550 205
rect 610 475 650 485
rect 610 205 620 475
rect 640 205 650 475
rect 610 195 650 205
rect 710 475 750 520
rect 710 205 720 475
rect 740 205 750 475
rect 710 195 750 205
rect 810 475 850 485
rect 810 205 820 475
rect 840 205 850 475
rect 810 195 850 205
rect 910 475 950 485
rect 910 205 920 475
rect 940 205 950 475
rect 910 175 950 205
rect 1010 475 1150 485
rect 1010 205 1020 475
rect 1040 205 1070 475
rect 1090 205 1120 475
rect 1140 205 1150 475
rect 1010 195 1150 205
rect 1210 475 1250 580
rect 1410 580 2220 620
rect 1210 205 1220 475
rect 1240 205 1250 475
rect 110 165 950 175
rect 110 145 170 165
rect 190 145 270 165
rect 290 145 370 165
rect 390 145 470 165
rect 490 145 570 165
rect 590 145 670 165
rect 690 145 770 165
rect 790 145 870 165
rect 890 145 950 165
rect 110 135 950 145
rect 1060 165 1100 195
rect 1060 145 1070 165
rect 1090 145 1100 165
rect 1060 135 1100 145
rect 1210 175 1250 205
rect 1310 475 1350 485
rect 1310 205 1320 475
rect 1340 205 1350 475
rect 1310 195 1350 205
rect 1410 475 1450 580
rect 1410 205 1420 475
rect 1440 205 1450 475
rect 1410 195 1450 205
rect 1510 475 1550 485
rect 1510 205 1520 475
rect 1540 205 1550 475
rect 1510 195 1550 205
rect 1610 475 1650 485
rect 1610 205 1620 475
rect 1640 205 1650 475
rect 1610 175 1650 205
rect 1710 475 1750 485
rect 1710 205 1720 475
rect 1740 205 1750 475
rect 1710 195 1750 205
rect 1810 475 1850 580
rect 1810 205 1820 475
rect 1840 205 1850 475
rect 1810 195 1850 205
rect 1910 475 1950 485
rect 1910 205 1920 475
rect 1940 205 1950 475
rect 1910 195 1950 205
rect 2010 475 2050 485
rect 2010 205 2020 475
rect 2040 205 2050 475
rect 2010 175 2050 205
rect 1210 165 2050 175
rect 1210 145 1270 165
rect 1290 145 1370 165
rect 1390 145 1470 165
rect 1490 145 1570 165
rect 1590 145 1670 165
rect 1690 145 1770 165
rect 1790 145 1870 165
rect 1890 145 1970 165
rect 1990 145 2050 165
rect 1210 135 2050 145
rect 2110 475 2200 485
rect 2110 205 2120 475
rect 2140 205 2170 475
rect 2190 205 2200 475
rect 2110 195 2200 205
rect 2110 165 2150 195
rect 2110 145 2120 165
rect 2140 145 2150 165
rect 2110 135 2150 145
<< viali >>
rect -30 1230 -10 1350
rect 20 1230 40 1350
rect 220 1230 240 1350
rect 420 1230 440 1350
rect 620 1230 640 1350
rect 820 1230 840 1350
rect 1020 1230 1040 1350
rect 1070 1230 1090 1350
rect 1120 1230 1140 1350
rect 1320 1230 1340 1350
rect 1520 1230 1540 1350
rect 1720 1230 1740 1350
rect 1920 1230 1940 1350
rect 2120 1230 2140 1350
rect 2170 1230 2190 1350
rect -30 730 -10 1000
rect 20 730 40 1000
rect 320 660 380 680
rect 680 660 740 680
rect 1020 730 1040 1000
rect 1070 730 1090 1000
rect 1120 730 1140 1000
rect 1320 730 1340 1000
rect 1180 660 1240 680
rect 1520 730 1540 1000
rect 1720 730 1740 1000
rect 1920 730 1940 1000
rect 2120 730 2140 1000
rect 2170 730 2190 1000
rect 120 530 180 550
rect 320 530 380 550
rect 680 530 740 550
rect -30 205 -10 475
rect 20 205 40 475
rect 220 205 240 475
rect 420 205 440 475
rect 620 205 640 475
rect 820 205 840 475
rect 1020 205 1040 475
rect 1070 205 1090 475
rect 1120 205 1140 475
rect 1320 205 1340 475
rect 1520 205 1540 475
rect 1720 205 1740 475
rect 1920 205 1940 475
rect 2120 205 2140 475
rect 2170 205 2190 475
<< metal1 >>
rect -65 1350 2225 1360
rect -65 1230 -30 1350
rect -10 1230 20 1350
rect 40 1230 220 1350
rect 240 1230 420 1350
rect 440 1230 620 1350
rect 640 1230 820 1350
rect 840 1230 1020 1350
rect 1040 1230 1070 1350
rect 1090 1230 1120 1350
rect 1140 1230 1320 1350
rect 1340 1230 1520 1350
rect 1540 1230 1720 1350
rect 1740 1230 1920 1350
rect 1940 1230 2120 1350
rect 2140 1230 2170 1350
rect 2190 1230 2225 1350
rect -65 1000 2225 1230
rect -65 730 -30 1000
rect -10 730 20 1000
rect 40 730 1020 1000
rect 1040 730 1070 1000
rect 1090 730 1120 1000
rect 1140 730 1320 1000
rect 1340 730 1520 1000
rect 1540 730 1720 1000
rect 1740 730 1920 1000
rect 1940 730 2120 1000
rect 2140 730 2170 1000
rect 2190 730 2225 1000
rect -65 720 2225 730
rect 210 680 750 690
rect 210 660 320 680
rect 380 660 680 680
rect 740 660 750 680
rect 210 650 750 660
rect 1060 680 1250 690
rect 1060 660 1180 680
rect 1240 660 1250 680
rect 1060 650 1250 660
rect 210 560 250 650
rect 1060 560 1100 650
rect 110 550 250 560
rect 110 530 120 550
rect 180 530 250 550
rect 110 520 250 530
rect 310 550 1100 560
rect 310 530 320 550
rect 380 530 680 550
rect 740 530 1100 550
rect 310 520 1100 530
rect -65 475 2225 485
rect -65 205 -30 475
rect -10 205 20 475
rect 40 205 220 475
rect 240 205 420 475
rect 440 205 620 475
rect 640 205 820 475
rect 840 205 1020 475
rect 1040 205 1070 475
rect 1090 205 1120 475
rect 1140 205 1320 475
rect 1340 205 1520 475
rect 1540 205 1720 475
rect 1740 205 1920 475
rect 1940 205 2120 475
rect 2140 205 2170 475
rect 2190 205 2225 475
rect -65 195 2225 205
<< labels >>
flabel locali 2220 600 2220 600 3 FreeSans 80 0 40 0 Vout
port 3 e
flabel locali -65 1400 -65 1400 7 FreeSans 80 0 -40 0 Vb
port 4 w
flabel locali -65 1090 -65 1090 7 FreeSans 80 0 -40 0 V1
port 1 w
flabel locali -65 655 -65 655 7 FreeSans 80 0 -40 0 V2
port 2 w
flabel metal1 -65 340 -65 340 7 FreeSans 80 0 -40 0 VN
port 6 w
flabel metal1 -65 1020 -65 1020 7 FreeSans 80 0 -80 0 VP
port 5 w
<< end >>
