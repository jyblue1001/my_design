* SPICE3 file created from mimcap_1pF.ext - technology: sky130A

X0 top bot sky130_fd_pr__cap_mim_m3_1 l=20 w=25
C0 bot VSUBS 10.1352f **FLOATING
