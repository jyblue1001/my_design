** sch_path: /foss/designs/my_design/projects/pll/charge_pump/xschem_ngspice/loop_filter_xschem.sch
**.subckt loop_filter_xschem VOUT GNDA
*.ipin GNDA
*.iopin VOUT
XC2 GNDA VOUT sky130_fd_pr__cap_mim_m3_1 W=13.8 L=60 MF=1 m=1
XC1 GNDA R1_C1 sky130_fd_pr__cap_mim_m3_1 W=69.8 L=60 MF=1 m=1
XR1 R1_C1 VOUT GNDA sky130_fd_pr__res_xhigh_po_0p35 L=7.52 mult=1 m=1
**.ends
.end
