* PEX produced on Thu Aug  7 12:18:39 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from two_stage_opamp_dummy_magic_24.ext - technology: sky130A

.subckt two_stage_opamp_dummy_magic_24 V_CMFB_S1 V_CMFB_S3 Vb3 Vb2 V_CMFB_S2 V_CMFB_S4
+ VOUT- VOUT+ V_tail_gate V_err_amp_ref V_err_gate
X0 VOUT-.t15 X.t25 w_109060_7290.t106 w_109060_7290.t105 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1 VOUT-.t1 V_b_2nd_stage.t2 a_109160_2280.t125 a_109160_2280.t124 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X2 VOUT+.t19 cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VOUT+.t20 cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 w_109060_7290.t104 X.t26 V_CMFB_S2.t10 a_109160_2280.t109 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X5 VOUT-.t19 cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT-.t20 cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VOUT-.t21 cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 w_109060_7290.t28 Vb3.t2 VD4.t25 w_109060_7290.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X9 V_source.t19 V_tail_gate.t4 a_109160_2280.t26 a_109160_2280.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X10 VD1.t18 VIN- V_source.t30 a_109160_2280.t206 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X11 VOUT+.t21 cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VOUT-.t22 cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 a_109160_2280.t228 V_tail_gate.t5 V_source.t18 a_109160_2280.t227 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X14 VD3.t35 Vb2.t3 X.t6 VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X15 VOUT-.t2 V_b_2nd_stage.t3 a_109160_2280.t123 a_109160_2280.t122 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X16 V_err_mir_p.t2 V_err_amp_ref.t0 V_err_gate.t0 w_109060_7290.t32 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X17 err_amp_mir.t3 w_109060_7290.t176 w_109060_7290.t178 w_109060_7290.t177 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X18 VOUT+.t22 cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VOUT+.t23 cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VOUT+.t24 cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT+.t25 cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 a_109160_2280.t196 a_109160_2280.t193 a_109160_2280.t195 a_109160_2280.t194 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X23 VOUT+.t26 cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 VOUT+.t27 cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VOUT-.t23 cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 VOUT+.t13 w_109060_7290.t173 w_109060_7290.t175 w_109060_7290.t174 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X27 VOUT-.t24 cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VOUT+.t28 cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VOUT-.t25 cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 a_109160_2280.t192 a_109160_2280.t190 VD2.t9 a_109160_2280.t191 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X31 VOUT-.t26 cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VOUT+.t29 cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 V_source.t17 V_tail_gate.t6 a_109160_2280.t2 a_109160_2280.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X34 VOUT+.t30 cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 w_109060_7290.t172 w_109060_7290.t170 VOUT+.t12 w_109060_7290.t171 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X36 VOUT-.t27 cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 Y.t18 Vb2.t4 VD4.t13 VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X38 V_CMFB_S3.t10 Y.t25 a_109160_2280.t81 w_109060_7290.t62 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X39 VD1.t21 Vb1.t10 X.t24 a_109160_2280.t232 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X40 VOUT+.t31 cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 a_109160_2280.t67 V_tail_gate.t7 V_source.t16 a_109160_2280.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X42 VOUT+.t32 cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VOUT+.t33 cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT+.t34 cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 VOUT+.t35 cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 X.t8 Vb2.t5 VD3.t33 VD3.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X47 VOUT-.t28 cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT+.t36 cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VOUT-.t29 cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 a_109160_2280.t108 X.t27 V_CMFB_S1.t10 w_109060_7290.t103 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X51 VOUT-.t30 cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VOUT-.t31 cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 w_109060_7290.t102 X.t28 V_CMFB_S2.t9 a_109160_2280.t107 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X54 Y.t17 Vb2.t6 VD4.t7 VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X55 Y.t2 Vb1.t11 VD2.t2 a_109160_2280.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X56 VOUT+.t37 cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VD4.t24 Vb3.t3 w_109060_7290.t53 w_109060_7290.t52 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X58 VOUT+.t38 cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VD1.t8 a_109160_2280.t187 a_109160_2280.t189 a_109160_2280.t188 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X60 VOUT+.t39 cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT+.t40 cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT+.t41 cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 VOUT+.t42 cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 VOUT-.t32 cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 VOUT-.t33 cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VOUT-.t34 cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VOUT-.t35 cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT-.t36 cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 VOUT-.t37 cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VOUT+.t43 cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VOUT-.t38 cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 V_CMFB_S2.t8 X.t29 w_109060_7290.t95 a_109160_2280.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X73 VOUT+.t44 cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 V_tail_gate.t2 VIN- V_p_mir.t2 a_109160_2280.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X75 V_source.t38 VIN+ VD2.t19 a_109160_2280.t220 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X76 VOUT-.t39 cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 w_109060_7290.t190 Y.t26 VOUT+.t16 w_109060_7290.t189 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X78 VOUT+.t45 cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VOUT+.t46 cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VD3.t15 Vb3.t4 w_109060_7290.t1 w_109060_7290.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X81 X.t0 Vb2.t7 VD3.t31 VD3.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X82 VOUT-.t40 cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VOUT+.t47 cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT+.t48 cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT-.t41 cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 a_109160_2280.t186 a_109160_2280.t184 Vb1.t9 a_109160_2280.t185 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X87 VOUT-.t42 cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT-.t43 cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VOUT-.t14 X.t30 w_109060_7290.t101 w_109060_7290.t100 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X90 VOUT+.t49 cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VOUT+.t50 cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 a_109160_2280.t105 X.t31 V_CMFB_S1.t9 w_109060_7290.t99 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X93 VOUT+.t51 cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VD4.t23 Vb3.t5 w_109060_7290.t108 w_109060_7290.t107 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X95 VOUT-.t44 cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT-.t45 cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT+.t52 cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 V_CMFB_S4.t10 Y.t27 w_109060_7290.t35 a_109160_2280.t38 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X99 w_109060_7290.t200 a_109160_2280.t181 a_109160_2280.t183 a_109160_2280.t182 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X100 Y.t23 Vb1.t12 VD2.t20 a_109160_2280.t226 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X101 VOUT-.t46 cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VOUT-.t47 cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 X.t17 Vb2.t8 VD3.t29 VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X104 VOUT-.t48 cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT-.t49 cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VOUT-.t50 cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 err_amp_out.t0 V_err_amp_ref.t1 V_err_p.t2 w_109060_7290.t36 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X108 VOUT-.t51 cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 V_CMFB_S1.t8 X.t32 a_109160_2280.t104 w_109060_7290.t98 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X110 VOUT+.t53 cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT+.t9 V_b_2nd_stage.t4 a_109160_2280.t121 a_109160_2280.t120 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X112 VD4.t5 Vb2.t9 Y.t16 VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X113 V_source.t35 VIN+ VD2.t18 a_109160_2280.t219 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X114 VOUT-.t52 cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 V_tail_gate.t1 a_109160_2280.t179 a_109160_2280.t180 a_109160_2280.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X116 a_118660_3088.t1 V_tot.t2 a_109160_2280.t73 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X117 VOUT-.t53 cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 a_109160_2280.t178 a_109160_2280.t176 VD1.t7 a_109160_2280.t177 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X119 VOUT+.t54 cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT+.t55 cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 Vb1_2.t3 Vb1.t0 Vb1.t1 a_109160_2280.t89 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X122 VOUT-.t13 X.t33 w_109060_7290.t97 w_109060_7290.t96 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X123 Vb2_Vb3.t6 Vb2_Vb3.t3 Vb2_Vb3.t5 Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X124 V_CMFB_S3.t9 Y.t28 a_109160_2280.t47 w_109060_7290.t47 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X125 a_109160_2280.t210 w_109060_7290.t164 w_109060_7290.t166 w_109060_7290.t165 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X126 VD4.t3 Vb2.t10 Y.t15 VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X127 VOUT-.t54 cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 w_109060_7290.t169 w_109060_7290.t167 VD4.t33 w_109060_7290.t168 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X129 VOUT-.t55 cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT-.t56 cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VOUT+.t56 cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 V_CMFB_S4.t9 Y.t29 w_109060_7290.t30 a_109160_2280.t33 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X133 Y.t24 Vb1.t13 VD2.t21 a_109160_2280.t230 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X134 VOUT+.t57 cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 X.t23 Vb1.t14 VD1.t20 a_109160_2280.t231 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X136 VOUT-.t57 cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 V_source.t0 Vb1.t15 Vb1_2.t4 a_109160_2280.t43 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X138 VOUT-.t58 cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT+.t58 cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VOUT+.t59 cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 w_109060_7290.t16 V_err_gate.t4 V_err_p.t1 w_109060_7290.t15 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X142 a_109160_2280.t175 a_109160_2280.t173 err_amp_out.t2 a_109160_2280.t174 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X143 VOUT+.t60 cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT+.t61 cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 w_109060_7290.t94 X.t34 VOUT-.t12 w_109060_7290.t93 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X146 VOUT+.t62 cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 Vb2_Vb3.t10 w_109060_7290.t161 w_109060_7290.t163 w_109060_7290.t162 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X148 VOUT-.t59 cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT-.t60 cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VOUT+.t63 cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VOUT-.t61 cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 V_source.t33 VIN+ VD2.t17 a_109160_2280.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X153 VOUT+.t64 cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 a_109160_2280.t172 a_109160_2280.t170 w_109060_7290.t179 a_109160_2280.t171 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X155 VD3.t27 Vb2.t11 X.t2 VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X156 w_109060_7290.t112 Vb3.t6 VD3.t14 w_109060_7290.t111 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X157 VOUT-.t62 cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 V_source.t23 VIN- VD1.t17 a_109160_2280.t205 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X159 VOUT-.t63 cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 V_source.t27 VIN- VD1.t16 a_109160_2280.t204 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X161 Vb2_Vb3.t2 Vb2_Vb3.t0 Vb3.t0 Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X162 cap_res_Y.t0 Y.t6 a_109160_2280.t65 sky130_fd_pr__res_high_po_1p41 l=1.41
X163 VOUT+.t65 cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 Vb1_2.t2 Vb1.t4 Vb1.t5 a_109160_2280.t64 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X165 V_CMFB_S4.t8 Y.t30 w_109060_7290.t26 a_109160_2280.t31 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X166 VD4.t31 VD4.t29 Y.t22 VD4.t30 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X167 VOUT+.t66 cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT-.t64 cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT+.t67 cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT-.t65 cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 w_109060_7290.t114 Vb3.t7 VD4.t22 w_109060_7290.t113 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X172 V_b_2nd_stage.t1 a_108650_n784.t1 a_109160_2280.t85 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X173 VOUT-.t66 cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 w_109060_7290.t56 Y.t31 VOUT+.t5 w_109060_7290.t55 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X175 VOUT-.t17 w_109060_7290.t158 w_109060_7290.t160 w_109060_7290.t159 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X176 VOUT-.t67 cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 V_CMFB_S3.t8 Y.t32 a_109160_2280.t233 w_109060_7290.t197 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X178 w_109060_7290.t49 Vb3.t8 VD3.t13 w_109060_7290.t48 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X179 VOUT-.t68 cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VD3.t5 VD3.t3 X.t14 VD3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X181 Y.t3 Vb1.t16 VD2.t3 a_109160_2280.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X182 VOUT+.t68 cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 V_CMFB_S4.t7 Y.t33 w_109060_7290.t46 a_109160_2280.t46 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X184 X.t20 Vb1.t17 VD1.t19 a_109160_2280.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X185 X.t4 Vb1.t18 VD1.t1 a_109160_2280.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X186 VOUT+.t69 cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VOUT+.t70 cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VOUT+.t71 cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VOUT+.t72 cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 V_source.t15 V_tail_gate.t8 a_109160_2280.t53 a_109160_2280.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X191 VOUT-.t69 cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VOUT+.t73 cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 a_109160_2280.t62 err_amp_mir.t0 err_amp_mir.t1 a_109160_2280.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X194 VOUT-.t70 cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT-.t71 cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT-.t72 cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 V_source.t14 V_tail_gate.t9 a_109160_2280.t4 a_109160_2280.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X198 Y.t14 Vb2.t12 VD4.t9 VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X199 w_109060_7290.t157 w_109060_7290.t155 a_109160_2280.t209 w_109060_7290.t156 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X200 VOUT+.t74 cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VD2.t0 Vb1.t19 Y.t0 a_109160_2280.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X202 V_source.t31 VIN+ VD2.t16 a_109160_2280.t217 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X203 VOUT-.t73 cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT-.t74 cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 a_109160_2280.t19 V_tail_gate.t10 V_source.t13 a_109160_2280.t18 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X206 V_CMFB_S2.t7 X.t35 w_109060_7290.t68 a_109160_2280.t103 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X207 V_source.t28 VIN- VD1.t15 a_109160_2280.t203 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X208 VOUT+.t75 cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT+.t76 cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 V_CMFB_S3.t7 Y.t34 a_109160_2280.t36 w_109060_7290.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X211 VOUT+.t77 cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+.t78 cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT-.t75 cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 V_source.t1 err_amp_out.t4 a_109160_2280.t51 a_109160_2280.t50 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X215 V_err_gate.t3 V_tot.t4 V_err_mir_p.t3 w_109060_7290.t191 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X216 VOUT-.t76 cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VOUT-.t77 cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT+.t79 cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT-.t78 cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 Vb3.t1 Vb2.t13 Vb2_Vb3.t9 Vb2_Vb3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X221 w_109060_7290.t154 w_109060_7290.t152 VD3.t37 w_109060_7290.t153 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X222 VOUT+.t80 cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 Y.t13 Vb2.t14 VD4.t1 VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X224 w_109060_7290.t45 Y.t35 VOUT+.t4 w_109060_7290.t44 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X225 a_108510_3088.t1 V_tot.t1 a_109160_2280.t71 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X226 VOUT+.t81 cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t82 cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 V_CMFB_S3.t6 Y.t36 a_109160_2280.t28 w_109060_7290.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X229 VOUT-.t79 cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VD2.t15 VIN+ V_source.t34 a_109160_2280.t216 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 VOUT+.t83 cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VOUT+.t84 cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 Y.t20 a_109160_2280.t167 a_109160_2280.t169 a_109160_2280.t168 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X234 X.t3 Vb1.t20 VD1.t0 a_109160_2280.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X235 VOUT-.t80 cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT+.t85 cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VOUT-.t81 cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 Y.t12 Vb2.t15 VD4.t15 VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X239 VOUT+.t86 cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT-.t82 cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT-.t83 cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 w_109060_7290.t10 Y.t37 V_CMFB_S4.t6 a_109160_2280.t10 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X243 a_109160_2280.t119 V_b_2nd_stage.t5 VOUT+.t8 a_109160_2280.t118 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X244 w_109060_7290.t7 Vb3.t9 Vb2_Vb3.t7 w_109060_7290.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X245 VOUT+.t87 cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT-.t84 cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 a_109160_2280.t87 V_tail_gate.t11 V_source.t12 a_109160_2280.t86 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X248 w_109060_7290.t151 w_109060_7290.t149 VOUT-.t16 w_109060_7290.t150 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X249 VOUT-.t85 cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VOUT+.t88 cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VD3.t12 Vb3.t10 w_109060_7290.t64 w_109060_7290.t63 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 VOUT+.t89 cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VOUT+.t90 cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 V_CMFB_S1.t7 X.t36 a_109160_2280.t102 w_109060_7290.t92 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X255 X.t15 Vb2.t16 VD3.t25 VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X256 VOUT-.t86 cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 V_CMFB_S2.t6 X.t37 w_109060_7290.t69 a_109160_2280.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X258 V_source.t11 V_tail_gate.t12 a_109160_2280.t224 a_109160_2280.t223 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X259 w_109060_7290.t188 Y.t38 VOUT+.t15 w_109060_7290.t187 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X260 VOUT-.t87 cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 a_109160_2280.t117 V_b_2nd_stage.t6 VOUT+.t7 a_109160_2280.t116 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X262 V_source.t29 VIN- VD1.t14 a_109160_2280.t202 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X263 VOUT-.t88 cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VOUT+.t91 cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 V_p_mir.t1 V_tail_gate.t13 a_109160_2280.t40 a_109160_2280.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X266 VOUT-.t89 cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 a_109160_2280.t115 V_b_2nd_stage.t7 VOUT-.t18 a_109160_2280.t114 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X268 w_109060_7290.t3 V_err_gate.t5 V_err_mir_p.t1 w_109060_7290.t2 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X269 VOUT+.t0 a_108650_n784.t0 a_109160_2280.t24 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X270 VD4.t21 Vb3.t11 w_109060_7290.t58 w_109060_7290.t57 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X271 VOUT+.t92 cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 a_109160_2280.t78 V_tail_gate.t14 V_source.t10 a_109160_2280.t77 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X273 VOUT+.t93 cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 Vb2_2.t2 Vb2.t17 w_109060_7290.t184 w_109060_7290.t183 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X275 VD3.t11 Vb3.t12 w_109060_7290.t199 w_109060_7290.t198 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X276 w_109060_7290.t34 Y.t39 VOUT+.t2 w_109060_7290.t33 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X277 VOUT-.t90 cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VOUT-.t91 cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VOUT-.t92 cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VOUT+.t94 cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 V_source.t9 V_tail_gate.t15 a_109160_2280.t84 a_109160_2280.t83 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X282 VOUT+.t95 cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VOUT-.t93 cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 a_109160_2280.t113 V_b_2nd_stage.t8 VOUT-.t3 a_109160_2280.t112 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X285 a_109160_2280.t42 Y.t40 V_CMFB_S3.t5 w_109060_7290.t40 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X286 X.t5 Vb1.t21 VD1.t2 a_109160_2280.t29 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X287 Vb1.t8 a_109160_2280.t164 a_109160_2280.t166 a_109160_2280.t165 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X288 w_109060_7290.t43 Y.t41 V_CMFB_S4.t5 a_109160_2280.t45 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X289 VD3.t10 Vb3.t13 w_109060_7290.t116 w_109060_7290.t115 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X290 VOUT+.t96 cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT+.t97 cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VD4.t11 Vb2.t18 Y.t11 VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X293 VOUT+.t98 cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT-.t94 cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VOUT-.t95 cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VOUT+.t99 cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 w_109060_7290.t91 X.t38 VOUT-.t11 w_109060_7290.t90 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X298 V_CMFB_S1.t6 X.t39 a_109160_2280.t100 w_109060_7290.t89 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X299 VOUT-.t96 cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t97 cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT-.t98 cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 VOUT-.t99 cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 V_CMFB_S2.t5 X.t40 w_109060_7290.t81 a_109160_2280.t99 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X304 a_109160_2280.t163 a_109160_2280.t161 Y.t19 a_109160_2280.t162 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X305 VOUT-.t100 cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 V_source.t24 VIN- VD1.t13 a_109160_2280.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X307 VOUT-.t101 cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 V_err_gate.t2 w_109060_7290.t146 w_109060_7290.t148 w_109060_7290.t147 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X309 VOUT-.t102 cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VOUT-.t103 cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 a_108630_3088.t0 V_tot.t0 a_109160_2280.t14 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X312 VOUT-.t104 cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VOUT-.t105 cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 w_109060_7290.t82 X.t41 V_CMFB_S2.t4 a_109160_2280.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X315 w_109060_7290.t145 w_109060_7290.t142 w_109060_7290.t144 w_109060_7290.t143 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X316 VOUT-.t106 cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 a_109160_2280.t160 a_109160_2280.t159 V_tail_gate.t0 a_109160_2280.t5 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X318 VD2.t14 VIN+ V_source.t40 a_109160_2280.t215 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X319 VOUT+.t14 Y.t42 w_109060_7290.t182 w_109060_7290.t181 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X320 VOUT+.t100 cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VD4.t37 Vb2.t19 Y.t10 VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X322 a_109160_2280.t27 Y.t43 V_CMFB_S3.t4 w_109060_7290.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X323 X.t12 a_109160_2280.t156 a_109160_2280.t158 a_109160_2280.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X324 VOUT+.t101 cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 a_109160_2280.t55 V_tail_gate.t16 V_source.t8 a_109160_2280.t54 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X326 w_109060_7290.t141 w_109060_7290.t139 w_109060_7290.t141 w_109060_7290.t140 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X327 VOUT+.t102 cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT-.t107 cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT-.t108 cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 w_109060_7290.t9 Vb3.t14 VD3.t9 w_109060_7290.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X331 w_109060_7290.t61 Vb3.t15 VD4.t20 w_109060_7290.t60 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X332 VD3.t23 Vb2.t20 X.t9 VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X333 w_109060_7290.t88 X.t42 VOUT-.t10 w_109060_7290.t87 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X334 V_CMFB_S1.t5 X.t43 a_109160_2280.t97 w_109060_7290.t86 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X335 VOUT+.t103 cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 Vb2.t2 Vb2_2.t7 Vb2_2.t9 Vb2_2.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X337 V_CMFB_S2.t3 X.t44 w_109060_7290.t83 a_109160_2280.t96 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X338 w_109060_7290.t29 Y.t44 V_CMFB_S4.t4 a_109160_2280.t32 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X339 VOUT+.t104 cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VD2.t5 Vb1.t22 Y.t5 a_109160_2280.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X341 VOUT+.t105 cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT+.t106 cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT+.t107 cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT-.t109 cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT+.t108 cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VOUT-.t110 cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VOUT-.t111 cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 w_109060_7290.t138 w_109060_7290.t136 Vb2_2.t3 w_109060_7290.t137 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X349 w_109060_7290.t135 w_109060_7290.t133 err_amp_out.t3 w_109060_7290.t134 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X350 VOUT-.t112 cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 a_118660_3088.t0 V_CMFB_S2.t0 a_109160_2280.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X352 VOUT+.t109 cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 a_109160_2280.t95 X.t45 V_CMFB_S1.t4 w_109060_7290.t85 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X354 VOUT+.t110 cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VOUT-.t113 cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT-.t114 cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 VOUT+.t111 cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 w_109060_7290.t84 X.t46 V_CMFB_S2.t2 a_109160_2280.t94 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X359 VOUT-.t115 cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 VOUT+.t112 cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 V_p_mir.t3 VIN+ V_tail_gate.t3 a_109160_2280.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X362 VD2.t13 VIN+ V_source.t39 a_109160_2280.t214 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X363 VOUT+.t1 Y.t45 w_109060_7290.t25 w_109060_7290.t24 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X364 VOUT+.t113 cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 w_109060_7290.t22 Vb3.t16 VD3.t8 w_109060_7290.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X366 VOUT+.t114 cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 VOUT-.t116 cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 VOUT-.t117 cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 VOUT+.t115 cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 VOUT-.t118 cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT-.t119 cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 Vb1.t7 Vb1.t6 Vb1_2.t1 a_109160_2280.t30 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X373 VOUT-.t120 cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 w_109060_7290.t80 X.t47 VOUT-.t9 w_109060_7290.t79 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X375 a_109160_2280.t74 Y.t46 V_CMFB_S3.t3 w_109060_7290.t59 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X376 V_CMFB_S1.t3 X.t48 a_109160_2280.t90 w_109060_7290.t78 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X377 VOUT+.t116 cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VOUT+.t117 cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 VOUT+.t118 cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VOUT+.t119 cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 VD2.t4 Vb1.t23 Y.t4 a_109160_2280.t58 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X382 w_109060_7290.t54 Y.t47 V_CMFB_S4.t3 a_109160_2280.t60 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X383 a_118780_3088.t1 V_tot.t3 a_109160_2280.t82 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X384 VOUT+.t120 cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VOUT-.t121 cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VOUT-.t122 cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 a_109160_2280.t155 a_109160_2280.t153 X.t18 a_109160_2280.t154 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X388 a_109160_2280.t152 a_109160_2280.t150 VOUT+.t11 a_109160_2280.t151 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X389 VOUT+.t121 cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 a_108630_3088.t1 V_CMFB_S3.t0 a_109160_2280.t70 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X391 VOUT-.t123 cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VD3.t36 w_109060_7290.t130 w_109060_7290.t132 w_109060_7290.t131 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X393 VOUT+.t122 cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 V_err_p.t0 V_err_gate.t6 w_109060_7290.t12 w_109060_7290.t11 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X395 VOUT-.t8 X.t49 w_109060_7290.t77 w_109060_7290.t76 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X396 VOUT+.t123 cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VOUT+.t124 cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 a_109160_2280.t91 X.t50 V_CMFB_S1.t2 w_109060_7290.t75 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X399 VOUT+.t125 cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VD2.t12 VIN+ V_source.t32 a_109160_2280.t213 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X401 VOUT-.t124 cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VOUT-.t125 cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 X.t13 VD3.t0 VD3.t2 VD3.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X404 VOUT-.t126 cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VOUT+.t126 cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VOUT-.t0 a_118760_n784.t0 a_109160_2280.t9 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X407 VD1.t12 VIN- V_source.t25 a_109160_2280.t200 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X408 VOUT-.t127 cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT+.t127 cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 Vb1.t3 Vb1.t2 Vb1_2.t0 a_109160_2280.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X411 VD4.t19 Vb3.t17 w_109060_7290.t110 w_109060_7290.t109 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 VOUT+.t128 cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT+.t129 cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT+.t130 cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT+.t131 cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT-.t128 cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VD4.t32 w_109060_7290.t127 w_109060_7290.t129 w_109060_7290.t128 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X418 VOUT-.t129 cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VOUT+.t18 Y.t48 w_109060_7290.t195 w_109060_7290.t194 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X420 VOUT+.t132 cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 w_109060_7290.t74 X.t51 VOUT-.t7 w_109060_7290.t73 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X422 Vb2_2.t1 Vb2.t0 Vb2.t1 Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X423 a_109160_2280.t225 Y.t49 V_CMFB_S3.t2 w_109060_7290.t185 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X424 VOUT-.t130 cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VOUT-.t131 cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT+.t133 cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VD2.t7 Vb1.t24 Y.t8 a_109160_2280.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X428 VOUT-.t132 cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 w_109060_7290.t186 Y.t50 V_CMFB_S4.t2 a_109160_2280.t229 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X430 VD1.t6 Vb1.t25 X.t19 a_109160_2280.t88 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X431 VD1.t5 Vb1.t26 X.t16 a_109160_2280.t63 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X432 VOUT+.t134 cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 a_118780_3088.t0 V_CMFB_S1.t0 a_109160_2280.t72 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X434 VOUT+.t135 cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 a_109160_2280.t80 V_tail_gate.t17 V_source.t7 a_109160_2280.t79 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X436 VOUT-.t133 cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT-.t134 cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 V_err_p.t3 V_tot.t5 err_amp_mir.t4 w_109060_7290.t196 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X439 cap_res_X.t0 X.t1 a_109160_2280.t8 sky130_fd_pr__res_high_po_1p41 l=1.41
X440 VOUT+.t136 cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 VOUT-.t135 cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 err_amp_out.t1 err_amp_mir.t5 a_109160_2280.t23 a_109160_2280.t22 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X443 VOUT-.t6 X.t52 w_109060_7290.t72 w_109060_7290.t71 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X444 VOUT-.t136 cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 V_source.t6 V_tail_gate.t18 a_109160_2280.t6 a_109160_2280.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X446 VOUT-.t137 cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 VOUT-.t138 cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VD2.t11 VIN+ V_source.t37 a_109160_2280.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X449 VOUT-.t139 cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 a_109160_2280.t149 a_109160_2280.t147 V_source.t20 a_109160_2280.t148 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X451 VD3.t7 Vb3.t18 w_109060_7290.t66 w_109060_7290.t65 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X452 VOUT-.t140 cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 w_109060_7290.t70 X.t53 V_CMFB_S2.t1 a_109160_2280.t93 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X454 VOUT+.t137 cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VD1.t11 VIN- V_source.t22 a_109160_2280.t199 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X456 VOUT+.t138 cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 VD1.t10 VIN- V_source.t21 a_109160_2280.t198 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X458 VD4.t18 Vb3.t19 w_109060_7290.t18 w_109060_7290.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X459 VOUT+.t139 cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 w_109060_7290.t126 w_109060_7290.t124 V_err_gate.t1 w_109060_7290.t125 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X461 VOUT-.t141 cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT-.t142 cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VOUT-.t143 cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 X.t21 Vb2.t21 VD3.t21 VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X465 VOUT-.t144 cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT+.t17 Y.t51 w_109060_7290.t193 w_109060_7290.t192 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X467 VOUT+.t140 cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 a_109160_2280.t41 Y.t52 V_CMFB_S3.t1 w_109060_7290.t39 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X469 a_109160_2280.t146 a_109160_2280.t144 VOUT-.t5 a_109160_2280.t145 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X470 V_source.t36 VIN+ VD2.t10 a_109160_2280.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X471 VOUT+.t141 cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT-.t145 cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VD2.t6 Vb1.t27 Y.t7 a_109160_2280.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X474 w_109060_7290.t23 a_109160_2280.t141 a_109160_2280.t143 a_109160_2280.t142 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X475 VOUT+.t142 cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VD1.t3 Vb1.t28 X.t7 a_109160_2280.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X477 a_108510_3088.t0 V_CMFB_S4.t0 a_109160_2280.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X478 VOUT+.t143 cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VD4.t35 Vb2.t22 Y.t9 VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X480 VOUT+.t144 cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT-.t146 cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 a_109160_2280.t140 a_109160_2280.t138 w_109060_7290.t117 a_109160_2280.t139 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X483 V_source.t5 V_tail_gate.t19 a_109160_2280.t235 a_109160_2280.t234 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X484 VOUT+.t145 cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT-.t147 cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 err_amp_mir.t2 a_109160_2280.t135 a_109160_2280.t137 a_109160_2280.t136 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X487 VOUT+.t146 cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 a_109160_2280.t21 V_tail_gate.t20 V_source.t4 a_109160_2280.t20 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X489 a_109160_2280.t92 X.t54 V_CMFB_S1.t1 w_109060_7290.t67 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X490 VD3.t19 Vb2.t23 X.t22 VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X491 VOUT+.t147 cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 V_b_2nd_stage.t0 a_118760_n784.t1 a_109160_2280.t13 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X493 VOUT-.t148 cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VOUT+.t148 cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 Y.t1 Vb1.t29 VD2.t1 a_109160_2280.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X496 VOUT-.t149 cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VD2.t8 a_109160_2280.t132 a_109160_2280.t134 a_109160_2280.t133 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X498 a_109160_2280.t69 V_tail_gate.t21 V_p_mir.t0 a_109160_2280.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X499 VD1.t9 VIN- V_source.t26 a_109160_2280.t197 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X500 VOUT-.t150 cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VOUT+.t10 a_109160_2280.t129 a_109160_2280.t131 a_109160_2280.t130 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X502 VOUT+.t149 cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 VOUT-.t151 cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VOUT-.t152 cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 VOUT-.t153 cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 w_109060_7290.t51 Vb3.t20 VD4.t17 w_109060_7290.t50 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X507 V_source.t3 V_tail_gate.t22 a_109160_2280.t35 a_109160_2280.t34 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X508 VOUT-.t154 cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 V_err_mir_p.t0 V_err_gate.t7 w_109060_7290.t38 w_109060_7290.t37 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X510 w_109060_7290.t14 Vb3.t21 VD4.t16 w_109060_7290.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X511 Vb2_2.t6 Vb2_2.t4 Vb2_2.t6 Vb2_2.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X512 a_109160_2280.t57 V_tail_gate.t23 V_source.t2 a_109160_2280.t56 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X513 VOUT+.t3 Y.t53 w_109060_7290.t42 w_109060_7290.t41 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X514 VOUT+.t150 cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VOUT+.t6 V_b_2nd_stage.t9 a_109160_2280.t111 a_109160_2280.t110 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X516 VOUT-.t155 cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VOUT+.t151 cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 a_109160_2280.t208 w_109060_7290.t121 w_109060_7290.t123 w_109060_7290.t122 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X519 VOUT+.t152 cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT-.t4 a_109160_2280.t126 a_109160_2280.t128 a_109160_2280.t127 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X521 w_109060_7290.t120 w_109060_7290.t118 a_109160_2280.t207 w_109060_7290.t119 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X522 VOUT-.t156 cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VD1.t4 Vb1.t30 X.t11 a_109160_2280.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X524 VOUT+.t153 cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 V_CMFB_S4.t1 Y.t54 w_109060_7290.t180 a_109160_2280.t221 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X526 w_109060_7290.t5 Vb3.t22 VD3.t6 w_109060_7290.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X527 VOUT+.t154 cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VD3.t17 Vb2.t24 X.t10 VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X529 Y.t21 VD4.t26 VD4.t28 VD4.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X530 VOUT+.t155 cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT+.t156 cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 X.n51 X.t25 1172.87
R1 X.n47 X.t51 1172.87
R2 X.n51 X.t38 996.134
R3 X.n52 X.t49 996.134
R4 X.n53 X.t34 996.134
R5 X.n54 X.t52 996.134
R6 X.n50 X.t42 996.134
R7 X.n49 X.t30 996.134
R8 X.n48 X.t47 996.134
R9 X.n47 X.t33 996.134
R10 X.n18 X.t53 690.867
R11 X.n17 X.t44 690.867
R12 X.n27 X.t54 530.201
R13 X.n26 X.t48 530.201
R14 X.n24 X.t40 514.134
R15 X.n23 X.t26 514.134
R16 X.n22 X.t37 514.134
R17 X.n21 X.t46 514.134
R18 X.n20 X.t29 514.134
R19 X.n19 X.t41 514.134
R20 X.n18 X.t35 514.134
R21 X.n17 X.t28 514.134
R22 X.n27 X.t36 353.467
R23 X.n28 X.t45 353.467
R24 X.n29 X.t32 353.467
R25 X.n30 X.t50 353.467
R26 X.n31 X.t39 353.467
R27 X.n32 X.t27 353.467
R28 X.n33 X.t43 353.467
R29 X.n26 X.t31 353.467
R30 X.n50 X.n49 176.733
R31 X.n49 X.n48 176.733
R32 X.n48 X.n47 176.733
R33 X.n52 X.n51 176.733
R34 X.n53 X.n52 176.733
R35 X.n54 X.n53 176.733
R36 X.n28 X.n27 176.733
R37 X.n29 X.n28 176.733
R38 X.n30 X.n29 176.733
R39 X.n31 X.n30 176.733
R40 X.n32 X.n31 176.733
R41 X.n33 X.n32 176.733
R42 X.n19 X.n18 176.733
R43 X.n20 X.n19 176.733
R44 X.n21 X.n20 176.733
R45 X.n22 X.n21 176.733
R46 X.n23 X.n22 176.733
R47 X.n24 X.n23 176.733
R48 X.n35 X.n34 165.472
R49 X.n35 X.n25 165.472
R50 X.n57 X.n56 152
R51 X.n58 X.n57 131.571
R52 X.n57 X.n55 124.517
R53 X.n125 X.n35 74.5362
R54 X.n79 X.n78 66.0338
R55 X.n77 X.n76 66.0338
R56 X.n89 X.n88 66.0338
R57 X.n85 X.n84 66.0338
R58 X.n82 X.n81 66.0338
R59 X.n75 X.n74 66.0338
R60 X.n6 X.n5 49.3505
R61 X.n10 X.n9 49.3505
R62 X.n134 X.n133 49.3505
R63 X.n140 X.n139 49.3505
R64 X.n143 X.n142 49.3505
R65 X.n147 X.n146 49.3505
R66 X.n41 X.t1 41.0384
R67 X.n55 X.n50 40.1672
R68 X.n55 X.n54 40.1672
R69 X.n34 X.n26 40.1672
R70 X.n34 X.n33 40.1672
R71 X.n25 X.n17 40.1672
R72 X.n25 X.n24 40.1672
R73 X.n59 X.n58 16.3217
R74 X.n5 X.t24 16.0005
R75 X.n5 X.t12 16.0005
R76 X.n9 X.t18 16.0005
R77 X.n9 X.t23 16.0005
R78 X.n133 X.t16 16.0005
R79 X.n133 X.t4 16.0005
R80 X.n139 X.t19 16.0005
R81 X.n139 X.t20 16.0005
R82 X.n142 X.t7 16.0005
R83 X.n142 X.t3 16.0005
R84 X.n146 X.t11 16.0005
R85 X.n146 X.t5 16.0005
R86 X.n56 X.n46 12.8005
R87 X.n78 X.t22 11.2576
R88 X.n78 X.t13 11.2576
R89 X.n76 X.t14 11.2576
R90 X.n76 X.t17 11.2576
R91 X.n88 X.t6 11.2576
R92 X.n88 X.t21 11.2576
R93 X.n84 X.t9 11.2576
R94 X.n84 X.t15 11.2576
R95 X.n81 X.t2 11.2576
R96 X.n81 X.t0 11.2576
R97 X.n74 X.t10 11.2576
R98 X.n74 X.t8 11.2576
R99 X.n56 X.n44 9.36264
R100 X.n46 X.n45 9.3005
R101 X.n87 X.n77 5.91717
R102 X.n80 X.n79 5.91717
R103 X.n10 X.n8 5.6255
R104 X.n145 X.n6 5.6255
R105 X.n58 X.n46 5.33141
R106 X.n89 X.n87 5.29217
R107 X.n86 X.n85 5.29217
R108 X.n83 X.n82 5.29217
R109 X.n80 X.n75 5.29217
R110 X.n94 X.n73 5.1255
R111 X.n91 X.n65 5.1255
R112 X.n134 X.n8 5.063
R113 X.n141 X.n140 5.063
R114 X.n144 X.n143 5.063
R115 X.n147 X.n145 5.063
R116 X.n150 X.n149 5.063
R117 X.n136 X.n11 5.063
R118 X.n95 X.n94 4.5005
R119 X.n93 X.n71 4.5005
R120 X.n92 X.n68 4.5005
R121 X.n91 X.n90 4.5005
R122 X.n119 X.n118 4.5005
R123 X.n149 X.n148 4.5005
R124 X.n7 X.n3 4.5005
R125 X.n138 X.n137 4.5005
R126 X.n136 X.n135 4.5005
R127 X.n124 X.n61 4.5005
R128 X.n126 X.n125 4.5005
R129 X.n125 X.n124 4.5005
R130 X.n60 X.n59 4.5005
R131 X.n38 X.n37 4.5005
R132 X.n120 X.n63 2.26187
R133 X.n40 X.n39 2.26187
R134 X.n39 X.n36 2.26187
R135 X.n117 X.n63 2.26187
R136 X.n121 X.n62 2.24063
R137 X.n126 X.n15 2.24063
R138 X.n16 X.n14 2.24063
R139 X.n117 X.n116 2.24063
R140 X.n123 X.n122 2.24063
R141 X.n41 X.n40 2.24063
R142 X.n43 X.n42 2.24063
R143 X.n60 X.n44 2.22018
R144 X.n98 X.n72 1.5005
R145 X.n100 X.n99 1.5005
R146 X.n101 X.n70 1.5005
R147 X.n103 X.n102 1.5005
R148 X.n104 X.n69 1.5005
R149 X.n106 X.n105 1.5005
R150 X.n107 X.n67 1.5005
R151 X.n109 X.n108 1.5005
R152 X.n110 X.n66 1.5005
R153 X.n112 X.n111 1.5005
R154 X.n113 X.n64 1.5005
R155 X.n115 X.n114 1.5005
R156 X.n153 X.n152 1.5005
R157 X.n154 X.n1 1.5005
R158 X.n156 X.n155 1.5005
R159 X.n2 X.n0 1.5005
R160 X.n130 X.n13 1.5005
R161 X.n132 X.n131 1.5005
R162 X.n129 X.n12 1.5005
R163 X.n128 X.n127 1.5005
R164 X.n151 X.n150 1.43397
R165 X.n135 X.n132 1.3755
R166 X.n138 X.n2 1.3755
R167 X.n154 X.n3 1.3755
R168 X.n148 X.n4 1.3755
R169 X.n127 X.n11 1.3755
R170 X.n122 X.n121 0.979667
R171 X.n90 X.n89 0.792167
R172 X.n85 X.n68 0.792167
R173 X.n82 X.n71 0.792167
R174 X.n95 X.n75 0.792167
R175 X.n77 X.n65 0.792167
R176 X.n79 X.n73 0.792167
R177 X.n60 X.n43 0.682792
R178 X.n128 X.n126 0.630708
R179 X.n94 X.n93 0.6255
R180 X.n93 X.n92 0.6255
R181 X.n92 X.n91 0.6255
R182 X.n87 X.n86 0.6255
R183 X.n86 X.n83 0.6255
R184 X.n83 X.n80 0.6255
R185 X.n116 X.n115 0.609875
R186 X.n152 X.n151 0.564601
R187 X.n149 X.n7 0.563
R188 X.n137 X.n7 0.563
R189 X.n137 X.n136 0.563
R190 X.n141 X.n8 0.563
R191 X.n144 X.n141 0.563
R192 X.n145 X.n144 0.563
R193 X.n97 X.n73 0.533638
R194 X.n90 X.n66 0.46925
R195 X.n106 X.n68 0.46925
R196 X.n101 X.n71 0.46925
R197 X.n96 X.n95 0.46925
R198 X.n114 X.n65 0.46925
R199 X.n124 X.n60 0.46925
R200 X.n98 X.n97 0.427973
R201 X.n135 X.n134 0.3755
R202 X.n140 X.n138 0.3755
R203 X.n143 X.n3 0.3755
R204 X.n148 X.n147 0.3755
R205 X.n11 X.n10 0.3755
R206 X.n150 X.n6 0.3755
R207 X.n59 X.n45 0.1255
R208 X.n45 X.n44 0.0626438
R209 X.n97 X.n96 0.0587394
R210 X.n127 X.n12 0.0577917
R211 X.n132 X.n12 0.0577917
R212 X.n132 X.n13 0.0577917
R213 X.n13 X.n2 0.0577917
R214 X.n155 X.n2 0.0577917
R215 X.n155 X.n154 0.0577917
R216 X.n154 X.n153 0.0577917
R217 X.n153 X.n4 0.0577917
R218 X.n129 X.n128 0.0577917
R219 X.n131 X.n129 0.0577917
R220 X.n131 X.n130 0.0577917
R221 X.n130 X.n0 0.0577917
R222 X.n156 X.n1 0.0577917
R223 X.n152 X.n1 0.0577917
R224 X.n151 X.n4 0.054517
R225 X.n114 X.n113 0.0421667
R226 X.n113 X.n112 0.0421667
R227 X.n112 X.n66 0.0421667
R228 X.n108 X.n66 0.0421667
R229 X.n108 X.n107 0.0421667
R230 X.n107 X.n106 0.0421667
R231 X.n106 X.n69 0.0421667
R232 X.n102 X.n69 0.0421667
R233 X.n102 X.n101 0.0421667
R234 X.n101 X.n100 0.0421667
R235 X.n100 X.n72 0.0421667
R236 X.n96 X.n72 0.0421667
R237 X.n115 X.n64 0.0421667
R238 X.n111 X.n64 0.0421667
R239 X.n111 X.n110 0.0421667
R240 X.n110 X.n109 0.0421667
R241 X.n109 X.n67 0.0421667
R242 X.n105 X.n67 0.0421667
R243 X.n105 X.n104 0.0421667
R244 X.n104 X.n103 0.0421667
R245 X.n103 X.n70 0.0421667
R246 X.n99 X.n70 0.0421667
R247 X.n99 X.n98 0.0421667
R248 X.n126 X.n14 0.0421667
R249 X X.n156 0.0369583
R250 X.n116 X.n62 0.0217373
R251 X.n120 X.n119 0.0217373
R252 X.n122 X.n15 0.0217373
R253 X.n125 X.n16 0.0217373
R254 X.n118 X.n62 0.0217373
R255 X.n121 X.n120 0.0217373
R256 X.n43 X.n36 0.0217373
R257 X.n61 X.n15 0.0217373
R258 X.n61 X.n16 0.0217373
R259 X.n39 X.n37 0.0217373
R260 X.n38 X.n36 0.0217373
R261 X.n118 X.n63 0.0217373
R262 X.n119 X.n117 0.0217373
R263 X.n40 X.n38 0.0217373
R264 X.n124 X.n123 0.0217373
R265 X.n123 X.n14 0.0217373
R266 X.n42 X.n37 0.0217373
R267 X.n42 X.n41 0.0217373
R268 X X.n0 0.0213333
R269 w_109060_7290.n173 w_109060_7290.t170 1231.74
R270 w_109060_7290.n176 w_109060_7290.t173 1231.74
R271 w_109060_7290.n48 w_109060_7290.t149 1231.74
R272 w_109060_7290.n51 w_109060_7290.t158 1231.74
R273 w_109060_7290.n121 w_109060_7290.t133 826.801
R274 w_109060_7290.n153 w_109060_7290.t146 826.801
R275 w_109060_7290.n127 w_109060_7290.t124 826.801
R276 w_109060_7290.n21 w_109060_7290.t176 826.801
R277 w_109060_7290.n73 w_109060_7290.t167 672.293
R278 w_109060_7290.n76 w_109060_7290.t127 672.293
R279 w_109060_7290.n57 w_109060_7290.t152 672.293
R280 w_109060_7290.n54 w_109060_7290.t130 672.293
R281 w_109060_7290.n100 w_109060_7290.t139 661.375
R282 w_109060_7290.n103 w_109060_7290.t161 661.375
R283 w_109060_7290.n33 w_109060_7290.t155 589.076
R284 w_109060_7290.n36 w_109060_7290.t164 589.076
R285 w_109060_7290.n169 w_109060_7290.t118 589.076
R286 w_109060_7290.n166 w_109060_7290.t121 589.076
R287 w_109060_7290.n152 w_109060_7290.n15 585
R288 w_109060_7290.n140 w_109060_7290.n139 585
R289 w_109060_7290.n137 w_109060_7290.n136 585
R290 w_109060_7290.n120 w_109060_7290.n119 585
R291 w_109060_7290.n96 w_109060_7290.t136 456.526
R292 w_109060_7290.n93 w_109060_7290.t142 456.526
R293 w_109060_7290.n95 w_109060_7290.t137 397.784
R294 w_109060_7290.t143 w_109060_7290.n94 397.784
R295 w_109060_7290.t156 w_109060_7290.n34 343.882
R296 w_109060_7290.n35 w_109060_7290.t165 343.882
R297 w_109060_7290.n168 w_109060_7290.t119 343.882
R298 w_109060_7290.t122 w_109060_7290.n167 343.882
R299 w_109060_7290.n139 w_109060_7290.n131 291.053
R300 w_109060_7290.n139 w_109060_7290.n138 291.053
R301 w_109060_7290.n136 w_109060_7290.n129 291.053
R302 w_109060_7290.n136 w_109060_7290.n135 291.053
R303 w_109060_7290.n145 w_109060_7290.n15 290.233
R304 w_109060_7290.n146 w_109060_7290.n15 290.233
R305 w_109060_7290.n119 w_109060_7290.n109 290.233
R306 w_109060_7290.n119 w_109060_7290.n118 290.233
R307 w_109060_7290.t137 w_109060_7290.t183 259.091
R308 w_109060_7290.t183 w_109060_7290.t143 259.091
R309 w_109060_7290.n146 w_109060_7290.n143 242.903
R310 w_109060_7290.n118 w_109060_7290.n117 242.903
R311 w_109060_7290.n152 w_109060_7290.n151 238.367
R312 w_109060_7290.n141 w_109060_7290.n140 238.367
R313 w_109060_7290.n137 w_109060_7290.n18 238.367
R314 w_109060_7290.n116 w_109060_7290.t134 221.121
R315 w_109060_7290.n142 w_109060_7290.t177 221.121
R316 w_109060_7290.t125 w_109060_7290.n142 221.121
R317 w_109060_7290.n150 w_109060_7290.t147 221.121
R318 w_109060_7290.t67 w_109060_7290.t156 217.708
R319 w_109060_7290.t92 w_109060_7290.t67 217.708
R320 w_109060_7290.t85 w_109060_7290.t92 217.708
R321 w_109060_7290.t98 w_109060_7290.t85 217.708
R322 w_109060_7290.t75 w_109060_7290.t98 217.708
R323 w_109060_7290.t89 w_109060_7290.t75 217.708
R324 w_109060_7290.t103 w_109060_7290.t89 217.708
R325 w_109060_7290.t86 w_109060_7290.t103 217.708
R326 w_109060_7290.t99 w_109060_7290.t86 217.708
R327 w_109060_7290.t78 w_109060_7290.t99 217.708
R328 w_109060_7290.t165 w_109060_7290.t78 217.708
R329 w_109060_7290.t119 w_109060_7290.t40 217.708
R330 w_109060_7290.t40 w_109060_7290.t62 217.708
R331 w_109060_7290.t62 w_109060_7290.t19 217.708
R332 w_109060_7290.t19 w_109060_7290.t31 217.708
R333 w_109060_7290.t31 w_109060_7290.t59 217.708
R334 w_109060_7290.t59 w_109060_7290.t47 217.708
R335 w_109060_7290.t47 w_109060_7290.t185 217.708
R336 w_109060_7290.t185 w_109060_7290.t197 217.708
R337 w_109060_7290.t197 w_109060_7290.t39 217.708
R338 w_109060_7290.t39 w_109060_7290.t20 217.708
R339 w_109060_7290.t20 w_109060_7290.t122 217.708
R340 w_109060_7290.n14 w_109060_7290.n13 216.677
R341 w_109060_7290.n124 w_109060_7290.n123 216.677
R342 w_109060_7290.t140 w_109060_7290.n101 213.131
R343 w_109060_7290.n102 w_109060_7290.t162 213.131
R344 w_109060_7290.t168 w_109060_7290.n74 213.131
R345 w_109060_7290.n75 w_109060_7290.t128 213.131
R346 w_109060_7290.n56 w_109060_7290.t153 213.131
R347 w_109060_7290.t131 w_109060_7290.n55 213.131
R348 w_109060_7290.n130 w_109060_7290.n20 185
R349 w_109060_7290.n134 w_109060_7290.n19 185
R350 w_109060_7290.n142 w_109060_7290.n19 185
R351 w_109060_7290.n133 w_109060_7290.n132 185
R352 w_109060_7290.n17 w_109060_7290.n16 185
R353 w_109060_7290.n149 w_109060_7290.n148 185
R354 w_109060_7290.n150 w_109060_7290.n149 185
R355 w_109060_7290.n147 w_109060_7290.n144 185
R356 w_109060_7290.n120 w_109060_7290.n107 185
R357 w_109060_7290.n116 w_109060_7290.n107 185
R358 w_109060_7290.n112 w_109060_7290.n108 185
R359 w_109060_7290.n114 w_109060_7290.n113 185
R360 w_109060_7290.n111 w_109060_7290.n110 185
R361 w_109060_7290.t134 w_109060_7290.t36 180.173
R362 w_109060_7290.t36 w_109060_7290.t11 180.173
R363 w_109060_7290.t11 w_109060_7290.t15 180.173
R364 w_109060_7290.t15 w_109060_7290.t196 180.173
R365 w_109060_7290.t196 w_109060_7290.t177 180.173
R366 w_109060_7290.t191 w_109060_7290.t125 180.173
R367 w_109060_7290.t37 w_109060_7290.t191 180.173
R368 w_109060_7290.t2 w_109060_7290.t37 180.173
R369 w_109060_7290.t32 w_109060_7290.t2 180.173
R370 w_109060_7290.t147 w_109060_7290.t32 180.173
R371 w_109060_7290.n95 w_109060_7290.t138 168.139
R372 w_109060_7290.n94 w_109060_7290.t145 168.139
R373 w_109060_7290.n92 w_109060_7290.n91 150.643
R374 w_109060_7290.n149 w_109060_7290.n17 150
R375 w_109060_7290.n149 w_109060_7290.n144 150
R376 w_109060_7290.n20 w_109060_7290.n19 150
R377 w_109060_7290.n132 w_109060_7290.n19 150
R378 w_109060_7290.n112 w_109060_7290.n107 150
R379 w_109060_7290.n114 w_109060_7290.n111 150
R380 w_109060_7290.t6 w_109060_7290.t140 146.155
R381 w_109060_7290.t162 w_109060_7290.t6 146.155
R382 w_109060_7290.t52 w_109060_7290.t168 146.155
R383 w_109060_7290.t50 w_109060_7290.t52 146.155
R384 w_109060_7290.t109 w_109060_7290.t50 146.155
R385 w_109060_7290.t60 w_109060_7290.t109 146.155
R386 w_109060_7290.t57 w_109060_7290.t60 146.155
R387 w_109060_7290.t113 w_109060_7290.t57 146.155
R388 w_109060_7290.t107 w_109060_7290.t113 146.155
R389 w_109060_7290.t27 w_109060_7290.t107 146.155
R390 w_109060_7290.t17 w_109060_7290.t27 146.155
R391 w_109060_7290.t13 w_109060_7290.t17 146.155
R392 w_109060_7290.t128 w_109060_7290.t13 146.155
R393 w_109060_7290.t153 w_109060_7290.t198 146.155
R394 w_109060_7290.t198 w_109060_7290.t48 146.155
R395 w_109060_7290.t48 w_109060_7290.t65 146.155
R396 w_109060_7290.t65 w_109060_7290.t21 146.155
R397 w_109060_7290.t21 w_109060_7290.t115 146.155
R398 w_109060_7290.t115 w_109060_7290.t8 146.155
R399 w_109060_7290.t8 w_109060_7290.t63 146.155
R400 w_109060_7290.t63 w_109060_7290.t111 146.155
R401 w_109060_7290.t111 w_109060_7290.t0 146.155
R402 w_109060_7290.t0 w_109060_7290.t4 146.155
R403 w_109060_7290.t4 w_109060_7290.t131 146.155
R404 w_109060_7290.n34 w_109060_7290.t157 136.701
R405 w_109060_7290.n35 w_109060_7290.t166 136.701
R406 w_109060_7290.n168 w_109060_7290.t120 136.701
R407 w_109060_7290.n167 w_109060_7290.t123 136.701
R408 w_109060_7290.t171 w_109060_7290.n174 122.829
R409 w_109060_7290.n175 w_109060_7290.t174 122.829
R410 w_109060_7290.t150 w_109060_7290.n49 122.829
R411 w_109060_7290.n50 w_109060_7290.t159 122.829
R412 w_109060_7290.t181 w_109060_7290.t171 81.6411
R413 w_109060_7290.t189 w_109060_7290.t181 81.6411
R414 w_109060_7290.t24 w_109060_7290.t189 81.6411
R415 w_109060_7290.t187 w_109060_7290.t24 81.6411
R416 w_109060_7290.t194 w_109060_7290.t187 81.6411
R417 w_109060_7290.t55 w_109060_7290.t194 81.6411
R418 w_109060_7290.t192 w_109060_7290.t55 81.6411
R419 w_109060_7290.t44 w_109060_7290.t192 81.6411
R420 w_109060_7290.t41 w_109060_7290.t44 81.6411
R421 w_109060_7290.t33 w_109060_7290.t41 81.6411
R422 w_109060_7290.t174 w_109060_7290.t33 81.6411
R423 w_109060_7290.t105 w_109060_7290.t150 81.6411
R424 w_109060_7290.t90 w_109060_7290.t105 81.6411
R425 w_109060_7290.t76 w_109060_7290.t90 81.6411
R426 w_109060_7290.t93 w_109060_7290.t76 81.6411
R427 w_109060_7290.t71 w_109060_7290.t93 81.6411
R428 w_109060_7290.t87 w_109060_7290.t71 81.6411
R429 w_109060_7290.t100 w_109060_7290.t87 81.6411
R430 w_109060_7290.t79 w_109060_7290.t100 81.6411
R431 w_109060_7290.t96 w_109060_7290.t79 81.6411
R432 w_109060_7290.t73 w_109060_7290.t96 81.6411
R433 w_109060_7290.t159 w_109060_7290.t73 81.6411
R434 w_109060_7290.n101 w_109060_7290.t141 76.2576
R435 w_109060_7290.n102 w_109060_7290.t163 76.2576
R436 w_109060_7290.n74 w_109060_7290.t169 76.2576
R437 w_109060_7290.n75 w_109060_7290.t129 76.2576
R438 w_109060_7290.n56 w_109060_7290.t154 76.2576
R439 w_109060_7290.n55 w_109060_7290.t132 76.2576
R440 w_109060_7290.n79 w_109060_7290.n78 71.3255
R441 w_109060_7290.n81 w_109060_7290.n80 71.3255
R442 w_109060_7290.n86 w_109060_7290.n85 71.3255
R443 w_109060_7290.n88 w_109060_7290.n87 71.3255
R444 w_109060_7290.n69 w_109060_7290.n68 71.3255
R445 w_109060_7290.n67 w_109060_7290.n66 71.3255
R446 w_109060_7290.n62 w_109060_7290.n61 71.3255
R447 w_109060_7290.n60 w_109060_7290.n59 71.3255
R448 w_109060_7290.n99 w_109060_7290.n98 68.4557
R449 w_109060_7290.n83 w_109060_7290.n82 66.8255
R450 w_109060_7290.n64 w_109060_7290.n63 66.8255
R451 w_109060_7290.n142 w_109060_7290.n141 65.8183
R452 w_109060_7290.n142 w_109060_7290.n18 65.8183
R453 w_109060_7290.n151 w_109060_7290.n150 65.8183
R454 w_109060_7290.n150 w_109060_7290.n143 65.8183
R455 w_109060_7290.n116 w_109060_7290.n115 65.8183
R456 w_109060_7290.n117 w_109060_7290.n116 65.8183
R457 w_109060_7290.n153 w_109060_7290.n152 58.0576
R458 w_109060_7290.n121 w_109060_7290.n120 58.0576
R459 w_109060_7290.n128 w_109060_7290.n127 54.4005
R460 w_109060_7290.n128 w_109060_7290.n21 54.4005
R461 w_109060_7290.n144 w_109060_7290.n143 53.3664
R462 w_109060_7290.n132 w_109060_7290.n18 53.3664
R463 w_109060_7290.n141 w_109060_7290.n20 53.3664
R464 w_109060_7290.n151 w_109060_7290.n17 53.3664
R465 w_109060_7290.n115 w_109060_7290.n112 53.3664
R466 w_109060_7290.n117 w_109060_7290.n111 53.3664
R467 w_109060_7290.n115 w_109060_7290.n114 53.3664
R468 w_109060_7290.n174 w_109060_7290.t172 40.9789
R469 w_109060_7290.n175 w_109060_7290.t175 40.9789
R470 w_109060_7290.n49 w_109060_7290.t151 40.9789
R471 w_109060_7290.n50 w_109060_7290.t160 40.9789
R472 w_109060_7290.n184 w_109060_7290.n183 38.2287
R473 w_109060_7290.n178 w_109060_7290.n177 38.2279
R474 w_109060_7290.n180 w_109060_7290.n179 38.2279
R475 w_109060_7290.n182 w_109060_7290.n181 38.2279
R476 w_109060_7290.n12 w_109060_7290.n11 38.2279
R477 w_109060_7290.n39 w_109060_7290.n38 38.2279
R478 w_109060_7290.n41 w_109060_7290.n40 38.2279
R479 w_109060_7290.n43 w_109060_7290.n42 38.2279
R480 w_109060_7290.n45 w_109060_7290.n44 38.2279
R481 w_109060_7290.n47 w_109060_7290.n46 38.2279
R482 w_109060_7290.n157 w_109060_7290.n155 26.9096
R483 w_109060_7290.n24 w_109060_7290.n22 26.8887
R484 w_109060_7290.n157 w_109060_7290.n156 26.795
R485 w_109060_7290.n159 w_109060_7290.n158 26.795
R486 w_109060_7290.n161 w_109060_7290.n160 26.795
R487 w_109060_7290.n163 w_109060_7290.n162 26.795
R488 w_109060_7290.n165 w_109060_7290.n164 26.795
R489 w_109060_7290.n32 w_109060_7290.n31 26.7741
R490 w_109060_7290.n30 w_109060_7290.n29 26.7741
R491 w_109060_7290.n28 w_109060_7290.n27 26.7741
R492 w_109060_7290.n26 w_109060_7290.n25 26.7741
R493 w_109060_7290.n24 w_109060_7290.n23 26.7741
R494 w_109060_7290.n91 w_109060_7290.t184 21.8894
R495 w_109060_7290.n91 w_109060_7290.t144 21.8894
R496 w_109060_7290.n119 w_109060_7290.t135 15.7605
R497 w_109060_7290.n15 w_109060_7290.t148 15.7605
R498 w_109060_7290.n136 w_109060_7290.t126 15.7605
R499 w_109060_7290.n139 w_109060_7290.t178 15.7605
R500 w_109060_7290.n13 w_109060_7290.t38 15.7605
R501 w_109060_7290.n13 w_109060_7290.t3 15.7605
R502 w_109060_7290.n123 w_109060_7290.t12 15.7605
R503 w_109060_7290.n123 w_109060_7290.t16 15.7605
R504 w_109060_7290.t141 w_109060_7290.n99 11.2576
R505 w_109060_7290.n99 w_109060_7290.t7 11.2576
R506 w_109060_7290.n78 w_109060_7290.t18 11.2576
R507 w_109060_7290.n78 w_109060_7290.t14 11.2576
R508 w_109060_7290.n80 w_109060_7290.t108 11.2576
R509 w_109060_7290.n80 w_109060_7290.t28 11.2576
R510 w_109060_7290.n82 w_109060_7290.t58 11.2576
R511 w_109060_7290.n82 w_109060_7290.t114 11.2576
R512 w_109060_7290.n85 w_109060_7290.t110 11.2576
R513 w_109060_7290.n85 w_109060_7290.t61 11.2576
R514 w_109060_7290.n87 w_109060_7290.t53 11.2576
R515 w_109060_7290.n87 w_109060_7290.t51 11.2576
R516 w_109060_7290.n68 w_109060_7290.t1 11.2576
R517 w_109060_7290.n68 w_109060_7290.t5 11.2576
R518 w_109060_7290.n66 w_109060_7290.t64 11.2576
R519 w_109060_7290.n66 w_109060_7290.t112 11.2576
R520 w_109060_7290.n63 w_109060_7290.t116 11.2576
R521 w_109060_7290.n63 w_109060_7290.t9 11.2576
R522 w_109060_7290.n61 w_109060_7290.t66 11.2576
R523 w_109060_7290.n61 w_109060_7290.t22 11.2576
R524 w_109060_7290.n59 w_109060_7290.t199 11.2576
R525 w_109060_7290.n59 w_109060_7290.t49 11.2576
R526 w_109060_7290.n122 w_109060_7290.n121 10.8696
R527 w_109060_7290.n125 w_109060_7290.n21 10.869
R528 w_109060_7290.n127 w_109060_7290.n126 10.869
R529 w_109060_7290.n154 w_109060_7290.n153 10.869
R530 w_109060_7290.n152 w_109060_7290.n16 9.14336
R531 w_109060_7290.n148 w_109060_7290.n147 9.14336
R532 w_109060_7290.n120 w_109060_7290.n108 9.14336
R533 w_109060_7290.n113 w_109060_7290.n110 9.14336
R534 w_109060_7290.n31 w_109060_7290.t83 8.0005
R535 w_109060_7290.n31 w_109060_7290.t200 8.0005
R536 w_109060_7290.n29 w_109060_7290.t81 8.0005
R537 w_109060_7290.n29 w_109060_7290.t102 8.0005
R538 w_109060_7290.n27 w_109060_7290.t69 8.0005
R539 w_109060_7290.n27 w_109060_7290.t104 8.0005
R540 w_109060_7290.n25 w_109060_7290.t95 8.0005
R541 w_109060_7290.n25 w_109060_7290.t84 8.0005
R542 w_109060_7290.n23 w_109060_7290.t68 8.0005
R543 w_109060_7290.n23 w_109060_7290.t82 8.0005
R544 w_109060_7290.n22 w_109060_7290.t179 8.0005
R545 w_109060_7290.n22 w_109060_7290.t70 8.0005
R546 w_109060_7290.n155 w_109060_7290.t46 8.0005
R547 w_109060_7290.n155 w_109060_7290.t23 8.0005
R548 w_109060_7290.n156 w_109060_7290.t30 8.0005
R549 w_109060_7290.n156 w_109060_7290.t186 8.0005
R550 w_109060_7290.n158 w_109060_7290.t35 8.0005
R551 w_109060_7290.n158 w_109060_7290.t54 8.0005
R552 w_109060_7290.n160 w_109060_7290.t26 8.0005
R553 w_109060_7290.n160 w_109060_7290.t29 8.0005
R554 w_109060_7290.n162 w_109060_7290.t180 8.0005
R555 w_109060_7290.n162 w_109060_7290.t43 8.0005
R556 w_109060_7290.n164 w_109060_7290.t117 8.0005
R557 w_109060_7290.n164 w_109060_7290.t10 8.0005
R558 w_109060_7290.n177 w_109060_7290.t42 6.56717
R559 w_109060_7290.n177 w_109060_7290.t34 6.56717
R560 w_109060_7290.n179 w_109060_7290.t193 6.56717
R561 w_109060_7290.n179 w_109060_7290.t45 6.56717
R562 w_109060_7290.n181 w_109060_7290.t195 6.56717
R563 w_109060_7290.n181 w_109060_7290.t56 6.56717
R564 w_109060_7290.n11 w_109060_7290.t182 6.56717
R565 w_109060_7290.n11 w_109060_7290.t190 6.56717
R566 w_109060_7290.n38 w_109060_7290.t97 6.56717
R567 w_109060_7290.n38 w_109060_7290.t74 6.56717
R568 w_109060_7290.n40 w_109060_7290.t101 6.56717
R569 w_109060_7290.n40 w_109060_7290.t80 6.56717
R570 w_109060_7290.n42 w_109060_7290.t72 6.56717
R571 w_109060_7290.n42 w_109060_7290.t88 6.56717
R572 w_109060_7290.n44 w_109060_7290.t77 6.56717
R573 w_109060_7290.n44 w_109060_7290.t94 6.56717
R574 w_109060_7290.n46 w_109060_7290.t106 6.56717
R575 w_109060_7290.n46 w_109060_7290.t91 6.56717
R576 w_109060_7290.t25 w_109060_7290.n184 6.56717
R577 w_109060_7290.n184 w_109060_7290.t188 6.56717
R578 w_109060_7290.n89 w_109060_7290.n88 5.1255
R579 w_109060_7290.n79 w_109060_7290.n77 5.1255
R580 w_109060_7290.n60 w_109060_7290.n58 5.1255
R581 w_109060_7290.n70 w_109060_7290.n69 5.1255
R582 w_109060_7290.n145 w_109060_7290.n16 4.53698
R583 w_109060_7290.n147 w_109060_7290.n146 4.53698
R584 w_109060_7290.n148 w_109060_7290.n145 4.53698
R585 w_109060_7290.n109 w_109060_7290.n108 4.53698
R586 w_109060_7290.n118 w_109060_7290.n110 4.53698
R587 w_109060_7290.n113 w_109060_7290.n109 4.53698
R588 w_109060_7290.n84 w_109060_7290.n83 4.5005
R589 w_109060_7290.n65 w_109060_7290.n64 4.5005
R590 w_109060_7290.n1 w_109060_7290.n0 0.499598
R591 w_109060_7290.n171 w_109060_7290.n6 0.0428468
R592 w_109060_7290.n5 w_109060_7290.n6 1.10813
R593 w_109060_7290.n9 w_109060_7290.n8 1.48724
R594 w_109060_7290.n106 w_109060_7290.n105 3.06776
R595 w_109060_7290.n37 w_109060_7290.n33 2.96402
R596 w_109060_7290.n170 w_109060_7290.n166 2.96402
R597 w_109060_7290.n130 w_109060_7290.n129 2.8957
R598 w_109060_7290.n131 w_109060_7290.n130 2.8957
R599 w_109060_7290.n135 w_109060_7290.n133 2.8957
R600 w_109060_7290.n138 w_109060_7290.n133 2.8957
R601 w_109060_7290.n134 w_109060_7290.n131 2.8957
R602 w_109060_7290.n138 w_109060_7290.n137 2.8957
R603 w_109060_7290.n140 w_109060_7290.n129 2.8957
R604 w_109060_7290.n135 w_109060_7290.n134 2.8957
R605 w_109060_7290.n94 w_109060_7290.n93 2.8255
R606 w_109060_7290.n96 w_109060_7290.n95 2.8255
R607 w_109060_7290.n58 w_109060_7290.n53 2.53694
R608 w_109060_7290.n77 w_109060_7290.n72 2.53694
R609 w_109060_7290.n36 w_109060_7290.n35 2.423
R610 w_109060_7290.n34 w_109060_7290.n33 2.423
R611 w_109060_7290.n167 w_109060_7290.n166 2.423
R612 w_109060_7290.n169 w_109060_7290.n168 2.423
R613 w_109060_7290.n140 w_109060_7290.n128 2.32777
R614 w_109060_7290.n37 w_109060_7290.n36 2.27652
R615 w_109060_7290.n170 w_109060_7290.n169 2.27652
R616 w_109060_7290.n71 w_109060_7290.n2 0.273728
R617 w_109060_7290.n171 w_109060_7290.n7 2.24063
R618 w_109060_7290.n8 w_109060_7290.n7 0.0150284
R619 w_109060_7290.n10 w_109060_7290.n170 0.772221
R620 w_109060_7290.n0 w_109060_7290.n2 1.46695
R621 w_109060_7290.n83 w_109060_7290.n72 2.16194
R622 w_109060_7290.n90 w_109060_7290.n89 2.16194
R623 w_109060_7290.n64 w_109060_7290.n53 2.16194
R624 w_109060_7290.n71 w_109060_7290.n70 2.16194
R625 w_109060_7290.n105 w_109060_7290.n104 2.12369
R626 w_109060_7290.n176 w_109060_7290.n175 1.97758
R627 w_109060_7290.n174 w_109060_7290.n173 1.97758
R628 w_109060_7290.n51 w_109060_7290.n50 1.97758
R629 w_109060_7290.n49 w_109060_7290.n48 1.97758
R630 w_109060_7290.n178 w_109060_7290.n176 1.95361
R631 w_109060_7290.n48 w_109060_7290.n47 1.95361
R632 w_109060_7290.n103 w_109060_7290.n102 1.888
R633 w_109060_7290.n101 w_109060_7290.n100 1.888
R634 w_109060_7290.n173 w_109060_7290.n172 1.83902
R635 w_109060_7290.n52 w_109060_7290.n51 1.83902
R636 w_109060_7290.n93 w_109060_7290.n92 1.63212
R637 w_109060_7290.n100 w_109060_7290.n98 1.63212
R638 w_109060_7290.n105 w_109060_7290.n97 1.59823
R639 w_109060_7290.n97 w_109060_7290.n96 1.56962
R640 w_109060_7290.n104 w_109060_7290.n103 1.56962
R641 w_109060_7290.n106 w_109060_7290.n3 1.36639
R642 w_109060_7290.n7 w_109060_7290.n10 1.17421
R643 w_109060_7290.n10 w_109060_7290.n165 1.98877
R644 w_109060_7290.n76 w_109060_7290.n75 1.03383
R645 w_109060_7290.n74 w_109060_7290.n73 1.03383
R646 w_109060_7290.n55 w_109060_7290.n54 1.03383
R647 w_109060_7290.n57 w_109060_7290.n56 1.03383
R648 w_109060_7290.n122 w_109060_7290.n1 0.971472
R649 w_109060_7290.n9 w_109060_7290.n154 0.932792
R650 w_109060_7290.n5 w_109060_7290.n3 1.43582
R651 w_109060_7290.n77 w_109060_7290.n76 0.792167
R652 w_109060_7290.n89 w_109060_7290.n73 0.792167
R653 w_109060_7290.n70 w_109060_7290.n54 0.792167
R654 w_109060_7290.n58 w_109060_7290.n57 0.792167
R655 w_109060_7290.n88 w_109060_7290.n86 0.6255
R656 w_109060_7290.n86 w_109060_7290.n84 0.6255
R657 w_109060_7290.n84 w_109060_7290.n81 0.6255
R658 w_109060_7290.n81 w_109060_7290.n79 0.6255
R659 w_109060_7290.n62 w_109060_7290.n60 0.6255
R660 w_109060_7290.n65 w_109060_7290.n62 0.6255
R661 w_109060_7290.n67 w_109060_7290.n65 0.6255
R662 w_109060_7290.n69 w_109060_7290.n67 0.6255
R663 w_109060_7290.n71 w_109060_7290.n53 0.3755
R664 w_109060_7290.n90 w_109060_7290.n72 0.3755
R665 w_109060_7290.n4 w_109060_7290.n32 1.97074
R666 w_109060_7290.n4 w_109060_7290.n37 0.764993
R667 w_109060_7290.n172 w_109060_7290.n171 0.266125
R668 w_109060_7290.n3 w_109060_7290.n90 0.273866
R669 w_109060_7290.n124 w_109060_7290.n122 0.172375
R670 w_109060_7290.n125 w_109060_7290.n124 0.172375
R671 w_109060_7290.n126 w_109060_7290.n14 0.172375
R672 w_109060_7290.n154 w_109060_7290.n14 0.172375
R673 w_109060_7290.n97 w_109060_7290.n92 0.1255
R674 w_109060_7290.n104 w_109060_7290.n98 0.1255
R675 w_109060_7290.n26 w_109060_7290.n24 0.115083
R676 w_109060_7290.n28 w_109060_7290.n26 0.115083
R677 w_109060_7290.n30 w_109060_7290.n28 0.115083
R678 w_109060_7290.n32 w_109060_7290.n30 0.115083
R679 w_109060_7290.n165 w_109060_7290.n163 0.115083
R680 w_109060_7290.n163 w_109060_7290.n161 0.115083
R681 w_109060_7290.n161 w_109060_7290.n159 0.115083
R682 w_109060_7290.n159 w_109060_7290.n157 0.115083
R683 w_109060_7290.n47 w_109060_7290.n45 0.115083
R684 w_109060_7290.n45 w_109060_7290.n43 0.115083
R685 w_109060_7290.n43 w_109060_7290.n41 0.115083
R686 w_109060_7290.n41 w_109060_7290.n39 0.115083
R687 w_109060_7290.n52 w_109060_7290.n39 0.115083
R688 w_109060_7290.n172 w_109060_7290.n12 0.115083
R689 w_109060_7290.n183 w_109060_7290.n12 0.115083
R690 w_109060_7290.n183 w_109060_7290.n182 0.115083
R691 w_109060_7290.n182 w_109060_7290.n180 0.115083
R692 w_109060_7290.n180 w_109060_7290.n178 0.115083
R693 w_109060_7290.n126 w_109060_7290.n125 0.0838333
R694 w_109060_7290.n106 w_109060_7290.n2 1.36571
R695 w_109060_7290.n1 w_109060_7290.n52 0.313661
R696 w_109060_7290.n8 w_109060_7290.n5 0.071655
R697 w_109060_7290.n9 w_109060_7290.n6 0.043506
R698 w_109060_7290.n4 w_109060_7290.n0 1.17842
R699 VOUT-.n193 VOUT-.t0 110.191
R700 VOUT-.n44 VOUT-.n43 34.9935
R701 VOUT-.n33 VOUT-.n32 34.9935
R702 VOUT-.n35 VOUT-.n34 34.9935
R703 VOUT-.n38 VOUT-.n37 34.9935
R704 VOUT-.n41 VOUT-.n40 34.9935
R705 VOUT-.n47 VOUT-.n46 34.9935
R706 VOUT-.n180 VOUT-.n179 9.73997
R707 VOUT-.n176 VOUT-.n175 9.73997
R708 VOUT-.n183 VOUT-.n182 9.73997
R709 VOUT-.n181 VOUT-.n176 6.64633
R710 VOUT-.n181 VOUT-.n180 6.64633
R711 VOUT-.n43 VOUT-.t7 6.56717
R712 VOUT-.n43 VOUT-.t17 6.56717
R713 VOUT-.n32 VOUT-.t16 6.56717
R714 VOUT-.n32 VOUT-.t15 6.56717
R715 VOUT-.n34 VOUT-.t11 6.56717
R716 VOUT-.n34 VOUT-.t8 6.56717
R717 VOUT-.n37 VOUT-.t12 6.56717
R718 VOUT-.n37 VOUT-.t6 6.56717
R719 VOUT-.n40 VOUT-.t10 6.56717
R720 VOUT-.n40 VOUT-.t14 6.56717
R721 VOUT-.n46 VOUT-.t9 6.56717
R722 VOUT-.n46 VOUT-.t13 6.56717
R723 VOUT-.n36 VOUT-.n33 6.3755
R724 VOUT-.n45 VOUT-.n44 6.3755
R725 VOUT-.n183 VOUT-.n181 6.02133
R726 VOUT-.n36 VOUT-.n35 5.813
R727 VOUT-.n39 VOUT-.n38 5.813
R728 VOUT-.n42 VOUT-.n41 5.813
R729 VOUT-.n47 VOUT-.n45 5.813
R730 VOUT-.n51 VOUT-.n31 5.063
R731 VOUT-.n48 VOUT-.n24 5.063
R732 VOUT-.n114 VOUT-.t114 4.8295
R733 VOUT-.n113 VOUT-.t148 4.8295
R734 VOUT-.n112 VOUT-.t45 4.8295
R735 VOUT-.n111 VOUT-.t94 4.8295
R736 VOUT-.n110 VOUT-.t129 4.8295
R737 VOUT-.n109 VOUT-.t32 4.8295
R738 VOUT-.n115 VOUT-.t58 4.8295
R739 VOUT-.n126 VOUT-.t69 4.8295
R740 VOUT-.n127 VOUT-.t120 4.8295
R741 VOUT-.n129 VOUT-.t105 4.8295
R742 VOUT-.n130 VOUT-.t86 4.8295
R743 VOUT-.n132 VOUT-.t60 4.8295
R744 VOUT-.n133 VOUT-.t46 4.8295
R745 VOUT-.n135 VOUT-.t21 4.8295
R746 VOUT-.n136 VOUT-.t146 4.8295
R747 VOUT-.n138 VOUT-.t55 4.8295
R748 VOUT-.n139 VOUT-.t40 4.8295
R749 VOUT-.n141 VOUT-.t156 4.8295
R750 VOUT-.n142 VOUT-.t141 4.8295
R751 VOUT-.n144 VOUT-.t118 4.8295
R752 VOUT-.n145 VOUT-.t103 4.8295
R753 VOUT-.n147 VOUT-.t152 4.8295
R754 VOUT-.n148 VOUT-.t135 4.8295
R755 VOUT-.n150 VOUT-.t110 4.8295
R756 VOUT-.n151 VOUT-.t95 4.8295
R757 VOUT-.n153 VOUT-.t71 4.8295
R758 VOUT-.n154 VOUT-.t54 4.8295
R759 VOUT-.n76 VOUT-.t155 4.8295
R760 VOUT-.n78 VOUT-.t115 4.8295
R761 VOUT-.n91 VOUT-.t149 4.8295
R762 VOUT-.n92 VOUT-.t57 4.8295
R763 VOUT-.n94 VOUT-.t132 4.8295
R764 VOUT-.n95 VOUT-.t116 4.8295
R765 VOUT-.n97 VOUT-.t109 4.8295
R766 VOUT-.n98 VOUT-.t80 4.8295
R767 VOUT-.n100 VOUT-.t75 4.8295
R768 VOUT-.n101 VOUT-.t48 4.8295
R769 VOUT-.n103 VOUT-.t25 4.8295
R770 VOUT-.n104 VOUT-.t150 4.8295
R771 VOUT-.n106 VOUT-.t67 4.8295
R772 VOUT-.n107 VOUT-.t52 4.8295
R773 VOUT-.n156 VOUT-.t107 4.8295
R774 VOUT-.n117 VOUT-.t68 4.8154
R775 VOUT-.n79 VOUT-.t38 4.806
R776 VOUT-.n80 VOUT-.t76 4.806
R777 VOUT-.n81 VOUT-.t113 4.806
R778 VOUT-.n82 VOUT-.t154 4.806
R779 VOUT-.n83 VOUT-.t128 4.806
R780 VOUT-.n84 VOUT-.t27 4.806
R781 VOUT-.n85 VOUT-.t65 4.806
R782 VOUT-.n86 VOUT-.t44 4.806
R783 VOUT-.n87 VOUT-.t82 4.806
R784 VOUT-.n88 VOUT-.t63 4.806
R785 VOUT-.n89 VOUT-.t41 4.806
R786 VOUT-.n114 VOUT-.t47 4.5005
R787 VOUT-.n113 VOUT-.t84 4.5005
R788 VOUT-.n112 VOUT-.t122 4.5005
R789 VOUT-.n111 VOUT-.t101 4.5005
R790 VOUT-.n110 VOUT-.t138 4.5005
R791 VOUT-.n109 VOUT-.t139 4.5005
R792 VOUT-.n125 VOUT-.t102 4.5005
R793 VOUT-.n124 VOUT-.t61 4.5005
R794 VOUT-.n123 VOUT-.t85 4.5005
R795 VOUT-.n122 VOUT-.t106 4.5005
R796 VOUT-.n121 VOUT-.t64 4.5005
R797 VOUT-.n120 VOUT-.t88 4.5005
R798 VOUT-.n119 VOUT-.t51 4.5005
R799 VOUT-.n118 VOUT-.t151 4.5005
R800 VOUT-.n117 VOUT-.t31 4.5005
R801 VOUT-.n116 VOUT-.t134 4.5005
R802 VOUT-.n115 VOUT-.t99 4.5005
R803 VOUT-.n126 VOUT-.t30 4.5005
R804 VOUT-.n128 VOUT-.t133 4.5005
R805 VOUT-.n127 VOUT-.t98 4.5005
R806 VOUT-.n129 VOUT-.t66 4.5005
R807 VOUT-.n131 VOUT-.t28 4.5005
R808 VOUT-.n130 VOUT-.t136 4.5005
R809 VOUT-.n132 VOUT-.t24 4.5005
R810 VOUT-.n134 VOUT-.t130 4.5005
R811 VOUT-.n133 VOUT-.t97 4.5005
R812 VOUT-.n135 VOUT-.t125 4.5005
R813 VOUT-.n137 VOUT-.t93 4.5005
R814 VOUT-.n136 VOUT-.t56 4.5005
R815 VOUT-.n138 VOUT-.t20 4.5005
R816 VOUT-.n140 VOUT-.t124 4.5005
R817 VOUT-.n139 VOUT-.t92 4.5005
R818 VOUT-.n141 VOUT-.t121 4.5005
R819 VOUT-.n143 VOUT-.t87 4.5005
R820 VOUT-.n142 VOUT-.t53 4.5005
R821 VOUT-.n144 VOUT-.t83 4.5005
R822 VOUT-.n146 VOUT-.t50 4.5005
R823 VOUT-.n145 VOUT-.t153 4.5005
R824 VOUT-.n147 VOUT-.t117 4.5005
R825 VOUT-.n149 VOUT-.t81 4.5005
R826 VOUT-.n148 VOUT-.t49 4.5005
R827 VOUT-.n150 VOUT-.t77 4.5005
R828 VOUT-.n152 VOUT-.t42 4.5005
R829 VOUT-.n151 VOUT-.t147 4.5005
R830 VOUT-.n153 VOUT-.t36 4.5005
R831 VOUT-.n155 VOUT-.t144 4.5005
R832 VOUT-.n154 VOUT-.t108 4.5005
R833 VOUT-.n76 VOUT-.t119 4.5005
R834 VOUT-.n77 VOUT-.t79 4.5005
R835 VOUT-.n78 VOUT-.t78 4.5005
R836 VOUT-.n90 VOUT-.t39 4.5005
R837 VOUT-.n89 VOUT-.t142 4.5005
R838 VOUT-.n88 VOUT-.t22 4.5005
R839 VOUT-.n87 VOUT-.t43 4.5005
R840 VOUT-.n86 VOUT-.t145 4.5005
R841 VOUT-.n85 VOUT-.t23 4.5005
R842 VOUT-.n84 VOUT-.t127 4.5005
R843 VOUT-.n83 VOUT-.t90 4.5005
R844 VOUT-.n82 VOUT-.t112 4.5005
R845 VOUT-.n81 VOUT-.t74 4.5005
R846 VOUT-.n80 VOUT-.t34 4.5005
R847 VOUT-.n79 VOUT-.t140 4.5005
R848 VOUT-.n91 VOUT-.t111 4.5005
R849 VOUT-.n93 VOUT-.t73 4.5005
R850 VOUT-.n92 VOUT-.t33 4.5005
R851 VOUT-.n94 VOUT-.t100 4.5005
R852 VOUT-.n96 VOUT-.t62 4.5005
R853 VOUT-.n95 VOUT-.t26 4.5005
R854 VOUT-.n97 VOUT-.t19 4.5005
R855 VOUT-.n99 VOUT-.t72 4.5005
R856 VOUT-.n98 VOUT-.t123 4.5005
R857 VOUT-.n100 VOUT-.t126 4.5005
R858 VOUT-.n102 VOUT-.t37 4.5005
R859 VOUT-.n101 VOUT-.t89 4.5005
R860 VOUT-.n103 VOUT-.t131 4.5005
R861 VOUT-.n105 VOUT-.t96 4.5005
R862 VOUT-.n104 VOUT-.t59 4.5005
R863 VOUT-.n106 VOUT-.t29 4.5005
R864 VOUT-.n108 VOUT-.t137 4.5005
R865 VOUT-.n107 VOUT-.t104 4.5005
R866 VOUT-.n156 VOUT-.t70 4.5005
R867 VOUT-.n157 VOUT-.t35 4.5005
R868 VOUT-.n158 VOUT-.t143 4.5005
R869 VOUT-.n159 VOUT-.t91 4.5005
R870 VOUT-.n52 VOUT-.n51 4.5005
R871 VOUT-.n50 VOUT-.n29 4.5005
R872 VOUT-.n49 VOUT-.n28 4.5005
R873 VOUT-.n48 VOUT-.n25 4.5005
R874 VOUT-.n70 VOUT-.n69 4.5005
R875 VOUT-.n21 VOUT-.n18 4.5005
R876 VOUT-.n70 VOUT-.n18 4.5005
R877 VOUT-.n71 VOUT-.n14 4.5005
R878 VOUT-.n71 VOUT-.n16 4.5005
R879 VOUT-.n71 VOUT-.n70 4.5005
R880 VOUT-.n168 VOUT-.n74 4.5005
R881 VOUT-.n169 VOUT-.n168 4.5005
R882 VOUT-.n169 VOUT-.n10 4.5005
R883 VOUT-.n170 VOUT-.n9 4.5005
R884 VOUT-.n170 VOUT-.n169 4.5005
R885 VOUT-.n197 VOUT-.n196 4.5005
R886 VOUT-.n172 VOUT-.n5 4.5005
R887 VOUT-.n197 VOUT-.n5 4.5005
R888 VOUT-.n198 VOUT-.n1 4.5005
R889 VOUT-.n198 VOUT-.n3 4.5005
R890 VOUT-.n198 VOUT-.n197 4.5005
R891 VOUT-.n179 VOUT-.t18 3.42907
R892 VOUT-.n179 VOUT-.t4 3.42907
R893 VOUT-.n175 VOUT-.t5 3.42907
R894 VOUT-.n175 VOUT-.t2 3.42907
R895 VOUT-.n182 VOUT-.t3 3.42907
R896 VOUT-.n182 VOUT-.t1 3.42907
R897 VOUT-.n68 VOUT-.n67 2.24601
R898 VOUT-.n19 VOUT-.n13 2.24601
R899 VOUT-.n195 VOUT-.n194 2.24601
R900 VOUT-.n6 VOUT-.n0 2.24601
R901 VOUT-.n167 VOUT-.n166 2.24477
R902 VOUT-.n12 VOUT-.n7 2.24477
R903 VOUT-.n71 VOUT-.n15 2.24063
R904 VOUT-.n170 VOUT-.n8 2.24063
R905 VOUT-.n198 VOUT-.n2 2.24063
R906 VOUT-.n18 VOUT-.n17 2.24063
R907 VOUT-.n168 VOUT-.n72 2.24063
R908 VOUT-.n73 VOUT-.n10 2.24063
R909 VOUT-.n5 VOUT-.n4 2.24063
R910 VOUT-.n69 VOUT-.n22 2.23934
R911 VOUT-.n69 VOUT-.n20 2.23934
R912 VOUT-.n196 VOUT-.n173 2.23934
R913 VOUT-.n196 VOUT-.n171 2.23934
R914 VOUT-.n180 VOUT-.n178 1.62886
R915 VOUT-.n191 VOUT-.n176 1.52133
R916 VOUT-.n184 VOUT-.n183 1.52133
R917 VOUT-.n186 VOUT-.n185 1.5005
R918 VOUT-.n187 VOUT-.n177 1.5005
R919 VOUT-.n189 VOUT-.n188 1.5005
R920 VOUT-.n190 VOUT-.n174 1.5005
R921 VOUT-.n192 VOUT-.n191 1.5005
R922 VOUT-.n55 VOUT-.n30 1.5005
R923 VOUT-.n57 VOUT-.n56 1.5005
R924 VOUT-.n58 VOUT-.n27 1.5005
R925 VOUT-.n60 VOUT-.n59 1.5005
R926 VOUT-.n61 VOUT-.n26 1.5005
R927 VOUT-.n63 VOUT-.n62 1.5005
R928 VOUT-.n64 VOUT-.n23 1.5005
R929 VOUT-.n66 VOUT-.n65 1.5005
R930 VOUT-.n35 VOUT-.n25 1.313
R931 VOUT-.n38 VOUT-.n28 1.313
R932 VOUT-.n41 VOUT-.n29 1.313
R933 VOUT-.n52 VOUT-.n47 1.313
R934 VOUT-.n33 VOUT-.n24 1.313
R935 VOUT-.n44 VOUT-.n31 1.313
R936 VOUT-.n166 VOUT-.n165 1.1455
R937 VOUT-.n160 VOUT-.n11 1.13717
R938 VOUT-.n162 VOUT-.n161 1.13717
R939 VOUT-.n164 VOUT-.n163 1.13717
R940 VOUT-.n169 VOUT-.n11 1.13717
R941 VOUT-.n162 VOUT-.n12 1.13717
R942 VOUT-.n163 VOUT-.n9 1.13717
R943 VOUT-.n75 VOUT-.n74 1.13717
R944 VOUT-.n54 VOUT-.n31 0.715216
R945 VOUT-.n63 VOUT-.n25 0.65675
R946 VOUT-.n59 VOUT-.n28 0.65675
R947 VOUT-.n57 VOUT-.n29 0.65675
R948 VOUT-.n53 VOUT-.n52 0.65675
R949 VOUT-.n65 VOUT-.n24 0.65675
R950 VOUT-.n165 VOUT-.n164 0.585
R951 VOUT-.n196 VOUT-.n170 0.5705
R952 VOUT-.n55 VOUT-.n54 0.564601
R953 VOUT-.n51 VOUT-.n50 0.563
R954 VOUT-.n50 VOUT-.n49 0.563
R955 VOUT-.n49 VOUT-.n48 0.563
R956 VOUT-.n39 VOUT-.n36 0.563
R957 VOUT-.n42 VOUT-.n39 0.563
R958 VOUT-.n45 VOUT-.n42 0.563
R959 VOUT-.n67 VOUT-.n66 0.495292
R960 VOUT-.n193 VOUT-.n192 0.380708
R961 VOUT-.n125 VOUT-.n109 0.3295
R962 VOUT-.n125 VOUT-.n124 0.3295
R963 VOUT-.n124 VOUT-.n123 0.3295
R964 VOUT-.n123 VOUT-.n122 0.3295
R965 VOUT-.n122 VOUT-.n121 0.3295
R966 VOUT-.n121 VOUT-.n120 0.3295
R967 VOUT-.n120 VOUT-.n119 0.3295
R968 VOUT-.n119 VOUT-.n118 0.3295
R969 VOUT-.n118 VOUT-.n117 0.3295
R970 VOUT-.n117 VOUT-.n116 0.3295
R971 VOUT-.n116 VOUT-.n115 0.3295
R972 VOUT-.n128 VOUT-.n126 0.3295
R973 VOUT-.n128 VOUT-.n127 0.3295
R974 VOUT-.n131 VOUT-.n129 0.3295
R975 VOUT-.n131 VOUT-.n130 0.3295
R976 VOUT-.n134 VOUT-.n132 0.3295
R977 VOUT-.n134 VOUT-.n133 0.3295
R978 VOUT-.n137 VOUT-.n135 0.3295
R979 VOUT-.n137 VOUT-.n136 0.3295
R980 VOUT-.n140 VOUT-.n138 0.3295
R981 VOUT-.n140 VOUT-.n139 0.3295
R982 VOUT-.n143 VOUT-.n141 0.3295
R983 VOUT-.n143 VOUT-.n142 0.3295
R984 VOUT-.n146 VOUT-.n144 0.3295
R985 VOUT-.n146 VOUT-.n145 0.3295
R986 VOUT-.n149 VOUT-.n147 0.3295
R987 VOUT-.n149 VOUT-.n148 0.3295
R988 VOUT-.n152 VOUT-.n150 0.3295
R989 VOUT-.n152 VOUT-.n151 0.3295
R990 VOUT-.n155 VOUT-.n153 0.3295
R991 VOUT-.n155 VOUT-.n154 0.3295
R992 VOUT-.n77 VOUT-.n76 0.3295
R993 VOUT-.n90 VOUT-.n78 0.3295
R994 VOUT-.n90 VOUT-.n89 0.3295
R995 VOUT-.n89 VOUT-.n88 0.3295
R996 VOUT-.n88 VOUT-.n87 0.3295
R997 VOUT-.n87 VOUT-.n86 0.3295
R998 VOUT-.n86 VOUT-.n85 0.3295
R999 VOUT-.n85 VOUT-.n84 0.3295
R1000 VOUT-.n84 VOUT-.n83 0.3295
R1001 VOUT-.n83 VOUT-.n82 0.3295
R1002 VOUT-.n82 VOUT-.n81 0.3295
R1003 VOUT-.n81 VOUT-.n80 0.3295
R1004 VOUT-.n80 VOUT-.n79 0.3295
R1005 VOUT-.n93 VOUT-.n91 0.3295
R1006 VOUT-.n93 VOUT-.n92 0.3295
R1007 VOUT-.n96 VOUT-.n94 0.3295
R1008 VOUT-.n96 VOUT-.n95 0.3295
R1009 VOUT-.n99 VOUT-.n97 0.3295
R1010 VOUT-.n99 VOUT-.n98 0.3295
R1011 VOUT-.n102 VOUT-.n100 0.3295
R1012 VOUT-.n102 VOUT-.n101 0.3295
R1013 VOUT-.n105 VOUT-.n103 0.3295
R1014 VOUT-.n105 VOUT-.n104 0.3295
R1015 VOUT-.n108 VOUT-.n106 0.3295
R1016 VOUT-.n108 VOUT-.n107 0.3295
R1017 VOUT-.n157 VOUT-.n156 0.3295
R1018 VOUT-.n158 VOUT-.n157 0.3295
R1019 VOUT-.n118 VOUT-.n114 0.3154
R1020 VOUT-.n186 VOUT-.n178 0.314966
R1021 VOUT-.n159 VOUT-.n158 0.3107
R1022 VOUT-.n119 VOUT-.n113 0.306
R1023 VOUT-.n120 VOUT-.n112 0.306
R1024 VOUT-.n121 VOUT-.n111 0.306
R1025 VOUT-.n122 VOUT-.n110 0.306
R1026 VOUT-.n128 VOUT-.n125 0.2825
R1027 VOUT-.n131 VOUT-.n128 0.2825
R1028 VOUT-.n134 VOUT-.n131 0.2825
R1029 VOUT-.n137 VOUT-.n134 0.2825
R1030 VOUT-.n140 VOUT-.n137 0.2825
R1031 VOUT-.n143 VOUT-.n140 0.2825
R1032 VOUT-.n146 VOUT-.n143 0.2825
R1033 VOUT-.n149 VOUT-.n146 0.2825
R1034 VOUT-.n152 VOUT-.n149 0.2825
R1035 VOUT-.n155 VOUT-.n152 0.2825
R1036 VOUT-.n90 VOUT-.n77 0.2825
R1037 VOUT-.n93 VOUT-.n90 0.2825
R1038 VOUT-.n96 VOUT-.n93 0.2825
R1039 VOUT-.n99 VOUT-.n96 0.2825
R1040 VOUT-.n102 VOUT-.n99 0.2825
R1041 VOUT-.n105 VOUT-.n102 0.2825
R1042 VOUT-.n108 VOUT-.n105 0.2825
R1043 VOUT-.n157 VOUT-.n108 0.2825
R1044 VOUT-.n157 VOUT-.n155 0.2825
R1045 VOUT-.n168 VOUT-.n71 0.2655
R1046 VOUT-.n194 VOUT-.n193 0.193208
R1047 VOUT-.n160 VOUT-.n159 0.138367
R1048 VOUT-.n184 VOUT-.n178 0.0891864
R1049 VOUT-.n65 VOUT-.n64 0.0577917
R1050 VOUT-.n64 VOUT-.n63 0.0577917
R1051 VOUT-.n63 VOUT-.n26 0.0577917
R1052 VOUT-.n59 VOUT-.n26 0.0577917
R1053 VOUT-.n59 VOUT-.n58 0.0577917
R1054 VOUT-.n58 VOUT-.n57 0.0577917
R1055 VOUT-.n57 VOUT-.n30 0.0577917
R1056 VOUT-.n53 VOUT-.n30 0.0577917
R1057 VOUT-.n66 VOUT-.n23 0.0577917
R1058 VOUT-.n62 VOUT-.n23 0.0577917
R1059 VOUT-.n62 VOUT-.n61 0.0577917
R1060 VOUT-.n61 VOUT-.n60 0.0577917
R1061 VOUT-.n60 VOUT-.n27 0.0577917
R1062 VOUT-.n56 VOUT-.n27 0.0577917
R1063 VOUT-.n56 VOUT-.n55 0.0577917
R1064 VOUT-.n54 VOUT-.n53 0.054517
R1065 VOUT-.n191 VOUT-.n190 0.0421667
R1066 VOUT-.n190 VOUT-.n189 0.0421667
R1067 VOUT-.n189 VOUT-.n177 0.0421667
R1068 VOUT-.n185 VOUT-.n177 0.0421667
R1069 VOUT-.n185 VOUT-.n184 0.0421667
R1070 VOUT-.n197 VOUT-.n6 0.0421667
R1071 VOUT-.n192 VOUT-.n174 0.0421667
R1072 VOUT-.n188 VOUT-.n174 0.0421667
R1073 VOUT-.n188 VOUT-.n187 0.0421667
R1074 VOUT-.n187 VOUT-.n186 0.0421667
R1075 VOUT-.n169 VOUT-.n12 0.0421667
R1076 VOUT-.n70 VOUT-.n19 0.0421667
R1077 VOUT-.n171 VOUT-.n6 0.0243161
R1078 VOUT-.n173 VOUT-.n1 0.0243161
R1079 VOUT-.n20 VOUT-.n19 0.0243161
R1080 VOUT-.n22 VOUT-.n14 0.0243161
R1081 VOUT-.n22 VOUT-.n21 0.0243161
R1082 VOUT-.n20 VOUT-.n16 0.0243161
R1083 VOUT-.n173 VOUT-.n172 0.0243161
R1084 VOUT-.n171 VOUT-.n3 0.0243161
R1085 VOUT-.n194 VOUT-.n2 0.0217373
R1086 VOUT-.n166 VOUT-.n8 0.0217373
R1087 VOUT-.n67 VOUT-.n15 0.0217373
R1088 VOUT-.n21 VOUT-.n15 0.0217373
R1089 VOUT-.n74 VOUT-.n8 0.0217373
R1090 VOUT-.n172 VOUT-.n2 0.0217373
R1091 VOUT-.n4 VOUT-.n1 0.0217373
R1092 VOUT-.n72 VOUT-.n12 0.0217373
R1093 VOUT-.n74 VOUT-.n73 0.0217373
R1094 VOUT-.n17 VOUT-.n14 0.0217373
R1095 VOUT-.n17 VOUT-.n16 0.0217373
R1096 VOUT-.n72 VOUT-.n9 0.0217373
R1097 VOUT-.n73 VOUT-.n9 0.0217373
R1098 VOUT-.n4 VOUT-.n3 0.0217373
R1099 VOUT-.n161 VOUT-.n160 0.0161667
R1100 VOUT-.n164 VOUT-.n161 0.0161667
R1101 VOUT-.n162 VOUT-.n11 0.0161667
R1102 VOUT-.n163 VOUT-.n162 0.0161667
R1103 VOUT-.n163 VOUT-.n75 0.0161667
R1104 VOUT-.n167 VOUT-.n10 0.0134654
R1105 VOUT-.n170 VOUT-.n7 0.0134654
R1106 VOUT-.n168 VOUT-.n167 0.0134654
R1107 VOUT-.n10 VOUT-.n7 0.0134654
R1108 VOUT-.n68 VOUT-.n18 0.0109778
R1109 VOUT-.n71 VOUT-.n13 0.0109778
R1110 VOUT-.n195 VOUT-.n5 0.0109778
R1111 VOUT-.n198 VOUT-.n0 0.0109778
R1112 VOUT-.n69 VOUT-.n68 0.0109778
R1113 VOUT-.n18 VOUT-.n13 0.0109778
R1114 VOUT-.n196 VOUT-.n195 0.0109778
R1115 VOUT-.n5 VOUT-.n0 0.0109778
R1116 VOUT- VOUT-.n198 0.0105
R1117 VOUT-.n165 VOUT-.n75 0.00872683
R1118 V_b_2nd_stage.n4 V_b_2nd_stage.t7 525.38
R1119 V_b_2nd_stage.n3 V_b_2nd_stage.t3 525.38
R1120 V_b_2nd_stage.n0 V_b_2nd_stage.t5 525.38
R1121 V_b_2nd_stage.n1 V_b_2nd_stage.t4 525.38
R1122 V_b_2nd_stage.n5 V_b_2nd_stage.n4 491.151
R1123 V_b_2nd_stage.n2 V_b_2nd_stage.n1 491.151
R1124 V_b_2nd_stage.n4 V_b_2nd_stage.t2 281.168
R1125 V_b_2nd_stage.n3 V_b_2nd_stage.t8 281.168
R1126 V_b_2nd_stage.n1 V_b_2nd_stage.t6 281.168
R1127 V_b_2nd_stage.n0 V_b_2nd_stage.t9 281.168
R1128 V_b_2nd_stage.n4 V_b_2nd_stage.n3 244.214
R1129 V_b_2nd_stage.n1 V_b_2nd_stage.n0 244.214
R1130 V_b_2nd_stage.n2 V_b_2nd_stage.t1 118.129
R1131 V_b_2nd_stage.t0 V_b_2nd_stage.n5 118.129
R1132 V_b_2nd_stage.n5 V_b_2nd_stage.n2 23.3755
R1133 a_109160_2280.n287 a_109160_2280.n2 13324.2
R1134 a_109160_2280.n285 a_109160_2280.n3 7587.98
R1135 a_109160_2280.n3 a_109160_2280.n2 7511.38
R1136 a_109160_2280.n125 a_109160_2280.n2 7511.38
R1137 a_109160_2280.t71 a_109160_2280.n288 5812.12
R1138 a_109160_2280.n287 a_109160_2280.n286 4034.11
R1139 a_109160_2280.n288 a_109160_2280.n1 3925.98
R1140 a_109160_2280.n289 a_109160_2280.n1 3882.89
R1141 a_109160_2280.n286 a_109160_2280.t8 3757.09
R1142 a_109160_2280.n286 a_109160_2280.n3 3080.82
R1143 a_109160_2280.n288 a_109160_2280.n287 2918.74
R1144 a_109160_2280.n285 a_109160_2280.t73 2321.39
R1145 a_109160_2280.t8 a_109160_2280.n285 1161.6
R1146 a_109160_2280.n277 a_109160_2280.n276 932.912
R1147 a_109160_2280.n255 a_109160_2280.n254 932.912
R1148 a_109160_2280.n282 a_109160_2280.t170 749.742
R1149 a_109160_2280.n203 a_109160_2280.t141 747.734
R1150 a_109160_2280.n252 a_109160_2280.t138 747.734
R1151 a_109160_2280.n279 a_109160_2280.t181 747.734
R1152 a_109160_2280.n271 a_109160_2280.t147 659.367
R1153 a_109160_2280.n186 a_109160_2280.t193 659.367
R1154 a_109160_2280.n147 a_109160_2280.t135 659.367
R1155 a_109160_2280.n117 a_109160_2280.t173 659.367
R1156 a_109160_2280.n125 a_109160_2280.n1 577.346
R1157 a_109160_2280.n239 a_109160_2280.t129 524.808
R1158 a_109160_2280.n249 a_109160_2280.t150 524.808
R1159 a_109160_2280.n11 a_109160_2280.t126 524.808
R1160 a_109160_2280.n69 a_109160_2280.t144 524.808
R1161 a_109160_2280.n161 a_109160_2280.t164 508.743
R1162 a_109160_2280.n268 a_109160_2280.t184 508.743
R1163 a_109160_2280.n123 a_109160_2280.t161 508.743
R1164 a_109160_2280.n121 a_109160_2280.t156 508.743
R1165 a_109160_2280.n28 a_109160_2280.t153 499.442
R1166 a_109160_2280.n257 a_109160_2280.t132 499.442
R1167 a_109160_2280.n274 a_109160_2280.t176 499.442
R1168 a_109160_2280.n128 a_109160_2280.t167 499.442
R1169 a_109160_2280.n260 a_109160_2280.t190 475.976
R1170 a_109160_2280.n260 a_109160_2280.t179 475.976
R1171 a_109160_2280.n155 a_109160_2280.t159 475.976
R1172 a_109160_2280.n155 a_109160_2280.t187 475.976
R1173 a_109160_2280.n30 a_109160_2280.n3 337.098
R1174 a_109160_2280.n126 a_109160_2280.n125 337.098
R1175 a_109160_2280.n163 a_109160_2280.n162 296.158
R1176 a_109160_2280.n267 a_109160_2280.n266 296.158
R1177 a_109160_2280.n149 a_109160_2280.n16 296.158
R1178 a_109160_2280.n120 a_109160_2280.n119 296.158
R1179 a_109160_2280.n30 a_109160_2280.n29 292.5
R1180 a_109160_2280.n127 a_109160_2280.n126 292.5
R1181 a_109160_2280.n276 a_109160_2280.n275 292.5
R1182 a_109160_2280.n152 a_109160_2280.n151 292.5
R1183 a_109160_2280.n265 a_109160_2280.n264 292.5
R1184 a_109160_2280.n256 a_109160_2280.n255 292.5
R1185 a_109160_2280.t154 a_109160_2280.n30 239.517
R1186 a_109160_2280.n119 a_109160_2280.t157 239.517
R1187 a_109160_2280.n119 a_109160_2280.t174 239.517
R1188 a_109160_2280.t136 a_109160_2280.n149 239.517
R1189 a_109160_2280.n149 a_109160_2280.t162 239.517
R1190 a_109160_2280.n126 a_109160_2280.t168 239.517
R1191 a_109160_2280.t0 a_109160_2280.n284 205.381
R1192 a_109160_2280.n165 a_109160_2280.n164 197.133
R1193 a_109160_2280.n273 a_109160_2280.n272 197.133
R1194 a_109160_2280.n149 a_109160_2280.n148 197.133
R1195 a_109160_2280.n119 a_109160_2280.n118 197.133
R1196 a_109160_2280.t231 a_109160_2280.t154 195.161
R1197 a_109160_2280.t63 a_109160_2280.t231 195.161
R1198 a_109160_2280.t15 a_109160_2280.t63 195.161
R1199 a_109160_2280.t88 a_109160_2280.t15 195.161
R1200 a_109160_2280.t222 a_109160_2280.t88 195.161
R1201 a_109160_2280.t37 a_109160_2280.t222 195.161
R1202 a_109160_2280.t12 a_109160_2280.t37 195.161
R1203 a_109160_2280.t48 a_109160_2280.t12 195.161
R1204 a_109160_2280.t29 a_109160_2280.t48 195.161
R1205 a_109160_2280.t232 a_109160_2280.t29 195.161
R1206 a_109160_2280.t157 a_109160_2280.t232 195.161
R1207 a_109160_2280.t174 a_109160_2280.t22 195.161
R1208 a_109160_2280.t61 a_109160_2280.t136 195.161
R1209 a_109160_2280.t17 a_109160_2280.t162 195.161
R1210 a_109160_2280.t59 a_109160_2280.t17 195.161
R1211 a_109160_2280.t226 a_109160_2280.t59 195.161
R1212 a_109160_2280.t7 a_109160_2280.t226 195.161
R1213 a_109160_2280.t11 a_109160_2280.t7 195.161
R1214 a_109160_2280.t58 a_109160_2280.t11 195.161
R1215 a_109160_2280.t230 a_109160_2280.t58 195.161
R1216 a_109160_2280.t76 a_109160_2280.t230 195.161
R1217 a_109160_2280.t49 a_109160_2280.t76 195.161
R1218 a_109160_2280.t75 a_109160_2280.t49 195.161
R1219 a_109160_2280.t168 a_109160_2280.t75 195.161
R1220 a_109160_2280.n261 a_109160_2280.n260 161.3
R1221 a_109160_2280.n156 a_109160_2280.n155 161.3
R1222 a_109160_2280.n202 a_109160_2280.n0 148.017
R1223 a_109160_2280.n254 a_109160_2280.n253 148.017
R1224 a_109160_2280.n278 a_109160_2280.n277 148.017
R1225 a_109160_2280.n284 a_109160_2280.n283 148.017
R1226 a_109160_2280.n210 a_109160_2280.n208 121.251
R1227 a_109160_2280.n104 a_109160_2280.n103 121.136
R1228 a_109160_2280.n102 a_109160_2280.n101 121.136
R1229 a_109160_2280.n100 a_109160_2280.n99 121.136
R1230 a_109160_2280.n98 a_109160_2280.n97 121.136
R1231 a_109160_2280.n96 a_109160_2280.n95 121.136
R1232 a_109160_2280.n94 a_109160_2280.n93 121.136
R1233 a_109160_2280.n218 a_109160_2280.n217 121.136
R1234 a_109160_2280.n216 a_109160_2280.n215 121.136
R1235 a_109160_2280.n214 a_109160_2280.n213 121.136
R1236 a_109160_2280.n212 a_109160_2280.n211 121.136
R1237 a_109160_2280.n210 a_109160_2280.n209 121.136
R1238 a_109160_2280.n150 a_109160_2280.t22 97.5812
R1239 a_109160_2280.n150 a_109160_2280.t61 97.5812
R1240 a_109160_2280.n276 a_109160_2280.t177 93.9878
R1241 a_109160_2280.n255 a_109160_2280.t133 93.9878
R1242 a_109160_2280.n289 a_109160_2280.t44 91.9344
R1243 a_109160_2280.t73 a_109160_2280.t82 83.5448
R1244 a_109160_2280.t103 a_109160_2280.t93 76.5828
R1245 a_109160_2280.t106 a_109160_2280.t98 76.5828
R1246 a_109160_2280.t101 a_109160_2280.t94 76.5828
R1247 a_109160_2280.t99 a_109160_2280.t109 76.5828
R1248 a_109160_2280.t96 a_109160_2280.t107 76.5828
R1249 a_109160_2280.t177 a_109160_2280.t200 76.5828
R1250 a_109160_2280.t200 a_109160_2280.t204 76.5828
R1251 a_109160_2280.t204 a_109160_2280.t198 76.5828
R1252 a_109160_2280.t227 a_109160_2280.t5 76.5828
R1253 a_109160_2280.t5 a_109160_2280.t18 76.5828
R1254 a_109160_2280.t77 a_109160_2280.t1 76.5828
R1255 a_109160_2280.t212 a_109160_2280.t217 76.5828
R1256 a_109160_2280.t217 a_109160_2280.t133 76.5828
R1257 a_109160_2280.t221 a_109160_2280.t10 76.5828
R1258 a_109160_2280.t31 a_109160_2280.t45 76.5828
R1259 a_109160_2280.t38 a_109160_2280.t32 76.5828
R1260 a_109160_2280.t33 a_109160_2280.t60 76.5828
R1261 a_109160_2280.t46 a_109160_2280.t229 76.5828
R1262 a_109160_2280.t145 a_109160_2280.t171 73.1018
R1263 a_109160_2280.t182 a_109160_2280.t127 73.1018
R1264 a_109160_2280.n266 a_109160_2280.t34 73.1018
R1265 a_109160_2280.t151 a_109160_2280.t139 73.1018
R1266 a_109160_2280.t142 a_109160_2280.t130 73.1018
R1267 a_109160_2280.t13 a_109160_2280.t72 69.6207
R1268 a_109160_2280.t9 a_109160_2280.t0 69.6207
R1269 a_109160_2280.n29 a_109160_2280.t155 62.2505
R1270 a_109160_2280.n162 a_109160_2280.t166 62.2505
R1271 a_109160_2280.n267 a_109160_2280.t186 62.2505
R1272 a_109160_2280.n263 a_109160_2280.t192 62.2505
R1273 a_109160_2280.n14 a_109160_2280.t180 62.2505
R1274 a_109160_2280.n153 a_109160_2280.t160 62.2505
R1275 a_109160_2280.n15 a_109160_2280.t189 62.2505
R1276 a_109160_2280.n256 a_109160_2280.t134 62.2505
R1277 a_109160_2280.n275 a_109160_2280.t178 62.2505
R1278 a_109160_2280.n16 a_109160_2280.t163 62.2505
R1279 a_109160_2280.n120 a_109160_2280.t158 62.2505
R1280 a_109160_2280.n127 a_109160_2280.t169 62.2505
R1281 a_109160_2280.n238 a_109160_2280.n237 59.2425
R1282 a_109160_2280.n251 a_109160_2280.n250 59.2425
R1283 a_109160_2280.n10 a_109160_2280.n7 59.2425
R1284 a_109160_2280.n68 a_109160_2280.n4 59.2425
R1285 a_109160_2280.t122 a_109160_2280.t103 59.1777
R1286 a_109160_2280.t107 a_109160_2280.t114 59.1777
R1287 a_109160_2280.n273 a_109160_2280.t205 59.1777
R1288 a_109160_2280.n265 a_109160_2280.t54 59.1777
R1289 a_109160_2280.n164 a_109160_2280.t218 59.1777
R1290 a_109160_2280.t120 a_109160_2280.t221 59.1777
R1291 a_109160_2280.t229 a_109160_2280.t118 59.1777
R1292 a_109160_2280.t171 a_109160_2280.n4 52.2157
R1293 a_109160_2280.n7 a_109160_2280.t182 52.2157
R1294 a_109160_2280.n251 a_109160_2280.t139 52.2157
R1295 a_109160_2280.n237 a_109160_2280.t142 52.2157
R1296 a_109160_2280.t14 a_109160_2280.t65 49.6021
R1297 a_109160_2280.t112 a_109160_2280.t106 45.2537
R1298 a_109160_2280.t109 a_109160_2280.t124 45.2537
R1299 a_109160_2280.t43 a_109160_2280.t223 45.2537
R1300 a_109160_2280.t116 a_109160_2280.t31 45.2537
R1301 a_109160_2280.t60 a_109160_2280.t110 45.2537
R1302 a_109160_2280.t44 a_109160_2280.t24 42.7605
R1303 a_109160_2280.t70 a_109160_2280.t85 42.7605
R1304 a_109160_2280.n284 a_109160_2280.n4 41.7727
R1305 a_109160_2280.n277 a_109160_2280.n7 41.7727
R1306 a_109160_2280.t199 a_109160_2280.t148 41.7727
R1307 a_109160_2280.t203 a_109160_2280.t50 41.7727
R1308 a_109160_2280.t197 a_109160_2280.t56 41.7727
R1309 a_109160_2280.t202 a_109160_2280.t83 41.7727
R1310 a_109160_2280.t206 a_109160_2280.t66 41.7727
R1311 a_109160_2280.t201 a_109160_2280.t52 41.7727
R1312 a_109160_2280.t188 a_109160_2280.t20 41.7727
R1313 a_109160_2280.t234 a_109160_2280.t191 41.7727
R1314 a_109160_2280.t86 a_109160_2280.t215 41.7727
R1315 a_109160_2280.t25 a_109160_2280.t220 41.7727
R1316 a_109160_2280.t79 a_109160_2280.t214 41.7727
R1317 a_109160_2280.t3 a_109160_2280.t211 41.7727
R1318 a_109160_2280.t68 a_109160_2280.t216 41.7727
R1319 a_109160_2280.t39 a_109160_2280.t219 41.7727
R1320 a_109160_2280.t194 a_109160_2280.t213 41.7727
R1321 a_109160_2280.n254 a_109160_2280.n251 41.7727
R1322 a_109160_2280.n237 a_109160_2280.n0 41.7727
R1323 a_109160_2280.n165 a_109160_2280.t196 40.4338
R1324 a_109160_2280.n272 a_109160_2280.t149 40.4338
R1325 a_109160_2280.n148 a_109160_2280.t137 40.4338
R1326 a_109160_2280.n118 a_109160_2280.t175 40.4338
R1327 a_109160_2280.t18 a_109160_2280.n150 38.2916
R1328 a_109160_2280.n150 a_109160_2280.t34 38.2916
R1329 a_109160_2280.n9 a_109160_2280.n8 37.5297
R1330 a_109160_2280.n167 a_109160_2280.n166 37.5297
R1331 a_109160_2280.n169 a_109160_2280.n168 37.5297
R1332 a_109160_2280.n171 a_109160_2280.n170 37.5297
R1333 a_109160_2280.n173 a_109160_2280.n172 37.5297
R1334 a_109160_2280.n175 a_109160_2280.n174 37.5297
R1335 a_109160_2280.n177 a_109160_2280.n176 37.5297
R1336 a_109160_2280.n179 a_109160_2280.n178 37.5297
R1337 a_109160_2280.n181 a_109160_2280.n180 37.5297
R1338 a_109160_2280.n183 a_109160_2280.n182 37.5297
R1339 a_109160_2280.n185 a_109160_2280.n184 37.5297
R1340 a_109160_2280.t148 a_109160_2280.t205 34.8106
R1341 a_109160_2280.t50 a_109160_2280.t199 34.8106
R1342 a_109160_2280.t56 a_109160_2280.t203 34.8106
R1343 a_109160_2280.t83 a_109160_2280.t197 34.8106
R1344 a_109160_2280.t66 a_109160_2280.t202 34.8106
R1345 a_109160_2280.t52 a_109160_2280.t206 34.8106
R1346 a_109160_2280.t20 a_109160_2280.t201 34.8106
R1347 a_109160_2280.t223 a_109160_2280.t188 34.8106
R1348 a_109160_2280.t219 a_109160_2280.t68 34.8106
R1349 a_109160_2280.t213 a_109160_2280.t39 34.8106
R1350 a_109160_2280.t218 a_109160_2280.t194 34.8106
R1351 a_109160_2280.n18 a_109160_2280.n17 34.5991
R1352 a_109160_2280.n257 a_109160_2280.n256 31.5738
R1353 a_109160_2280.t94 a_109160_2280.t112 31.3296
R1354 a_109160_2280.t124 a_109160_2280.t101 31.3296
R1355 a_109160_2280.n163 a_109160_2280.t3 31.3296
R1356 a_109160_2280.t32 a_109160_2280.t116 31.3296
R1357 a_109160_2280.t110 a_109160_2280.t38 31.3296
R1358 a_109160_2280.n202 a_109160_2280.t143 31.1255
R1359 a_109160_2280.n253 a_109160_2280.t140 31.1255
R1360 a_109160_2280.n278 a_109160_2280.t183 31.1255
R1361 a_109160_2280.n283 a_109160_2280.t172 31.1255
R1362 a_109160_2280.n275 a_109160_2280.n274 29.8672
R1363 a_109160_2280.n128 a_109160_2280.n127 29.8672
R1364 a_109160_2280.n29 a_109160_2280.n28 29.8672
R1365 a_109160_2280.n290 a_109160_2280.n0 27.8486
R1366 a_109160_2280.n290 a_109160_2280.n289 27.8486
R1367 a_109160_2280.t191 a_109160_2280.t30 20.8866
R1368 a_109160_2280.t215 a_109160_2280.t89 20.8866
R1369 a_109160_2280.t220 a_109160_2280.t16 20.8866
R1370 a_109160_2280.t214 a_109160_2280.t64 20.8866
R1371 a_109160_2280.t211 a_109160_2280.t165 20.8866
R1372 a_109160_2280.n103 a_109160_2280.t90 19.7005
R1373 a_109160_2280.n103 a_109160_2280.t210 19.7005
R1374 a_109160_2280.n101 a_109160_2280.t97 19.7005
R1375 a_109160_2280.n101 a_109160_2280.t105 19.7005
R1376 a_109160_2280.n99 a_109160_2280.t100 19.7005
R1377 a_109160_2280.n99 a_109160_2280.t108 19.7005
R1378 a_109160_2280.n97 a_109160_2280.t104 19.7005
R1379 a_109160_2280.n97 a_109160_2280.t91 19.7005
R1380 a_109160_2280.n95 a_109160_2280.t102 19.7005
R1381 a_109160_2280.n95 a_109160_2280.t95 19.7005
R1382 a_109160_2280.n93 a_109160_2280.t209 19.7005
R1383 a_109160_2280.n93 a_109160_2280.t92 19.7005
R1384 a_109160_2280.n217 a_109160_2280.t28 19.7005
R1385 a_109160_2280.n217 a_109160_2280.t208 19.7005
R1386 a_109160_2280.n215 a_109160_2280.t233 19.7005
R1387 a_109160_2280.n215 a_109160_2280.t41 19.7005
R1388 a_109160_2280.n213 a_109160_2280.t47 19.7005
R1389 a_109160_2280.n213 a_109160_2280.t225 19.7005
R1390 a_109160_2280.n211 a_109160_2280.t36 19.7005
R1391 a_109160_2280.n211 a_109160_2280.t74 19.7005
R1392 a_109160_2280.n209 a_109160_2280.t81 19.7005
R1393 a_109160_2280.n209 a_109160_2280.t27 19.7005
R1394 a_109160_2280.n208 a_109160_2280.t207 19.7005
R1395 a_109160_2280.n208 a_109160_2280.t42 19.7005
R1396 a_109160_2280.t98 a_109160_2280.t122 17.4056
R1397 a_109160_2280.t114 a_109160_2280.t99 17.4056
R1398 a_109160_2280.t198 a_109160_2280.n273 17.4056
R1399 a_109160_2280.n151 a_109160_2280.t227 17.4056
R1400 a_109160_2280.n164 a_109160_2280.t212 17.4056
R1401 a_109160_2280.t45 a_109160_2280.t120 17.4056
R1402 a_109160_2280.t118 a_109160_2280.t33 17.4056
R1403 a_109160_2280.t82 a_109160_2280.t13 13.9246
R1404 a_109160_2280.t72 a_109160_2280.t9 13.9246
R1405 a_109160_2280.n151 a_109160_2280.t43 13.9246
R1406 a_109160_2280.t1 a_109160_2280.t185 13.9246
R1407 a_109160_2280.t30 a_109160_2280.t54 13.9246
R1408 a_109160_2280.t89 a_109160_2280.t234 13.9246
R1409 a_109160_2280.t16 a_109160_2280.t86 13.9246
R1410 a_109160_2280.t64 a_109160_2280.t25 13.9246
R1411 a_109160_2280.t165 a_109160_2280.t79 13.9246
R1412 a_109160_2280.n238 a_109160_2280.t131 12.6791
R1413 a_109160_2280.n250 a_109160_2280.t152 12.6791
R1414 a_109160_2280.n10 a_109160_2280.t128 12.6791
R1415 a_109160_2280.n68 a_109160_2280.t146 12.6791
R1416 a_109160_2280.n61 a_109160_2280.n60 12.641
R1417 a_109160_2280.n247 a_109160_2280.n193 12.641
R1418 a_109160_2280.n242 a_109160_2280.n241 12.1114
R1419 a_109160_2280.n63 a_109160_2280.n62 12.1114
R1420 a_109160_2280.n258 a_109160_2280.n257 11.4533
R1421 a_109160_2280.n274 a_109160_2280.n6 11.4533
R1422 a_109160_2280.n129 a_109160_2280.n128 11.2033
R1423 a_109160_2280.n28 a_109160_2280.n27 11.2029
R1424 a_109160_2280.n8 a_109160_2280.t51 9.6005
R1425 a_109160_2280.n8 a_109160_2280.t57 9.6005
R1426 a_109160_2280.n166 a_109160_2280.t84 9.6005
R1427 a_109160_2280.n166 a_109160_2280.t67 9.6005
R1428 a_109160_2280.n168 a_109160_2280.t53 9.6005
R1429 a_109160_2280.n168 a_109160_2280.t21 9.6005
R1430 a_109160_2280.n170 a_109160_2280.t224 9.6005
R1431 a_109160_2280.n170 a_109160_2280.t228 9.6005
R1432 a_109160_2280.n172 a_109160_2280.t6 9.6005
R1433 a_109160_2280.n172 a_109160_2280.t19 9.6005
R1434 a_109160_2280.n174 a_109160_2280.t35 9.6005
R1435 a_109160_2280.n174 a_109160_2280.t78 9.6005
R1436 a_109160_2280.n176 a_109160_2280.t2 9.6005
R1437 a_109160_2280.n176 a_109160_2280.t55 9.6005
R1438 a_109160_2280.n178 a_109160_2280.t235 9.6005
R1439 a_109160_2280.n178 a_109160_2280.t87 9.6005
R1440 a_109160_2280.n180 a_109160_2280.t26 9.6005
R1441 a_109160_2280.n180 a_109160_2280.t80 9.6005
R1442 a_109160_2280.n182 a_109160_2280.t4 9.6005
R1443 a_109160_2280.n182 a_109160_2280.t69 9.6005
R1444 a_109160_2280.n184 a_109160_2280.t40 9.6005
R1445 a_109160_2280.n184 a_109160_2280.t195 9.6005
R1446 a_109160_2280.n17 a_109160_2280.t23 9.6005
R1447 a_109160_2280.n17 a_109160_2280.t62 9.6005
R1448 a_109160_2280.t24 a_109160_2280.t70 8.55249
R1449 a_109160_2280.t85 a_109160_2280.t14 8.55249
R1450 a_109160_2280.n271 a_109160_2280.n9 5.063
R1451 a_109160_2280.n186 a_109160_2280.n185 4.71925
R1452 a_109160_2280.n74 a_109160_2280.n52 4.5005
R1453 a_109160_2280.n73 a_109160_2280.n72 4.5005
R1454 a_109160_2280.n74 a_109160_2280.n73 4.5005
R1455 a_109160_2280.n67 a_109160_2280.n56 4.5005
R1456 a_109160_2280.n66 a_109160_2280.n65 4.5005
R1457 a_109160_2280.n67 a_109160_2280.n66 4.5005
R1458 a_109160_2280.n246 a_109160_2280.n194 4.5005
R1459 a_109160_2280.n245 a_109160_2280.n244 4.5005
R1460 a_109160_2280.n246 a_109160_2280.n245 4.5005
R1461 a_109160_2280.n192 a_109160_2280.n191 4.5005
R1462 a_109160_2280.n191 a_109160_2280.n190 4.5005
R1463 a_109160_2280.n190 a_109160_2280.n188 4.5005
R1464 a_109160_2280.n223 a_109160_2280.n222 4.5005
R1465 a_109160_2280.n231 a_109160_2280.n199 4.5005
R1466 a_109160_2280.n229 a_109160_2280.n205 4.5005
R1467 a_109160_2280.n230 a_109160_2280.n201 4.5005
R1468 a_109160_2280.n230 a_109160_2280.n229 4.5005
R1469 a_109160_2280.n85 a_109160_2280.n50 4.5005
R1470 a_109160_2280.n81 a_109160_2280.n75 4.5005
R1471 a_109160_2280.n81 a_109160_2280.n80 4.5005
R1472 a_109160_2280.n80 a_109160_2280.n76 4.5005
R1473 a_109160_2280.n90 a_109160_2280.n88 4.5005
R1474 a_109160_2280.n92 a_109160_2280.n91 4.5005
R1475 a_109160_2280.n91 a_109160_2280.n90 4.5005
R1476 a_109160_2280.n24 a_109160_2280.n23 4.5005
R1477 a_109160_2280.n145 a_109160_2280.n19 4.5005
R1478 a_109160_2280.n144 a_109160_2280.n143 4.5005
R1479 a_109160_2280.n145 a_109160_2280.n144 4.5005
R1480 a_109160_2280.n33 a_109160_2280.n32 4.5005
R1481 a_109160_2280.n36 a_109160_2280.n35 4.5005
R1482 a_109160_2280.n41 a_109160_2280.n38 4.5005
R1483 a_109160_2280.n43 a_109160_2280.n42 4.5005
R1484 a_109160_2280.n42 a_109160_2280.n41 4.5005
R1485 a_109160_2280.n135 a_109160_2280.n26 4.5005
R1486 a_109160_2280.n135 a_109160_2280.n134 4.5005
R1487 a_109160_2280.n134 a_109160_2280.n130 4.5005
R1488 a_109160_2280.n271 a_109160_2280.n270 3.85122
R1489 a_109160_2280.n264 a_109160_2280.n14 3.65764
R1490 a_109160_2280.n264 a_109160_2280.n263 3.65764
R1491 a_109160_2280.n152 a_109160_2280.n15 3.65764
R1492 a_109160_2280.n153 a_109160_2280.n152 3.65764
R1493 a_109160_2280.t93 a_109160_2280.t145 3.48151
R1494 a_109160_2280.t127 a_109160_2280.t96 3.48151
R1495 a_109160_2280.n266 a_109160_2280.t77 3.48151
R1496 a_109160_2280.t185 a_109160_2280.n265 3.48151
R1497 a_109160_2280.t216 a_109160_2280.n163 3.48151
R1498 a_109160_2280.t10 a_109160_2280.t151 3.48151
R1499 a_109160_2280.t130 a_109160_2280.t46 3.48151
R1500 a_109160_2280.n241 a_109160_2280.t111 3.42907
R1501 a_109160_2280.n241 a_109160_2280.t119 3.42907
R1502 a_109160_2280.n193 a_109160_2280.t121 3.42907
R1503 a_109160_2280.n193 a_109160_2280.t117 3.42907
R1504 a_109160_2280.n60 a_109160_2280.t125 3.42907
R1505 a_109160_2280.n60 a_109160_2280.t115 3.42907
R1506 a_109160_2280.n62 a_109160_2280.t123 3.42907
R1507 a_109160_2280.n62 a_109160_2280.t113 3.42907
R1508 a_109160_2280.n162 a_109160_2280.n161 3.39217
R1509 a_109160_2280.n268 a_109160_2280.n267 3.39217
R1510 a_109160_2280.n123 a_109160_2280.n16 3.39217
R1511 a_109160_2280.n121 a_109160_2280.n120 3.39217
R1512 a_109160_2280.n262 a_109160_2280.n14 3.13621
R1513 a_109160_2280.n263 a_109160_2280.n262 3.13621
R1514 a_109160_2280.n154 a_109160_2280.n15 3.13621
R1515 a_109160_2280.n154 a_109160_2280.n153 3.13621
R1516 a_109160_2280.n240 a_109160_2280.n239 2.38247
R1517 a_109160_2280.n249 a_109160_2280.n248 2.38247
R1518 a_109160_2280.n12 a_109160_2280.n11 2.38247
R1519 a_109160_2280.n70 a_109160_2280.n69 2.38247
R1520 a_109160_2280.n204 a_109160_2280.n203 2.29914
R1521 a_109160_2280.n252 a_109160_2280.n158 2.29914
R1522 a_109160_2280.n280 a_109160_2280.n279 2.29914
R1523 a_109160_2280.n282 a_109160_2280.n281 2.29914
R1524 a_109160_2280.n189 a_109160_2280.n160 2.26187
R1525 a_109160_2280.n232 a_109160_2280.n198 2.26187
R1526 a_109160_2280.n84 a_109160_2280.n49 2.26187
R1527 a_109160_2280.n79 a_109160_2280.n77 2.26187
R1528 a_109160_2280.n136 a_109160_2280.n22 2.26187
R1529 a_109160_2280.n113 a_109160_2280.n112 2.26187
R1530 a_109160_2280.n133 a_109160_2280.n131 2.26187
R1531 a_109160_2280.n233 a_109160_2280.n232 2.26187
R1532 a_109160_2280.n71 a_109160_2280.n53 2.26187
R1533 a_109160_2280.n220 a_109160_2280.n207 2.26187
R1534 a_109160_2280.n221 a_109160_2280.n220 2.26187
R1535 a_109160_2280.n109 a_109160_2280.n108 2.26187
R1536 a_109160_2280.n89 a_109160_2280.n47 2.26187
R1537 a_109160_2280.n139 a_109160_2280.n138 2.26187
R1538 a_109160_2280.n142 a_109160_2280.n20 2.26187
R1539 a_109160_2280.n114 a_109160_2280.n113 2.26187
R1540 a_109160_2280.n65 a_109160_2280.n64 2.24241
R1541 a_109160_2280.n59 a_109160_2280.n58 2.24241
R1542 a_109160_2280.n244 a_109160_2280.n243 2.24241
R1543 a_109160_2280.n197 a_109160_2280.n196 2.24241
R1544 a_109160_2280.n72 a_109160_2280.n71 2.24063
R1545 a_109160_2280.n55 a_109160_2280.n54 2.24063
R1546 a_109160_2280.n192 a_109160_2280.n160 2.24063
R1547 a_109160_2280.n187 a_109160_2280.n159 2.24063
R1548 a_109160_2280.n224 a_109160_2280.n219 2.24063
R1549 a_109160_2280.n225 a_109160_2280.n207 2.24063
R1550 a_109160_2280.n236 a_109160_2280.n198 2.24063
R1551 a_109160_2280.n226 a_109160_2280.n201 2.24063
R1552 a_109160_2280.n206 a_109160_2280.n200 2.24063
R1553 a_109160_2280.n83 a_109160_2280.n82 2.24063
R1554 a_109160_2280.n77 a_109160_2280.n75 2.24063
R1555 a_109160_2280.n78 a_109160_2280.n51 2.24063
R1556 a_109160_2280.n92 a_109160_2280.n47 2.24063
R1557 a_109160_2280.n48 a_109160_2280.n46 2.24063
R1558 a_109160_2280.n138 a_109160_2280.n137 2.24063
R1559 a_109160_2280.n143 a_109160_2280.n142 2.24063
R1560 a_109160_2280.n141 a_109160_2280.n21 2.24063
R1561 a_109160_2280.n111 a_109160_2280.n31 2.24063
R1562 a_109160_2280.n106 a_109160_2280.n105 2.24063
R1563 a_109160_2280.n108 a_109160_2280.n107 2.24063
R1564 a_109160_2280.n44 a_109160_2280.n43 2.24063
R1565 a_109160_2280.n40 a_109160_2280.n39 2.24063
R1566 a_109160_2280.n131 a_109160_2280.n26 2.24063
R1567 a_109160_2280.n132 a_109160_2280.n25 2.24063
R1568 a_109160_2280.n63 a_109160_2280.n57 2.24063
R1569 a_109160_2280.n242 a_109160_2280.n195 2.24063
R1570 a_109160_2280.n235 a_109160_2280.n234 2.24063
R1571 a_109160_2280.n228 a_109160_2280.n227 2.24063
R1572 a_109160_2280.n87 a_109160_2280.n49 2.24063
R1573 a_109160_2280.n86 a_109160_2280.n5 2.24063
R1574 a_109160_2280.n140 a_109160_2280.n22 2.24063
R1575 a_109160_2280.n115 a_109160_2280.n114 2.24063
R1576 a_109160_2280.n110 a_109160_2280.n34 2.24063
R1577 a_109160_2280.n45 a_109160_2280.n37 2.24063
R1578 a_109160_2280.n191 a_109160_2280.n186 2.24008
R1579 a_109160_2280.n272 a_109160_2280.n271 2.19633
R1580 a_109160_2280.n148 a_109160_2280.n147 2.19633
R1581 a_109160_2280.n118 a_109160_2280.n117 2.19633
R1582 a_109160_2280.n261 a_109160_2280.n259 2.15331
R1583 a_109160_2280.n157 a_109160_2280.n156 2.15331
R1584 a_109160_2280.n239 a_109160_2280.n238 2.09414
R1585 a_109160_2280.n250 a_109160_2280.n249 2.09414
R1586 a_109160_2280.n11 a_109160_2280.n10 2.09414
R1587 a_109160_2280.n69 a_109160_2280.n68 2.09414
R1588 a_109160_2280.n161 a_109160_2280.n13 2.00747
R1589 a_109160_2280.n269 a_109160_2280.n268 2.00747
R1590 a_109160_2280.n203 a_109160_2280.n202 1.93383
R1591 a_109160_2280.n253 a_109160_2280.n252 1.93383
R1592 a_109160_2280.n279 a_109160_2280.n278 1.93383
R1593 a_109160_2280.n283 a_109160_2280.n282 1.93383
R1594 a_109160_2280.n186 a_109160_2280.n165 1.91062
R1595 a_109160_2280.n124 a_109160_2280.n123 1.90331
R1596 a_109160_2280.n122 a_109160_2280.n121 1.90331
R1597 a_109160_2280.t65 a_109160_2280.t71 1.7109
R1598 a_109160_2280.n117 a_109160_2280.n116 1.56997
R1599 a_109160_2280.n147 a_109160_2280.n146 1.56997
R1600 a_109160_2280.n234 a_109160_2280.n230 1.5005
R1601 a_109160_2280.n83 a_109160_2280.n81 1.5005
R1602 a_109160_2280.n227 a_109160_2280.n225 1.07342
R1603 a_109160_2280.n91 a_109160_2280.n87 1.07342
R1604 a_109160_2280.n270 a_109160_2280.n12 1.07324
R1605 a_109160_2280.n116 a_109160_2280.n115 1.063
R1606 a_109160_2280.n146 a_109160_2280.n145 1.063
R1607 a_109160_2280.n248 a_109160_2280.n192 0.930936
R1608 a_109160_2280.n219 a_109160_2280.n218 0.786958
R1609 a_109160_2280.n94 a_109160_2280.n92 0.786958
R1610 a_109160_2280.n280 a_109160_2280.n6 0.78175
R1611 a_109160_2280.n258 a_109160_2280.n158 0.78175
R1612 a_109160_2280.n240 a_109160_2280.n236 0.764269
R1613 a_109160_2280.n270 a_109160_2280.n269 0.759061
R1614 a_109160_2280.n281 a_109160_2280.n5 0.729667
R1615 a_109160_2280.n157 a_109160_2280.n6 0.729667
R1616 a_109160_2280.n259 a_109160_2280.n258 0.729667
R1617 a_109160_2280.n229 a_109160_2280.n204 0.729667
R1618 a_109160_2280.n281 a_109160_2280.n280 0.688
R1619 a_109160_2280.n204 a_109160_2280.n158 0.688
R1620 a_109160_2280.n122 a_109160_2280.n27 0.688
R1621 a_109160_2280.n129 a_109160_2280.n124 0.688
R1622 a_109160_2280.n185 a_109160_2280.n183 0.563
R1623 a_109160_2280.n183 a_109160_2280.n181 0.563
R1624 a_109160_2280.n181 a_109160_2280.n179 0.563
R1625 a_109160_2280.n179 a_109160_2280.n177 0.563
R1626 a_109160_2280.n177 a_109160_2280.n175 0.563
R1627 a_109160_2280.n175 a_109160_2280.n173 0.563
R1628 a_109160_2280.n173 a_109160_2280.n171 0.563
R1629 a_109160_2280.n171 a_109160_2280.n169 0.563
R1630 a_109160_2280.n169 a_109160_2280.n167 0.563
R1631 a_109160_2280.n167 a_109160_2280.n9 0.563
R1632 a_109160_2280.n105 a_109160_2280.n104 0.464042
R1633 a_109160_2280.n75 a_109160_2280.n74 0.408426
R1634 a_109160_2280.n124 a_109160_2280.n122 0.396333
R1635 a_109160_2280.n269 a_109160_2280.n13 0.345926
R1636 a_109160_2280.n137 a_109160_2280.n135 0.34425
R1637 a_109160_2280.n107 a_109160_2280.n45 0.34425
R1638 a_109160_2280.n65 a_109160_2280.n61 0.322473
R1639 a_109160_2280.n247 a_109160_2280.n246 0.322025
R1640 a_109160_2280.n259 a_109160_2280.n157 0.313
R1641 a_109160_2280.n43 a_109160_2280.n27 0.292167
R1642 a_109160_2280.n134 a_109160_2280.n129 0.292167
R1643 a_109160_2280.n72 a_109160_2280.n70 0.271333
R1644 a_109160_2280.n190 a_109160_2280.n13 0.21925
R1645 a_109160_2280.n262 a_109160_2280.n261 0.208833
R1646 a_109160_2280.n156 a_109160_2280.n154 0.208833
R1647 a_109160_2280.n144 a_109160_2280.n140 0.172375
R1648 a_109160_2280.n111 a_109160_2280.n110 0.172375
R1649 a_109160_2280.n61 a_109160_2280.n12 0.128173
R1650 a_109160_2280.n248 a_109160_2280.n247 0.126673
R1651 a_109160_2280.n212 a_109160_2280.n210 0.115083
R1652 a_109160_2280.n214 a_109160_2280.n212 0.115083
R1653 a_109160_2280.n216 a_109160_2280.n214 0.115083
R1654 a_109160_2280.n218 a_109160_2280.n216 0.115083
R1655 a_109160_2280.n96 a_109160_2280.n94 0.115083
R1656 a_109160_2280.n98 a_109160_2280.n96 0.115083
R1657 a_109160_2280.n100 a_109160_2280.n98 0.115083
R1658 a_109160_2280.n102 a_109160_2280.n100 0.115083
R1659 a_109160_2280.n104 a_109160_2280.n102 0.115083
R1660 a_109160_2280.n116 a_109160_2280.n18 0.115083
R1661 a_109160_2280.n146 a_109160_2280.n18 0.115083
R1662 a_109160_2280.n70 a_109160_2280.n67 0.09425
R1663 a_109160_2280.n244 a_109160_2280.n240 0.09425
R1664 a_109160_2280.n78 a_109160_2280.n75 0.0421667
R1665 a_109160_2280.n72 a_109160_2280.n55 0.0421667
R1666 a_109160_2280.n65 a_109160_2280.n59 0.0421667
R1667 a_109160_2280.n192 a_109160_2280.n159 0.0421667
R1668 a_109160_2280.n244 a_109160_2280.n197 0.0421667
R1669 a_109160_2280.n206 a_109160_2280.n201 0.0421667
R1670 a_109160_2280.n92 a_109160_2280.n46 0.0421667
R1671 a_109160_2280.n143 a_109160_2280.n141 0.0421667
R1672 a_109160_2280.n43 a_109160_2280.n39 0.0421667
R1673 a_109160_2280.n132 a_109160_2280.n26 0.0421667
R1674 a_109160_2280.n188 a_109160_2280.n187 0.0217373
R1675 a_109160_2280.n188 a_109160_2280.n160 0.0217373
R1676 a_109160_2280.n73 a_109160_2280.n54 0.0217373
R1677 a_109160_2280.n79 a_109160_2280.n78 0.0217373
R1678 a_109160_2280.n189 a_109160_2280.n159 0.0217373
R1679 a_109160_2280.n71 a_109160_2280.n52 0.0217373
R1680 a_109160_2280.n54 a_109160_2280.n52 0.0217373
R1681 a_109160_2280.n191 a_109160_2280.n187 0.0217373
R1682 a_109160_2280.n190 a_109160_2280.n189 0.0217373
R1683 a_109160_2280.n224 a_109160_2280.n223 0.0217373
R1684 a_109160_2280.n227 a_109160_2280.n226 0.0217373
R1685 a_109160_2280.n230 a_109160_2280.n200 0.0217373
R1686 a_109160_2280.n231 a_109160_2280.n198 0.0217373
R1687 a_109160_2280.n222 a_109160_2280.n207 0.0217373
R1688 a_109160_2280.n225 a_109160_2280.n224 0.0217373
R1689 a_109160_2280.n232 a_109160_2280.n199 0.0217373
R1690 a_109160_2280.n82 a_109160_2280.n5 0.0217373
R1691 a_109160_2280.n226 a_109160_2280.n205 0.0217373
R1692 a_109160_2280.n205 a_109160_2280.n200 0.0217373
R1693 a_109160_2280.n91 a_109160_2280.n48 0.0217373
R1694 a_109160_2280.n85 a_109160_2280.n84 0.0217373
R1695 a_109160_2280.n76 a_109160_2280.n51 0.0217373
R1696 a_109160_2280.n77 a_109160_2280.n76 0.0217373
R1697 a_109160_2280.n82 a_109160_2280.n50 0.0217373
R1698 a_109160_2280.n84 a_109160_2280.n83 0.0217373
R1699 a_109160_2280.n81 a_109160_2280.n51 0.0217373
R1700 a_109160_2280.n80 a_109160_2280.n79 0.0217373
R1701 a_109160_2280.n88 a_109160_2280.n47 0.0217373
R1702 a_109160_2280.n88 a_109160_2280.n48 0.0217373
R1703 a_109160_2280.n144 a_109160_2280.n21 0.0217373
R1704 a_109160_2280.n136 a_109160_2280.n23 0.0217373
R1705 a_109160_2280.n130 a_109160_2280.n25 0.0217373
R1706 a_109160_2280.n131 a_109160_2280.n130 0.0217373
R1707 a_109160_2280.n138 a_109160_2280.n24 0.0217373
R1708 a_109160_2280.n137 a_109160_2280.n136 0.0217373
R1709 a_109160_2280.n115 a_109160_2280.n31 0.0217373
R1710 a_109160_2280.n142 a_109160_2280.n19 0.0217373
R1711 a_109160_2280.n21 a_109160_2280.n19 0.0217373
R1712 a_109160_2280.n112 a_109160_2280.n32 0.0217373
R1713 a_109160_2280.n106 a_109160_2280.n35 0.0217373
R1714 a_109160_2280.n45 a_109160_2280.n44 0.0217373
R1715 a_109160_2280.n42 a_109160_2280.n40 0.0217373
R1716 a_109160_2280.n33 a_109160_2280.n31 0.0217373
R1717 a_109160_2280.n112 a_109160_2280.n111 0.0217373
R1718 a_109160_2280.n108 a_109160_2280.n36 0.0217373
R1719 a_109160_2280.n107 a_109160_2280.n106 0.0217373
R1720 a_109160_2280.n133 a_109160_2280.n132 0.0217373
R1721 a_109160_2280.n44 a_109160_2280.n38 0.0217373
R1722 a_109160_2280.n40 a_109160_2280.n38 0.0217373
R1723 a_109160_2280.n135 a_109160_2280.n25 0.0217373
R1724 a_109160_2280.n134 a_109160_2280.n133 0.0217373
R1725 a_109160_2280.n74 a_109160_2280.n53 0.0217373
R1726 a_109160_2280.n67 a_109160_2280.n57 0.0217373
R1727 a_109160_2280.n246 a_109160_2280.n195 0.0217373
R1728 a_109160_2280.n235 a_109160_2280.n199 0.0217373
R1729 a_109160_2280.n55 a_109160_2280.n53 0.0217373
R1730 a_109160_2280.n59 a_109160_2280.n57 0.0217373
R1731 a_109160_2280.n197 a_109160_2280.n195 0.0217373
R1732 a_109160_2280.n222 a_109160_2280.n221 0.0217373
R1733 a_109160_2280.n223 a_109160_2280.n220 0.0217373
R1734 a_109160_2280.n233 a_109160_2280.n231 0.0217373
R1735 a_109160_2280.n221 a_109160_2280.n219 0.0217373
R1736 a_109160_2280.n234 a_109160_2280.n233 0.0217373
R1737 a_109160_2280.n236 a_109160_2280.n235 0.0217373
R1738 a_109160_2280.n50 a_109160_2280.n49 0.0217373
R1739 a_109160_2280.n229 a_109160_2280.n228 0.0217373
R1740 a_109160_2280.n228 a_109160_2280.n206 0.0217373
R1741 a_109160_2280.n86 a_109160_2280.n85 0.0217373
R1742 a_109160_2280.n87 a_109160_2280.n86 0.0217373
R1743 a_109160_2280.n90 a_109160_2280.n89 0.0217373
R1744 a_109160_2280.n36 a_109160_2280.n34 0.0217373
R1745 a_109160_2280.n89 a_109160_2280.n46 0.0217373
R1746 a_109160_2280.n24 a_109160_2280.n22 0.0217373
R1747 a_109160_2280.n139 a_109160_2280.n23 0.0217373
R1748 a_109160_2280.n140 a_109160_2280.n139 0.0217373
R1749 a_109160_2280.n113 a_109160_2280.n33 0.0217373
R1750 a_109160_2280.n145 a_109160_2280.n20 0.0217373
R1751 a_109160_2280.n141 a_109160_2280.n20 0.0217373
R1752 a_109160_2280.n114 a_109160_2280.n32 0.0217373
R1753 a_109160_2280.n109 a_109160_2280.n35 0.0217373
R1754 a_109160_2280.n110 a_109160_2280.n109 0.0217373
R1755 a_109160_2280.n105 a_109160_2280.n34 0.0217373
R1756 a_109160_2280.n41 a_109160_2280.n37 0.0217373
R1757 a_109160_2280.n39 a_109160_2280.n37 0.0217373
R1758 a_109160_2280.n243 a_109160_2280.n242 0.0181756
R1759 a_109160_2280.n245 a_109160_2280.n196 0.0181756
R1760 a_109160_2280.n64 a_109160_2280.n63 0.0181756
R1761 a_109160_2280.n66 a_109160_2280.n58 0.0181756
R1762 a_109160_2280.n64 a_109160_2280.n56 0.0181756
R1763 a_109160_2280.n58 a_109160_2280.n56 0.0181756
R1764 a_109160_2280.n243 a_109160_2280.n194 0.0181756
R1765 a_109160_2280.n196 a_109160_2280.n194 0.0181756
R1766 VOUT+.n27 VOUT+.t0 110.191
R1767 VOUT+.n51 VOUT+.n50 34.9935
R1768 VOUT+.n49 VOUT+.n48 34.9935
R1769 VOUT+.n63 VOUT+.n62 34.9935
R1770 VOUT+.n59 VOUT+.n58 34.9935
R1771 VOUT+.n56 VOUT+.n55 34.9935
R1772 VOUT+.n53 VOUT+.n52 34.9935
R1773 VOUT+.n10 VOUT+.n9 9.73997
R1774 VOUT+.n14 VOUT+.n13 9.73997
R1775 VOUT+.n17 VOUT+.n16 9.73997
R1776 VOUT+.n15 VOUT+.n14 6.64633
R1777 VOUT+.n15 VOUT+.n10 6.64633
R1778 VOUT+.n50 VOUT+.t2 6.56717
R1779 VOUT+.n50 VOUT+.t13 6.56717
R1780 VOUT+.n48 VOUT+.t12 6.56717
R1781 VOUT+.n48 VOUT+.t14 6.56717
R1782 VOUT+.n62 VOUT+.t16 6.56717
R1783 VOUT+.n62 VOUT+.t1 6.56717
R1784 VOUT+.n58 VOUT+.t15 6.56717
R1785 VOUT+.n58 VOUT+.t18 6.56717
R1786 VOUT+.n55 VOUT+.t5 6.56717
R1787 VOUT+.n55 VOUT+.t17 6.56717
R1788 VOUT+.n52 VOUT+.t4 6.56717
R1789 VOUT+.n52 VOUT+.t3 6.56717
R1790 VOUT+.n61 VOUT+.n49 6.3755
R1791 VOUT+.n54 VOUT+.n51 6.3755
R1792 VOUT+.n17 VOUT+.n15 6.02133
R1793 VOUT+.n63 VOUT+.n61 5.813
R1794 VOUT+.n60 VOUT+.n59 5.813
R1795 VOUT+.n57 VOUT+.n56 5.813
R1796 VOUT+.n54 VOUT+.n53 5.813
R1797 VOUT+.n64 VOUT+.n40 5.063
R1798 VOUT+.n67 VOUT+.n47 5.063
R1799 VOUT+.n134 VOUT+.t99 4.8295
R1800 VOUT+.n135 VOUT+.t132 4.8295
R1801 VOUT+.n136 VOUT+.t27 4.8295
R1802 VOUT+.n137 VOUT+.t79 4.8295
R1803 VOUT+.n138 VOUT+.t36 4.8295
R1804 VOUT+.n139 VOUT+.t85 4.8295
R1805 VOUT+.n149 VOUT+.t24 4.8295
R1806 VOUT+.n151 VOUT+.t94 4.8295
R1807 VOUT+.n152 VOUT+.t59 4.8295
R1808 VOUT+.n154 VOUT+.t62 4.8295
R1809 VOUT+.n155 VOUT+.t31 4.8295
R1810 VOUT+.n157 VOUT+.t20 4.8295
R1811 VOUT+.n158 VOUT+.t127 4.8295
R1812 VOUT+.n160 VOUT+.t119 4.8295
R1813 VOUT+.n161 VOUT+.t92 4.8295
R1814 VOUT+.n163 VOUT+.t152 4.8295
R1815 VOUT+.n164 VOUT+.t122 4.8295
R1816 VOUT+.n166 VOUT+.t113 4.8295
R1817 VOUT+.n167 VOUT+.t87 4.8295
R1818 VOUT+.n169 VOUT+.t78 4.8295
R1819 VOUT+.n170 VOUT+.t51 4.8295
R1820 VOUT+.n172 VOUT+.t106 4.8295
R1821 VOUT+.n173 VOUT+.t82 4.8295
R1822 VOUT+.n175 VOUT+.t72 4.8295
R1823 VOUT+.n176 VOUT+.t44 4.8295
R1824 VOUT+.n178 VOUT+.t35 4.8295
R1825 VOUT+.n179 VOUT+.t138 4.8295
R1826 VOUT+.n101 VOUT+.t141 4.8295
R1827 VOUT+.n114 VOUT+.t100 4.8295
R1828 VOUT+.n116 VOUT+.t33 4.8295
R1829 VOUT+.n117 VOUT+.t137 4.8295
R1830 VOUT+.n119 VOUT+.t95 4.8295
R1831 VOUT+.n120 VOUT+.t60 4.8295
R1832 VOUT+.n122 VOUT+.t55 4.8295
R1833 VOUT+.n123 VOUT+.t71 4.8295
R1834 VOUT+.n125 VOUT+.t154 4.8295
R1835 VOUT+.n126 VOUT+.t41 4.8295
R1836 VOUT+.n128 VOUT+.t125 4.8295
R1837 VOUT+.n129 VOUT+.t96 4.8295
R1838 VOUT+.n131 VOUT+.t26 4.8295
R1839 VOUT+.n132 VOUT+.t134 4.8295
R1840 VOUT+.n181 VOUT+.t38 4.8295
R1841 VOUT+.n141 VOUT+.t64 4.8154
R1842 VOUT+.n113 VOUT+.t57 4.806
R1843 VOUT+.n112 VOUT+.t42 4.806
R1844 VOUT+.n111 VOUT+.t74 4.806
R1845 VOUT+.n110 VOUT+.t108 4.806
R1846 VOUT+.n109 VOUT+.t147 4.806
R1847 VOUT+.n108 VOUT+.t126 4.806
R1848 VOUT+.n107 VOUT+.t103 4.806
R1849 VOUT+.n106 VOUT+.t145 4.806
R1850 VOUT+.n105 VOUT+.t123 4.806
R1851 VOUT+.n104 VOUT+.t21 4.806
R1852 VOUT+.n103 VOUT+.t61 4.806
R1853 VOUT+.n134 VOUT+.t128 4.5005
R1854 VOUT+.n135 VOUT+.t29 4.5005
R1855 VOUT+.n136 VOUT+.t66 4.5005
R1856 VOUT+.n137 VOUT+.t49 4.5005
R1857 VOUT+.n138 VOUT+.t22 4.5005
R1858 VOUT+.n139 VOUT+.t50 4.5005
R1859 VOUT+.n140 VOUT+.t143 4.5005
R1860 VOUT+.n141 VOUT+.t30 4.5005
R1861 VOUT+.n142 VOUT+.t130 4.5005
R1862 VOUT+.n143 VOUT+.t146 4.5005
R1863 VOUT+.n144 VOUT+.t34 4.5005
R1864 VOUT+.n145 VOUT+.t133 4.5005
R1865 VOUT+.n146 VOUT+.t97 4.5005
R1866 VOUT+.n147 VOUT+.t56 4.5005
R1867 VOUT+.n148 VOUT+.t81 4.5005
R1868 VOUT+.n150 VOUT+.t48 4.5005
R1869 VOUT+.n149 VOUT+.t140 4.5005
R1870 VOUT+.n151 VOUT+.t110 4.5005
R1871 VOUT+.n153 VOUT+.t77 4.5005
R1872 VOUT+.n152 VOUT+.t43 4.5005
R1873 VOUT+.n154 VOUT+.t148 4.5005
R1874 VOUT+.n156 VOUT+.t111 4.5005
R1875 VOUT+.n155 VOUT+.t83 4.5005
R1876 VOUT+.n157 VOUT+.t105 4.5005
R1877 VOUT+.n159 VOUT+.t75 4.5005
R1878 VOUT+.n158 VOUT+.t45 4.5005
R1879 VOUT+.n160 VOUT+.t70 4.5005
R1880 VOUT+.n162 VOUT+.t40 4.5005
R1881 VOUT+.n161 VOUT+.t139 4.5005
R1882 VOUT+.n163 VOUT+.t101 4.5005
R1883 VOUT+.n165 VOUT+.t69 4.5005
R1884 VOUT+.n164 VOUT+.t39 4.5005
R1885 VOUT+.n166 VOUT+.t65 4.5005
R1886 VOUT+.n168 VOUT+.t32 4.5005
R1887 VOUT+.n167 VOUT+.t135 4.5005
R1888 VOUT+.n169 VOUT+.t25 4.5005
R1889 VOUT+.n171 VOUT+.t131 4.5005
R1890 VOUT+.n170 VOUT+.t98 4.5005
R1891 VOUT+.n172 VOUT+.t58 4.5005
R1892 VOUT+.n174 VOUT+.t23 4.5005
R1893 VOUT+.n173 VOUT+.t129 4.5005
R1894 VOUT+.n175 VOUT+.t156 4.5005
R1895 VOUT+.n177 VOUT+.t124 4.5005
R1896 VOUT+.n176 VOUT+.t93 4.5005
R1897 VOUT+.n178 VOUT+.t118 4.5005
R1898 VOUT+.n180 VOUT+.t90 4.5005
R1899 VOUT+.n179 VOUT+.t53 4.5005
R1900 VOUT+.n102 VOUT+.t155 4.5005
R1901 VOUT+.n101 VOUT+.t120 4.5005
R1902 VOUT+.n103 VOUT+.t19 4.5005
R1903 VOUT+.n104 VOUT+.t121 4.5005
R1904 VOUT+.n105 VOUT+.t88 4.5005
R1905 VOUT+.n106 VOUT+.t102 4.5005
R1906 VOUT+.n107 VOUT+.t68 4.5005
R1907 VOUT+.n108 VOUT+.t91 4.5005
R1908 VOUT+.n109 VOUT+.t104 4.5005
R1909 VOUT+.n110 VOUT+.t73 4.5005
R1910 VOUT+.n111 VOUT+.t37 4.5005
R1911 VOUT+.n112 VOUT+.t136 4.5005
R1912 VOUT+.n113 VOUT+.t153 4.5005
R1913 VOUT+.n115 VOUT+.t116 4.5005
R1914 VOUT+.n114 VOUT+.t86 4.5005
R1915 VOUT+.n116 VOUT+.t54 4.5005
R1916 VOUT+.n118 VOUT+.t150 4.5005
R1917 VOUT+.n117 VOUT+.t115 4.5005
R1918 VOUT+.n119 VOUT+.t47 4.5005
R1919 VOUT+.n121 VOUT+.t144 4.5005
R1920 VOUT+.n120 VOUT+.t107 4.5005
R1921 VOUT+.n122 VOUT+.t149 4.5005
R1922 VOUT+.n124 VOUT+.t63 4.5005
R1923 VOUT+.n123 VOUT+.t109 4.5005
R1924 VOUT+.n125 VOUT+.t114 4.5005
R1925 VOUT+.n127 VOUT+.t28 4.5005
R1926 VOUT+.n126 VOUT+.t80 4.5005
R1927 VOUT+.n128 VOUT+.t76 4.5005
R1928 VOUT+.n130 VOUT+.t46 4.5005
R1929 VOUT+.n129 VOUT+.t142 4.5005
R1930 VOUT+.n131 VOUT+.t112 4.5005
R1931 VOUT+.n133 VOUT+.t84 4.5005
R1932 VOUT+.n132 VOUT+.t52 4.5005
R1933 VOUT+.n183 VOUT+.t151 4.5005
R1934 VOUT+.n182 VOUT+.t117 4.5005
R1935 VOUT+.n181 VOUT+.t89 4.5005
R1936 VOUT+.n184 VOUT+.t67 4.5005
R1937 VOUT+.n64 VOUT+.n41 4.5005
R1938 VOUT+.n65 VOUT+.n44 4.5005
R1939 VOUT+.n66 VOUT+.n45 4.5005
R1940 VOUT+.n68 VOUT+.n67 4.5005
R1941 VOUT+.n91 VOUT+.n90 4.5005
R1942 VOUT+.n87 VOUT+.n84 4.5005
R1943 VOUT+.n91 VOUT+.n84 4.5005
R1944 VOUT+.n92 VOUT+.n36 4.5005
R1945 VOUT+.n92 VOUT+.n38 4.5005
R1946 VOUT+.n92 VOUT+.n91 4.5005
R1947 VOUT+.n189 VOUT+.n95 4.5005
R1948 VOUT+.n190 VOUT+.n189 4.5005
R1949 VOUT+.n190 VOUT+.n32 4.5005
R1950 VOUT+.n191 VOUT+.n31 4.5005
R1951 VOUT+.n191 VOUT+.n190 4.5005
R1952 VOUT+.n192 VOUT+.n6 4.5005
R1953 VOUT+.n195 VOUT+.n6 4.5005
R1954 VOUT+ VOUT+.n195 4.5005
R1955 VOUT+.n195 VOUT+.n7 4.5005
R1956 VOUT+.n195 VOUT+.n194 4.5005
R1957 VOUT+ VOUT+.n0 4.5005
R1958 VOUT+.n7 VOUT+.n0 4.5005
R1959 VOUT+.n194 VOUT+.n0 4.5005
R1960 VOUT+.n9 VOUT+.t8 3.42907
R1961 VOUT+.n9 VOUT+.t10 3.42907
R1962 VOUT+.n13 VOUT+.t11 3.42907
R1963 VOUT+.n13 VOUT+.t9 3.42907
R1964 VOUT+.n16 VOUT+.t7 3.42907
R1965 VOUT+.n16 VOUT+.t6 3.42907
R1966 VOUT+.n89 VOUT+.n37 2.26725
R1967 VOUT+.n85 VOUT+.n35 2.24601
R1968 VOUT+.n3 VOUT+.n2 2.24601
R1969 VOUT+.n28 VOUT+.n4 2.24601
R1970 VOUT+.n188 VOUT+.n187 2.24477
R1971 VOUT+.n34 VOUT+.n29 2.24477
R1972 VOUT+.n92 VOUT+.n37 2.24063
R1973 VOUT+.n191 VOUT+.n30 2.24063
R1974 VOUT+.n5 VOUT+.n0 2.24063
R1975 VOUT+.n84 VOUT+.n83 2.24063
R1976 VOUT+.n189 VOUT+.n93 2.24063
R1977 VOUT+.n94 VOUT+.n32 2.24063
R1978 VOUT+.n192 VOUT+.n1 2.24063
R1979 VOUT+.n193 VOUT+.n192 2.24063
R1980 VOUT+.n90 VOUT+.n88 2.23934
R1981 VOUT+.n90 VOUT+.n86 2.23934
R1982 VOUT+.n14 VOUT+.n12 1.62886
R1983 VOUT+.n18 VOUT+.n17 1.52133
R1984 VOUT+.n25 VOUT+.n10 1.52133
R1985 VOUT+.n82 VOUT+.n81 1.5005
R1986 VOUT+.n80 VOUT+.n39 1.5005
R1987 VOUT+.n79 VOUT+.n78 1.5005
R1988 VOUT+.n77 VOUT+.n42 1.5005
R1989 VOUT+.n76 VOUT+.n75 1.5005
R1990 VOUT+.n74 VOUT+.n43 1.5005
R1991 VOUT+.n73 VOUT+.n72 1.5005
R1992 VOUT+.n71 VOUT+.n46 1.5005
R1993 VOUT+.n26 VOUT+.n25 1.5005
R1994 VOUT+.n24 VOUT+.n8 1.5005
R1995 VOUT+.n23 VOUT+.n22 1.5005
R1996 VOUT+.n21 VOUT+.n11 1.5005
R1997 VOUT+.n20 VOUT+.n19 1.5005
R1998 VOUT+.n68 VOUT+.n63 1.313
R1999 VOUT+.n59 VOUT+.n45 1.313
R2000 VOUT+.n56 VOUT+.n44 1.313
R2001 VOUT+.n53 VOUT+.n41 1.313
R2002 VOUT+.n49 VOUT+.n47 1.313
R2003 VOUT+.n51 VOUT+.n40 1.313
R2004 VOUT+.n190 VOUT+.n33 1.1455
R2005 VOUT+.n99 VOUT+.n98 1.13717
R2006 VOUT+.n100 VOUT+.n96 1.13717
R2007 VOUT+.n186 VOUT+.n185 1.13717
R2008 VOUT+.n97 VOUT+.n34 1.13717
R2009 VOUT+.n98 VOUT+.n31 1.13717
R2010 VOUT+.n96 VOUT+.n95 1.13717
R2011 VOUT+.n187 VOUT+.n186 1.13717
R2012 VOUT+.n70 VOUT+.n47 0.715216
R2013 VOUT+.n69 VOUT+.n68 0.65675
R2014 VOUT+.n73 VOUT+.n45 0.65675
R2015 VOUT+.n75 VOUT+.n44 0.65675
R2016 VOUT+.n79 VOUT+.n41 0.65675
R2017 VOUT+.n81 VOUT+.n40 0.65675
R2018 VOUT+.n99 VOUT+.n33 0.585
R2019 VOUT+.n192 VOUT+.n191 0.5705
R2020 VOUT+.n71 VOUT+.n70 0.564601
R2021 VOUT+.n65 VOUT+.n64 0.563
R2022 VOUT+.n66 VOUT+.n65 0.563
R2023 VOUT+.n67 VOUT+.n66 0.563
R2024 VOUT+.n61 VOUT+.n60 0.563
R2025 VOUT+.n60 VOUT+.n57 0.563
R2026 VOUT+.n57 VOUT+.n54 0.563
R2027 VOUT+.n91 VOUT+.n82 0.495292
R2028 VOUT+.n27 VOUT+.n26 0.380708
R2029 VOUT+.n140 VOUT+.n139 0.3295
R2030 VOUT+.n141 VOUT+.n140 0.3295
R2031 VOUT+.n142 VOUT+.n141 0.3295
R2032 VOUT+.n143 VOUT+.n142 0.3295
R2033 VOUT+.n144 VOUT+.n143 0.3295
R2034 VOUT+.n145 VOUT+.n144 0.3295
R2035 VOUT+.n146 VOUT+.n145 0.3295
R2036 VOUT+.n147 VOUT+.n146 0.3295
R2037 VOUT+.n148 VOUT+.n147 0.3295
R2038 VOUT+.n150 VOUT+.n148 0.3295
R2039 VOUT+.n150 VOUT+.n149 0.3295
R2040 VOUT+.n153 VOUT+.n151 0.3295
R2041 VOUT+.n153 VOUT+.n152 0.3295
R2042 VOUT+.n156 VOUT+.n154 0.3295
R2043 VOUT+.n156 VOUT+.n155 0.3295
R2044 VOUT+.n159 VOUT+.n157 0.3295
R2045 VOUT+.n159 VOUT+.n158 0.3295
R2046 VOUT+.n162 VOUT+.n160 0.3295
R2047 VOUT+.n162 VOUT+.n161 0.3295
R2048 VOUT+.n165 VOUT+.n163 0.3295
R2049 VOUT+.n165 VOUT+.n164 0.3295
R2050 VOUT+.n168 VOUT+.n166 0.3295
R2051 VOUT+.n168 VOUT+.n167 0.3295
R2052 VOUT+.n171 VOUT+.n169 0.3295
R2053 VOUT+.n171 VOUT+.n170 0.3295
R2054 VOUT+.n174 VOUT+.n172 0.3295
R2055 VOUT+.n174 VOUT+.n173 0.3295
R2056 VOUT+.n177 VOUT+.n175 0.3295
R2057 VOUT+.n177 VOUT+.n176 0.3295
R2058 VOUT+.n180 VOUT+.n178 0.3295
R2059 VOUT+.n180 VOUT+.n179 0.3295
R2060 VOUT+.n102 VOUT+.n101 0.3295
R2061 VOUT+.n104 VOUT+.n103 0.3295
R2062 VOUT+.n105 VOUT+.n104 0.3295
R2063 VOUT+.n106 VOUT+.n105 0.3295
R2064 VOUT+.n107 VOUT+.n106 0.3295
R2065 VOUT+.n108 VOUT+.n107 0.3295
R2066 VOUT+.n109 VOUT+.n108 0.3295
R2067 VOUT+.n110 VOUT+.n109 0.3295
R2068 VOUT+.n111 VOUT+.n110 0.3295
R2069 VOUT+.n112 VOUT+.n111 0.3295
R2070 VOUT+.n113 VOUT+.n112 0.3295
R2071 VOUT+.n115 VOUT+.n113 0.3295
R2072 VOUT+.n115 VOUT+.n114 0.3295
R2073 VOUT+.n118 VOUT+.n116 0.3295
R2074 VOUT+.n118 VOUT+.n117 0.3295
R2075 VOUT+.n121 VOUT+.n119 0.3295
R2076 VOUT+.n121 VOUT+.n120 0.3295
R2077 VOUT+.n124 VOUT+.n122 0.3295
R2078 VOUT+.n124 VOUT+.n123 0.3295
R2079 VOUT+.n127 VOUT+.n125 0.3295
R2080 VOUT+.n127 VOUT+.n126 0.3295
R2081 VOUT+.n130 VOUT+.n128 0.3295
R2082 VOUT+.n130 VOUT+.n129 0.3295
R2083 VOUT+.n133 VOUT+.n131 0.3295
R2084 VOUT+.n133 VOUT+.n132 0.3295
R2085 VOUT+.n183 VOUT+.n182 0.3295
R2086 VOUT+.n182 VOUT+.n181 0.3295
R2087 VOUT+.n142 VOUT+.n138 0.3154
R2088 VOUT+.n20 VOUT+.n12 0.314966
R2089 VOUT+.n184 VOUT+.n183 0.313833
R2090 VOUT+.n146 VOUT+.n134 0.306
R2091 VOUT+.n145 VOUT+.n135 0.306
R2092 VOUT+.n144 VOUT+.n136 0.306
R2093 VOUT+.n143 VOUT+.n137 0.306
R2094 VOUT+.n153 VOUT+.n150 0.2825
R2095 VOUT+.n156 VOUT+.n153 0.2825
R2096 VOUT+.n159 VOUT+.n156 0.2825
R2097 VOUT+.n162 VOUT+.n159 0.2825
R2098 VOUT+.n165 VOUT+.n162 0.2825
R2099 VOUT+.n168 VOUT+.n165 0.2825
R2100 VOUT+.n171 VOUT+.n168 0.2825
R2101 VOUT+.n174 VOUT+.n171 0.2825
R2102 VOUT+.n177 VOUT+.n174 0.2825
R2103 VOUT+.n180 VOUT+.n177 0.2825
R2104 VOUT+.n115 VOUT+.n102 0.2825
R2105 VOUT+.n118 VOUT+.n115 0.2825
R2106 VOUT+.n121 VOUT+.n118 0.2825
R2107 VOUT+.n124 VOUT+.n121 0.2825
R2108 VOUT+.n127 VOUT+.n124 0.2825
R2109 VOUT+.n130 VOUT+.n127 0.2825
R2110 VOUT+.n133 VOUT+.n130 0.2825
R2111 VOUT+.n182 VOUT+.n133 0.2825
R2112 VOUT+.n182 VOUT+.n180 0.2825
R2113 VOUT+.n189 VOUT+.n92 0.2655
R2114 VOUT+.n194 VOUT+.n27 0.193208
R2115 VOUT+.n185 VOUT+.n184 0.138367
R2116 VOUT+.n18 VOUT+.n12 0.0891864
R2117 VOUT+.n69 VOUT+.n46 0.0577917
R2118 VOUT+.n73 VOUT+.n46 0.0577917
R2119 VOUT+.n74 VOUT+.n73 0.0577917
R2120 VOUT+.n75 VOUT+.n74 0.0577917
R2121 VOUT+.n75 VOUT+.n42 0.0577917
R2122 VOUT+.n79 VOUT+.n42 0.0577917
R2123 VOUT+.n80 VOUT+.n79 0.0577917
R2124 VOUT+.n81 VOUT+.n80 0.0577917
R2125 VOUT+.n72 VOUT+.n71 0.0577917
R2126 VOUT+.n72 VOUT+.n43 0.0577917
R2127 VOUT+.n76 VOUT+.n43 0.0577917
R2128 VOUT+.n77 VOUT+.n76 0.0577917
R2129 VOUT+.n78 VOUT+.n77 0.0577917
R2130 VOUT+.n78 VOUT+.n39 0.0577917
R2131 VOUT+.n82 VOUT+.n39 0.0577917
R2132 VOUT+.n70 VOUT+.n69 0.054517
R2133 VOUT+.n28 VOUT+.n7 0.047375
R2134 VOUT+ VOUT+.n2 0.047375
R2135 VOUT+.n190 VOUT+.n34 0.0421667
R2136 VOUT+.n91 VOUT+.n85 0.0421667
R2137 VOUT+.n19 VOUT+.n18 0.0421667
R2138 VOUT+.n19 VOUT+.n11 0.0421667
R2139 VOUT+.n23 VOUT+.n11 0.0421667
R2140 VOUT+.n24 VOUT+.n23 0.0421667
R2141 VOUT+.n25 VOUT+.n24 0.0421667
R2142 VOUT+.n21 VOUT+.n20 0.0421667
R2143 VOUT+.n22 VOUT+.n21 0.0421667
R2144 VOUT+.n22 VOUT+.n8 0.0421667
R2145 VOUT+.n26 VOUT+.n8 0.0421667
R2146 VOUT+.n86 VOUT+.n85 0.0243161
R2147 VOUT+.n88 VOUT+.n36 0.0243161
R2148 VOUT+.n88 VOUT+.n87 0.0243161
R2149 VOUT+.n86 VOUT+.n38 0.0243161
R2150 VOUT+.n187 VOUT+.n30 0.0217373
R2151 VOUT+.n87 VOUT+.n37 0.0217373
R2152 VOUT+.n95 VOUT+.n30 0.0217373
R2153 VOUT+.n6 VOUT+.n5 0.0217373
R2154 VOUT+.n5 VOUT+.n2 0.0217373
R2155 VOUT+.n93 VOUT+.n34 0.0217373
R2156 VOUT+.n95 VOUT+.n94 0.0217373
R2157 VOUT+.n83 VOUT+.n36 0.0217373
R2158 VOUT+.n83 VOUT+.n38 0.0217373
R2159 VOUT+.n93 VOUT+.n31 0.0217373
R2160 VOUT+.n94 VOUT+.n31 0.0217373
R2161 VOUT+.n194 VOUT+.n193 0.0217373
R2162 VOUT+.n7 VOUT+.n1 0.0217373
R2163 VOUT+ VOUT+.n1 0.0217373
R2164 VOUT+.n193 VOUT+.n28 0.0217373
R2165 VOUT+.n100 VOUT+.n99 0.0161667
R2166 VOUT+.n185 VOUT+.n100 0.0161667
R2167 VOUT+.n98 VOUT+.n97 0.0161667
R2168 VOUT+.n98 VOUT+.n96 0.0161667
R2169 VOUT+.n186 VOUT+.n96 0.0161667
R2170 VOUT+.n188 VOUT+.n32 0.0134654
R2171 VOUT+.n191 VOUT+.n29 0.0134654
R2172 VOUT+.n189 VOUT+.n188 0.0134654
R2173 VOUT+.n32 VOUT+.n29 0.0134654
R2174 VOUT+.n89 VOUT+.n84 0.0109778
R2175 VOUT+.n92 VOUT+.n35 0.0109778
R2176 VOUT+.n195 VOUT+.n3 0.0109778
R2177 VOUT+.n4 VOUT+.n0 0.0109778
R2178 VOUT+.n90 VOUT+.n89 0.0109778
R2179 VOUT+.n84 VOUT+.n35 0.0109778
R2180 VOUT+.n192 VOUT+.n3 0.0109778
R2181 VOUT+.n195 VOUT+.n4 0.0109778
R2182 VOUT+.n97 VOUT+.n33 0.00872683
R2183 cap_res_Y cap_res_Y.t0 49.4263
R2184 cap_res_Y cap_res_Y.t25 1.481
R2185 cap_res_Y.t17 cap_res_Y.t133 0.1603
R2186 cap_res_Y.t114 cap_res_Y.t98 0.1603
R2187 cap_res_Y.t47 cap_res_Y.t63 0.1603
R2188 cap_res_Y.t74 cap_res_Y.t126 0.1603
R2189 cap_res_Y.t9 cap_res_Y.t95 0.1603
R2190 cap_res_Y.t112 cap_res_Y.t30 0.1603
R2191 cap_res_Y.t52 cap_res_Y.t137 0.1603
R2192 cap_res_Y.t18 cap_res_Y.t65 0.1603
R2193 cap_res_Y.t87 cap_res_Y.t38 0.1603
R2194 cap_res_Y.t118 cap_res_Y.t35 0.1603
R2195 cap_res_Y.t56 cap_res_Y.t5 0.1603
R2196 cap_res_Y.t22 cap_res_Y.t70 0.1603
R2197 cap_res_Y.t92 cap_res_Y.t44 0.1603
R2198 cap_res_Y.t59 cap_res_Y.t106 0.1603
R2199 cap_res_Y.t132 cap_res_Y.t79 0.1603
R2200 cap_res_Y.t28 cap_res_Y.t75 0.1603
R2201 cap_res_Y.t99 cap_res_Y.t51 0.1603
R2202 cap_res_Y.t64 cap_res_Y.t113 0.1603
R2203 cap_res_Y.t1 cap_res_Y.t85 0.1603
R2204 cap_res_Y.t104 cap_res_Y.t19 0.1603
R2205 cap_res_Y.t39 cap_res_Y.t122 0.1603
R2206 cap_res_Y.t68 cap_res_Y.t119 0.1603
R2207 cap_res_Y.t6 cap_res_Y.t90 0.1603
R2208 cap_res_Y.t105 cap_res_Y.t23 0.1603
R2209 cap_res_Y.t45 cap_res_Y.t131 0.1603
R2210 cap_res_Y.t15 cap_res_Y.t61 0.1603
R2211 cap_res_Y.t81 cap_res_Y.t32 0.1603
R2212 cap_res_Y.t77 cap_res_Y.t116 0.1603
R2213 cap_res_Y.t43 cap_res_Y.t3 0.1603
R2214 cap_res_Y.t48 cap_res_Y.t86 0.1603
R2215 cap_res_Y.t8 cap_res_Y.t102 0.1603
R2216 cap_res_Y.t50 cap_res_Y.t97 0.1603
R2217 cap_res_Y.t110 cap_res_Y.t62 0.1603
R2218 cap_res_Y.t42 cap_res_Y.t20 0.1603
R2219 cap_res_Y.t103 cap_res_Y.t124 0.1603
R2220 cap_res_Y.t71 cap_res_Y.t57 0.1603
R2221 cap_res_Y.t138 cap_res_Y.t96 0.1603
R2222 cap_res_Y.t36 cap_res_Y.t136 0.1603
R2223 cap_res_Y.t69 cap_res_Y.t34 0.1603
R2224 cap_res_Y.t55 cap_res_Y.t12 0.1603
R2225 cap_res_Y.t89 cap_res_Y.t54 0.1603
R2226 cap_res_Y.t66 cap_res_Y.t31 0.1603
R2227 cap_res_Y.t53 cap_res_Y.t10 0.1603
R2228 cap_res_Y.t84 cap_res_Y.t49 0.1603
R2229 cap_res_Y.t120 cap_res_Y.t83 0.1603
R2230 cap_res_Y.t21 cap_res_Y.t115 0.1603
R2231 cap_res_Y.t4 cap_res_Y.t100 0.1603
R2232 cap_res_Y.t37 cap_res_Y.t16 0.1603
R2233 cap_res_Y.t101 cap_res_Y.t76 0.1603
R2234 cap_res_Y.t29 cap_res_Y.t58 0.1603
R2235 cap_res_Y.t60 cap_res_Y.t29 0.1603
R2236 cap_res_Y.t107 cap_res_Y.t72 0.1603
R2237 cap_res_Y.t14 cap_res_Y.t107 0.1603
R2238 cap_res_Y.t127 cap_res_Y.t93 0.1603
R2239 cap_res_Y.t135 cap_res_Y.t121 0.1603
R2240 cap_res_Y.t27 cap_res_Y.t135 0.1603
R2241 cap_res_Y.t108 cap_res_Y.t78 0.1603
R2242 cap_res_Y.t11 cap_res_Y.t108 0.1603
R2243 cap_res_Y.t91 cap_res_Y.t130 0.1603
R2244 cap_res_Y.t123 cap_res_Y.t91 0.1603
R2245 cap_res_Y.t128 cap_res_Y.t24 0.1603
R2246 cap_res_Y.t25 cap_res_Y.t128 0.1603
R2247 cap_res_Y.t41 cap_res_Y.n14 0.159278
R2248 cap_res_Y.t7 cap_res_Y.n15 0.159278
R2249 cap_res_Y.t13 cap_res_Y.n16 0.159278
R2250 cap_res_Y.t94 cap_res_Y.n17 0.159278
R2251 cap_res_Y.t129 cap_res_Y.n18 0.159278
R2252 cap_res_Y.t111 cap_res_Y.n19 0.159278
R2253 cap_res_Y.t73 cap_res_Y.n20 0.159278
R2254 cap_res_Y.t40 cap_res_Y.n21 0.159278
R2255 cap_res_Y.t67 cap_res_Y.n22 0.159278
R2256 cap_res_Y.t33 cap_res_Y.n23 0.159278
R2257 cap_res_Y.t134 cap_res_Y.n24 0.159278
R2258 cap_res_Y.t26 cap_res_Y.n25 0.159278
R2259 cap_res_Y.t125 cap_res_Y.n26 0.159278
R2260 cap_res_Y.t88 cap_res_Y.n27 0.159278
R2261 cap_res_Y.t117 cap_res_Y.n28 0.159278
R2262 cap_res_Y.t82 cap_res_Y.n29 0.159278
R2263 cap_res_Y.t46 cap_res_Y.n30 0.159278
R2264 cap_res_Y.t80 cap_res_Y.n31 0.159278
R2265 cap_res_Y.t109 cap_res_Y.n32 0.159278
R2266 cap_res_Y.n33 cap_res_Y.t17 0.1368
R2267 cap_res_Y.n32 cap_res_Y.t114 0.1368
R2268 cap_res_Y.n32 cap_res_Y.t47 0.1368
R2269 cap_res_Y.n31 cap_res_Y.t74 0.1368
R2270 cap_res_Y.n31 cap_res_Y.t9 0.1368
R2271 cap_res_Y.n30 cap_res_Y.t112 0.1368
R2272 cap_res_Y.n30 cap_res_Y.t52 0.1368
R2273 cap_res_Y.n29 cap_res_Y.t18 0.1368
R2274 cap_res_Y.n29 cap_res_Y.t87 0.1368
R2275 cap_res_Y.n28 cap_res_Y.t118 0.1368
R2276 cap_res_Y.n28 cap_res_Y.t56 0.1368
R2277 cap_res_Y.n27 cap_res_Y.t22 0.1368
R2278 cap_res_Y.n27 cap_res_Y.t92 0.1368
R2279 cap_res_Y.n26 cap_res_Y.t59 0.1368
R2280 cap_res_Y.n26 cap_res_Y.t132 0.1368
R2281 cap_res_Y.n25 cap_res_Y.t28 0.1368
R2282 cap_res_Y.n25 cap_res_Y.t99 0.1368
R2283 cap_res_Y.n24 cap_res_Y.t64 0.1368
R2284 cap_res_Y.n24 cap_res_Y.t1 0.1368
R2285 cap_res_Y.n23 cap_res_Y.t104 0.1368
R2286 cap_res_Y.n23 cap_res_Y.t39 0.1368
R2287 cap_res_Y.n22 cap_res_Y.t68 0.1368
R2288 cap_res_Y.n22 cap_res_Y.t6 0.1368
R2289 cap_res_Y.n21 cap_res_Y.t105 0.1368
R2290 cap_res_Y.n21 cap_res_Y.t45 0.1368
R2291 cap_res_Y.n20 cap_res_Y.t15 0.1368
R2292 cap_res_Y.n20 cap_res_Y.t81 0.1368
R2293 cap_res_Y.n19 cap_res_Y.t77 0.1368
R2294 cap_res_Y.n19 cap_res_Y.t43 0.1368
R2295 cap_res_Y.n18 cap_res_Y.t48 0.1368
R2296 cap_res_Y.n18 cap_res_Y.t8 0.1368
R2297 cap_res_Y.n17 cap_res_Y.t50 0.1368
R2298 cap_res_Y.n17 cap_res_Y.t110 0.1368
R2299 cap_res_Y.n16 cap_res_Y.t42 0.1368
R2300 cap_res_Y.n16 cap_res_Y.t103 0.1368
R2301 cap_res_Y.n15 cap_res_Y.t71 0.1368
R2302 cap_res_Y.n14 cap_res_Y.t37 0.1368
R2303 cap_res_Y.t76 cap_res_Y.n33 0.1368
R2304 cap_res_Y.n34 cap_res_Y.t101 0.1368
R2305 cap_res_Y.n0 cap_res_Y.t14 0.1368
R2306 cap_res_Y.n4 cap_res_Y.t138 0.114322
R2307 cap_res_Y.n5 cap_res_Y.n4 0.1133
R2308 cap_res_Y.n6 cap_res_Y.n5 0.1133
R2309 cap_res_Y.n7 cap_res_Y.n6 0.1133
R2310 cap_res_Y.n8 cap_res_Y.n7 0.1133
R2311 cap_res_Y.n9 cap_res_Y.n8 0.1133
R2312 cap_res_Y.n10 cap_res_Y.n9 0.1133
R2313 cap_res_Y.n11 cap_res_Y.n10 0.1133
R2314 cap_res_Y.n12 cap_res_Y.n11 0.1133
R2315 cap_res_Y.n13 cap_res_Y.n12 0.1133
R2316 cap_res_Y.n15 cap_res_Y.n13 0.1133
R2317 cap_res_Y.n1 cap_res_Y.n0 0.1133
R2318 cap_res_Y.n2 cap_res_Y.n1 0.1133
R2319 cap_res_Y.n3 cap_res_Y.n2 0.1133
R2320 cap_res_Y.n35 cap_res_Y.n3 0.1133
R2321 cap_res_Y.n35 cap_res_Y.n34 0.1133
R2322 cap_res_Y.n4 cap_res_Y.t36 0.00152174
R2323 cap_res_Y.n5 cap_res_Y.t69 0.00152174
R2324 cap_res_Y.n6 cap_res_Y.t55 0.00152174
R2325 cap_res_Y.n7 cap_res_Y.t89 0.00152174
R2326 cap_res_Y.n8 cap_res_Y.t66 0.00152174
R2327 cap_res_Y.n9 cap_res_Y.t53 0.00152174
R2328 cap_res_Y.n10 cap_res_Y.t84 0.00152174
R2329 cap_res_Y.n11 cap_res_Y.t120 0.00152174
R2330 cap_res_Y.n12 cap_res_Y.t21 0.00152174
R2331 cap_res_Y.n13 cap_res_Y.t4 0.00152174
R2332 cap_res_Y.n14 cap_res_Y.t2 0.00152174
R2333 cap_res_Y.n15 cap_res_Y.t41 0.00152174
R2334 cap_res_Y.n16 cap_res_Y.t7 0.00152174
R2335 cap_res_Y.n17 cap_res_Y.t13 0.00152174
R2336 cap_res_Y.n18 cap_res_Y.t94 0.00152174
R2337 cap_res_Y.n19 cap_res_Y.t129 0.00152174
R2338 cap_res_Y.n20 cap_res_Y.t111 0.00152174
R2339 cap_res_Y.n21 cap_res_Y.t73 0.00152174
R2340 cap_res_Y.n22 cap_res_Y.t40 0.00152174
R2341 cap_res_Y.n23 cap_res_Y.t67 0.00152174
R2342 cap_res_Y.n24 cap_res_Y.t33 0.00152174
R2343 cap_res_Y.n25 cap_res_Y.t134 0.00152174
R2344 cap_res_Y.n26 cap_res_Y.t26 0.00152174
R2345 cap_res_Y.n27 cap_res_Y.t125 0.00152174
R2346 cap_res_Y.n28 cap_res_Y.t88 0.00152174
R2347 cap_res_Y.n29 cap_res_Y.t117 0.00152174
R2348 cap_res_Y.n30 cap_res_Y.t82 0.00152174
R2349 cap_res_Y.n31 cap_res_Y.t46 0.00152174
R2350 cap_res_Y.n32 cap_res_Y.t80 0.00152174
R2351 cap_res_Y.n33 cap_res_Y.t109 0.00152174
R2352 cap_res_Y.n34 cap_res_Y.t60 0.00152174
R2353 cap_res_Y.n0 cap_res_Y.t127 0.00152174
R2354 cap_res_Y.n1 cap_res_Y.t27 0.00152174
R2355 cap_res_Y.n2 cap_res_Y.t11 0.00152174
R2356 cap_res_Y.n3 cap_res_Y.t123 0.00152174
R2357 cap_res_Y.t24 cap_res_Y.n35 0.00152174
R2358 V_CMFB_S2.n19 V_CMFB_S2.t0 119.785
R2359 V_CMFB_S2.n17 V_CMFB_S2.n16 24.288
R2360 V_CMFB_S2.n14 V_CMFB_S2.n13 24.288
R2361 V_CMFB_S2.n11 V_CMFB_S2.n10 24.288
R2362 V_CMFB_S2.n7 V_CMFB_S2.n6 24.288
R2363 V_CMFB_S2.n3 V_CMFB_S2.n2 24.288
R2364 V_CMFB_S2.n16 V_CMFB_S2.t1 8.0005
R2365 V_CMFB_S2.n16 V_CMFB_S2.t7 8.0005
R2366 V_CMFB_S2.n13 V_CMFB_S2.t4 8.0005
R2367 V_CMFB_S2.n13 V_CMFB_S2.t8 8.0005
R2368 V_CMFB_S2.n10 V_CMFB_S2.t2 8.0005
R2369 V_CMFB_S2.n10 V_CMFB_S2.t6 8.0005
R2370 V_CMFB_S2.n6 V_CMFB_S2.t10 8.0005
R2371 V_CMFB_S2.n6 V_CMFB_S2.t5 8.0005
R2372 V_CMFB_S2.n2 V_CMFB_S2.t9 8.0005
R2373 V_CMFB_S2.n2 V_CMFB_S2.t3 8.0005
R2374 V_CMFB_S2.n3 V_CMFB_S2.n1 5.7505
R2375 V_CMFB_S2.n17 V_CMFB_S2.n15 5.7505
R2376 V_CMFB_S2.n19 V_CMFB_S2.n18 5.6255
R2377 V_CMFB_S2.n14 V_CMFB_S2.n0 5.188
R2378 V_CMFB_S2.n15 V_CMFB_S2.n14 5.188
R2379 V_CMFB_S2.n11 V_CMFB_S2.n9 5.188
R2380 V_CMFB_S2.n12 V_CMFB_S2.n11 5.188
R2381 V_CMFB_S2.n8 V_CMFB_S2.n7 5.188
R2382 V_CMFB_S2.n7 V_CMFB_S2.n1 5.188
R2383 V_CMFB_S2.n18 V_CMFB_S2.n17 5.188
R2384 V_CMFB_S2.n8 V_CMFB_S2.n5 5.063
R2385 V_CMFB_S2.n5 V_CMFB_S2.n4 2.0005
R2386 V_CMFB_S2.n5 V_CMFB_S2.n3 0.6255
R2387 V_CMFB_S2.n12 V_CMFB_S2.n1 0.563
R2388 V_CMFB_S2.n15 V_CMFB_S2.n12 0.563
R2389 V_CMFB_S2.n18 V_CMFB_S2.n0 0.563
R2390 V_CMFB_S2.n9 V_CMFB_S2.n0 0.563
R2391 V_CMFB_S2.n9 V_CMFB_S2.n8 0.563
R2392 V_CMFB_S2 V_CMFB_S2.n19 0.063
R2393 cap_res_X cap_res_X.t0 49.4254
R2394 cap_res_X cap_res_X.t63 1.481
R2395 cap_res_X.t58 cap_res_X.t99 0.1603
R2396 cap_res_X.t23 cap_res_X.t58 0.1603
R2397 cap_res_X.t126 cap_res_X.t89 0.1603
R2398 cap_res_X.t110 cap_res_X.t43 0.1603
R2399 cap_res_X.t6 cap_res_X.t110 0.1603
R2400 cap_res_X.t73 cap_res_X.t9 0.1603
R2401 cap_res_X.t106 cap_res_X.t73 0.1603
R2402 cap_res_X.t35 cap_res_X.t112 0.1603
R2403 cap_res_X.t69 cap_res_X.t35 0.1603
R2404 cap_res_X.t18 cap_res_X.t125 0.1603
R2405 cap_res_X.t59 cap_res_X.t37 0.1603
R2406 cap_res_X.t127 cap_res_X.t88 0.1603
R2407 cap_res_X.t21 cap_res_X.t71 0.1603
R2408 cap_res_X.t91 cap_res_X.t52 0.1603
R2409 cap_res_X.t60 cap_res_X.t111 0.1603
R2410 cap_res_X.t133 cap_res_X.t97 0.1603
R2411 cap_res_X.t101 cap_res_X.t11 0.1603
R2412 cap_res_X.t32 cap_res_X.t136 0.1603
R2413 cap_res_X.t65 cap_res_X.t117 0.1603
R2414 cap_res_X.t137 cap_res_X.t102 0.1603
R2415 cap_res_X.t104 cap_res_X.t16 0.1603
R2416 cap_res_X.t36 cap_res_X.t1 0.1603
R2417 cap_res_X.t4 cap_res_X.t54 0.1603
R2418 cap_res_X.t74 cap_res_X.t39 0.1603
R2419 cap_res_X.t108 cap_res_X.t22 0.1603
R2420 cap_res_X.t40 cap_res_X.t5 0.1603
R2421 cap_res_X.t10 cap_res_X.t62 0.1603
R2422 cap_res_X.t80 cap_res_X.t47 0.1603
R2423 cap_res_X.t49 cap_res_X.t103 0.1603
R2424 cap_res_X.t121 cap_res_X.t86 0.1603
R2425 cap_res_X.t14 cap_res_X.t66 0.1603
R2426 cap_res_X.t87 cap_res_X.t50 0.1603
R2427 cap_res_X.t53 cap_res_X.t105 0.1603
R2428 cap_res_X.t128 cap_res_X.t90 0.1603
R2429 cap_res_X.t98 cap_res_X.t7 0.1603
R2430 cap_res_X.t26 cap_res_X.t132 0.1603
R2431 cap_res_X.t68 cap_res_X.t109 0.1603
R2432 cap_res_X.t31 cap_res_X.t82 0.1603
R2433 cap_res_X.t34 cap_res_X.t77 0.1603
R2434 cap_res_X.t138 cap_res_X.t48 0.1603
R2435 cap_res_X.t131 cap_res_X.t41 0.1603
R2436 cap_res_X.t57 cap_res_X.t25 0.1603
R2437 cap_res_X.t124 cap_res_X.t100 0.1603
R2438 cap_res_X.t46 cap_res_X.t8 0.1603
R2439 cap_res_X.t17 cap_res_X.t119 0.1603
R2440 cap_res_X.t123 cap_res_X.t81 0.1603
R2441 cap_res_X.t83 cap_res_X.t44 0.1603
R2442 cap_res_X.t45 cap_res_X.t3 0.1603
R2443 cap_res_X.t67 cap_res_X.t29 0.1603
R2444 cap_res_X.t30 cap_res_X.t130 0.1603
R2445 cap_res_X.t134 cap_res_X.t92 0.1603
R2446 cap_res_X.t12 cap_res_X.t113 0.1603
R2447 cap_res_X.t114 cap_res_X.t75 0.1603
R2448 cap_res_X.t135 cap_res_X.t94 0.1603
R2449 cap_res_X.t15 cap_res_X.t116 0.1603
R2450 cap_res_X.t79 cap_res_X.t42 0.1603
R2451 cap_res_X.t38 cap_res_X.t2 0.1603
R2452 cap_res_X.t72 cap_res_X.t96 0.1603
R2453 cap_res_X.t19 cap_res_X.t28 0.1603
R2454 cap_res_X.t51 cap_res_X.t19 0.1603
R2455 cap_res_X.t56 cap_res_X.t93 0.1603
R2456 cap_res_X.t63 cap_res_X.t56 0.1603
R2457 cap_res_X.t118 cap_res_X.n10 0.159278
R2458 cap_res_X.t84 cap_res_X.n11 0.159278
R2459 cap_res_X.t95 cap_res_X.n12 0.159278
R2460 cap_res_X.t85 cap_res_X.n13 0.159278
R2461 cap_res_X.t120 cap_res_X.n14 0.159278
R2462 cap_res_X.t61 cap_res_X.n15 0.159278
R2463 cap_res_X.t20 cap_res_X.n16 0.159278
R2464 cap_res_X.t122 cap_res_X.n17 0.159278
R2465 cap_res_X.t13 cap_res_X.n18 0.159278
R2466 cap_res_X.t115 cap_res_X.n19 0.159278
R2467 cap_res_X.t76 cap_res_X.n20 0.159278
R2468 cap_res_X.t107 cap_res_X.n21 0.159278
R2469 cap_res_X.t70 cap_res_X.n22 0.159278
R2470 cap_res_X.t33 cap_res_X.n23 0.159278
R2471 cap_res_X.t64 cap_res_X.n24 0.159278
R2472 cap_res_X.t27 cap_res_X.n25 0.159278
R2473 cap_res_X.t129 cap_res_X.n26 0.159278
R2474 cap_res_X.t24 cap_res_X.n27 0.159278
R2475 cap_res_X.t55 cap_res_X.n28 0.159278
R2476 cap_res_X.n31 cap_res_X.t23 0.1368
R2477 cap_res_X.n29 cap_res_X.t18 0.1368
R2478 cap_res_X.n28 cap_res_X.t59 0.1368
R2479 cap_res_X.n28 cap_res_X.t127 0.1368
R2480 cap_res_X.n27 cap_res_X.t21 0.1368
R2481 cap_res_X.n27 cap_res_X.t91 0.1368
R2482 cap_res_X.n26 cap_res_X.t60 0.1368
R2483 cap_res_X.n26 cap_res_X.t133 0.1368
R2484 cap_res_X.n25 cap_res_X.t101 0.1368
R2485 cap_res_X.n25 cap_res_X.t32 0.1368
R2486 cap_res_X.n24 cap_res_X.t65 0.1368
R2487 cap_res_X.n24 cap_res_X.t137 0.1368
R2488 cap_res_X.n23 cap_res_X.t104 0.1368
R2489 cap_res_X.n23 cap_res_X.t36 0.1368
R2490 cap_res_X.n22 cap_res_X.t4 0.1368
R2491 cap_res_X.n22 cap_res_X.t74 0.1368
R2492 cap_res_X.n21 cap_res_X.t108 0.1368
R2493 cap_res_X.n21 cap_res_X.t40 0.1368
R2494 cap_res_X.n20 cap_res_X.t10 0.1368
R2495 cap_res_X.n20 cap_res_X.t80 0.1368
R2496 cap_res_X.n19 cap_res_X.t49 0.1368
R2497 cap_res_X.n19 cap_res_X.t121 0.1368
R2498 cap_res_X.n18 cap_res_X.t14 0.1368
R2499 cap_res_X.n18 cap_res_X.t87 0.1368
R2500 cap_res_X.n17 cap_res_X.t53 0.1368
R2501 cap_res_X.n17 cap_res_X.t128 0.1368
R2502 cap_res_X.n16 cap_res_X.t98 0.1368
R2503 cap_res_X.n16 cap_res_X.t26 0.1368
R2504 cap_res_X.n15 cap_res_X.t68 0.1368
R2505 cap_res_X.n15 cap_res_X.t31 0.1368
R2506 cap_res_X.n14 cap_res_X.t34 0.1368
R2507 cap_res_X.n14 cap_res_X.t138 0.1368
R2508 cap_res_X.n13 cap_res_X.t131 0.1368
R2509 cap_res_X.n13 cap_res_X.t57 0.1368
R2510 cap_res_X.n12 cap_res_X.t124 0.1368
R2511 cap_res_X.n12 cap_res_X.t46 0.1368
R2512 cap_res_X.n11 cap_res_X.t79 0.1368
R2513 cap_res_X.n10 cap_res_X.t38 0.1368
R2514 cap_res_X.t96 cap_res_X.n29 0.1368
R2515 cap_res_X.n30 cap_res_X.t72 0.1368
R2516 cap_res_X.n0 cap_res_X.t17 0.114322
R2517 cap_res_X.n32 cap_res_X.n31 0.1133
R2518 cap_res_X.n33 cap_res_X.n32 0.1133
R2519 cap_res_X.n34 cap_res_X.n33 0.1133
R2520 cap_res_X.n1 cap_res_X.n0 0.1133
R2521 cap_res_X.n2 cap_res_X.n1 0.1133
R2522 cap_res_X.n3 cap_res_X.n2 0.1133
R2523 cap_res_X.n4 cap_res_X.n3 0.1133
R2524 cap_res_X.n5 cap_res_X.n4 0.1133
R2525 cap_res_X.n6 cap_res_X.n5 0.1133
R2526 cap_res_X.n7 cap_res_X.n6 0.1133
R2527 cap_res_X.n8 cap_res_X.n7 0.1133
R2528 cap_res_X.n9 cap_res_X.n8 0.1133
R2529 cap_res_X.n11 cap_res_X.n9 0.1133
R2530 cap_res_X.n35 cap_res_X.n30 0.1133
R2531 cap_res_X.n35 cap_res_X.n34 0.1133
R2532 cap_res_X.n31 cap_res_X.t126 0.00152174
R2533 cap_res_X.n32 cap_res_X.t6 0.00152174
R2534 cap_res_X.n33 cap_res_X.t106 0.00152174
R2535 cap_res_X.n34 cap_res_X.t69 0.00152174
R2536 cap_res_X.n0 cap_res_X.t123 0.00152174
R2537 cap_res_X.n1 cap_res_X.t83 0.00152174
R2538 cap_res_X.n2 cap_res_X.t45 0.00152174
R2539 cap_res_X.n3 cap_res_X.t67 0.00152174
R2540 cap_res_X.n4 cap_res_X.t30 0.00152174
R2541 cap_res_X.n5 cap_res_X.t134 0.00152174
R2542 cap_res_X.n6 cap_res_X.t12 0.00152174
R2543 cap_res_X.n7 cap_res_X.t114 0.00152174
R2544 cap_res_X.n8 cap_res_X.t135 0.00152174
R2545 cap_res_X.n9 cap_res_X.t15 0.00152174
R2546 cap_res_X.n10 cap_res_X.t78 0.00152174
R2547 cap_res_X.n11 cap_res_X.t118 0.00152174
R2548 cap_res_X.n12 cap_res_X.t84 0.00152174
R2549 cap_res_X.n13 cap_res_X.t95 0.00152174
R2550 cap_res_X.n14 cap_res_X.t85 0.00152174
R2551 cap_res_X.n15 cap_res_X.t120 0.00152174
R2552 cap_res_X.n16 cap_res_X.t61 0.00152174
R2553 cap_res_X.n17 cap_res_X.t20 0.00152174
R2554 cap_res_X.n18 cap_res_X.t122 0.00152174
R2555 cap_res_X.n19 cap_res_X.t13 0.00152174
R2556 cap_res_X.n20 cap_res_X.t115 0.00152174
R2557 cap_res_X.n21 cap_res_X.t76 0.00152174
R2558 cap_res_X.n22 cap_res_X.t107 0.00152174
R2559 cap_res_X.n23 cap_res_X.t70 0.00152174
R2560 cap_res_X.n24 cap_res_X.t33 0.00152174
R2561 cap_res_X.n25 cap_res_X.t64 0.00152174
R2562 cap_res_X.n26 cap_res_X.t27 0.00152174
R2563 cap_res_X.n27 cap_res_X.t129 0.00152174
R2564 cap_res_X.n28 cap_res_X.t24 0.00152174
R2565 cap_res_X.n29 cap_res_X.t55 0.00152174
R2566 cap_res_X.n30 cap_res_X.t51 0.00152174
R2567 cap_res_X.t93 cap_res_X.n35 0.00152174
R2568 Vb3.n19 Vb3.t9 768.551
R2569 Vb3.n13 Vb3.t3 611.739
R2570 Vb3.n9 Vb3.t21 611.739
R2571 Vb3.n4 Vb3.t12 611.739
R2572 Vb3.n0 Vb3.t22 611.739
R2573 Vb3.n20 Vb3.n17 431.07
R2574 Vb3 Vb3.n8 430.226
R2575 Vb3.n13 Vb3.t20 421.75
R2576 Vb3.n14 Vb3.t17 421.75
R2577 Vb3.n15 Vb3.t15 421.75
R2578 Vb3.n16 Vb3.t11 421.75
R2579 Vb3.n9 Vb3.t19 421.75
R2580 Vb3.n10 Vb3.t2 421.75
R2581 Vb3.n11 Vb3.t5 421.75
R2582 Vb3.n12 Vb3.t7 421.75
R2583 Vb3.n4 Vb3.t8 421.75
R2584 Vb3.n5 Vb3.t18 421.75
R2585 Vb3.n6 Vb3.t16 421.75
R2586 Vb3.n7 Vb3.t13 421.75
R2587 Vb3.n0 Vb3.t4 421.75
R2588 Vb3.n1 Vb3.t6 421.75
R2589 Vb3.n2 Vb3.t10 421.75
R2590 Vb3.n3 Vb3.t14 421.75
R2591 Vb3.n14 Vb3.n13 167.094
R2592 Vb3.n15 Vb3.n14 167.094
R2593 Vb3.n16 Vb3.n15 167.094
R2594 Vb3.n10 Vb3.n9 167.094
R2595 Vb3.n11 Vb3.n10 167.094
R2596 Vb3.n12 Vb3.n11 167.094
R2597 Vb3.n5 Vb3.n4 167.094
R2598 Vb3.n6 Vb3.n5 167.094
R2599 Vb3.n7 Vb3.n6 167.094
R2600 Vb3.n1 Vb3.n0 167.094
R2601 Vb3.n2 Vb3.n1 167.094
R2602 Vb3.n3 Vb3.n2 167.094
R2603 Vb3.n19 Vb3.n18 74.6588
R2604 Vb3.n17 Vb3.n16 35.3472
R2605 Vb3.n17 Vb3.n12 35.3472
R2606 Vb3.n8 Vb3.n7 35.3472
R2607 Vb3.n8 Vb3.n3 35.3472
R2608 Vb3.n20 Vb3.n19 15.563
R2609 Vb3.n18 Vb3.t0 11.2576
R2610 Vb3.n18 Vb3.t1 11.2576
R2611 Vb3 Vb3.n20 0.28175
R2612 VD4.n16 VD4.t26 672.293
R2613 VD4.n31 VD4.t29 672.293
R2614 VD4.n30 VD4.t30 213.131
R2615 VD4.t27 VD4.n29 213.131
R2616 VD4.t30 VD4.t0 146.155
R2617 VD4.t0 VD4.t2 146.155
R2618 VD4.t2 VD4.t6 146.155
R2619 VD4.t6 VD4.t36 146.155
R2620 VD4.t36 VD4.t14 146.155
R2621 VD4.t14 VD4.t10 146.155
R2622 VD4.t10 VD4.t8 146.155
R2623 VD4.t8 VD4.t4 146.155
R2624 VD4.t4 VD4.t12 146.155
R2625 VD4.t12 VD4.t34 146.155
R2626 VD4.t34 VD4.t27 146.155
R2627 VD4.n30 VD4.t31 76.2576
R2628 VD4.n29 VD4.t28 76.2576
R2629 VD4.n28 VD4.n27 66.9922
R2630 VD4.n36 VD4.n26 66.9922
R2631 VD4.n41 VD4.n23 66.9922
R2632 VD4.n46 VD4.n20 66.9922
R2633 VD4.n18 VD4.n17 66.9922
R2634 VD4.n62 VD4.n61 66.0338
R2635 VD4.n59 VD4.n58 66.0338
R2636 VD4.n14 VD4.n13 66.0338
R2637 VD4.n12 VD4.n11 66.0338
R2638 VD4.n67 VD4.n66 66.0338
R2639 VD4.n70 VD4.n69 66.0338
R2640 VD4.n61 VD4.t33 11.2576
R2641 VD4.n61 VD4.t24 11.2576
R2642 VD4.n58 VD4.t17 11.2576
R2643 VD4.n58 VD4.t19 11.2576
R2644 VD4.n13 VD4.t20 11.2576
R2645 VD4.n13 VD4.t21 11.2576
R2646 VD4.n11 VD4.t22 11.2576
R2647 VD4.n11 VD4.t23 11.2576
R2648 VD4.n66 VD4.t16 11.2576
R2649 VD4.n66 VD4.t32 11.2576
R2650 VD4.n27 VD4.t1 11.2576
R2651 VD4.n27 VD4.t3 11.2576
R2652 VD4.n26 VD4.t7 11.2576
R2653 VD4.n26 VD4.t37 11.2576
R2654 VD4.n23 VD4.t15 11.2576
R2655 VD4.n23 VD4.t11 11.2576
R2656 VD4.n20 VD4.t9 11.2576
R2657 VD4.n20 VD4.t5 11.2576
R2658 VD4.n17 VD4.t13 11.2576
R2659 VD4.n17 VD4.t35 11.2576
R2660 VD4.t25 VD4.n70 11.2576
R2661 VD4.n70 VD4.t18 11.2576
R2662 VD4.n68 VD4.n67 5.91717
R2663 VD4.n62 VD4.n60 5.91717
R2664 VD4.n60 VD4.n59 5.29217
R2665 VD4.n57 VD4.n14 5.29217
R2666 VD4.n12 VD4.n10 5.29217
R2667 VD4.n69 VD4.n68 5.29217
R2668 VD4.n55 VD4.n54 1.5005
R2669 VD4.n53 VD4.n15 1.5005
R2670 VD4.n52 VD4.n51 1.5005
R2671 VD4.n50 VD4.n18 1.5005
R2672 VD4.n49 VD4.n48 1.5005
R2673 VD4.n47 VD4.n19 1.5005
R2674 VD4.n46 VD4.n45 1.5005
R2675 VD4.n44 VD4.n21 1.5005
R2676 VD4.n43 VD4.n42 1.5005
R2677 VD4.n41 VD4.n22 1.5005
R2678 VD4.n40 VD4.n39 1.5005
R2679 VD4.n38 VD4.n24 1.5005
R2680 VD4.n37 VD4.n36 1.5005
R2681 VD4.n35 VD4.n25 1.5005
R2682 VD4.n34 VD4.n33 1.5005
R2683 VD4.n0 VD4.n1 0.740726
R2684 VD4.n64 VD4.n63 1.5005
R2685 VD4.n8 VD4.n7 0.740726
R2686 VD4.n2 VD4.n6 0.740726
R2687 VD4.n5 VD4.n4 0.740726
R2688 VD4.n3 VD4.n56 1.5005
R2689 VD4.n31 VD4.n30 1.03383
R2690 VD4.n29 VD4.n16 1.03383
R2691 VD4.n32 VD4.n31 1.02322
R2692 VD4.n67 VD4.n65 1.02322
R2693 VD4.n59 VD4.n2 0.958833
R2694 VD4.n7 VD4.n14 0.958833
R2695 VD4.n64 VD4.n12 0.958833
R2696 VD4.n54 VD4.n16 0.958833
R2697 VD4.n3 VD4.n62 0.958833
R2698 VD4.n69 VD4.n9 0.958833
R2699 VD4.n56 VD4.n55 0.786958
R2700 VD4.n60 VD4.n57 0.6255
R2701 VD4.n57 VD4.n10 0.6255
R2702 VD4.n68 VD4.n10 0.6255
R2703 VD4.n33 VD4.n32 0.427973
R2704 VD4.n65 VD4.n0 0.427973
R2705 VD4.n7 VD4.n2 0.0838333
R2706 VD4.n32 VD4.n28 0.0587394
R2707 VD4.n65 VD4.n9 0.0587394
R2708 VD4.n1 VD4.n64 0.0632146
R2709 VD4.n9 VD4.n1 0.0632146
R2710 VD4.n34 VD4.n28 0.0421667
R2711 VD4.n35 VD4.n34 0.0421667
R2712 VD4.n36 VD4.n35 0.0421667
R2713 VD4.n36 VD4.n24 0.0421667
R2714 VD4.n40 VD4.n24 0.0421667
R2715 VD4.n41 VD4.n40 0.0421667
R2716 VD4.n42 VD4.n41 0.0421667
R2717 VD4.n42 VD4.n21 0.0421667
R2718 VD4.n46 VD4.n21 0.0421667
R2719 VD4.n47 VD4.n46 0.0421667
R2720 VD4.n48 VD4.n47 0.0421667
R2721 VD4.n48 VD4.n18 0.0421667
R2722 VD4.n52 VD4.n18 0.0421667
R2723 VD4.n53 VD4.n52 0.0421667
R2724 VD4.n54 VD4.n53 0.0421667
R2725 VD4.n33 VD4.n25 0.0421667
R2726 VD4.n37 VD4.n25 0.0421667
R2727 VD4.n38 VD4.n37 0.0421667
R2728 VD4.n39 VD4.n38 0.0421667
R2729 VD4.n39 VD4.n22 0.0421667
R2730 VD4.n43 VD4.n22 0.0421667
R2731 VD4.n44 VD4.n43 0.0421667
R2732 VD4.n45 VD4.n44 0.0421667
R2733 VD4.n45 VD4.n19 0.0421667
R2734 VD4.n49 VD4.n19 0.0421667
R2735 VD4.n50 VD4.n49 0.0421667
R2736 VD4.n51 VD4.n50 0.0421667
R2737 VD4.n51 VD4.n15 0.0421667
R2738 VD4.n55 VD4.n15 0.0421667
R2739 VD4.n56 VD4.n5 0.0632146
R2740 VD4.n6 VD4.n5 0.0842626
R2741 VD4.n8 VD4.n6 0.0842626
R2742 VD4.n63 VD4.n8 0.146548
R2743 VD4.n4 VD4.n2 0.0838333
R2744 VD4.n4 VD4.n3 0.0838333
R2745 VD4.n63 VD4.n0 0.0838333
R2746 V_tail_gate.n9 V_tail_gate.t13 610.534
R2747 V_tail_gate.n2 V_tail_gate.t23 610.534
R2748 V_tail_gate.n9 V_tail_gate.t21 433.8
R2749 V_tail_gate.n10 V_tail_gate.t9 433.8
R2750 V_tail_gate.n11 V_tail_gate.t17 433.8
R2751 V_tail_gate.n12 V_tail_gate.t4 433.8
R2752 V_tail_gate.n13 V_tail_gate.t11 433.8
R2753 V_tail_gate.n14 V_tail_gate.t19 433.8
R2754 V_tail_gate.n15 V_tail_gate.t16 433.8
R2755 V_tail_gate.n16 V_tail_gate.t6 433.8
R2756 V_tail_gate.n17 V_tail_gate.t14 433.8
R2757 V_tail_gate.n8 V_tail_gate.t18 433.8
R2758 V_tail_gate.n7 V_tail_gate.t5 433.8
R2759 V_tail_gate.n6 V_tail_gate.t12 433.8
R2760 V_tail_gate.n5 V_tail_gate.t20 433.8
R2761 V_tail_gate.n4 V_tail_gate.t8 433.8
R2762 V_tail_gate.n3 V_tail_gate.t7 433.8
R2763 V_tail_gate.n2 V_tail_gate.t15 433.8
R2764 V_tail_gate.n21 V_tail_gate.t22 433.8
R2765 V_tail_gate.n22 V_tail_gate.t10 433.8
R2766 V_tail_gate.n17 V_tail_gate.n16 176.733
R2767 V_tail_gate.n16 V_tail_gate.n15 176.733
R2768 V_tail_gate.n15 V_tail_gate.n14 176.733
R2769 V_tail_gate.n14 V_tail_gate.n13 176.733
R2770 V_tail_gate.n13 V_tail_gate.n12 176.733
R2771 V_tail_gate.n12 V_tail_gate.n11 176.733
R2772 V_tail_gate.n11 V_tail_gate.n10 176.733
R2773 V_tail_gate.n10 V_tail_gate.n9 176.733
R2774 V_tail_gate.n3 V_tail_gate.n2 176.733
R2775 V_tail_gate.n4 V_tail_gate.n3 176.733
R2776 V_tail_gate.n5 V_tail_gate.n4 176.733
R2777 V_tail_gate.n6 V_tail_gate.n5 176.733
R2778 V_tail_gate.n7 V_tail_gate.n6 176.733
R2779 V_tail_gate.n8 V_tail_gate.n7 176.733
R2780 V_tail_gate.n22 V_tail_gate.n21 176.733
R2781 V_tail_gate.n20 V_tail_gate.n19 163.16
R2782 V_tail_gate V_tail_gate.n23 161.925
R2783 V_tail_gate.n19 V_tail_gate.n18 49.7255
R2784 V_tail_gate.n1 V_tail_gate.n0 49.7255
R2785 V_tail_gate.n20 V_tail_gate.n17 45.5227
R2786 V_tail_gate.n23 V_tail_gate.n8 45.5227
R2787 V_tail_gate.n23 V_tail_gate.n22 45.5227
R2788 V_tail_gate.n21 V_tail_gate.n20 45.5227
R2789 V_tail_gate.n18 V_tail_gate.t3 16.0005
R2790 V_tail_gate.n18 V_tail_gate.t1 16.0005
R2791 V_tail_gate.n0 V_tail_gate.t0 16.0005
R2792 V_tail_gate.n0 V_tail_gate.t2 16.0005
R2793 V_tail_gate.n19 V_tail_gate.n1 9.563
R2794 V_tail_gate V_tail_gate.n1 1.23488
R2795 V_source.n12 V_source.t0 82.6422
R2796 V_source.n34 V_source.n33 49.3505
R2797 V_source.n32 V_source.n31 49.3505
R2798 V_source.n22 V_source.n21 49.3505
R2799 V_source.n40 V_source.n39 49.3505
R2800 V_source.n37 V_source.n36 49.3505
R2801 V_source.n49 V_source.n48 49.3505
R2802 V_source.n45 V_source.n44 49.3505
R2803 V_source.n43 V_source.n42 49.3505
R2804 V_source.n28 V_source.n27 49.3505
R2805 V_source.n24 V_source.n23 49.3505
R2806 V_source.n53 V_source.n52 32.3838
R2807 V_source.n55 V_source.n54 32.3838
R2808 V_source.n5 V_source.n4 32.3838
R2809 V_source.n11 V_source.n10 32.3838
R2810 V_source.n8 V_source.n7 32.3838
R2811 V_source.n15 V_source.n14 32.3838
R2812 V_source.n61 V_source.n60 32.3838
R2813 V_source.n64 V_source.n63 32.3838
R2814 V_source.n68 V_source.n67 32.3838
R2815 V_source.n58 V_source.n57 32.3838
R2816 V_source.n33 V_source.t30 16.0005
R2817 V_source.n33 V_source.t24 16.0005
R2818 V_source.n31 V_source.t26 16.0005
R2819 V_source.n31 V_source.t29 16.0005
R2820 V_source.n21 V_source.t25 16.0005
R2821 V_source.n21 V_source.t27 16.0005
R2822 V_source.n39 V_source.t39 16.0005
R2823 V_source.n39 V_source.t36 16.0005
R2824 V_source.n36 V_source.t40 16.0005
R2825 V_source.n36 V_source.t38 16.0005
R2826 V_source.n48 V_source.t34 16.0005
R2827 V_source.n48 V_source.t35 16.0005
R2828 V_source.n44 V_source.t32 16.0005
R2829 V_source.n44 V_source.t33 16.0005
R2830 V_source.n42 V_source.t37 16.0005
R2831 V_source.n42 V_source.t31 16.0005
R2832 V_source.n27 V_source.t22 16.0005
R2833 V_source.n27 V_source.t28 16.0005
R2834 V_source.n23 V_source.t21 16.0005
R2835 V_source.n23 V_source.t23 16.0005
R2836 V_source.n52 V_source.t8 9.6005
R2837 V_source.n52 V_source.t5 9.6005
R2838 V_source.n54 V_source.t7 9.6005
R2839 V_source.n54 V_source.t14 9.6005
R2840 V_source.n4 V_source.t20 9.6005
R2841 V_source.n4 V_source.t1 9.6005
R2842 V_source.n10 V_source.t16 9.6005
R2843 V_source.n10 V_source.t15 9.6005
R2844 V_source.n7 V_source.t2 9.6005
R2845 V_source.n7 V_source.t9 9.6005
R2846 V_source.n14 V_source.t4 9.6005
R2847 V_source.n14 V_source.t11 9.6005
R2848 V_source.n60 V_source.t10 9.6005
R2849 V_source.n60 V_source.t17 9.6005
R2850 V_source.n63 V_source.t13 9.6005
R2851 V_source.n63 V_source.t3 9.6005
R2852 V_source.n67 V_source.t18 9.6005
R2853 V_source.n67 V_source.t6 9.6005
R2854 V_source.n57 V_source.t12 9.6005
R2855 V_source.n57 V_source.t19 9.6005
R2856 V_source.n70 V_source.n5 5.85227
R2857 V_source.n56 V_source.n55 5.71925
R2858 V_source.n9 V_source.n5 5.71925
R2859 V_source.n43 V_source.n19 5.51092
R2860 V_source.n25 V_source.n22 5.51092
R2861 V_source.n46 V_source.n43 5.45883
R2862 V_source.n22 V_source.n20 5.45883
R2863 V_source.n53 V_source.n17 5.3755
R2864 V_source.n9 V_source.n8 5.3755
R2865 V_source.n16 V_source.n15 5.3755
R2866 V_source.n62 V_source.n61 5.3755
R2867 V_source.n65 V_source.n64 5.3755
R2868 V_source.n68 V_source.n66 5.3755
R2869 V_source.n58 V_source.n56 5.3755
R2870 V_source.n61 V_source.n59 5.188
R2871 V_source.n64 V_source.n6 5.188
R2872 V_source.n69 V_source.n68 5.188
R2873 V_source.n50 V_source.n49 5.16717
R2874 V_source.n45 V_source.n19 5.16717
R2875 V_source.n28 V_source.n26 5.16717
R2876 V_source.n25 V_source.n24 5.16717
R2877 V_source.n41 V_source.n40 4.89633
R2878 V_source.n49 V_source.n47 4.89633
R2879 V_source.n46 V_source.n45 4.89633
R2880 V_source.n35 V_source.n34 4.89633
R2881 V_source.n38 V_source.n37 4.89633
R2882 V_source.n29 V_source.n28 4.89633
R2883 V_source.n24 V_source.n20 4.89633
R2884 V_source.n32 V_source.n30 4.89633
R2885 V_source.n13 V_source.n12 4.5005
R2886 V_source.n38 V_source.n35 3.6255
R2887 V_source.n51 V_source.n18 2.2076
R2888 V_source.n0 V_source.n51 2.16822
R2889 V_source.n18 V_source.n2 2.16822
R2890 V_source.n59 V_source.n1 2.02255
R2891 V_source.n3 V_source.n70 1.36007
R2892 V_source.n12 V_source.n11 0.8755
R2893 V_source.n70 V_source.n69 0.664374
R2894 V_source.n1 V_source.n53 0.6255
R2895 V_source.n1 V_source.n55 0.6255
R2896 V_source.n15 V_source.n3 0.6255
R2897 V_source.n8 V_source.n3 0.6255
R2898 V_source.n11 V_source.n3 0.6255
R2899 V_source.n1 V_source.n58 0.6255
R2900 V_source.n37 V_source.n0 0.604667
R2901 V_source.n40 V_source.n0 0.604667
R2902 V_source.n2 V_source.n32 0.604667
R2903 V_source.n34 V_source.n2 0.604667
R2904 V_source.n47 V_source.n46 0.563
R2905 V_source.n47 V_source.n41 0.563
R2906 V_source.n41 V_source.n38 0.563
R2907 V_source.n35 V_source.n30 0.563
R2908 V_source.n29 V_source.n20 0.563
R2909 V_source.n30 V_source.n29 0.563
R2910 V_source.n26 V_source.n18 0.510302
R2911 V_source.n51 V_source.n50 0.510302
R2912 V_source.n26 V_source.n25 0.34425
R2913 V_source.n50 V_source.n19 0.34425
R2914 V_source.n69 V_source.n6 0.34425
R2915 V_source.n59 V_source.n6 0.34425
R2916 V_source.n13 V_source.n9 0.34425
R2917 V_source.n16 V_source.n13 0.34425
R2918 V_source.n66 V_source.n16 0.34425
R2919 V_source.n66 V_source.n65 0.34425
R2920 V_source.n65 V_source.n62 0.34425
R2921 V_source.n62 V_source.n17 0.34425
R2922 V_source.n56 V_source.n17 0.34425
R2923 V_source.n1 V_source.n0 0.267327
R2924 V_source V_source.n2 0.226462
R2925 V_source V_source.n3 0.0413654
R2926 VD1.n15 VD1.n14 49.3505
R2927 VD1.n18 VD1.n17 49.3505
R2928 VD1.n4 VD1.n3 49.3505
R2929 VD1.n43 VD1.n42 49.3505
R2930 VD1.n9 VD1.n8 49.3505
R2931 VD1.n12 VD1.n11 49.3505
R2932 VD1.n25 VD1.n24 49.3505
R2933 VD1.n28 VD1.n27 49.3505
R2934 VD1.n32 VD1.n31 49.3505
R2935 VD1.n7 VD1.n6 49.3505
R2936 VD1.n39 VD1.n38 49.3505
R2937 VD1.n14 VD1.t7 16.0005
R2938 VD1.n14 VD1.t12 16.0005
R2939 VD1.n17 VD1.t16 16.0005
R2940 VD1.n17 VD1.t10 16.0005
R2941 VD1.n3 VD1.t17 16.0005
R2942 VD1.n3 VD1.t11 16.0005
R2943 VD1.n42 VD1.t15 16.0005
R2944 VD1.n42 VD1.t9 16.0005
R2945 VD1.n8 VD1.t2 16.0005
R2946 VD1.n8 VD1.t21 16.0005
R2947 VD1.n11 VD1.t20 16.0005
R2948 VD1.n11 VD1.t5 16.0005
R2949 VD1.n24 VD1.t1 16.0005
R2950 VD1.n24 VD1.t6 16.0005
R2951 VD1.n27 VD1.t19 16.0005
R2952 VD1.n27 VD1.t3 16.0005
R2953 VD1.n31 VD1.t0 16.0005
R2954 VD1.n31 VD1.t4 16.0005
R2955 VD1.n6 VD1.t13 16.0005
R2956 VD1.n6 VD1.t8 16.0005
R2957 VD1.n38 VD1.t14 16.0005
R2958 VD1.n38 VD1.t18 16.0005
R2959 VD1.n23 VD1.n13 6.2505
R2960 VD1.n33 VD1.n2 6.2505
R2961 VD1.n21 VD1.n20 6.2505
R2962 VD1.n36 VD1.n35 6.2505
R2963 VD1.n26 VD1.n12 5.6255
R2964 VD1.n30 VD1.n9 5.6255
R2965 VD1.n40 VD1.n7 5.438
R2966 VD1.n16 VD1.n15 5.438
R2967 VD1.n36 VD1.n7 5.31821
R2968 VD1.n20 VD1.n15 5.31821
R2969 VD1.n19 VD1.n18 5.08383
R2970 VD1.n4 VD1.n1 5.08383
R2971 VD1.n44 VD1.n43 5.08383
R2972 VD1.n39 VD1.n37 5.08383
R2973 VD1.n26 VD1.n25 5.063
R2974 VD1.n29 VD1.n28 5.063
R2975 VD1.n32 VD1.n30 5.063
R2976 VD1.n35 VD1.n34 5.063
R2977 VD1.n22 VD1.n21 5.063
R2978 VD1.n18 VD1.n16 4.8755
R2979 VD1.n5 VD1.n4 4.8755
R2980 VD1.n43 VD1.n41 4.8755
R2981 VD1.n40 VD1.n39 4.8755
R2982 VD1 VD1.n45 4.60467
R2983 VD1.n34 VD1.n33 4.5005
R2984 VD1.n10 VD1.n0 4.5005
R2985 VD1.n23 VD1.n22 4.5005
R2986 VD1 VD1.n0 1.64633
R2987 VD1.n34 VD1.n10 0.563
R2988 VD1.n22 VD1.n10 0.563
R2989 VD1.n29 VD1.n26 0.563
R2990 VD1.n30 VD1.n29 0.563
R2991 VD1.n16 VD1.n5 0.563
R2992 VD1.n41 VD1.n5 0.563
R2993 VD1.n41 VD1.n40 0.563
R2994 VD1.n25 VD1.n23 0.3755
R2995 VD1.n28 VD1.n0 0.3755
R2996 VD1.n33 VD1.n32 0.3755
R2997 VD1.n21 VD1.n12 0.3755
R2998 VD1.n35 VD1.n9 0.3755
R2999 VD1.n37 VD1.n36 0.234875
R3000 VD1.n37 VD1.n2 0.234875
R3001 VD1.n44 VD1.n2 0.234875
R3002 VD1.n45 VD1.n44 0.234875
R3003 VD1.n45 VD1.n1 0.234875
R3004 VD1.n13 VD1.n1 0.234875
R3005 VD1.n19 VD1.n13 0.234875
R3006 VD1.n20 VD1.n19 0.234875
R3007 Vb2.n3 Vb2.t13 751.226
R3008 Vb2.n1 Vb2.t0 721.625
R3009 Vb2.n17 Vb2.t14 611.739
R3010 Vb2.n13 Vb2.t22 611.739
R3011 Vb2.n8 Vb2.t8 611.739
R3012 Vb2.n4 Vb2.t23 611.739
R3013 Vb2.n2 Vb2.t17 563.451
R3014 Vb2.n17 Vb2.t10 421.75
R3015 Vb2.n18 Vb2.t6 421.75
R3016 Vb2.n19 Vb2.t19 421.75
R3017 Vb2.n20 Vb2.t15 421.75
R3018 Vb2.n13 Vb2.t4 421.75
R3019 Vb2.n14 Vb2.t9 421.75
R3020 Vb2.n15 Vb2.t12 421.75
R3021 Vb2.n16 Vb2.t18 421.75
R3022 Vb2.n8 Vb2.t3 421.75
R3023 Vb2.n9 Vb2.t21 421.75
R3024 Vb2.n10 Vb2.t20 421.75
R3025 Vb2.n11 Vb2.t16 421.75
R3026 Vb2.n4 Vb2.t5 421.75
R3027 Vb2.n5 Vb2.t24 421.75
R3028 Vb2.n6 Vb2.t7 421.75
R3029 Vb2.n7 Vb2.t11 421.75
R3030 Vb2.n22 Vb2.n12 313.776
R3031 Vb2.n22 Vb2.n21 313.212
R3032 Vb2.n18 Vb2.n17 167.094
R3033 Vb2.n19 Vb2.n18 167.094
R3034 Vb2.n20 Vb2.n19 167.094
R3035 Vb2.n14 Vb2.n13 167.094
R3036 Vb2.n15 Vb2.n14 167.094
R3037 Vb2.n16 Vb2.n15 167.094
R3038 Vb2.n9 Vb2.n8 167.094
R3039 Vb2.n10 Vb2.n9 167.094
R3040 Vb2.n11 Vb2.n10 167.094
R3041 Vb2.n5 Vb2.n4 167.094
R3042 Vb2.n6 Vb2.n5 167.094
R3043 Vb2.n7 Vb2.n6 167.094
R3044 Vb2.n1 Vb2.n0 67.013
R3045 Vb2.n21 Vb2.n20 35.3472
R3046 Vb2.n21 Vb2.n16 35.3472
R3047 Vb2.n12 Vb2.n11 35.3472
R3048 Vb2.n12 Vb2.n7 35.3472
R3049 Vb2.n0 Vb2.t1 11.2576
R3050 Vb2.n0 Vb2.t2 11.2576
R3051 Vb2.n23 Vb2.n3 10.0005
R3052 Vb2.n2 Vb2.n1 7.35988
R3053 Vb2.n23 Vb2.n22 4.5005
R3054 Vb2.n3 Vb2.n2 1.14112
R3055 Vb2 Vb2.n23 0.063
R3056 VD3.n53 VD3.t3 672.293
R3057 VD3.n56 VD3.t0 672.293
R3058 VD3.t4 VD3.n54 213.131
R3059 VD3.n55 VD3.t1 213.131
R3060 VD3.t28 VD3.t4 146.155
R3061 VD3.t34 VD3.t28 146.155
R3062 VD3.t20 VD3.t34 146.155
R3063 VD3.t22 VD3.t20 146.155
R3064 VD3.t24 VD3.t22 146.155
R3065 VD3.t26 VD3.t24 146.155
R3066 VD3.t30 VD3.t26 146.155
R3067 VD3.t16 VD3.t30 146.155
R3068 VD3.t32 VD3.t16 146.155
R3069 VD3.t18 VD3.t32 146.155
R3070 VD3.t1 VD3.t18 146.155
R3071 VD3.n54 VD3.t5 76.2576
R3072 VD3.n55 VD3.t2 76.2576
R3073 VD3.n72 VD3.n4 66.9922
R3074 VD3.n6 VD3.n5 66.9922
R3075 VD3.n64 VD3.n8 66.9922
R3076 VD3.n59 VD3.n58 66.9922
R3077 VD3.n78 VD3.n77 66.9922
R3078 VD3.n18 VD3.n17 66.0338
R3079 VD3.n34 VD3.n33 66.0338
R3080 VD3.n43 VD3.n42 66.0338
R3081 VD3.n46 VD3.n45 66.0338
R3082 VD3.n22 VD3.n21 66.0338
R3083 VD3.n25 VD3.n24 66.0338
R3084 VD3.n4 VD3.t21 11.2576
R3085 VD3.n4 VD3.t23 11.2576
R3086 VD3.n5 VD3.t25 11.2576
R3087 VD3.n5 VD3.t27 11.2576
R3088 VD3.n8 VD3.t31 11.2576
R3089 VD3.n8 VD3.t17 11.2576
R3090 VD3.n58 VD3.t33 11.2576
R3091 VD3.n58 VD3.t19 11.2576
R3092 VD3.n17 VD3.t8 11.2576
R3093 VD3.n17 VD3.t10 11.2576
R3094 VD3.n33 VD3.t9 11.2576
R3095 VD3.n33 VD3.t12 11.2576
R3096 VD3.n42 VD3.t14 11.2576
R3097 VD3.n42 VD3.t15 11.2576
R3098 VD3.n45 VD3.t6 11.2576
R3099 VD3.n45 VD3.t36 11.2576
R3100 VD3.n21 VD3.t13 11.2576
R3101 VD3.n21 VD3.t7 11.2576
R3102 VD3.n24 VD3.t37 11.2576
R3103 VD3.n24 VD3.t11 11.2576
R3104 VD3.n78 VD3.t29 11.2576
R3105 VD3.t35 VD3.n78 11.2576
R3106 VD3.n46 VD3.n44 5.91717
R3107 VD3.n25 VD3.n23 5.91717
R3108 VD3.n34 VD3.n13 5.29217
R3109 VD3.n44 VD3.n43 5.29217
R3110 VD3.n23 VD3.n22 5.29217
R3111 VD3.n20 VD3.n18 5.29217
R3112 VD3.n31 VD3.n30 1.5005
R3113 VD3.n29 VD3.n16 1.5005
R3114 VD3.n28 VD3.n27 1.5005
R3115 VD3.n48 VD3.n47 1.5005
R3116 VD3.n12 VD3.n11 1.5005
R3117 VD3.n39 VD3.n15 1.5005
R3118 VD3.n41 VD3.n40 1.5005
R3119 VD3.n38 VD3.n14 1.5005
R3120 VD3.n37 VD3.n36 1.5005
R3121 VD3.n35 VD3.n32 1.5005
R3122 VD3.n61 VD3.n60 1.5005
R3123 VD3.n62 VD3.n9 1.5005
R3124 VD3.n64 VD3.n63 1.5005
R3125 VD3.n65 VD3.n7 1.5005
R3126 VD3.n67 VD3.n66 1.5005
R3127 VD3.n68 VD3.n6 1.5005
R3128 VD3.n70 VD3.n69 1.5005
R3129 VD3.n71 VD3.n3 1.5005
R3130 VD3.n73 VD3.n72 1.5005
R3131 VD3.n74 VD3.n2 1.5005
R3132 VD3.n76 VD3.n75 1.5005
R3133 VD3.n77 VD3.n1 1.5005
R3134 VD3.n49 VD3.n0 1.5005
R3135 VD3.n50 VD3.n10 1.5005
R3136 VD3.n52 VD3.n51 1.5005
R3137 VD3.n54 VD3.n53 1.03383
R3138 VD3.n56 VD3.n55 1.03383
R3139 VD3.n57 VD3.n56 1.02405
R3140 VD3.n26 VD3.n25 1.02322
R3141 VD3.n53 VD3.n52 0.958833
R3142 VD3.n35 VD3.n34 0.958833
R3143 VD3.n43 VD3.n41 0.958833
R3144 VD3.n47 VD3.n46 0.958833
R3145 VD3.n22 VD3.n19 0.958833
R3146 VD3.n30 VD3.n18 0.958833
R3147 VD3.n51 VD3.n48 0.786958
R3148 VD3.n44 VD3.n13 0.6255
R3149 VD3.n20 VD3.n13 0.6255
R3150 VD3.n23 VD3.n20 0.6255
R3151 VD3.n27 VD3.n26 0.427973
R3152 VD3.n61 VD3.n57 0.427925
R3153 VD3.n32 VD3.n31 0.1255
R3154 VD3.n59 VD3.n57 0.0588743
R3155 VD3.n26 VD3.n19 0.0587394
R3156 VD3.n36 VD3.n35 0.0421667
R3157 VD3.n36 VD3.n14 0.0421667
R3158 VD3.n41 VD3.n14 0.0421667
R3159 VD3.n41 VD3.n15 0.0421667
R3160 VD3.n15 VD3.n12 0.0421667
R3161 VD3.n47 VD3.n12 0.0421667
R3162 VD3.n28 VD3.n19 0.0421667
R3163 VD3.n29 VD3.n28 0.0421667
R3164 VD3.n30 VD3.n29 0.0421667
R3165 VD3.n27 VD3.n16 0.0421667
R3166 VD3.n31 VD3.n16 0.0421667
R3167 VD3.n37 VD3.n32 0.0421667
R3168 VD3.n38 VD3.n37 0.0421667
R3169 VD3.n40 VD3.n38 0.0421667
R3170 VD3.n40 VD3.n39 0.0421667
R3171 VD3.n39 VD3.n11 0.0421667
R3172 VD3.n48 VD3.n11 0.0421667
R3173 VD3.n51 VD3.n50 0.0421667
R3174 VD3.n50 VD3.n49 0.0421667
R3175 VD3.n49 VD3.n1 0.0421667
R3176 VD3.n75 VD3.n1 0.0421667
R3177 VD3.n75 VD3.n74 0.0421667
R3178 VD3.n74 VD3.n73 0.0421667
R3179 VD3.n73 VD3.n3 0.0421667
R3180 VD3.n69 VD3.n3 0.0421667
R3181 VD3.n69 VD3.n68 0.0421667
R3182 VD3.n68 VD3.n67 0.0421667
R3183 VD3.n67 VD3.n7 0.0421667
R3184 VD3.n63 VD3.n7 0.0421667
R3185 VD3.n63 VD3.n62 0.0421667
R3186 VD3.n62 VD3.n61 0.0421667
R3187 VD3.n52 VD3.n10 0.0421667
R3188 VD3.n10 VD3.n0 0.0421667
R3189 VD3.n77 VD3.n0 0.0421667
R3190 VD3.n77 VD3.n76 0.0421667
R3191 VD3.n76 VD3.n2 0.0421667
R3192 VD3.n72 VD3.n2 0.0421667
R3193 VD3.n72 VD3.n71 0.0421667
R3194 VD3.n71 VD3.n70 0.0421667
R3195 VD3.n70 VD3.n6 0.0421667
R3196 VD3.n66 VD3.n6 0.0421667
R3197 VD3.n66 VD3.n65 0.0421667
R3198 VD3.n65 VD3.n64 0.0421667
R3199 VD3.n64 VD3.n9 0.0421667
R3200 VD3.n60 VD3.n9 0.0421667
R3201 VD3.n60 VD3.n59 0.0421667
R3202 V_err_amp_ref.n0 V_err_amp_ref.t1 651.405
R3203 V_err_amp_ref.n0 V_err_amp_ref.t0 648.03
R3204 V_err_amp_ref V_err_amp_ref.n0 1.53175
R3205 V_err_gate.n5 V_err_gate.t4 479.322
R3206 V_err_gate.n5 V_err_gate.t6 479.322
R3207 V_err_gate.n1 V_err_gate.t5 479.322
R3208 V_err_gate.n1 V_err_gate.t7 479.322
R3209 V_err_gate.n2 V_err_gate.n0 178.627
R3210 V_err_gate.n4 V_err_gate.n3 177.987
R3211 V_err_gate.n6 V_err_gate.n5 165.8
R3212 V_err_gate.n2 V_err_gate.n1 165.8
R3213 V_err_gate.n3 V_err_gate.t1 15.7605
R3214 V_err_gate.n3 V_err_gate.t3 15.7605
R3215 V_err_gate.n0 V_err_gate.t0 15.7605
R3216 V_err_gate.n0 V_err_gate.t2 15.7605
R3217 V_err_gate.n6 V_err_gate.n4 1.70362
R3218 V_err_gate.n4 V_err_gate.n2 0.641125
R3219 V_err_gate V_err_gate.n6 0.063
R3220 V_err_mir_p V_err_mir_p.n0 187.315
R3221 V_err_mir_p V_err_mir_p.n1 177.755
R3222 V_err_mir_p.n0 V_err_mir_p.t3 15.7605
R3223 V_err_mir_p.n0 V_err_mir_p.t0 15.7605
R3224 V_err_mir_p.n1 V_err_mir_p.t1 15.7605
R3225 V_err_mir_p.n1 V_err_mir_p.t2 15.7605
R3226 err_amp_mir.n1 err_amp_mir.t5 573.044
R3227 err_amp_mir.n1 err_amp_mir.t0 433.8
R3228 err_amp_mir.n2 err_amp_mir.n0 184.643
R3229 err_amp_mir.n2 err_amp_mir.n1 163.978
R3230 err_amp_mir.n3 err_amp_mir.n2 33.0088
R3231 err_amp_mir.n0 err_amp_mir.t4 15.7605
R3232 err_amp_mir.n0 err_amp_mir.t3 15.7605
R3233 err_amp_mir.t1 err_amp_mir.n3 9.6005
R3234 err_amp_mir.n3 err_amp_mir.t2 9.6005
R3235 VD2.n15 VD2.n14 49.3505
R3236 VD2.n9 VD2.n8 49.3505
R3237 VD2.n12 VD2.n11 49.3505
R3238 VD2.n25 VD2.n24 49.3505
R3239 VD2.n28 VD2.n27 49.3505
R3240 VD2.n32 VD2.n31 49.3505
R3241 VD2.n7 VD2.n6 49.3505
R3242 VD2.n39 VD2.n38 49.3505
R3243 VD2.n43 VD2.n42 49.3505
R3244 VD2.n4 VD2.n3 49.3505
R3245 VD2.n18 VD2.n17 49.3505
R3246 VD2.n14 VD2.t9 16.0005
R3247 VD2.n14 VD2.t14 16.0005
R3248 VD2.n8 VD2.t3 16.0005
R3249 VD2.n8 VD2.t6 16.0005
R3250 VD2.n11 VD2.t2 16.0005
R3251 VD2.n11 VD2.t5 16.0005
R3252 VD2.n24 VD2.t20 16.0005
R3253 VD2.n24 VD2.t0 16.0005
R3254 VD2.n27 VD2.t1 16.0005
R3255 VD2.n27 VD2.t4 16.0005
R3256 VD2.n31 VD2.t21 16.0005
R3257 VD2.n31 VD2.t7 16.0005
R3258 VD2.n6 VD2.t16 16.0005
R3259 VD2.n6 VD2.t8 16.0005
R3260 VD2.n38 VD2.t17 16.0005
R3261 VD2.n38 VD2.t11 16.0005
R3262 VD2.n42 VD2.t18 16.0005
R3263 VD2.n42 VD2.t12 16.0005
R3264 VD2.n3 VD2.t10 16.0005
R3265 VD2.n3 VD2.t15 16.0005
R3266 VD2.n17 VD2.t19 16.0005
R3267 VD2.n17 VD2.t13 16.0005
R3268 VD2.n23 VD2.n13 6.2505
R3269 VD2.n33 VD2.n2 6.2505
R3270 VD2.n21 VD2.n20 6.2505
R3271 VD2.n36 VD2.n35 6.2505
R3272 VD2.n26 VD2.n12 5.6255
R3273 VD2.n30 VD2.n9 5.6255
R3274 VD2.n40 VD2.n7 5.438
R3275 VD2.n16 VD2.n15 5.438
R3276 VD2.n36 VD2.n7 5.31821
R3277 VD2.n20 VD2.n15 5.31821
R3278 VD2.n19 VD2.n18 5.08383
R3279 VD2.n39 VD2.n37 5.08383
R3280 VD2.n44 VD2.n43 5.08383
R3281 VD2.n4 VD2.n1 5.08383
R3282 VD2.n26 VD2.n25 5.063
R3283 VD2.n29 VD2.n28 5.063
R3284 VD2.n32 VD2.n30 5.063
R3285 VD2.n35 VD2.n34 5.063
R3286 VD2.n22 VD2.n21 5.063
R3287 VD2.n40 VD2.n39 4.8755
R3288 VD2.n43 VD2.n41 4.8755
R3289 VD2.n5 VD2.n4 4.8755
R3290 VD2.n18 VD2.n16 4.8755
R3291 VD2 VD2.n45 4.60467
R3292 VD2.n34 VD2.n33 4.5005
R3293 VD2.n10 VD2.n0 4.5005
R3294 VD2.n23 VD2.n22 4.5005
R3295 VD2 VD2.n0 1.64633
R3296 VD2.n34 VD2.n10 0.563
R3297 VD2.n22 VD2.n10 0.563
R3298 VD2.n29 VD2.n26 0.563
R3299 VD2.n30 VD2.n29 0.563
R3300 VD2.n16 VD2.n5 0.563
R3301 VD2.n41 VD2.n5 0.563
R3302 VD2.n41 VD2.n40 0.563
R3303 VD2.n25 VD2.n23 0.3755
R3304 VD2.n28 VD2.n0 0.3755
R3305 VD2.n33 VD2.n32 0.3755
R3306 VD2.n21 VD2.n12 0.3755
R3307 VD2.n35 VD2.n9 0.3755
R3308 VD2.n37 VD2.n36 0.234875
R3309 VD2.n37 VD2.n2 0.234875
R3310 VD2.n44 VD2.n2 0.234875
R3311 VD2.n45 VD2.n44 0.234875
R3312 VD2.n45 VD2.n1 0.234875
R3313 VD2.n13 VD2.n1 0.234875
R3314 VD2.n19 VD2.n13 0.234875
R3315 VD2.n20 VD2.n19 0.234875
R3316 Y.n74 Y.t42 1172.87
R3317 Y.n70 Y.t39 1172.87
R3318 Y.n74 Y.t26 996.134
R3319 Y.n75 Y.t45 996.134
R3320 Y.n76 Y.t38 996.134
R3321 Y.n77 Y.t48 996.134
R3322 Y.n73 Y.t31 996.134
R3323 Y.n72 Y.t51 996.134
R3324 Y.n71 Y.t35 996.134
R3325 Y.n70 Y.t53 996.134
R3326 Y.n46 Y.t37 690.867
R3327 Y.n39 Y.t33 690.867
R3328 Y.n55 Y.t40 530.201
R3329 Y.n48 Y.t36 530.201
R3330 Y.n46 Y.t54 514.134
R3331 Y.n39 Y.t50 514.134
R3332 Y.n40 Y.t29 514.134
R3333 Y.n41 Y.t47 514.134
R3334 Y.n42 Y.t27 514.134
R3335 Y.n43 Y.t44 514.134
R3336 Y.n44 Y.t30 514.134
R3337 Y.n45 Y.t41 514.134
R3338 Y.n55 Y.t25 353.467
R3339 Y.n54 Y.t43 353.467
R3340 Y.n53 Y.t34 353.467
R3341 Y.n52 Y.t46 353.467
R3342 Y.n51 Y.t28 353.467
R3343 Y.n50 Y.t49 353.467
R3344 Y.n49 Y.t32 353.467
R3345 Y.n48 Y.t52 353.467
R3346 Y.n73 Y.n72 176.733
R3347 Y.n72 Y.n71 176.733
R3348 Y.n71 Y.n70 176.733
R3349 Y.n75 Y.n74 176.733
R3350 Y.n76 Y.n75 176.733
R3351 Y.n77 Y.n76 176.733
R3352 Y.n54 Y.n53 176.733
R3353 Y.n53 Y.n52 176.733
R3354 Y.n52 Y.n51 176.733
R3355 Y.n51 Y.n50 176.733
R3356 Y.n50 Y.n49 176.733
R3357 Y.n49 Y.n48 176.733
R3358 Y.n45 Y.n44 176.733
R3359 Y.n44 Y.n43 176.733
R3360 Y.n43 Y.n42 176.733
R3361 Y.n42 Y.n41 176.733
R3362 Y.n41 Y.n40 176.733
R3363 Y.n40 Y.n39 176.733
R3364 Y.n57 Y.n56 165.472
R3365 Y.n57 Y.n47 165.472
R3366 Y.n80 Y.n79 152
R3367 Y.n81 Y.n80 131.571
R3368 Y.n80 Y.n78 124.517
R3369 Y.n147 Y.n57 74.5372
R3370 Y.n107 Y.n106 66.0338
R3371 Y.n98 Y.n97 66.0338
R3372 Y.n96 Y.n95 66.0338
R3373 Y.n101 Y.n100 66.0338
R3374 Y.n104 Y.n103 66.0338
R3375 Y.n110 Y.n109 66.0338
R3376 Y.n7 Y.n6 49.3505
R3377 Y.n11 Y.n10 49.3505
R3378 Y.n20 Y.n19 49.3505
R3379 Y.n30 Y.n29 49.3505
R3380 Y.n26 Y.n25 49.3505
R3381 Y.n23 Y.n22 49.3505
R3382 Y.n64 Y.t6 41.0384
R3383 Y.n78 Y.n73 40.1672
R3384 Y.n78 Y.n77 40.1672
R3385 Y.n56 Y.n54 40.1672
R3386 Y.n56 Y.n55 40.1672
R3387 Y.n47 Y.n45 40.1672
R3388 Y.n47 Y.n46 40.1672
R3389 Y.n82 Y.n81 16.3217
R3390 Y.n6 Y.t7 16.0005
R3391 Y.n6 Y.t20 16.0005
R3392 Y.n10 Y.t19 16.0005
R3393 Y.n10 Y.t2 16.0005
R3394 Y.n19 Y.t5 16.0005
R3395 Y.n19 Y.t23 16.0005
R3396 Y.n29 Y.t0 16.0005
R3397 Y.n29 Y.t1 16.0005
R3398 Y.n25 Y.t4 16.0005
R3399 Y.n25 Y.t24 16.0005
R3400 Y.n22 Y.t8 16.0005
R3401 Y.n22 Y.t3 16.0005
R3402 Y.n79 Y.n69 12.8005
R3403 Y.n106 Y.t9 11.2576
R3404 Y.n106 Y.t21 11.2576
R3405 Y.n97 Y.t22 11.2576
R3406 Y.n97 Y.t13 11.2576
R3407 Y.n95 Y.t15 11.2576
R3408 Y.n95 Y.t17 11.2576
R3409 Y.n100 Y.t10 11.2576
R3410 Y.n100 Y.t12 11.2576
R3411 Y.n103 Y.t11 11.2576
R3412 Y.n103 Y.t14 11.2576
R3413 Y.n109 Y.t16 11.2576
R3414 Y.n109 Y.t18 11.2576
R3415 Y.n79 Y.n67 9.36264
R3416 Y.n69 Y.n68 9.3005
R3417 Y.n99 Y.n98 5.91717
R3418 Y.n108 Y.n107 5.91717
R3419 Y.n21 Y.n11 5.6255
R3420 Y.n24 Y.n7 5.6255
R3421 Y.n81 Y.n69 5.33141
R3422 Y.n99 Y.n96 5.29217
R3423 Y.n102 Y.n101 5.29217
R3424 Y.n105 Y.n104 5.29217
R3425 Y.n110 Y.n108 5.29217
R3426 Y.n112 Y.n86 5.1255
R3427 Y.n115 Y.n94 5.1255
R3428 Y.n21 Y.n20 5.063
R3429 Y.n30 Y.n28 5.063
R3430 Y.n27 Y.n26 5.063
R3431 Y.n24 Y.n23 5.063
R3432 Y.n35 Y.n34 5.063
R3433 Y.n12 Y.n8 5.063
R3434 Y.n112 Y.n111 4.5005
R3435 Y.n113 Y.n89 4.5005
R3436 Y.n114 Y.n92 4.5005
R3437 Y.n116 Y.n115 4.5005
R3438 Y.n141 Y.n140 4.5005
R3439 Y.n34 Y.n5 4.5005
R3440 Y.n33 Y.n1 4.5005
R3441 Y.n32 Y.n31 4.5005
R3442 Y.n18 Y.n8 4.5005
R3443 Y.n148 Y.n36 4.5005
R3444 Y.n147 Y.n146 4.5005
R3445 Y.n148 Y.n147 4.5005
R3446 Y.n83 Y.n82 4.5005
R3447 Y.n61 Y.n60 4.5005
R3448 Y.n62 Y.n59 2.26187
R3449 Y.n138 Y.n84 2.26187
R3450 Y.n139 Y.n138 2.26187
R3451 Y.n63 Y.n62 2.26187
R3452 Y.n142 Y.n137 2.24063
R3453 Y.n143 Y.n84 2.24063
R3454 Y.n146 Y.n145 2.24063
R3455 Y.n58 Y.n38 2.24063
R3456 Y.n66 Y.n59 2.24063
R3457 Y.n144 Y.n37 2.24063
R3458 Y.n65 Y.n64 2.24063
R3459 Y.n83 Y.n67 2.22018
R3460 Y.n136 Y.n135 1.5005
R3461 Y.n134 Y.n85 1.5005
R3462 Y.n133 Y.n132 1.5005
R3463 Y.n131 Y.n87 1.5005
R3464 Y.n130 Y.n129 1.5005
R3465 Y.n128 Y.n88 1.5005
R3466 Y.n127 Y.n126 1.5005
R3467 Y.n125 Y.n90 1.5005
R3468 Y.n124 Y.n123 1.5005
R3469 Y.n122 Y.n91 1.5005
R3470 Y.n121 Y.n120 1.5005
R3471 Y.n119 Y.n93 1.5005
R3472 Y.n150 Y.n149 1.5005
R3473 Y.n151 Y.n4 1.5005
R3474 Y.n153 Y.n152 1.5005
R3475 Y.n154 Y.n2 1.5005
R3476 Y.n156 Y.n155 1.5005
R3477 Y.n3 Y.n0 1.5005
R3478 Y.n14 Y.n9 1.5005
R3479 Y.n16 Y.n15 1.5005
R3480 Y.n13 Y.n12 1.43397
R3481 Y.n18 Y.n17 1.3755
R3482 Y.n31 Y.n9 1.3755
R3483 Y.n156 Y.n1 1.3755
R3484 Y.n152 Y.n5 1.3755
R3485 Y.n150 Y.n35 1.3755
R3486 Y.n144 Y.n143 0.979667
R3487 Y.n116 Y.n96 0.792167
R3488 Y.n101 Y.n92 0.792167
R3489 Y.n104 Y.n89 0.792167
R3490 Y.n111 Y.n110 0.792167
R3491 Y.n98 Y.n94 0.792167
R3492 Y.n107 Y.n86 0.792167
R3493 Y.n83 Y.n66 0.682792
R3494 Y.n149 Y.n148 0.630708
R3495 Y.n113 Y.n112 0.6255
R3496 Y.n114 Y.n113 0.6255
R3497 Y.n115 Y.n114 0.6255
R3498 Y.n102 Y.n99 0.6255
R3499 Y.n105 Y.n102 0.6255
R3500 Y.n108 Y.n105 0.6255
R3501 Y.n137 Y.n136 0.609875
R3502 Y.n15 Y.n13 0.564601
R3503 Y.n34 Y.n33 0.563
R3504 Y.n33 Y.n32 0.563
R3505 Y.n32 Y.n8 0.563
R3506 Y.n28 Y.n21 0.563
R3507 Y.n28 Y.n27 0.563
R3508 Y.n27 Y.n24 0.563
R3509 Y.n118 Y.n94 0.533638
R3510 Y.n117 Y.n116 0.46925
R3511 Y.n122 Y.n92 0.46925
R3512 Y.n127 Y.n89 0.46925
R3513 Y.n111 Y.n87 0.46925
R3514 Y.n135 Y.n86 0.46925
R3515 Y.n146 Y.n83 0.46925
R3516 Y.n119 Y.n118 0.427973
R3517 Y.n20 Y.n18 0.3755
R3518 Y.n31 Y.n30 0.3755
R3519 Y.n26 Y.n1 0.3755
R3520 Y.n23 Y.n5 0.3755
R3521 Y.n12 Y.n11 0.3755
R3522 Y.n35 Y.n7 0.3755
R3523 Y.n82 Y.n68 0.1255
R3524 Y.n68 Y.n67 0.0626438
R3525 Y.n118 Y.n117 0.0587394
R3526 Y.n17 Y.n16 0.0577917
R3527 Y.n16 Y.n9 0.0577917
R3528 Y.n9 Y.n0 0.0577917
R3529 Y.n156 Y.n2 0.0577917
R3530 Y.n152 Y.n2 0.0577917
R3531 Y.n152 Y.n151 0.0577917
R3532 Y.n151 Y.n150 0.0577917
R3533 Y.n15 Y.n14 0.0577917
R3534 Y.n14 Y.n3 0.0577917
R3535 Y.n155 Y.n3 0.0577917
R3536 Y.n155 Y.n154 0.0577917
R3537 Y.n154 Y.n153 0.0577917
R3538 Y.n153 Y.n4 0.0577917
R3539 Y.n149 Y.n4 0.0577917
R3540 Y.n17 Y.n13 0.054517
R3541 Y.n117 Y.n93 0.0421667
R3542 Y.n121 Y.n93 0.0421667
R3543 Y.n122 Y.n121 0.0421667
R3544 Y.n123 Y.n122 0.0421667
R3545 Y.n123 Y.n90 0.0421667
R3546 Y.n127 Y.n90 0.0421667
R3547 Y.n128 Y.n127 0.0421667
R3548 Y.n129 Y.n128 0.0421667
R3549 Y.n129 Y.n87 0.0421667
R3550 Y.n133 Y.n87 0.0421667
R3551 Y.n134 Y.n133 0.0421667
R3552 Y.n135 Y.n134 0.0421667
R3553 Y.n120 Y.n119 0.0421667
R3554 Y.n120 Y.n91 0.0421667
R3555 Y.n124 Y.n91 0.0421667
R3556 Y.n125 Y.n124 0.0421667
R3557 Y.n126 Y.n125 0.0421667
R3558 Y.n126 Y.n88 0.0421667
R3559 Y.n130 Y.n88 0.0421667
R3560 Y.n131 Y.n130 0.0421667
R3561 Y.n132 Y.n131 0.0421667
R3562 Y.n132 Y.n85 0.0421667
R3563 Y.n136 Y.n85 0.0421667
R3564 Y.n146 Y.n58 0.0421667
R3565 Y Y.n0 0.0369583
R3566 Y.n142 Y.n141 0.0217373
R3567 Y.n145 Y.n144 0.0217373
R3568 Y.n147 Y.n38 0.0217373
R3569 Y.n140 Y.n84 0.0217373
R3570 Y.n143 Y.n142 0.0217373
R3571 Y.n145 Y.n36 0.0217373
R3572 Y.n38 Y.n36 0.0217373
R3573 Y.n61 Y.n59 0.0217373
R3574 Y.n62 Y.n60 0.0217373
R3575 Y.n140 Y.n139 0.0217373
R3576 Y.n141 Y.n138 0.0217373
R3577 Y.n139 Y.n137 0.0217373
R3578 Y.n148 Y.n37 0.0217373
R3579 Y.n65 Y.n60 0.0217373
R3580 Y.n58 Y.n37 0.0217373
R3581 Y.n63 Y.n61 0.0217373
R3582 Y.n64 Y.n63 0.0217373
R3583 Y.n66 Y.n65 0.0217373
R3584 Y Y.n156 0.0213333
R3585 V_CMFB_S3 V_CMFB_S3.t0 126.431
R3586 V_CMFB_S3.n3 V_CMFB_S3.n2 118.861
R3587 V_CMFB_S3.n5 V_CMFB_S3.n4 118.861
R3588 V_CMFB_S3.n9 V_CMFB_S3.n8 118.861
R3589 V_CMFB_S3.n12 V_CMFB_S3.n11 118.861
R3590 V_CMFB_S3.n15 V_CMFB_S3.n14 118.861
R3591 V_CMFB_S3.n2 V_CMFB_S3.t5 19.7005
R3592 V_CMFB_S3.n2 V_CMFB_S3.t10 19.7005
R3593 V_CMFB_S3.n4 V_CMFB_S3.t4 19.7005
R3594 V_CMFB_S3.n4 V_CMFB_S3.t7 19.7005
R3595 V_CMFB_S3.n8 V_CMFB_S3.t3 19.7005
R3596 V_CMFB_S3.n8 V_CMFB_S3.t9 19.7005
R3597 V_CMFB_S3.n11 V_CMFB_S3.t2 19.7005
R3598 V_CMFB_S3.n11 V_CMFB_S3.t8 19.7005
R3599 V_CMFB_S3.n14 V_CMFB_S3.t1 19.7005
R3600 V_CMFB_S3.n14 V_CMFB_S3.t6 19.7005
R3601 V_CMFB_S3.n6 V_CMFB_S3.n3 5.60467
R3602 V_CMFB_S3.n15 V_CMFB_S3.n13 5.54217
R3603 V_CMFB_S3.n3 V_CMFB_S3.n1 5.54217
R3604 V_CMFB_S3.n6 V_CMFB_S3.n5 5.04217
R3605 V_CMFB_S3.n9 V_CMFB_S3.n7 5.04217
R3606 V_CMFB_S3.n12 V_CMFB_S3.n0 5.04217
R3607 V_CMFB_S3.n16 V_CMFB_S3.n15 5.04217
R3608 V_CMFB_S3.n5 V_CMFB_S3.n1 4.97967
R3609 V_CMFB_S3.n10 V_CMFB_S3.n9 4.97967
R3610 V_CMFB_S3.n13 V_CMFB_S3.n12 4.97967
R3611 V_CMFB_S3 V_CMFB_S3.n16 1.40675
R3612 V_CMFB_S3.n13 V_CMFB_S3.n10 0.563
R3613 V_CMFB_S3.n10 V_CMFB_S3.n1 0.563
R3614 V_CMFB_S3.n7 V_CMFB_S3.n6 0.563
R3615 V_CMFB_S3.n7 V_CMFB_S3.n0 0.563
R3616 V_CMFB_S3.n16 V_CMFB_S3.n0 0.563
R3617 Vb1.n16 Vb1.t4 449.868
R3618 Vb1.n15 Vb1.t6 449.868
R3619 Vb1.n6 Vb1.t14 449.868
R3620 Vb1.n22 Vb1.n1 440.565
R3621 Vb1 Vb1.n14 433.519
R3622 Vb1 Vb1.n31 433.519
R3623 Vb1.n16 Vb1.t2 273.134
R3624 Vb1.n15 Vb1.t0 273.134
R3625 Vb1.n22 Vb1.t27 273.134
R3626 Vb1.n31 Vb1.t11 273.134
R3627 Vb1.n14 Vb1.t10 273.134
R3628 Vb1.n13 Vb1.t21 273.134
R3629 Vb1.n12 Vb1.t30 273.134
R3630 Vb1.n11 Vb1.t20 273.134
R3631 Vb1.n10 Vb1.t28 273.134
R3632 Vb1.n9 Vb1.t17 273.134
R3633 Vb1.n8 Vb1.t25 273.134
R3634 Vb1.n7 Vb1.t18 273.134
R3635 Vb1.n6 Vb1.t26 273.134
R3636 Vb1.n23 Vb1.t16 273.134
R3637 Vb1.n24 Vb1.t24 273.134
R3638 Vb1.n25 Vb1.t13 273.134
R3639 Vb1.n26 Vb1.t23 273.134
R3640 Vb1.n27 Vb1.t29 273.134
R3641 Vb1.n28 Vb1.t19 273.134
R3642 Vb1.n29 Vb1.t12 273.134
R3643 Vb1.n30 Vb1.t22 273.134
R3644 Vb1.n7 Vb1.n6 176.733
R3645 Vb1.n8 Vb1.n7 176.733
R3646 Vb1.n9 Vb1.n8 176.733
R3647 Vb1.n10 Vb1.n9 176.733
R3648 Vb1.n11 Vb1.n10 176.733
R3649 Vb1.n12 Vb1.n11 176.733
R3650 Vb1.n13 Vb1.n12 176.733
R3651 Vb1.n14 Vb1.n13 176.733
R3652 Vb1.n31 Vb1.n30 176.733
R3653 Vb1.n30 Vb1.n29 176.733
R3654 Vb1.n29 Vb1.n28 176.733
R3655 Vb1.n28 Vb1.n27 176.733
R3656 Vb1.n27 Vb1.n26 176.733
R3657 Vb1.n26 Vb1.n25 176.733
R3658 Vb1.n25 Vb1.n24 176.733
R3659 Vb1.n24 Vb1.n23 176.733
R3660 Vb1.n23 Vb1.n22 176.733
R3661 Vb1.n3 Vb1.t15 166.847
R3662 Vb1.t15 Vb1.n5 166.847
R3663 Vb1.n0 Vb1.n17 161.3
R3664 Vb1.n0 Vb1.n20 49.3505
R3665 Vb1.n19 Vb1.n18 49.3505
R3666 Vb1.n17 Vb1.n16 45.5227
R3667 Vb1.n17 Vb1.n15 45.5227
R3668 Vb1.n20 Vb1.t1 16.0005
R3669 Vb1.n20 Vb1.t3 16.0005
R3670 Vb1.n21 Vb1.t5 16.0005
R3671 Vb1.n21 Vb1.t8 16.0005
R3672 Vb1.n18 Vb1.t9 16.0005
R3673 Vb1.n18 Vb1.t7 16.0005
R3674 Vb1.n1 Vb1.n0 4.938
R3675 Vb1.n1 Vb1.n2 0.376365
R3676 Vb1.n21 Vb1.n2 51.6321
R3677 Vb1.n3 Vb1.n19 4.938
R3678 Vb1.n19 Vb1.n5 4.938
R3679 Vb1.n0 Vb1.n4 4.938
R3680 Vb1.n2 Vb1.n4 0.376365
R3681 Vb1.n1 Vb1.n5 0.688
R3682 Vb1.n4 Vb1.n3 0.688
R3683 V_CMFB_S1.n19 V_CMFB_S1.t0 121.785
R3684 V_CMFB_S1.n3 V_CMFB_S1.n2 118.861
R3685 V_CMFB_S1.n5 V_CMFB_S1.n4 118.861
R3686 V_CMFB_S1.n9 V_CMFB_S1.n8 118.861
R3687 V_CMFB_S1.n12 V_CMFB_S1.n11 118.861
R3688 V_CMFB_S1.n15 V_CMFB_S1.n14 118.861
R3689 V_CMFB_S1.n2 V_CMFB_S1.t9 19.7005
R3690 V_CMFB_S1.n2 V_CMFB_S1.t3 19.7005
R3691 V_CMFB_S1.n4 V_CMFB_S1.t10 19.7005
R3692 V_CMFB_S1.n4 V_CMFB_S1.t5 19.7005
R3693 V_CMFB_S1.n8 V_CMFB_S1.t2 19.7005
R3694 V_CMFB_S1.n8 V_CMFB_S1.t6 19.7005
R3695 V_CMFB_S1.n11 V_CMFB_S1.t4 19.7005
R3696 V_CMFB_S1.n11 V_CMFB_S1.t8 19.7005
R3697 V_CMFB_S1.n14 V_CMFB_S1.t1 19.7005
R3698 V_CMFB_S1.n14 V_CMFB_S1.t7 19.7005
R3699 V_CMFB_S1.n19 V_CMFB_S1.n18 5.90675
R3700 V_CMFB_S1.n6 V_CMFB_S1.n3 5.60467
R3701 V_CMFB_S1.n15 V_CMFB_S1.n13 5.54217
R3702 V_CMFB_S1.n3 V_CMFB_S1.n1 5.54217
R3703 V_CMFB_S1.n6 V_CMFB_S1.n5 5.04217
R3704 V_CMFB_S1.n9 V_CMFB_S1.n7 5.04217
R3705 V_CMFB_S1.n12 V_CMFB_S1.n0 5.04217
R3706 V_CMFB_S1.n5 V_CMFB_S1.n1 4.97967
R3707 V_CMFB_S1.n10 V_CMFB_S1.n9 4.97967
R3708 V_CMFB_S1.n13 V_CMFB_S1.n12 4.97967
R3709 V_CMFB_S1.n18 V_CMFB_S1.n17 4.5005
R3710 V_CMFB_S1.n17 V_CMFB_S1.n16 0.766125
R3711 V_CMFB_S1.n13 V_CMFB_S1.n10 0.563
R3712 V_CMFB_S1.n10 V_CMFB_S1.n1 0.563
R3713 V_CMFB_S1.n7 V_CMFB_S1.n6 0.563
R3714 V_CMFB_S1.n7 V_CMFB_S1.n0 0.563
R3715 V_CMFB_S1.n18 V_CMFB_S1.n0 0.563
R3716 V_CMFB_S1.n17 V_CMFB_S1.n15 0.479667
R3717 V_CMFB_S1 V_CMFB_S1.n19 0.063
R3718 V_p_mir.n0 V_p_mir.t2 16.0005
R3719 V_p_mir.n0 V_p_mir.t3 16.0005
R3720 V_p_mir.n1 V_p_mir.t0 9.6005
R3721 V_p_mir.t1 V_p_mir.n1 9.6005
R3722 V_p_mir.n1 V_p_mir.n0 89.8428
R3723 V_CMFB_S4 V_CMFB_S4.t0 124.285
R3724 V_CMFB_S4.n3 V_CMFB_S4.n2 24.288
R3725 V_CMFB_S4.n5 V_CMFB_S4.n4 24.288
R3726 V_CMFB_S4.n9 V_CMFB_S4.n8 24.288
R3727 V_CMFB_S4.n12 V_CMFB_S4.n11 24.288
R3728 V_CMFB_S4.n15 V_CMFB_S4.n14 24.288
R3729 V_CMFB_S4.n2 V_CMFB_S4.t6 8.0005
R3730 V_CMFB_S4.n2 V_CMFB_S4.t1 8.0005
R3731 V_CMFB_S4.n4 V_CMFB_S4.t5 8.0005
R3732 V_CMFB_S4.n4 V_CMFB_S4.t8 8.0005
R3733 V_CMFB_S4.n8 V_CMFB_S4.t4 8.0005
R3734 V_CMFB_S4.n8 V_CMFB_S4.t10 8.0005
R3735 V_CMFB_S4.n11 V_CMFB_S4.t3 8.0005
R3736 V_CMFB_S4.n11 V_CMFB_S4.t9 8.0005
R3737 V_CMFB_S4.n14 V_CMFB_S4.t2 8.0005
R3738 V_CMFB_S4.n14 V_CMFB_S4.t7 8.0005
R3739 V_CMFB_S4.n15 V_CMFB_S4.n13 5.7505
R3740 V_CMFB_S4.n3 V_CMFB_S4.n1 5.7505
R3741 V_CMFB_S4.n6 V_CMFB_S4.n3 5.7505
R3742 V_CMFB_S4.n6 V_CMFB_S4.n5 5.188
R3743 V_CMFB_S4.n5 V_CMFB_S4.n1 5.188
R3744 V_CMFB_S4.n9 V_CMFB_S4.n7 5.188
R3745 V_CMFB_S4.n10 V_CMFB_S4.n9 5.188
R3746 V_CMFB_S4.n12 V_CMFB_S4.n0 5.188
R3747 V_CMFB_S4.n13 V_CMFB_S4.n12 5.188
R3748 V_CMFB_S4.n16 V_CMFB_S4.n15 5.188
R3749 V_CMFB_S4 V_CMFB_S4.n16 1.1255
R3750 V_CMFB_S4.n13 V_CMFB_S4.n10 0.563
R3751 V_CMFB_S4.n10 V_CMFB_S4.n1 0.563
R3752 V_CMFB_S4.n7 V_CMFB_S4.n6 0.563
R3753 V_CMFB_S4.n7 V_CMFB_S4.n0 0.563
R3754 V_CMFB_S4.n16 V_CMFB_S4.n0 0.563
R3755 V_err_p.n1 V_err_p.n0 365.07
R3756 V_err_p.n0 V_err_p.t2 15.7605
R3757 V_err_p.n0 V_err_p.t0 15.7605
R3758 V_err_p.t1 V_err_p.n1 15.7605
R3759 V_err_p.n1 V_err_p.t3 15.7605
R3760 err_amp_out.n1 err_amp_out.t4 1025.2
R3761 err_amp_out.n1 err_amp_out.n0 179.382
R3762 err_amp_out.n2 err_amp_out.n1 39.3422
R3763 err_amp_out.n0 err_amp_out.t3 15.7605
R3764 err_amp_out.n0 err_amp_out.t0 15.7605
R3765 err_amp_out.n2 err_amp_out.t2 9.6005
R3766 err_amp_out.t1 err_amp_out.n2 9.6005
R3767 a_118660_3088.t0 a_118660_3088.t1 294.339
R3768 V_tot.n2 V_tot.t4 648.343
R3769 V_tot.n1 V_tot.t5 648.343
R3770 V_tot.n0 V_tot.t3 117.591
R3771 V_tot.t0 V_tot.n3 117.591
R3772 V_tot.n3 V_tot.t1 108.424
R3773 V_tot.n0 V_tot.t2 108.424
R3774 V_tot.n1 V_tot.n0 43.0496
R3775 V_tot.n3 V_tot.n2 43.0496
R3776 V_tot.n2 V_tot.n1 1.563
R3777 Vb1_2.n1 Vb1_2.t4 65.3505
R3778 Vb1_2.n3 Vb1_2.n2 49.3505
R3779 Vb1_2.n6 Vb1_2.n5 49.3505
R3780 Vb1_2.n2 Vb1_2.t0 16.0005
R3781 Vb1_2.n2 Vb1_2.t2 16.0005
R3782 Vb1_2.n6 Vb1_2.t1 16.0005
R3783 Vb1_2.t3 Vb1_2.n6 16.0005
R3784 Vb1_2.n1 Vb1_2.n0 6.41717
R3785 Vb1_2.n4 Vb1_2.n1 5.85467
R3786 Vb1_2.n3 Vb1_2.n0 5.72967
R3787 Vb1_2.n4 Vb1_2.n3 5.51092
R3788 Vb1_2.n5 Vb1_2.n0 5.16717
R3789 Vb1_2.n5 Vb1_2.n4 5.16717
R3790 Vb2_Vb3.n0 Vb2_Vb3.t3 661.375
R3791 Vb2_Vb3.n5 Vb2_Vb3.t0 661.375
R3792 Vb2_Vb3.t1 Vb2_Vb3.n6 213.131
R3793 Vb2_Vb3.n7 Vb2_Vb3.t4 213.131
R3794 Vb2_Vb3.t8 Vb2_Vb3.t1 146.155
R3795 Vb2_Vb3.t4 Vb2_Vb3.t8 146.155
R3796 Vb2_Vb3.n6 Vb2_Vb3.t2 76.2576
R3797 Vb2_Vb3.t6 Vb2_Vb3.n7 76.2576
R3798 Vb2_Vb3.n3 Vb2_Vb3.n1 72.5885
R3799 Vb2_Vb3.n3 Vb2_Vb3.n2 66.4444
R3800 Vb2_Vb3.n2 Vb2_Vb3.t9 11.2576
R3801 Vb2_Vb3.n2 Vb2_Vb3.t5 11.2576
R3802 Vb2_Vb3.n1 Vb2_Vb3.t7 11.2576
R3803 Vb2_Vb3.n1 Vb2_Vb3.t10 11.2576
R3804 Vb2_Vb3.n5 Vb2_Vb3.n4 5.1255
R3805 Vb2_Vb3.n4 Vb2_Vb3.n3 4.91892
R3806 Vb2_Vb3.n4 Vb2_Vb3.n0 4.7505
R3807 Vb2_Vb3.n6 Vb2_Vb3.n5 1.888
R3808 Vb2_Vb3.n7 Vb2_Vb3.n0 1.888
R3809 a_108650_n784.t0 a_108650_n784.t1 169.905
R3810 a_108510_3088.t0 a_108510_3088.t1 294.339
R3811 Vb2_2.n2 Vb2_2.t4 661.375
R3812 Vb2_2.n4 Vb2_2.t7 661.375
R3813 Vb2_2.t5 Vb2_2.n0 213.131
R3814 Vb2_2.n3 Vb2_2.t8 213.131
R3815 Vb2_2.n6 Vb2_2.n1 155.123
R3816 Vb2_2.t0 Vb2_2.t5 146.155
R3817 Vb2_2.t8 Vb2_2.t0 146.155
R3818 Vb2_2.t6 Vb2_2.n0 76.2576
R3819 Vb2_2.n3 Vb2_2.t9 76.2576
R3820 Vb2_2.n7 Vb2_2.n6 66.4336
R3821 Vb2_2.n1 Vb2_2.t3 21.8894
R3822 Vb2_2.n1 Vb2_2.t2 21.8894
R3823 Vb2_2.t6 Vb2_2.n7 11.2576
R3824 Vb2_2.n7 Vb2_2.t1 11.2576
R3825 Vb2_2.n5 Vb2_2.n4 5.1255
R3826 Vb2_2.n6 Vb2_2.n5 4.92976
R3827 Vb2_2.n5 Vb2_2.n2 4.7505
R3828 Vb2_2.n4 Vb2_2.n3 1.888
R3829 Vb2_2.n2 Vb2_2.n0 1.888
R3830 a_108630_3088.t0 a_108630_3088.t1 169.905
R3831 a_118780_3088.t0 a_118780_3088.t1 169.905
R3832 a_118760_n784.t0 a_118760_n784.t1 169.905
C0 V_err_gate V_err_mir_p 0.429395f
C1 cap_res_X Vb1 0.05001f
C2 VIN+ V_source 0.526392f
C3 V_tail_gate VIN+ 0.056217f
C4 V_CMFB_S2 V_CMFB_S1 1.15612f
C5 Vb3 cap_res_X 0.033116f
C6 cap_res_X cap_res_Y 0.345243f
C7 V_CMFB_S2 X 0.660498f
C8 VOUT+ Vb1 0.072817f
C9 VIN- V_source 0.526856f
C10 V_tail_gate VIN- 0.053799f
C11 VOUT+ Y 3.9238f
C12 cap_res_X X 0.05802f
C13 VOUT+ cap_res_Y 50.931602f
C14 V_tail_gate V_source 1.80219f
C15 VOUT- cap_res_Y 0.011897f
C16 VOUT+ V_CMFB_S4 0.015752f
C17 VOUT- V_CMFB_S1 0.139418f
C18 V_CMFB_S3 Y 0.674709f
C19 VOUT- X 3.9238f
C20 V_err_gate Y 0.013749f
C21 V_err_mir_p Y 0.013108f
C22 Vb1 VD2 0.357086f
C23 Y VD2 6.06356f
C24 V_err_amp_ref V_err_gate 0.665266f
C25 V_err_amp_ref V_err_mir_p 0.047104f
C26 VOUT+ cap_res_X 0.011897f
C27 V_CMFB_S3 V_CMFB_S4 1.15311f
C28 VIN+ VD2 0.533286f
C29 VOUT- V_CMFB_S2 0.015752f
C30 Vb2 Y 1.42469f
C31 Vb3 Vb2 2.03131f
C32 Vb1 VD1 0.329453f
C33 VOUT- cap_res_X 50.9331f
C34 Vb2 X 1.40695f
C35 VOUT+ VOUT- 0.118487f
C36 V_source VD2 5.03831f
C37 V_tail_gate VD2 0.01273f
C38 Vb1 Y 0.479502f
C39 VD1 X 6.06356f
C40 Vb1 cap_res_Y 0.072182f
C41 Vb3 Y 1.92012f
C42 VOUT+ V_CMFB_S3 0.139415f
C43 Vb1 VIN+ 0.020671f
C44 VD1 VIN- 0.533286f
C45 cap_res_Y Y 0.05802f
C46 Vb3 cap_res_Y 0.028593f
C47 Vb1 X 0.40038f
C48 Y X 0.081053f
C49 Vb3 X 1.94309f
C50 Vb1 VIN- 0.015071f
C51 VD1 V_source 5.03986f
C52 V_tail_gate VD1 0.012216f
C53 V_CMFB_S1 X 0.674709f
C54 V_CMFB_S4 Y 0.660498f
C55 Vb1 V_source 0.163912f
C56 Vb1 V_tail_gate 0.016424f
C57 VIN+ VIN- 0.075694f
C58 V_CMFB_S2 0 1.011331f
C59 V_tail_gate 0 4.57934f
C60 V_CMFB_S4 0 1.570256f
C61 V_CMFB_S1 0 5.22673f
C62 V_CMFB_S3 0 5.22768f
C63 VOUT- 0 26.588573f
C64 VOUT+ 0 26.559055f
C65 V_err_gate 0 0.519198f
C66 V_err_amp_ref 0 0.513289f
C67 Vb3 0 4.238993f
C68 Vb2 0 3.189286f
C69 V_source 0 18.610468f
C70 VIN- 0 1.83054f
C71 VIN+ 0 1.82624f
C72 VD1 0 3.177854f
C73 VD2 0 3.163864f
C74 Vb1 0 9.850801f
C75 cap_res_X 0 41.763683f
C76 V_err_mir_p 0 0.109531f
C77 cap_res_Y 0 41.743282f
C78 X 0 12.286777f
C79 Y 0 11.989277f
C80 Vb1_2.t1 0 0.046205f
C81 Vb1_2.n0 0 0.312531f
C82 Vb1_2.t4 0 0.157018f
C83 Vb1_2.n1 0 0.539239f
C84 Vb1_2.t0 0 0.046205f
C85 Vb1_2.t2 0 0.046205f
C86 Vb1_2.n2 0 0.100536f
C87 Vb1_2.n3 0 0.474689f
C88 Vb1_2.n4 0 0.470919f
C89 Vb1_2.n5 0 0.459714f
C90 Vb1_2.n6 0 0.100536f
C91 Vb1_2.t3 0 0.046205f
C92 V_tot.t1 0 0.07817f
C93 V_tot.t3 0 0.08327f
C94 V_tot.t2 0 0.07817f
C95 V_tot.n0 0 0.472359f
C96 V_tot.t5 0 0.023685f
C97 V_tot.n1 0 0.442517f
C98 V_tot.t4 0 0.023685f
C99 V_tot.n2 0 0.442517f
C100 V_tot.n3 0 0.472359f
C101 V_tot.t0 0 0.08327f
C102 err_amp_out.t2 0 0.036496f
C103 err_amp_out.t4 0 0.08233f
C104 err_amp_out.t3 0 0.036496f
C105 err_amp_out.t0 0 0.036496f
C106 err_amp_out.n0 0 0.114419f
C107 err_amp_out.n1 0 1.7352f
C108 err_amp_out.n2 0 0.122064f
C109 err_amp_out.t1 0 0.036496f
C110 V_CMFB_S4.n0 0 0.08992f
C111 V_CMFB_S4.n1 0 0.154718f
C112 V_CMFB_S4.t6 0 0.077555f
C113 V_CMFB_S4.t1 0 0.077555f
C114 V_CMFB_S4.n2 0 0.165875f
C115 V_CMFB_S4.n3 0 0.518857f
C116 V_CMFB_S4.t5 0 0.077555f
C117 V_CMFB_S4.t8 0 0.077555f
C118 V_CMFB_S4.n4 0 0.165875f
C119 V_CMFB_S4.n5 0 0.504805f
C120 V_CMFB_S4.n6 0 0.154718f
C121 V_CMFB_S4.n7 0 0.08992f
C122 V_CMFB_S4.t4 0 0.077555f
C123 V_CMFB_S4.t10 0 0.077555f
C124 V_CMFB_S4.n8 0 0.165875f
C125 V_CMFB_S4.n9 0 0.504805f
C126 V_CMFB_S4.n10 0 0.08992f
C127 V_CMFB_S4.t3 0 0.077555f
C128 V_CMFB_S4.t9 0 0.077555f
C129 V_CMFB_S4.n11 0 0.165875f
C130 V_CMFB_S4.n12 0 0.504805f
C131 V_CMFB_S4.n13 0 0.154718f
C132 V_CMFB_S4.t2 0 0.077555f
C133 V_CMFB_S4.t7 0 0.077555f
C134 V_CMFB_S4.n14 0 0.165875f
C135 V_CMFB_S4.n15 0 0.511831f
C136 V_CMFB_S4.n16 0 0.113187f
C137 V_CMFB_S4.t0 0 0.335044f
C138 Vb1.n0 0 0.061744f
C139 Vb1.n1 0 1.61865f
C140 Vb1.n2 0 0.051547f
C141 Vb1.n3 0 0.087649f
C142 Vb1.n4 0 0.042219f
C143 Vb1.n5 0 0.087649f
C144 Vb1.n14 0 0.011739f
C145 Vb1.t15 0 0.258007f
C146 Vb1.n18 0 0.014598f
C147 Vb1.n19 0 0.05393f
C148 Vb1.n20 0 0.014598f
C149 Vb1.n21 0 0.016981f
C150 Vb1.n22 0 0.018868f
C151 Vb1.n31 0 0.011739f
C152 Y.n0 0 0.083909f
C153 Y.n1 0 0.162703f
C154 Y.n2 0 0.102555f
C155 Y.n3 0 0.102555f
C156 Y.n4 0 0.102555f
C157 Y.n5 0 0.162703f
C158 Y.t7 0 0.023308f
C159 Y.t20 0 0.023308f
C160 Y.n6 0 0.050716f
C161 Y.n7 0 0.162065f
C162 Y.n8 0 0.078384f
C163 Y.n9 0 0.239296f
C164 Y.t19 0 0.023308f
C165 Y.t2 0 0.023308f
C166 Y.n10 0 0.050716f
C167 Y.n11 0 0.162065f
C168 Y.n12 0 0.177677f
C169 Y.n13 0 0.327848f
C170 Y.n14 0 0.102555f
C171 Y.n15 0 0.351511f
C172 Y.n16 0 0.102555f
C173 Y.n17 0 0.273038f
C174 Y.n18 0 0.162703f
C175 Y.t5 0 0.023308f
C176 Y.t23 0 0.023308f
C177 Y.n19 0 0.050716f
C178 Y.n20 0 0.157946f
C179 Y.n21 0 0.089133f
C180 Y.t8 0 0.023308f
C181 Y.t3 0 0.023308f
C182 Y.n22 0 0.050716f
C183 Y.n23 0 0.157946f
C184 Y.n24 0 0.089133f
C185 Y.t4 0 0.023308f
C186 Y.t24 0 0.023308f
C187 Y.n25 0 0.050716f
C188 Y.n26 0 0.157946f
C189 Y.n27 0 0.052064f
C190 Y.n28 0 0.052064f
C191 Y.t0 0 0.023308f
C192 Y.t1 0 0.023308f
C193 Y.n29 0 0.050716f
C194 Y.n30 0 0.157946f
C195 Y.n31 0 0.162703f
C196 Y.n32 0 0.046616f
C197 Y.n33 0 0.046616f
C198 Y.n34 0 0.078384f
C199 Y.n35 0 0.166674f
C200 Y.n36 0 0.074586f
C201 Y.t41 0 0.050112f
C202 Y.t30 0 0.050112f
C203 Y.t44 0 0.050112f
C204 Y.t27 0 0.050112f
C205 Y.t47 0 0.050112f
C206 Y.t29 0 0.050112f
C207 Y.t50 0 0.050112f
C208 Y.t33 0 0.056969f
C209 Y.n39 0 0.051413f
C210 Y.n40 0 0.031466f
C211 Y.n41 0 0.031466f
C212 Y.n42 0 0.031466f
C213 Y.n43 0 0.031466f
C214 Y.n44 0 0.031466f
C215 Y.n45 0 0.026513f
C216 Y.t54 0 0.050112f
C217 Y.t37 0 0.056969f
C218 Y.n46 0 0.04646f
C219 Y.n47 0 0.012874f
C220 Y.t43 0 0.032631f
C221 Y.t34 0 0.032631f
C222 Y.t46 0 0.032631f
C223 Y.t28 0 0.032631f
C224 Y.t49 0 0.032631f
C225 Y.t32 0 0.032631f
C226 Y.t52 0 0.032631f
C227 Y.t36 0 0.039624f
C228 Y.n48 0 0.039624f
C229 Y.n49 0 0.025639f
C230 Y.n50 0 0.025639f
C231 Y.n51 0 0.025639f
C232 Y.n52 0 0.025639f
C233 Y.n53 0 0.025639f
C234 Y.n54 0 0.020686f
C235 Y.t25 0 0.032631f
C236 Y.t40 0 0.039624f
C237 Y.n55 0 0.034671f
C238 Y.n56 0 0.012874f
C239 Y.n57 0 0.080313f
C240 Y.n58 0 0.074586f
C241 Y.n59 0 0.073885f
C242 Y.n60 0 0.074586f
C243 Y.t6 0 0.644946f
C244 Y.n61 0 0.074586f
C245 Y.n62 0 0.074586f
C246 Y.n64 0 0.692003f
C247 Y.n66 0 0.647964f
C248 Y.n67 0 0.024697f
C249 Y.n68 0 0.024862f
C250 Y.n69 0 0.024862f
C251 Y.t31 0 0.102555f
C252 Y.t51 0 0.102555f
C253 Y.t35 0 0.102555f
C254 Y.t53 0 0.102555f
C255 Y.t39 0 0.109229f
C256 Y.n70 0 0.086559f
C257 Y.n71 0 0.048947f
C258 Y.n72 0 0.048947f
C259 Y.n73 0 0.043994f
C260 Y.t48 0 0.102555f
C261 Y.t38 0 0.102555f
C262 Y.t45 0 0.102555f
C263 Y.t26 0 0.102555f
C264 Y.t42 0 0.109229f
C265 Y.n74 0 0.086559f
C266 Y.n75 0 0.048947f
C267 Y.n76 0 0.048947f
C268 Y.n77 0 0.043994f
C269 Y.n78 0 0.010564f
C270 Y.n79 0 0.025027f
C271 Y.n80 0 0.058911f
C272 Y.n81 0 0.0336f
C273 Y.n82 0 0.038132f
C274 Y.n83 0 1.03022f
C275 Y.n84 0 0.073885f
C276 Y.n85 0 0.074586f
C277 Y.n86 0 0.100673f
C278 Y.n87 0 0.121202f
C279 Y.n88 0 0.074586f
C280 Y.n89 0 0.096125f
C281 Y.n90 0 0.074586f
C282 Y.n91 0 0.074586f
C283 Y.n92 0 0.096125f
C284 Y.n93 0 0.074586f
C285 Y.n94 0 0.122901f
C286 Y.t15 0 0.054385f
C287 Y.t17 0 0.054385f
C288 Y.n95 0 0.111251f
C289 Y.n96 0 0.297688f
C290 Y.t22 0 0.054385f
C291 Y.t13 0 0.054385f
C292 Y.n97 0 0.111251f
C293 Y.n98 0 0.302606f
C294 Y.n99 0 0.100632f
C295 Y.t10 0 0.054385f
C296 Y.t12 0 0.054385f
C297 Y.n100 0 0.111251f
C298 Y.n101 0 0.297688f
C299 Y.n102 0 0.058991f
C300 Y.t11 0 0.054385f
C301 Y.t14 0 0.054385f
C302 Y.n103 0 0.111251f
C303 Y.n104 0 0.297688f
C304 Y.n105 0 0.058991f
C305 Y.t9 0 0.054385f
C306 Y.t21 0 0.054385f
C307 Y.n106 0 0.111251f
C308 Y.n107 0 0.302606f
C309 Y.n108 0 0.100632f
C310 Y.t16 0 0.054385f
C311 Y.t18 0 0.054385f
C312 Y.n109 0 0.111251f
C313 Y.n110 0 0.297688f
C314 Y.n111 0 0.096125f
C315 Y.n112 0 0.082469f
C316 Y.n113 0 0.049724f
C317 Y.n114 0 0.049724f
C318 Y.n115 0 0.082469f
C319 Y.n116 0 0.096125f
C320 Y.n117 0 0.170057f
C321 Y.n118 0 0.251893f
C322 Y.n119 0 0.320326f
C323 Y.n120 0 0.074586f
C324 Y.n121 0 0.074586f
C325 Y.n122 0 0.121202f
C326 Y.n123 0 0.074586f
C327 Y.n124 0 0.074586f
C328 Y.n125 0 0.074586f
C329 Y.n126 0 0.074586f
C330 Y.n127 0 0.121202f
C331 Y.n128 0 0.074586f
C332 Y.n129 0 0.074586f
C333 Y.n130 0 0.074586f
C334 Y.n131 0 0.074586f
C335 Y.n132 0 0.074586f
C336 Y.n133 0 0.074586f
C337 Y.n134 0 0.074586f
C338 Y.n135 0 0.121202f
C339 Y.n136 0 0.582701f
C340 Y.n137 0 0.582701f
C341 Y.n138 0 0.074586f
C342 Y.n140 0 0.074586f
C343 Y.n141 0 0.074586f
C344 Y.n143 0 0.913675f
C345 Y.n144 0 0.913675f
C346 Y.n146 0 0.456838f
C347 Y.n147 0 2.20415f
C348 Y.n148 0 0.601348f
C349 Y.n149 0 0.615332f
C350 Y.n150 0 0.225311f
C351 Y.n151 0 0.102555f
C352 Y.n152 0 0.239296f
C353 Y.n153 0 0.102555f
C354 Y.n154 0 0.102555f
C355 Y.n155 0 0.102555f
C356 Y.n156 0 0.206665f
C357 VD2.n0 0 0.259344f
C358 VD2.n1 0 0.073525f
C359 VD2.n2 0 0.119354f
C360 VD2.t10 0 0.048999f
C361 VD2.t15 0 0.048999f
C362 VD2.n3 0 0.106617f
C363 VD2.n4 0 0.410788f
C364 VD2.n5 0 0.104208f
C365 VD2.t16 0 0.048999f
C366 VD2.t8 0 0.048999f
C367 VD2.n6 0 0.106617f
C368 VD2.n7 0 0.422242f
C369 VD2.t3 0 0.048999f
C370 VD2.t6 0 0.048999f
C371 VD2.n8 0 0.106617f
C372 VD2.n9 0 0.340702f
C373 VD2.n10 0 0.097999f
C374 VD2.t2 0 0.048999f
C375 VD2.t5 0 0.048999f
C376 VD2.n11 0 0.106617f
C377 VD2.n12 0 0.340702f
C378 VD2.n13 0 0.119354f
C379 VD2.t9 0 0.048999f
C380 VD2.t14 0 0.048999f
C381 VD2.n14 0 0.106617f
C382 VD2.n15 0 0.422242f
C383 VD2.n16 0 0.177134f
C384 VD2.t19 0 0.048999f
C385 VD2.t13 0 0.048999f
C386 VD2.n17 0 0.106617f
C387 VD2.n18 0 0.410788f
C388 VD2.n19 0 0.073525f
C389 VD2.n20 0 0.185267f
C390 VD2.n21 0 0.442388f
C391 VD2.n22 0 0.164783f
C392 VD2.n23 0 0.434039f
C393 VD2.t20 0 0.048999f
C394 VD2.t0 0 0.048999f
C395 VD2.n24 0 0.106617f
C396 VD2.n25 0 0.332044f
C397 VD2.n26 0 0.187379f
C398 VD2.t1 0 0.048999f
C399 VD2.t4 0 0.048999f
C400 VD2.n27 0 0.106617f
C401 VD2.n28 0 0.332044f
C402 VD2.n29 0 0.109452f
C403 VD2.n30 0 0.187379f
C404 VD2.t21 0 0.048999f
C405 VD2.t7 0 0.048999f
C406 VD2.n31 0 0.106617f
C407 VD2.n32 0 0.332044f
C408 VD2.n33 0 0.434039f
C409 VD2.n34 0 0.164783f
C410 VD2.n35 0 0.442388f
C411 VD2.n36 0 0.185267f
C412 VD2.n37 0 0.073525f
C413 VD2.t17 0 0.048999f
C414 VD2.t11 0 0.048999f
C415 VD2.n38 0 0.106617f
C416 VD2.n39 0 0.410788f
C417 VD2.n40 0 0.177134f
C418 VD2.n41 0 0.104208f
C419 VD2.t18 0 0.048999f
C420 VD2.t12 0 0.048999f
C421 VD2.n42 0 0.106617f
C422 VD2.n43 0 0.410788f
C423 VD2.n44 0 0.073525f
C424 VD2.n45 0 0.056907f
C425 VD3.t29 0 0.055114f
C426 VD3.n0 0 0.075585f
C427 VD3.n1 0 0.075585f
C428 VD3.n2 0 0.075585f
C429 VD3.n3 0 0.075585f
C430 VD3.t21 0 0.055114f
C431 VD3.t23 0 0.055114f
C432 VD3.n4 0 0.116929f
C433 VD3.t25 0 0.055114f
C434 VD3.t27 0 0.055114f
C435 VD3.n5 0 0.116929f
C436 VD3.n6 0 0.418462f
C437 VD3.n7 0 0.075585f
C438 VD3.t31 0 0.055114f
C439 VD3.t17 0 0.055114f
C440 VD3.n8 0 0.116929f
C441 VD3.n9 0 0.075585f
C442 VD3.t0 0 0.09664f
C443 VD3.t2 0 0.196047f
C444 VD3.n10 0 0.075585f
C445 VD3.n11 0 0.075585f
C446 VD3.n12 0 0.075585f
C447 VD3.n13 0 0.059781f
C448 VD3.n14 0 0.075585f
C449 VD3.n15 0 0.075585f
C450 VD3.n16 0 0.075585f
C451 VD3.t8 0 0.055114f
C452 VD3.t10 0 0.055114f
C453 VD3.n17 0 0.112741f
C454 VD3.n18 0 0.310905f
C455 VD3.n19 0 0.17942f
C456 VD3.n20 0 0.059781f
C457 VD3.t13 0 0.055114f
C458 VD3.t7 0 0.055114f
C459 VD3.n21 0 0.112741f
C460 VD3.n22 0 0.310905f
C461 VD3.n23 0 0.101979f
C462 VD3.t37 0 0.055114f
C463 VD3.t11 0 0.055114f
C464 VD3.n24 0 0.112741f
C465 VD3.n25 0 0.328078f
C466 VD3.n26 0 0.272689f
C467 VD3.n27 0 0.324616f
C468 VD3.n28 0 0.075585f
C469 VD3.n29 0 0.075585f
C470 VD3.n30 0 0.129911f
C471 VD3.n31 0 0.151169f
C472 VD3.n32 0 0.151169f
C473 VD3.t9 0 0.055114f
C474 VD3.t12 0 0.055114f
C475 VD3.n33 0 0.112741f
C476 VD3.n34 0 0.310905f
C477 VD3.n35 0 0.129911f
C478 VD3.n36 0 0.075585f
C479 VD3.n37 0 0.075585f
C480 VD3.n38 0 0.075585f
C481 VD3.n39 0 0.075585f
C482 VD3.n40 0 0.075585f
C483 VD3.n41 0 0.129911f
C484 VD3.t14 0 0.055114f
C485 VD3.t15 0 0.055114f
C486 VD3.n42 0 0.112741f
C487 VD3.n43 0 0.310905f
C488 VD3.n44 0 0.101979f
C489 VD3.t6 0 0.055114f
C490 VD3.t36 0 0.055114f
C491 VD3.n45 0 0.112741f
C492 VD3.n46 0 0.315889f
C493 VD3.n47 0 0.129911f
C494 VD3.n48 0 0.751122f
C495 VD3.n49 0 0.075585f
C496 VD3.n50 0 0.075585f
C497 VD3.n51 0 0.751122f
C498 VD3.n52 0 0.129911f
C499 VD3.t3 0 0.09664f
C500 VD3.n53 0 0.220264f
C501 VD3.t5 0 0.196047f
C502 VD3.n54 0 0.568717f
C503 VD3.t4 0 0.469785f
C504 VD3.t28 0 0.368475f
C505 VD3.t34 0 0.368475f
C506 VD3.t20 0 0.368475f
C507 VD3.t22 0 0.368475f
C508 VD3.t24 0 0.368475f
C509 VD3.t26 0 0.368475f
C510 VD3.t30 0 0.368475f
C511 VD3.t16 0 0.368475f
C512 VD3.t32 0 0.368475f
C513 VD3.t18 0 0.368475f
C514 VD3.t1 0 0.469785f
C515 VD3.n55 0 0.568717f
C516 VD3.n56 0 0.232551f
C517 VD3.n57 0 0.272343f
C518 VD3.t33 0 0.055114f
C519 VD3.t19 0 0.055114f
C520 VD3.n58 0 0.116929f
C521 VD3.n59 0 0.468223f
C522 VD3.n60 0 0.075585f
C523 VD3.n61 0 0.324614f
C524 VD3.n62 0 0.075585f
C525 VD3.n63 0 0.075585f
C526 VD3.n64 0 0.418462f
C527 VD3.n65 0 0.075585f
C528 VD3.n66 0 0.075585f
C529 VD3.n67 0 0.075585f
C530 VD3.n68 0 0.075585f
C531 VD3.n69 0 0.075585f
C532 VD3.n70 0 0.075585f
C533 VD3.n71 0 0.075585f
C534 VD3.n72 0 0.418462f
C535 VD3.n73 0 0.075585f
C536 VD3.n74 0 0.075585f
C537 VD3.n75 0 0.075585f
C538 VD3.n76 0 0.075585f
C539 VD3.n77 0 0.418462f
C540 VD3.n78 0 0.116929f
C541 VD3.t35 0 0.055114f
C542 Vb2.t13 0 0.042112f
C543 Vb2.t1 0 0.022626f
C544 Vb2.t2 0 0.022626f
C545 Vb2.n0 0 0.048048f
C546 Vb2.t0 0 0.042236f
C547 Vb2.n1 0 0.19558f
C548 Vb2.t17 0 0.025365f
C549 Vb2.n2 0 0.097376f
C550 Vb2.n3 0 0.189208f
C551 Vb2.t11 0 0.032f
C552 Vb2.t7 0 0.032f
C553 Vb2.t24 0 0.032f
C554 Vb2.t5 0 0.032f
C555 Vb2.t23 0 0.036927f
C556 Vb2.n4 0 0.029981f
C557 Vb2.n5 0 0.018424f
C558 Vb2.n6 0 0.018424f
C559 Vb2.n7 0 0.016154f
C560 Vb2.t16 0 0.032f
C561 Vb2.t20 0 0.032f
C562 Vb2.t21 0 0.032f
C563 Vb2.t3 0 0.032f
C564 Vb2.t8 0 0.036927f
C565 Vb2.n8 0 0.029981f
C566 Vb2.n9 0 0.018424f
C567 Vb2.n10 0 0.018424f
C568 Vb2.n11 0 0.016154f
C569 Vb2.n12 0 0.011973f
C570 Vb2.t18 0 0.032f
C571 Vb2.t12 0 0.032f
C572 Vb2.t9 0 0.032f
C573 Vb2.t4 0 0.032f
C574 Vb2.t22 0 0.036927f
C575 Vb2.n13 0 0.029981f
C576 Vb2.n14 0 0.018424f
C577 Vb2.n15 0 0.018424f
C578 Vb2.n16 0 0.016154f
C579 Vb2.t15 0 0.032f
C580 Vb2.t19 0 0.032f
C581 Vb2.t6 0 0.032f
C582 Vb2.t10 0 0.032f
C583 Vb2.t14 0 0.036927f
C584 Vb2.n17 0 0.029981f
C585 Vb2.n18 0 0.018424f
C586 Vb2.n19 0 0.018424f
C587 Vb2.n20 0 0.016154f
C588 Vb2.n21 0 0.011797f
C589 Vb2.n22 0 0.203812f
C590 Vb2.n23 0 0.093025f
C591 VD1.n0 0 0.259344f
C592 VD1.n1 0 0.073525f
C593 VD1.n2 0 0.119354f
C594 VD1.t17 0 0.048999f
C595 VD1.t11 0 0.048999f
C596 VD1.n3 0 0.106617f
C597 VD1.n4 0 0.410788f
C598 VD1.n5 0 0.104207f
C599 VD1.t13 0 0.048999f
C600 VD1.t8 0 0.048999f
C601 VD1.n6 0 0.106617f
C602 VD1.n7 0 0.422242f
C603 VD1.t2 0 0.048999f
C604 VD1.t21 0 0.048999f
C605 VD1.n8 0 0.106617f
C606 VD1.n9 0 0.340702f
C607 VD1.n10 0 0.097999f
C608 VD1.t20 0 0.048999f
C609 VD1.t5 0 0.048999f
C610 VD1.n11 0 0.106617f
C611 VD1.n12 0 0.340702f
C612 VD1.n13 0 0.119354f
C613 VD1.t7 0 0.048999f
C614 VD1.t12 0 0.048999f
C615 VD1.n14 0 0.106617f
C616 VD1.n15 0 0.422242f
C617 VD1.n16 0 0.177134f
C618 VD1.t16 0 0.048999f
C619 VD1.t10 0 0.048999f
C620 VD1.n17 0 0.106617f
C621 VD1.n18 0 0.410788f
C622 VD1.n19 0 0.073525f
C623 VD1.n20 0 0.185267f
C624 VD1.n21 0 0.442387f
C625 VD1.n22 0 0.164783f
C626 VD1.n23 0 0.434039f
C627 VD1.t1 0 0.048999f
C628 VD1.t6 0 0.048999f
C629 VD1.n24 0 0.106617f
C630 VD1.n25 0 0.332043f
C631 VD1.n26 0 0.187379f
C632 VD1.t19 0 0.048999f
C633 VD1.t3 0 0.048999f
C634 VD1.n27 0 0.106617f
C635 VD1.n28 0 0.332043f
C636 VD1.n29 0 0.109452f
C637 VD1.n30 0 0.187379f
C638 VD1.t0 0 0.048999f
C639 VD1.t4 0 0.048999f
C640 VD1.n31 0 0.106617f
C641 VD1.n32 0 0.332043f
C642 VD1.n33 0 0.434039f
C643 VD1.n34 0 0.164783f
C644 VD1.n35 0 0.442387f
C645 VD1.n36 0 0.185267f
C646 VD1.n37 0 0.073525f
C647 VD1.t14 0 0.048999f
C648 VD1.t18 0 0.048999f
C649 VD1.n38 0 0.106617f
C650 VD1.n39 0 0.410788f
C651 VD1.n40 0 0.177134f
C652 VD1.n41 0 0.104207f
C653 VD1.t15 0 0.048999f
C654 VD1.t9 0 0.048999f
C655 VD1.n42 0 0.106617f
C656 VD1.n43 0 0.410788f
C657 VD1.n44 0 0.073525f
C658 VD1.n45 0 0.056907f
C659 V_source.n0 0 0.774331f
C660 V_source.n1 0 0.828472f
C661 V_source.n2 0 0.6888f
C662 V_source.n3 0 0.206488f
C663 V_source.t20 0 0.025305f
C664 V_source.t1 0 0.025305f
C665 V_source.n4 0 0.054098f
C666 V_source.n5 0 0.204115f
C667 V_source.n6 0 0.049378f
C668 V_source.t2 0 0.025305f
C669 V_source.t9 0 0.025305f
C670 V_source.n7 0 0.054098f
C671 V_source.n8 0 0.160508f
C672 V_source.n9 0 0.086782f
C673 V_source.t16 0 0.025305f
C674 V_source.t15 0 0.025305f
C675 V_source.n10 0 0.054098f
C676 V_source.n11 0 0.124175f
C677 V_source.t0 0 0.056141f
C678 V_source.n12 0 0.237776f
C679 V_source.n13 0 0.044537f
C680 V_source.t4 0 0.025305f
C681 V_source.t11 0 0.025305f
C682 V_source.n14 0 0.054098f
C683 V_source.n15 0 0.160508f
C684 V_source.n16 0 0.051601f
C685 V_source.n17 0 0.051601f
C686 V_source.n18 0 0.173762f
C687 V_source.n19 0 0.081951f
C688 V_source.n20 0 0.055202f
C689 V_source.t25 0 0.015183f
C690 V_source.t27 0 0.015183f
C691 V_source.n21 0 0.033036f
C692 V_source.n22 0 0.138652f
C693 V_source.t21 0 0.015183f
C694 V_source.t23 0 0.015183f
C695 V_source.n23 0 0.033036f
C696 V_source.n24 0 0.133856f
C697 V_source.n25 0 0.081951f
C698 V_source.n26 0 0.063658f
C699 V_source.t22 0 0.015183f
C700 V_source.t28 0 0.015183f
C701 V_source.n27 0 0.033036f
C702 V_source.n28 0 0.133856f
C703 V_source.n29 0 0.032451f
C704 V_source.n30 0 0.032451f
C705 V_source.t26 0 0.015183f
C706 V_source.t29 0 0.015183f
C707 V_source.n31 0 0.033036f
C708 V_source.n32 0 0.10026f
C709 V_source.t30 0 0.015183f
C710 V_source.t24 0 0.015183f
C711 V_source.n33 0 0.033036f
C712 V_source.n34 0 0.10026f
C713 V_source.n35 0 0.082048f
C714 V_source.t40 0 0.015183f
C715 V_source.t38 0 0.015183f
C716 V_source.n36 0 0.033036f
C717 V_source.n37 0 0.10026f
C718 V_source.n38 0 0.082048f
C719 V_source.t39 0 0.015183f
C720 V_source.t36 0 0.015183f
C721 V_source.n39 0 0.033036f
C722 V_source.n40 0 0.10026f
C723 V_source.n41 0 0.032451f
C724 V_source.t37 0 0.015183f
C725 V_source.t31 0 0.015183f
C726 V_source.n42 0 0.033036f
C727 V_source.n43 0 0.138652f
C728 V_source.t32 0 0.015183f
C729 V_source.t33 0 0.015183f
C730 V_source.n44 0 0.033036f
C731 V_source.n45 0 0.133856f
C732 V_source.n46 0 0.055202f
C733 V_source.n47 0 0.032451f
C734 V_source.t34 0 0.015183f
C735 V_source.t35 0 0.015183f
C736 V_source.n48 0 0.033036f
C737 V_source.n49 0 0.133856f
C738 V_source.n50 0 0.063658f
C739 V_source.n51 0 0.173762f
C740 V_source.t8 0 0.025305f
C741 V_source.t5 0 0.025305f
C742 V_source.n52 0 0.054098f
C743 V_source.n53 0 0.160508f
C744 V_source.t7 0 0.025305f
C745 V_source.t14 0 0.025305f
C746 V_source.n54 0 0.054098f
C747 V_source.n55 0 0.162758f
C748 V_source.n56 0 0.086782f
C749 V_source.t12 0 0.025305f
C750 V_source.t19 0 0.025305f
C751 V_source.n57 0 0.054098f
C752 V_source.n58 0 0.160508f
C753 V_source.n59 0 0.138969f
C754 V_source.t10 0 0.025305f
C755 V_source.t17 0 0.025305f
C756 V_source.n60 0 0.054098f
C757 V_source.n61 0 0.194636f
C758 V_source.n62 0 0.051601f
C759 V_source.t13 0 0.025305f
C760 V_source.t3 0 0.025305f
C761 V_source.n63 0 0.054098f
C762 V_source.n64 0 0.194636f
C763 V_source.n65 0 0.051601f
C764 V_source.n66 0 0.051601f
C765 V_source.t18 0 0.025305f
C766 V_source.t6 0 0.025305f
C767 V_source.n67 0 0.054098f
C768 V_source.n68 0 0.194636f
C769 V_source.n69 0 0.077849f
C770 V_source.n70 0 0.133118f
C771 VD4.n0 0 0.400201f
C772 VD4.n1 0 0.100435f
C773 VD4.n2 0 0.205496f
C774 VD4.n3 0 0.129911f
C775 VD4.n4 0 0.151169f
C776 VD4.n5 0 0.125802f
C777 VD4.n6 0 0.151169f
C778 VD4.n7 0 0.205496f
C779 VD4.n8 0 0.204968f
C780 VD4.t18 0 0.055114f
C781 VD4.n9 0 0.204788f
C782 VD4.n10 0 0.059781f
C783 VD4.t22 0 0.055114f
C784 VD4.t23 0 0.055114f
C785 VD4.n11 0 0.112741f
C786 VD4.n12 0 0.310905f
C787 VD4.t20 0 0.055114f
C788 VD4.t21 0 0.055114f
C789 VD4.n13 0 0.112741f
C790 VD4.n14 0 0.310905f
C791 VD4.n15 0 0.075585f
C792 VD4.t26 0 0.09664f
C793 VD4.n16 0 0.220264f
C794 VD4.t13 0 0.055114f
C795 VD4.t35 0 0.055114f
C796 VD4.n17 0 0.116929f
C797 VD4.n18 0 0.418462f
C798 VD4.n19 0 0.075585f
C799 VD4.t9 0 0.055114f
C800 VD4.t5 0 0.055114f
C801 VD4.n20 0 0.116929f
C802 VD4.n21 0 0.075585f
C803 VD4.n22 0 0.075585f
C804 VD4.t15 0 0.055114f
C805 VD4.t11 0 0.055114f
C806 VD4.n23 0 0.116929f
C807 VD4.n24 0 0.075585f
C808 VD4.n25 0 0.075585f
C809 VD4.t7 0 0.055114f
C810 VD4.t37 0 0.055114f
C811 VD4.n26 0 0.116929f
C812 VD4.t1 0 0.055114f
C813 VD4.t3 0 0.055114f
C814 VD4.n27 0 0.116929f
C815 VD4.n28 0 0.467972f
C816 VD4.t29 0 0.09664f
C817 VD4.t28 0 0.196047f
C818 VD4.n29 0 0.568717f
C819 VD4.t27 0 0.469785f
C820 VD4.t34 0 0.368475f
C821 VD4.t12 0 0.368475f
C822 VD4.t4 0 0.368475f
C823 VD4.t8 0 0.368475f
C824 VD4.t10 0 0.368475f
C825 VD4.t14 0 0.368475f
C826 VD4.t36 0 0.368475f
C827 VD4.t6 0 0.368475f
C828 VD4.t2 0 0.368475f
C829 VD4.t0 0 0.368475f
C830 VD4.t30 0 0.469785f
C831 VD4.t31 0 0.196047f
C832 VD4.n30 0 0.568717f
C833 VD4.n31 0 0.232453f
C834 VD4.n32 0 0.272689f
C835 VD4.n33 0 0.324616f
C836 VD4.n34 0 0.075585f
C837 VD4.n35 0 0.075585f
C838 VD4.n36 0 0.418462f
C839 VD4.n37 0 0.075585f
C840 VD4.n38 0 0.075585f
C841 VD4.n39 0 0.075585f
C842 VD4.n40 0 0.075585f
C843 VD4.n41 0 0.418462f
C844 VD4.n42 0 0.075585f
C845 VD4.n43 0 0.075585f
C846 VD4.n44 0 0.075585f
C847 VD4.n45 0 0.075585f
C848 VD4.n46 0 0.418462f
C849 VD4.n47 0 0.075585f
C850 VD4.n48 0 0.075585f
C851 VD4.n49 0 0.075585f
C852 VD4.n50 0 0.075585f
C853 VD4.n51 0 0.075585f
C854 VD4.n52 0 0.075585f
C855 VD4.n53 0 0.075585f
C856 VD4.n54 0 0.129911f
C857 VD4.n55 0 0.751122f
C858 VD4.n56 0 0.77649f
C859 VD4.n57 0 0.059781f
C860 VD4.t17 0 0.055114f
C861 VD4.t19 0 0.055114f
C862 VD4.n58 0 0.112741f
C863 VD4.n59 0 0.310905f
C864 VD4.n60 0 0.101979f
C865 VD4.t33 0 0.055114f
C866 VD4.t24 0 0.055114f
C867 VD4.n61 0 0.112741f
C868 VD4.n62 0 0.315889f
C869 VD4.n63 0 0.172955f
C870 VD4.n64 0 0.155278f
C871 VD4.n65 0 0.272689f
C872 VD4.t16 0 0.055114f
C873 VD4.t32 0 0.055114f
C874 VD4.n66 0 0.112741f
C875 VD4.n67 0 0.328078f
C876 VD4.n68 0 0.101979f
C877 VD4.n69 0 0.310905f
C878 VD4.n70 0 0.112741f
C879 VD4.t25 0 0.055114f
C880 Vb3.t14 0 0.091008f
C881 Vb3.t10 0 0.091008f
C882 Vb3.t6 0 0.091008f
C883 Vb3.t4 0 0.091008f
C884 Vb3.t22 0 0.105022f
C885 Vb3.n0 0 0.085266f
C886 Vb3.n1 0 0.052398f
C887 Vb3.n2 0 0.052398f
C888 Vb3.n3 0 0.045943f
C889 Vb3.t13 0 0.091008f
C890 Vb3.t16 0 0.091008f
C891 Vb3.t18 0 0.091008f
C892 Vb3.t8 0 0.091008f
C893 Vb3.t12 0 0.105022f
C894 Vb3.n4 0 0.085266f
C895 Vb3.n5 0 0.052398f
C896 Vb3.n6 0 0.052398f
C897 Vb3.n7 0 0.045943f
C898 Vb3.n8 0 0.049338f
C899 Vb3.t7 0 0.091008f
C900 Vb3.t5 0 0.091008f
C901 Vb3.t2 0 0.091008f
C902 Vb3.t19 0 0.091008f
C903 Vb3.t21 0 0.105022f
C904 Vb3.n9 0 0.085266f
C905 Vb3.n10 0 0.052398f
C906 Vb3.n11 0 0.052398f
C907 Vb3.n12 0 0.045943f
C908 Vb3.t11 0 0.091008f
C909 Vb3.t15 0 0.091008f
C910 Vb3.t17 0 0.091008f
C911 Vb3.t20 0 0.091008f
C912 Vb3.t3 0 0.105022f
C913 Vb3.n13 0 0.085266f
C914 Vb3.n14 0 0.052398f
C915 Vb3.n15 0 0.052398f
C916 Vb3.n16 0 0.045943f
C917 Vb3.n17 0 0.050888f
C918 Vb3.t0 0 0.064349f
C919 Vb3.t1 0 0.064349f
C920 Vb3.n18 0 0.18786f
C921 Vb3.t9 0 0.118885f
C922 Vb3.n19 0 1.02001f
C923 Vb3.n20 0 1.04758f
C924 cap_res_X.t125 0 0.398042f
C925 cap_res_X.t18 0 0.399485f
C926 cap_res_X.t88 0 0.398042f
C927 cap_res_X.t127 0 0.399485f
C928 cap_res_X.t37 0 0.398042f
C929 cap_res_X.t59 0 0.399485f
C930 cap_res_X.t52 0 0.398042f
C931 cap_res_X.t91 0 0.399485f
C932 cap_res_X.t71 0 0.398042f
C933 cap_res_X.t21 0 0.399485f
C934 cap_res_X.t97 0 0.398042f
C935 cap_res_X.t133 0 0.399485f
C936 cap_res_X.t111 0 0.398042f
C937 cap_res_X.t60 0 0.399485f
C938 cap_res_X.t136 0 0.398042f
C939 cap_res_X.t32 0 0.399485f
C940 cap_res_X.t11 0 0.398042f
C941 cap_res_X.t101 0 0.399485f
C942 cap_res_X.t102 0 0.398042f
C943 cap_res_X.t137 0 0.399485f
C944 cap_res_X.t117 0 0.398042f
C945 cap_res_X.t65 0 0.399485f
C946 cap_res_X.t1 0 0.398042f
C947 cap_res_X.t36 0 0.399485f
C948 cap_res_X.t16 0 0.398042f
C949 cap_res_X.t104 0 0.399485f
C950 cap_res_X.t39 0 0.398042f
C951 cap_res_X.t74 0 0.399485f
C952 cap_res_X.t54 0 0.398042f
C953 cap_res_X.t4 0 0.399485f
C954 cap_res_X.t5 0 0.398042f
C955 cap_res_X.t40 0 0.399485f
C956 cap_res_X.t22 0 0.398042f
C957 cap_res_X.t108 0 0.399485f
C958 cap_res_X.t47 0 0.398042f
C959 cap_res_X.t80 0 0.399485f
C960 cap_res_X.t62 0 0.398042f
C961 cap_res_X.t10 0 0.399485f
C962 cap_res_X.t86 0 0.398042f
C963 cap_res_X.t121 0 0.399485f
C964 cap_res_X.t103 0 0.398042f
C965 cap_res_X.t49 0 0.399485f
C966 cap_res_X.t50 0 0.398042f
C967 cap_res_X.t87 0 0.399485f
C968 cap_res_X.t66 0 0.398042f
C969 cap_res_X.t14 0 0.399485f
C970 cap_res_X.t90 0 0.398042f
C971 cap_res_X.t128 0 0.399485f
C972 cap_res_X.t105 0 0.398042f
C973 cap_res_X.t53 0 0.399485f
C974 cap_res_X.t132 0 0.398042f
C975 cap_res_X.t26 0 0.399485f
C976 cap_res_X.t7 0 0.398042f
C977 cap_res_X.t98 0 0.399485f
C978 cap_res_X.t82 0 0.398042f
C979 cap_res_X.t31 0 0.399485f
C980 cap_res_X.t109 0 0.398042f
C981 cap_res_X.t68 0 0.399485f
C982 cap_res_X.t48 0 0.398042f
C983 cap_res_X.t138 0 0.399485f
C984 cap_res_X.t77 0 0.398042f
C985 cap_res_X.t34 0 0.399485f
C986 cap_res_X.t25 0 0.398042f
C987 cap_res_X.t57 0 0.399485f
C988 cap_res_X.t41 0 0.398042f
C989 cap_res_X.t131 0 0.399485f
C990 cap_res_X.t8 0 0.398042f
C991 cap_res_X.t46 0 0.399485f
C992 cap_res_X.t100 0 0.398042f
C993 cap_res_X.t124 0 0.399485f
C994 cap_res_X.t42 0 0.398042f
C995 cap_res_X.t79 0 0.399485f
C996 cap_res_X.t119 0 0.398042f
C997 cap_res_X.t17 0 0.417559f
C998 cap_res_X.t81 0 0.398042f
C999 cap_res_X.t123 0 0.213796f
C1000 cap_res_X.n0 0 0.228815f
C1001 cap_res_X.t44 0 0.398042f
C1002 cap_res_X.t83 0 0.213796f
C1003 cap_res_X.n1 0 0.22697f
C1004 cap_res_X.t3 0 0.398042f
C1005 cap_res_X.t45 0 0.213796f
C1006 cap_res_X.n2 0 0.22697f
C1007 cap_res_X.t29 0 0.398042f
C1008 cap_res_X.t67 0 0.213796f
C1009 cap_res_X.n3 0 0.22697f
C1010 cap_res_X.t130 0 0.398042f
C1011 cap_res_X.t30 0 0.213796f
C1012 cap_res_X.n4 0 0.22697f
C1013 cap_res_X.t92 0 0.398042f
C1014 cap_res_X.t134 0 0.213796f
C1015 cap_res_X.n5 0 0.22697f
C1016 cap_res_X.t113 0 0.398042f
C1017 cap_res_X.t12 0 0.213796f
C1018 cap_res_X.n6 0 0.22697f
C1019 cap_res_X.t75 0 0.398042f
C1020 cap_res_X.t114 0 0.213796f
C1021 cap_res_X.n7 0 0.22697f
C1022 cap_res_X.t94 0 0.398042f
C1023 cap_res_X.t135 0 0.213796f
C1024 cap_res_X.n8 0 0.22697f
C1025 cap_res_X.t116 0 0.398042f
C1026 cap_res_X.t15 0 0.213796f
C1027 cap_res_X.n9 0 0.22697f
C1028 cap_res_X.t2 0 0.398042f
C1029 cap_res_X.t38 0 0.399485f
C1030 cap_res_X.t78 0 0.192435f
C1031 cap_res_X.n10 0 0.248212f
C1032 cap_res_X.t118 0 0.212473f
C1033 cap_res_X.n11 0 0.269574f
C1034 cap_res_X.t84 0 0.212473f
C1035 cap_res_X.n12 0 0.289493f
C1036 cap_res_X.t95 0 0.212473f
C1037 cap_res_X.n13 0 0.289493f
C1038 cap_res_X.t85 0 0.212473f
C1039 cap_res_X.n14 0 0.289493f
C1040 cap_res_X.t120 0 0.212473f
C1041 cap_res_X.n15 0 0.289493f
C1042 cap_res_X.t61 0 0.212473f
C1043 cap_res_X.n16 0 0.289493f
C1044 cap_res_X.t20 0 0.212473f
C1045 cap_res_X.n17 0 0.289493f
C1046 cap_res_X.t122 0 0.212473f
C1047 cap_res_X.n18 0 0.289493f
C1048 cap_res_X.t13 0 0.212473f
C1049 cap_res_X.n19 0 0.289493f
C1050 cap_res_X.t115 0 0.212473f
C1051 cap_res_X.n20 0 0.289493f
C1052 cap_res_X.t76 0 0.212473f
C1053 cap_res_X.n21 0 0.289493f
C1054 cap_res_X.t107 0 0.212473f
C1055 cap_res_X.n22 0 0.289493f
C1056 cap_res_X.t70 0 0.212473f
C1057 cap_res_X.n23 0 0.289493f
C1058 cap_res_X.t33 0 0.212473f
C1059 cap_res_X.n24 0 0.289493f
C1060 cap_res_X.t64 0 0.212473f
C1061 cap_res_X.n25 0 0.289493f
C1062 cap_res_X.t27 0 0.212473f
C1063 cap_res_X.n26 0 0.289493f
C1064 cap_res_X.t129 0 0.212473f
C1065 cap_res_X.n27 0 0.289493f
C1066 cap_res_X.t24 0 0.212473f
C1067 cap_res_X.n28 0 0.289493f
C1068 cap_res_X.t55 0 0.212473f
C1069 cap_res_X.n29 0 0.266808f
C1070 cap_res_X.t96 0 0.399485f
C1071 cap_res_X.t72 0 0.399485f
C1072 cap_res_X.t28 0 0.398042f
C1073 cap_res_X.t19 0 0.419404f
C1074 cap_res_X.t51 0 0.213796f
C1075 cap_res_X.n30 0 0.246889f
C1076 cap_res_X.t99 0 0.398042f
C1077 cap_res_X.t58 0 0.419404f
C1078 cap_res_X.t23 0 0.399485f
C1079 cap_res_X.t89 0 0.398042f
C1080 cap_res_X.t126 0 0.213796f
C1081 cap_res_X.n31 0 0.246889f
C1082 cap_res_X.t43 0 0.398042f
C1083 cap_res_X.t110 0 0.419404f
C1084 cap_res_X.t6 0 0.213796f
C1085 cap_res_X.n32 0 0.22697f
C1086 cap_res_X.t9 0 0.398042f
C1087 cap_res_X.t73 0 0.419404f
C1088 cap_res_X.t106 0 0.213796f
C1089 cap_res_X.n33 0 0.22697f
C1090 cap_res_X.t112 0 0.398042f
C1091 cap_res_X.t35 0 0.419404f
C1092 cap_res_X.t69 0 0.213796f
C1093 cap_res_X.n34 0 0.22697f
C1094 cap_res_X.n35 0 0.22697f
C1095 cap_res_X.t93 0 0.213796f
C1096 cap_res_X.t56 0 0.419404f
C1097 cap_res_X.t63 0 0.570336f
C1098 cap_res_X.t0 0 0.343308f
C1099 V_CMFB_S2.t0 0 0.31682f
C1100 V_CMFB_S2.n0 0 0.08992f
C1101 V_CMFB_S2.n1 0 0.154718f
C1102 V_CMFB_S2.t9 0 0.077555f
C1103 V_CMFB_S2.t3 0 0.077555f
C1104 V_CMFB_S2.n2 0 0.165875f
C1105 V_CMFB_S2.n3 0 0.424667f
C1106 V_CMFB_S2.n4 0 -0.31022f
C1107 V_CMFB_S2.n5 0 0.416356f
C1108 V_CMFB_S2.t10 0 0.077555f
C1109 V_CMFB_S2.t5 0 0.077555f
C1110 V_CMFB_S2.n6 0 0.165875f
C1111 V_CMFB_S2.n7 0 0.504805f
C1112 V_CMFB_S2.n8 0 0.142773f
C1113 V_CMFB_S2.n9 0 0.08992f
C1114 V_CMFB_S2.t2 0 0.077555f
C1115 V_CMFB_S2.t6 0 0.077555f
C1116 V_CMFB_S2.n10 0 0.165875f
C1117 V_CMFB_S2.n11 0 0.504805f
C1118 V_CMFB_S2.n12 0 0.08992f
C1119 V_CMFB_S2.t4 0 0.077555f
C1120 V_CMFB_S2.t8 0 0.077555f
C1121 V_CMFB_S2.n13 0 0.165875f
C1122 V_CMFB_S2.n14 0 0.504805f
C1123 V_CMFB_S2.n15 0 0.154718f
C1124 V_CMFB_S2.t1 0 0.077555f
C1125 V_CMFB_S2.t7 0 0.077555f
C1126 V_CMFB_S2.n16 0 0.165875f
C1127 V_CMFB_S2.n17 0 0.511831f
C1128 V_CMFB_S2.n18 0 0.179367f
C1129 V_CMFB_S2.n19 0 0.509529f
C1130 cap_res_Y.t72 0 0.398042f
C1131 cap_res_Y.t107 0 0.419404f
C1132 cap_res_Y.t14 0 0.399485f
C1133 cap_res_Y.t93 0 0.398042f
C1134 cap_res_Y.t127 0 0.213796f
C1135 cap_res_Y.n0 0 0.246889f
C1136 cap_res_Y.t121 0 0.398042f
C1137 cap_res_Y.t135 0 0.419404f
C1138 cap_res_Y.t27 0 0.213796f
C1139 cap_res_Y.n1 0 0.22697f
C1140 cap_res_Y.t78 0 0.398042f
C1141 cap_res_Y.t108 0 0.419404f
C1142 cap_res_Y.t11 0 0.213796f
C1143 cap_res_Y.n2 0 0.22697f
C1144 cap_res_Y.t130 0 0.398042f
C1145 cap_res_Y.t91 0 0.419404f
C1146 cap_res_Y.t123 0 0.213796f
C1147 cap_res_Y.n3 0 0.22697f
C1148 cap_res_Y.t133 0 0.398042f
C1149 cap_res_Y.t17 0 0.399485f
C1150 cap_res_Y.t63 0 0.398042f
C1151 cap_res_Y.t47 0 0.399485f
C1152 cap_res_Y.t98 0 0.398042f
C1153 cap_res_Y.t114 0 0.399485f
C1154 cap_res_Y.t95 0 0.398042f
C1155 cap_res_Y.t9 0 0.399485f
C1156 cap_res_Y.t126 0 0.398042f
C1157 cap_res_Y.t74 0 0.399485f
C1158 cap_res_Y.t137 0 0.398042f
C1159 cap_res_Y.t52 0 0.399485f
C1160 cap_res_Y.t30 0 0.398042f
C1161 cap_res_Y.t112 0 0.399485f
C1162 cap_res_Y.t38 0 0.398042f
C1163 cap_res_Y.t87 0 0.399485f
C1164 cap_res_Y.t65 0 0.398042f
C1165 cap_res_Y.t18 0 0.399485f
C1166 cap_res_Y.t5 0 0.398042f
C1167 cap_res_Y.t56 0 0.399485f
C1168 cap_res_Y.t35 0 0.398042f
C1169 cap_res_Y.t118 0 0.399485f
C1170 cap_res_Y.t44 0 0.398042f
C1171 cap_res_Y.t92 0 0.399485f
C1172 cap_res_Y.t70 0 0.398042f
C1173 cap_res_Y.t22 0 0.399485f
C1174 cap_res_Y.t79 0 0.398042f
C1175 cap_res_Y.t132 0 0.399485f
C1176 cap_res_Y.t106 0 0.398042f
C1177 cap_res_Y.t59 0 0.399485f
C1178 cap_res_Y.t51 0 0.398042f
C1179 cap_res_Y.t99 0 0.399485f
C1180 cap_res_Y.t75 0 0.398042f
C1181 cap_res_Y.t28 0 0.399485f
C1182 cap_res_Y.t85 0 0.398042f
C1183 cap_res_Y.t1 0 0.399485f
C1184 cap_res_Y.t113 0 0.398042f
C1185 cap_res_Y.t64 0 0.399485f
C1186 cap_res_Y.t122 0 0.398042f
C1187 cap_res_Y.t39 0 0.399485f
C1188 cap_res_Y.t19 0 0.398042f
C1189 cap_res_Y.t104 0 0.399485f
C1190 cap_res_Y.t90 0 0.398042f
C1191 cap_res_Y.t6 0 0.399485f
C1192 cap_res_Y.t119 0 0.398042f
C1193 cap_res_Y.t68 0 0.399485f
C1194 cap_res_Y.t131 0 0.398042f
C1195 cap_res_Y.t45 0 0.399485f
C1196 cap_res_Y.t23 0 0.398042f
C1197 cap_res_Y.t105 0 0.399485f
C1198 cap_res_Y.t32 0 0.398042f
C1199 cap_res_Y.t81 0 0.399485f
C1200 cap_res_Y.t61 0 0.398042f
C1201 cap_res_Y.t15 0 0.399485f
C1202 cap_res_Y.t3 0 0.398042f
C1203 cap_res_Y.t43 0 0.399485f
C1204 cap_res_Y.t116 0 0.398042f
C1205 cap_res_Y.t77 0 0.399485f
C1206 cap_res_Y.t102 0 0.398042f
C1207 cap_res_Y.t8 0 0.399485f
C1208 cap_res_Y.t86 0 0.398042f
C1209 cap_res_Y.t48 0 0.399485f
C1210 cap_res_Y.t62 0 0.398042f
C1211 cap_res_Y.t110 0 0.399485f
C1212 cap_res_Y.t97 0 0.398042f
C1213 cap_res_Y.t50 0 0.399485f
C1214 cap_res_Y.t124 0 0.398042f
C1215 cap_res_Y.t103 0 0.399485f
C1216 cap_res_Y.t20 0 0.398042f
C1217 cap_res_Y.t42 0 0.399485f
C1218 cap_res_Y.t96 0 0.398042f
C1219 cap_res_Y.t138 0 0.417559f
C1220 cap_res_Y.t136 0 0.398042f
C1221 cap_res_Y.t36 0 0.213796f
C1222 cap_res_Y.n4 0 0.228815f
C1223 cap_res_Y.t34 0 0.398042f
C1224 cap_res_Y.t69 0 0.213796f
C1225 cap_res_Y.n5 0 0.22697f
C1226 cap_res_Y.t12 0 0.398042f
C1227 cap_res_Y.t55 0 0.213796f
C1228 cap_res_Y.n6 0 0.22697f
C1229 cap_res_Y.t54 0 0.398042f
C1230 cap_res_Y.t89 0 0.213796f
C1231 cap_res_Y.n7 0 0.22697f
C1232 cap_res_Y.t31 0 0.398042f
C1233 cap_res_Y.t66 0 0.213796f
C1234 cap_res_Y.n8 0 0.22697f
C1235 cap_res_Y.t10 0 0.398042f
C1236 cap_res_Y.t53 0 0.213796f
C1237 cap_res_Y.n9 0 0.22697f
C1238 cap_res_Y.t49 0 0.398042f
C1239 cap_res_Y.t84 0 0.213796f
C1240 cap_res_Y.n10 0 0.22697f
C1241 cap_res_Y.t83 0 0.398042f
C1242 cap_res_Y.t120 0 0.213796f
C1243 cap_res_Y.n11 0 0.22697f
C1244 cap_res_Y.t115 0 0.398042f
C1245 cap_res_Y.t21 0 0.213796f
C1246 cap_res_Y.n12 0 0.22697f
C1247 cap_res_Y.t100 0 0.398042f
C1248 cap_res_Y.t4 0 0.213796f
C1249 cap_res_Y.n13 0 0.22697f
C1250 cap_res_Y.t57 0 0.398042f
C1251 cap_res_Y.t71 0 0.399485f
C1252 cap_res_Y.t16 0 0.398042f
C1253 cap_res_Y.t37 0 0.399485f
C1254 cap_res_Y.t2 0 0.192435f
C1255 cap_res_Y.n14 0 0.248212f
C1256 cap_res_Y.t41 0 0.212473f
C1257 cap_res_Y.n15 0 0.269574f
C1258 cap_res_Y.t7 0 0.212473f
C1259 cap_res_Y.n16 0 0.289493f
C1260 cap_res_Y.t13 0 0.212473f
C1261 cap_res_Y.n17 0 0.289493f
C1262 cap_res_Y.t94 0 0.212473f
C1263 cap_res_Y.n18 0 0.289493f
C1264 cap_res_Y.t129 0 0.212473f
C1265 cap_res_Y.n19 0 0.289493f
C1266 cap_res_Y.t111 0 0.212473f
C1267 cap_res_Y.n20 0 0.289493f
C1268 cap_res_Y.t73 0 0.212473f
C1269 cap_res_Y.n21 0 0.289493f
C1270 cap_res_Y.t40 0 0.212473f
C1271 cap_res_Y.n22 0 0.289493f
C1272 cap_res_Y.t67 0 0.212473f
C1273 cap_res_Y.n23 0 0.289493f
C1274 cap_res_Y.t33 0 0.212473f
C1275 cap_res_Y.n24 0 0.289493f
C1276 cap_res_Y.t134 0 0.212473f
C1277 cap_res_Y.n25 0 0.289493f
C1278 cap_res_Y.t26 0 0.212473f
C1279 cap_res_Y.n26 0 0.289493f
C1280 cap_res_Y.t125 0 0.212473f
C1281 cap_res_Y.n27 0 0.289493f
C1282 cap_res_Y.t88 0 0.212473f
C1283 cap_res_Y.n28 0 0.289493f
C1284 cap_res_Y.t117 0 0.212473f
C1285 cap_res_Y.n29 0 0.289493f
C1286 cap_res_Y.t82 0 0.212473f
C1287 cap_res_Y.n30 0 0.289493f
C1288 cap_res_Y.t46 0 0.212473f
C1289 cap_res_Y.n31 0 0.289493f
C1290 cap_res_Y.t80 0 0.212473f
C1291 cap_res_Y.n32 0 0.289493f
C1292 cap_res_Y.t109 0 0.212473f
C1293 cap_res_Y.n33 0 0.266808f
C1294 cap_res_Y.t76 0 0.399485f
C1295 cap_res_Y.t101 0 0.399485f
C1296 cap_res_Y.t58 0 0.398042f
C1297 cap_res_Y.t29 0 0.419404f
C1298 cap_res_Y.t60 0 0.213796f
C1299 cap_res_Y.n34 0 0.246889f
C1300 cap_res_Y.n35 0 0.22697f
C1301 cap_res_Y.t24 0 0.213796f
C1302 cap_res_Y.t128 0 0.419404f
C1303 cap_res_Y.t25 0 0.570336f
C1304 cap_res_Y.t0 0 0.34331f
C1305 VOUT+.n0 0 0.0754f
C1306 VOUT+.n2 0 0.038454f
C1307 VOUT+.n6 0 0.036192f
C1308 VOUT+.n7 0 0.038454f
C1309 VOUT+.n8 0 0.036192f
C1310 VOUT+.t8 0 0.05278f
C1311 VOUT+.t10 0 0.05278f
C1312 VOUT+.n9 0 0.113404f
C1313 VOUT+.n10 0 0.272735f
C1314 VOUT+.n11 0 0.036192f
C1315 VOUT+.n12 0 0.23372f
C1316 VOUT+.t11 0 0.05278f
C1317 VOUT+.t9 0 0.05278f
C1318 VOUT+.n13 0 0.113404f
C1319 VOUT+.n14 0 0.282262f
C1320 VOUT+.n15 0 0.161339f
C1321 VOUT+.t7 0 0.05278f
C1322 VOUT+.t6 0 0.05278f
C1323 VOUT+.n16 0 0.113404f
C1324 VOUT+.n17 0 0.268146f
C1325 VOUT+.n18 0 0.12306f
C1326 VOUT+.n19 0 0.036192f
C1327 VOUT+.n20 0 0.186755f
C1328 VOUT+.n21 0 0.036192f
C1329 VOUT+.n22 0 0.036192f
C1330 VOUT+.n23 0 0.036192f
C1331 VOUT+.n24 0 0.036192f
C1332 VOUT+.n25 0 0.077474f
C1333 VOUT+.n26 0 0.183223f
C1334 VOUT+.t0 0 0.086088f
C1335 VOUT+.n27 0 0.330876f
C1336 VOUT+.n28 0 0.038454f
C1337 VOUT+.n31 0 0.05655f
C1338 VOUT+.n32 0 0.09425f
C1339 VOUT+.n33 0 0.059913f
C1340 VOUT+.n34 0 0.05655f
C1341 VOUT+.n36 0 0.038454f
C1342 VOUT+.n37 0 0.035853f
C1343 VOUT+.n38 0 0.038454f
C1344 VOUT+.n39 0 0.049764f
C1345 VOUT+.n40 0 0.071798f
C1346 VOUT+.n41 0 0.069871f
C1347 VOUT+.n42 0 0.049764f
C1348 VOUT+.n43 0 0.049764f
C1349 VOUT+.n44 0 0.069871f
C1350 VOUT+.n45 0 0.069871f
C1351 VOUT+.n46 0 0.049764f
C1352 VOUT+.n47 0 0.079669f
C1353 VOUT+.t12 0 0.04524f
C1354 VOUT+.t14 0 0.04524f
C1355 VOUT+.n48 0 0.092697f
C1356 VOUT+.n49 0 0.239278f
C1357 VOUT+.t2 0 0.04524f
C1358 VOUT+.t13 0 0.04524f
C1359 VOUT+.n50 0 0.092697f
C1360 VOUT+.n51 0 0.239278f
C1361 VOUT+.t4 0 0.04524f
C1362 VOUT+.t3 0 0.04524f
C1363 VOUT+.n52 0 0.092697f
C1364 VOUT+.n53 0 0.236867f
C1365 VOUT+.n54 0 0.057528f
C1366 VOUT+.t5 0 0.04524f
C1367 VOUT+.t17 0 0.04524f
C1368 VOUT+.n55 0 0.092697f
C1369 VOUT+.n56 0 0.236867f
C1370 VOUT+.n57 0 0.032609f
C1371 VOUT+.t15 0 0.04524f
C1372 VOUT+.t18 0 0.04524f
C1373 VOUT+.n58 0 0.092697f
C1374 VOUT+.n59 0 0.236867f
C1375 VOUT+.n60 0 0.032609f
C1376 VOUT+.n61 0 0.057528f
C1377 VOUT+.t16 0 0.04524f
C1378 VOUT+.t1 0 0.04524f
C1379 VOUT+.n62 0 0.092697f
C1380 VOUT+.n63 0 0.236867f
C1381 VOUT+.n64 0 0.038035f
C1382 VOUT+.n65 0 0.02262f
C1383 VOUT+.n66 0 0.02262f
C1384 VOUT+.n67 0 0.038035f
C1385 VOUT+.n68 0 0.069871f
C1386 VOUT+.n69 0 0.097805f
C1387 VOUT+.n70 0 0.12187f
C1388 VOUT+.n71 0 0.170568f
C1389 VOUT+.n72 0 0.049764f
C1390 VOUT+.n73 0 0.081432f
C1391 VOUT+.n74 0 0.049764f
C1392 VOUT+.n75 0 0.081432f
C1393 VOUT+.n76 0 0.049764f
C1394 VOUT+.n77 0 0.049764f
C1395 VOUT+.n78 0 0.049764f
C1396 VOUT+.n79 0 0.081432f
C1397 VOUT+.n80 0 0.049764f
C1398 VOUT+.n81 0 0.074646f
C1399 VOUT+.n82 0 0.239773f
C1400 VOUT+.n84 0 0.0754f
C1401 VOUT+.n85 0 0.038454f
C1402 VOUT+.n87 0 0.038454f
C1403 VOUT+.n90 0 0.0754f
C1404 VOUT+.n91 0 0.232987f
C1405 VOUT+.n92 0 0.537227f
C1406 VOUT+.n95 0 0.05655f
C1407 VOUT+.n96 0 0.05655f
C1408 VOUT+.n97 0 0.05655f
C1409 VOUT+.n98 0 0.05655f
C1410 VOUT+.n99 0 0.165871f
C1411 VOUT+.n100 0 0.05655f
C1412 VOUT+.t155 0 0.301601f
C1413 VOUT+.t141 0 0.306738f
C1414 VOUT+.t120 0 0.301601f
C1415 VOUT+.n101 0 0.202214f
C1416 VOUT+.n102 0 0.13195f
C1417 VOUT+.t57 0 0.306095f
C1418 VOUT+.t42 0 0.306095f
C1419 VOUT+.t74 0 0.306095f
C1420 VOUT+.t108 0 0.306095f
C1421 VOUT+.t147 0 0.306095f
C1422 VOUT+.t126 0 0.306095f
C1423 VOUT+.t103 0 0.306095f
C1424 VOUT+.t145 0 0.306095f
C1425 VOUT+.t123 0 0.306095f
C1426 VOUT+.t21 0 0.306095f
C1427 VOUT+.t61 0 0.306095f
C1428 VOUT+.t19 0 0.301601f
C1429 VOUT+.n103 0 0.202857f
C1430 VOUT+.t121 0 0.301601f
C1431 VOUT+.n104 0 0.259407f
C1432 VOUT+.t88 0 0.301601f
C1433 VOUT+.n105 0 0.259407f
C1434 VOUT+.t102 0 0.301601f
C1435 VOUT+.n106 0 0.259407f
C1436 VOUT+.t68 0 0.301601f
C1437 VOUT+.n107 0 0.259407f
C1438 VOUT+.t91 0 0.301601f
C1439 VOUT+.n108 0 0.259407f
C1440 VOUT+.t104 0 0.301601f
C1441 VOUT+.n109 0 0.259407f
C1442 VOUT+.t73 0 0.301601f
C1443 VOUT+.n110 0 0.259407f
C1444 VOUT+.t37 0 0.301601f
C1445 VOUT+.n111 0 0.259407f
C1446 VOUT+.t136 0 0.301601f
C1447 VOUT+.n112 0 0.259407f
C1448 VOUT+.t153 0 0.301601f
C1449 VOUT+.n113 0 0.259407f
C1450 VOUT+.t116 0 0.301601f
C1451 VOUT+.t100 0 0.306738f
C1452 VOUT+.t86 0 0.301601f
C1453 VOUT+.n114 0 0.202214f
C1454 VOUT+.n115 0 0.245051f
C1455 VOUT+.t33 0 0.306738f
C1456 VOUT+.t54 0 0.301601f
C1457 VOUT+.n116 0 0.202214f
C1458 VOUT+.t150 0 0.301601f
C1459 VOUT+.t137 0 0.306738f
C1460 VOUT+.t115 0 0.301601f
C1461 VOUT+.n117 0 0.202214f
C1462 VOUT+.n118 0 0.245051f
C1463 VOUT+.t95 0 0.306738f
C1464 VOUT+.t47 0 0.301601f
C1465 VOUT+.n119 0 0.202214f
C1466 VOUT+.t144 0 0.301601f
C1467 VOUT+.t60 0 0.306738f
C1468 VOUT+.t107 0 0.301601f
C1469 VOUT+.n120 0 0.202214f
C1470 VOUT+.n121 0 0.245051f
C1471 VOUT+.t55 0 0.306738f
C1472 VOUT+.t149 0 0.301601f
C1473 VOUT+.n122 0 0.202214f
C1474 VOUT+.t63 0 0.301601f
C1475 VOUT+.t71 0 0.306738f
C1476 VOUT+.t109 0 0.301601f
C1477 VOUT+.n123 0 0.202214f
C1478 VOUT+.n124 0 0.245051f
C1479 VOUT+.t154 0 0.306738f
C1480 VOUT+.t114 0 0.301601f
C1481 VOUT+.n125 0 0.202214f
C1482 VOUT+.t28 0 0.301601f
C1483 VOUT+.t41 0 0.306738f
C1484 VOUT+.t80 0 0.301601f
C1485 VOUT+.n126 0 0.202214f
C1486 VOUT+.n127 0 0.245051f
C1487 VOUT+.t125 0 0.306738f
C1488 VOUT+.t76 0 0.301601f
C1489 VOUT+.n128 0 0.202214f
C1490 VOUT+.t46 0 0.301601f
C1491 VOUT+.t96 0 0.306738f
C1492 VOUT+.t142 0 0.301601f
C1493 VOUT+.n129 0 0.202214f
C1494 VOUT+.n130 0 0.245051f
C1495 VOUT+.t26 0 0.306738f
C1496 VOUT+.t112 0 0.301601f
C1497 VOUT+.n131 0 0.202214f
C1498 VOUT+.t84 0 0.301601f
C1499 VOUT+.t134 0 0.306738f
C1500 VOUT+.t52 0 0.301601f
C1501 VOUT+.n132 0 0.202214f
C1502 VOUT+.n133 0 0.245051f
C1503 VOUT+.t99 0 0.306738f
C1504 VOUT+.t128 0 0.301601f
C1505 VOUT+.n134 0 0.197501f
C1506 VOUT+.t132 0 0.306738f
C1507 VOUT+.t29 0 0.301601f
C1508 VOUT+.n135 0 0.197501f
C1509 VOUT+.t27 0 0.306738f
C1510 VOUT+.t66 0 0.301601f
C1511 VOUT+.n136 0 0.197501f
C1512 VOUT+.t79 0 0.306738f
C1513 VOUT+.t49 0 0.301601f
C1514 VOUT+.n137 0 0.197501f
C1515 VOUT+.t36 0 0.306738f
C1516 VOUT+.t22 0 0.301601f
C1517 VOUT+.n138 0 0.199386f
C1518 VOUT+.t64 0 0.306347f
C1519 VOUT+.t85 0 0.306738f
C1520 VOUT+.t50 0 0.301601f
C1521 VOUT+.n139 0 0.202214f
C1522 VOUT+.t143 0 0.301601f
C1523 VOUT+.n140 0 0.13195f
C1524 VOUT+.t30 0 0.301601f
C1525 VOUT+.n141 0 0.262925f
C1526 VOUT+.t130 0 0.301601f
C1527 VOUT+.n142 0 0.195098f
C1528 VOUT+.t146 0 0.301601f
C1529 VOUT+.n143 0 0.193213f
C1530 VOUT+.t34 0 0.301601f
C1531 VOUT+.n144 0 0.193213f
C1532 VOUT+.t133 0 0.301601f
C1533 VOUT+.n145 0 0.193213f
C1534 VOUT+.t97 0 0.301601f
C1535 VOUT+.n146 0 0.193213f
C1536 VOUT+.t56 0 0.301601f
C1537 VOUT+.n147 0 0.13195f
C1538 VOUT+.t81 0 0.301601f
C1539 VOUT+.n148 0 0.13195f
C1540 VOUT+.t48 0 0.301601f
C1541 VOUT+.t24 0 0.306738f
C1542 VOUT+.t140 0 0.301601f
C1543 VOUT+.n149 0 0.202214f
C1544 VOUT+.n150 0 0.188501f
C1545 VOUT+.t94 0 0.306738f
C1546 VOUT+.t110 0 0.301601f
C1547 VOUT+.n151 0 0.202214f
C1548 VOUT+.t77 0 0.301601f
C1549 VOUT+.t59 0 0.306738f
C1550 VOUT+.t43 0 0.301601f
C1551 VOUT+.n152 0 0.202214f
C1552 VOUT+.n153 0 0.245051f
C1553 VOUT+.t62 0 0.306738f
C1554 VOUT+.t148 0 0.301601f
C1555 VOUT+.n154 0 0.202214f
C1556 VOUT+.t111 0 0.301601f
C1557 VOUT+.t31 0 0.306738f
C1558 VOUT+.t83 0 0.301601f
C1559 VOUT+.n155 0 0.202214f
C1560 VOUT+.n156 0 0.245051f
C1561 VOUT+.t20 0 0.306738f
C1562 VOUT+.t105 0 0.301601f
C1563 VOUT+.n157 0 0.202214f
C1564 VOUT+.t75 0 0.301601f
C1565 VOUT+.t127 0 0.306738f
C1566 VOUT+.t45 0 0.301601f
C1567 VOUT+.n158 0 0.202214f
C1568 VOUT+.n159 0 0.245051f
C1569 VOUT+.t119 0 0.306738f
C1570 VOUT+.t70 0 0.301601f
C1571 VOUT+.n160 0 0.202214f
C1572 VOUT+.t40 0 0.301601f
C1573 VOUT+.t92 0 0.306738f
C1574 VOUT+.t139 0 0.301601f
C1575 VOUT+.n161 0 0.202214f
C1576 VOUT+.n162 0 0.245051f
C1577 VOUT+.t152 0 0.306738f
C1578 VOUT+.t101 0 0.301601f
C1579 VOUT+.n163 0 0.202214f
C1580 VOUT+.t69 0 0.301601f
C1581 VOUT+.t122 0 0.306738f
C1582 VOUT+.t39 0 0.301601f
C1583 VOUT+.n164 0 0.202214f
C1584 VOUT+.n165 0 0.245051f
C1585 VOUT+.t113 0 0.306738f
C1586 VOUT+.t65 0 0.301601f
C1587 VOUT+.n166 0 0.202214f
C1588 VOUT+.t32 0 0.301601f
C1589 VOUT+.t87 0 0.306738f
C1590 VOUT+.t135 0 0.301601f
C1591 VOUT+.n167 0 0.202214f
C1592 VOUT+.n168 0 0.245051f
C1593 VOUT+.t78 0 0.306738f
C1594 VOUT+.t25 0 0.301601f
C1595 VOUT+.n169 0 0.202214f
C1596 VOUT+.t131 0 0.301601f
C1597 VOUT+.t51 0 0.306738f
C1598 VOUT+.t98 0 0.301601f
C1599 VOUT+.n170 0 0.202214f
C1600 VOUT+.n171 0 0.245051f
C1601 VOUT+.t106 0 0.306738f
C1602 VOUT+.t58 0 0.301601f
C1603 VOUT+.n172 0 0.202214f
C1604 VOUT+.t23 0 0.301601f
C1605 VOUT+.t82 0 0.306738f
C1606 VOUT+.t129 0 0.301601f
C1607 VOUT+.n173 0 0.202214f
C1608 VOUT+.n174 0 0.245051f
C1609 VOUT+.t72 0 0.306738f
C1610 VOUT+.t156 0 0.301601f
C1611 VOUT+.n175 0 0.202214f
C1612 VOUT+.t124 0 0.301601f
C1613 VOUT+.t44 0 0.306738f
C1614 VOUT+.t93 0 0.301601f
C1615 VOUT+.n176 0 0.202214f
C1616 VOUT+.n177 0 0.245051f
C1617 VOUT+.t35 0 0.306738f
C1618 VOUT+.t118 0 0.301601f
C1619 VOUT+.n178 0 0.202214f
C1620 VOUT+.t90 0 0.301601f
C1621 VOUT+.t138 0 0.306738f
C1622 VOUT+.t53 0 0.301601f
C1623 VOUT+.n179 0 0.202214f
C1624 VOUT+.n180 0 0.245051f
C1625 VOUT+.t38 0 0.306738f
C1626 VOUT+.t89 0 0.301601f
C1627 VOUT+.n181 0 0.202214f
C1628 VOUT+.t117 0 0.301601f
C1629 VOUT+.n182 0 0.245051f
C1630 VOUT+.t151 0 0.301601f
C1631 VOUT+.n183 0 0.129123f
C1632 VOUT+.t67 0 0.301601f
C1633 VOUT+.n184 0 0.336474f
C1634 VOUT+.n185 0 0.277096f
C1635 VOUT+.n186 0 0.05655f
C1636 VOUT+.n187 0 0.05655f
C1637 VOUT+.n189 0 0.546652f
C1638 VOUT+.n190 0 0.056967f
C1639 VOUT+.n191 0 1.12158f
C1640 VOUT+.n192 0 1.11215f
C1641 VOUT+.n194 0 0.10179f
C1642 VOUT+.n195 0 0.0754f
C1643 V_b_2nd_stage.t1 0 0.155439f
C1644 V_b_2nd_stage.t6 0 0.385095f
C1645 V_b_2nd_stage.t4 0 0.457048f
C1646 V_b_2nd_stage.t9 0 0.385095f
C1647 V_b_2nd_stage.t5 0 0.457048f
C1648 V_b_2nd_stage.n0 0 0.241409f
C1649 V_b_2nd_stage.n1 0 0.271017f
C1650 V_b_2nd_stage.n2 0 0.847851f
C1651 V_b_2nd_stage.t2 0 0.385095f
C1652 V_b_2nd_stage.t8 0 0.385095f
C1653 V_b_2nd_stage.t3 0 0.457048f
C1654 V_b_2nd_stage.n3 0 0.241409f
C1655 V_b_2nd_stage.t7 0 0.457048f
C1656 V_b_2nd_stage.n4 0 0.271017f
C1657 V_b_2nd_stage.n5 0 0.847851f
C1658 V_b_2nd_stage.t0 0 0.155439f
C1659 VOUT-.n1 0 0.038505f
C1660 VOUT-.n3 0 0.038505f
C1661 VOUT-.n5 0 0.075499f
C1662 VOUT-.n6 0 0.038505f
C1663 VOUT-.n9 0 0.056624f
C1664 VOUT-.n10 0 0.094374f
C1665 VOUT-.n11 0 0.056624f
C1666 VOUT-.n12 0 0.056624f
C1667 VOUT-.n14 0 0.038505f
C1668 VOUT-.n16 0 0.038505f
C1669 VOUT-.n18 0 0.075499f
C1670 VOUT-.n19 0 0.038505f
C1671 VOUT-.n21 0 0.038505f
C1672 VOUT-.n23 0 0.049829f
C1673 VOUT-.n24 0 0.071892f
C1674 VOUT-.n25 0 0.069963f
C1675 VOUT-.n26 0 0.049829f
C1676 VOUT-.n27 0 0.049829f
C1677 VOUT-.n28 0 0.069963f
C1678 VOUT-.n29 0 0.069963f
C1679 VOUT-.n30 0 0.049829f
C1680 VOUT-.n31 0 0.079773f
C1681 VOUT-.t16 0 0.0453f
C1682 VOUT-.t15 0 0.0453f
C1683 VOUT-.n32 0 0.092819f
C1684 VOUT-.n33 0 0.239593f
C1685 VOUT-.t11 0 0.0453f
C1686 VOUT-.t8 0 0.0453f
C1687 VOUT-.n34 0 0.092819f
C1688 VOUT-.n35 0 0.237178f
C1689 VOUT-.n36 0 0.057603f
C1690 VOUT-.t12 0 0.0453f
C1691 VOUT-.t6 0 0.0453f
C1692 VOUT-.n37 0 0.092819f
C1693 VOUT-.n38 0 0.237178f
C1694 VOUT-.n39 0 0.032651f
C1695 VOUT-.t10 0 0.0453f
C1696 VOUT-.t14 0 0.0453f
C1697 VOUT-.n40 0 0.092819f
C1698 VOUT-.n41 0 0.237178f
C1699 VOUT-.n42 0 0.032651f
C1700 VOUT-.t7 0 0.0453f
C1701 VOUT-.t17 0 0.0453f
C1702 VOUT-.n43 0 0.092819f
C1703 VOUT-.n44 0 0.239593f
C1704 VOUT-.n45 0 0.057603f
C1705 VOUT-.t9 0 0.0453f
C1706 VOUT-.t13 0 0.0453f
C1707 VOUT-.n46 0 0.092819f
C1708 VOUT-.n47 0 0.237178f
C1709 VOUT-.n48 0 0.038085f
C1710 VOUT-.n49 0 0.02265f
C1711 VOUT-.n50 0 0.02265f
C1712 VOUT-.n51 0 0.038085f
C1713 VOUT-.n52 0 0.069963f
C1714 VOUT-.n53 0 0.097934f
C1715 VOUT-.n54 0 0.12203f
C1716 VOUT-.n55 0 0.170792f
C1717 VOUT-.n56 0 0.049829f
C1718 VOUT-.n57 0 0.081539f
C1719 VOUT-.n58 0 0.049829f
C1720 VOUT-.n59 0 0.081539f
C1721 VOUT-.n60 0 0.049829f
C1722 VOUT-.n61 0 0.049829f
C1723 VOUT-.n62 0 0.049829f
C1724 VOUT-.n63 0 0.081539f
C1725 VOUT-.n64 0 0.049829f
C1726 VOUT-.n65 0 0.074744f
C1727 VOUT-.n66 0 0.240088f
C1728 VOUT-.n67 0 0.233293f
C1729 VOUT-.n69 0 0.075499f
C1730 VOUT-.n70 0 0.03624f
C1731 VOUT-.n71 0 0.537932f
C1732 VOUT-.n74 0 0.056624f
C1733 VOUT-.n75 0 0.056624f
C1734 VOUT-.t155 0 0.307141f
C1735 VOUT-.t119 0 0.301997f
C1736 VOUT-.n76 0 0.202479f
C1737 VOUT-.t79 0 0.301997f
C1738 VOUT-.n77 0 0.132124f
C1739 VOUT-.t115 0 0.307141f
C1740 VOUT-.t78 0 0.301997f
C1741 VOUT-.n78 0 0.202479f
C1742 VOUT-.t39 0 0.301997f
C1743 VOUT-.t41 0 0.306497f
C1744 VOUT-.t63 0 0.306497f
C1745 VOUT-.t82 0 0.306497f
C1746 VOUT-.t44 0 0.306497f
C1747 VOUT-.t65 0 0.306497f
C1748 VOUT-.t27 0 0.306497f
C1749 VOUT-.t128 0 0.306497f
C1750 VOUT-.t154 0 0.306497f
C1751 VOUT-.t113 0 0.306497f
C1752 VOUT-.t76 0 0.306497f
C1753 VOUT-.t38 0 0.306497f
C1754 VOUT-.t140 0 0.301997f
C1755 VOUT-.n79 0 0.203123f
C1756 VOUT-.t34 0 0.301997f
C1757 VOUT-.n80 0 0.259748f
C1758 VOUT-.t74 0 0.301997f
C1759 VOUT-.n81 0 0.259748f
C1760 VOUT-.t112 0 0.301997f
C1761 VOUT-.n82 0 0.259748f
C1762 VOUT-.t90 0 0.301997f
C1763 VOUT-.n83 0 0.259748f
C1764 VOUT-.t127 0 0.301997f
C1765 VOUT-.n84 0 0.259748f
C1766 VOUT-.t23 0 0.301997f
C1767 VOUT-.n85 0 0.259748f
C1768 VOUT-.t145 0 0.301997f
C1769 VOUT-.n86 0 0.259748f
C1770 VOUT-.t43 0 0.301997f
C1771 VOUT-.n87 0 0.259748f
C1772 VOUT-.t22 0 0.301997f
C1773 VOUT-.n88 0 0.259748f
C1774 VOUT-.t142 0 0.301997f
C1775 VOUT-.n89 0 0.259748f
C1776 VOUT-.n90 0 0.245373f
C1777 VOUT-.t149 0 0.307141f
C1778 VOUT-.t111 0 0.301997f
C1779 VOUT-.n91 0 0.202479f
C1780 VOUT-.t73 0 0.301997f
C1781 VOUT-.t57 0 0.307141f
C1782 VOUT-.t33 0 0.301997f
C1783 VOUT-.n92 0 0.202479f
C1784 VOUT-.n93 0 0.245373f
C1785 VOUT-.t132 0 0.307141f
C1786 VOUT-.t100 0 0.301997f
C1787 VOUT-.n94 0 0.202479f
C1788 VOUT-.t62 0 0.301997f
C1789 VOUT-.t116 0 0.307141f
C1790 VOUT-.t26 0 0.301997f
C1791 VOUT-.n95 0 0.202479f
C1792 VOUT-.n96 0 0.245373f
C1793 VOUT-.t109 0 0.307141f
C1794 VOUT-.t19 0 0.301997f
C1795 VOUT-.n97 0 0.202479f
C1796 VOUT-.t72 0 0.301997f
C1797 VOUT-.t80 0 0.307141f
C1798 VOUT-.t123 0 0.301997f
C1799 VOUT-.n98 0 0.202479f
C1800 VOUT-.n99 0 0.245373f
C1801 VOUT-.t75 0 0.307141f
C1802 VOUT-.t126 0 0.301997f
C1803 VOUT-.n100 0 0.202479f
C1804 VOUT-.t37 0 0.301997f
C1805 VOUT-.t48 0 0.307141f
C1806 VOUT-.t89 0 0.301997f
C1807 VOUT-.n101 0 0.202479f
C1808 VOUT-.n102 0 0.245373f
C1809 VOUT-.t25 0 0.307141f
C1810 VOUT-.t131 0 0.301997f
C1811 VOUT-.n103 0 0.202479f
C1812 VOUT-.t96 0 0.301997f
C1813 VOUT-.t150 0 0.307141f
C1814 VOUT-.t59 0 0.301997f
C1815 VOUT-.n104 0 0.202479f
C1816 VOUT-.n105 0 0.245373f
C1817 VOUT-.t67 0 0.307141f
C1818 VOUT-.t29 0 0.301997f
C1819 VOUT-.n106 0 0.202479f
C1820 VOUT-.t137 0 0.301997f
C1821 VOUT-.t52 0 0.307141f
C1822 VOUT-.t104 0 0.301997f
C1823 VOUT-.n107 0 0.202479f
C1824 VOUT-.n108 0 0.245373f
C1825 VOUT-.t32 0 0.307141f
C1826 VOUT-.t139 0 0.301997f
C1827 VOUT-.n109 0 0.202479f
C1828 VOUT-.t102 0 0.301997f
C1829 VOUT-.t129 0 0.307141f
C1830 VOUT-.t138 0 0.301997f
C1831 VOUT-.n110 0 0.19776f
C1832 VOUT-.t94 0 0.307141f
C1833 VOUT-.t101 0 0.301997f
C1834 VOUT-.n111 0 0.19776f
C1835 VOUT-.t45 0 0.307141f
C1836 VOUT-.t122 0 0.301997f
C1837 VOUT-.n112 0 0.19776f
C1838 VOUT-.t148 0 0.307141f
C1839 VOUT-.t84 0 0.301997f
C1840 VOUT-.n113 0 0.19776f
C1841 VOUT-.t114 0 0.307141f
C1842 VOUT-.t47 0 0.301997f
C1843 VOUT-.n114 0 0.199648f
C1844 VOUT-.t68 0 0.30675f
C1845 VOUT-.t58 0 0.307141f
C1846 VOUT-.t99 0 0.301997f
C1847 VOUT-.n115 0 0.202479f
C1848 VOUT-.t134 0 0.301997f
C1849 VOUT-.n116 0 0.132124f
C1850 VOUT-.t31 0 0.301997f
C1851 VOUT-.n117 0 0.26327f
C1852 VOUT-.t151 0 0.301997f
C1853 VOUT-.n118 0 0.195354f
C1854 VOUT-.t51 0 0.301997f
C1855 VOUT-.n119 0 0.193467f
C1856 VOUT-.t88 0 0.301997f
C1857 VOUT-.n120 0 0.193467f
C1858 VOUT-.t64 0 0.301997f
C1859 VOUT-.n121 0 0.193467f
C1860 VOUT-.t106 0 0.301997f
C1861 VOUT-.n122 0 0.193467f
C1862 VOUT-.t85 0 0.301997f
C1863 VOUT-.n123 0 0.132124f
C1864 VOUT-.t61 0 0.301997f
C1865 VOUT-.n124 0 0.132124f
C1866 VOUT-.n125 0 0.188748f
C1867 VOUT-.t69 0 0.307141f
C1868 VOUT-.t30 0 0.301997f
C1869 VOUT-.n126 0 0.202479f
C1870 VOUT-.t133 0 0.301997f
C1871 VOUT-.t120 0 0.307141f
C1872 VOUT-.t98 0 0.301997f
C1873 VOUT-.n127 0 0.202479f
C1874 VOUT-.n128 0 0.245373f
C1875 VOUT-.t105 0 0.307141f
C1876 VOUT-.t66 0 0.301997f
C1877 VOUT-.n129 0 0.202479f
C1878 VOUT-.t28 0 0.301997f
C1879 VOUT-.t86 0 0.307141f
C1880 VOUT-.t136 0 0.301997f
C1881 VOUT-.n130 0 0.202479f
C1882 VOUT-.n131 0 0.245373f
C1883 VOUT-.t60 0 0.307141f
C1884 VOUT-.t24 0 0.301997f
C1885 VOUT-.n132 0 0.202479f
C1886 VOUT-.t130 0 0.301997f
C1887 VOUT-.t46 0 0.307141f
C1888 VOUT-.t97 0 0.301997f
C1889 VOUT-.n133 0 0.202479f
C1890 VOUT-.n134 0 0.245373f
C1891 VOUT-.t21 0 0.307141f
C1892 VOUT-.t125 0 0.301997f
C1893 VOUT-.n135 0 0.202479f
C1894 VOUT-.t93 0 0.301997f
C1895 VOUT-.t146 0 0.307141f
C1896 VOUT-.t56 0 0.301997f
C1897 VOUT-.n136 0 0.202479f
C1898 VOUT-.n137 0 0.245373f
C1899 VOUT-.t55 0 0.307141f
C1900 VOUT-.t20 0 0.301997f
C1901 VOUT-.n138 0 0.202479f
C1902 VOUT-.t124 0 0.301997f
C1903 VOUT-.t40 0 0.307141f
C1904 VOUT-.t92 0 0.301997f
C1905 VOUT-.n139 0 0.202479f
C1906 VOUT-.n140 0 0.245373f
C1907 VOUT-.t156 0 0.307141f
C1908 VOUT-.t121 0 0.301997f
C1909 VOUT-.n141 0 0.202479f
C1910 VOUT-.t87 0 0.301997f
C1911 VOUT-.t141 0 0.307141f
C1912 VOUT-.t53 0 0.301997f
C1913 VOUT-.n142 0 0.202479f
C1914 VOUT-.n143 0 0.245373f
C1915 VOUT-.t118 0 0.307141f
C1916 VOUT-.t83 0 0.301997f
C1917 VOUT-.n144 0 0.202479f
C1918 VOUT-.t50 0 0.301997f
C1919 VOUT-.t103 0 0.307141f
C1920 VOUT-.t153 0 0.301997f
C1921 VOUT-.n145 0 0.202479f
C1922 VOUT-.n146 0 0.245373f
C1923 VOUT-.t152 0 0.307141f
C1924 VOUT-.t117 0 0.301997f
C1925 VOUT-.n147 0 0.202479f
C1926 VOUT-.t81 0 0.301997f
C1927 VOUT-.t135 0 0.307141f
C1928 VOUT-.t49 0 0.301997f
C1929 VOUT-.n148 0 0.202479f
C1930 VOUT-.n149 0 0.245373f
C1931 VOUT-.t110 0 0.307141f
C1932 VOUT-.t77 0 0.301997f
C1933 VOUT-.n150 0 0.202479f
C1934 VOUT-.t42 0 0.301997f
C1935 VOUT-.t95 0 0.307141f
C1936 VOUT-.t147 0 0.301997f
C1937 VOUT-.n151 0 0.202479f
C1938 VOUT-.n152 0 0.245373f
C1939 VOUT-.t71 0 0.307141f
C1940 VOUT-.t36 0 0.301997f
C1941 VOUT-.n153 0 0.202479f
C1942 VOUT-.t144 0 0.301997f
C1943 VOUT-.t54 0 0.307141f
C1944 VOUT-.t108 0 0.301997f
C1945 VOUT-.n154 0 0.202479f
C1946 VOUT-.n155 0 0.245373f
C1947 VOUT-.t107 0 0.307141f
C1948 VOUT-.t70 0 0.301997f
C1949 VOUT-.n156 0 0.202479f
C1950 VOUT-.t35 0 0.301997f
C1951 VOUT-.n157 0 0.245373f
C1952 VOUT-.t143 0 0.301997f
C1953 VOUT-.n158 0 0.128806f
C1954 VOUT-.t91 0 0.301997f
C1955 VOUT-.n159 0 0.341177f
C1956 VOUT-.n160 0 0.27746f
C1957 VOUT-.n161 0 0.056624f
C1958 VOUT-.n162 0 0.056624f
C1959 VOUT-.n163 0 0.056624f
C1960 VOUT-.n164 0 0.166089f
C1961 VOUT-.n165 0 0.059991f
C1962 VOUT-.n166 0 0.057042f
C1963 VOUT-.n168 0 0.54737f
C1964 VOUT-.n169 0 0.056624f
C1965 VOUT-.n170 0 1.12305f
C1966 VOUT-.n172 0 0.038505f
C1967 VOUT-.n174 0 0.03624f
C1968 VOUT-.t5 0 0.052849f
C1969 VOUT-.t2 0 0.052849f
C1970 VOUT-.n175 0 0.113553f
C1971 VOUT-.n176 0 0.273093f
C1972 VOUT-.n177 0 0.03624f
C1973 VOUT-.n178 0 0.234026f
C1974 VOUT-.t18 0 0.052849f
C1975 VOUT-.t4 0 0.052849f
C1976 VOUT-.n179 0 0.113553f
C1977 VOUT-.n180 0 0.282633f
C1978 VOUT-.n181 0 0.161551f
C1979 VOUT-.t3 0 0.052849f
C1980 VOUT-.t1 0 0.052849f
C1981 VOUT-.n182 0 0.113553f
C1982 VOUT-.n183 0 0.268498f
C1983 VOUT-.n184 0 0.123221f
C1984 VOUT-.n185 0 0.03624f
C1985 VOUT-.n186 0 0.187f
C1986 VOUT-.n187 0 0.03624f
C1987 VOUT-.n188 0 0.03624f
C1988 VOUT-.n189 0 0.03624f
C1989 VOUT-.n190 0 0.03624f
C1990 VOUT-.n191 0 0.077575f
C1991 VOUT-.n192 0 0.183463f
C1992 VOUT-.t0 0 0.086201f
C1993 VOUT-.n193 0 0.33131f
C1994 VOUT-.n194 0 0.101924f
C1995 VOUT-.n196 0 1.11361f
C1996 VOUT-.n197 0 0.03624f
C1997 VOUT-.n198 0 0.056624f
C1998 w_109060_7290.n0 0 1.49009f
C1999 w_109060_7290.n1 0 0.719844f
C2000 w_109060_7290.n2 0 1.34784f
C2001 w_109060_7290.n3 0 1.33146f
C2002 w_109060_7290.n4 0 1.76138f
C2003 w_109060_7290.n5 0 0.797054f
C2004 w_109060_7290.n6 0 0.023274f
C2005 w_109060_7290.n7 0 0.687131f
C2006 w_109060_7290.n8 0 0.020024f
C2007 w_109060_7290.n9 0 0.561718f
C2008 w_109060_7290.n10 0 1.76538f
C2009 w_109060_7290.t188 0 0.058833f
C2010 w_109060_7290.t182 0 0.058833f
C2011 w_109060_7290.t190 0 0.058833f
C2012 w_109060_7290.n11 0 0.151392f
C2013 w_109060_7290.n12 0 0.516368f
C2014 w_109060_7290.t172 0 0.20705f
C2015 w_109060_7290.t38 0 0.024514f
C2016 w_109060_7290.t3 0 0.024514f
C2017 w_109060_7290.n13 0 0.085345f
C2018 w_109060_7290.n14 0 0.290209f
C2019 w_109060_7290.t148 0 0.024514f
C2020 w_109060_7290.n15 0 0.073542f
C2021 w_109060_7290.n16 0 0.034319f
C2022 w_109060_7290.n17 0 0.019611f
C2023 w_109060_7290.t177 0 0.174172f
C2024 w_109060_7290.n18 0 0.015221f
C2025 w_109060_7290.n19 0 0.019611f
C2026 w_109060_7290.n20 0 0.019611f
C2027 w_109060_7290.t176 0 0.037477f
C2028 w_109060_7290.n21 0 0.053493f
C2029 w_109060_7290.t179 0 0.029417f
C2030 w_109060_7290.t70 0 0.029417f
C2031 w_109060_7290.n22 0 0.082987f
C2032 w_109060_7290.t68 0 0.029417f
C2033 w_109060_7290.t82 0 0.029417f
C2034 w_109060_7290.n23 0 0.081706f
C2035 w_109060_7290.n24 0 0.641326f
C2036 w_109060_7290.t95 0 0.029417f
C2037 w_109060_7290.t84 0 0.029417f
C2038 w_109060_7290.n25 0 0.081706f
C2039 w_109060_7290.n26 0 0.341896f
C2040 w_109060_7290.t69 0 0.029417f
C2041 w_109060_7290.t104 0 0.029417f
C2042 w_109060_7290.n27 0 0.081706f
C2043 w_109060_7290.n28 0 0.341896f
C2044 w_109060_7290.t81 0 0.029417f
C2045 w_109060_7290.t102 0 0.029417f
C2046 w_109060_7290.n29 0 0.081706f
C2047 w_109060_7290.n30 0 0.341896f
C2048 w_109060_7290.t83 0 0.029417f
C2049 w_109060_7290.t200 0 0.029417f
C2050 w_109060_7290.n31 0 0.081706f
C2051 w_109060_7290.n32 0 1.13007f
C2052 w_109060_7290.t155 0 0.028643f
C2053 w_109060_7290.n33 0 0.2548f
C2054 w_109060_7290.t157 0 0.069966f
C2055 w_109060_7290.n34 0 0.214942f
C2056 w_109060_7290.t156 0 0.174306f
C2057 w_109060_7290.t67 0 0.129434f
C2058 w_109060_7290.t92 0 0.129434f
C2059 w_109060_7290.t85 0 0.129434f
C2060 w_109060_7290.t98 0 0.129434f
C2061 w_109060_7290.t75 0 0.129434f
C2062 w_109060_7290.t89 0 0.129434f
C2063 w_109060_7290.t103 0 0.129434f
C2064 w_109060_7290.t86 0 0.129434f
C2065 w_109060_7290.t99 0 0.129434f
C2066 w_109060_7290.t78 0 0.129434f
C2067 w_109060_7290.t165 0 0.174306f
C2068 w_109060_7290.t166 0 0.069966f
C2069 w_109060_7290.n35 0 0.214942f
C2070 w_109060_7290.t164 0 0.028643f
C2071 w_109060_7290.n36 0 0.154061f
C2072 w_109060_7290.n37 0 1.06445f
C2073 w_109060_7290.t97 0 0.058833f
C2074 w_109060_7290.t74 0 0.058833f
C2075 w_109060_7290.n38 0 0.151392f
C2076 w_109060_7290.n39 0 0.516368f
C2077 w_109060_7290.t151 0 0.20705f
C2078 w_109060_7290.t101 0 0.058833f
C2079 w_109060_7290.t80 0 0.058833f
C2080 w_109060_7290.n40 0 0.151392f
C2081 w_109060_7290.n41 0 0.516368f
C2082 w_109060_7290.t72 0 0.058833f
C2083 w_109060_7290.t88 0 0.058833f
C2084 w_109060_7290.n42 0 0.151392f
C2085 w_109060_7290.n43 0 0.516368f
C2086 w_109060_7290.t77 0 0.058833f
C2087 w_109060_7290.t94 0 0.058833f
C2088 w_109060_7290.n44 0 0.151392f
C2089 w_109060_7290.n45 0 0.516368f
C2090 w_109060_7290.t106 0 0.058833f
C2091 w_109060_7290.t91 0 0.058833f
C2092 w_109060_7290.n46 0 0.151392f
C2093 w_109060_7290.n47 0 0.608258f
C2094 w_109060_7290.t149 0 0.071381f
C2095 w_109060_7290.n48 0 0.190752f
C2096 w_109060_7290.n49 0 0.692599f
C2097 w_109060_7290.t150 0 0.448577f
C2098 w_109060_7290.t105 0 0.345157f
C2099 w_109060_7290.t90 0 0.342973f
C2100 w_109060_7290.t76 0 0.340477f
C2101 w_109060_7290.t93 0 0.345157f
C2102 w_109060_7290.t71 0 0.345157f
C2103 w_109060_7290.t87 0 0.345157f
C2104 w_109060_7290.t100 0 0.345157f
C2105 w_109060_7290.t79 0 0.345157f
C2106 w_109060_7290.t96 0 0.345157f
C2107 w_109060_7290.t73 0 0.345157f
C2108 w_109060_7290.t159 0 0.448577f
C2109 w_109060_7290.t160 0 0.20705f
C2110 w_109060_7290.n50 0 0.692599f
C2111 w_109060_7290.t158 0 0.071381f
C2112 w_109060_7290.n51 0 0.185025f
C2113 w_109060_7290.n52 0 0.252585f
C2114 w_109060_7290.n53 0 12.5228f
C2115 w_109060_7290.t130 0 0.060178f
C2116 w_109060_7290.n54 0 0.131412f
C2117 w_109060_7290.t152 0 0.060178f
C2118 w_109060_7290.t132 0 0.122079f
C2119 w_109060_7290.n55 0 0.354142f
C2120 w_109060_7290.t131 0 0.292537f
C2121 w_109060_7290.t4 0 0.229451f
C2122 w_109060_7290.t0 0 0.229451f
C2123 w_109060_7290.t111 0 0.229451f
C2124 w_109060_7290.t63 0 0.229451f
C2125 w_109060_7290.t8 0 0.229451f
C2126 w_109060_7290.t115 0 0.229451f
C2127 w_109060_7290.t21 0 0.229451f
C2128 w_109060_7290.t65 0 0.229451f
C2129 w_109060_7290.t48 0 0.229451f
C2130 w_109060_7290.t198 0 0.229451f
C2131 w_109060_7290.t153 0 0.292537f
C2132 w_109060_7290.t154 0 0.122079f
C2133 w_109060_7290.n56 0 0.354142f
C2134 w_109060_7290.n57 0 0.131412f
C2135 w_109060_7290.n58 0 2.22062f
C2136 w_109060_7290.t199 0 0.034319f
C2137 w_109060_7290.t49 0 0.034319f
C2138 w_109060_7290.n59 0 0.085768f
C2139 w_109060_7290.n60 0 0.252106f
C2140 w_109060_7290.t66 0 0.034319f
C2141 w_109060_7290.t22 0 0.034319f
C2142 w_109060_7290.n61 0 0.085768f
C2143 w_109060_7290.n62 0 0.231443f
C2144 w_109060_7290.t116 0 0.034319f
C2145 w_109060_7290.t9 0 0.034319f
C2146 w_109060_7290.n63 0 0.072296f
C2147 w_109060_7290.n64 0 0.296953f
C2148 w_109060_7290.n65 0 0.031378f
C2149 w_109060_7290.t64 0 0.034319f
C2150 w_109060_7290.t112 0 0.034319f
C2151 w_109060_7290.n66 0 0.085768f
C2152 w_109060_7290.n67 0 0.231443f
C2153 w_109060_7290.t1 0 0.034319f
C2154 w_109060_7290.t5 0 0.034319f
C2155 w_109060_7290.n68 0 0.085768f
C2156 w_109060_7290.n69 0 0.252106f
C2157 w_109060_7290.n70 0 0.125373f
C2158 w_109060_7290.n71 0 0.391366f
C2159 w_109060_7290.n72 0 12.5228f
C2160 w_109060_7290.t167 0 0.060178f
C2161 w_109060_7290.n73 0 0.131412f
C2162 w_109060_7290.t127 0 0.060178f
C2163 w_109060_7290.t169 0 0.122079f
C2164 w_109060_7290.n74 0 0.354142f
C2165 w_109060_7290.t168 0 0.292537f
C2166 w_109060_7290.t52 0 0.229451f
C2167 w_109060_7290.t50 0 0.229451f
C2168 w_109060_7290.t109 0 0.229451f
C2169 w_109060_7290.t60 0 0.229451f
C2170 w_109060_7290.t57 0 0.229451f
C2171 w_109060_7290.t113 0 0.229451f
C2172 w_109060_7290.t107 0 0.229451f
C2173 w_109060_7290.t27 0 0.229451f
C2174 w_109060_7290.t17 0 0.229451f
C2175 w_109060_7290.t13 0 0.229451f
C2176 w_109060_7290.t128 0 0.292537f
C2177 w_109060_7290.t129 0 0.122079f
C2178 w_109060_7290.n75 0 0.354142f
C2179 w_109060_7290.n76 0 0.131412f
C2180 w_109060_7290.n77 0 2.22062f
C2181 w_109060_7290.t18 0 0.034319f
C2182 w_109060_7290.t14 0 0.034319f
C2183 w_109060_7290.n78 0 0.085768f
C2184 w_109060_7290.n79 0 0.252106f
C2185 w_109060_7290.t108 0 0.034319f
C2186 w_109060_7290.t28 0 0.034319f
C2187 w_109060_7290.n80 0 0.085768f
C2188 w_109060_7290.n81 0 0.231443f
C2189 w_109060_7290.t58 0 0.034319f
C2190 w_109060_7290.t114 0 0.034319f
C2191 w_109060_7290.n82 0 0.072296f
C2192 w_109060_7290.n83 0 0.296953f
C2193 w_109060_7290.n84 0 0.031378f
C2194 w_109060_7290.t110 0 0.034319f
C2195 w_109060_7290.t61 0 0.034319f
C2196 w_109060_7290.n85 0 0.085768f
C2197 w_109060_7290.n86 0 0.231443f
C2198 w_109060_7290.t53 0 0.034319f
C2199 w_109060_7290.t51 0 0.034319f
C2200 w_109060_7290.n87 0 0.085768f
C2201 w_109060_7290.n88 0 0.252106f
C2202 w_109060_7290.n89 0 0.125373f
C2203 w_109060_7290.n90 0 0.39088f
C2204 w_109060_7290.t184 0 0.01765f
C2205 w_109060_7290.t144 0 0.01765f
C2206 w_109060_7290.n91 0 0.037951f
C2207 w_109060_7290.n92 0 0.31476f
C2208 w_109060_7290.t136 0 0.036887f
C2209 w_109060_7290.t142 0 0.036887f
C2210 w_109060_7290.n93 0 0.128394f
C2211 w_109060_7290.t145 0 0.063707f
C2212 w_109060_7290.n94 0 0.191813f
C2213 w_109060_7290.t143 0 0.170766f
C2214 w_109060_7290.t183 0 0.129434f
C2215 w_109060_7290.t137 0 0.170766f
C2216 w_109060_7290.t138 0 0.063707f
C2217 w_109060_7290.n95 0 0.191813f
C2218 w_109060_7290.n96 0 0.126062f
C2219 w_109060_7290.n97 0 0.256503f
C2220 w_109060_7290.n98 0 0.407921f
C2221 w_109060_7290.t161 0 0.060775f
C2222 w_109060_7290.t7 0 0.034319f
C2223 w_109060_7290.n99 0 0.078146f
C2224 w_109060_7290.t141 0 0.156399f
C2225 w_109060_7290.t139 0 0.060775f
C2226 w_109060_7290.n100 0 0.159108f
C2227 w_109060_7290.n101 0 0.390474f
C2228 w_109060_7290.t140 0 0.292537f
C2229 w_109060_7290.t6 0 0.229451f
C2230 w_109060_7290.t162 0 0.292537f
C2231 w_109060_7290.t163 0 0.122079f
C2232 w_109060_7290.n102 0 0.390474f
C2233 w_109060_7290.n103 0 0.156777f
C2234 w_109060_7290.n104 0 0.273144f
C2235 w_109060_7290.n105 0 0.255326f
C2236 w_109060_7290.n106 0 1.60979f
C2237 w_109060_7290.t133 0 0.037477f
C2238 w_109060_7290.n107 0 0.019611f
C2239 w_109060_7290.n108 0 0.034319f
C2240 w_109060_7290.n110 0 0.034319f
C2241 w_109060_7290.n111 0 0.019611f
C2242 w_109060_7290.n112 0 0.019611f
C2243 w_109060_7290.n113 0 0.034319f
C2244 w_109060_7290.n114 0 0.019611f
C2245 w_109060_7290.t196 0 0.156399f
C2246 w_109060_7290.t15 0 0.156399f
C2247 w_109060_7290.t11 0 0.156399f
C2248 w_109060_7290.t36 0 0.156399f
C2249 w_109060_7290.t134 0 0.174172f
C2250 w_109060_7290.n116 0 0.209717f
C2251 w_109060_7290.n117 0 0.015879f
C2252 w_109060_7290.n118 0 0.034619f
C2253 w_109060_7290.t135 0 0.024514f
C2254 w_109060_7290.n119 0 0.073542f
C2255 w_109060_7290.n120 0 0.038589f
C2256 w_109060_7290.n121 0 0.054475f
C2257 w_109060_7290.n122 0 0.686601f
C2258 w_109060_7290.t12 0 0.024514f
C2259 w_109060_7290.t16 0 0.024514f
C2260 w_109060_7290.n123 0 0.085345f
C2261 w_109060_7290.n124 0 0.290209f
C2262 w_109060_7290.n125 0 0.184712f
C2263 w_109060_7290.n126 0 0.184712f
C2264 w_109060_7290.t124 0 0.037477f
C2265 w_109060_7290.n127 0 0.053493f
C2266 w_109060_7290.n128 0 0.028148f
C2267 w_109060_7290.t178 0 0.024514f
C2268 w_109060_7290.n130 0 0.053931f
C2269 w_109060_7290.n132 0 0.019611f
C2270 w_109060_7290.n133 0 0.053931f
C2271 w_109060_7290.n134 0 0.053931f
C2272 w_109060_7290.t126 0 0.024514f
C2273 w_109060_7290.n136 0 0.073542f
C2274 w_109060_7290.n137 0 0.052928f
C2275 w_109060_7290.n139 0 0.073542f
C2276 w_109060_7290.n140 0 0.042142f
C2277 w_109060_7290.n141 0 0.015221f
C2278 w_109060_7290.n142 0 0.191944f
C2279 w_109060_7290.t125 0 0.174172f
C2280 w_109060_7290.t191 0 0.156399f
C2281 w_109060_7290.t37 0 0.156399f
C2282 w_109060_7290.t2 0 0.156399f
C2283 w_109060_7290.t32 0 0.156399f
C2284 w_109060_7290.t147 0 0.174172f
C2285 w_109060_7290.n143 0 0.015879f
C2286 w_109060_7290.n144 0 0.019611f
C2287 w_109060_7290.n146 0 0.034619f
C2288 w_109060_7290.n147 0 0.034319f
C2289 w_109060_7290.n148 0 0.034319f
C2290 w_109060_7290.n149 0 0.019611f
C2291 w_109060_7290.n150 0 0.209717f
C2292 w_109060_7290.n151 0 0.015221f
C2293 w_109060_7290.n152 0 0.04298f
C2294 w_109060_7290.t146 0 0.037477f
C2295 w_109060_7290.n153 0 0.054472f
C2296 w_109060_7290.n154 0 0.664205f
C2297 w_109060_7290.t46 0 0.029417f
C2298 w_109060_7290.t23 0 0.029417f
C2299 w_109060_7290.n155 0 0.08321f
C2300 w_109060_7290.t30 0 0.029417f
C2301 w_109060_7290.t186 0 0.029417f
C2302 w_109060_7290.n156 0 0.081924f
C2303 w_109060_7290.n157 0 0.643826f
C2304 w_109060_7290.t35 0 0.029417f
C2305 w_109060_7290.t54 0 0.029417f
C2306 w_109060_7290.n158 0 0.081924f
C2307 w_109060_7290.n159 0 0.343148f
C2308 w_109060_7290.t26 0 0.029417f
C2309 w_109060_7290.t29 0 0.029417f
C2310 w_109060_7290.n160 0 0.081924f
C2311 w_109060_7290.n161 0 0.343148f
C2312 w_109060_7290.t180 0 0.029417f
C2313 w_109060_7290.t43 0 0.029417f
C2314 w_109060_7290.n162 0 0.081924f
C2315 w_109060_7290.n163 0 0.343148f
C2316 w_109060_7290.t117 0 0.029417f
C2317 w_109060_7290.t10 0 0.029417f
C2318 w_109060_7290.n164 0 0.081924f
C2319 w_109060_7290.n165 0 1.13534f
C2320 w_109060_7290.t121 0 0.028643f
C2321 w_109060_7290.n166 0 0.2548f
C2322 w_109060_7290.t123 0 0.069966f
C2323 w_109060_7290.n167 0 0.214942f
C2324 w_109060_7290.t122 0 0.174306f
C2325 w_109060_7290.t20 0 0.129434f
C2326 w_109060_7290.t39 0 0.129434f
C2327 w_109060_7290.t197 0 0.129434f
C2328 w_109060_7290.t185 0 0.129434f
C2329 w_109060_7290.t47 0 0.129434f
C2330 w_109060_7290.t59 0 0.129434f
C2331 w_109060_7290.t31 0 0.129434f
C2332 w_109060_7290.t19 0 0.129434f
C2333 w_109060_7290.t62 0 0.129434f
C2334 w_109060_7290.t40 0 0.129434f
C2335 w_109060_7290.t119 0 0.174306f
C2336 w_109060_7290.t120 0 0.069966f
C2337 w_109060_7290.n168 0 0.214942f
C2338 w_109060_7290.t118 0 0.028643f
C2339 w_109060_7290.n169 0 0.154061f
C2340 w_109060_7290.n170 0 1.06483f
C2341 w_109060_7290.n171 0 0.185727f
C2342 w_109060_7290.n172 0 0.224109f
C2343 w_109060_7290.t170 0 0.071381f
C2344 w_109060_7290.n173 0 0.185025f
C2345 w_109060_7290.n174 0 0.692599f
C2346 w_109060_7290.t171 0 0.448577f
C2347 w_109060_7290.t181 0 0.345157f
C2348 w_109060_7290.t189 0 0.345157f
C2349 w_109060_7290.t24 0 0.345157f
C2350 w_109060_7290.t187 0 0.345157f
C2351 w_109060_7290.t194 0 0.345157f
C2352 w_109060_7290.t55 0 0.345157f
C2353 w_109060_7290.t192 0 0.345157f
C2354 w_109060_7290.t44 0 0.345157f
C2355 w_109060_7290.t41 0 0.345157f
C2356 w_109060_7290.t33 0 0.345157f
C2357 w_109060_7290.t174 0 0.448577f
C2358 w_109060_7290.t175 0 0.20705f
C2359 w_109060_7290.n175 0 0.692599f
C2360 w_109060_7290.t173 0 0.071381f
C2361 w_109060_7290.n176 0 0.190752f
C2362 w_109060_7290.t42 0 0.058833f
C2363 w_109060_7290.t34 0 0.058833f
C2364 w_109060_7290.n177 0 0.151392f
C2365 w_109060_7290.n178 0 0.608258f
C2366 w_109060_7290.t193 0 0.058833f
C2367 w_109060_7290.t45 0 0.058833f
C2368 w_109060_7290.n179 0 0.151392f
C2369 w_109060_7290.n180 0 0.516368f
C2370 w_109060_7290.t195 0 0.058833f
C2371 w_109060_7290.t56 0 0.058833f
C2372 w_109060_7290.n181 0 0.151392f
C2373 w_109060_7290.n182 0 0.516368f
C2374 w_109060_7290.n183 0 0.516361f
C2375 w_109060_7290.n184 0 0.151399f
C2376 w_109060_7290.t25 0 0.058833f
C2377 X.n0 0 0.069924f
C2378 X.n1 0 0.102555f
C2379 X.n2 0 0.239296f
C2380 X.n3 0 0.162703f
C2381 X.n4 0 0.273038f
C2382 X.t24 0 0.023308f
C2383 X.t12 0 0.023308f
C2384 X.n5 0 0.050716f
C2385 X.n6 0 0.162065f
C2386 X.n7 0 0.046616f
C2387 X.n8 0 0.089133f
C2388 X.t18 0 0.023308f
C2389 X.t23 0 0.023308f
C2390 X.n9 0 0.050716f
C2391 X.n10 0 0.162065f
C2392 X.n11 0 0.166674f
C2393 X.n12 0 0.102555f
C2394 X.n13 0 0.102555f
C2395 X.n14 0 0.074586f
C2396 X.t28 0 0.050112f
C2397 X.t44 0 0.056969f
C2398 X.n17 0 0.04646f
C2399 X.t40 0 0.050112f
C2400 X.t26 0 0.050112f
C2401 X.t37 0 0.050112f
C2402 X.t46 0 0.050112f
C2403 X.t29 0 0.050112f
C2404 X.t41 0 0.050112f
C2405 X.t35 0 0.050112f
C2406 X.t53 0 0.056969f
C2407 X.n18 0 0.051413f
C2408 X.n19 0 0.031466f
C2409 X.n20 0 0.031466f
C2410 X.n21 0 0.031466f
C2411 X.n22 0 0.031466f
C2412 X.n23 0 0.031466f
C2413 X.n24 0 0.026513f
C2414 X.n25 0 0.012874f
C2415 X.t31 0 0.032631f
C2416 X.t48 0 0.039624f
C2417 X.n26 0 0.034671f
C2418 X.t43 0 0.032631f
C2419 X.t27 0 0.032631f
C2420 X.t39 0 0.032631f
C2421 X.t50 0 0.032631f
C2422 X.t32 0 0.032631f
C2423 X.t45 0 0.032631f
C2424 X.t36 0 0.032631f
C2425 X.t54 0 0.039624f
C2426 X.n27 0 0.039624f
C2427 X.n28 0 0.025639f
C2428 X.n29 0 0.025639f
C2429 X.n30 0 0.025639f
C2430 X.n31 0 0.025639f
C2431 X.n32 0 0.025639f
C2432 X.n33 0 0.020686f
C2433 X.n34 0 0.012874f
C2434 X.n35 0 0.080307f
C2435 X.n37 0 0.074586f
C2436 X.t1 0 0.644946f
C2437 X.n38 0 0.074586f
C2438 X.n39 0 0.074586f
C2439 X.n40 0 0.073885f
C2440 X.n41 0 0.692003f
C2441 X.n43 0 0.647964f
C2442 X.n44 0 0.024697f
C2443 X.n45 0 0.024862f
C2444 X.n46 0 0.024862f
C2445 X.t42 0 0.102555f
C2446 X.t30 0 0.102555f
C2447 X.t47 0 0.102555f
C2448 X.t33 0 0.102555f
C2449 X.t51 0 0.109229f
C2450 X.n47 0 0.086559f
C2451 X.n48 0 0.048947f
C2452 X.n49 0 0.048947f
C2453 X.n50 0 0.043994f
C2454 X.t52 0 0.102555f
C2455 X.t34 0 0.102555f
C2456 X.t49 0 0.102555f
C2457 X.t38 0 0.102555f
C2458 X.t25 0 0.109229f
C2459 X.n51 0 0.086559f
C2460 X.n52 0 0.048947f
C2461 X.n53 0 0.048947f
C2462 X.n54 0 0.043994f
C2463 X.n55 0 0.010564f
C2464 X.n56 0 0.025027f
C2465 X.n57 0 0.058911f
C2466 X.n58 0 0.0336f
C2467 X.n59 0 0.038132f
C2468 X.n60 0 1.03022f
C2469 X.n61 0 0.074586f
C2470 X.n63 0 0.074586f
C2471 X.n64 0 0.074586f
C2472 X.n65 0 0.100673f
C2473 X.n66 0 0.121202f
C2474 X.n67 0 0.074586f
C2475 X.n68 0 0.096125f
C2476 X.n69 0 0.074586f
C2477 X.n70 0 0.074586f
C2478 X.n71 0 0.096125f
C2479 X.n72 0 0.074586f
C2480 X.n73 0 0.122901f
C2481 X.t10 0 0.054385f
C2482 X.t8 0 0.054385f
C2483 X.n74 0 0.111251f
C2484 X.n75 0 0.297688f
C2485 X.t14 0 0.054385f
C2486 X.t17 0 0.054385f
C2487 X.n76 0 0.111251f
C2488 X.n77 0 0.302606f
C2489 X.t22 0 0.054385f
C2490 X.t13 0 0.054385f
C2491 X.n78 0 0.111251f
C2492 X.n79 0 0.302606f
C2493 X.n80 0 0.100632f
C2494 X.t2 0 0.054385f
C2495 X.t0 0 0.054385f
C2496 X.n81 0 0.111251f
C2497 X.n82 0 0.297688f
C2498 X.n83 0 0.058991f
C2499 X.t9 0 0.054385f
C2500 X.t15 0 0.054385f
C2501 X.n84 0 0.111251f
C2502 X.n85 0 0.297688f
C2503 X.n86 0 0.058991f
C2504 X.n87 0 0.100632f
C2505 X.t6 0 0.054385f
C2506 X.t21 0 0.054385f
C2507 X.n88 0 0.111251f
C2508 X.n89 0 0.297688f
C2509 X.n90 0 0.096125f
C2510 X.n91 0 0.082469f
C2511 X.n92 0 0.049724f
C2512 X.n93 0 0.049724f
C2513 X.n94 0 0.082469f
C2514 X.n95 0 0.096125f
C2515 X.n96 0 0.170057f
C2516 X.n97 0 0.251893f
C2517 X.n98 0 0.320326f
C2518 X.n99 0 0.074586f
C2519 X.n100 0 0.074586f
C2520 X.n101 0 0.121202f
C2521 X.n102 0 0.074586f
C2522 X.n103 0 0.074586f
C2523 X.n104 0 0.074586f
C2524 X.n105 0 0.074586f
C2525 X.n106 0 0.121202f
C2526 X.n107 0 0.074586f
C2527 X.n108 0 0.074586f
C2528 X.n109 0 0.074586f
C2529 X.n110 0 0.074586f
C2530 X.n111 0 0.074586f
C2531 X.n112 0 0.074586f
C2532 X.n113 0 0.074586f
C2533 X.n114 0 0.121202f
C2534 X.n115 0 0.582701f
C2535 X.n116 0 0.582701f
C2536 X.n117 0 0.073885f
C2537 X.n118 0 0.074586f
C2538 X.n119 0 0.074586f
C2539 X.n121 0 0.913675f
C2540 X.n122 0 0.913675f
C2541 X.n124 0 0.456838f
C2542 X.n125 0 2.20416f
C2543 X.n126 0 0.601348f
C2544 X.n127 0 0.225311f
C2545 X.n128 0 0.615332f
C2546 X.n129 0 0.102555f
C2547 X.n130 0 0.102555f
C2548 X.n131 0 0.102555f
C2549 X.n132 0 0.239296f
C2550 X.t16 0 0.023308f
C2551 X.t4 0 0.023308f
C2552 X.n133 0 0.050716f
C2553 X.n134 0 0.157946f
C2554 X.n135 0 0.162703f
C2555 X.n136 0 0.078384f
C2556 X.n137 0 0.046616f
C2557 X.n138 0 0.162703f
C2558 X.t19 0 0.023308f
C2559 X.t20 0 0.023308f
C2560 X.n139 0 0.050716f
C2561 X.n140 0 0.157946f
C2562 X.n141 0 0.052064f
C2563 X.t7 0 0.023308f
C2564 X.t3 0 0.023308f
C2565 X.n142 0 0.050716f
C2566 X.n143 0 0.157946f
C2567 X.n144 0 0.052064f
C2568 X.n145 0 0.089133f
C2569 X.t11 0 0.023308f
C2570 X.t5 0 0.023308f
C2571 X.n146 0 0.050716f
C2572 X.n147 0 0.157946f
C2573 X.n148 0 0.162703f
C2574 X.n149 0 0.078384f
C2575 X.n150 0 0.177677f
C2576 X.n151 0 0.327848f
C2577 X.n152 0 0.351511f
C2578 X.n153 0 0.102555f
C2579 X.n154 0 0.239296f
C2580 X.n155 0 0.102555f
C2581 X.n156 0 0.083909f
.ends

