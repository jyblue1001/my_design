* PEX produced on Mon Feb  3 03:52:54 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from TSPC_FF_ratioed_divide24_magic.ext - technology: sky130A

.subckt TSPC_FF_ratioed_divide24_magic VOUT VIN VDDA GNDA
X0 VDDA.t45 div2.t2 div2_3_1.A.t1 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1 div2_3_0.C.t3 div2_3_0.CLK.t3 GNDA.t63 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 div2.t1 div2_3_1.C.t4 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X3 div2_3_0.A.t1 div2_3_0.CLK.t4 div2_3_0.B.t1 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 GNDA.t60 div2_3_0.CLK.t5 div2_3_0.C.t2 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X5 VDDA.t43 div2.t3 div2_3_2.CLK.t1 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 GNDA.t14 div3_2_0.I.t2 div3_2_0.G.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X7 VDDA.t9 div3_2_0.I.t3 VOUT.t1 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 div2_3_0.CLK.t2 div4.t2 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 div2_3_0.B.t0 div8.t2 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X10 div3_2_0.G.t1 div3_2_0.D.t2 div3_2_0.F.t0 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VDDA.t25 div3_2_0.E.t3 div3_2_0.H.t1 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 GNDA.t36 div2_3_1.CLK.t3 div2_3_1.C.t1 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X13 GNDA.t31 div4.t3 div2_3_0.CLK.t1 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 div3_2_0.D.t1 div3_2_0.C.t4 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 VOUT.t2 div3_2_0.I.t4 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X16 div3_2_0.F.t1 div3_2_0.CLK.t3 div3_2_0.E.t2 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 div2_3_1.C.t0 div2_3_1.CLK.t4 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X18 VDDA.t33 div8.t3 div2_3_0.A.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X19 GNDA.t16 div3_2_0.CLK.t4 div3_2_0.C.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X20 VDDA.t23 div8.t4 div3_2_0.CLK.t1 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X21 div2_3_2.C.t0 div2_3_2.A.t2 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X22 div3_2_0.C.t3 div3_2_0.A.t2 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 GNDA.t46 div2_3_1.CLK.t5 div2_3_1.C.t2 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X24 VDDA.t39 VIN.t0 div2_3_1.CLK.t2 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X25 div2_3_1.C.t3 div2_3_1.A.t2 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X26 GNDA.t9 div2_3_2.CLK.t3 div2_3_2.C.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 div3_2_0.C.t0 div3_2_0.CLK.t5 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X28 div3_2_0.D.t0 div3_2_0.CLK.t6 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X29 VDDA.t1 div3_2_0.D.t3 div3_2_0.E.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X30 div4.t0 div2_3_2.C.t4 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X31 div4.t1 div2_3_2.CLK.t4 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X32 GNDA.t28 div2_3_2.CLK.t5 div2_3_2.C.t2 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X33 GNDA.t26 div3_2_0.CLK.t7 div3_2_0.C.t2 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X34 div3_2_0.CLK.t0 div8.t5 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X35 div2_3_1.A.t0 div2_3_1.CLK.t6 div2_3_1.B.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X36 div2_3_2.C.t1 div2_3_2.CLK.t6 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X37 div2_3_2.A.t0 div2_3_2.CLK.t7 div2_3_2.B.t0 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X38 GNDA.t22 div8.t6 div3_2_0.CLK.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X39 VDDA.t49 VOUT.t3 div3_2_0.A.t1 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X40 div2_3_1.B.t1 div2.t4 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X41 GNDA.t34 div3_2_0.CLK.t8 div3_2_0.H.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X42 VOUT.t0 div3_2_0.I.t5 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X43 VDDA.t13 div4.t4 div2_3_0.CLK.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X44 div2_3_2.B.t1 div4.t5 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X45 div3_2_0.A.t0 div3_2_0.CLK.t9 div3_2_0.B.t0 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 div2.t0 div2_3_1.CLK.t7 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X47 div2_3_0.C.t0 div2_3_0.A.t2 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X48 GNDA.t52 VIN.t1 div2_3_1.CLK.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X49 div3_2_0.H.t0 div3_2_0.CLK.t10 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 div2_3_2.CLK.t0 div2.t5 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X51 div8.t1 div2_3_0.CLK.t6 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X52 GNDA.t54 div2.t6 div2_3_2.CLK.t2 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X53 div8.t0 div2_3_0.C.t4 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X54 div3_2_0.B.t1 VOUT.t4 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X55 div2_3_1.CLK.t0 VIN.t2 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X56 div3_2_0.I.t1 div3_2_0.H.t4 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X57 GNDA.t48 div3_2_0.CLK.t11 div3_2_0.H.t3 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X58 div3_2_0.E.t0 div3_2_0.I.t6 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X59 GNDA.t58 div2_3_0.CLK.t7 div2_3_0.C.t1 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X60 VDDA.t15 div4.t6 div2_3_2.A.t1 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X61 div3_2_0.I.t0 div3_2_0.CLK.t12 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
R0 div2.t2 div2.t4 819.4
R1 div2.n0 div2.t0 663.801
R2 div2.n0 div2.t2 489.168
R3 div2.t3 div2.t5 401.668
R4 div2.n1 div2.t1 270.12
R5 div2.n2 div2.t3 257.067
R6 div2_3_2.VIN div2.n2 216.9
R7 div2.n2 div2.t6 208.868
R8 div2.n3 div2_3_2.VIN 192.167
R9 div2.n1 div2.n0 67.2005
R10 div2.n3 div2.n1 25.6005
R11 div2_3_1.VOUT div2.n3 4.8005
R12 div2_3_1.A.n0 div2_3_1.A.t1 713.933
R13 div2_3_1.A.n0 div2_3_1.A.t2 314.233
R14 div2_3_1.A.t0 div2_3_1.A.n0 308.2
R15 VDDA.t4 VDDA.t0 2307.14
R16 VDDA.t2 VDDA.t18 2126.19
R17 VDDA.t16 VDDA.t22 2080.95
R18 VDDA.t12 VDDA.t6 2080.95
R19 VDDA.t30 VDDA.t42 2080.95
R20 VDDA.t10 VDDA.t24 1492.86
R21 VDDA.t50 VDDA.t48 1130.95
R22 VDDA.t32 VDDA.t26 1130.95
R23 VDDA.t40 VDDA.t14 1130.95
R24 VDDA.t44 VDDA.t36 1130.95
R25 VDDA.t28 VDDA.n18 927.381
R26 VDDA.n19 VDDA.t20 927.381
R27 VDDA.t34 VDDA.n33 927.381
R28 VDDA.n34 VDDA.t46 927.381
R29 VDDA.n6 VDDA.t9 673.375
R30 VDDA.n6 VDDA.t19 673.101
R31 VDDA.n1 VDDA.t31 663.801
R32 VDDA.n2 VDDA.t7 663.801
R33 VDDA.n4 VDDA.t17 663.801
R34 VDDA.n5 VDDA.t5 663.801
R35 VDDA.n18 VDDA.t4 610.715
R36 VDDA.n19 VDDA.t16 610.715
R37 VDDA.n33 VDDA.t6 610.715
R38 VDDA.n34 VDDA.t30 610.715
R39 VDDA.n40 VDDA.n39 594.301
R40 VDDA.n38 VDDA.n37 594.301
R41 VDDA.n28 VDDA.n27 594.301
R42 VDDA.n30 VDDA.n29 594.301
R43 VDDA.n25 VDDA.n24 594.301
R44 VDDA.n23 VDDA.n22 594.301
R45 VDDA.n13 VDDA.n12 594.301
R46 VDDA.n15 VDDA.n14 594.301
R47 VDDA.n10 VDDA.n9 594.301
R48 VDDA.n8 VDDA.n7 594.301
R49 VDDA.t18 VDDA.t8 497.62
R50 VDDA.t24 VDDA.t2 497.62
R51 VDDA.t0 VDDA.t10 497.62
R52 VDDA.t48 VDDA.t28 497.62
R53 VDDA.t22 VDDA.t50 497.62
R54 VDDA.t20 VDDA.t32 497.62
R55 VDDA.t26 VDDA.t12 497.62
R56 VDDA.t14 VDDA.t34 497.62
R57 VDDA.t42 VDDA.t40 497.62
R58 VDDA.t46 VDDA.t44 497.62
R59 VDDA.t36 VDDA.t38 497.62
R60 VDDA.n20 VDDA.n19 370
R61 VDDA.n33 VDDA.n32 370
R62 VDDA.n35 VDDA.n34 370
R63 VDDA.n18 VDDA.n17 370
R64 VDDA.n39 VDDA.t37 78.8005
R65 VDDA.n39 VDDA.t39 78.8005
R66 VDDA.n37 VDDA.t47 78.8005
R67 VDDA.n37 VDDA.t45 78.8005
R68 VDDA.n27 VDDA.t41 78.8005
R69 VDDA.n27 VDDA.t43 78.8005
R70 VDDA.n29 VDDA.t35 78.8005
R71 VDDA.n29 VDDA.t15 78.8005
R72 VDDA.n24 VDDA.t27 78.8005
R73 VDDA.n24 VDDA.t13 78.8005
R74 VDDA.n22 VDDA.t21 78.8005
R75 VDDA.n22 VDDA.t33 78.8005
R76 VDDA.n12 VDDA.t51 78.8005
R77 VDDA.n12 VDDA.t23 78.8005
R78 VDDA.n14 VDDA.t29 78.8005
R79 VDDA.n14 VDDA.t49 78.8005
R80 VDDA.n9 VDDA.t11 78.8005
R81 VDDA.n9 VDDA.t1 78.8005
R82 VDDA.n7 VDDA.t3 78.8005
R83 VDDA.n7 VDDA.t25 78.8005
R84 VDDA.n35 VDDA.n1 12.8005
R85 VDDA.n32 VDDA.n2 12.8005
R86 VDDA.n20 VDDA.n4 12.8005
R87 VDDA.n17 VDDA.n5 12.8005
R88 VDDA.n11 VDDA.n5 9.3005
R89 VDDA.n17 VDDA.n16 9.3005
R90 VDDA.n4 VDDA.n3 9.3005
R91 VDDA.n21 VDDA.n20 9.3005
R92 VDDA.n26 VDDA.n2 9.3005
R93 VDDA.n32 VDDA.n31 9.3005
R94 VDDA.n1 VDDA.n0 9.3005
R95 VDDA.n36 VDDA.n35 9.3005
R96 VDDA.n11 VDDA.n10 0.7755
R97 VDDA.n8 VDDA.n6 0.588
R98 VDDA.n10 VDDA.n8 0.5505
R99 VDDA VDDA.n3 0.4755
R100 VDDA.n26 VDDA 0.4755
R101 VDDA VDDA.n0 0.4755
R102 VDDA.n15 VDDA.n13 0.4505
R103 VDDA.n25 VDDA.n23 0.4505
R104 VDDA.n30 VDDA.n28 0.4505
R105 VDDA.n40 VDDA.n38 0.4505
R106 VDDA.n16 VDDA.n15 0.3255
R107 VDDA.n23 VDDA.n21 0.3255
R108 VDDA.n31 VDDA.n30 0.3255
R109 VDDA.n38 VDDA.n36 0.3255
R110 VDDA.n13 VDDA 0.238
R111 VDDA VDDA.n25 0.238
R112 VDDA.n28 VDDA 0.238
R113 VDDA VDDA.n40 0.238
R114 VDDA.n16 VDDA.n11 0.1005
R115 VDDA.n21 VDDA.n3 0.1005
R116 VDDA.n31 VDDA.n26 0.1005
R117 VDDA.n36 VDDA.n0 0.1005
R118 div2_3_0.CLK.n5 div2_3_0.CLK.t0 723.534
R119 div2_3_0.CLK.n4 div2_3_0.CLK.t2 723.534
R120 div2_3_0.CLK.n0 div2_3_0.CLK.t6 369.534
R121 div2_3_0.CLK.n3 div2_3_0.CLK.n2 366.856
R122 div2_3_0.CLK.t1 div2_3_0.CLK.n5 254.333
R123 div2_3_0.CLK.n3 div2_3_0.CLK.t4 190.123
R124 div2_3_0.CLK.n4 div2_3_0.CLK.n3 187.201
R125 div2_3_0.CLK.n1 div2_3_0.CLK.n0 176.733
R126 div2_3_0.CLK.n2 div2_3_0.CLK.n1 176.733
R127 div2_3_0.CLK.n0 div2_3_0.CLK.t7 112.468
R128 div2_3_0.CLK.n2 div2_3_0.CLK.t5 112.468
R129 div2_3_0.CLK.n1 div2_3_0.CLK.t3 112.468
R130 div2_3_0.CLK.n5 div2_3_0.CLK.n4 70.4005
R131 GNDA.t51 GNDA.t19 719016
R132 GNDA.t23 GNDA.t38 3723.08
R133 GNDA.t37 GNDA.t25 3723.08
R134 GNDA.t59 GNDA.t61 3723.08
R135 GNDA.t8 GNDA.t29 3723.08
R136 GNDA.t45 GNDA.t10 3723.08
R137 GNDA.t19 GNDA.t17 2820.51
R138 GNDA.t47 GNDA.n30 2200
R139 GNDA.n19 GNDA.t21 2200
R140 GNDA.n19 GNDA.t64 2200
R141 GNDA.t30 GNDA.n18 2200
R142 GNDA.n18 GNDA.t11 2200
R143 GNDA.n31 GNDA.t53 2200
R144 GNDA.n31 GNDA.t41 2200
R145 GNDA.n30 GNDA.t13 1523.08
R146 GNDA.t17 GNDA.t33 1241.03
R147 GNDA.t33 GNDA.t4 1241.03
R148 GNDA.t4 GNDA.t47 1241.03
R149 GNDA.t32 GNDA.t13 1241.03
R150 GNDA.t38 GNDA.t32 1241.03
R151 GNDA.t15 GNDA.t23 1241.03
R152 GNDA.t6 GNDA.t15 1241.03
R153 GNDA.t25 GNDA.t6 1241.03
R154 GNDA.t49 GNDA.t37 1241.03
R155 GNDA.t21 GNDA.t49 1241.03
R156 GNDA.t64 GNDA.t57 1241.03
R157 GNDA.t57 GNDA.t62 1241.03
R158 GNDA.t62 GNDA.t59 1241.03
R159 GNDA.t61 GNDA.t0 1241.03
R160 GNDA.t0 GNDA.t30 1241.03
R161 GNDA.t11 GNDA.t27 1241.03
R162 GNDA.t27 GNDA.t39 1241.03
R163 GNDA.t39 GNDA.t8 1241.03
R164 GNDA.t29 GNDA.t43 1241.03
R165 GNDA.t43 GNDA.t53 1241.03
R166 GNDA.t41 GNDA.t35 1241.03
R167 GNDA.t35 GNDA.t2 1241.03
R168 GNDA.t2 GNDA.t45 1241.03
R169 GNDA.t10 GNDA.t55 1241.03
R170 GNDA.t55 GNDA.t51 1241.03
R171 GNDA.n20 GNDA.n19 1179.3
R172 GNDA.n18 GNDA.n17 1179.3
R173 GNDA.n32 GNDA.n31 1179.3
R174 GNDA.n30 GNDA.n29 1170
R175 GNDA.n2 GNDA.t20 242.613
R176 GNDA.n0 GNDA.t14 233
R177 GNDA.n38 GNDA.n37 194.3
R178 GNDA.n36 GNDA.n35 194.3
R179 GNDA.n34 GNDA.n33 194.3
R180 GNDA.n12 GNDA.n11 194.3
R181 GNDA.n14 GNDA.n13 194.3
R182 GNDA.n16 GNDA.n15 194.3
R183 GNDA.n10 GNDA.n9 194.3
R184 GNDA.n8 GNDA.n7 194.3
R185 GNDA.n6 GNDA.n5 194.3
R186 GNDA.n22 GNDA.n21 194.3
R187 GNDA.n24 GNDA.n23 194.3
R188 GNDA.n26 GNDA.n25 194.3
R189 GNDA.n4 GNDA.n3 194.3
R190 GNDA.n2 GNDA.n1 194.3
R191 GNDA.n37 GNDA.t56 48.0005
R192 GNDA.n37 GNDA.t52 48.0005
R193 GNDA.n35 GNDA.t3 48.0005
R194 GNDA.n35 GNDA.t46 48.0005
R195 GNDA.n33 GNDA.t42 48.0005
R196 GNDA.n33 GNDA.t36 48.0005
R197 GNDA.n11 GNDA.t44 48.0005
R198 GNDA.n11 GNDA.t54 48.0005
R199 GNDA.n13 GNDA.t40 48.0005
R200 GNDA.n13 GNDA.t9 48.0005
R201 GNDA.n15 GNDA.t12 48.0005
R202 GNDA.n15 GNDA.t28 48.0005
R203 GNDA.n9 GNDA.t1 48.0005
R204 GNDA.n9 GNDA.t31 48.0005
R205 GNDA.n7 GNDA.t63 48.0005
R206 GNDA.n7 GNDA.t60 48.0005
R207 GNDA.n5 GNDA.t65 48.0005
R208 GNDA.n5 GNDA.t58 48.0005
R209 GNDA.n21 GNDA.t50 48.0005
R210 GNDA.n21 GNDA.t22 48.0005
R211 GNDA.n23 GNDA.t7 48.0005
R212 GNDA.n23 GNDA.t26 48.0005
R213 GNDA.n25 GNDA.t24 48.0005
R214 GNDA.n25 GNDA.t16 48.0005
R215 GNDA.n3 GNDA.t5 48.0005
R216 GNDA.n3 GNDA.t48 48.0005
R217 GNDA.n1 GNDA.t18 48.0005
R218 GNDA.n1 GNDA.t34 48.0005
R219 GNDA.n29 GNDA.n0 12.8005
R220 GNDA.n29 GNDA.n28 9.3005
R221 GNDA.n27 GNDA.n0 9.3005
R222 GNDA.n27 GNDA.n26 0.8255
R223 GNDA.n24 GNDA.n22 0.688
R224 GNDA.n10 GNDA.n8 0.688
R225 GNDA.n14 GNDA.n12 0.688
R226 GNDA.n38 GNDA.n36 0.688
R227 GNDA.n28 GNDA.n4 0.313
R228 GNDA.n20 GNDA.n6 0.313
R229 GNDA.n17 GNDA.n16 0.313
R230 GNDA.n34 GNDA.n32 0.313
R231 GNDA.n4 GNDA.n2 0.2755
R232 GNDA.n26 GNDA.n24 0.2755
R233 GNDA.n8 GNDA.n6 0.2755
R234 GNDA.n16 GNDA.n14 0.2755
R235 GNDA.n36 GNDA.n34 0.2755
R236 GNDA.n22 GNDA 0.238
R237 GNDA GNDA.n10 0.238
R238 GNDA.n12 GNDA 0.238
R239 GNDA GNDA.n38 0.238
R240 GNDA.n28 GNDA.n27 0.1005
R241 GNDA GNDA.n20 0.0755
R242 GNDA.n17 GNDA 0.0755
R243 GNDA.n32 GNDA 0.0755
R244 div2_3_0.C.n0 div2_3_0.C.t0 721.4
R245 div2_3_0.C.n1 div2_3_0.C.t4 349.433
R246 div2_3_0.C.n0 div2_3_0.C.t2 276.733
R247 div2_3_0.C.n2 div2_3_0.C.n1 206.333
R248 div2_3_0.C.n1 div2_3_0.C.n0 48.0005
R249 div2_3_0.C.n2 div2_3_0.C.t1 48.0005
R250 div2_3_0.C.t3 div2_3_0.C.n2 48.0005
R251 div2_3_1.C.n0 div2_3_1.C.t3 721.4
R252 div2_3_1.C.n1 div2_3_1.C.t4 349.433
R253 div2_3_1.C.n0 div2_3_1.C.t2 276.733
R254 div2_3_1.C.n2 div2_3_1.C.n1 206.333
R255 div2_3_1.C.n1 div2_3_1.C.n0 48.0005
R256 div2_3_1.C.n2 div2_3_1.C.t1 48.0005
R257 div2_3_1.C.t0 div2_3_1.C.n2 48.0005
R258 div2_3_0.B.t0 div2_3_0.B.t1 96.0005
R259 div2_3_0.A.n0 div2_3_0.A.t0 713.933
R260 div2_3_0.A.n0 div2_3_0.A.t2 314.233
R261 div2_3_0.A.t1 div2_3_0.A.n0 308.2
R262 div2_3_2.CLK.n4 div2_3_2.CLK.t0 723.534
R263 div2_3_2.CLK.t1 div2_3_2.CLK.n5 723.534
R264 div2_3_2.CLK.n0 div2_3_2.CLK.t4 369.534
R265 div2_3_2.CLK.n3 div2_3_2.CLK.n2 366.856
R266 div2_3_2.CLK.n5 div2_3_2.CLK.t2 254.333
R267 div2_3_2.CLK.n3 div2_3_2.CLK.t7 190.123
R268 div2_3_2.CLK.n4 div2_3_2.CLK.n3 187.201
R269 div2_3_2.CLK.n1 div2_3_2.CLK.n0 176.733
R270 div2_3_2.CLK.n2 div2_3_2.CLK.n1 176.733
R271 div2_3_2.CLK.n0 div2_3_2.CLK.t5 112.468
R272 div2_3_2.CLK.n2 div2_3_2.CLK.t3 112.468
R273 div2_3_2.CLK.n1 div2_3_2.CLK.t6 112.468
R274 div2_3_2.CLK.n5 div2_3_2.CLK.n4 70.4005
R275 div3_2_0.I.n0 div3_2_0.I.t0 663.801
R276 div3_2_0.I.n0 div3_2_0.I.t6 568.067
R277 div3_2_0.I.t6 div3_2_0.I.t2 514.134
R278 div3_2_0.I.n3 div3_2_0.I.n2 344.8
R279 div3_2_0.I.n1 div3_2_0.I.t3 289.2
R280 div3_2_0.I.t1 div3_2_0.I.n3 275.454
R281 div3_2_0.I.n2 div3_2_0.I.t4 241
R282 div3_2_0.I.n1 div3_2_0.I.t5 112.468
R283 div3_2_0.I.n3 div3_2_0.I.n0 97.9205
R284 div3_2_0.I.n2 div3_2_0.I.n1 64.2672
R285 div3_2_0.G.t0 div3_2_0.G.t1 96.0005
R286 VOUT.n2 VOUT.t4 4546.23
R287 VOUT.t4 VOUT.t3 819.4
R288 VOUT.n1 VOUT.n0 628.734
R289 VOUT.n1 VOUT.t2 257.534
R290 VOUT.n0 VOUT.t1 78.8005
R291 VOUT.n0 VOUT.t0 78.8005
R292 VOUT VOUT.n2 35.2005
R293 VOUT.n2 VOUT.n1 9.6005
R294 div4.t6 div4.t5 819.4
R295 div4.n0 div4.t1 663.801
R296 div4.n0 div4.t6 489.168
R297 div4.t4 div4.t2 401.668
R298 div4.n1 div4.t0 270.12
R299 div4.n2 div4.t4 257.067
R300 div2_3_0.VIN div4.n2 216.9
R301 div4.n2 div4.t3 208.868
R302 div4.n3 div2_3_0.VIN 192.167
R303 div4.n1 div4.n0 67.2005
R304 div4.n3 div4.n1 25.6005
R305 div2_3_2.VOUT div4.n3 4.8005
R306 div8.t3 div8.t2 819.4
R307 div8.n0 div8.t1 663.801
R308 div8.n0 div8.t3 489.168
R309 div8.t4 div8.t5 401.668
R310 div8.n1 div8.t0 270.12
R311 div8.n2 div8.t4 257.067
R312 div3_2_0.VIN div8.n2 216.9
R313 div8.n2 div8.t6 208.868
R314 div8.n3 div3_2_0.VIN 192.167
R315 div8.n1 div8.n0 67.2005
R316 div8.n3 div8.n1 25.6005
R317 div2_3_0.VOUT div8.n3 4.8005
R318 div3_2_0.D.n1 div3_2_0.D.n0 701.467
R319 div3_2_0.D.n1 div3_2_0.D.t0 694.201
R320 div3_2_0.D.n0 div3_2_0.D.t2 321.334
R321 div3_2_0.D.t1 div3_2_0.D.n1 314.921
R322 div3_2_0.D.n0 div3_2_0.D.t3 144.601
R323 div3_2_0.F.t0 div3_2_0.F.t1 96.0005
R324 div3_2_0.E.n0 div3_2_0.E.t0 685.134
R325 div3_2_0.E.n1 div3_2_0.E.t1 663.801
R326 div3_2_0.E.n0 div3_2_0.E.t3 534.268
R327 div3_2_0.E.t2 div3_2_0.E.n1 362.921
R328 div3_2_0.E.n1 div3_2_0.E.n0 91.7338
R329 div3_2_0.H.n0 div3_2_0.H.t1 723.534
R330 div3_2_0.H.n1 div3_2_0.H.t4 553.534
R331 div3_2_0.H.n0 div3_2_0.H.t3 254.333
R332 div3_2_0.H.n2 div3_2_0.H.n1 206.333
R333 div3_2_0.H.n1 div3_2_0.H.n0 70.4005
R334 div3_2_0.H.n2 div3_2_0.H.t2 48.0005
R335 div3_2_0.H.t0 div3_2_0.H.n2 48.0005
R336 div2_3_1.CLK.n5 div2_3_1.CLK.t2 723.534
R337 div2_3_1.CLK.n4 div2_3_1.CLK.t0 723.534
R338 div2_3_1.CLK.n0 div2_3_1.CLK.t7 369.534
R339 div2_3_1.CLK.n3 div2_3_1.CLK.n2 366.856
R340 div2_3_1.CLK.t1 div2_3_1.CLK.n5 254.333
R341 div2_3_1.CLK.n3 div2_3_1.CLK.t6 190.123
R342 div2_3_1.CLK.n4 div2_3_1.CLK.n3 187.201
R343 div2_3_1.CLK.n1 div2_3_1.CLK.n0 176.733
R344 div2_3_1.CLK.n2 div2_3_1.CLK.n1 176.733
R345 div2_3_1.CLK.n0 div2_3_1.CLK.t3 112.468
R346 div2_3_1.CLK.n2 div2_3_1.CLK.t5 112.468
R347 div2_3_1.CLK.n1 div2_3_1.CLK.t4 112.468
R348 div2_3_1.CLK.n5 div2_3_1.CLK.n4 70.4005
R349 div3_2_0.C.n0 div3_2_0.C.t3 721.4
R350 div3_2_0.C.n1 div3_2_0.C.t4 350.349
R351 div3_2_0.C.n0 div3_2_0.C.t2 276.733
R352 div3_2_0.C.n2 div3_2_0.C.n1 206.333
R353 div3_2_0.C.n1 div3_2_0.C.n0 48.0005
R354 div3_2_0.C.n2 div3_2_0.C.t1 48.0005
R355 div3_2_0.C.t0 div3_2_0.C.n2 48.0005
R356 div3_2_0.CLK.n3 div3_2_0.CLK.n2 742.51
R357 div3_2_0.CLK.n8 div3_2_0.CLK.t0 723.534
R358 div3_2_0.CLK.t1 div3_2_0.CLK.n9 723.534
R359 div3_2_0.CLK.n2 div3_2_0.CLK.n1 684.806
R360 div3_2_0.CLK.n7 div3_2_0.CLK.n6 366.856
R361 div3_2_0.CLK.n0 div3_2_0.CLK.t12 337.401
R362 div3_2_0.CLK.n0 div3_2_0.CLK.t8 305.267
R363 div3_2_0.CLK.n9 div3_2_0.CLK.t2 254.333
R364 div3_2_0.CLK.n4 div3_2_0.CLK.n3 224.934
R365 div3_2_0.CLK.n7 div3_2_0.CLK.t9 190.123
R366 div3_2_0.CLK.n8 div3_2_0.CLK.n7 187.201
R367 div3_2_0.CLK.n1 div3_2_0.CLK.n0 176.733
R368 div3_2_0.CLK.n5 div3_2_0.CLK.n4 176.733
R369 div3_2_0.CLK.n6 div3_2_0.CLK.n5 176.733
R370 div3_2_0.CLK.n3 div3_2_0.CLK.t6 144.601
R371 div3_2_0.CLK.n2 div3_2_0.CLK.t3 131.976
R372 div3_2_0.CLK.n0 div3_2_0.CLK.t10 128.534
R373 div3_2_0.CLK.n1 div3_2_0.CLK.t11 128.534
R374 div3_2_0.CLK.n4 div3_2_0.CLK.t4 112.468
R375 div3_2_0.CLK.n6 div3_2_0.CLK.t7 112.468
R376 div3_2_0.CLK.n5 div3_2_0.CLK.t5 112.468
R377 div3_2_0.CLK.n9 div3_2_0.CLK.n8 70.4005
R378 div2_3_2.A.n0 div2_3_2.A.t1 713.933
R379 div2_3_2.A.n0 div2_3_2.A.t2 314.233
R380 div2_3_2.A.t0 div2_3_2.A.n0 308.2
R381 div2_3_2.C.n2 div2_3_2.C.t0 721.4
R382 div2_3_2.C.n1 div2_3_2.C.t4 349.433
R383 div2_3_2.C.t3 div2_3_2.C.n2 276.733
R384 div2_3_2.C.n1 div2_3_2.C.n0 206.333
R385 div2_3_2.C.n0 div2_3_2.C.t2 48.0005
R386 div2_3_2.C.n0 div2_3_2.C.t1 48.0005
R387 div2_3_2.C.n2 div2_3_2.C.n1 48.0005
R388 div3_2_0.A.n0 div3_2_0.A.t1 713.933
R389 div3_2_0.A.n0 div3_2_0.A.t2 314.233
R390 div3_2_0.A.t0 div3_2_0.A.n0 308.2
R391 VIN.t0 VIN.t2 401.668
R392 VIN.n0 VIN.t0 257.067
R393 VIN VIN.n0 216.9
R394 VIN.n0 VIN.t1 208.868
R395 div2_3_1.B.t0 div2_3_1.B.t1 96.0005
R396 div2_3_2.B.t0 div2_3_2.B.t1 96.0005
R397 div3_2_0.B.t0 div3_2_0.B.t1 96.0005
C0 VIN VDDA 0.125773f
C1 VOUT VDDA 0.231994f
C2 VOUT GNDA 2.08651f
C3 VIN GNDA 0.304628f
C4 VDDA GNDA 6.63616f
.ends

