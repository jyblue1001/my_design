magic
tech sky130A
timestamp 1739119761
<< error_p >>
rect 0 14 1 21
rect -12 1 1 14
rect 15 1 16 15
rect -13 0 27 1
rect -25 -24 26 0
rect 2775 -160 3355 -158
rect 3895 -160 3935 -158
rect 3905 -175 3925 -160
rect 2775 -4160 3355 -4158
rect 3895 -4160 3935 -4158
rect 3905 -4175 3925 -4160
<< nwell >>
rect -60 140 2525 280
rect 2775 65 4200 355
rect -60 -1480 1325 -1340
rect -60 -1860 1315 -1720
rect -150 -3460 1290 -2840
rect 1475 -3215 2230 -2840
rect 1475 -3460 2095 -3215
rect 2775 -3935 4200 -3645
rect 1475 -5555 2230 -5310
rect 1475 -5940 2230 -5690
<< nmos >>
rect 0 1 15 50
rect 1 0 15 1
rect 55 0 70 50
rect 260 0 275 50
rect 315 0 330 50
rect 440 0 455 50
rect 495 0 510 50
rect 700 0 715 50
rect 755 0 770 50
rect 880 0 895 50
rect 935 0 950 50
rect 1140 0 1155 50
rect 1195 0 1210 50
rect 1330 0 1345 50
rect 1385 0 1400 50
rect 1590 0 1605 50
rect 1645 0 1660 50
rect 1770 0 1785 50
rect 1825 0 1840 50
rect 1950 0 1965 50
rect 2075 0 2090 50
rect 2200 0 2215 50
rect 2325 0 2340 50
rect 2450 0 2465 50
rect 2865 -145 2880 -45
rect 3010 -145 3025 -45
rect 3155 -145 3170 -45
rect 3300 -145 3315 -45
rect 3445 -145 3460 -45
rect 3590 -145 3605 -45
rect 3735 -145 3750 -45
rect 3880 -145 3895 -45
rect 4025 -145 4040 -45
rect 0 -1250 15 -1200
rect 55 -1250 70 -1200
rect 260 -1250 275 -1200
rect 315 -1250 330 -1200
rect 440 -1250 455 -1200
rect 495 -1250 510 -1200
rect 700 -1250 715 -1200
rect 755 -1250 770 -1200
rect 940 -1250 955 -1200
rect 995 -1250 1010 -1200
rect 1120 -1250 1135 -1200
rect 1245 -1250 1260 -1200
rect 0 -2000 15 -1950
rect 55 -2000 70 -1950
rect 260 -2000 275 -1950
rect 315 -2000 330 -1950
rect 440 -2000 455 -1950
rect 495 -2000 510 -1950
rect 700 -2000 715 -1950
rect 755 -2000 770 -1950
rect 990 -2000 1005 -1950
rect 1115 -2000 1130 -1950
rect 1240 -2000 1255 -1950
rect -90 -2750 -75 -2650
rect -35 -2750 -20 -2650
rect 170 -2750 185 -2650
rect 225 -2750 240 -2650
rect 360 -2750 375 -2650
rect 415 -2750 430 -2650
rect 620 -2750 635 -2650
rect 675 -2750 690 -2650
rect 825 -2750 840 -2650
rect 880 -2750 895 -2650
rect 1045 -2750 1060 -2650
rect 1210 -2750 1225 -2650
rect 1565 -2750 1580 -2650
rect 1710 -2750 1725 -2650
rect 1855 -2750 1870 -2650
rect 2000 -2750 2015 -2650
rect -90 -3650 -75 -3550
rect -35 -3650 -20 -3550
rect 170 -3650 185 -3550
rect 225 -3650 240 -3550
rect 360 -3650 375 -3550
rect 415 -3650 430 -3550
rect 620 -3650 635 -3550
rect 675 -3650 690 -3550
rect 875 -3650 890 -3550
rect 1040 -3650 1055 -3550
rect 1205 -3650 1220 -3550
rect 1565 -3650 1580 -3550
rect 1710 -3650 1725 -3550
rect 1855 -3650 1870 -3550
rect 2000 -3650 2015 -3550
rect 2145 -3650 2160 -3550
rect 2865 -4145 2880 -4045
rect 3010 -4145 3025 -4045
rect 3155 -4145 3170 -4045
rect 3300 -4145 3315 -4045
rect 3445 -4145 3460 -4045
rect 3590 -4145 3605 -4045
rect 3735 -4145 3750 -4045
rect 3880 -4145 3895 -4045
rect 4025 -4145 4040 -4045
rect 1565 -5200 1580 -5100
rect 1710 -5200 1725 -5100
rect 1855 -5200 1870 -5100
rect 2000 -5200 2015 -5100
rect 1565 -6150 1580 -6050
rect 1710 -6150 1725 -6050
rect 1855 -6150 1870 -6050
rect 2000 -6150 2015 -6050
rect 2145 -6150 2160 -6050
<< pmos >>
rect 0 160 15 260
rect 55 160 70 260
rect 260 160 275 260
rect 315 160 330 260
rect 440 160 455 260
rect 495 160 510 260
rect 700 160 715 260
rect 755 160 770 260
rect 880 160 895 260
rect 935 160 950 260
rect 1140 160 1155 260
rect 1195 160 1210 260
rect 1330 160 1345 260
rect 1385 160 1400 260
rect 1590 160 1605 260
rect 1645 160 1660 260
rect 1770 160 1785 260
rect 1825 160 1840 260
rect 1950 160 1965 260
rect 2075 160 2090 260
rect 2200 160 2215 260
rect 2325 160 2340 260
rect 2450 160 2465 260
rect 2865 85 2880 285
rect 3010 85 3025 285
rect 3155 85 3170 285
rect 3300 85 3315 285
rect 3445 85 3460 285
rect 3590 85 3605 285
rect 3735 85 3750 285
rect 3880 85 3895 285
rect 4025 85 4040 285
rect 0 -1460 15 -1360
rect 55 -1460 70 -1360
rect 260 -1460 275 -1360
rect 315 -1460 330 -1360
rect 440 -1460 455 -1360
rect 495 -1460 510 -1360
rect 700 -1460 715 -1360
rect 755 -1460 770 -1360
rect 940 -1460 955 -1360
rect 995 -1460 1010 -1360
rect 1120 -1460 1135 -1360
rect 1245 -1460 1260 -1360
rect 0 -1840 15 -1740
rect 55 -1840 70 -1740
rect 260 -1840 275 -1740
rect 315 -1840 330 -1740
rect 440 -1840 455 -1740
rect 495 -1840 510 -1740
rect 700 -1840 715 -1740
rect 755 -1840 770 -1740
rect 990 -1840 1005 -1740
rect 1115 -1840 1130 -1740
rect 1240 -1840 1255 -1740
rect -90 -3060 -75 -2860
rect -35 -3060 -20 -2860
rect 170 -3060 185 -2860
rect 225 -3060 240 -2860
rect 360 -3060 375 -2860
rect 415 -3060 430 -2860
rect 620 -3060 635 -2860
rect 675 -3060 690 -2860
rect 825 -3060 840 -2860
rect 880 -3060 895 -2860
rect 1045 -3060 1060 -2860
rect 1210 -3060 1225 -2860
rect 1565 -3060 1580 -2860
rect 1710 -3060 1725 -2860
rect 1855 -3060 1870 -2860
rect 2000 -3060 2015 -2860
rect 2145 -3060 2160 -2860
rect -90 -3440 -75 -3240
rect -35 -3440 -20 -3240
rect 170 -3440 185 -3240
rect 225 -3440 240 -3240
rect 360 -3440 375 -3240
rect 415 -3440 430 -3240
rect 620 -3440 635 -3240
rect 675 -3440 690 -3240
rect 875 -3440 890 -3240
rect 1040 -3440 1055 -3240
rect 1205 -3440 1220 -3240
rect 1565 -3440 1580 -3240
rect 1710 -3440 1725 -3240
rect 1855 -3440 1870 -3240
rect 2000 -3440 2015 -3240
rect 2865 -3915 2880 -3715
rect 3010 -3915 3025 -3715
rect 3155 -3915 3170 -3715
rect 3300 -3915 3315 -3715
rect 3445 -3915 3460 -3715
rect 3590 -3915 3605 -3715
rect 3735 -3915 3750 -3715
rect 3880 -3915 3895 -3715
rect 4025 -3915 4040 -3715
rect 1565 -5530 1580 -5330
rect 1710 -5530 1725 -5330
rect 1855 -5530 1870 -5330
rect 2000 -5530 2015 -5330
rect 1565 -5920 1580 -5720
rect 1710 -5920 1725 -5720
rect 1855 -5920 1870 -5720
rect 2000 -5920 2015 -5720
rect 2145 -5920 2160 -5720
<< ndiff >>
rect -40 35 0 50
rect -40 15 -30 35
rect -10 15 0 35
rect -40 0 0 15
rect 15 35 55 50
rect 15 15 25 35
rect 45 15 55 35
rect 15 0 55 15
rect 70 35 110 50
rect 70 15 80 35
rect 100 15 110 35
rect 70 0 110 15
rect 220 35 260 50
rect 220 15 230 35
rect 250 15 260 35
rect 220 0 260 15
rect 275 35 315 50
rect 275 15 285 35
rect 305 15 315 35
rect 275 0 315 15
rect 330 35 370 50
rect 330 15 340 35
rect 360 15 370 35
rect 330 0 370 15
rect 400 35 440 50
rect 400 15 410 35
rect 430 15 440 35
rect 400 0 440 15
rect 455 35 495 50
rect 455 15 465 35
rect 485 15 495 35
rect 455 0 495 15
rect 510 35 550 50
rect 510 15 520 35
rect 540 15 550 35
rect 510 0 550 15
rect 660 35 700 50
rect 660 15 670 35
rect 690 15 700 35
rect 660 0 700 15
rect 715 35 755 50
rect 715 15 725 35
rect 745 15 755 35
rect 715 0 755 15
rect 770 35 810 50
rect 770 15 780 35
rect 800 15 810 35
rect 770 0 810 15
rect 840 35 880 50
rect 840 15 850 35
rect 870 15 880 35
rect 840 0 880 15
rect 895 35 935 50
rect 895 15 905 35
rect 925 15 935 35
rect 895 0 935 15
rect 950 35 990 50
rect 950 15 960 35
rect 980 15 990 35
rect 950 0 990 15
rect 1100 35 1140 50
rect 1100 15 1110 35
rect 1130 15 1140 35
rect 1100 0 1140 15
rect 1155 35 1195 50
rect 1155 15 1165 35
rect 1185 15 1195 35
rect 1155 0 1195 15
rect 1210 35 1250 50
rect 1290 35 1330 50
rect 1210 15 1220 35
rect 1240 15 1250 35
rect 1290 15 1300 35
rect 1320 15 1330 35
rect 1210 0 1250 15
rect 1290 0 1330 15
rect 1345 35 1385 50
rect 1345 15 1355 35
rect 1375 15 1385 35
rect 1345 0 1385 15
rect 1400 35 1440 50
rect 1400 15 1410 35
rect 1430 15 1440 35
rect 1400 0 1440 15
rect 1550 35 1590 50
rect 1550 15 1560 35
rect 1580 15 1590 35
rect 1550 0 1590 15
rect 1605 35 1645 50
rect 1605 15 1615 35
rect 1635 15 1645 35
rect 1605 0 1645 15
rect 1660 35 1700 50
rect 1660 15 1670 35
rect 1690 15 1700 35
rect 1660 0 1700 15
rect 1730 35 1770 50
rect 1730 15 1740 35
rect 1760 15 1770 35
rect 1730 0 1770 15
rect 1785 35 1825 50
rect 1785 15 1795 35
rect 1815 15 1825 35
rect 1785 0 1825 15
rect 1840 35 1880 50
rect 1840 15 1850 35
rect 1870 15 1880 35
rect 1840 0 1880 15
rect 1910 35 1950 50
rect 1910 15 1920 35
rect 1940 15 1950 35
rect 1910 0 1950 15
rect 1965 35 2005 50
rect 1965 15 1975 35
rect 1995 15 2005 35
rect 1965 0 2005 15
rect 2035 35 2075 50
rect 2035 15 2045 35
rect 2065 15 2075 35
rect 2035 0 2075 15
rect 2090 35 2130 50
rect 2090 15 2100 35
rect 2120 15 2130 35
rect 2090 0 2130 15
rect 2160 35 2200 50
rect 2160 15 2170 35
rect 2190 15 2200 35
rect 2160 0 2200 15
rect 2215 35 2255 50
rect 2215 15 2225 35
rect 2245 15 2255 35
rect 2215 0 2255 15
rect 2285 35 2325 50
rect 2285 15 2295 35
rect 2315 15 2325 35
rect 2285 0 2325 15
rect 2340 35 2380 50
rect 2340 15 2350 35
rect 2370 15 2380 35
rect 2340 0 2380 15
rect 2410 35 2450 50
rect 2410 15 2420 35
rect 2440 15 2450 35
rect 2410 0 2450 15
rect 2465 35 2505 50
rect 2465 15 2475 35
rect 2495 15 2505 35
rect 2465 0 2505 15
rect 2815 -60 2865 -45
rect 2815 -130 2830 -60
rect 2850 -130 2865 -60
rect 2815 -145 2865 -130
rect 2880 -60 2930 -45
rect 2880 -130 2895 -60
rect 2915 -130 2930 -60
rect 2880 -145 2930 -130
rect 2960 -60 3010 -45
rect 2960 -130 2975 -60
rect 2995 -130 3010 -60
rect 2960 -145 3010 -130
rect 3025 -60 3075 -45
rect 3025 -130 3040 -60
rect 3060 -130 3075 -60
rect 3025 -145 3075 -130
rect 3105 -60 3155 -45
rect 3105 -130 3120 -60
rect 3140 -130 3155 -60
rect 3105 -145 3155 -130
rect 3170 -60 3220 -45
rect 3170 -130 3185 -60
rect 3205 -130 3220 -60
rect 3170 -145 3220 -130
rect 3250 -60 3300 -45
rect 3250 -130 3265 -60
rect 3285 -130 3300 -60
rect 3250 -145 3300 -130
rect 3315 -60 3365 -45
rect 3315 -130 3330 -60
rect 3350 -130 3365 -60
rect 3315 -145 3365 -130
rect 3395 -60 3445 -45
rect 3395 -130 3410 -60
rect 3430 -130 3445 -60
rect 3395 -145 3445 -130
rect 3460 -60 3510 -45
rect 3460 -130 3475 -60
rect 3495 -130 3510 -60
rect 3460 -145 3510 -130
rect 3540 -60 3590 -45
rect 3540 -130 3555 -60
rect 3575 -130 3590 -60
rect 3540 -145 3590 -130
rect 3605 -60 3655 -45
rect 3605 -130 3620 -60
rect 3640 -130 3655 -60
rect 3605 -145 3655 -130
rect 3685 -60 3735 -45
rect 3685 -130 3700 -60
rect 3720 -130 3735 -60
rect 3685 -145 3735 -130
rect 3750 -60 3800 -45
rect 3750 -130 3765 -60
rect 3785 -130 3800 -60
rect 3750 -145 3800 -130
rect 3830 -60 3880 -45
rect 3830 -130 3845 -60
rect 3865 -130 3880 -60
rect 3830 -145 3880 -130
rect 3895 -60 3945 -45
rect 3895 -130 3910 -60
rect 3930 -130 3945 -60
rect 3895 -145 3945 -130
rect 3975 -60 4025 -45
rect 3975 -130 3990 -60
rect 4010 -130 4025 -60
rect 3975 -145 4025 -130
rect 4040 -60 4090 -45
rect 4040 -130 4055 -60
rect 4075 -130 4090 -60
rect 4040 -145 4090 -130
rect -40 -1215 0 -1200
rect -40 -1235 -30 -1215
rect -10 -1235 0 -1215
rect -40 -1250 0 -1235
rect 15 -1215 55 -1200
rect 15 -1235 25 -1215
rect 45 -1235 55 -1215
rect 15 -1250 55 -1235
rect 70 -1215 110 -1200
rect 70 -1235 80 -1215
rect 100 -1235 110 -1215
rect 70 -1250 110 -1235
rect 220 -1215 260 -1200
rect 220 -1235 230 -1215
rect 250 -1235 260 -1215
rect 220 -1250 260 -1235
rect 275 -1215 315 -1200
rect 275 -1235 285 -1215
rect 305 -1235 315 -1215
rect 275 -1250 315 -1235
rect 330 -1215 370 -1200
rect 330 -1235 340 -1215
rect 360 -1235 370 -1215
rect 330 -1250 370 -1235
rect 400 -1215 440 -1200
rect 400 -1235 410 -1215
rect 430 -1235 440 -1215
rect 400 -1250 440 -1235
rect 455 -1215 495 -1200
rect 455 -1235 465 -1215
rect 485 -1235 495 -1215
rect 455 -1250 495 -1235
rect 510 -1215 550 -1200
rect 510 -1235 520 -1215
rect 540 -1235 550 -1215
rect 510 -1250 550 -1235
rect 660 -1215 700 -1200
rect 660 -1235 670 -1215
rect 690 -1235 700 -1215
rect 660 -1250 700 -1235
rect 715 -1215 755 -1200
rect 715 -1235 725 -1215
rect 745 -1235 755 -1215
rect 715 -1250 755 -1235
rect 770 -1215 810 -1200
rect 770 -1235 780 -1215
rect 800 -1235 810 -1215
rect 770 -1250 810 -1235
rect 900 -1215 940 -1200
rect 900 -1235 910 -1215
rect 930 -1235 940 -1215
rect 900 -1250 940 -1235
rect 955 -1215 995 -1200
rect 955 -1235 965 -1215
rect 985 -1235 995 -1215
rect 955 -1250 995 -1235
rect 1010 -1215 1050 -1200
rect 1010 -1235 1020 -1215
rect 1040 -1235 1050 -1215
rect 1010 -1250 1050 -1235
rect 1080 -1215 1120 -1200
rect 1080 -1235 1090 -1215
rect 1110 -1235 1120 -1215
rect 1080 -1250 1120 -1235
rect 1135 -1215 1175 -1200
rect 1135 -1235 1145 -1215
rect 1165 -1235 1175 -1215
rect 1135 -1250 1175 -1235
rect 1205 -1215 1245 -1200
rect 1205 -1235 1215 -1215
rect 1235 -1235 1245 -1215
rect 1205 -1250 1245 -1235
rect 1260 -1215 1300 -1200
rect 1260 -1235 1270 -1215
rect 1290 -1235 1300 -1215
rect 1260 -1250 1300 -1235
rect -40 -1965 0 -1950
rect -40 -1985 -30 -1965
rect -10 -1985 0 -1965
rect -40 -2000 0 -1985
rect 15 -1965 55 -1950
rect 15 -1985 25 -1965
rect 45 -1985 55 -1965
rect 15 -2000 55 -1985
rect 70 -1965 110 -1950
rect 70 -1985 80 -1965
rect 100 -1985 110 -1965
rect 70 -2000 110 -1985
rect 220 -1965 260 -1950
rect 220 -1985 230 -1965
rect 250 -1985 260 -1965
rect 220 -2000 260 -1985
rect 275 -1965 315 -1950
rect 275 -1985 285 -1965
rect 305 -1985 315 -1965
rect 275 -2000 315 -1985
rect 330 -1965 370 -1950
rect 330 -1985 340 -1965
rect 360 -1985 370 -1965
rect 330 -2000 370 -1985
rect 400 -1965 440 -1950
rect 400 -1985 410 -1965
rect 430 -1985 440 -1965
rect 400 -2000 440 -1985
rect 455 -1965 495 -1950
rect 455 -1985 465 -1965
rect 485 -1985 495 -1965
rect 455 -2000 495 -1985
rect 510 -1965 550 -1950
rect 510 -1985 520 -1965
rect 540 -1985 550 -1965
rect 510 -2000 550 -1985
rect 660 -1965 700 -1950
rect 660 -1985 670 -1965
rect 690 -1985 700 -1965
rect 660 -2000 700 -1985
rect 715 -1965 755 -1950
rect 715 -1985 725 -1965
rect 745 -1985 755 -1965
rect 715 -2000 755 -1985
rect 770 -1965 810 -1950
rect 770 -1985 780 -1965
rect 800 -1985 810 -1965
rect 770 -2000 810 -1985
rect 950 -1965 990 -1950
rect 950 -1985 960 -1965
rect 980 -1985 990 -1965
rect 950 -2000 990 -1985
rect 1005 -1965 1045 -1950
rect 1005 -1985 1015 -1965
rect 1035 -1985 1045 -1965
rect 1005 -2000 1045 -1985
rect 1075 -1965 1115 -1950
rect 1075 -1985 1085 -1965
rect 1105 -1985 1115 -1965
rect 1075 -2000 1115 -1985
rect 1130 -1965 1170 -1950
rect 1130 -1985 1140 -1965
rect 1160 -1985 1170 -1965
rect 1130 -2000 1170 -1985
rect 1200 -1965 1240 -1950
rect 1200 -1985 1210 -1965
rect 1230 -1985 1240 -1965
rect 1200 -2000 1240 -1985
rect 1255 -1965 1295 -1950
rect 1255 -1985 1265 -1965
rect 1285 -1985 1295 -1965
rect 1255 -2000 1295 -1985
rect -130 -2665 -90 -2650
rect -130 -2735 -120 -2665
rect -100 -2735 -90 -2665
rect -130 -2750 -90 -2735
rect -75 -2665 -35 -2650
rect -75 -2735 -65 -2665
rect -45 -2735 -35 -2665
rect -75 -2750 -35 -2735
rect -20 -2665 20 -2650
rect -20 -2735 -10 -2665
rect 10 -2735 20 -2665
rect -20 -2750 20 -2735
rect 130 -2665 170 -2650
rect 130 -2735 140 -2665
rect 160 -2735 170 -2665
rect 130 -2750 170 -2735
rect 185 -2665 225 -2650
rect 185 -2735 195 -2665
rect 215 -2735 225 -2665
rect 185 -2750 225 -2735
rect 240 -2665 280 -2650
rect 240 -2735 250 -2665
rect 270 -2735 280 -2665
rect 240 -2750 280 -2735
rect 320 -2665 360 -2650
rect 320 -2735 330 -2665
rect 350 -2735 360 -2665
rect 320 -2750 360 -2735
rect 375 -2665 415 -2650
rect 375 -2735 385 -2665
rect 405 -2735 415 -2665
rect 375 -2750 415 -2735
rect 430 -2665 470 -2650
rect 430 -2735 440 -2665
rect 460 -2735 470 -2665
rect 430 -2750 470 -2735
rect 580 -2665 620 -2650
rect 580 -2735 590 -2665
rect 610 -2735 620 -2665
rect 580 -2750 620 -2735
rect 635 -2665 675 -2650
rect 635 -2735 645 -2665
rect 665 -2735 675 -2665
rect 635 -2750 675 -2735
rect 690 -2665 730 -2650
rect 690 -2735 700 -2665
rect 720 -2735 730 -2665
rect 690 -2750 730 -2735
rect 785 -2665 825 -2650
rect 785 -2735 795 -2665
rect 815 -2735 825 -2665
rect 785 -2750 825 -2735
rect 840 -2665 880 -2650
rect 840 -2735 850 -2665
rect 870 -2735 880 -2665
rect 840 -2750 880 -2735
rect 895 -2665 935 -2650
rect 895 -2735 905 -2665
rect 925 -2735 935 -2665
rect 895 -2750 935 -2735
rect 1005 -2665 1045 -2650
rect 1005 -2735 1015 -2665
rect 1035 -2735 1045 -2665
rect 1005 -2750 1045 -2735
rect 1060 -2665 1100 -2650
rect 1060 -2735 1070 -2665
rect 1090 -2735 1100 -2665
rect 1060 -2750 1100 -2735
rect 1170 -2665 1210 -2650
rect 1170 -2735 1180 -2665
rect 1200 -2735 1210 -2665
rect 1170 -2750 1210 -2735
rect 1225 -2665 1265 -2650
rect 1225 -2735 1235 -2665
rect 1255 -2735 1265 -2665
rect 1225 -2750 1265 -2735
rect 1515 -2665 1565 -2650
rect 1515 -2685 1530 -2665
rect 1550 -2685 1565 -2665
rect 1515 -2715 1565 -2685
rect 1515 -2735 1530 -2715
rect 1550 -2735 1565 -2715
rect 1515 -2750 1565 -2735
rect 1580 -2665 1630 -2650
rect 1580 -2685 1595 -2665
rect 1615 -2685 1630 -2665
rect 1580 -2715 1630 -2685
rect 1580 -2735 1595 -2715
rect 1615 -2735 1630 -2715
rect 1580 -2750 1630 -2735
rect 1660 -2665 1710 -2650
rect 1660 -2685 1675 -2665
rect 1695 -2685 1710 -2665
rect 1660 -2715 1710 -2685
rect 1660 -2735 1675 -2715
rect 1695 -2735 1710 -2715
rect 1660 -2750 1710 -2735
rect 1725 -2665 1775 -2650
rect 1725 -2685 1740 -2665
rect 1760 -2685 1775 -2665
rect 1725 -2715 1775 -2685
rect 1725 -2735 1740 -2715
rect 1760 -2735 1775 -2715
rect 1725 -2750 1775 -2735
rect 1805 -2665 1855 -2650
rect 1805 -2685 1820 -2665
rect 1840 -2685 1855 -2665
rect 1805 -2715 1855 -2685
rect 1805 -2735 1820 -2715
rect 1840 -2735 1855 -2715
rect 1805 -2750 1855 -2735
rect 1870 -2665 1920 -2650
rect 1870 -2685 1885 -2665
rect 1905 -2685 1920 -2665
rect 1870 -2715 1920 -2685
rect 1870 -2735 1885 -2715
rect 1905 -2735 1920 -2715
rect 1870 -2750 1920 -2735
rect 1950 -2665 2000 -2650
rect 1950 -2685 1965 -2665
rect 1985 -2685 2000 -2665
rect 1950 -2715 2000 -2685
rect 1950 -2735 1965 -2715
rect 1985 -2735 2000 -2715
rect 1950 -2750 2000 -2735
rect 2015 -2665 2065 -2650
rect 2015 -2685 2030 -2665
rect 2050 -2685 2065 -2665
rect 2015 -2715 2065 -2685
rect 2015 -2735 2030 -2715
rect 2050 -2735 2065 -2715
rect 2015 -2750 2065 -2735
rect -130 -3565 -90 -3550
rect -130 -3585 -120 -3565
rect -100 -3585 -90 -3565
rect -130 -3615 -90 -3585
rect -130 -3635 -120 -3615
rect -100 -3635 -90 -3615
rect -130 -3650 -90 -3635
rect -75 -3565 -35 -3550
rect -75 -3585 -65 -3565
rect -45 -3585 -35 -3565
rect -75 -3615 -35 -3585
rect -75 -3635 -65 -3615
rect -45 -3635 -35 -3615
rect -75 -3650 -35 -3635
rect -20 -3565 20 -3550
rect -20 -3585 -10 -3565
rect 10 -3585 20 -3565
rect -20 -3615 20 -3585
rect -20 -3635 -10 -3615
rect 10 -3635 20 -3615
rect -20 -3650 20 -3635
rect 130 -3565 170 -3550
rect 130 -3585 140 -3565
rect 160 -3585 170 -3565
rect 130 -3615 170 -3585
rect 130 -3635 140 -3615
rect 160 -3635 170 -3615
rect 130 -3650 170 -3635
rect 185 -3565 225 -3550
rect 185 -3585 195 -3565
rect 215 -3585 225 -3565
rect 185 -3615 225 -3585
rect 185 -3635 195 -3615
rect 215 -3635 225 -3615
rect 185 -3650 225 -3635
rect 240 -3565 280 -3550
rect 320 -3565 360 -3550
rect 240 -3585 250 -3565
rect 270 -3585 280 -3565
rect 320 -3585 330 -3565
rect 350 -3585 360 -3565
rect 240 -3615 280 -3585
rect 320 -3615 360 -3585
rect 240 -3635 250 -3615
rect 270 -3635 280 -3615
rect 320 -3635 330 -3615
rect 350 -3635 360 -3615
rect 240 -3650 280 -3635
rect 320 -3650 360 -3635
rect 375 -3565 415 -3550
rect 375 -3585 385 -3565
rect 405 -3585 415 -3565
rect 375 -3615 415 -3585
rect 375 -3635 385 -3615
rect 405 -3635 415 -3615
rect 375 -3650 415 -3635
rect 430 -3565 470 -3550
rect 430 -3585 440 -3565
rect 460 -3585 470 -3565
rect 430 -3615 470 -3585
rect 430 -3635 440 -3615
rect 460 -3635 470 -3615
rect 430 -3650 470 -3635
rect 580 -3565 620 -3550
rect 580 -3585 590 -3565
rect 610 -3585 620 -3565
rect 580 -3615 620 -3585
rect 580 -3635 590 -3615
rect 610 -3635 620 -3615
rect 580 -3650 620 -3635
rect 635 -3565 675 -3550
rect 635 -3585 645 -3565
rect 665 -3585 675 -3565
rect 635 -3615 675 -3585
rect 635 -3635 645 -3615
rect 665 -3635 675 -3615
rect 635 -3650 675 -3635
rect 690 -3565 730 -3550
rect 690 -3585 700 -3565
rect 720 -3585 730 -3565
rect 690 -3615 730 -3585
rect 690 -3635 700 -3615
rect 720 -3635 730 -3615
rect 690 -3650 730 -3635
rect 835 -3565 875 -3550
rect 835 -3585 845 -3565
rect 865 -3585 875 -3565
rect 835 -3615 875 -3585
rect 835 -3635 845 -3615
rect 865 -3635 875 -3615
rect 835 -3650 875 -3635
rect 890 -3565 930 -3550
rect 890 -3585 900 -3565
rect 920 -3585 930 -3565
rect 890 -3615 930 -3585
rect 890 -3635 900 -3615
rect 920 -3635 930 -3615
rect 890 -3650 930 -3635
rect 1000 -3565 1040 -3550
rect 1000 -3585 1010 -3565
rect 1030 -3585 1040 -3565
rect 1000 -3615 1040 -3585
rect 1000 -3635 1010 -3615
rect 1030 -3635 1040 -3615
rect 1000 -3650 1040 -3635
rect 1055 -3565 1095 -3550
rect 1055 -3585 1065 -3565
rect 1085 -3585 1095 -3565
rect 1055 -3615 1095 -3585
rect 1055 -3635 1065 -3615
rect 1085 -3635 1095 -3615
rect 1055 -3650 1095 -3635
rect 1165 -3565 1205 -3550
rect 1165 -3585 1175 -3565
rect 1195 -3585 1205 -3565
rect 1165 -3615 1205 -3585
rect 1165 -3635 1175 -3615
rect 1195 -3635 1205 -3615
rect 1165 -3650 1205 -3635
rect 1220 -3565 1260 -3550
rect 1220 -3585 1230 -3565
rect 1250 -3585 1260 -3565
rect 1220 -3615 1260 -3585
rect 1220 -3635 1230 -3615
rect 1250 -3635 1260 -3615
rect 1220 -3650 1260 -3635
rect 1515 -3565 1565 -3550
rect 1515 -3585 1530 -3565
rect 1550 -3585 1565 -3565
rect 1515 -3615 1565 -3585
rect 1515 -3635 1530 -3615
rect 1550 -3635 1565 -3615
rect 1515 -3650 1565 -3635
rect 1580 -3565 1630 -3550
rect 1580 -3585 1595 -3565
rect 1615 -3585 1630 -3565
rect 1580 -3615 1630 -3585
rect 1580 -3635 1595 -3615
rect 1615 -3635 1630 -3615
rect 1580 -3650 1630 -3635
rect 1660 -3565 1710 -3550
rect 1660 -3585 1675 -3565
rect 1695 -3585 1710 -3565
rect 1660 -3615 1710 -3585
rect 1660 -3635 1675 -3615
rect 1695 -3635 1710 -3615
rect 1660 -3650 1710 -3635
rect 1725 -3565 1775 -3550
rect 1725 -3585 1740 -3565
rect 1760 -3585 1775 -3565
rect 1725 -3615 1775 -3585
rect 1725 -3635 1740 -3615
rect 1760 -3635 1775 -3615
rect 1725 -3650 1775 -3635
rect 1805 -3565 1855 -3550
rect 1805 -3585 1820 -3565
rect 1840 -3585 1855 -3565
rect 1805 -3615 1855 -3585
rect 1805 -3635 1820 -3615
rect 1840 -3635 1855 -3615
rect 1805 -3650 1855 -3635
rect 1870 -3565 1920 -3550
rect 1870 -3585 1885 -3565
rect 1905 -3585 1920 -3565
rect 1870 -3615 1920 -3585
rect 1870 -3635 1885 -3615
rect 1905 -3635 1920 -3615
rect 1870 -3650 1920 -3635
rect 1950 -3565 2000 -3550
rect 1950 -3585 1965 -3565
rect 1985 -3585 2000 -3565
rect 1950 -3615 2000 -3585
rect 1950 -3635 1965 -3615
rect 1985 -3635 2000 -3615
rect 1950 -3650 2000 -3635
rect 2015 -3565 2065 -3550
rect 2015 -3585 2030 -3565
rect 2050 -3585 2065 -3565
rect 2015 -3615 2065 -3585
rect 2015 -3635 2030 -3615
rect 2050 -3635 2065 -3615
rect 2015 -3650 2065 -3635
rect 2095 -3565 2145 -3550
rect 2095 -3585 2110 -3565
rect 2130 -3585 2145 -3565
rect 2095 -3615 2145 -3585
rect 2095 -3635 2110 -3615
rect 2130 -3635 2145 -3615
rect 2095 -3650 2145 -3635
rect 2160 -3565 2210 -3550
rect 2160 -3585 2175 -3565
rect 2195 -3585 2210 -3565
rect 2160 -3615 2210 -3585
rect 2160 -3635 2175 -3615
rect 2195 -3635 2210 -3615
rect 2160 -3650 2210 -3635
rect 2815 -4060 2865 -4045
rect 2815 -4130 2830 -4060
rect 2850 -4130 2865 -4060
rect 2815 -4145 2865 -4130
rect 2880 -4060 2930 -4045
rect 2880 -4130 2895 -4060
rect 2915 -4130 2930 -4060
rect 2880 -4145 2930 -4130
rect 2960 -4060 3010 -4045
rect 2960 -4130 2975 -4060
rect 2995 -4130 3010 -4060
rect 2960 -4145 3010 -4130
rect 3025 -4060 3075 -4045
rect 3025 -4130 3040 -4060
rect 3060 -4130 3075 -4060
rect 3025 -4145 3075 -4130
rect 3105 -4060 3155 -4045
rect 3105 -4130 3120 -4060
rect 3140 -4130 3155 -4060
rect 3105 -4145 3155 -4130
rect 3170 -4060 3220 -4045
rect 3170 -4130 3185 -4060
rect 3205 -4130 3220 -4060
rect 3170 -4145 3220 -4130
rect 3250 -4060 3300 -4045
rect 3250 -4130 3265 -4060
rect 3285 -4130 3300 -4060
rect 3250 -4145 3300 -4130
rect 3315 -4060 3365 -4045
rect 3315 -4130 3330 -4060
rect 3350 -4130 3365 -4060
rect 3315 -4145 3365 -4130
rect 3395 -4060 3445 -4045
rect 3395 -4130 3410 -4060
rect 3430 -4130 3445 -4060
rect 3395 -4145 3445 -4130
rect 3460 -4060 3510 -4045
rect 3460 -4130 3475 -4060
rect 3495 -4130 3510 -4060
rect 3460 -4145 3510 -4130
rect 3540 -4060 3590 -4045
rect 3540 -4130 3555 -4060
rect 3575 -4130 3590 -4060
rect 3540 -4145 3590 -4130
rect 3605 -4060 3655 -4045
rect 3605 -4130 3620 -4060
rect 3640 -4130 3655 -4060
rect 3605 -4145 3655 -4130
rect 3685 -4060 3735 -4045
rect 3685 -4130 3700 -4060
rect 3720 -4130 3735 -4060
rect 3685 -4145 3735 -4130
rect 3750 -4060 3800 -4045
rect 3750 -4130 3765 -4060
rect 3785 -4130 3800 -4060
rect 3750 -4145 3800 -4130
rect 3830 -4060 3880 -4045
rect 3830 -4130 3845 -4060
rect 3865 -4130 3880 -4060
rect 3830 -4145 3880 -4130
rect 3895 -4060 3945 -4045
rect 3895 -4130 3910 -4060
rect 3930 -4130 3945 -4060
rect 3895 -4145 3945 -4130
rect 3975 -4060 4025 -4045
rect 3975 -4130 3990 -4060
rect 4010 -4130 4025 -4060
rect 3975 -4145 4025 -4130
rect 4040 -4060 4090 -4045
rect 4040 -4130 4055 -4060
rect 4075 -4130 4090 -4060
rect 4040 -4145 4090 -4130
rect 1515 -5115 1565 -5100
rect 1515 -5135 1530 -5115
rect 1550 -5135 1565 -5115
rect 1515 -5165 1565 -5135
rect 1515 -5185 1530 -5165
rect 1550 -5185 1565 -5165
rect 1515 -5200 1565 -5185
rect 1580 -5115 1630 -5100
rect 1580 -5135 1595 -5115
rect 1615 -5135 1630 -5115
rect 1580 -5165 1630 -5135
rect 1580 -5185 1595 -5165
rect 1615 -5185 1630 -5165
rect 1580 -5200 1630 -5185
rect 1660 -5115 1710 -5100
rect 1660 -5135 1675 -5115
rect 1695 -5135 1710 -5115
rect 1660 -5165 1710 -5135
rect 1660 -5185 1675 -5165
rect 1695 -5185 1710 -5165
rect 1660 -5200 1710 -5185
rect 1725 -5115 1775 -5100
rect 1725 -5135 1740 -5115
rect 1760 -5135 1775 -5115
rect 1725 -5165 1775 -5135
rect 1725 -5185 1740 -5165
rect 1760 -5185 1775 -5165
rect 1725 -5200 1775 -5185
rect 1805 -5115 1855 -5100
rect 1805 -5135 1820 -5115
rect 1840 -5135 1855 -5115
rect 1805 -5165 1855 -5135
rect 1805 -5185 1820 -5165
rect 1840 -5185 1855 -5165
rect 1805 -5200 1855 -5185
rect 1870 -5115 1920 -5100
rect 1870 -5135 1885 -5115
rect 1905 -5135 1920 -5115
rect 1870 -5165 1920 -5135
rect 1870 -5185 1885 -5165
rect 1905 -5185 1920 -5165
rect 1870 -5200 1920 -5185
rect 1950 -5115 2000 -5100
rect 1950 -5135 1965 -5115
rect 1985 -5135 2000 -5115
rect 1950 -5165 2000 -5135
rect 1950 -5185 1965 -5165
rect 1985 -5185 2000 -5165
rect 1950 -5200 2000 -5185
rect 2015 -5115 2065 -5100
rect 2015 -5135 2030 -5115
rect 2050 -5135 2065 -5115
rect 2015 -5165 2065 -5135
rect 2015 -5185 2030 -5165
rect 2050 -5185 2065 -5165
rect 2015 -5200 2065 -5185
rect 1515 -6065 1565 -6050
rect 1515 -6085 1530 -6065
rect 1550 -6085 1565 -6065
rect 1515 -6115 1565 -6085
rect 1515 -6135 1530 -6115
rect 1550 -6135 1565 -6115
rect 1515 -6150 1565 -6135
rect 1580 -6065 1630 -6050
rect 1580 -6085 1595 -6065
rect 1615 -6085 1630 -6065
rect 1580 -6115 1630 -6085
rect 1580 -6135 1595 -6115
rect 1615 -6135 1630 -6115
rect 1580 -6150 1630 -6135
rect 1660 -6065 1710 -6050
rect 1660 -6085 1675 -6065
rect 1695 -6085 1710 -6065
rect 1660 -6115 1710 -6085
rect 1660 -6135 1675 -6115
rect 1695 -6135 1710 -6115
rect 1660 -6150 1710 -6135
rect 1725 -6065 1775 -6050
rect 1725 -6085 1740 -6065
rect 1760 -6085 1775 -6065
rect 1725 -6115 1775 -6085
rect 1725 -6135 1740 -6115
rect 1760 -6135 1775 -6115
rect 1725 -6150 1775 -6135
rect 1805 -6065 1855 -6050
rect 1805 -6085 1820 -6065
rect 1840 -6085 1855 -6065
rect 1805 -6115 1855 -6085
rect 1805 -6135 1820 -6115
rect 1840 -6135 1855 -6115
rect 1805 -6150 1855 -6135
rect 1870 -6065 1920 -6050
rect 1870 -6085 1885 -6065
rect 1905 -6085 1920 -6065
rect 1870 -6115 1920 -6085
rect 1870 -6135 1885 -6115
rect 1905 -6135 1920 -6115
rect 1870 -6150 1920 -6135
rect 1950 -6065 2000 -6050
rect 1950 -6085 1965 -6065
rect 1985 -6085 2000 -6065
rect 1950 -6115 2000 -6085
rect 1950 -6135 1965 -6115
rect 1985 -6135 2000 -6115
rect 1950 -6150 2000 -6135
rect 2015 -6065 2065 -6050
rect 2015 -6085 2030 -6065
rect 2050 -6085 2065 -6065
rect 2015 -6115 2065 -6085
rect 2015 -6135 2030 -6115
rect 2050 -6135 2065 -6115
rect 2015 -6150 2065 -6135
rect 2095 -6065 2145 -6050
rect 2095 -6085 2110 -6065
rect 2130 -6085 2145 -6065
rect 2095 -6115 2145 -6085
rect 2095 -6135 2110 -6115
rect 2130 -6135 2145 -6115
rect 2095 -6150 2145 -6135
rect 2160 -6065 2210 -6050
rect 2160 -6085 2175 -6065
rect 2195 -6085 2210 -6065
rect 2160 -6115 2210 -6085
rect 2160 -6135 2175 -6115
rect 2195 -6135 2210 -6115
rect 2160 -6150 2210 -6135
<< pdiff >>
rect -40 245 0 260
rect -40 175 -30 245
rect -10 175 0 245
rect -40 160 0 175
rect 15 245 55 260
rect 15 175 25 245
rect 45 175 55 245
rect 15 160 55 175
rect 70 245 110 260
rect 70 175 80 245
rect 100 175 110 245
rect 70 160 110 175
rect 220 245 260 260
rect 220 175 230 245
rect 250 175 260 245
rect 220 160 260 175
rect 275 245 315 260
rect 275 175 285 245
rect 305 175 315 245
rect 275 160 315 175
rect 330 245 370 260
rect 330 175 340 245
rect 360 175 370 245
rect 330 160 370 175
rect 400 245 440 260
rect 400 175 410 245
rect 430 175 440 245
rect 400 160 440 175
rect 455 245 495 260
rect 455 175 465 245
rect 485 175 495 245
rect 455 160 495 175
rect 510 245 550 260
rect 510 175 520 245
rect 540 175 550 245
rect 510 160 550 175
rect 660 245 700 260
rect 660 175 670 245
rect 690 175 700 245
rect 660 160 700 175
rect 715 245 755 260
rect 715 175 725 245
rect 745 175 755 245
rect 715 160 755 175
rect 770 245 810 260
rect 770 175 780 245
rect 800 175 810 245
rect 770 160 810 175
rect 840 245 880 260
rect 840 175 850 245
rect 870 175 880 245
rect 840 160 880 175
rect 895 245 935 260
rect 895 175 905 245
rect 925 175 935 245
rect 895 160 935 175
rect 950 245 990 260
rect 950 175 960 245
rect 980 175 990 245
rect 950 160 990 175
rect 1100 245 1140 260
rect 1100 175 1110 245
rect 1130 175 1140 245
rect 1100 160 1140 175
rect 1155 245 1195 260
rect 1155 175 1165 245
rect 1185 175 1195 245
rect 1155 160 1195 175
rect 1210 245 1250 260
rect 1290 245 1330 260
rect 1210 175 1220 245
rect 1240 175 1250 245
rect 1290 175 1300 245
rect 1320 175 1330 245
rect 1210 160 1250 175
rect 1290 160 1330 175
rect 1345 245 1385 260
rect 1345 175 1355 245
rect 1375 175 1385 245
rect 1345 160 1385 175
rect 1400 245 1440 260
rect 1400 175 1410 245
rect 1430 175 1440 245
rect 1400 160 1440 175
rect 1550 245 1590 260
rect 1550 175 1560 245
rect 1580 175 1590 245
rect 1550 160 1590 175
rect 1605 245 1645 260
rect 1605 175 1615 245
rect 1635 175 1645 245
rect 1605 160 1645 175
rect 1660 245 1700 260
rect 1660 175 1670 245
rect 1690 175 1700 245
rect 1660 160 1700 175
rect 1730 245 1770 260
rect 1730 175 1740 245
rect 1760 175 1770 245
rect 1730 160 1770 175
rect 1785 245 1825 260
rect 1785 175 1795 245
rect 1815 175 1825 245
rect 1785 160 1825 175
rect 1840 245 1880 260
rect 1840 175 1850 245
rect 1870 175 1880 245
rect 1840 160 1880 175
rect 1910 245 1950 260
rect 1910 175 1920 245
rect 1940 175 1950 245
rect 1910 160 1950 175
rect 1965 245 2005 260
rect 1965 175 1975 245
rect 1995 175 2005 245
rect 1965 160 2005 175
rect 2035 245 2075 260
rect 2035 175 2045 245
rect 2065 175 2075 245
rect 2035 160 2075 175
rect 2090 245 2130 260
rect 2090 175 2100 245
rect 2120 175 2130 245
rect 2090 160 2130 175
rect 2160 245 2200 260
rect 2160 175 2170 245
rect 2190 175 2200 245
rect 2160 160 2200 175
rect 2215 245 2255 260
rect 2215 175 2225 245
rect 2245 175 2255 245
rect 2215 160 2255 175
rect 2285 245 2325 260
rect 2285 175 2295 245
rect 2315 175 2325 245
rect 2285 160 2325 175
rect 2340 245 2380 260
rect 2340 175 2350 245
rect 2370 175 2380 245
rect 2340 160 2380 175
rect 2410 245 2450 260
rect 2410 175 2420 245
rect 2440 175 2450 245
rect 2410 160 2450 175
rect 2465 245 2505 260
rect 2465 175 2475 245
rect 2495 175 2505 245
rect 2465 160 2505 175
rect 2815 270 2865 285
rect 2815 100 2830 270
rect 2850 100 2865 270
rect 2815 85 2865 100
rect 2880 270 2930 285
rect 2880 100 2895 270
rect 2915 100 2930 270
rect 2880 85 2930 100
rect 2960 270 3010 285
rect 2960 100 2975 270
rect 2995 100 3010 270
rect 2960 85 3010 100
rect 3025 270 3075 285
rect 3025 100 3040 270
rect 3060 100 3075 270
rect 3025 85 3075 100
rect 3105 270 3155 285
rect 3105 100 3120 270
rect 3140 100 3155 270
rect 3105 85 3155 100
rect 3170 270 3220 285
rect 3170 100 3185 270
rect 3205 100 3220 270
rect 3170 85 3220 100
rect 3250 270 3300 285
rect 3250 100 3265 270
rect 3285 100 3300 270
rect 3250 85 3300 100
rect 3315 270 3365 285
rect 3315 100 3330 270
rect 3350 100 3365 270
rect 3315 85 3365 100
rect 3395 270 3445 285
rect 3395 100 3410 270
rect 3430 100 3445 270
rect 3395 85 3445 100
rect 3460 270 3510 285
rect 3460 100 3475 270
rect 3495 100 3510 270
rect 3460 85 3510 100
rect 3540 270 3590 285
rect 3540 100 3555 270
rect 3575 100 3590 270
rect 3540 85 3590 100
rect 3605 270 3655 285
rect 3605 100 3620 270
rect 3640 100 3655 270
rect 3605 85 3655 100
rect 3685 270 3735 285
rect 3685 100 3700 270
rect 3720 100 3735 270
rect 3685 85 3735 100
rect 3750 270 3800 285
rect 3750 100 3765 270
rect 3785 100 3800 270
rect 3750 85 3800 100
rect 3830 270 3880 285
rect 3830 100 3845 270
rect 3865 100 3880 270
rect 3830 85 3880 100
rect 3895 270 3945 285
rect 3895 100 3910 270
rect 3930 100 3945 270
rect 3895 85 3945 100
rect 3975 270 4025 285
rect 3975 100 3990 270
rect 4010 100 4025 270
rect 3975 85 4025 100
rect 4040 270 4090 285
rect 4040 100 4055 270
rect 4075 100 4090 270
rect 4040 85 4090 100
rect -40 -1375 0 -1360
rect -40 -1445 -30 -1375
rect -10 -1445 0 -1375
rect -40 -1460 0 -1445
rect 15 -1375 55 -1360
rect 15 -1445 25 -1375
rect 45 -1445 55 -1375
rect 15 -1460 55 -1445
rect 70 -1375 110 -1360
rect 70 -1445 80 -1375
rect 100 -1445 110 -1375
rect 70 -1460 110 -1445
rect 220 -1375 260 -1360
rect 220 -1445 230 -1375
rect 250 -1445 260 -1375
rect 220 -1460 260 -1445
rect 275 -1375 315 -1360
rect 275 -1445 285 -1375
rect 305 -1445 315 -1375
rect 275 -1460 315 -1445
rect 330 -1375 370 -1360
rect 330 -1445 340 -1375
rect 360 -1445 370 -1375
rect 330 -1460 370 -1445
rect 400 -1375 440 -1360
rect 400 -1445 410 -1375
rect 430 -1445 440 -1375
rect 400 -1460 440 -1445
rect 455 -1375 495 -1360
rect 455 -1445 465 -1375
rect 485 -1445 495 -1375
rect 455 -1460 495 -1445
rect 510 -1375 550 -1360
rect 510 -1445 520 -1375
rect 540 -1445 550 -1375
rect 510 -1460 550 -1445
rect 660 -1375 700 -1360
rect 660 -1445 670 -1375
rect 690 -1445 700 -1375
rect 660 -1460 700 -1445
rect 715 -1375 755 -1360
rect 715 -1445 725 -1375
rect 745 -1445 755 -1375
rect 715 -1460 755 -1445
rect 770 -1375 810 -1360
rect 770 -1445 780 -1375
rect 800 -1445 810 -1375
rect 770 -1460 810 -1445
rect 900 -1375 940 -1360
rect 900 -1445 910 -1375
rect 930 -1445 940 -1375
rect 900 -1460 940 -1445
rect 955 -1375 995 -1360
rect 955 -1445 965 -1375
rect 985 -1445 995 -1375
rect 955 -1460 995 -1445
rect 1010 -1375 1050 -1360
rect 1010 -1445 1020 -1375
rect 1040 -1445 1050 -1375
rect 1010 -1460 1050 -1445
rect 1080 -1375 1120 -1360
rect 1080 -1445 1090 -1375
rect 1110 -1445 1120 -1375
rect 1080 -1460 1120 -1445
rect 1135 -1375 1175 -1360
rect 1135 -1445 1145 -1375
rect 1165 -1445 1175 -1375
rect 1135 -1460 1175 -1445
rect 1205 -1375 1245 -1360
rect 1205 -1445 1215 -1375
rect 1235 -1445 1245 -1375
rect 1205 -1460 1245 -1445
rect 1260 -1375 1300 -1360
rect 1260 -1445 1270 -1375
rect 1290 -1445 1300 -1375
rect 1260 -1460 1300 -1445
rect -40 -1755 0 -1740
rect -40 -1825 -30 -1755
rect -10 -1825 0 -1755
rect -40 -1840 0 -1825
rect 15 -1755 55 -1740
rect 15 -1825 25 -1755
rect 45 -1825 55 -1755
rect 15 -1840 55 -1825
rect 70 -1755 110 -1740
rect 70 -1825 80 -1755
rect 100 -1825 110 -1755
rect 70 -1840 110 -1825
rect 220 -1755 260 -1740
rect 220 -1825 230 -1755
rect 250 -1825 260 -1755
rect 220 -1840 260 -1825
rect 275 -1755 315 -1740
rect 275 -1825 285 -1755
rect 305 -1825 315 -1755
rect 275 -1840 315 -1825
rect 330 -1755 370 -1740
rect 330 -1825 340 -1755
rect 360 -1825 370 -1755
rect 330 -1840 370 -1825
rect 400 -1755 440 -1740
rect 400 -1825 410 -1755
rect 430 -1825 440 -1755
rect 400 -1840 440 -1825
rect 455 -1755 495 -1740
rect 455 -1825 465 -1755
rect 485 -1825 495 -1755
rect 455 -1840 495 -1825
rect 510 -1755 550 -1740
rect 510 -1825 520 -1755
rect 540 -1825 550 -1755
rect 510 -1840 550 -1825
rect 660 -1755 700 -1740
rect 660 -1825 670 -1755
rect 690 -1825 700 -1755
rect 660 -1840 700 -1825
rect 715 -1755 755 -1740
rect 715 -1825 725 -1755
rect 745 -1825 755 -1755
rect 715 -1840 755 -1825
rect 770 -1755 810 -1740
rect 770 -1825 780 -1755
rect 800 -1825 810 -1755
rect 770 -1840 810 -1825
rect 950 -1755 990 -1740
rect 950 -1825 960 -1755
rect 980 -1825 990 -1755
rect 950 -1840 990 -1825
rect 1005 -1755 1045 -1740
rect 1005 -1825 1015 -1755
rect 1035 -1825 1045 -1755
rect 1005 -1840 1045 -1825
rect 1075 -1755 1115 -1740
rect 1075 -1825 1085 -1755
rect 1105 -1825 1115 -1755
rect 1075 -1840 1115 -1825
rect 1130 -1755 1170 -1740
rect 1130 -1825 1140 -1755
rect 1160 -1825 1170 -1755
rect 1130 -1840 1170 -1825
rect 1200 -1755 1240 -1740
rect 1200 -1825 1210 -1755
rect 1230 -1825 1240 -1755
rect 1200 -1840 1240 -1825
rect 1255 -1755 1295 -1740
rect 1255 -1825 1265 -1755
rect 1285 -1825 1295 -1755
rect 1255 -1840 1295 -1825
rect -130 -2875 -90 -2860
rect -130 -2895 -120 -2875
rect -100 -2895 -90 -2875
rect -130 -2925 -90 -2895
rect -130 -2945 -120 -2925
rect -100 -2945 -90 -2925
rect -130 -2975 -90 -2945
rect -130 -2995 -120 -2975
rect -100 -2995 -90 -2975
rect -130 -3025 -90 -2995
rect -130 -3045 -120 -3025
rect -100 -3045 -90 -3025
rect -130 -3060 -90 -3045
rect -75 -2875 -35 -2860
rect -75 -2895 -65 -2875
rect -45 -2895 -35 -2875
rect -75 -2925 -35 -2895
rect -75 -2945 -65 -2925
rect -45 -2945 -35 -2925
rect -75 -2975 -35 -2945
rect -75 -2995 -65 -2975
rect -45 -2995 -35 -2975
rect -75 -3025 -35 -2995
rect -75 -3045 -65 -3025
rect -45 -3045 -35 -3025
rect -75 -3060 -35 -3045
rect -20 -2875 20 -2860
rect -20 -2895 -10 -2875
rect 10 -2895 20 -2875
rect -20 -2925 20 -2895
rect -20 -2945 -10 -2925
rect 10 -2945 20 -2925
rect -20 -2975 20 -2945
rect -20 -2995 -10 -2975
rect 10 -2995 20 -2975
rect -20 -3025 20 -2995
rect -20 -3045 -10 -3025
rect 10 -3045 20 -3025
rect -20 -3060 20 -3045
rect 130 -2875 170 -2860
rect 130 -2895 140 -2875
rect 160 -2895 170 -2875
rect 130 -2925 170 -2895
rect 130 -2945 140 -2925
rect 160 -2945 170 -2925
rect 130 -2975 170 -2945
rect 130 -2995 140 -2975
rect 160 -2995 170 -2975
rect 130 -3025 170 -2995
rect 130 -3045 140 -3025
rect 160 -3045 170 -3025
rect 130 -3060 170 -3045
rect 185 -2875 225 -2860
rect 185 -2895 195 -2875
rect 215 -2895 225 -2875
rect 185 -2925 225 -2895
rect 185 -2945 195 -2925
rect 215 -2945 225 -2925
rect 185 -2975 225 -2945
rect 185 -2995 195 -2975
rect 215 -2995 225 -2975
rect 185 -3025 225 -2995
rect 185 -3045 195 -3025
rect 215 -3045 225 -3025
rect 185 -3060 225 -3045
rect 240 -2875 280 -2860
rect 240 -2895 250 -2875
rect 270 -2895 280 -2875
rect 240 -2925 280 -2895
rect 240 -2945 250 -2925
rect 270 -2945 280 -2925
rect 240 -2975 280 -2945
rect 240 -2995 250 -2975
rect 270 -2995 280 -2975
rect 240 -3025 280 -2995
rect 240 -3045 250 -3025
rect 270 -3045 280 -3025
rect 240 -3060 280 -3045
rect 320 -2875 360 -2860
rect 320 -2895 330 -2875
rect 350 -2895 360 -2875
rect 320 -2925 360 -2895
rect 320 -2945 330 -2925
rect 350 -2945 360 -2925
rect 320 -2975 360 -2945
rect 320 -2995 330 -2975
rect 350 -2995 360 -2975
rect 320 -3025 360 -2995
rect 320 -3045 330 -3025
rect 350 -3045 360 -3025
rect 320 -3060 360 -3045
rect 375 -2875 415 -2860
rect 375 -2895 385 -2875
rect 405 -2895 415 -2875
rect 375 -2925 415 -2895
rect 375 -2945 385 -2925
rect 405 -2945 415 -2925
rect 375 -2975 415 -2945
rect 375 -2995 385 -2975
rect 405 -2995 415 -2975
rect 375 -3025 415 -2995
rect 375 -3045 385 -3025
rect 405 -3045 415 -3025
rect 375 -3060 415 -3045
rect 430 -2875 470 -2860
rect 430 -2895 440 -2875
rect 460 -2895 470 -2875
rect 430 -2925 470 -2895
rect 430 -2945 440 -2925
rect 460 -2945 470 -2925
rect 430 -2975 470 -2945
rect 430 -2995 440 -2975
rect 460 -2995 470 -2975
rect 430 -3025 470 -2995
rect 430 -3045 440 -3025
rect 460 -3045 470 -3025
rect 430 -3060 470 -3045
rect 580 -2875 620 -2860
rect 580 -2895 590 -2875
rect 610 -2895 620 -2875
rect 580 -2925 620 -2895
rect 580 -2945 590 -2925
rect 610 -2945 620 -2925
rect 580 -2975 620 -2945
rect 580 -2995 590 -2975
rect 610 -2995 620 -2975
rect 580 -3025 620 -2995
rect 580 -3045 590 -3025
rect 610 -3045 620 -3025
rect 580 -3060 620 -3045
rect 635 -2875 675 -2860
rect 635 -2895 645 -2875
rect 665 -2895 675 -2875
rect 635 -2925 675 -2895
rect 635 -2945 645 -2925
rect 665 -2945 675 -2925
rect 635 -2975 675 -2945
rect 635 -2995 645 -2975
rect 665 -2995 675 -2975
rect 635 -3025 675 -2995
rect 635 -3045 645 -3025
rect 665 -3045 675 -3025
rect 635 -3060 675 -3045
rect 690 -2875 730 -2860
rect 690 -2895 700 -2875
rect 720 -2895 730 -2875
rect 690 -2925 730 -2895
rect 690 -2945 700 -2925
rect 720 -2945 730 -2925
rect 690 -2975 730 -2945
rect 690 -2995 700 -2975
rect 720 -2995 730 -2975
rect 690 -3025 730 -2995
rect 690 -3045 700 -3025
rect 720 -3045 730 -3025
rect 690 -3060 730 -3045
rect 785 -2875 825 -2860
rect 785 -2895 795 -2875
rect 815 -2895 825 -2875
rect 785 -2925 825 -2895
rect 785 -2945 795 -2925
rect 815 -2945 825 -2925
rect 785 -2975 825 -2945
rect 785 -2995 795 -2975
rect 815 -2995 825 -2975
rect 785 -3025 825 -2995
rect 785 -3045 795 -3025
rect 815 -3045 825 -3025
rect 785 -3060 825 -3045
rect 840 -2875 880 -2860
rect 840 -2895 850 -2875
rect 870 -2895 880 -2875
rect 840 -2925 880 -2895
rect 840 -2945 850 -2925
rect 870 -2945 880 -2925
rect 840 -2975 880 -2945
rect 840 -2995 850 -2975
rect 870 -2995 880 -2975
rect 840 -3025 880 -2995
rect 840 -3045 850 -3025
rect 870 -3045 880 -3025
rect 840 -3060 880 -3045
rect 895 -2875 935 -2860
rect 895 -2895 905 -2875
rect 925 -2895 935 -2875
rect 895 -2925 935 -2895
rect 895 -2945 905 -2925
rect 925 -2945 935 -2925
rect 895 -2975 935 -2945
rect 895 -2995 905 -2975
rect 925 -2995 935 -2975
rect 895 -3025 935 -2995
rect 895 -3045 905 -3025
rect 925 -3045 935 -3025
rect 895 -3060 935 -3045
rect 1005 -2875 1045 -2860
rect 1005 -2895 1015 -2875
rect 1035 -2895 1045 -2875
rect 1005 -2925 1045 -2895
rect 1005 -2945 1015 -2925
rect 1035 -2945 1045 -2925
rect 1005 -2975 1045 -2945
rect 1005 -2995 1015 -2975
rect 1035 -2995 1045 -2975
rect 1005 -3025 1045 -2995
rect 1005 -3045 1015 -3025
rect 1035 -3045 1045 -3025
rect 1005 -3060 1045 -3045
rect 1060 -2875 1100 -2860
rect 1060 -2895 1070 -2875
rect 1090 -2895 1100 -2875
rect 1060 -2925 1100 -2895
rect 1060 -2945 1070 -2925
rect 1090 -2945 1100 -2925
rect 1060 -2975 1100 -2945
rect 1060 -2995 1070 -2975
rect 1090 -2995 1100 -2975
rect 1060 -3025 1100 -2995
rect 1060 -3045 1070 -3025
rect 1090 -3045 1100 -3025
rect 1060 -3060 1100 -3045
rect 1170 -2875 1210 -2860
rect 1170 -2895 1180 -2875
rect 1200 -2895 1210 -2875
rect 1170 -2925 1210 -2895
rect 1170 -2945 1180 -2925
rect 1200 -2945 1210 -2925
rect 1170 -2975 1210 -2945
rect 1170 -2995 1180 -2975
rect 1200 -2995 1210 -2975
rect 1170 -3025 1210 -2995
rect 1170 -3045 1180 -3025
rect 1200 -3045 1210 -3025
rect 1170 -3060 1210 -3045
rect 1225 -2875 1265 -2860
rect 1225 -2895 1235 -2875
rect 1255 -2895 1265 -2875
rect 1225 -2925 1265 -2895
rect 1225 -2945 1235 -2925
rect 1255 -2945 1265 -2925
rect 1225 -2975 1265 -2945
rect 1225 -2995 1235 -2975
rect 1255 -2995 1265 -2975
rect 1225 -3025 1265 -2995
rect 1225 -3045 1235 -3025
rect 1255 -3045 1265 -3025
rect 1225 -3060 1265 -3045
rect 1515 -2875 1565 -2860
rect 1515 -2895 1530 -2875
rect 1550 -2895 1565 -2875
rect 1515 -2925 1565 -2895
rect 1515 -2945 1530 -2925
rect 1550 -2945 1565 -2925
rect 1515 -2975 1565 -2945
rect 1515 -2995 1530 -2975
rect 1550 -2995 1565 -2975
rect 1515 -3025 1565 -2995
rect 1515 -3045 1530 -3025
rect 1550 -3045 1565 -3025
rect 1515 -3060 1565 -3045
rect 1580 -2875 1630 -2860
rect 1580 -2895 1595 -2875
rect 1615 -2895 1630 -2875
rect 1580 -2925 1630 -2895
rect 1580 -2945 1595 -2925
rect 1615 -2945 1630 -2925
rect 1580 -2975 1630 -2945
rect 1580 -2995 1595 -2975
rect 1615 -2995 1630 -2975
rect 1580 -3025 1630 -2995
rect 1580 -3045 1595 -3025
rect 1615 -3045 1630 -3025
rect 1580 -3060 1630 -3045
rect 1660 -2875 1710 -2860
rect 1660 -2895 1675 -2875
rect 1695 -2895 1710 -2875
rect 1660 -2925 1710 -2895
rect 1660 -2945 1675 -2925
rect 1695 -2945 1710 -2925
rect 1660 -2975 1710 -2945
rect 1660 -2995 1675 -2975
rect 1695 -2995 1710 -2975
rect 1660 -3025 1710 -2995
rect 1660 -3045 1675 -3025
rect 1695 -3045 1710 -3025
rect 1660 -3060 1710 -3045
rect 1725 -2875 1775 -2860
rect 1725 -2895 1740 -2875
rect 1760 -2895 1775 -2875
rect 1725 -2925 1775 -2895
rect 1725 -2945 1740 -2925
rect 1760 -2945 1775 -2925
rect 1725 -2975 1775 -2945
rect 1725 -2995 1740 -2975
rect 1760 -2995 1775 -2975
rect 1725 -3025 1775 -2995
rect 1725 -3045 1740 -3025
rect 1760 -3045 1775 -3025
rect 1725 -3060 1775 -3045
rect 1805 -2875 1855 -2860
rect 1805 -2895 1820 -2875
rect 1840 -2895 1855 -2875
rect 1805 -2925 1855 -2895
rect 1805 -2945 1820 -2925
rect 1840 -2945 1855 -2925
rect 1805 -2975 1855 -2945
rect 1805 -2995 1820 -2975
rect 1840 -2995 1855 -2975
rect 1805 -3025 1855 -2995
rect 1805 -3045 1820 -3025
rect 1840 -3045 1855 -3025
rect 1805 -3060 1855 -3045
rect 1870 -2875 1920 -2860
rect 1870 -2895 1885 -2875
rect 1905 -2895 1920 -2875
rect 1870 -2925 1920 -2895
rect 1870 -2945 1885 -2925
rect 1905 -2945 1920 -2925
rect 1870 -2975 1920 -2945
rect 1870 -2995 1885 -2975
rect 1905 -2995 1920 -2975
rect 1870 -3025 1920 -2995
rect 1870 -3045 1885 -3025
rect 1905 -3045 1920 -3025
rect 1870 -3060 1920 -3045
rect 1950 -2875 2000 -2860
rect 1950 -2895 1965 -2875
rect 1985 -2895 2000 -2875
rect 1950 -2925 2000 -2895
rect 1950 -2945 1965 -2925
rect 1985 -2945 2000 -2925
rect 1950 -2975 2000 -2945
rect 1950 -2995 1965 -2975
rect 1985 -2995 2000 -2975
rect 1950 -3025 2000 -2995
rect 1950 -3045 1965 -3025
rect 1985 -3045 2000 -3025
rect 1950 -3060 2000 -3045
rect 2015 -2875 2065 -2860
rect 2015 -2895 2030 -2875
rect 2050 -2895 2065 -2875
rect 2015 -2925 2065 -2895
rect 2015 -2945 2030 -2925
rect 2050 -2945 2065 -2925
rect 2015 -2975 2065 -2945
rect 2015 -2995 2030 -2975
rect 2050 -2995 2065 -2975
rect 2015 -3025 2065 -2995
rect 2015 -3045 2030 -3025
rect 2050 -3045 2065 -3025
rect 2015 -3060 2065 -3045
rect 2095 -2875 2145 -2860
rect 2095 -2895 2110 -2875
rect 2130 -2895 2145 -2875
rect 2095 -2925 2145 -2895
rect 2095 -2945 2110 -2925
rect 2130 -2945 2145 -2925
rect 2095 -2975 2145 -2945
rect 2095 -2995 2110 -2975
rect 2130 -2995 2145 -2975
rect 2095 -3025 2145 -2995
rect 2095 -3045 2110 -3025
rect 2130 -3045 2145 -3025
rect 2095 -3060 2145 -3045
rect 2160 -2875 2210 -2860
rect 2160 -2895 2175 -2875
rect 2195 -2895 2210 -2875
rect 2160 -2925 2210 -2895
rect 2160 -2945 2175 -2925
rect 2195 -2945 2210 -2925
rect 2160 -2975 2210 -2945
rect 2160 -2995 2175 -2975
rect 2195 -2995 2210 -2975
rect 2160 -3025 2210 -2995
rect 2160 -3045 2175 -3025
rect 2195 -3045 2210 -3025
rect 2160 -3060 2210 -3045
rect -130 -3255 -90 -3240
rect -130 -3275 -120 -3255
rect -100 -3275 -90 -3255
rect -130 -3305 -90 -3275
rect -130 -3325 -120 -3305
rect -100 -3325 -90 -3305
rect -130 -3355 -90 -3325
rect -130 -3375 -120 -3355
rect -100 -3375 -90 -3355
rect -130 -3405 -90 -3375
rect -130 -3425 -120 -3405
rect -100 -3425 -90 -3405
rect -130 -3440 -90 -3425
rect -75 -3255 -35 -3240
rect -75 -3275 -65 -3255
rect -45 -3275 -35 -3255
rect -75 -3305 -35 -3275
rect -75 -3325 -65 -3305
rect -45 -3325 -35 -3305
rect -75 -3355 -35 -3325
rect -75 -3375 -65 -3355
rect -45 -3375 -35 -3355
rect -75 -3405 -35 -3375
rect -75 -3425 -65 -3405
rect -45 -3425 -35 -3405
rect -75 -3440 -35 -3425
rect -20 -3255 20 -3240
rect -20 -3275 -10 -3255
rect 10 -3275 20 -3255
rect -20 -3305 20 -3275
rect -20 -3325 -10 -3305
rect 10 -3325 20 -3305
rect -20 -3355 20 -3325
rect -20 -3375 -10 -3355
rect 10 -3375 20 -3355
rect -20 -3405 20 -3375
rect -20 -3425 -10 -3405
rect 10 -3425 20 -3405
rect -20 -3440 20 -3425
rect 130 -3255 170 -3240
rect 130 -3275 140 -3255
rect 160 -3275 170 -3255
rect 130 -3305 170 -3275
rect 130 -3325 140 -3305
rect 160 -3325 170 -3305
rect 130 -3355 170 -3325
rect 130 -3375 140 -3355
rect 160 -3375 170 -3355
rect 130 -3405 170 -3375
rect 130 -3425 140 -3405
rect 160 -3425 170 -3405
rect 130 -3440 170 -3425
rect 185 -3255 225 -3240
rect 185 -3275 195 -3255
rect 215 -3275 225 -3255
rect 185 -3305 225 -3275
rect 185 -3325 195 -3305
rect 215 -3325 225 -3305
rect 185 -3355 225 -3325
rect 185 -3375 195 -3355
rect 215 -3375 225 -3355
rect 185 -3405 225 -3375
rect 185 -3425 195 -3405
rect 215 -3425 225 -3405
rect 185 -3440 225 -3425
rect 240 -3255 280 -3240
rect 240 -3275 250 -3255
rect 270 -3275 280 -3255
rect 240 -3305 280 -3275
rect 240 -3325 250 -3305
rect 270 -3325 280 -3305
rect 240 -3355 280 -3325
rect 240 -3375 250 -3355
rect 270 -3375 280 -3355
rect 240 -3405 280 -3375
rect 240 -3425 250 -3405
rect 270 -3425 280 -3405
rect 240 -3440 280 -3425
rect 320 -3255 360 -3240
rect 320 -3275 330 -3255
rect 350 -3275 360 -3255
rect 320 -3305 360 -3275
rect 320 -3325 330 -3305
rect 350 -3325 360 -3305
rect 320 -3355 360 -3325
rect 320 -3375 330 -3355
rect 350 -3375 360 -3355
rect 320 -3405 360 -3375
rect 320 -3425 330 -3405
rect 350 -3425 360 -3405
rect 320 -3440 360 -3425
rect 375 -3255 415 -3240
rect 375 -3275 385 -3255
rect 405 -3275 415 -3255
rect 375 -3305 415 -3275
rect 375 -3325 385 -3305
rect 405 -3325 415 -3305
rect 375 -3355 415 -3325
rect 375 -3375 385 -3355
rect 405 -3375 415 -3355
rect 375 -3405 415 -3375
rect 375 -3425 385 -3405
rect 405 -3425 415 -3405
rect 375 -3440 415 -3425
rect 430 -3255 470 -3240
rect 430 -3275 440 -3255
rect 460 -3275 470 -3255
rect 430 -3305 470 -3275
rect 430 -3325 440 -3305
rect 460 -3325 470 -3305
rect 430 -3355 470 -3325
rect 430 -3375 440 -3355
rect 460 -3375 470 -3355
rect 430 -3405 470 -3375
rect 430 -3425 440 -3405
rect 460 -3425 470 -3405
rect 430 -3440 470 -3425
rect 580 -3255 620 -3240
rect 580 -3275 590 -3255
rect 610 -3275 620 -3255
rect 580 -3305 620 -3275
rect 580 -3325 590 -3305
rect 610 -3325 620 -3305
rect 580 -3355 620 -3325
rect 580 -3375 590 -3355
rect 610 -3375 620 -3355
rect 580 -3405 620 -3375
rect 580 -3425 590 -3405
rect 610 -3425 620 -3405
rect 580 -3440 620 -3425
rect 635 -3255 675 -3240
rect 635 -3275 645 -3255
rect 665 -3275 675 -3255
rect 635 -3305 675 -3275
rect 635 -3325 645 -3305
rect 665 -3325 675 -3305
rect 635 -3355 675 -3325
rect 635 -3375 645 -3355
rect 665 -3375 675 -3355
rect 635 -3405 675 -3375
rect 635 -3425 645 -3405
rect 665 -3425 675 -3405
rect 635 -3440 675 -3425
rect 690 -3255 730 -3240
rect 690 -3275 700 -3255
rect 720 -3275 730 -3255
rect 690 -3305 730 -3275
rect 690 -3325 700 -3305
rect 720 -3325 730 -3305
rect 690 -3355 730 -3325
rect 690 -3375 700 -3355
rect 720 -3375 730 -3355
rect 690 -3405 730 -3375
rect 690 -3425 700 -3405
rect 720 -3425 730 -3405
rect 690 -3440 730 -3425
rect 835 -3255 875 -3240
rect 835 -3275 845 -3255
rect 865 -3275 875 -3255
rect 835 -3305 875 -3275
rect 835 -3325 845 -3305
rect 865 -3325 875 -3305
rect 835 -3355 875 -3325
rect 835 -3375 845 -3355
rect 865 -3375 875 -3355
rect 835 -3405 875 -3375
rect 835 -3425 845 -3405
rect 865 -3425 875 -3405
rect 835 -3440 875 -3425
rect 890 -3255 930 -3240
rect 890 -3275 900 -3255
rect 920 -3275 930 -3255
rect 890 -3305 930 -3275
rect 890 -3325 900 -3305
rect 920 -3325 930 -3305
rect 890 -3355 930 -3325
rect 890 -3375 900 -3355
rect 920 -3375 930 -3355
rect 890 -3405 930 -3375
rect 890 -3425 900 -3405
rect 920 -3425 930 -3405
rect 890 -3440 930 -3425
rect 1000 -3255 1040 -3240
rect 1000 -3275 1010 -3255
rect 1030 -3275 1040 -3255
rect 1000 -3305 1040 -3275
rect 1000 -3325 1010 -3305
rect 1030 -3325 1040 -3305
rect 1000 -3355 1040 -3325
rect 1000 -3375 1010 -3355
rect 1030 -3375 1040 -3355
rect 1000 -3405 1040 -3375
rect 1000 -3425 1010 -3405
rect 1030 -3425 1040 -3405
rect 1000 -3440 1040 -3425
rect 1055 -3255 1095 -3240
rect 1055 -3275 1065 -3255
rect 1085 -3275 1095 -3255
rect 1055 -3305 1095 -3275
rect 1055 -3325 1065 -3305
rect 1085 -3325 1095 -3305
rect 1055 -3355 1095 -3325
rect 1055 -3375 1065 -3355
rect 1085 -3375 1095 -3355
rect 1055 -3405 1095 -3375
rect 1055 -3425 1065 -3405
rect 1085 -3425 1095 -3405
rect 1055 -3440 1095 -3425
rect 1165 -3255 1205 -3240
rect 1165 -3275 1175 -3255
rect 1195 -3275 1205 -3255
rect 1165 -3305 1205 -3275
rect 1165 -3325 1175 -3305
rect 1195 -3325 1205 -3305
rect 1165 -3355 1205 -3325
rect 1165 -3375 1175 -3355
rect 1195 -3375 1205 -3355
rect 1165 -3405 1205 -3375
rect 1165 -3425 1175 -3405
rect 1195 -3425 1205 -3405
rect 1165 -3440 1205 -3425
rect 1220 -3255 1260 -3240
rect 1220 -3275 1230 -3255
rect 1250 -3275 1260 -3255
rect 1220 -3305 1260 -3275
rect 1220 -3325 1230 -3305
rect 1250 -3325 1260 -3305
rect 1220 -3355 1260 -3325
rect 1220 -3375 1230 -3355
rect 1250 -3375 1260 -3355
rect 1220 -3405 1260 -3375
rect 1220 -3425 1230 -3405
rect 1250 -3425 1260 -3405
rect 1220 -3440 1260 -3425
rect 1515 -3255 1565 -3240
rect 1515 -3275 1530 -3255
rect 1550 -3275 1565 -3255
rect 1515 -3305 1565 -3275
rect 1515 -3325 1530 -3305
rect 1550 -3325 1565 -3305
rect 1515 -3355 1565 -3325
rect 1515 -3375 1530 -3355
rect 1550 -3375 1565 -3355
rect 1515 -3405 1565 -3375
rect 1515 -3425 1530 -3405
rect 1550 -3425 1565 -3405
rect 1515 -3440 1565 -3425
rect 1580 -3255 1630 -3240
rect 1580 -3275 1595 -3255
rect 1615 -3275 1630 -3255
rect 1580 -3305 1630 -3275
rect 1580 -3325 1595 -3305
rect 1615 -3325 1630 -3305
rect 1580 -3355 1630 -3325
rect 1580 -3375 1595 -3355
rect 1615 -3375 1630 -3355
rect 1580 -3405 1630 -3375
rect 1580 -3425 1595 -3405
rect 1615 -3425 1630 -3405
rect 1580 -3440 1630 -3425
rect 1660 -3255 1710 -3240
rect 1660 -3275 1675 -3255
rect 1695 -3275 1710 -3255
rect 1660 -3305 1710 -3275
rect 1660 -3325 1675 -3305
rect 1695 -3325 1710 -3305
rect 1660 -3355 1710 -3325
rect 1660 -3375 1675 -3355
rect 1695 -3375 1710 -3355
rect 1660 -3405 1710 -3375
rect 1660 -3425 1675 -3405
rect 1695 -3425 1710 -3405
rect 1660 -3440 1710 -3425
rect 1725 -3255 1775 -3240
rect 1725 -3275 1740 -3255
rect 1760 -3275 1775 -3255
rect 1725 -3305 1775 -3275
rect 1725 -3325 1740 -3305
rect 1760 -3325 1775 -3305
rect 1725 -3355 1775 -3325
rect 1725 -3375 1740 -3355
rect 1760 -3375 1775 -3355
rect 1725 -3405 1775 -3375
rect 1725 -3425 1740 -3405
rect 1760 -3425 1775 -3405
rect 1725 -3440 1775 -3425
rect 1805 -3255 1855 -3240
rect 1805 -3275 1820 -3255
rect 1840 -3275 1855 -3255
rect 1805 -3305 1855 -3275
rect 1805 -3325 1820 -3305
rect 1840 -3325 1855 -3305
rect 1805 -3355 1855 -3325
rect 1805 -3375 1820 -3355
rect 1840 -3375 1855 -3355
rect 1805 -3405 1855 -3375
rect 1805 -3425 1820 -3405
rect 1840 -3425 1855 -3405
rect 1805 -3440 1855 -3425
rect 1870 -3255 1920 -3240
rect 1870 -3275 1885 -3255
rect 1905 -3275 1920 -3255
rect 1870 -3305 1920 -3275
rect 1870 -3325 1885 -3305
rect 1905 -3325 1920 -3305
rect 1870 -3355 1920 -3325
rect 1870 -3375 1885 -3355
rect 1905 -3375 1920 -3355
rect 1870 -3405 1920 -3375
rect 1870 -3425 1885 -3405
rect 1905 -3425 1920 -3405
rect 1870 -3440 1920 -3425
rect 1950 -3255 2000 -3240
rect 1950 -3275 1965 -3255
rect 1985 -3275 2000 -3255
rect 1950 -3305 2000 -3275
rect 1950 -3325 1965 -3305
rect 1985 -3325 2000 -3305
rect 1950 -3355 2000 -3325
rect 1950 -3375 1965 -3355
rect 1985 -3375 2000 -3355
rect 1950 -3405 2000 -3375
rect 1950 -3425 1965 -3405
rect 1985 -3425 2000 -3405
rect 1950 -3440 2000 -3425
rect 2015 -3255 2065 -3240
rect 2015 -3275 2030 -3255
rect 2050 -3275 2065 -3255
rect 2015 -3305 2065 -3275
rect 2015 -3325 2030 -3305
rect 2050 -3325 2065 -3305
rect 2015 -3355 2065 -3325
rect 2015 -3375 2030 -3355
rect 2050 -3375 2065 -3355
rect 2015 -3405 2065 -3375
rect 2015 -3425 2030 -3405
rect 2050 -3425 2065 -3405
rect 2015 -3440 2065 -3425
rect 2815 -3730 2865 -3715
rect 2815 -3900 2830 -3730
rect 2850 -3900 2865 -3730
rect 2815 -3915 2865 -3900
rect 2880 -3730 2930 -3715
rect 2880 -3900 2895 -3730
rect 2915 -3900 2930 -3730
rect 2880 -3915 2930 -3900
rect 2960 -3730 3010 -3715
rect 2960 -3900 2975 -3730
rect 2995 -3900 3010 -3730
rect 2960 -3915 3010 -3900
rect 3025 -3730 3075 -3715
rect 3025 -3900 3040 -3730
rect 3060 -3900 3075 -3730
rect 3025 -3915 3075 -3900
rect 3105 -3730 3155 -3715
rect 3105 -3900 3120 -3730
rect 3140 -3900 3155 -3730
rect 3105 -3915 3155 -3900
rect 3170 -3730 3220 -3715
rect 3170 -3900 3185 -3730
rect 3205 -3900 3220 -3730
rect 3170 -3915 3220 -3900
rect 3250 -3730 3300 -3715
rect 3250 -3900 3265 -3730
rect 3285 -3900 3300 -3730
rect 3250 -3915 3300 -3900
rect 3315 -3730 3365 -3715
rect 3315 -3900 3330 -3730
rect 3350 -3900 3365 -3730
rect 3315 -3915 3365 -3900
rect 3395 -3730 3445 -3715
rect 3395 -3900 3410 -3730
rect 3430 -3900 3445 -3730
rect 3395 -3915 3445 -3900
rect 3460 -3730 3510 -3715
rect 3460 -3900 3475 -3730
rect 3495 -3900 3510 -3730
rect 3460 -3915 3510 -3900
rect 3540 -3730 3590 -3715
rect 3540 -3900 3555 -3730
rect 3575 -3900 3590 -3730
rect 3540 -3915 3590 -3900
rect 3605 -3730 3655 -3715
rect 3605 -3900 3620 -3730
rect 3640 -3900 3655 -3730
rect 3605 -3915 3655 -3900
rect 3685 -3730 3735 -3715
rect 3685 -3900 3700 -3730
rect 3720 -3900 3735 -3730
rect 3685 -3915 3735 -3900
rect 3750 -3730 3800 -3715
rect 3750 -3900 3765 -3730
rect 3785 -3900 3800 -3730
rect 3750 -3915 3800 -3900
rect 3830 -3730 3880 -3715
rect 3830 -3900 3845 -3730
rect 3865 -3900 3880 -3730
rect 3830 -3915 3880 -3900
rect 3895 -3730 3945 -3715
rect 3895 -3900 3910 -3730
rect 3930 -3900 3945 -3730
rect 3895 -3915 3945 -3900
rect 3975 -3730 4025 -3715
rect 3975 -3900 3990 -3730
rect 4010 -3900 4025 -3730
rect 3975 -3915 4025 -3900
rect 4040 -3730 4090 -3715
rect 4040 -3900 4055 -3730
rect 4075 -3900 4090 -3730
rect 4040 -3915 4090 -3900
rect 1515 -5345 1565 -5330
rect 1515 -5365 1530 -5345
rect 1550 -5365 1565 -5345
rect 1515 -5395 1565 -5365
rect 1515 -5415 1530 -5395
rect 1550 -5415 1565 -5395
rect 1515 -5445 1565 -5415
rect 1515 -5465 1530 -5445
rect 1550 -5465 1565 -5445
rect 1515 -5495 1565 -5465
rect 1515 -5515 1530 -5495
rect 1550 -5515 1565 -5495
rect 1515 -5530 1565 -5515
rect 1580 -5345 1630 -5330
rect 1580 -5365 1595 -5345
rect 1615 -5365 1630 -5345
rect 1580 -5395 1630 -5365
rect 1580 -5415 1595 -5395
rect 1615 -5415 1630 -5395
rect 1580 -5445 1630 -5415
rect 1580 -5465 1595 -5445
rect 1615 -5465 1630 -5445
rect 1580 -5495 1630 -5465
rect 1580 -5515 1595 -5495
rect 1615 -5515 1630 -5495
rect 1580 -5530 1630 -5515
rect 1660 -5345 1710 -5330
rect 1660 -5365 1675 -5345
rect 1695 -5365 1710 -5345
rect 1660 -5395 1710 -5365
rect 1660 -5415 1675 -5395
rect 1695 -5415 1710 -5395
rect 1660 -5445 1710 -5415
rect 1660 -5465 1675 -5445
rect 1695 -5465 1710 -5445
rect 1660 -5495 1710 -5465
rect 1660 -5515 1675 -5495
rect 1695 -5515 1710 -5495
rect 1660 -5530 1710 -5515
rect 1725 -5345 1775 -5330
rect 1725 -5365 1740 -5345
rect 1760 -5365 1775 -5345
rect 1725 -5395 1775 -5365
rect 1725 -5415 1740 -5395
rect 1760 -5415 1775 -5395
rect 1725 -5445 1775 -5415
rect 1725 -5465 1740 -5445
rect 1760 -5465 1775 -5445
rect 1725 -5495 1775 -5465
rect 1725 -5515 1740 -5495
rect 1760 -5515 1775 -5495
rect 1725 -5530 1775 -5515
rect 1805 -5345 1855 -5330
rect 1805 -5365 1820 -5345
rect 1840 -5365 1855 -5345
rect 1805 -5395 1855 -5365
rect 1805 -5415 1820 -5395
rect 1840 -5415 1855 -5395
rect 1805 -5445 1855 -5415
rect 1805 -5465 1820 -5445
rect 1840 -5465 1855 -5445
rect 1805 -5495 1855 -5465
rect 1805 -5515 1820 -5495
rect 1840 -5515 1855 -5495
rect 1805 -5530 1855 -5515
rect 1870 -5345 1920 -5330
rect 1870 -5365 1885 -5345
rect 1905 -5365 1920 -5345
rect 1870 -5395 1920 -5365
rect 1870 -5415 1885 -5395
rect 1905 -5415 1920 -5395
rect 1870 -5445 1920 -5415
rect 1870 -5465 1885 -5445
rect 1905 -5465 1920 -5445
rect 1870 -5495 1920 -5465
rect 1870 -5515 1885 -5495
rect 1905 -5515 1920 -5495
rect 1870 -5530 1920 -5515
rect 1950 -5345 2000 -5330
rect 1950 -5365 1965 -5345
rect 1985 -5365 2000 -5345
rect 1950 -5395 2000 -5365
rect 1950 -5415 1965 -5395
rect 1985 -5415 2000 -5395
rect 1950 -5445 2000 -5415
rect 1950 -5465 1965 -5445
rect 1985 -5465 2000 -5445
rect 1950 -5495 2000 -5465
rect 1950 -5515 1965 -5495
rect 1985 -5515 2000 -5495
rect 1950 -5530 2000 -5515
rect 2015 -5345 2065 -5330
rect 2015 -5365 2030 -5345
rect 2050 -5365 2065 -5345
rect 2015 -5395 2065 -5365
rect 2015 -5415 2030 -5395
rect 2050 -5415 2065 -5395
rect 2015 -5445 2065 -5415
rect 2015 -5465 2030 -5445
rect 2050 -5465 2065 -5445
rect 2015 -5495 2065 -5465
rect 2015 -5515 2030 -5495
rect 2050 -5515 2065 -5495
rect 2015 -5530 2065 -5515
rect 1515 -5735 1565 -5720
rect 1515 -5755 1530 -5735
rect 1550 -5755 1565 -5735
rect 1515 -5785 1565 -5755
rect 1515 -5805 1530 -5785
rect 1550 -5805 1565 -5785
rect 1515 -5835 1565 -5805
rect 1515 -5855 1530 -5835
rect 1550 -5855 1565 -5835
rect 1515 -5885 1565 -5855
rect 1515 -5905 1530 -5885
rect 1550 -5905 1565 -5885
rect 1515 -5920 1565 -5905
rect 1580 -5735 1630 -5720
rect 1580 -5755 1595 -5735
rect 1615 -5755 1630 -5735
rect 1580 -5785 1630 -5755
rect 1580 -5805 1595 -5785
rect 1615 -5805 1630 -5785
rect 1580 -5835 1630 -5805
rect 1580 -5855 1595 -5835
rect 1615 -5855 1630 -5835
rect 1580 -5885 1630 -5855
rect 1580 -5905 1595 -5885
rect 1615 -5905 1630 -5885
rect 1580 -5920 1630 -5905
rect 1660 -5735 1710 -5720
rect 1660 -5755 1675 -5735
rect 1695 -5755 1710 -5735
rect 1660 -5785 1710 -5755
rect 1660 -5805 1675 -5785
rect 1695 -5805 1710 -5785
rect 1660 -5835 1710 -5805
rect 1660 -5855 1675 -5835
rect 1695 -5855 1710 -5835
rect 1660 -5885 1710 -5855
rect 1660 -5905 1675 -5885
rect 1695 -5905 1710 -5885
rect 1660 -5920 1710 -5905
rect 1725 -5735 1775 -5720
rect 1725 -5755 1740 -5735
rect 1760 -5755 1775 -5735
rect 1725 -5785 1775 -5755
rect 1725 -5805 1740 -5785
rect 1760 -5805 1775 -5785
rect 1725 -5835 1775 -5805
rect 1725 -5855 1740 -5835
rect 1760 -5855 1775 -5835
rect 1725 -5885 1775 -5855
rect 1725 -5905 1740 -5885
rect 1760 -5905 1775 -5885
rect 1725 -5920 1775 -5905
rect 1805 -5735 1855 -5720
rect 1805 -5755 1820 -5735
rect 1840 -5755 1855 -5735
rect 1805 -5785 1855 -5755
rect 1805 -5805 1820 -5785
rect 1840 -5805 1855 -5785
rect 1805 -5835 1855 -5805
rect 1805 -5855 1820 -5835
rect 1840 -5855 1855 -5835
rect 1805 -5885 1855 -5855
rect 1805 -5905 1820 -5885
rect 1840 -5905 1855 -5885
rect 1805 -5920 1855 -5905
rect 1870 -5735 1920 -5720
rect 1870 -5755 1885 -5735
rect 1905 -5755 1920 -5735
rect 1870 -5785 1920 -5755
rect 1870 -5805 1885 -5785
rect 1905 -5805 1920 -5785
rect 1870 -5835 1920 -5805
rect 1870 -5855 1885 -5835
rect 1905 -5855 1920 -5835
rect 1870 -5885 1920 -5855
rect 1870 -5905 1885 -5885
rect 1905 -5905 1920 -5885
rect 1870 -5920 1920 -5905
rect 1950 -5735 2000 -5720
rect 1950 -5755 1965 -5735
rect 1985 -5755 2000 -5735
rect 1950 -5785 2000 -5755
rect 1950 -5805 1965 -5785
rect 1985 -5805 2000 -5785
rect 1950 -5835 2000 -5805
rect 1950 -5855 1965 -5835
rect 1985 -5855 2000 -5835
rect 1950 -5885 2000 -5855
rect 1950 -5905 1965 -5885
rect 1985 -5905 2000 -5885
rect 1950 -5920 2000 -5905
rect 2015 -5735 2065 -5720
rect 2015 -5755 2030 -5735
rect 2050 -5755 2065 -5735
rect 2015 -5785 2065 -5755
rect 2015 -5805 2030 -5785
rect 2050 -5805 2065 -5785
rect 2015 -5835 2065 -5805
rect 2015 -5855 2030 -5835
rect 2050 -5855 2065 -5835
rect 2015 -5885 2065 -5855
rect 2015 -5905 2030 -5885
rect 2050 -5905 2065 -5885
rect 2015 -5920 2065 -5905
rect 2095 -5735 2145 -5720
rect 2095 -5755 2110 -5735
rect 2130 -5755 2145 -5735
rect 2095 -5785 2145 -5755
rect 2095 -5805 2110 -5785
rect 2130 -5805 2145 -5785
rect 2095 -5835 2145 -5805
rect 2095 -5855 2110 -5835
rect 2130 -5855 2145 -5835
rect 2095 -5885 2145 -5855
rect 2095 -5905 2110 -5885
rect 2130 -5905 2145 -5885
rect 2095 -5920 2145 -5905
rect 2160 -5735 2210 -5720
rect 2160 -5755 2175 -5735
rect 2195 -5755 2210 -5735
rect 2160 -5785 2210 -5755
rect 2160 -5805 2175 -5785
rect 2195 -5805 2210 -5785
rect 2160 -5835 2210 -5805
rect 2160 -5855 2175 -5835
rect 2195 -5855 2210 -5835
rect 2160 -5885 2210 -5855
rect 2160 -5905 2175 -5885
rect 2195 -5905 2210 -5885
rect 2160 -5920 2210 -5905
<< ndiffc >>
rect -30 15 -10 35
rect 25 15 45 35
rect 80 15 100 35
rect 230 15 250 35
rect 285 15 305 35
rect 340 15 360 35
rect 410 15 430 35
rect 465 15 485 35
rect 520 15 540 35
rect 670 15 690 35
rect 725 15 745 35
rect 780 15 800 35
rect 850 15 870 35
rect 905 15 925 35
rect 960 15 980 35
rect 1110 15 1130 35
rect 1165 15 1185 35
rect 1220 15 1240 35
rect 1300 15 1320 35
rect 1355 15 1375 35
rect 1410 15 1430 35
rect 1560 15 1580 35
rect 1615 15 1635 35
rect 1670 15 1690 35
rect 1740 15 1760 35
rect 1795 15 1815 35
rect 1850 15 1870 35
rect 1920 15 1940 35
rect 1975 15 1995 35
rect 2045 15 2065 35
rect 2100 15 2120 35
rect 2170 15 2190 35
rect 2225 15 2245 35
rect 2295 15 2315 35
rect 2350 15 2370 35
rect 2420 15 2440 35
rect 2475 15 2495 35
rect 2830 -130 2850 -60
rect 2895 -130 2915 -60
rect 2975 -130 2995 -60
rect 3040 -130 3060 -60
rect 3120 -130 3140 -60
rect 3185 -130 3205 -60
rect 3265 -130 3285 -60
rect 3330 -130 3350 -60
rect 3410 -130 3430 -60
rect 3475 -130 3495 -60
rect 3555 -130 3575 -60
rect 3620 -130 3640 -60
rect 3700 -130 3720 -60
rect 3765 -130 3785 -60
rect 3845 -130 3865 -60
rect 3910 -130 3930 -60
rect 3990 -130 4010 -60
rect 4055 -130 4075 -60
rect -30 -1235 -10 -1215
rect 25 -1235 45 -1215
rect 80 -1235 100 -1215
rect 230 -1235 250 -1215
rect 285 -1235 305 -1215
rect 340 -1235 360 -1215
rect 410 -1235 430 -1215
rect 465 -1235 485 -1215
rect 520 -1235 540 -1215
rect 670 -1235 690 -1215
rect 725 -1235 745 -1215
rect 780 -1235 800 -1215
rect 910 -1235 930 -1215
rect 965 -1235 985 -1215
rect 1020 -1235 1040 -1215
rect 1090 -1235 1110 -1215
rect 1145 -1235 1165 -1215
rect 1215 -1235 1235 -1215
rect 1270 -1235 1290 -1215
rect -30 -1985 -10 -1965
rect 25 -1985 45 -1965
rect 80 -1985 100 -1965
rect 230 -1985 250 -1965
rect 285 -1985 305 -1965
rect 340 -1985 360 -1965
rect 410 -1985 430 -1965
rect 465 -1985 485 -1965
rect 520 -1985 540 -1965
rect 670 -1985 690 -1965
rect 725 -1985 745 -1965
rect 780 -1985 800 -1965
rect 960 -1985 980 -1965
rect 1015 -1985 1035 -1965
rect 1085 -1985 1105 -1965
rect 1140 -1985 1160 -1965
rect 1210 -1985 1230 -1965
rect 1265 -1985 1285 -1965
rect -120 -2735 -100 -2665
rect -65 -2735 -45 -2665
rect -10 -2735 10 -2665
rect 140 -2735 160 -2665
rect 195 -2735 215 -2665
rect 250 -2735 270 -2665
rect 330 -2735 350 -2665
rect 385 -2735 405 -2665
rect 440 -2735 460 -2665
rect 590 -2735 610 -2665
rect 645 -2735 665 -2665
rect 700 -2735 720 -2665
rect 795 -2735 815 -2665
rect 850 -2735 870 -2665
rect 905 -2735 925 -2665
rect 1015 -2735 1035 -2665
rect 1070 -2735 1090 -2665
rect 1180 -2735 1200 -2665
rect 1235 -2735 1255 -2665
rect 1530 -2685 1550 -2665
rect 1530 -2735 1550 -2715
rect 1595 -2685 1615 -2665
rect 1595 -2735 1615 -2715
rect 1675 -2685 1695 -2665
rect 1675 -2735 1695 -2715
rect 1740 -2685 1760 -2665
rect 1740 -2735 1760 -2715
rect 1820 -2685 1840 -2665
rect 1820 -2735 1840 -2715
rect 1885 -2685 1905 -2665
rect 1885 -2735 1905 -2715
rect 1965 -2685 1985 -2665
rect 1965 -2735 1985 -2715
rect 2030 -2685 2050 -2665
rect 2030 -2735 2050 -2715
rect -120 -3585 -100 -3565
rect -120 -3635 -100 -3615
rect -65 -3585 -45 -3565
rect -65 -3635 -45 -3615
rect -10 -3585 10 -3565
rect -10 -3635 10 -3615
rect 140 -3585 160 -3565
rect 140 -3635 160 -3615
rect 195 -3585 215 -3565
rect 195 -3635 215 -3615
rect 250 -3585 270 -3565
rect 330 -3585 350 -3565
rect 250 -3635 270 -3615
rect 330 -3635 350 -3615
rect 385 -3585 405 -3565
rect 385 -3635 405 -3615
rect 440 -3585 460 -3565
rect 440 -3635 460 -3615
rect 590 -3585 610 -3565
rect 590 -3635 610 -3615
rect 645 -3585 665 -3565
rect 645 -3635 665 -3615
rect 700 -3585 720 -3565
rect 700 -3635 720 -3615
rect 845 -3585 865 -3565
rect 845 -3635 865 -3615
rect 900 -3585 920 -3565
rect 900 -3635 920 -3615
rect 1010 -3585 1030 -3565
rect 1010 -3635 1030 -3615
rect 1065 -3585 1085 -3565
rect 1065 -3635 1085 -3615
rect 1175 -3585 1195 -3565
rect 1175 -3635 1195 -3615
rect 1230 -3585 1250 -3565
rect 1230 -3635 1250 -3615
rect 1530 -3585 1550 -3565
rect 1530 -3635 1550 -3615
rect 1595 -3585 1615 -3565
rect 1595 -3635 1615 -3615
rect 1675 -3585 1695 -3565
rect 1675 -3635 1695 -3615
rect 1740 -3585 1760 -3565
rect 1740 -3635 1760 -3615
rect 1820 -3585 1840 -3565
rect 1820 -3635 1840 -3615
rect 1885 -3585 1905 -3565
rect 1885 -3635 1905 -3615
rect 1965 -3585 1985 -3565
rect 1965 -3635 1985 -3615
rect 2030 -3585 2050 -3565
rect 2030 -3635 2050 -3615
rect 2110 -3585 2130 -3565
rect 2110 -3635 2130 -3615
rect 2175 -3585 2195 -3565
rect 2175 -3635 2195 -3615
rect 2830 -4130 2850 -4060
rect 2895 -4130 2915 -4060
rect 2975 -4130 2995 -4060
rect 3040 -4130 3060 -4060
rect 3120 -4130 3140 -4060
rect 3185 -4130 3205 -4060
rect 3265 -4130 3285 -4060
rect 3330 -4130 3350 -4060
rect 3410 -4130 3430 -4060
rect 3475 -4130 3495 -4060
rect 3555 -4130 3575 -4060
rect 3620 -4130 3640 -4060
rect 3700 -4130 3720 -4060
rect 3765 -4130 3785 -4060
rect 3845 -4130 3865 -4060
rect 3910 -4130 3930 -4060
rect 3990 -4130 4010 -4060
rect 4055 -4130 4075 -4060
rect 1530 -5135 1550 -5115
rect 1530 -5185 1550 -5165
rect 1595 -5135 1615 -5115
rect 1595 -5185 1615 -5165
rect 1675 -5135 1695 -5115
rect 1675 -5185 1695 -5165
rect 1740 -5135 1760 -5115
rect 1740 -5185 1760 -5165
rect 1820 -5135 1840 -5115
rect 1820 -5185 1840 -5165
rect 1885 -5135 1905 -5115
rect 1885 -5185 1905 -5165
rect 1965 -5135 1985 -5115
rect 1965 -5185 1985 -5165
rect 2030 -5135 2050 -5115
rect 2030 -5185 2050 -5165
rect 1530 -6085 1550 -6065
rect 1530 -6135 1550 -6115
rect 1595 -6085 1615 -6065
rect 1595 -6135 1615 -6115
rect 1675 -6085 1695 -6065
rect 1675 -6135 1695 -6115
rect 1740 -6085 1760 -6065
rect 1740 -6135 1760 -6115
rect 1820 -6085 1840 -6065
rect 1820 -6135 1840 -6115
rect 1885 -6085 1905 -6065
rect 1885 -6135 1905 -6115
rect 1965 -6085 1985 -6065
rect 1965 -6135 1985 -6115
rect 2030 -6085 2050 -6065
rect 2030 -6135 2050 -6115
rect 2110 -6085 2130 -6065
rect 2110 -6135 2130 -6115
rect 2175 -6085 2195 -6065
rect 2175 -6135 2195 -6115
<< pdiffc >>
rect -30 175 -10 245
rect 25 175 45 245
rect 80 175 100 245
rect 230 175 250 245
rect 285 175 305 245
rect 340 175 360 245
rect 410 175 430 245
rect 465 175 485 245
rect 520 175 540 245
rect 670 175 690 245
rect 725 175 745 245
rect 780 175 800 245
rect 850 175 870 245
rect 905 175 925 245
rect 960 175 980 245
rect 1110 175 1130 245
rect 1165 175 1185 245
rect 1220 175 1240 245
rect 1300 175 1320 245
rect 1355 175 1375 245
rect 1410 175 1430 245
rect 1560 175 1580 245
rect 1615 175 1635 245
rect 1670 175 1690 245
rect 1740 175 1760 245
rect 1795 175 1815 245
rect 1850 175 1870 245
rect 1920 175 1940 245
rect 1975 175 1995 245
rect 2045 175 2065 245
rect 2100 175 2120 245
rect 2170 175 2190 245
rect 2225 175 2245 245
rect 2295 175 2315 245
rect 2350 175 2370 245
rect 2420 175 2440 245
rect 2475 175 2495 245
rect 2830 100 2850 270
rect 2895 100 2915 270
rect 2975 100 2995 270
rect 3040 100 3060 270
rect 3120 100 3140 270
rect 3185 100 3205 270
rect 3265 100 3285 270
rect 3330 100 3350 270
rect 3410 100 3430 270
rect 3475 100 3495 270
rect 3555 100 3575 270
rect 3620 100 3640 270
rect 3700 100 3720 270
rect 3765 100 3785 270
rect 3845 100 3865 270
rect 3910 100 3930 270
rect 3990 100 4010 270
rect 4055 100 4075 270
rect -30 -1445 -10 -1375
rect 25 -1445 45 -1375
rect 80 -1445 100 -1375
rect 230 -1445 250 -1375
rect 285 -1445 305 -1375
rect 340 -1445 360 -1375
rect 410 -1445 430 -1375
rect 465 -1445 485 -1375
rect 520 -1445 540 -1375
rect 670 -1445 690 -1375
rect 725 -1445 745 -1375
rect 780 -1445 800 -1375
rect 910 -1445 930 -1375
rect 965 -1445 985 -1375
rect 1020 -1445 1040 -1375
rect 1090 -1445 1110 -1375
rect 1145 -1445 1165 -1375
rect 1215 -1445 1235 -1375
rect 1270 -1445 1290 -1375
rect -30 -1825 -10 -1755
rect 25 -1825 45 -1755
rect 80 -1825 100 -1755
rect 230 -1825 250 -1755
rect 285 -1825 305 -1755
rect 340 -1825 360 -1755
rect 410 -1825 430 -1755
rect 465 -1825 485 -1755
rect 520 -1825 540 -1755
rect 670 -1825 690 -1755
rect 725 -1825 745 -1755
rect 780 -1825 800 -1755
rect 960 -1825 980 -1755
rect 1015 -1825 1035 -1755
rect 1085 -1825 1105 -1755
rect 1140 -1825 1160 -1755
rect 1210 -1825 1230 -1755
rect 1265 -1825 1285 -1755
rect -120 -2895 -100 -2875
rect -120 -2945 -100 -2925
rect -120 -2995 -100 -2975
rect -120 -3045 -100 -3025
rect -65 -2895 -45 -2875
rect -65 -2945 -45 -2925
rect -65 -2995 -45 -2975
rect -65 -3045 -45 -3025
rect -10 -2895 10 -2875
rect -10 -2945 10 -2925
rect -10 -2995 10 -2975
rect -10 -3045 10 -3025
rect 140 -2895 160 -2875
rect 140 -2945 160 -2925
rect 140 -2995 160 -2975
rect 140 -3045 160 -3025
rect 195 -2895 215 -2875
rect 195 -2945 215 -2925
rect 195 -2995 215 -2975
rect 195 -3045 215 -3025
rect 250 -2895 270 -2875
rect 250 -2945 270 -2925
rect 250 -2995 270 -2975
rect 250 -3045 270 -3025
rect 330 -2895 350 -2875
rect 330 -2945 350 -2925
rect 330 -2995 350 -2975
rect 330 -3045 350 -3025
rect 385 -2895 405 -2875
rect 385 -2945 405 -2925
rect 385 -2995 405 -2975
rect 385 -3045 405 -3025
rect 440 -2895 460 -2875
rect 440 -2945 460 -2925
rect 440 -2995 460 -2975
rect 440 -3045 460 -3025
rect 590 -2895 610 -2875
rect 590 -2945 610 -2925
rect 590 -2995 610 -2975
rect 590 -3045 610 -3025
rect 645 -2895 665 -2875
rect 645 -2945 665 -2925
rect 645 -2995 665 -2975
rect 645 -3045 665 -3025
rect 700 -2895 720 -2875
rect 700 -2945 720 -2925
rect 700 -2995 720 -2975
rect 700 -3045 720 -3025
rect 795 -2895 815 -2875
rect 795 -2945 815 -2925
rect 795 -2995 815 -2975
rect 795 -3045 815 -3025
rect 850 -2895 870 -2875
rect 850 -2945 870 -2925
rect 850 -2995 870 -2975
rect 850 -3045 870 -3025
rect 905 -2895 925 -2875
rect 905 -2945 925 -2925
rect 905 -2995 925 -2975
rect 905 -3045 925 -3025
rect 1015 -2895 1035 -2875
rect 1015 -2945 1035 -2925
rect 1015 -2995 1035 -2975
rect 1015 -3045 1035 -3025
rect 1070 -2895 1090 -2875
rect 1070 -2945 1090 -2925
rect 1070 -2995 1090 -2975
rect 1070 -3045 1090 -3025
rect 1180 -2895 1200 -2875
rect 1180 -2945 1200 -2925
rect 1180 -2995 1200 -2975
rect 1180 -3045 1200 -3025
rect 1235 -2895 1255 -2875
rect 1235 -2945 1255 -2925
rect 1235 -2995 1255 -2975
rect 1235 -3045 1255 -3025
rect 1530 -2895 1550 -2875
rect 1530 -2945 1550 -2925
rect 1530 -2995 1550 -2975
rect 1530 -3045 1550 -3025
rect 1595 -2895 1615 -2875
rect 1595 -2945 1615 -2925
rect 1595 -2995 1615 -2975
rect 1595 -3045 1615 -3025
rect 1675 -2895 1695 -2875
rect 1675 -2945 1695 -2925
rect 1675 -2995 1695 -2975
rect 1675 -3045 1695 -3025
rect 1740 -2895 1760 -2875
rect 1740 -2945 1760 -2925
rect 1740 -2995 1760 -2975
rect 1740 -3045 1760 -3025
rect 1820 -2895 1840 -2875
rect 1820 -2945 1840 -2925
rect 1820 -2995 1840 -2975
rect 1820 -3045 1840 -3025
rect 1885 -2895 1905 -2875
rect 1885 -2945 1905 -2925
rect 1885 -2995 1905 -2975
rect 1885 -3045 1905 -3025
rect 1965 -2895 1985 -2875
rect 1965 -2945 1985 -2925
rect 1965 -2995 1985 -2975
rect 1965 -3045 1985 -3025
rect 2030 -2895 2050 -2875
rect 2030 -2945 2050 -2925
rect 2030 -2995 2050 -2975
rect 2030 -3045 2050 -3025
rect 2110 -2895 2130 -2875
rect 2110 -2945 2130 -2925
rect 2110 -2995 2130 -2975
rect 2110 -3045 2130 -3025
rect 2175 -2895 2195 -2875
rect 2175 -2945 2195 -2925
rect 2175 -2995 2195 -2975
rect 2175 -3045 2195 -3025
rect -120 -3275 -100 -3255
rect -120 -3325 -100 -3305
rect -120 -3375 -100 -3355
rect -120 -3425 -100 -3405
rect -65 -3275 -45 -3255
rect -65 -3325 -45 -3305
rect -65 -3375 -45 -3355
rect -65 -3425 -45 -3405
rect -10 -3275 10 -3255
rect -10 -3325 10 -3305
rect -10 -3375 10 -3355
rect -10 -3425 10 -3405
rect 140 -3275 160 -3255
rect 140 -3325 160 -3305
rect 140 -3375 160 -3355
rect 140 -3425 160 -3405
rect 195 -3275 215 -3255
rect 195 -3325 215 -3305
rect 195 -3375 215 -3355
rect 195 -3425 215 -3405
rect 250 -3275 270 -3255
rect 250 -3325 270 -3305
rect 250 -3375 270 -3355
rect 250 -3425 270 -3405
rect 330 -3275 350 -3255
rect 330 -3325 350 -3305
rect 330 -3375 350 -3355
rect 330 -3425 350 -3405
rect 385 -3275 405 -3255
rect 385 -3325 405 -3305
rect 385 -3375 405 -3355
rect 385 -3425 405 -3405
rect 440 -3275 460 -3255
rect 440 -3325 460 -3305
rect 440 -3375 460 -3355
rect 440 -3425 460 -3405
rect 590 -3275 610 -3255
rect 590 -3325 610 -3305
rect 590 -3375 610 -3355
rect 590 -3425 610 -3405
rect 645 -3275 665 -3255
rect 645 -3325 665 -3305
rect 645 -3375 665 -3355
rect 645 -3425 665 -3405
rect 700 -3275 720 -3255
rect 700 -3325 720 -3305
rect 700 -3375 720 -3355
rect 700 -3425 720 -3405
rect 845 -3275 865 -3255
rect 845 -3325 865 -3305
rect 845 -3375 865 -3355
rect 845 -3425 865 -3405
rect 900 -3275 920 -3255
rect 900 -3325 920 -3305
rect 900 -3375 920 -3355
rect 900 -3425 920 -3405
rect 1010 -3275 1030 -3255
rect 1010 -3325 1030 -3305
rect 1010 -3375 1030 -3355
rect 1010 -3425 1030 -3405
rect 1065 -3275 1085 -3255
rect 1065 -3325 1085 -3305
rect 1065 -3375 1085 -3355
rect 1065 -3425 1085 -3405
rect 1175 -3275 1195 -3255
rect 1175 -3325 1195 -3305
rect 1175 -3375 1195 -3355
rect 1175 -3425 1195 -3405
rect 1230 -3275 1250 -3255
rect 1230 -3325 1250 -3305
rect 1230 -3375 1250 -3355
rect 1230 -3425 1250 -3405
rect 1530 -3275 1550 -3255
rect 1530 -3325 1550 -3305
rect 1530 -3375 1550 -3355
rect 1530 -3425 1550 -3405
rect 1595 -3275 1615 -3255
rect 1595 -3325 1615 -3305
rect 1595 -3375 1615 -3355
rect 1595 -3425 1615 -3405
rect 1675 -3275 1695 -3255
rect 1675 -3325 1695 -3305
rect 1675 -3375 1695 -3355
rect 1675 -3425 1695 -3405
rect 1740 -3275 1760 -3255
rect 1740 -3325 1760 -3305
rect 1740 -3375 1760 -3355
rect 1740 -3425 1760 -3405
rect 1820 -3275 1840 -3255
rect 1820 -3325 1840 -3305
rect 1820 -3375 1840 -3355
rect 1820 -3425 1840 -3405
rect 1885 -3275 1905 -3255
rect 1885 -3325 1905 -3305
rect 1885 -3375 1905 -3355
rect 1885 -3425 1905 -3405
rect 1965 -3275 1985 -3255
rect 1965 -3325 1985 -3305
rect 1965 -3375 1985 -3355
rect 1965 -3425 1985 -3405
rect 2030 -3275 2050 -3255
rect 2030 -3325 2050 -3305
rect 2030 -3375 2050 -3355
rect 2030 -3425 2050 -3405
rect 2830 -3900 2850 -3730
rect 2895 -3900 2915 -3730
rect 2975 -3900 2995 -3730
rect 3040 -3900 3060 -3730
rect 3120 -3900 3140 -3730
rect 3185 -3900 3205 -3730
rect 3265 -3900 3285 -3730
rect 3330 -3900 3350 -3730
rect 3410 -3900 3430 -3730
rect 3475 -3900 3495 -3730
rect 3555 -3900 3575 -3730
rect 3620 -3900 3640 -3730
rect 3700 -3900 3720 -3730
rect 3765 -3900 3785 -3730
rect 3845 -3900 3865 -3730
rect 3910 -3900 3930 -3730
rect 3990 -3900 4010 -3730
rect 4055 -3900 4075 -3730
rect 1530 -5365 1550 -5345
rect 1530 -5415 1550 -5395
rect 1530 -5465 1550 -5445
rect 1530 -5515 1550 -5495
rect 1595 -5365 1615 -5345
rect 1595 -5415 1615 -5395
rect 1595 -5465 1615 -5445
rect 1595 -5515 1615 -5495
rect 1675 -5365 1695 -5345
rect 1675 -5415 1695 -5395
rect 1675 -5465 1695 -5445
rect 1675 -5515 1695 -5495
rect 1740 -5365 1760 -5345
rect 1740 -5415 1760 -5395
rect 1740 -5465 1760 -5445
rect 1740 -5515 1760 -5495
rect 1820 -5365 1840 -5345
rect 1820 -5415 1840 -5395
rect 1820 -5465 1840 -5445
rect 1820 -5515 1840 -5495
rect 1885 -5365 1905 -5345
rect 1885 -5415 1905 -5395
rect 1885 -5465 1905 -5445
rect 1885 -5515 1905 -5495
rect 1965 -5365 1985 -5345
rect 1965 -5415 1985 -5395
rect 1965 -5465 1985 -5445
rect 1965 -5515 1985 -5495
rect 2030 -5365 2050 -5345
rect 2030 -5415 2050 -5395
rect 2030 -5465 2050 -5445
rect 2030 -5515 2050 -5495
rect 1530 -5755 1550 -5735
rect 1530 -5805 1550 -5785
rect 1530 -5855 1550 -5835
rect 1530 -5905 1550 -5885
rect 1595 -5755 1615 -5735
rect 1595 -5805 1615 -5785
rect 1595 -5855 1615 -5835
rect 1595 -5905 1615 -5885
rect 1675 -5755 1695 -5735
rect 1675 -5805 1695 -5785
rect 1675 -5855 1695 -5835
rect 1675 -5905 1695 -5885
rect 1740 -5755 1760 -5735
rect 1740 -5805 1760 -5785
rect 1740 -5855 1760 -5835
rect 1740 -5905 1760 -5885
rect 1820 -5755 1840 -5735
rect 1820 -5805 1840 -5785
rect 1820 -5855 1840 -5835
rect 1820 -5905 1840 -5885
rect 1885 -5755 1905 -5735
rect 1885 -5805 1905 -5785
rect 1885 -5855 1905 -5835
rect 1885 -5905 1905 -5885
rect 1965 -5755 1985 -5735
rect 1965 -5805 1985 -5785
rect 1965 -5855 1985 -5835
rect 1965 -5905 1985 -5885
rect 2030 -5755 2050 -5735
rect 2030 -5805 2050 -5785
rect 2030 -5855 2050 -5835
rect 2030 -5905 2050 -5885
rect 2110 -5755 2130 -5735
rect 2110 -5805 2130 -5785
rect 2110 -5855 2130 -5835
rect 2110 -5905 2130 -5885
rect 2175 -5755 2195 -5735
rect 2175 -5805 2195 -5785
rect 2175 -5855 2195 -5835
rect 2175 -5905 2195 -5885
<< psubdiff >>
rect 1250 35 1290 50
rect 1250 15 1260 35
rect 1280 15 1290 35
rect 1250 0 1290 15
rect 4120 -60 4170 -45
rect 4120 -130 4135 -60
rect 4155 -130 4170 -60
rect 4120 -145 4170 -130
rect -170 -3565 -130 -3550
rect -170 -3585 -160 -3565
rect -140 -3585 -130 -3565
rect -170 -3615 -130 -3585
rect -170 -3635 -160 -3615
rect -140 -3635 -130 -3615
rect -170 -3650 -130 -3635
rect 280 -3565 320 -3550
rect 280 -3585 290 -3565
rect 310 -3585 320 -3565
rect 280 -3615 320 -3585
rect 280 -3635 290 -3615
rect 310 -3635 320 -3615
rect 280 -3650 320 -3635
rect 730 -3565 770 -3550
rect 730 -3585 740 -3565
rect 760 -3585 770 -3565
rect 730 -3615 770 -3585
rect 730 -3635 740 -3615
rect 760 -3635 770 -3615
rect 730 -3650 770 -3635
rect 930 -3565 970 -3550
rect 930 -3585 940 -3565
rect 960 -3585 970 -3565
rect 930 -3615 970 -3585
rect 930 -3635 940 -3615
rect 960 -3635 970 -3615
rect 930 -3650 970 -3635
rect 1095 -3565 1135 -3550
rect 1095 -3585 1105 -3565
rect 1125 -3585 1135 -3565
rect 1095 -3615 1135 -3585
rect 1095 -3635 1105 -3615
rect 1125 -3635 1135 -3615
rect 1095 -3650 1135 -3635
rect 1260 -3565 1300 -3550
rect 1260 -3585 1270 -3565
rect 1290 -3585 1300 -3565
rect 1260 -3615 1300 -3585
rect 1260 -3635 1270 -3615
rect 1290 -3635 1300 -3615
rect 1260 -3650 1300 -3635
rect 4120 -4060 4170 -4045
rect 4120 -4130 4135 -4060
rect 4155 -4130 4170 -4060
rect 4120 -4145 4170 -4130
<< nsubdiff >>
rect 1250 245 1290 260
rect 1250 175 1260 245
rect 1280 175 1290 245
rect 1250 160 1290 175
rect 4120 270 4170 285
rect 4120 100 4135 270
rect 4155 100 4170 270
rect 4120 85 4170 100
rect 4120 -3730 4170 -3715
rect 4120 -3900 4135 -3730
rect 4155 -3900 4170 -3730
rect 4120 -3915 4170 -3900
<< psubdiffcont >>
rect 1260 15 1280 35
rect 4135 -130 4155 -60
rect -160 -3585 -140 -3565
rect -160 -3635 -140 -3615
rect 290 -3585 310 -3565
rect 290 -3635 310 -3615
rect 740 -3585 760 -3565
rect 740 -3635 760 -3615
rect 940 -3585 960 -3565
rect 940 -3635 960 -3615
rect 1105 -3585 1125 -3565
rect 1105 -3635 1125 -3615
rect 1270 -3585 1290 -3565
rect 1270 -3635 1290 -3615
rect 4135 -4130 4155 -4060
<< nsubdiffcont >>
rect 1260 175 1280 245
rect 4135 100 4155 270
rect 4135 -3900 4155 -3730
<< poly >>
rect 755 340 2530 355
rect 185 305 225 315
rect 185 285 195 305
rect 215 285 225 305
rect 185 275 225 285
rect 0 260 15 275
rect 55 260 70 275
rect 260 260 275 275
rect 315 260 330 275
rect 440 260 455 275
rect 495 260 510 275
rect 700 260 715 275
rect 755 260 770 340
rect 880 260 895 275
rect 935 260 950 275
rect 1140 260 1155 275
rect 1195 260 1210 275
rect 1330 260 1345 275
rect 1385 260 1400 275
rect 1590 260 1605 275
rect 1645 260 1660 340
rect 1745 305 1785 315
rect 1745 285 1755 305
rect 1775 285 1785 305
rect 1745 275 1785 285
rect 1770 260 1785 275
rect 1825 260 1840 275
rect 1950 260 1965 275
rect 2075 260 2090 275
rect 2200 260 2215 275
rect 2325 260 2340 275
rect 2450 260 2465 275
rect 125 245 165 255
rect 125 225 135 245
rect 155 225 165 245
rect 125 215 165 225
rect 0 100 15 160
rect -60 85 15 100
rect 0 50 15 85
rect 55 105 70 160
rect 55 95 105 105
rect 55 75 75 95
rect 95 75 105 95
rect 55 65 105 75
rect 150 85 165 215
rect 565 245 605 255
rect 565 225 575 245
rect 595 225 605 245
rect 565 215 605 225
rect 260 85 275 160
rect 150 70 275 85
rect 55 50 70 65
rect 260 50 275 70
rect 315 145 330 160
rect 315 135 365 145
rect 315 115 335 135
rect 355 115 365 135
rect 315 105 365 115
rect 315 50 330 105
rect 440 50 455 160
rect 495 105 510 160
rect 495 95 545 105
rect 495 75 515 95
rect 535 75 545 95
rect 495 65 545 75
rect 590 85 605 215
rect 1005 245 1045 255
rect 1005 225 1015 245
rect 1035 225 1045 245
rect 1005 215 1045 225
rect 700 85 715 160
rect 590 70 715 85
rect 495 50 510 65
rect 700 50 715 70
rect 755 50 770 160
rect 880 50 895 160
rect 935 105 950 160
rect 935 95 985 105
rect 935 75 955 95
rect 975 75 985 95
rect 935 65 985 75
rect 1030 85 1045 215
rect 1455 245 1495 255
rect 1455 225 1465 245
rect 1485 225 1495 245
rect 1455 215 1495 225
rect 1140 85 1155 160
rect 1030 70 1155 85
rect 935 50 950 65
rect 1140 50 1155 70
rect 1195 145 1210 160
rect 1195 135 1245 145
rect 1195 115 1215 135
rect 1235 115 1245 135
rect 1195 105 1245 115
rect 1195 50 1210 105
rect 1330 50 1345 160
rect 1385 105 1400 160
rect 1385 95 1435 105
rect 1385 75 1405 95
rect 1425 75 1435 95
rect 1385 65 1435 75
rect 1480 85 1495 215
rect 1590 85 1605 160
rect 1480 70 1605 85
rect 1385 50 1400 65
rect 1590 50 1605 70
rect 1645 50 1660 160
rect 1770 50 1785 160
rect 1825 50 1840 160
rect 1865 120 1905 130
rect 1865 100 1875 120
rect 1895 115 1905 120
rect 1950 115 1965 160
rect 1895 100 1965 115
rect 1865 90 1905 100
rect 1950 50 1965 100
rect 1990 120 2030 130
rect 1990 100 2000 120
rect 2020 115 2030 120
rect 2075 115 2090 160
rect 2020 100 2090 115
rect 1990 90 2030 100
rect 2075 50 2090 100
rect 2115 120 2155 130
rect 2115 100 2125 120
rect 2145 115 2155 120
rect 2200 115 2215 160
rect 2145 100 2215 115
rect 2115 90 2155 100
rect 2200 50 2215 100
rect 2240 120 2280 130
rect 2240 100 2250 120
rect 2270 115 2280 120
rect 2325 115 2340 160
rect 2270 100 2340 115
rect 2240 90 2280 100
rect 2325 50 2340 100
rect 2365 120 2405 130
rect 2365 100 2375 120
rect 2395 115 2405 120
rect 2450 115 2465 160
rect 2515 130 2530 340
rect 3155 335 4040 350
rect 2865 285 2880 300
rect 3010 285 3025 300
rect 3155 285 3170 335
rect 3300 285 3315 300
rect 3445 285 3460 300
rect 3590 285 3605 300
rect 3735 285 3750 300
rect 3880 285 3895 300
rect 4025 285 4040 335
rect 2395 100 2465 115
rect 2365 90 2405 100
rect 2450 50 2465 100
rect 2490 120 2530 130
rect 2490 100 2500 120
rect 2520 100 2530 120
rect 2490 90 2530 100
rect 2865 30 2880 85
rect 3010 45 3025 85
rect 3155 45 3170 85
rect 3300 70 3315 85
rect 2775 15 2880 30
rect 0 -15 15 0
rect 55 -15 70 0
rect 260 -40 275 0
rect 315 -15 330 0
rect 440 -40 455 0
rect 495 -15 510 0
rect 700 -15 715 0
rect 755 -15 770 0
rect 260 -55 455 -40
rect 880 -80 895 0
rect 935 -15 950 0
rect 1140 -40 1155 0
rect 1195 -15 1210 0
rect 1330 -40 1345 0
rect 1385 -15 1400 0
rect 1590 -15 1605 0
rect 1645 -15 1660 0
rect 1770 -15 1785 0
rect 1825 -15 1840 0
rect 1950 -15 1965 0
rect 2075 -15 2090 0
rect 2200 -15 2215 0
rect 2325 -15 2340 0
rect 2450 -15 2465 0
rect 1140 -55 1345 -40
rect 1825 -25 1865 -15
rect 1825 -45 1835 -25
rect 1855 -45 1865 -25
rect 2865 -45 2880 15
rect 2985 35 3025 45
rect 2985 15 2995 35
rect 3015 15 3025 35
rect 2985 5 3025 15
rect 3130 35 3170 45
rect 3130 15 3140 35
rect 3160 15 3170 35
rect 3195 60 3315 70
rect 3195 40 3205 60
rect 3225 55 3315 60
rect 3225 40 3235 55
rect 3195 30 3235 40
rect 3130 5 3170 15
rect 3010 -45 3025 5
rect 3155 -20 3170 5
rect 3155 -35 3315 -20
rect 3155 -45 3170 -35
rect 3300 -45 3315 -35
rect 3445 -45 3460 85
rect 3590 75 3605 85
rect 3510 60 3605 75
rect 3630 60 3670 70
rect 3735 60 3750 85
rect 3880 60 3895 85
rect 4025 70 4040 85
rect 3510 10 3525 60
rect 3630 40 3640 60
rect 3660 45 4005 60
rect 3660 40 3670 45
rect 3630 35 3670 40
rect 3485 0 3525 10
rect 3670 5 3710 10
rect 3485 -20 3495 0
rect 3515 -20 3525 0
rect 3485 -30 3525 -20
rect 3590 0 3710 5
rect 3590 -10 3680 0
rect 3590 -45 3605 -10
rect 3670 -20 3680 -10
rect 3700 -20 3710 0
rect 3670 -30 3710 -20
rect 3735 -45 3750 45
rect 3990 25 4005 45
rect 3990 10 4040 25
rect 3775 -5 3815 5
rect 3775 -25 3785 -5
rect 3805 -20 3815 -5
rect 3805 -25 3895 -20
rect 3775 -35 3895 -25
rect 3880 -45 3895 -35
rect 4025 -45 4040 10
rect 1825 -55 1865 -45
rect -60 -95 895 -80
rect 2865 -160 2880 -145
rect 3010 -160 3025 -145
rect 3155 -160 3170 -145
rect 3300 -160 3315 -145
rect 3445 -175 3460 -145
rect 3590 -160 3605 -145
rect 3735 -175 3750 -145
rect 3880 -160 3895 -145
rect 3880 -170 3935 -160
rect 3880 -175 3905 -170
rect 3925 -175 3935 -170
rect 4025 -175 4040 -145
rect 260 -1160 455 -1145
rect 0 -1200 15 -1185
rect 55 -1200 70 -1185
rect 260 -1200 275 -1160
rect 315 -1200 330 -1185
rect 440 -1200 455 -1160
rect 915 -1155 955 -1145
rect 915 -1175 925 -1155
rect 945 -1175 955 -1155
rect 915 -1185 955 -1175
rect 495 -1200 510 -1185
rect 700 -1200 715 -1185
rect 755 -1200 770 -1185
rect 940 -1200 955 -1185
rect 995 -1200 1010 -1185
rect 1120 -1200 1135 -1185
rect 1245 -1200 1260 -1185
rect 0 -1285 15 -1250
rect -60 -1300 15 -1285
rect 0 -1360 15 -1300
rect 55 -1265 70 -1250
rect 55 -1275 105 -1265
rect 260 -1270 275 -1250
rect 55 -1295 75 -1275
rect 95 -1295 105 -1275
rect 55 -1305 105 -1295
rect 150 -1285 275 -1270
rect 55 -1360 70 -1305
rect 150 -1415 165 -1285
rect 260 -1360 275 -1285
rect 315 -1305 330 -1250
rect 315 -1315 365 -1305
rect 315 -1335 335 -1315
rect 355 -1335 365 -1315
rect 315 -1345 365 -1335
rect 315 -1360 330 -1345
rect 440 -1360 455 -1250
rect 495 -1265 510 -1250
rect 495 -1275 545 -1265
rect 700 -1270 715 -1250
rect 495 -1295 515 -1275
rect 535 -1295 545 -1275
rect 495 -1305 545 -1295
rect 590 -1285 715 -1270
rect 495 -1360 510 -1305
rect 125 -1425 165 -1415
rect 125 -1445 135 -1425
rect 155 -1445 165 -1425
rect 125 -1455 165 -1445
rect 590 -1415 605 -1285
rect 700 -1360 715 -1285
rect 755 -1270 770 -1250
rect 755 -1280 880 -1270
rect 755 -1285 850 -1280
rect 755 -1360 770 -1285
rect 840 -1300 850 -1285
rect 870 -1300 880 -1280
rect 840 -1310 880 -1300
rect 940 -1360 955 -1250
rect 995 -1360 1010 -1250
rect 1035 -1300 1075 -1290
rect 1120 -1300 1135 -1250
rect 1035 -1320 1045 -1300
rect 1065 -1315 1135 -1300
rect 1065 -1320 1075 -1315
rect 1035 -1330 1075 -1320
rect 1120 -1360 1135 -1315
rect 1160 -1300 1200 -1290
rect 1245 -1300 1260 -1250
rect 1160 -1320 1170 -1300
rect 1190 -1315 1260 -1300
rect 1190 -1320 1200 -1315
rect 1160 -1330 1200 -1320
rect 1245 -1360 1260 -1315
rect 1285 -1300 1325 -1290
rect 1285 -1320 1295 -1300
rect 1315 -1320 1325 -1300
rect 1285 -1330 1325 -1320
rect 565 -1425 605 -1415
rect 565 -1445 575 -1425
rect 595 -1445 605 -1425
rect 565 -1455 605 -1445
rect 0 -1475 15 -1460
rect 55 -1475 70 -1460
rect 260 -1475 275 -1460
rect 315 -1475 330 -1460
rect 440 -1475 455 -1460
rect 495 -1475 510 -1460
rect 700 -1475 715 -1460
rect 755 -1475 770 -1460
rect 940 -1475 955 -1460
rect 995 -1475 1010 -1460
rect 1120 -1475 1135 -1460
rect 1245 -1475 1260 -1460
rect 995 -1485 1035 -1475
rect 995 -1505 1005 -1485
rect 1025 -1505 1035 -1485
rect 995 -1515 1035 -1505
rect 860 -1655 900 -1645
rect 860 -1675 870 -1655
rect 890 -1675 900 -1655
rect 860 -1685 900 -1675
rect 0 -1740 15 -1725
rect 55 -1740 70 -1725
rect 260 -1740 275 -1725
rect 315 -1740 330 -1725
rect 440 -1740 455 -1725
rect 495 -1740 510 -1725
rect 700 -1740 715 -1725
rect 755 -1740 770 -1725
rect 125 -1755 165 -1745
rect 125 -1775 135 -1755
rect 155 -1775 165 -1755
rect 125 -1785 165 -1775
rect 0 -1900 15 -1840
rect -60 -1915 15 -1900
rect 0 -1950 15 -1915
rect 55 -1895 70 -1840
rect 55 -1905 105 -1895
rect 55 -1925 75 -1905
rect 95 -1925 105 -1905
rect 55 -1935 105 -1925
rect 150 -1915 165 -1785
rect 565 -1755 605 -1745
rect 565 -1775 575 -1755
rect 595 -1775 605 -1755
rect 565 -1785 605 -1775
rect 260 -1915 275 -1840
rect 150 -1930 275 -1915
rect 55 -1950 70 -1935
rect 260 -1950 275 -1930
rect 315 -1855 330 -1840
rect 315 -1865 365 -1855
rect 315 -1885 335 -1865
rect 355 -1885 365 -1865
rect 315 -1895 365 -1885
rect 315 -1950 330 -1895
rect 440 -1950 455 -1840
rect 495 -1895 510 -1840
rect 495 -1905 545 -1895
rect 495 -1925 515 -1905
rect 535 -1925 545 -1905
rect 495 -1935 545 -1925
rect 590 -1915 605 -1785
rect 700 -1915 715 -1840
rect 590 -1930 715 -1915
rect 495 -1950 510 -1935
rect 700 -1950 715 -1930
rect 755 -1870 770 -1840
rect 860 -1870 875 -1685
rect 990 -1740 1005 -1725
rect 1115 -1740 1130 -1725
rect 1240 -1740 1255 -1725
rect 755 -1880 965 -1870
rect 755 -1885 935 -1880
rect 755 -1950 770 -1885
rect 925 -1900 935 -1885
rect 955 -1900 965 -1880
rect 925 -1910 965 -1900
rect 990 -1885 1005 -1840
rect 1050 -1880 1090 -1870
rect 1050 -1885 1060 -1880
rect 990 -1900 1060 -1885
rect 1080 -1900 1090 -1880
rect 990 -1950 1005 -1900
rect 1050 -1910 1090 -1900
rect 1115 -1885 1130 -1840
rect 1175 -1880 1215 -1870
rect 1175 -1885 1185 -1880
rect 1115 -1900 1185 -1885
rect 1205 -1900 1215 -1880
rect 1115 -1950 1130 -1900
rect 1175 -1910 1215 -1900
rect 1240 -1885 1255 -1840
rect 1305 -1880 1345 -1870
rect 1305 -1885 1315 -1880
rect 1240 -1900 1315 -1885
rect 1335 -1900 1345 -1880
rect 1240 -1950 1255 -1900
rect 1305 -1910 1345 -1900
rect 0 -2015 15 -2000
rect 55 -2015 70 -2000
rect 260 -2040 275 -2000
rect 315 -2015 330 -2000
rect 440 -2040 455 -2000
rect 495 -2015 510 -2000
rect 700 -2015 715 -2000
rect 755 -2015 770 -2000
rect 990 -2015 1005 -2000
rect 1115 -2015 1130 -2000
rect 1240 -2015 1255 -2000
rect 260 -2055 455 -2040
rect 170 -2610 375 -2595
rect -90 -2650 -75 -2635
rect -35 -2650 -20 -2635
rect 170 -2650 185 -2610
rect 225 -2650 240 -2635
rect 360 -2650 375 -2610
rect 880 -2605 920 -2595
rect 880 -2625 890 -2605
rect 910 -2625 920 -2605
rect 880 -2635 920 -2625
rect 415 -2650 430 -2635
rect 620 -2650 635 -2635
rect 675 -2650 690 -2635
rect 825 -2650 840 -2635
rect 880 -2650 895 -2635
rect 1045 -2650 1060 -2635
rect 1210 -2650 1225 -2635
rect 1565 -2650 1580 -2635
rect 1710 -2650 1725 -2635
rect 1855 -2650 1870 -2635
rect 2000 -2650 2015 -2635
rect -90 -2785 -75 -2750
rect -150 -2800 -75 -2785
rect -90 -2860 -75 -2800
rect -35 -2765 -20 -2750
rect -35 -2775 15 -2765
rect 170 -2770 185 -2750
rect -35 -2795 -15 -2775
rect 5 -2795 15 -2775
rect -35 -2805 15 -2795
rect 60 -2785 185 -2770
rect -35 -2860 -20 -2805
rect 60 -3015 75 -2785
rect 170 -2860 185 -2785
rect 225 -2805 240 -2750
rect 225 -2815 275 -2805
rect 225 -2835 245 -2815
rect 265 -2835 275 -2815
rect 225 -2845 275 -2835
rect 225 -2860 240 -2845
rect 360 -2860 375 -2750
rect 415 -2765 430 -2750
rect 415 -2775 465 -2765
rect 620 -2770 635 -2750
rect 415 -2795 435 -2775
rect 455 -2795 465 -2775
rect 415 -2805 465 -2795
rect 510 -2785 635 -2770
rect 415 -2860 430 -2805
rect 35 -3025 75 -3015
rect 35 -3045 45 -3025
rect 65 -3045 75 -3025
rect 35 -3055 75 -3045
rect 510 -3015 525 -2785
rect 620 -2860 635 -2785
rect 675 -2770 690 -2750
rect 675 -2780 760 -2770
rect 675 -2785 730 -2780
rect 675 -2860 690 -2785
rect 720 -2800 730 -2785
rect 750 -2800 760 -2780
rect 720 -2810 760 -2800
rect 825 -2860 840 -2750
rect 880 -2860 895 -2750
rect 920 -2800 960 -2790
rect 1045 -2800 1060 -2750
rect 920 -2820 930 -2800
rect 950 -2815 1060 -2800
rect 950 -2820 960 -2815
rect 920 -2830 960 -2820
rect 1045 -2860 1060 -2815
rect 1085 -2800 1165 -2790
rect 1210 -2800 1225 -2750
rect 1085 -2820 1095 -2800
rect 1155 -2815 1225 -2800
rect 1155 -2820 1165 -2815
rect 1085 -2830 1165 -2820
rect 1210 -2860 1225 -2815
rect 1250 -2800 1290 -2790
rect 1565 -2800 1580 -2750
rect 1710 -2790 1725 -2750
rect 1855 -2760 1870 -2750
rect 2000 -2760 2015 -2750
rect 1855 -2775 2160 -2760
rect 1855 -2790 1870 -2775
rect 1250 -2820 1260 -2800
rect 1280 -2820 1290 -2800
rect 1530 -2815 1580 -2800
rect 1250 -2830 1290 -2820
rect 1565 -2860 1580 -2815
rect 1685 -2800 1725 -2790
rect 1685 -2820 1695 -2800
rect 1715 -2820 1725 -2800
rect 1685 -2830 1725 -2820
rect 1830 -2800 1870 -2790
rect 1830 -2820 1840 -2800
rect 1860 -2820 1870 -2800
rect 1830 -2830 1870 -2820
rect 1710 -2860 1725 -2830
rect 1855 -2860 1870 -2830
rect 1895 -2815 1935 -2805
rect 1895 -2835 1905 -2815
rect 1925 -2830 1935 -2815
rect 1925 -2835 2015 -2830
rect 1895 -2845 2015 -2835
rect 2000 -2860 2015 -2845
rect 2145 -2860 2160 -2775
rect 485 -3025 525 -3015
rect 485 -3045 495 -3025
rect 515 -3045 525 -3025
rect 485 -3055 525 -3045
rect -90 -3075 -75 -3060
rect -35 -3075 -20 -3060
rect 170 -3075 185 -3060
rect 225 -3075 240 -3060
rect 360 -3075 375 -3060
rect 415 -3075 430 -3060
rect 620 -3075 635 -3060
rect 675 -3075 690 -3060
rect 825 -3075 840 -3060
rect 880 -3075 895 -3060
rect 1045 -3075 1060 -3060
rect 1210 -3075 1225 -3060
rect 1565 -3075 1580 -3060
rect 1710 -3075 1725 -3060
rect 1855 -3075 1870 -3060
rect 2000 -3075 2015 -3060
rect 2145 -3075 2160 -3060
rect 795 -3085 840 -3075
rect 795 -3105 805 -3085
rect 825 -3105 840 -3085
rect 795 -3115 840 -3105
rect 1685 -3225 1725 -3185
rect 1975 -3225 2015 -3185
rect -90 -3240 -75 -3225
rect -35 -3240 -20 -3225
rect 170 -3240 185 -3225
rect 225 -3240 240 -3225
rect 360 -3240 375 -3225
rect 415 -3240 430 -3225
rect 620 -3240 635 -3225
rect 675 -3240 690 -3225
rect 875 -3240 890 -3225
rect 1040 -3240 1055 -3225
rect 1205 -3240 1220 -3225
rect 1565 -3240 1580 -3225
rect 1710 -3240 1725 -3225
rect 1855 -3240 1870 -3225
rect 2000 -3240 2015 -3225
rect 35 -3255 75 -3245
rect 35 -3275 45 -3255
rect 65 -3275 75 -3255
rect 35 -3285 75 -3275
rect -90 -3500 -75 -3440
rect -150 -3515 -75 -3500
rect -90 -3550 -75 -3515
rect -35 -3495 -20 -3440
rect -35 -3505 15 -3495
rect -35 -3525 -15 -3505
rect 5 -3525 15 -3505
rect -35 -3535 15 -3525
rect 60 -3515 75 -3285
rect 485 -3255 525 -3245
rect 485 -3275 495 -3255
rect 515 -3275 525 -3255
rect 485 -3285 525 -3275
rect 170 -3515 185 -3440
rect 60 -3530 185 -3515
rect -35 -3550 -20 -3535
rect 170 -3550 185 -3530
rect 225 -3455 240 -3440
rect 225 -3465 275 -3455
rect 225 -3485 245 -3465
rect 265 -3485 275 -3465
rect 225 -3495 275 -3485
rect 225 -3550 240 -3495
rect 360 -3550 375 -3440
rect 415 -3495 430 -3440
rect 415 -3505 465 -3495
rect 415 -3525 435 -3505
rect 455 -3525 465 -3505
rect 415 -3535 465 -3525
rect 510 -3515 525 -3285
rect 620 -3515 635 -3440
rect 510 -3530 635 -3515
rect 415 -3550 430 -3535
rect 620 -3550 635 -3530
rect 675 -3470 690 -3440
rect 675 -3480 850 -3470
rect 675 -3485 740 -3480
rect 675 -3550 690 -3485
rect 730 -3500 740 -3485
rect 760 -3485 820 -3480
rect 760 -3500 770 -3485
rect 730 -3510 770 -3500
rect 810 -3500 820 -3485
rect 840 -3500 850 -3480
rect 810 -3510 850 -3500
rect 875 -3485 890 -3440
rect 975 -3480 1015 -3470
rect 975 -3485 985 -3480
rect 875 -3500 985 -3485
rect 1005 -3500 1015 -3480
rect 875 -3550 890 -3500
rect 975 -3510 1015 -3500
rect 1040 -3485 1055 -3440
rect 1140 -3480 1180 -3470
rect 1140 -3485 1150 -3480
rect 1040 -3500 1150 -3485
rect 1170 -3500 1180 -3480
rect 1040 -3550 1055 -3500
rect 1140 -3510 1180 -3500
rect 1205 -3485 1220 -3440
rect 1270 -3480 1310 -3470
rect 1270 -3485 1280 -3480
rect 1205 -3500 1280 -3485
rect 1300 -3500 1310 -3480
rect 1565 -3500 1580 -3440
rect 1710 -3455 1725 -3440
rect 1750 -3465 1790 -3455
rect 1855 -3465 1870 -3440
rect 2000 -3465 2015 -3440
rect 1750 -3485 1760 -3465
rect 1780 -3480 2160 -3465
rect 1780 -3485 1790 -3480
rect 1750 -3495 1790 -3485
rect 1205 -3550 1220 -3500
rect 1270 -3510 1310 -3500
rect 1475 -3515 1580 -3500
rect 1565 -3550 1580 -3515
rect 1710 -3550 1725 -3535
rect 1855 -3550 1870 -3480
rect 1895 -3510 1935 -3505
rect 1895 -3530 1905 -3510
rect 1925 -3525 1935 -3510
rect 2000 -3525 2015 -3480
rect 1925 -3530 2015 -3525
rect 1895 -3540 2015 -3530
rect 2000 -3550 2015 -3540
rect 2145 -3550 2160 -3480
rect -90 -3665 -75 -3650
rect -35 -3665 -20 -3650
rect 170 -3690 185 -3650
rect 225 -3665 240 -3650
rect 360 -3690 375 -3650
rect 415 -3665 430 -3650
rect 620 -3665 635 -3650
rect 675 -3665 690 -3650
rect 875 -3665 890 -3650
rect 1040 -3665 1055 -3650
rect 1205 -3665 1220 -3650
rect 1565 -3665 1580 -3650
rect 1710 -3665 1725 -3650
rect 1855 -3665 1870 -3650
rect 2000 -3665 2015 -3650
rect 2145 -3665 2160 -3650
rect 3155 -3665 4040 -3650
rect 170 -3705 375 -3690
rect 1710 -3675 1765 -3665
rect 1710 -3695 1735 -3675
rect 1755 -3695 1765 -3675
rect 1710 -3705 1765 -3695
rect 2000 -3675 2055 -3665
rect 2000 -3695 2025 -3675
rect 2045 -3695 2055 -3675
rect 2000 -3705 2055 -3695
rect 2865 -3715 2880 -3700
rect 3010 -3715 3025 -3700
rect 3155 -3715 3170 -3665
rect 3300 -3715 3315 -3700
rect 3445 -3715 3460 -3700
rect 3590 -3715 3605 -3700
rect 3735 -3715 3750 -3700
rect 3880 -3715 3895 -3700
rect 4025 -3715 4040 -3665
rect 2865 -3970 2880 -3915
rect 3010 -3955 3025 -3915
rect 3155 -3955 3170 -3915
rect 3300 -3930 3315 -3915
rect 2775 -3985 2880 -3970
rect 2865 -4045 2880 -3985
rect 2985 -3965 3025 -3955
rect 2985 -3985 2995 -3965
rect 3015 -3985 3025 -3965
rect 2985 -3995 3025 -3985
rect 3130 -3965 3170 -3955
rect 3130 -3985 3140 -3965
rect 3160 -3985 3170 -3965
rect 3195 -3940 3315 -3930
rect 3195 -3960 3205 -3940
rect 3225 -3945 3315 -3940
rect 3225 -3960 3235 -3945
rect 3195 -3970 3235 -3960
rect 3130 -3995 3170 -3985
rect 3010 -4045 3025 -3995
rect 3155 -4020 3170 -3995
rect 3155 -4035 3315 -4020
rect 3155 -4045 3170 -4035
rect 3300 -4045 3315 -4035
rect 3445 -4045 3460 -3915
rect 3590 -3925 3605 -3915
rect 3510 -3940 3605 -3925
rect 3630 -3940 3670 -3930
rect 3735 -3940 3750 -3915
rect 3880 -3940 3895 -3915
rect 4025 -3930 4040 -3915
rect 3510 -3990 3525 -3940
rect 3630 -3960 3640 -3940
rect 3660 -3955 4005 -3940
rect 3660 -3960 3670 -3955
rect 3630 -3965 3670 -3960
rect 3485 -4000 3525 -3990
rect 3670 -3995 3710 -3990
rect 3485 -4020 3495 -4000
rect 3515 -4020 3525 -4000
rect 3485 -4030 3525 -4020
rect 3590 -4000 3710 -3995
rect 3590 -4010 3680 -4000
rect 3590 -4045 3605 -4010
rect 3670 -4020 3680 -4010
rect 3700 -4020 3710 -4000
rect 3670 -4030 3710 -4020
rect 3735 -4045 3750 -3955
rect 3990 -3975 4005 -3955
rect 3990 -3990 4040 -3975
rect 3775 -4005 3815 -3995
rect 3775 -4025 3785 -4005
rect 3805 -4020 3815 -4005
rect 3805 -4025 3895 -4020
rect 3775 -4035 3895 -4025
rect 3880 -4045 3895 -4035
rect 4025 -4045 4040 -3990
rect 2865 -4160 2880 -4145
rect 3010 -4160 3025 -4145
rect 3155 -4160 3170 -4145
rect 3300 -4160 3315 -4145
rect 3445 -4175 3460 -4145
rect 3590 -4160 3605 -4145
rect 3735 -4175 3750 -4145
rect 3880 -4160 3895 -4145
rect 3880 -4170 3935 -4160
rect 3880 -4175 3905 -4170
rect 3925 -4175 3935 -4170
rect 4025 -4175 4040 -4145
rect 1565 -5100 1580 -5085
rect 1710 -5100 1725 -5085
rect 1855 -5100 1870 -5085
rect 2000 -5100 2015 -5085
rect 1565 -5260 1580 -5200
rect 1710 -5250 1725 -5200
rect 1855 -5210 1870 -5200
rect 2000 -5210 2015 -5200
rect 1855 -5225 2015 -5210
rect 1855 -5250 1870 -5225
rect 1475 -5275 1580 -5260
rect 1565 -5330 1580 -5275
rect 1685 -5260 1725 -5250
rect 1685 -5280 1695 -5260
rect 1715 -5280 1725 -5260
rect 1685 -5290 1725 -5280
rect 1830 -5260 1870 -5250
rect 1830 -5280 1840 -5260
rect 1860 -5280 1870 -5260
rect 1830 -5290 1870 -5280
rect 1710 -5330 1725 -5290
rect 1855 -5330 1870 -5290
rect 1895 -5285 1935 -5275
rect 1895 -5305 1905 -5285
rect 1925 -5300 1935 -5285
rect 1925 -5305 2015 -5300
rect 1895 -5315 2015 -5305
rect 2000 -5330 2015 -5315
rect 1565 -5545 1580 -5530
rect 1710 -5545 1725 -5530
rect 1855 -5545 1870 -5530
rect 2000 -5545 2015 -5530
rect 1565 -5720 1580 -5705
rect 1710 -5720 1725 -5705
rect 1855 -5720 1870 -5705
rect 2000 -5720 2015 -5705
rect 2145 -5720 2160 -5705
rect 1565 -6050 1580 -5920
rect 1710 -5930 1725 -5920
rect 1630 -5945 1725 -5930
rect 1750 -5945 1790 -5935
rect 1855 -5945 1870 -5920
rect 2000 -5945 2015 -5920
rect 2145 -5935 2160 -5920
rect 1630 -5995 1645 -5945
rect 1750 -5965 1760 -5945
rect 1780 -5960 2125 -5945
rect 1780 -5965 1790 -5960
rect 1750 -5970 1790 -5965
rect 1605 -6005 1645 -5995
rect 1790 -6000 1830 -5995
rect 1605 -6025 1615 -6005
rect 1635 -6025 1645 -6005
rect 1605 -6035 1645 -6025
rect 1710 -6005 1830 -6000
rect 1710 -6015 1800 -6005
rect 1710 -6050 1725 -6015
rect 1790 -6025 1800 -6015
rect 1820 -6025 1830 -6005
rect 1790 -6035 1830 -6025
rect 1855 -6050 1870 -5960
rect 2110 -5980 2125 -5960
rect 2110 -5995 2160 -5980
rect 1895 -6010 1935 -6000
rect 1895 -6030 1905 -6010
rect 1925 -6025 1935 -6010
rect 1925 -6030 2015 -6025
rect 1895 -6040 2015 -6030
rect 2000 -6050 2015 -6040
rect 2145 -6050 2160 -5995
rect 1565 -6165 1580 -6150
rect 1710 -6165 1725 -6150
rect 1855 -6165 1870 -6150
rect 2000 -6165 2015 -6150
rect 2145 -6165 2160 -6150
<< polycont >>
rect 195 285 215 305
rect 1755 285 1775 305
rect 135 225 155 245
rect 75 75 95 95
rect 575 225 595 245
rect 335 115 355 135
rect 515 75 535 95
rect 1015 225 1035 245
rect 955 75 975 95
rect 1465 225 1485 245
rect 1215 115 1235 135
rect 1405 75 1425 95
rect 1875 100 1895 120
rect 2000 100 2020 120
rect 2125 100 2145 120
rect 2250 100 2270 120
rect 2375 100 2395 120
rect 2500 100 2520 120
rect 1835 -45 1855 -25
rect 2995 15 3015 35
rect 3140 15 3160 35
rect 3205 40 3225 60
rect 3640 40 3660 60
rect 3495 -20 3515 0
rect 3680 -20 3700 0
rect 3785 -25 3805 -5
rect 3905 -175 3925 -170
rect 925 -1175 945 -1155
rect 75 -1295 95 -1275
rect 335 -1335 355 -1315
rect 515 -1295 535 -1275
rect 135 -1445 155 -1425
rect 850 -1300 870 -1280
rect 1045 -1320 1065 -1300
rect 1170 -1320 1190 -1300
rect 1295 -1320 1315 -1300
rect 575 -1445 595 -1425
rect 1005 -1505 1025 -1485
rect 870 -1675 890 -1655
rect 135 -1775 155 -1755
rect 75 -1925 95 -1905
rect 575 -1775 595 -1755
rect 335 -1885 355 -1865
rect 515 -1925 535 -1905
rect 935 -1900 955 -1880
rect 1060 -1900 1080 -1880
rect 1185 -1900 1205 -1880
rect 1315 -1900 1335 -1880
rect 890 -2625 910 -2605
rect -15 -2795 5 -2775
rect 245 -2835 265 -2815
rect 435 -2795 455 -2775
rect 45 -3045 65 -3025
rect 730 -2800 750 -2780
rect 930 -2820 950 -2800
rect 1095 -2820 1155 -2800
rect 1260 -2820 1280 -2800
rect 1695 -2820 1715 -2800
rect 1840 -2820 1860 -2800
rect 1905 -2835 1925 -2815
rect 495 -3045 515 -3025
rect 805 -3105 825 -3085
rect 45 -3275 65 -3255
rect -15 -3525 5 -3505
rect 495 -3275 515 -3255
rect 245 -3485 265 -3465
rect 435 -3525 455 -3505
rect 740 -3500 760 -3480
rect 820 -3500 840 -3480
rect 985 -3500 1005 -3480
rect 1150 -3500 1170 -3480
rect 1280 -3500 1300 -3480
rect 1760 -3485 1780 -3465
rect 1905 -3530 1925 -3510
rect 1735 -3695 1755 -3675
rect 2025 -3695 2045 -3675
rect 2995 -3985 3015 -3965
rect 3140 -3985 3160 -3965
rect 3205 -3960 3225 -3940
rect 3640 -3960 3660 -3940
rect 3495 -4020 3515 -4000
rect 3680 -4020 3700 -4000
rect 3785 -4025 3805 -4005
rect 3905 -4175 3925 -4170
rect 1695 -5280 1715 -5260
rect 1840 -5280 1860 -5260
rect 1905 -5305 1925 -5285
rect 1760 -5965 1780 -5945
rect 1615 -6025 1635 -6005
rect 1800 -6025 1820 -6005
rect 1905 -6030 1925 -6010
<< locali >>
rect 185 305 225 315
rect 185 285 195 305
rect 215 295 225 305
rect 1745 305 1785 315
rect 1745 295 1755 305
rect 215 285 1755 295
rect 1775 295 1785 305
rect 1775 285 2530 295
rect 185 275 2530 285
rect 3185 280 3205 355
rect 3265 280 3285 355
rect 3330 300 4200 320
rect 3330 280 3350 300
rect 4055 280 4075 300
rect 185 255 205 275
rect 2820 270 2860 280
rect -35 245 -5 255
rect -35 175 -30 245
rect -10 175 -5 245
rect -35 165 -5 175
rect 20 245 50 255
rect 20 175 25 245
rect 45 175 50 245
rect 20 165 50 175
rect 75 245 165 255
rect 75 175 80 245
rect 100 230 135 245
rect 100 175 105 230
rect 125 225 135 230
rect 155 225 165 245
rect 125 215 165 225
rect 185 245 255 255
rect 185 235 230 245
rect 75 165 105 175
rect 80 145 100 165
rect 20 125 100 145
rect 20 45 40 125
rect 185 105 205 235
rect 225 175 230 235
rect 250 175 255 245
rect 225 165 255 175
rect 280 245 310 255
rect 280 175 285 245
rect 305 175 310 245
rect 280 165 310 175
rect 335 245 365 255
rect 335 175 340 245
rect 360 175 365 245
rect 335 165 365 175
rect 405 245 435 255
rect 405 175 410 245
rect 430 175 435 245
rect 405 165 435 175
rect 460 245 490 255
rect 460 175 465 245
rect 485 175 490 245
rect 460 165 490 175
rect 515 245 605 255
rect 515 175 520 245
rect 540 230 575 245
rect 540 175 545 230
rect 565 225 575 230
rect 595 225 605 245
rect 565 215 605 225
rect 625 245 695 255
rect 625 235 670 245
rect 515 165 545 175
rect 230 145 250 165
rect 520 145 540 165
rect 230 125 305 145
rect 65 95 205 105
rect 65 75 75 95
rect 95 85 205 95
rect 95 75 105 85
rect 65 65 105 75
rect 285 45 305 125
rect 325 135 540 145
rect 325 115 335 135
rect 355 125 540 135
rect 355 115 365 125
rect 325 105 365 115
rect 460 45 480 125
rect 625 105 645 235
rect 665 175 670 235
rect 690 175 695 245
rect 665 165 695 175
rect 720 245 750 255
rect 720 175 725 245
rect 745 175 750 245
rect 720 165 750 175
rect 775 245 805 255
rect 775 175 780 245
rect 800 175 805 245
rect 775 165 805 175
rect 845 245 875 255
rect 845 175 850 245
rect 870 175 875 245
rect 845 165 875 175
rect 900 245 930 255
rect 900 175 905 245
rect 925 175 930 245
rect 900 165 930 175
rect 955 245 1045 255
rect 955 175 960 245
rect 980 230 1015 245
rect 980 175 985 230
rect 1005 225 1015 230
rect 1035 225 1045 245
rect 1005 215 1045 225
rect 1065 245 1135 255
rect 1065 235 1110 245
rect 955 165 985 175
rect 670 145 690 165
rect 960 145 980 165
rect 670 125 745 145
rect 505 95 645 105
rect 505 75 515 95
rect 535 85 645 95
rect 535 75 545 85
rect 505 65 545 75
rect 725 45 745 125
rect 900 125 980 145
rect 900 45 920 125
rect 1065 105 1085 235
rect 1105 175 1110 235
rect 1130 175 1135 245
rect 1105 165 1135 175
rect 1160 245 1190 255
rect 1160 175 1165 245
rect 1185 175 1190 245
rect 1160 165 1190 175
rect 1215 245 1325 255
rect 1215 175 1220 245
rect 1240 175 1260 245
rect 1280 175 1300 245
rect 1320 175 1325 245
rect 1215 165 1325 175
rect 1350 245 1380 255
rect 1350 175 1355 245
rect 1375 175 1380 245
rect 1350 165 1380 175
rect 1405 245 1495 255
rect 1405 175 1410 245
rect 1430 230 1465 245
rect 1430 175 1435 230
rect 1455 225 1465 230
rect 1485 225 1495 245
rect 1455 215 1495 225
rect 1515 245 1585 255
rect 1515 235 1560 245
rect 1405 165 1435 175
rect 1110 145 1130 165
rect 1410 145 1430 165
rect 1110 125 1185 145
rect 945 95 1085 105
rect 945 75 955 95
rect 975 85 1085 95
rect 975 75 985 85
rect 945 65 985 75
rect 1165 45 1185 125
rect 1205 135 1430 145
rect 1205 115 1215 135
rect 1235 125 1430 135
rect 1235 115 1245 125
rect 1205 105 1245 115
rect 1350 45 1370 125
rect 1515 105 1535 235
rect 1555 175 1560 235
rect 1580 175 1585 245
rect 1555 165 1585 175
rect 1610 245 1640 255
rect 1610 175 1615 245
rect 1635 175 1640 245
rect 1610 165 1640 175
rect 1665 245 1695 255
rect 1665 175 1670 245
rect 1690 175 1695 245
rect 1665 165 1695 175
rect 1735 245 1765 255
rect 1735 175 1740 245
rect 1760 175 1765 245
rect 1735 165 1765 175
rect 1790 245 1820 255
rect 1790 175 1795 245
rect 1815 175 1820 245
rect 1790 165 1820 175
rect 1845 245 1875 255
rect 1845 175 1850 245
rect 1870 175 1875 245
rect 1845 165 1875 175
rect 1915 245 1945 255
rect 1915 175 1920 245
rect 1940 175 1945 245
rect 1915 165 1945 175
rect 1970 245 2000 255
rect 1970 175 1975 245
rect 1995 175 2000 245
rect 1970 165 2000 175
rect 2040 245 2070 255
rect 2040 175 2045 245
rect 2065 175 2070 245
rect 2040 165 2070 175
rect 2095 245 2125 255
rect 2095 175 2100 245
rect 2120 175 2125 245
rect 2095 165 2125 175
rect 2165 245 2195 255
rect 2165 175 2170 245
rect 2190 175 2195 245
rect 2165 165 2195 175
rect 2220 245 2250 255
rect 2220 175 2225 245
rect 2245 175 2250 245
rect 2220 165 2250 175
rect 2290 245 2320 255
rect 2290 175 2295 245
rect 2315 175 2320 245
rect 2290 165 2320 175
rect 2345 245 2375 255
rect 2345 175 2350 245
rect 2370 175 2375 245
rect 2345 165 2375 175
rect 2415 245 2445 255
rect 2415 175 2420 245
rect 2440 175 2445 245
rect 2415 165 2445 175
rect 2470 245 2500 255
rect 2470 175 2475 245
rect 2495 175 2500 245
rect 2470 165 2500 175
rect 1560 145 1580 165
rect 1740 145 1760 165
rect 1850 145 1870 165
rect 1560 125 1635 145
rect 1740 130 1870 145
rect 1980 130 2000 165
rect 2105 130 2125 165
rect 2230 130 2250 165
rect 2355 130 2375 165
rect 2480 130 2500 165
rect 1740 125 1905 130
rect 1395 95 1535 105
rect 1395 75 1405 95
rect 1425 85 1535 95
rect 1425 75 1435 85
rect 1395 65 1435 75
rect 1615 45 1635 125
rect 1850 120 1905 125
rect 1850 100 1875 120
rect 1895 100 1905 120
rect 1850 90 1905 100
rect 1980 120 2030 130
rect 1980 100 2000 120
rect 2020 100 2030 120
rect 1980 90 2030 100
rect 2105 120 2155 130
rect 2105 100 2125 120
rect 2145 100 2155 120
rect 2105 90 2155 100
rect 2230 120 2280 130
rect 2230 100 2250 120
rect 2270 100 2280 120
rect 2230 90 2280 100
rect 2355 120 2405 130
rect 2355 100 2375 120
rect 2395 100 2405 120
rect 2355 90 2405 100
rect 2480 120 2530 130
rect 2480 100 2500 120
rect 2520 100 2530 120
rect 2480 90 2530 100
rect 2820 100 2830 270
rect 2850 100 2860 270
rect 2820 90 2860 100
rect 2885 270 2925 280
rect 2885 100 2895 270
rect 2915 100 2925 270
rect 2885 90 2925 100
rect 2965 270 3005 280
rect 2965 100 2975 270
rect 2995 100 3005 270
rect 2965 90 3005 100
rect 3030 270 3070 280
rect 3030 100 3040 270
rect 3060 100 3070 270
rect 3030 90 3070 100
rect 3110 270 3150 280
rect 3110 100 3120 270
rect 3140 100 3150 270
rect 3110 90 3150 100
rect 3175 270 3215 280
rect 3175 100 3185 270
rect 3205 100 3215 270
rect 3175 90 3215 100
rect 3255 270 3295 280
rect 3255 100 3265 270
rect 3285 100 3295 270
rect 3255 90 3295 100
rect 3320 270 3360 280
rect 3320 100 3330 270
rect 3350 100 3360 270
rect 3320 90 3360 100
rect 3400 270 3440 280
rect 3400 100 3410 270
rect 3430 100 3440 270
rect 3400 90 3440 100
rect 3465 270 3505 280
rect 3465 100 3475 270
rect 3495 120 3505 270
rect 3545 270 3585 280
rect 3495 100 3510 120
rect 3465 90 3510 100
rect 3545 100 3555 270
rect 3575 100 3585 270
rect 3545 90 3585 100
rect 3610 270 3650 280
rect 3610 100 3620 270
rect 3640 100 3650 270
rect 3610 90 3650 100
rect 3690 270 3730 280
rect 3690 100 3700 270
rect 3720 100 3730 270
rect 3690 90 3730 100
rect 3755 270 3795 280
rect 3755 100 3765 270
rect 3785 100 3795 270
rect 3755 90 3795 100
rect 3835 270 3875 280
rect 3835 100 3845 270
rect 3865 100 3875 270
rect 3835 90 3875 100
rect 3900 270 3940 280
rect 3900 100 3910 270
rect 3930 100 3940 270
rect 3900 90 3940 100
rect 3980 270 4020 280
rect 3980 100 3990 270
rect 4010 100 4020 270
rect 3980 90 4020 100
rect 4045 270 4085 280
rect 4045 100 4055 270
rect 4075 100 4085 270
rect 4045 90 4085 100
rect 4125 270 4165 280
rect 4125 100 4135 270
rect 4155 100 4165 270
rect 4125 90 4165 100
rect 1850 45 1870 90
rect 1980 45 2000 90
rect 2105 45 2125 90
rect 2230 45 2250 90
rect 2355 45 2375 90
rect 2480 45 2500 90
rect -35 35 -5 45
rect -35 15 -30 35
rect -10 15 -5 35
rect -35 5 -5 15
rect 20 35 50 45
rect 20 15 25 35
rect 45 15 50 35
rect 20 5 50 15
rect 75 35 105 45
rect 75 15 80 35
rect 100 15 105 35
rect 75 5 105 15
rect 225 35 255 45
rect 225 15 230 35
rect 250 15 255 35
rect 225 5 255 15
rect 280 35 310 45
rect 280 15 285 35
rect 305 15 310 35
rect 280 5 310 15
rect 335 35 365 45
rect 335 15 340 35
rect 360 15 365 35
rect 335 5 365 15
rect 405 35 435 45
rect 405 15 410 35
rect 430 15 435 35
rect 405 5 435 15
rect 460 35 490 45
rect 460 15 465 35
rect 485 15 490 35
rect 460 5 490 15
rect 515 35 545 45
rect 515 15 520 35
rect 540 15 545 35
rect 515 5 545 15
rect 665 35 695 45
rect 665 15 670 35
rect 690 15 695 35
rect 665 5 695 15
rect 720 35 750 45
rect 720 15 725 35
rect 745 15 750 35
rect 720 5 750 15
rect 775 35 805 45
rect 775 15 780 35
rect 800 15 805 35
rect 775 5 805 15
rect 845 35 875 45
rect 845 15 850 35
rect 870 15 875 35
rect 845 5 875 15
rect 900 35 930 45
rect 900 15 905 35
rect 925 15 930 35
rect 900 5 930 15
rect 955 35 985 45
rect 955 15 960 35
rect 980 15 985 35
rect 955 5 985 15
rect 1105 35 1135 45
rect 1105 15 1110 35
rect 1130 15 1135 35
rect 1105 5 1135 15
rect 1160 35 1190 45
rect 1160 15 1165 35
rect 1185 15 1190 35
rect 1160 5 1190 15
rect 1215 35 1325 45
rect 1215 15 1220 35
rect 1240 15 1260 35
rect 1280 15 1300 35
rect 1320 15 1325 35
rect 1215 5 1325 15
rect 1350 35 1380 45
rect 1350 15 1355 35
rect 1375 15 1380 35
rect 1350 5 1380 15
rect 1405 35 1435 45
rect 1405 15 1410 35
rect 1430 15 1435 35
rect 1405 5 1435 15
rect 1555 35 1585 45
rect 1555 15 1560 35
rect 1580 15 1585 35
rect 1555 5 1585 15
rect 1610 35 1640 45
rect 1610 15 1615 35
rect 1635 15 1640 35
rect 1610 5 1640 15
rect 1665 35 1695 45
rect 1665 15 1670 35
rect 1690 15 1695 35
rect 1665 5 1695 15
rect 1735 35 1765 45
rect 1735 15 1740 35
rect 1760 15 1765 35
rect 1735 5 1765 15
rect 1790 35 1820 45
rect 1790 15 1795 35
rect 1815 15 1820 35
rect 1790 5 1820 15
rect 1845 35 1875 45
rect 1845 15 1850 35
rect 1870 15 1875 35
rect 1845 5 1875 15
rect 1915 35 1945 45
rect 1915 15 1920 35
rect 1940 15 1945 35
rect 1915 5 1945 15
rect 1970 35 2000 45
rect 1970 15 1975 35
rect 1995 15 2000 35
rect 1970 5 2000 15
rect 2040 35 2070 45
rect 2040 15 2045 35
rect 2065 15 2070 35
rect 2040 5 2070 15
rect 2095 35 2125 45
rect 2095 15 2100 35
rect 2120 15 2125 35
rect 2095 5 2125 15
rect 2165 35 2195 45
rect 2165 15 2170 35
rect 2190 15 2195 35
rect 2165 5 2195 15
rect 2220 35 2250 45
rect 2220 15 2225 35
rect 2245 15 2250 35
rect 2220 5 2250 15
rect 2290 35 2320 45
rect 2290 15 2295 35
rect 2315 15 2320 35
rect 2290 5 2320 15
rect 2345 35 2375 45
rect 2345 15 2350 35
rect 2370 15 2375 35
rect 2345 5 2375 15
rect 2415 35 2445 45
rect 2415 15 2420 35
rect 2440 15 2445 35
rect 2415 5 2445 15
rect 2470 35 2500 45
rect 2470 15 2475 35
rect 2495 15 2500 35
rect 2470 5 2500 15
rect 2905 35 2925 90
rect 2985 35 3025 45
rect 2905 15 2995 35
rect 3015 15 3025 35
rect 1165 -15 1185 5
rect 1165 -25 2530 -15
rect 1165 -35 1835 -25
rect 1825 -45 1835 -35
rect 1855 -35 2530 -25
rect 1855 -45 1865 -35
rect 1825 -55 1865 -45
rect 2905 -50 2925 15
rect 2985 5 3025 15
rect 3050 35 3070 90
rect 3195 70 3215 90
rect 3195 60 3235 70
rect 3130 35 3170 45
rect 3050 15 3140 35
rect 3160 15 3170 35
rect 3050 -50 3070 15
rect 3130 5 3170 15
rect 3195 40 3205 60
rect 3225 40 3235 60
rect 3195 30 3235 40
rect 3195 -50 3215 30
rect 3265 -50 3285 90
rect 3320 -50 3340 90
rect 3420 70 3440 90
rect 3555 70 3575 90
rect 3420 50 3575 70
rect 3420 -50 3440 50
rect 3485 0 3525 10
rect 3485 -20 3495 0
rect 3515 -20 3525 0
rect 3485 -30 3525 -20
rect 3485 -50 3505 -30
rect 3555 -50 3575 50
rect 3620 70 3640 90
rect 3620 60 3670 70
rect 3620 40 3640 60
rect 3660 40 3670 60
rect 3620 35 3670 40
rect 3620 -50 3640 35
rect 3695 10 3715 90
rect 3670 0 3715 10
rect 3670 -20 3680 0
rect 3700 -20 3715 0
rect 3670 -30 3715 -20
rect 3775 5 3795 90
rect 3775 -5 3815 5
rect 3775 -25 3785 -5
rect 3805 -25 3815 -5
rect 3775 -35 3815 -25
rect 3775 -50 3795 -35
rect 3845 -50 3865 90
rect 3910 10 3930 90
rect 3910 -10 4200 10
rect 3910 -50 3930 -10
rect 4055 -50 4075 -10
rect 2820 -60 2860 -50
rect 2820 -130 2830 -60
rect 2850 -130 2860 -60
rect 2820 -140 2860 -130
rect 2885 -60 2925 -50
rect 2885 -130 2895 -60
rect 2915 -130 2925 -60
rect 2885 -140 2925 -130
rect 2965 -60 3005 -50
rect 2965 -130 2975 -60
rect 2995 -130 3005 -60
rect 2965 -140 3005 -130
rect 3030 -60 3070 -50
rect 3030 -130 3040 -60
rect 3060 -130 3070 -60
rect 3030 -140 3070 -130
rect 3110 -60 3150 -50
rect 3110 -130 3120 -60
rect 3140 -130 3150 -60
rect 3110 -140 3150 -130
rect 3175 -60 3215 -50
rect 3175 -130 3185 -60
rect 3205 -130 3215 -60
rect 3175 -140 3215 -130
rect 3255 -60 3295 -50
rect 3255 -130 3265 -60
rect 3285 -130 3295 -60
rect 3255 -140 3295 -130
rect 3320 -60 3360 -50
rect 3320 -130 3330 -60
rect 3350 -130 3360 -60
rect 3320 -140 3360 -130
rect 3400 -60 3440 -50
rect 3400 -130 3410 -60
rect 3430 -130 3440 -60
rect 3400 -140 3440 -130
rect 3465 -60 3505 -50
rect 3465 -130 3475 -60
rect 3495 -130 3505 -60
rect 3465 -140 3505 -130
rect 3545 -60 3585 -50
rect 3545 -130 3555 -60
rect 3575 -130 3585 -60
rect 3545 -140 3585 -130
rect 3610 -60 3650 -50
rect 3610 -130 3620 -60
rect 3640 -130 3650 -60
rect 3610 -140 3650 -130
rect 3690 -60 3730 -50
rect 3690 -130 3700 -60
rect 3720 -130 3730 -60
rect 3690 -140 3730 -130
rect 3755 -60 3795 -50
rect 3755 -130 3765 -60
rect 3785 -130 3795 -60
rect 3755 -140 3795 -130
rect 3835 -60 3875 -50
rect 3835 -130 3845 -60
rect 3865 -130 3875 -60
rect 3835 -140 3875 -130
rect 3900 -60 3945 -50
rect 3900 -130 3910 -60
rect 3930 -130 3945 -60
rect 3900 -140 3945 -130
rect 3980 -60 4020 -50
rect 3980 -130 3990 -60
rect 4010 -130 4020 -60
rect 3980 -140 4020 -130
rect 4045 -60 4085 -50
rect 4045 -130 4055 -60
rect 4075 -130 4085 -60
rect 4045 -140 4085 -130
rect 4125 -60 4165 -50
rect 4125 -130 4135 -60
rect 4155 -130 4165 -60
rect 4125 -140 4165 -130
rect 2775 -175 3355 -160
rect 3845 -175 3865 -140
rect 3895 -170 3935 -160
rect 3895 -175 3905 -170
rect 3925 -175 3935 -170
rect 915 -1155 955 -1145
rect 915 -1165 925 -1155
rect 185 -1175 925 -1165
rect 945 -1165 955 -1155
rect 945 -1175 1325 -1165
rect 185 -1185 1325 -1175
rect -35 -1215 -5 -1205
rect -35 -1235 -30 -1215
rect -10 -1235 -5 -1215
rect -35 -1245 -5 -1235
rect 20 -1215 50 -1205
rect 20 -1235 25 -1215
rect 45 -1235 50 -1215
rect 20 -1245 50 -1235
rect 75 -1215 105 -1205
rect 75 -1235 80 -1215
rect 100 -1235 105 -1215
rect 75 -1245 105 -1235
rect 20 -1325 40 -1245
rect 65 -1275 105 -1265
rect 65 -1295 75 -1275
rect 95 -1285 105 -1275
rect 185 -1285 205 -1185
rect 225 -1215 255 -1205
rect 225 -1235 230 -1215
rect 250 -1235 255 -1215
rect 225 -1245 255 -1235
rect 280 -1215 310 -1205
rect 280 -1235 285 -1215
rect 305 -1235 310 -1215
rect 280 -1245 310 -1235
rect 335 -1215 365 -1205
rect 335 -1235 340 -1215
rect 360 -1235 365 -1215
rect 335 -1245 365 -1235
rect 405 -1215 435 -1205
rect 405 -1235 410 -1215
rect 430 -1235 435 -1215
rect 405 -1245 435 -1235
rect 460 -1215 490 -1205
rect 460 -1235 465 -1215
rect 485 -1235 490 -1215
rect 460 -1245 490 -1235
rect 515 -1215 545 -1205
rect 515 -1235 520 -1215
rect 540 -1235 545 -1215
rect 515 -1245 545 -1235
rect 665 -1215 695 -1205
rect 665 -1235 670 -1215
rect 690 -1235 695 -1215
rect 665 -1245 695 -1235
rect 720 -1215 750 -1205
rect 720 -1235 725 -1215
rect 745 -1235 750 -1215
rect 720 -1245 750 -1235
rect 775 -1215 805 -1205
rect 775 -1235 780 -1215
rect 800 -1235 805 -1215
rect 775 -1245 805 -1235
rect 905 -1215 935 -1205
rect 905 -1235 910 -1215
rect 930 -1235 935 -1215
rect 905 -1245 935 -1235
rect 960 -1215 990 -1205
rect 960 -1235 965 -1215
rect 985 -1235 990 -1215
rect 960 -1245 990 -1235
rect 1015 -1215 1045 -1205
rect 1015 -1235 1020 -1215
rect 1040 -1235 1045 -1215
rect 1015 -1245 1045 -1235
rect 1085 -1215 1115 -1205
rect 1085 -1235 1090 -1215
rect 1110 -1235 1115 -1215
rect 1085 -1245 1115 -1235
rect 1140 -1215 1170 -1205
rect 1140 -1235 1145 -1215
rect 1165 -1235 1170 -1215
rect 1140 -1245 1170 -1235
rect 1210 -1215 1240 -1205
rect 1210 -1235 1215 -1215
rect 1235 -1235 1240 -1215
rect 1210 -1245 1240 -1235
rect 1265 -1215 1295 -1205
rect 1265 -1235 1270 -1215
rect 1290 -1235 1295 -1215
rect 1265 -1245 1295 -1235
rect 95 -1295 205 -1285
rect 65 -1305 205 -1295
rect 20 -1345 100 -1325
rect 80 -1365 100 -1345
rect -35 -1375 -5 -1365
rect -35 -1445 -30 -1375
rect -10 -1445 -5 -1375
rect -35 -1455 -5 -1445
rect 20 -1375 50 -1365
rect 20 -1445 25 -1375
rect 45 -1445 50 -1375
rect 20 -1455 50 -1445
rect 75 -1375 105 -1365
rect 75 -1445 80 -1375
rect 100 -1430 105 -1375
rect 125 -1425 165 -1415
rect 125 -1430 135 -1425
rect 100 -1445 135 -1430
rect 155 -1445 165 -1425
rect 75 -1455 165 -1445
rect 185 -1435 205 -1305
rect 285 -1325 305 -1245
rect 230 -1345 305 -1325
rect 325 -1315 365 -1305
rect 325 -1335 335 -1315
rect 355 -1325 365 -1315
rect 460 -1325 480 -1245
rect 505 -1275 545 -1265
rect 505 -1295 515 -1275
rect 535 -1285 545 -1275
rect 535 -1295 645 -1285
rect 505 -1305 645 -1295
rect 355 -1335 540 -1325
rect 325 -1345 540 -1335
rect 230 -1365 250 -1345
rect 520 -1365 540 -1345
rect 225 -1375 255 -1365
rect 225 -1435 230 -1375
rect 185 -1445 230 -1435
rect 250 -1445 255 -1375
rect 185 -1455 255 -1445
rect 280 -1375 310 -1365
rect 280 -1445 285 -1375
rect 305 -1445 310 -1375
rect 280 -1455 310 -1445
rect 335 -1375 365 -1365
rect 335 -1445 340 -1375
rect 360 -1445 365 -1375
rect 335 -1455 365 -1445
rect 405 -1375 435 -1365
rect 405 -1445 410 -1375
rect 430 -1445 435 -1375
rect 405 -1455 435 -1445
rect 460 -1375 490 -1365
rect 460 -1445 465 -1375
rect 485 -1445 490 -1375
rect 460 -1455 490 -1445
rect 515 -1375 545 -1365
rect 515 -1445 520 -1375
rect 540 -1430 545 -1375
rect 565 -1425 605 -1415
rect 565 -1430 575 -1425
rect 540 -1445 575 -1430
rect 595 -1445 605 -1425
rect 515 -1455 605 -1445
rect 625 -1435 645 -1305
rect 725 -1325 745 -1245
rect 840 -1280 880 -1270
rect 840 -1300 850 -1280
rect 870 -1300 880 -1280
rect 840 -1310 880 -1300
rect 670 -1345 745 -1325
rect 670 -1365 690 -1345
rect 665 -1375 695 -1365
rect 665 -1435 670 -1375
rect 625 -1445 670 -1435
rect 690 -1445 695 -1375
rect 625 -1455 695 -1445
rect 720 -1375 750 -1365
rect 720 -1445 725 -1375
rect 745 -1445 750 -1375
rect 720 -1455 750 -1445
rect 775 -1375 805 -1365
rect 775 -1445 780 -1375
rect 800 -1445 805 -1375
rect 775 -1455 805 -1445
rect 860 -1645 880 -1310
rect 1020 -1290 1040 -1245
rect 1150 -1290 1170 -1245
rect 1275 -1290 1295 -1245
rect 1020 -1300 1075 -1290
rect 1020 -1320 1045 -1300
rect 1065 -1320 1075 -1300
rect 1020 -1325 1075 -1320
rect 910 -1330 1075 -1325
rect 1150 -1300 1200 -1290
rect 1150 -1320 1170 -1300
rect 1190 -1320 1200 -1300
rect 1150 -1330 1200 -1320
rect 1275 -1300 1345 -1290
rect 1275 -1320 1295 -1300
rect 1315 -1320 1345 -1300
rect 1275 -1330 1345 -1320
rect 910 -1345 1040 -1330
rect 910 -1365 930 -1345
rect 1020 -1365 1040 -1345
rect 1150 -1365 1170 -1330
rect 1275 -1365 1295 -1330
rect 905 -1375 935 -1365
rect 905 -1445 910 -1375
rect 930 -1445 935 -1375
rect 905 -1455 935 -1445
rect 960 -1375 990 -1365
rect 960 -1445 965 -1375
rect 985 -1445 990 -1375
rect 960 -1455 990 -1445
rect 1015 -1375 1045 -1365
rect 1015 -1445 1020 -1375
rect 1040 -1445 1045 -1375
rect 1015 -1455 1045 -1445
rect 1085 -1375 1115 -1365
rect 1085 -1445 1090 -1375
rect 1110 -1445 1115 -1375
rect 1085 -1455 1115 -1445
rect 1140 -1375 1170 -1365
rect 1140 -1445 1145 -1375
rect 1165 -1445 1170 -1375
rect 1140 -1455 1170 -1445
rect 1210 -1375 1240 -1365
rect 1210 -1445 1215 -1375
rect 1235 -1445 1240 -1375
rect 1210 -1455 1240 -1445
rect 1265 -1375 1295 -1365
rect 1265 -1445 1270 -1375
rect 1290 -1445 1295 -1375
rect 1265 -1455 1295 -1445
rect 995 -1485 1035 -1475
rect 995 -1505 1005 -1485
rect 1025 -1505 1035 -1485
rect 995 -1515 1035 -1505
rect 860 -1655 900 -1645
rect 860 -1675 870 -1655
rect 890 -1675 900 -1655
rect 860 -1685 900 -1675
rect 995 -1705 1015 -1515
rect 185 -1725 1015 -1705
rect 185 -1745 205 -1725
rect -35 -1755 -5 -1745
rect -35 -1825 -30 -1755
rect -10 -1825 -5 -1755
rect -35 -1835 -5 -1825
rect 20 -1755 50 -1745
rect 20 -1825 25 -1755
rect 45 -1825 50 -1755
rect 20 -1835 50 -1825
rect 75 -1755 165 -1745
rect 75 -1825 80 -1755
rect 100 -1770 135 -1755
rect 100 -1825 105 -1770
rect 125 -1775 135 -1770
rect 155 -1775 165 -1755
rect 125 -1785 165 -1775
rect 185 -1755 255 -1745
rect 185 -1765 230 -1755
rect 75 -1835 105 -1825
rect 80 -1855 100 -1835
rect 20 -1875 100 -1855
rect 20 -1955 40 -1875
rect 185 -1895 205 -1765
rect 225 -1825 230 -1765
rect 250 -1825 255 -1755
rect 225 -1835 255 -1825
rect 280 -1755 310 -1745
rect 280 -1825 285 -1755
rect 305 -1825 310 -1755
rect 280 -1835 310 -1825
rect 335 -1755 365 -1745
rect 335 -1825 340 -1755
rect 360 -1825 365 -1755
rect 335 -1835 365 -1825
rect 405 -1755 435 -1745
rect 405 -1825 410 -1755
rect 430 -1825 435 -1755
rect 405 -1835 435 -1825
rect 460 -1755 490 -1745
rect 460 -1825 465 -1755
rect 485 -1825 490 -1755
rect 460 -1835 490 -1825
rect 515 -1755 605 -1745
rect 515 -1825 520 -1755
rect 540 -1770 575 -1755
rect 540 -1825 545 -1770
rect 565 -1775 575 -1770
rect 595 -1775 605 -1755
rect 565 -1785 605 -1775
rect 625 -1755 695 -1745
rect 625 -1765 670 -1755
rect 515 -1835 545 -1825
rect 230 -1855 250 -1835
rect 520 -1855 540 -1835
rect 230 -1875 305 -1855
rect 65 -1905 205 -1895
rect 65 -1925 75 -1905
rect 95 -1915 205 -1905
rect 95 -1925 105 -1915
rect 65 -1935 105 -1925
rect 285 -1955 305 -1875
rect 325 -1865 540 -1855
rect 325 -1885 335 -1865
rect 355 -1875 540 -1865
rect 355 -1885 365 -1875
rect 325 -1895 365 -1885
rect 460 -1955 480 -1875
rect 625 -1895 645 -1765
rect 665 -1825 670 -1765
rect 690 -1825 695 -1755
rect 665 -1835 695 -1825
rect 720 -1755 750 -1745
rect 720 -1825 725 -1755
rect 745 -1825 750 -1755
rect 720 -1835 750 -1825
rect 775 -1755 805 -1745
rect 775 -1825 780 -1755
rect 800 -1825 805 -1755
rect 775 -1835 805 -1825
rect 955 -1755 985 -1745
rect 955 -1825 960 -1755
rect 980 -1825 985 -1755
rect 955 -1835 985 -1825
rect 1010 -1755 1040 -1745
rect 1010 -1825 1015 -1755
rect 1035 -1825 1040 -1755
rect 1010 -1835 1040 -1825
rect 1080 -1755 1110 -1745
rect 1080 -1825 1085 -1755
rect 1105 -1825 1110 -1755
rect 1080 -1835 1110 -1825
rect 1135 -1755 1165 -1745
rect 1135 -1825 1140 -1755
rect 1160 -1825 1165 -1755
rect 1135 -1835 1165 -1825
rect 1205 -1755 1235 -1745
rect 1205 -1825 1210 -1755
rect 1230 -1825 1235 -1755
rect 1205 -1835 1235 -1825
rect 1260 -1755 1290 -1745
rect 1260 -1825 1265 -1755
rect 1285 -1825 1290 -1755
rect 1260 -1835 1290 -1825
rect 670 -1855 690 -1835
rect 670 -1875 745 -1855
rect 955 -1870 975 -1835
rect 1080 -1870 1100 -1835
rect 1205 -1870 1225 -1835
rect 1325 -1870 1345 -1330
rect 505 -1905 645 -1895
rect 505 -1925 515 -1905
rect 535 -1915 645 -1905
rect 535 -1925 545 -1915
rect 505 -1935 545 -1925
rect 725 -1955 745 -1875
rect 925 -1880 975 -1870
rect 925 -1900 935 -1880
rect 955 -1900 975 -1880
rect 925 -1910 975 -1900
rect 1050 -1880 1100 -1870
rect 1050 -1900 1060 -1880
rect 1080 -1900 1100 -1880
rect 1050 -1910 1100 -1900
rect 1175 -1880 1225 -1870
rect 1175 -1900 1185 -1880
rect 1205 -1900 1225 -1880
rect 1175 -1910 1225 -1900
rect 1305 -1880 1345 -1870
rect 1305 -1900 1315 -1880
rect 1335 -1900 1345 -1880
rect 1305 -1910 1345 -1900
rect 955 -1955 975 -1910
rect 1080 -1955 1100 -1910
rect 1205 -1955 1225 -1910
rect -35 -1965 -5 -1955
rect -35 -1985 -30 -1965
rect -10 -1985 -5 -1965
rect -35 -1995 -5 -1985
rect 20 -1965 50 -1955
rect 20 -1985 25 -1965
rect 45 -1985 50 -1965
rect 20 -1995 50 -1985
rect 75 -1965 105 -1955
rect 75 -1985 80 -1965
rect 100 -1985 105 -1965
rect 75 -1995 105 -1985
rect 225 -1965 255 -1955
rect 225 -1985 230 -1965
rect 250 -1985 255 -1965
rect 225 -1995 255 -1985
rect 280 -1965 310 -1955
rect 280 -1985 285 -1965
rect 305 -1985 310 -1965
rect 280 -1995 310 -1985
rect 335 -1965 365 -1955
rect 335 -1985 340 -1965
rect 360 -1985 365 -1965
rect 335 -1995 365 -1985
rect 405 -1965 435 -1955
rect 405 -1985 410 -1965
rect 430 -1985 435 -1965
rect 405 -1995 435 -1985
rect 460 -1965 490 -1955
rect 460 -1985 465 -1965
rect 485 -1985 490 -1965
rect 460 -1995 490 -1985
rect 515 -1965 545 -1955
rect 515 -1985 520 -1965
rect 540 -1985 545 -1965
rect 515 -1995 545 -1985
rect 665 -1965 695 -1955
rect 665 -1985 670 -1965
rect 690 -1985 695 -1965
rect 665 -1995 695 -1985
rect 720 -1965 750 -1955
rect 720 -1985 725 -1965
rect 745 -1985 750 -1965
rect 720 -1995 750 -1985
rect 775 -1965 805 -1955
rect 775 -1985 780 -1965
rect 800 -1985 805 -1965
rect 775 -1995 805 -1985
rect 955 -1965 985 -1955
rect 955 -1985 960 -1965
rect 980 -1985 985 -1965
rect 955 -1995 985 -1985
rect 1010 -1965 1040 -1955
rect 1010 -1985 1015 -1965
rect 1035 -1985 1040 -1965
rect 1010 -1995 1040 -1985
rect 1080 -1965 1110 -1955
rect 1080 -1985 1085 -1965
rect 1105 -1985 1110 -1965
rect 1080 -1995 1110 -1985
rect 1135 -1965 1165 -1955
rect 1135 -1985 1140 -1965
rect 1160 -1985 1165 -1965
rect 1135 -1995 1165 -1985
rect 1205 -1965 1235 -1955
rect 1205 -1985 1210 -1965
rect 1230 -1985 1235 -1965
rect 1205 -1995 1235 -1985
rect 1260 -1965 1290 -1955
rect 1260 -1985 1265 -1965
rect 1285 -1985 1290 -1965
rect 1260 -1995 1290 -1985
rect 935 -2035 1300 -2015
rect -190 -2570 -170 -2550
rect -150 -2570 -120 -2550
rect -100 -2570 -70 -2550
rect -50 -2570 -20 -2550
rect 0 -2570 30 -2550
rect 50 -2570 80 -2550
rect 100 -2570 130 -2550
rect 150 -2570 180 -2550
rect 200 -2570 230 -2550
rect 250 -2570 280 -2550
rect 300 -2570 340 -2550
rect 360 -2570 390 -2550
rect 410 -2570 440 -2550
rect 460 -2570 490 -2550
rect 510 -2570 540 -2550
rect 560 -2570 590 -2550
rect 610 -2570 640 -2550
rect 660 -2570 690 -2550
rect 710 -2570 740 -2550
rect 760 -2570 790 -2550
rect 810 -2570 840 -2550
rect 860 -2570 890 -2550
rect 910 -2570 980 -2550
rect 1000 -2570 1030 -2550
rect 1050 -2570 1080 -2550
rect 1100 -2570 1170 -2550
rect 1190 -2570 1220 -2550
rect 1240 -2570 1270 -2550
rect 1290 -2570 1350 -2550
rect 1450 -2570 1470 -2550
rect 1490 -2570 1520 -2550
rect 1540 -2570 1570 -2550
rect 1590 -2570 1620 -2550
rect 1640 -2570 1670 -2550
rect 1690 -2570 1720 -2550
rect 1740 -2570 1770 -2550
rect 1790 -2570 1820 -2550
rect 1840 -2570 1870 -2550
rect 1890 -2570 1920 -2550
rect 1940 -2570 1970 -2550
rect 1990 -2570 2020 -2550
rect 2040 -2570 2070 -2550
rect 2090 -2570 2120 -2550
rect 2140 -2570 2170 -2550
rect 2190 -2570 2220 -2550
rect 2240 -2570 2270 -2550
rect -120 -2655 -100 -2570
rect -10 -2655 10 -2570
rect 75 -2605 115 -2595
rect 75 -2625 85 -2605
rect 105 -2625 115 -2605
rect 75 -2635 115 -2625
rect -125 -2665 -95 -2655
rect -125 -2735 -120 -2665
rect -100 -2735 -95 -2665
rect -125 -2745 -95 -2735
rect -70 -2665 -40 -2655
rect -70 -2735 -65 -2665
rect -45 -2735 -40 -2665
rect -70 -2745 -40 -2735
rect -15 -2665 15 -2655
rect -15 -2735 -10 -2665
rect 10 -2735 15 -2665
rect -15 -2745 15 -2735
rect -70 -2825 -50 -2745
rect -25 -2775 15 -2765
rect -25 -2795 -15 -2775
rect 5 -2785 15 -2775
rect 95 -2785 115 -2635
rect 140 -2655 160 -2570
rect 250 -2655 270 -2570
rect 330 -2655 350 -2570
rect 440 -2655 460 -2570
rect 590 -2655 610 -2570
rect 700 -2655 720 -2570
rect 795 -2655 815 -2570
rect 880 -2605 920 -2595
rect 880 -2625 890 -2605
rect 910 -2625 920 -2605
rect 880 -2635 920 -2625
rect 1180 -2655 1200 -2570
rect 1530 -2655 1550 -2570
rect 1675 -2655 1695 -2570
rect 1820 -2655 1840 -2570
rect 135 -2665 165 -2655
rect 135 -2735 140 -2665
rect 160 -2735 165 -2665
rect 135 -2745 165 -2735
rect 190 -2665 220 -2655
rect 190 -2735 195 -2665
rect 215 -2735 220 -2665
rect 190 -2745 220 -2735
rect 245 -2665 275 -2655
rect 245 -2735 250 -2665
rect 270 -2735 275 -2665
rect 245 -2745 275 -2735
rect 325 -2665 355 -2655
rect 325 -2735 330 -2665
rect 350 -2735 355 -2665
rect 325 -2745 355 -2735
rect 380 -2665 410 -2655
rect 380 -2735 385 -2665
rect 405 -2735 410 -2665
rect 380 -2745 410 -2735
rect 435 -2665 465 -2655
rect 435 -2735 440 -2665
rect 460 -2735 465 -2665
rect 435 -2745 465 -2735
rect 585 -2665 615 -2655
rect 585 -2735 590 -2665
rect 610 -2735 615 -2665
rect 585 -2745 615 -2735
rect 640 -2665 670 -2655
rect 640 -2735 645 -2665
rect 665 -2735 670 -2665
rect 640 -2745 670 -2735
rect 695 -2665 725 -2655
rect 695 -2735 700 -2665
rect 720 -2735 725 -2665
rect 695 -2745 725 -2735
rect 790 -2665 820 -2655
rect 790 -2735 795 -2665
rect 815 -2735 820 -2665
rect 790 -2745 820 -2735
rect 845 -2665 875 -2655
rect 845 -2735 850 -2665
rect 870 -2735 875 -2665
rect 845 -2745 875 -2735
rect 900 -2665 930 -2655
rect 900 -2735 905 -2665
rect 925 -2735 930 -2665
rect 900 -2745 930 -2735
rect 1010 -2665 1040 -2655
rect 1010 -2735 1015 -2665
rect 1035 -2735 1040 -2665
rect 1010 -2745 1040 -2735
rect 1065 -2665 1095 -2655
rect 1065 -2735 1070 -2665
rect 1090 -2735 1095 -2665
rect 1065 -2745 1095 -2735
rect 1175 -2665 1205 -2655
rect 1175 -2735 1180 -2665
rect 1200 -2735 1205 -2665
rect 1175 -2745 1205 -2735
rect 1230 -2665 1260 -2655
rect 1230 -2735 1235 -2665
rect 1255 -2735 1260 -2665
rect 1230 -2745 1260 -2735
rect 1520 -2665 1560 -2655
rect 1520 -2685 1530 -2665
rect 1550 -2685 1560 -2665
rect 1520 -2715 1560 -2685
rect 1520 -2735 1530 -2715
rect 1550 -2735 1560 -2715
rect 1520 -2745 1560 -2735
rect 1585 -2665 1625 -2655
rect 1585 -2685 1595 -2665
rect 1615 -2685 1625 -2665
rect 1585 -2715 1625 -2685
rect 1585 -2735 1595 -2715
rect 1615 -2735 1625 -2715
rect 1585 -2745 1625 -2735
rect 1665 -2665 1705 -2655
rect 1665 -2685 1675 -2665
rect 1695 -2685 1705 -2665
rect 1665 -2715 1705 -2685
rect 1665 -2735 1675 -2715
rect 1695 -2735 1705 -2715
rect 1665 -2745 1705 -2735
rect 1730 -2665 1770 -2655
rect 1730 -2685 1740 -2665
rect 1760 -2685 1770 -2665
rect 1730 -2715 1770 -2685
rect 1730 -2735 1740 -2715
rect 1760 -2735 1770 -2715
rect 1730 -2745 1770 -2735
rect 1810 -2665 1850 -2655
rect 1810 -2685 1820 -2665
rect 1840 -2685 1850 -2665
rect 1810 -2715 1850 -2685
rect 1810 -2735 1820 -2715
rect 1840 -2735 1850 -2715
rect 1810 -2745 1850 -2735
rect 1875 -2665 1915 -2655
rect 1875 -2685 1885 -2665
rect 1905 -2685 1915 -2665
rect 1875 -2715 1915 -2685
rect 1875 -2735 1885 -2715
rect 1905 -2735 1915 -2715
rect 1875 -2745 1915 -2735
rect 1955 -2665 1995 -2655
rect 1955 -2685 1965 -2665
rect 1985 -2685 1995 -2665
rect 1955 -2715 1995 -2685
rect 1955 -2735 1965 -2715
rect 1985 -2735 1995 -2715
rect 1955 -2745 1995 -2735
rect 2020 -2665 2060 -2655
rect 2020 -2685 2030 -2665
rect 2050 -2685 2060 -2665
rect 2020 -2715 2060 -2685
rect 2020 -2735 2030 -2715
rect 2050 -2735 2060 -2715
rect 2020 -2745 2060 -2735
rect 5 -2795 115 -2785
rect -25 -2805 115 -2795
rect -70 -2845 10 -2825
rect -10 -2865 10 -2845
rect -125 -2875 -95 -2865
rect -125 -2895 -120 -2875
rect -100 -2895 -95 -2875
rect -125 -2925 -95 -2895
rect -125 -2945 -120 -2925
rect -100 -2945 -95 -2925
rect -125 -2975 -95 -2945
rect -125 -2995 -120 -2975
rect -100 -2995 -95 -2975
rect -125 -3025 -95 -2995
rect -125 -3045 -120 -3025
rect -100 -3045 -95 -3025
rect -125 -3055 -95 -3045
rect -70 -2875 -40 -2865
rect -70 -2895 -65 -2875
rect -45 -2895 -40 -2875
rect -70 -2925 -40 -2895
rect -70 -2945 -65 -2925
rect -45 -2945 -40 -2925
rect -70 -2975 -40 -2945
rect -70 -2995 -65 -2975
rect -45 -2995 -40 -2975
rect -70 -3025 -40 -2995
rect -70 -3045 -65 -3025
rect -45 -3045 -40 -3025
rect -70 -3055 -40 -3045
rect -15 -2875 15 -2865
rect -15 -2895 -10 -2875
rect 10 -2895 15 -2875
rect -15 -2925 15 -2895
rect -15 -2945 -10 -2925
rect 10 -2945 15 -2925
rect -15 -2975 15 -2945
rect -15 -2995 -10 -2975
rect 10 -2995 15 -2975
rect -15 -3025 15 -2995
rect -15 -3045 -10 -3025
rect 10 -3030 15 -3025
rect 35 -3025 75 -3015
rect 35 -3030 45 -3025
rect 10 -3045 45 -3030
rect 65 -3045 75 -3025
rect -15 -3055 75 -3045
rect 95 -3035 115 -2805
rect 195 -2825 215 -2745
rect 140 -2845 215 -2825
rect 235 -2815 275 -2805
rect 235 -2835 245 -2815
rect 265 -2825 275 -2815
rect 380 -2825 400 -2745
rect 425 -2775 465 -2765
rect 425 -2795 435 -2775
rect 455 -2785 465 -2775
rect 455 -2795 565 -2785
rect 425 -2805 565 -2795
rect 265 -2835 460 -2825
rect 235 -2845 460 -2835
rect 140 -2865 160 -2845
rect 440 -2865 460 -2845
rect 135 -2875 165 -2865
rect 135 -2895 140 -2875
rect 160 -2895 165 -2875
rect 135 -2925 165 -2895
rect 135 -2945 140 -2925
rect 160 -2945 165 -2925
rect 135 -2975 165 -2945
rect 135 -2995 140 -2975
rect 160 -2995 165 -2975
rect 135 -3025 165 -2995
rect 135 -3035 140 -3025
rect 95 -3045 140 -3035
rect 160 -3045 165 -3025
rect 95 -3055 165 -3045
rect 190 -2875 220 -2865
rect 190 -2895 195 -2875
rect 215 -2895 220 -2875
rect 190 -2925 220 -2895
rect 190 -2945 195 -2925
rect 215 -2945 220 -2925
rect 190 -2975 220 -2945
rect 190 -2995 195 -2975
rect 215 -2995 220 -2975
rect 190 -3025 220 -2995
rect 190 -3045 195 -3025
rect 215 -3045 220 -3025
rect 190 -3055 220 -3045
rect 245 -2875 275 -2865
rect 245 -2895 250 -2875
rect 270 -2895 275 -2875
rect 245 -2925 275 -2895
rect 245 -2945 250 -2925
rect 270 -2945 275 -2925
rect 245 -2975 275 -2945
rect 245 -2995 250 -2975
rect 270 -2995 275 -2975
rect 245 -3025 275 -2995
rect 245 -3045 250 -3025
rect 270 -3045 275 -3025
rect 245 -3055 275 -3045
rect 325 -2875 355 -2865
rect 325 -2895 330 -2875
rect 350 -2895 355 -2875
rect 325 -2925 355 -2895
rect 325 -2945 330 -2925
rect 350 -2945 355 -2925
rect 325 -2975 355 -2945
rect 325 -2995 330 -2975
rect 350 -2995 355 -2975
rect 325 -3025 355 -2995
rect 325 -3045 330 -3025
rect 350 -3045 355 -3025
rect 325 -3055 355 -3045
rect 380 -2875 410 -2865
rect 380 -2895 385 -2875
rect 405 -2895 410 -2875
rect 380 -2925 410 -2895
rect 380 -2945 385 -2925
rect 405 -2945 410 -2925
rect 380 -2975 410 -2945
rect 380 -2995 385 -2975
rect 405 -2995 410 -2975
rect 380 -3025 410 -2995
rect 380 -3045 385 -3025
rect 405 -3045 410 -3025
rect 380 -3055 410 -3045
rect 435 -2875 465 -2865
rect 435 -2895 440 -2875
rect 460 -2895 465 -2875
rect 435 -2925 465 -2895
rect 435 -2945 440 -2925
rect 460 -2945 465 -2925
rect 435 -2975 465 -2945
rect 435 -2995 440 -2975
rect 460 -2995 465 -2975
rect 435 -3025 465 -2995
rect 435 -3045 440 -3025
rect 460 -3030 465 -3025
rect 485 -3025 525 -3015
rect 485 -3030 495 -3025
rect 460 -3045 495 -3030
rect 515 -3045 525 -3025
rect 435 -3055 525 -3045
rect 545 -3035 565 -2805
rect 645 -2825 665 -2745
rect 720 -2780 760 -2770
rect 720 -2800 730 -2780
rect 750 -2800 760 -2780
rect 720 -2810 760 -2800
rect 905 -2790 925 -2745
rect 1075 -2790 1095 -2745
rect 1240 -2790 1260 -2745
rect 905 -2800 960 -2790
rect 905 -2820 930 -2800
rect 950 -2820 960 -2800
rect 905 -2825 960 -2820
rect 590 -2845 665 -2825
rect 795 -2830 960 -2825
rect 1075 -2800 1165 -2790
rect 1075 -2820 1095 -2800
rect 1155 -2820 1165 -2800
rect 1075 -2830 1165 -2820
rect 1240 -2800 1290 -2790
rect 1240 -2820 1260 -2800
rect 1280 -2820 1290 -2800
rect 1240 -2830 1290 -2820
rect 1605 -2800 1625 -2745
rect 1685 -2800 1725 -2790
rect 1605 -2820 1695 -2800
rect 1715 -2820 1725 -2800
rect 795 -2845 925 -2830
rect 590 -2865 610 -2845
rect 795 -2865 815 -2845
rect 905 -2865 925 -2845
rect 1075 -2865 1095 -2830
rect 1240 -2865 1260 -2830
rect 1605 -2865 1625 -2820
rect 1685 -2830 1725 -2820
rect 1750 -2800 1770 -2745
rect 1830 -2800 1870 -2790
rect 1750 -2820 1840 -2800
rect 1860 -2820 1870 -2800
rect 1750 -2865 1770 -2820
rect 1830 -2830 1870 -2820
rect 1895 -2805 1915 -2745
rect 1895 -2815 1935 -2805
rect 1895 -2835 1905 -2815
rect 1925 -2835 1935 -2815
rect 1895 -2845 1935 -2835
rect 1895 -2865 1915 -2845
rect 1965 -2865 1985 -2745
rect 2030 -2865 2050 -2745
rect 585 -2875 615 -2865
rect 585 -2895 590 -2875
rect 610 -2895 615 -2875
rect 585 -2925 615 -2895
rect 585 -2945 590 -2925
rect 610 -2945 615 -2925
rect 585 -2975 615 -2945
rect 585 -2995 590 -2975
rect 610 -2995 615 -2975
rect 585 -3025 615 -2995
rect 585 -3035 590 -3025
rect 545 -3045 590 -3035
rect 610 -3045 615 -3025
rect 545 -3055 615 -3045
rect 640 -2875 670 -2865
rect 640 -2895 645 -2875
rect 665 -2895 670 -2875
rect 640 -2925 670 -2895
rect 640 -2945 645 -2925
rect 665 -2945 670 -2925
rect 640 -2975 670 -2945
rect 640 -2995 645 -2975
rect 665 -2995 670 -2975
rect 640 -3025 670 -2995
rect 640 -3045 645 -3025
rect 665 -3045 670 -3025
rect 640 -3055 670 -3045
rect 695 -2875 725 -2865
rect 695 -2895 700 -2875
rect 720 -2895 725 -2875
rect 695 -2925 725 -2895
rect 695 -2945 700 -2925
rect 720 -2945 725 -2925
rect 695 -2975 725 -2945
rect 695 -2995 700 -2975
rect 720 -2995 725 -2975
rect 695 -3025 725 -2995
rect 695 -3045 700 -3025
rect 720 -3045 725 -3025
rect 695 -3055 725 -3045
rect 790 -2875 820 -2865
rect 790 -2895 795 -2875
rect 815 -2895 820 -2875
rect 790 -2925 820 -2895
rect 790 -2945 795 -2925
rect 815 -2945 820 -2925
rect 790 -2975 820 -2945
rect 790 -2995 795 -2975
rect 815 -2995 820 -2975
rect 790 -3025 820 -2995
rect 790 -3045 795 -3025
rect 815 -3045 820 -3025
rect 790 -3055 820 -3045
rect 845 -2875 875 -2865
rect 845 -2895 850 -2875
rect 870 -2895 875 -2875
rect 845 -2925 875 -2895
rect 845 -2945 850 -2925
rect 870 -2945 875 -2925
rect 845 -2975 875 -2945
rect 845 -2995 850 -2975
rect 870 -2995 875 -2975
rect 845 -3025 875 -2995
rect 845 -3045 850 -3025
rect 870 -3045 875 -3025
rect 845 -3055 875 -3045
rect 900 -2875 930 -2865
rect 900 -2895 905 -2875
rect 925 -2895 930 -2875
rect 900 -2925 930 -2895
rect 900 -2945 905 -2925
rect 925 -2945 930 -2925
rect 900 -2975 930 -2945
rect 900 -2995 905 -2975
rect 925 -2995 930 -2975
rect 900 -3025 930 -2995
rect 900 -3045 905 -3025
rect 925 -3045 930 -3025
rect 900 -3055 930 -3045
rect 1010 -2875 1040 -2865
rect 1010 -2895 1015 -2875
rect 1035 -2895 1040 -2875
rect 1010 -2925 1040 -2895
rect 1010 -2945 1015 -2925
rect 1035 -2945 1040 -2925
rect 1010 -2975 1040 -2945
rect 1010 -2995 1015 -2975
rect 1035 -2995 1040 -2975
rect 1010 -3025 1040 -2995
rect 1010 -3045 1015 -3025
rect 1035 -3045 1040 -3025
rect 1010 -3055 1040 -3045
rect 1065 -2875 1095 -2865
rect 1065 -2895 1070 -2875
rect 1090 -2895 1095 -2875
rect 1065 -2925 1095 -2895
rect 1065 -2945 1070 -2925
rect 1090 -2945 1095 -2925
rect 1065 -2975 1095 -2945
rect 1065 -2995 1070 -2975
rect 1090 -2995 1095 -2975
rect 1065 -3025 1095 -2995
rect 1065 -3045 1070 -3025
rect 1090 -3045 1095 -3025
rect 1065 -3055 1095 -3045
rect 1175 -2875 1205 -2865
rect 1175 -2895 1180 -2875
rect 1200 -2895 1205 -2875
rect 1175 -2925 1205 -2895
rect 1175 -2945 1180 -2925
rect 1200 -2945 1205 -2925
rect 1175 -2975 1205 -2945
rect 1175 -2995 1180 -2975
rect 1200 -2995 1205 -2975
rect 1175 -3025 1205 -2995
rect 1175 -3045 1180 -3025
rect 1200 -3045 1205 -3025
rect 1175 -3055 1205 -3045
rect 1230 -2875 1260 -2865
rect 1230 -2895 1235 -2875
rect 1255 -2895 1260 -2875
rect 1230 -2925 1260 -2895
rect 1230 -2945 1235 -2925
rect 1255 -2945 1260 -2925
rect 1230 -2975 1260 -2945
rect 1230 -2995 1235 -2975
rect 1255 -2995 1260 -2975
rect 1230 -3025 1260 -2995
rect 1230 -3045 1235 -3025
rect 1255 -3045 1260 -3025
rect 1230 -3055 1260 -3045
rect 1520 -2875 1560 -2865
rect 1520 -2895 1530 -2875
rect 1550 -2895 1560 -2875
rect 1520 -2925 1560 -2895
rect 1520 -2945 1530 -2925
rect 1550 -2945 1560 -2925
rect 1520 -2975 1560 -2945
rect 1520 -2995 1530 -2975
rect 1550 -2995 1560 -2975
rect 1520 -3025 1560 -2995
rect 1520 -3045 1530 -3025
rect 1550 -3045 1560 -3025
rect 1520 -3055 1560 -3045
rect 1585 -2875 1625 -2865
rect 1585 -2895 1595 -2875
rect 1615 -2895 1625 -2875
rect 1585 -2925 1625 -2895
rect 1585 -2945 1595 -2925
rect 1615 -2945 1625 -2925
rect 1585 -2975 1625 -2945
rect 1585 -2995 1595 -2975
rect 1615 -2995 1625 -2975
rect 1585 -3025 1625 -2995
rect 1585 -3045 1595 -3025
rect 1615 -3045 1625 -3025
rect 1585 -3055 1625 -3045
rect 1665 -2875 1705 -2865
rect 1665 -2895 1675 -2875
rect 1695 -2895 1705 -2875
rect 1665 -2925 1705 -2895
rect 1665 -2945 1675 -2925
rect 1695 -2945 1705 -2925
rect 1665 -2975 1705 -2945
rect 1665 -2995 1675 -2975
rect 1695 -2995 1705 -2975
rect 1665 -3025 1705 -2995
rect 1665 -3045 1675 -3025
rect 1695 -3045 1705 -3025
rect 1665 -3055 1705 -3045
rect 1730 -2875 1770 -2865
rect 1730 -2895 1740 -2875
rect 1760 -2895 1770 -2875
rect 1730 -2925 1770 -2895
rect 1730 -2945 1740 -2925
rect 1760 -2945 1770 -2925
rect 1730 -2975 1770 -2945
rect 1730 -2995 1740 -2975
rect 1760 -2995 1770 -2975
rect 1730 -3025 1770 -2995
rect 1730 -3045 1740 -3025
rect 1760 -3045 1770 -3025
rect 1730 -3055 1770 -3045
rect 1810 -2875 1850 -2865
rect 1810 -2895 1820 -2875
rect 1840 -2895 1850 -2875
rect 1810 -2925 1850 -2895
rect 1810 -2945 1820 -2925
rect 1840 -2945 1850 -2925
rect 1810 -2975 1850 -2945
rect 1810 -2995 1820 -2975
rect 1840 -2995 1850 -2975
rect 1810 -3025 1850 -2995
rect 1810 -3045 1820 -3025
rect 1840 -3045 1850 -3025
rect 1810 -3055 1850 -3045
rect 1875 -2875 1915 -2865
rect 1875 -2895 1885 -2875
rect 1905 -2895 1915 -2875
rect 1875 -2925 1915 -2895
rect 1875 -2945 1885 -2925
rect 1905 -2945 1915 -2925
rect 1875 -2975 1915 -2945
rect 1875 -2995 1885 -2975
rect 1905 -2995 1915 -2975
rect 1875 -3025 1915 -2995
rect 1875 -3045 1885 -3025
rect 1905 -3045 1915 -3025
rect 1875 -3055 1915 -3045
rect 1955 -2875 1995 -2865
rect 1955 -2895 1965 -2875
rect 1985 -2895 1995 -2875
rect 1955 -2925 1995 -2895
rect 1955 -2945 1965 -2925
rect 1985 -2945 1995 -2925
rect 1955 -2975 1995 -2945
rect 1955 -2995 1965 -2975
rect 1985 -2995 1995 -2975
rect 1955 -3025 1995 -2995
rect 1955 -3045 1965 -3025
rect 1985 -3045 1995 -3025
rect 1955 -3055 1995 -3045
rect 2020 -2875 2060 -2865
rect 2020 -2895 2030 -2875
rect 2050 -2895 2060 -2875
rect 2020 -2925 2060 -2895
rect 2020 -2945 2030 -2925
rect 2050 -2945 2060 -2925
rect 2020 -2975 2060 -2945
rect 2020 -2995 2030 -2975
rect 2050 -2995 2060 -2975
rect 2020 -3025 2060 -2995
rect 2020 -3045 2030 -3025
rect 2050 -3045 2060 -3025
rect 2020 -3055 2060 -3045
rect 2100 -2875 2140 -2865
rect 2100 -2895 2110 -2875
rect 2130 -2895 2140 -2875
rect 2100 -2925 2140 -2895
rect 2100 -2945 2110 -2925
rect 2130 -2945 2140 -2925
rect 2100 -2975 2140 -2945
rect 2100 -2995 2110 -2975
rect 2130 -2995 2140 -2975
rect 2100 -3025 2140 -2995
rect 2100 -3045 2110 -3025
rect 2130 -3045 2140 -3025
rect 2100 -3055 2140 -3045
rect 2165 -2875 2205 -2865
rect 2165 -2895 2175 -2875
rect 2195 -2895 2205 -2875
rect 2165 -2925 2205 -2895
rect 2165 -2945 2175 -2925
rect 2195 -2945 2205 -2925
rect 2165 -2975 2205 -2945
rect 2165 -2995 2175 -2975
rect 2195 -2995 2205 -2975
rect 2165 -3025 2205 -2995
rect 2165 -3045 2175 -3025
rect 2195 -3045 2205 -3025
rect 2165 -3055 2205 -3045
rect -120 -3140 -100 -3055
rect 250 -3140 270 -3055
rect 330 -3140 350 -3055
rect 700 -3140 720 -3055
rect 795 -3085 835 -3075
rect 795 -3105 805 -3085
rect 825 -3105 835 -3085
rect 795 -3115 835 -3105
rect 855 -3140 875 -3055
rect 1015 -3140 1035 -3055
rect 1180 -3140 1200 -3055
rect 1530 -3140 1550 -3055
rect 1675 -3140 1695 -3055
rect 1820 -3140 1840 -3055
rect 2110 -3140 2130 -3055
rect -190 -3160 -170 -3140
rect -150 -3160 -120 -3140
rect -100 -3160 -70 -3140
rect -50 -3160 -20 -3140
rect 0 -3160 30 -3140
rect 50 -3160 80 -3140
rect 100 -3160 130 -3140
rect 150 -3160 180 -3140
rect 200 -3160 230 -3140
rect 250 -3160 280 -3140
rect 300 -3160 340 -3140
rect 360 -3160 390 -3140
rect 410 -3160 440 -3140
rect 460 -3160 490 -3140
rect 510 -3160 540 -3140
rect 560 -3160 590 -3140
rect 610 -3160 640 -3140
rect 660 -3160 690 -3140
rect 710 -3160 740 -3140
rect 760 -3160 790 -3140
rect 810 -3160 840 -3140
rect 860 -3160 890 -3140
rect 910 -3160 980 -3140
rect 1000 -3160 1030 -3140
rect 1050 -3160 1080 -3140
rect 1100 -3160 1170 -3140
rect 1190 -3160 1220 -3140
rect 1240 -3160 1270 -3140
rect 1290 -3160 1345 -3140
rect 1450 -3160 1470 -3140
rect 1490 -3160 1520 -3140
rect 1540 -3160 1570 -3140
rect 1590 -3160 1620 -3140
rect 1640 -3160 1670 -3140
rect 1690 -3160 1720 -3140
rect 1740 -3160 1770 -3140
rect 1790 -3160 1820 -3140
rect 1840 -3160 1870 -3140
rect 1890 -3160 1920 -3140
rect 1940 -3160 1970 -3140
rect 1990 -3160 2020 -3140
rect 2040 -3160 2070 -3140
rect 2090 -3160 2120 -3140
rect 2140 -3160 2170 -3140
rect 2190 -3160 2220 -3140
rect 2240 -3160 2270 -3140
rect -120 -3245 -100 -3160
rect 95 -3195 135 -3185
rect 95 -3215 105 -3195
rect 125 -3215 135 -3195
rect 95 -3225 135 -3215
rect 95 -3245 115 -3225
rect 250 -3245 270 -3160
rect 330 -3245 350 -3160
rect 700 -3245 720 -3160
rect 900 -3245 920 -3160
rect 1065 -3245 1085 -3160
rect 1230 -3245 1250 -3160
rect 1595 -3245 1615 -3160
rect 1685 -3195 1725 -3185
rect 1685 -3215 1695 -3195
rect 1715 -3215 1725 -3195
rect 1685 -3225 1725 -3215
rect 1820 -3245 1840 -3160
rect 1975 -3195 2015 -3185
rect 1975 -3215 1985 -3195
rect 2005 -3215 2015 -3195
rect 1975 -3225 2015 -3215
rect -125 -3255 -95 -3245
rect -125 -3275 -120 -3255
rect -100 -3275 -95 -3255
rect -125 -3305 -95 -3275
rect -125 -3325 -120 -3305
rect -100 -3325 -95 -3305
rect -125 -3355 -95 -3325
rect -125 -3375 -120 -3355
rect -100 -3375 -95 -3355
rect -125 -3405 -95 -3375
rect -125 -3425 -120 -3405
rect -100 -3425 -95 -3405
rect -125 -3435 -95 -3425
rect -70 -3255 -40 -3245
rect -70 -3275 -65 -3255
rect -45 -3275 -40 -3255
rect -70 -3305 -40 -3275
rect -70 -3325 -65 -3305
rect -45 -3325 -40 -3305
rect -70 -3355 -40 -3325
rect -70 -3375 -65 -3355
rect -45 -3375 -40 -3355
rect -70 -3405 -40 -3375
rect -70 -3425 -65 -3405
rect -45 -3425 -40 -3405
rect -70 -3435 -40 -3425
rect -15 -3255 75 -3245
rect -15 -3275 -10 -3255
rect 10 -3270 45 -3255
rect 10 -3275 15 -3270
rect -15 -3305 15 -3275
rect 35 -3275 45 -3270
rect 65 -3275 75 -3255
rect 35 -3285 75 -3275
rect 95 -3255 165 -3245
rect 95 -3265 140 -3255
rect -15 -3325 -10 -3305
rect 10 -3325 15 -3305
rect -15 -3355 15 -3325
rect -15 -3375 -10 -3355
rect 10 -3375 15 -3355
rect -15 -3405 15 -3375
rect -15 -3425 -10 -3405
rect 10 -3425 15 -3405
rect -15 -3435 15 -3425
rect -10 -3455 10 -3435
rect -70 -3475 10 -3455
rect -70 -3555 -50 -3475
rect 95 -3495 115 -3265
rect 135 -3275 140 -3265
rect 160 -3275 165 -3255
rect 135 -3305 165 -3275
rect 135 -3325 140 -3305
rect 160 -3325 165 -3305
rect 135 -3355 165 -3325
rect 135 -3375 140 -3355
rect 160 -3375 165 -3355
rect 135 -3405 165 -3375
rect 135 -3425 140 -3405
rect 160 -3425 165 -3405
rect 135 -3435 165 -3425
rect 190 -3255 220 -3245
rect 190 -3275 195 -3255
rect 215 -3275 220 -3255
rect 190 -3305 220 -3275
rect 190 -3325 195 -3305
rect 215 -3325 220 -3305
rect 190 -3355 220 -3325
rect 190 -3375 195 -3355
rect 215 -3375 220 -3355
rect 190 -3405 220 -3375
rect 190 -3425 195 -3405
rect 215 -3425 220 -3405
rect 190 -3435 220 -3425
rect 245 -3255 275 -3245
rect 245 -3275 250 -3255
rect 270 -3275 275 -3255
rect 245 -3305 275 -3275
rect 245 -3325 250 -3305
rect 270 -3325 275 -3305
rect 245 -3355 275 -3325
rect 245 -3375 250 -3355
rect 270 -3375 275 -3355
rect 245 -3405 275 -3375
rect 245 -3425 250 -3405
rect 270 -3425 275 -3405
rect 245 -3435 275 -3425
rect 325 -3255 355 -3245
rect 325 -3275 330 -3255
rect 350 -3275 355 -3255
rect 325 -3305 355 -3275
rect 325 -3325 330 -3305
rect 350 -3325 355 -3305
rect 325 -3355 355 -3325
rect 325 -3375 330 -3355
rect 350 -3375 355 -3355
rect 325 -3405 355 -3375
rect 325 -3425 330 -3405
rect 350 -3425 355 -3405
rect 325 -3435 355 -3425
rect 380 -3255 410 -3245
rect 380 -3275 385 -3255
rect 405 -3275 410 -3255
rect 380 -3305 410 -3275
rect 380 -3325 385 -3305
rect 405 -3325 410 -3305
rect 380 -3355 410 -3325
rect 380 -3375 385 -3355
rect 405 -3375 410 -3355
rect 380 -3405 410 -3375
rect 380 -3425 385 -3405
rect 405 -3425 410 -3405
rect 380 -3435 410 -3425
rect 435 -3255 525 -3245
rect 435 -3275 440 -3255
rect 460 -3270 495 -3255
rect 460 -3275 465 -3270
rect 435 -3305 465 -3275
rect 485 -3275 495 -3270
rect 515 -3275 525 -3255
rect 485 -3285 525 -3275
rect 545 -3255 615 -3245
rect 545 -3265 590 -3255
rect 435 -3325 440 -3305
rect 460 -3325 465 -3305
rect 435 -3355 465 -3325
rect 435 -3375 440 -3355
rect 460 -3375 465 -3355
rect 435 -3405 465 -3375
rect 435 -3425 440 -3405
rect 460 -3425 465 -3405
rect 435 -3435 465 -3425
rect 140 -3455 160 -3435
rect 440 -3455 460 -3435
rect 140 -3475 215 -3455
rect -25 -3505 115 -3495
rect -25 -3525 -15 -3505
rect 5 -3515 115 -3505
rect 5 -3525 15 -3515
rect -25 -3535 15 -3525
rect 195 -3555 215 -3475
rect 235 -3465 460 -3455
rect 235 -3485 245 -3465
rect 265 -3475 460 -3465
rect 265 -3485 275 -3475
rect 235 -3495 275 -3485
rect 380 -3555 400 -3475
rect 545 -3495 565 -3265
rect 585 -3275 590 -3265
rect 610 -3275 615 -3255
rect 585 -3305 615 -3275
rect 585 -3325 590 -3305
rect 610 -3325 615 -3305
rect 585 -3355 615 -3325
rect 585 -3375 590 -3355
rect 610 -3375 615 -3355
rect 585 -3405 615 -3375
rect 585 -3425 590 -3405
rect 610 -3425 615 -3405
rect 585 -3435 615 -3425
rect 640 -3255 670 -3245
rect 640 -3275 645 -3255
rect 665 -3275 670 -3255
rect 640 -3305 670 -3275
rect 640 -3325 645 -3305
rect 665 -3325 670 -3305
rect 640 -3355 670 -3325
rect 640 -3375 645 -3355
rect 665 -3375 670 -3355
rect 640 -3405 670 -3375
rect 640 -3425 645 -3405
rect 665 -3425 670 -3405
rect 640 -3435 670 -3425
rect 695 -3255 725 -3245
rect 695 -3275 700 -3255
rect 720 -3275 725 -3255
rect 695 -3305 725 -3275
rect 695 -3325 700 -3305
rect 720 -3325 725 -3305
rect 695 -3355 725 -3325
rect 695 -3375 700 -3355
rect 720 -3375 725 -3355
rect 695 -3405 725 -3375
rect 695 -3425 700 -3405
rect 720 -3425 725 -3405
rect 695 -3435 725 -3425
rect 840 -3255 870 -3245
rect 840 -3275 845 -3255
rect 865 -3275 870 -3255
rect 840 -3305 870 -3275
rect 840 -3325 845 -3305
rect 865 -3325 870 -3305
rect 840 -3355 870 -3325
rect 840 -3375 845 -3355
rect 865 -3375 870 -3355
rect 840 -3405 870 -3375
rect 840 -3425 845 -3405
rect 865 -3425 870 -3405
rect 840 -3435 870 -3425
rect 895 -3255 925 -3245
rect 895 -3275 900 -3255
rect 920 -3275 925 -3255
rect 895 -3305 925 -3275
rect 895 -3325 900 -3305
rect 920 -3325 925 -3305
rect 895 -3355 925 -3325
rect 895 -3375 900 -3355
rect 920 -3375 925 -3355
rect 895 -3405 925 -3375
rect 895 -3425 900 -3405
rect 920 -3425 925 -3405
rect 895 -3435 925 -3425
rect 1005 -3255 1035 -3245
rect 1005 -3275 1010 -3255
rect 1030 -3275 1035 -3255
rect 1005 -3305 1035 -3275
rect 1005 -3325 1010 -3305
rect 1030 -3325 1035 -3305
rect 1005 -3355 1035 -3325
rect 1005 -3375 1010 -3355
rect 1030 -3375 1035 -3355
rect 1005 -3405 1035 -3375
rect 1005 -3425 1010 -3405
rect 1030 -3425 1035 -3405
rect 1005 -3435 1035 -3425
rect 1060 -3255 1090 -3245
rect 1060 -3275 1065 -3255
rect 1085 -3275 1090 -3255
rect 1060 -3305 1090 -3275
rect 1060 -3325 1065 -3305
rect 1085 -3325 1090 -3305
rect 1060 -3355 1090 -3325
rect 1060 -3375 1065 -3355
rect 1085 -3375 1090 -3355
rect 1060 -3405 1090 -3375
rect 1060 -3425 1065 -3405
rect 1085 -3425 1090 -3405
rect 1060 -3435 1090 -3425
rect 1170 -3255 1200 -3245
rect 1170 -3275 1175 -3255
rect 1195 -3275 1200 -3255
rect 1170 -3305 1200 -3275
rect 1170 -3325 1175 -3305
rect 1195 -3325 1200 -3305
rect 1170 -3355 1200 -3325
rect 1170 -3375 1175 -3355
rect 1195 -3375 1200 -3355
rect 1170 -3405 1200 -3375
rect 1170 -3425 1175 -3405
rect 1195 -3425 1200 -3405
rect 1170 -3435 1200 -3425
rect 1225 -3255 1255 -3245
rect 1225 -3275 1230 -3255
rect 1250 -3275 1255 -3255
rect 1225 -3305 1255 -3275
rect 1225 -3325 1230 -3305
rect 1250 -3325 1255 -3305
rect 1225 -3355 1255 -3325
rect 1225 -3375 1230 -3355
rect 1250 -3375 1255 -3355
rect 1225 -3405 1255 -3375
rect 1225 -3425 1230 -3405
rect 1250 -3425 1255 -3405
rect 1225 -3435 1255 -3425
rect 1520 -3255 1560 -3245
rect 1520 -3275 1530 -3255
rect 1550 -3275 1560 -3255
rect 1520 -3305 1560 -3275
rect 1520 -3325 1530 -3305
rect 1550 -3325 1560 -3305
rect 1520 -3355 1560 -3325
rect 1520 -3375 1530 -3355
rect 1550 -3375 1560 -3355
rect 1520 -3405 1560 -3375
rect 1520 -3425 1530 -3405
rect 1550 -3425 1560 -3405
rect 1520 -3435 1560 -3425
rect 1585 -3255 1625 -3245
rect 1585 -3275 1595 -3255
rect 1615 -3275 1625 -3255
rect 1585 -3305 1625 -3275
rect 1585 -3325 1595 -3305
rect 1615 -3325 1625 -3305
rect 1585 -3355 1625 -3325
rect 1585 -3375 1595 -3355
rect 1615 -3375 1625 -3355
rect 1585 -3405 1625 -3375
rect 1585 -3425 1595 -3405
rect 1615 -3425 1625 -3405
rect 1585 -3435 1625 -3425
rect 1665 -3255 1705 -3245
rect 1665 -3275 1675 -3255
rect 1695 -3275 1705 -3255
rect 1665 -3305 1705 -3275
rect 1665 -3325 1675 -3305
rect 1695 -3325 1705 -3305
rect 1665 -3355 1705 -3325
rect 1665 -3375 1675 -3355
rect 1695 -3375 1705 -3355
rect 1665 -3405 1705 -3375
rect 1665 -3425 1675 -3405
rect 1695 -3425 1705 -3405
rect 1665 -3435 1705 -3425
rect 1730 -3255 1770 -3245
rect 1730 -3275 1740 -3255
rect 1760 -3275 1770 -3255
rect 1730 -3305 1770 -3275
rect 1730 -3325 1740 -3305
rect 1760 -3325 1770 -3305
rect 1730 -3355 1770 -3325
rect 1730 -3375 1740 -3355
rect 1760 -3375 1770 -3355
rect 1730 -3405 1770 -3375
rect 1730 -3425 1740 -3405
rect 1760 -3425 1770 -3405
rect 1730 -3435 1770 -3425
rect 1810 -3255 1850 -3245
rect 1810 -3275 1820 -3255
rect 1840 -3275 1850 -3255
rect 1810 -3305 1850 -3275
rect 1810 -3325 1820 -3305
rect 1840 -3325 1850 -3305
rect 1810 -3355 1850 -3325
rect 1810 -3375 1820 -3355
rect 1840 -3375 1850 -3355
rect 1810 -3405 1850 -3375
rect 1810 -3425 1820 -3405
rect 1840 -3425 1850 -3405
rect 1810 -3435 1850 -3425
rect 1875 -3255 1915 -3245
rect 1875 -3275 1885 -3255
rect 1905 -3275 1915 -3255
rect 1875 -3305 1915 -3275
rect 1875 -3325 1885 -3305
rect 1905 -3325 1915 -3305
rect 1875 -3355 1915 -3325
rect 1875 -3375 1885 -3355
rect 1905 -3375 1915 -3355
rect 1875 -3405 1915 -3375
rect 1875 -3425 1885 -3405
rect 1905 -3425 1915 -3405
rect 1875 -3435 1915 -3425
rect 1955 -3255 1995 -3245
rect 1955 -3275 1965 -3255
rect 1985 -3275 1995 -3255
rect 1955 -3305 1995 -3275
rect 1955 -3325 1965 -3305
rect 1985 -3325 1995 -3305
rect 1955 -3355 1995 -3325
rect 1955 -3375 1965 -3355
rect 1985 -3375 1995 -3355
rect 1955 -3405 1995 -3375
rect 1955 -3425 1965 -3405
rect 1985 -3425 1995 -3405
rect 1955 -3435 1995 -3425
rect 2020 -3255 2060 -3245
rect 2020 -3275 2030 -3255
rect 2050 -3275 2060 -3255
rect 2020 -3305 2060 -3275
rect 2020 -3325 2030 -3305
rect 2050 -3325 2060 -3305
rect 2020 -3355 2060 -3325
rect 2020 -3375 2030 -3355
rect 2050 -3375 2060 -3355
rect 2020 -3405 2060 -3375
rect 2020 -3425 2030 -3405
rect 2050 -3425 2060 -3405
rect 2020 -3435 2060 -3425
rect 590 -3455 610 -3435
rect 590 -3475 665 -3455
rect 840 -3470 860 -3435
rect 1005 -3470 1025 -3435
rect 1170 -3470 1190 -3435
rect 1595 -3455 1615 -3435
rect 1675 -3455 1695 -3435
rect 425 -3505 565 -3495
rect 425 -3525 435 -3505
rect 455 -3515 565 -3505
rect 455 -3525 465 -3515
rect 425 -3535 465 -3525
rect 645 -3555 665 -3475
rect 730 -3480 770 -3470
rect 730 -3500 740 -3480
rect 760 -3500 770 -3480
rect 730 -3510 770 -3500
rect 810 -3480 860 -3470
rect 810 -3500 820 -3480
rect 840 -3500 860 -3480
rect 810 -3510 860 -3500
rect 975 -3480 1025 -3470
rect 975 -3500 985 -3480
rect 1005 -3500 1025 -3480
rect 975 -3510 1025 -3500
rect 1140 -3480 1190 -3470
rect 1140 -3500 1150 -3480
rect 1170 -3500 1190 -3480
rect 1140 -3510 1190 -3500
rect 1270 -3480 1310 -3470
rect 1270 -3500 1280 -3480
rect 1300 -3500 1310 -3480
rect 1270 -3510 1310 -3500
rect 1595 -3475 1695 -3455
rect 840 -3555 860 -3510
rect 1005 -3555 1025 -3510
rect 1170 -3555 1190 -3510
rect 1595 -3555 1615 -3475
rect 1675 -3555 1695 -3475
rect 1740 -3455 1760 -3435
rect 1740 -3465 1790 -3455
rect 1740 -3485 1760 -3465
rect 1780 -3485 1790 -3465
rect 1740 -3495 1790 -3485
rect 1740 -3555 1760 -3495
rect 1895 -3505 1915 -3435
rect 1895 -3510 1935 -3505
rect 1895 -3530 1905 -3510
rect 1925 -3530 1935 -3510
rect 1895 -3540 1935 -3530
rect 1895 -3555 1915 -3540
rect 1965 -3555 1985 -3435
rect 2030 -3495 2050 -3435
rect 2030 -3515 2195 -3495
rect 2030 -3555 2050 -3515
rect 2175 -3555 2195 -3515
rect -165 -3565 -95 -3555
rect -165 -3585 -160 -3565
rect -140 -3585 -120 -3565
rect -100 -3585 -95 -3565
rect -165 -3615 -95 -3585
rect -165 -3635 -160 -3615
rect -140 -3635 -120 -3615
rect -100 -3635 -95 -3615
rect -165 -3645 -95 -3635
rect -70 -3565 -40 -3555
rect -70 -3585 -65 -3565
rect -45 -3585 -40 -3565
rect -70 -3615 -40 -3585
rect -70 -3635 -65 -3615
rect -45 -3635 -40 -3615
rect -70 -3645 -40 -3635
rect -15 -3565 15 -3555
rect -15 -3585 -10 -3565
rect 10 -3585 15 -3565
rect -15 -3615 15 -3585
rect -15 -3635 -10 -3615
rect 10 -3635 15 -3615
rect -15 -3645 15 -3635
rect 135 -3565 165 -3555
rect 135 -3585 140 -3565
rect 160 -3585 165 -3565
rect 135 -3615 165 -3585
rect 135 -3635 140 -3615
rect 160 -3635 165 -3615
rect 135 -3645 165 -3635
rect 190 -3565 220 -3555
rect 190 -3585 195 -3565
rect 215 -3585 220 -3565
rect 190 -3615 220 -3585
rect 190 -3635 195 -3615
rect 215 -3635 220 -3615
rect 190 -3645 220 -3635
rect 245 -3565 355 -3555
rect 245 -3585 250 -3565
rect 270 -3585 290 -3565
rect 310 -3585 330 -3565
rect 350 -3585 355 -3565
rect 245 -3615 355 -3585
rect 245 -3635 250 -3615
rect 270 -3635 290 -3615
rect 310 -3635 330 -3615
rect 350 -3635 355 -3615
rect 245 -3645 355 -3635
rect 380 -3565 410 -3555
rect 380 -3585 385 -3565
rect 405 -3585 410 -3565
rect 380 -3615 410 -3585
rect 380 -3635 385 -3615
rect 405 -3635 410 -3615
rect 380 -3645 410 -3635
rect 435 -3565 465 -3555
rect 435 -3585 440 -3565
rect 460 -3585 465 -3565
rect 435 -3615 465 -3585
rect 435 -3635 440 -3615
rect 460 -3635 465 -3615
rect 435 -3645 465 -3635
rect 585 -3565 615 -3555
rect 585 -3585 590 -3565
rect 610 -3585 615 -3565
rect 585 -3615 615 -3585
rect 585 -3635 590 -3615
rect 610 -3635 615 -3615
rect 585 -3645 615 -3635
rect 640 -3565 670 -3555
rect 640 -3585 645 -3565
rect 665 -3585 670 -3565
rect 640 -3615 670 -3585
rect 640 -3635 645 -3615
rect 665 -3635 670 -3615
rect 640 -3645 670 -3635
rect 695 -3565 765 -3555
rect 695 -3585 700 -3565
rect 720 -3585 740 -3565
rect 760 -3585 765 -3565
rect 695 -3615 765 -3585
rect 695 -3635 700 -3615
rect 720 -3635 740 -3615
rect 760 -3635 765 -3615
rect 695 -3645 765 -3635
rect 840 -3565 870 -3555
rect 840 -3585 845 -3565
rect 865 -3585 870 -3565
rect 840 -3615 870 -3585
rect 840 -3635 845 -3615
rect 865 -3635 870 -3615
rect 840 -3645 870 -3635
rect 895 -3565 965 -3555
rect 895 -3585 900 -3565
rect 920 -3585 940 -3565
rect 960 -3585 965 -3565
rect 895 -3615 965 -3585
rect 895 -3635 900 -3615
rect 920 -3635 940 -3615
rect 960 -3635 965 -3615
rect 895 -3645 965 -3635
rect 1005 -3565 1035 -3555
rect 1005 -3585 1010 -3565
rect 1030 -3585 1035 -3565
rect 1005 -3615 1035 -3585
rect 1005 -3635 1010 -3615
rect 1030 -3635 1035 -3615
rect 1005 -3645 1035 -3635
rect 1060 -3565 1130 -3555
rect 1060 -3585 1065 -3565
rect 1085 -3585 1105 -3565
rect 1125 -3585 1130 -3565
rect 1060 -3615 1130 -3585
rect 1060 -3635 1065 -3615
rect 1085 -3635 1105 -3615
rect 1125 -3635 1130 -3615
rect 1060 -3645 1130 -3635
rect 1170 -3565 1200 -3555
rect 1170 -3585 1175 -3565
rect 1195 -3585 1200 -3565
rect 1170 -3615 1200 -3585
rect 1170 -3635 1175 -3615
rect 1195 -3635 1200 -3615
rect 1170 -3645 1200 -3635
rect 1225 -3565 1295 -3555
rect 1225 -3585 1230 -3565
rect 1250 -3585 1270 -3565
rect 1290 -3585 1295 -3565
rect 1225 -3615 1295 -3585
rect 1225 -3635 1230 -3615
rect 1250 -3635 1270 -3615
rect 1290 -3635 1295 -3615
rect 1225 -3645 1295 -3635
rect 1520 -3565 1560 -3555
rect 1520 -3585 1530 -3565
rect 1550 -3585 1560 -3565
rect 1520 -3615 1560 -3585
rect 1520 -3635 1530 -3615
rect 1550 -3635 1560 -3615
rect 1520 -3645 1560 -3635
rect 1585 -3565 1625 -3555
rect 1585 -3585 1595 -3565
rect 1615 -3585 1625 -3565
rect 1585 -3615 1625 -3585
rect 1585 -3635 1595 -3615
rect 1615 -3635 1625 -3615
rect 1585 -3645 1625 -3635
rect 1665 -3565 1705 -3555
rect 1665 -3585 1675 -3565
rect 1695 -3585 1705 -3565
rect 1665 -3615 1705 -3585
rect 1665 -3635 1675 -3615
rect 1695 -3635 1705 -3615
rect 1665 -3645 1705 -3635
rect 1730 -3565 1770 -3555
rect 1730 -3585 1740 -3565
rect 1760 -3585 1770 -3565
rect 1730 -3615 1770 -3585
rect 1730 -3635 1740 -3615
rect 1760 -3635 1770 -3615
rect 1730 -3645 1770 -3635
rect 1810 -3565 1850 -3555
rect 1810 -3585 1820 -3565
rect 1840 -3585 1850 -3565
rect 1810 -3615 1850 -3585
rect 1810 -3635 1820 -3615
rect 1840 -3635 1850 -3615
rect 1810 -3645 1850 -3635
rect 1875 -3565 1915 -3555
rect 1875 -3585 1885 -3565
rect 1905 -3585 1915 -3565
rect 1875 -3615 1915 -3585
rect 1875 -3635 1885 -3615
rect 1905 -3635 1915 -3615
rect 1875 -3645 1915 -3635
rect 1955 -3565 1995 -3555
rect 1955 -3585 1965 -3565
rect 1985 -3585 1995 -3565
rect 1955 -3615 1995 -3585
rect 1955 -3635 1965 -3615
rect 1985 -3635 1995 -3615
rect 1955 -3645 1995 -3635
rect 2020 -3565 2060 -3555
rect 2020 -3585 2030 -3565
rect 2050 -3585 2060 -3565
rect 2020 -3615 2060 -3585
rect 2020 -3635 2030 -3615
rect 2050 -3635 2060 -3615
rect 2020 -3645 2060 -3635
rect 2100 -3565 2140 -3555
rect 2100 -3585 2110 -3565
rect 2130 -3585 2140 -3565
rect 2100 -3615 2140 -3585
rect 2100 -3635 2110 -3615
rect 2130 -3635 2140 -3615
rect 2100 -3645 2140 -3635
rect 2165 -3565 2205 -3555
rect 2165 -3585 2175 -3565
rect 2195 -3585 2205 -3565
rect 2165 -3615 2205 -3585
rect 2165 -3635 2175 -3615
rect 2195 -3635 2205 -3615
rect 2165 -3645 2205 -3635
rect -120 -3730 -100 -3645
rect -10 -3730 10 -3645
rect 140 -3730 160 -3645
rect 255 -3730 275 -3645
rect 330 -3730 350 -3645
rect 440 -3730 460 -3645
rect 590 -3730 610 -3645
rect 700 -3730 720 -3645
rect 900 -3730 920 -3645
rect 1065 -3730 1085 -3645
rect 1230 -3730 1250 -3645
rect 1595 -3730 1615 -3645
rect 1725 -3675 1765 -3665
rect 1725 -3695 1735 -3675
rect 1755 -3695 1765 -3675
rect 1725 -3705 1765 -3695
rect 1820 -3730 1840 -3645
rect 2015 -3675 2055 -3665
rect 2015 -3695 2025 -3675
rect 2045 -3695 2055 -3675
rect 2015 -3705 2055 -3695
rect 2110 -3730 2130 -3645
rect 3185 -3720 3205 -3645
rect 3265 -3720 3285 -3645
rect 3330 -3700 4200 -3680
rect 3330 -3720 3350 -3700
rect 4055 -3720 4075 -3700
rect 2820 -3730 2860 -3720
rect -190 -3750 -170 -3730
rect -150 -3750 -120 -3730
rect -100 -3750 -70 -3730
rect -50 -3750 -20 -3730
rect 0 -3750 30 -3730
rect 50 -3750 80 -3730
rect 100 -3750 130 -3730
rect 150 -3750 180 -3730
rect 200 -3750 230 -3730
rect 250 -3750 280 -3730
rect 300 -3750 340 -3730
rect 360 -3750 390 -3730
rect 410 -3750 440 -3730
rect 460 -3750 490 -3730
rect 510 -3750 540 -3730
rect 560 -3750 590 -3730
rect 610 -3750 640 -3730
rect 660 -3750 690 -3730
rect 710 -3750 740 -3730
rect 760 -3750 790 -3730
rect 810 -3750 840 -3730
rect 860 -3750 890 -3730
rect 910 -3750 980 -3730
rect 1000 -3750 1030 -3730
rect 1050 -3750 1080 -3730
rect 1100 -3750 1170 -3730
rect 1190 -3750 1220 -3730
rect 1240 -3750 1270 -3730
rect 1290 -3750 1320 -3730
rect 1450 -3750 1470 -3730
rect 1490 -3750 1520 -3730
rect 1540 -3750 1570 -3730
rect 1590 -3750 1620 -3730
rect 1640 -3750 1670 -3730
rect 1690 -3750 1720 -3730
rect 1740 -3750 1770 -3730
rect 1790 -3750 1820 -3730
rect 1840 -3750 1870 -3730
rect 1890 -3750 1920 -3730
rect 1940 -3750 1970 -3730
rect 1990 -3750 2020 -3730
rect 2040 -3750 2070 -3730
rect 2090 -3750 2120 -3730
rect 2140 -3750 2170 -3730
rect 2190 -3750 2220 -3730
rect 2240 -3750 2270 -3730
rect 2820 -3900 2830 -3730
rect 2850 -3900 2860 -3730
rect 2820 -3910 2860 -3900
rect 2885 -3730 2925 -3720
rect 2885 -3900 2895 -3730
rect 2915 -3900 2925 -3730
rect 2885 -3910 2925 -3900
rect 2965 -3730 3005 -3720
rect 2965 -3900 2975 -3730
rect 2995 -3900 3005 -3730
rect 2965 -3910 3005 -3900
rect 3030 -3730 3070 -3720
rect 3030 -3900 3040 -3730
rect 3060 -3900 3070 -3730
rect 3030 -3910 3070 -3900
rect 3110 -3730 3150 -3720
rect 3110 -3900 3120 -3730
rect 3140 -3900 3150 -3730
rect 3110 -3910 3150 -3900
rect 3175 -3730 3215 -3720
rect 3175 -3900 3185 -3730
rect 3205 -3900 3215 -3730
rect 3175 -3910 3215 -3900
rect 3255 -3730 3295 -3720
rect 3255 -3900 3265 -3730
rect 3285 -3900 3295 -3730
rect 3255 -3910 3295 -3900
rect 3320 -3730 3360 -3720
rect 3320 -3900 3330 -3730
rect 3350 -3900 3360 -3730
rect 3320 -3910 3360 -3900
rect 3400 -3730 3440 -3720
rect 3400 -3900 3410 -3730
rect 3430 -3900 3440 -3730
rect 3400 -3910 3440 -3900
rect 3465 -3730 3505 -3720
rect 3465 -3900 3475 -3730
rect 3495 -3880 3505 -3730
rect 3545 -3730 3585 -3720
rect 3495 -3900 3510 -3880
rect 3465 -3910 3510 -3900
rect 3545 -3900 3555 -3730
rect 3575 -3900 3585 -3730
rect 3545 -3910 3585 -3900
rect 3610 -3730 3650 -3720
rect 3610 -3900 3620 -3730
rect 3640 -3900 3650 -3730
rect 3610 -3910 3650 -3900
rect 3690 -3730 3730 -3720
rect 3690 -3900 3700 -3730
rect 3720 -3900 3730 -3730
rect 3690 -3910 3730 -3900
rect 3755 -3730 3795 -3720
rect 3755 -3900 3765 -3730
rect 3785 -3900 3795 -3730
rect 3755 -3910 3795 -3900
rect 3835 -3730 3875 -3720
rect 3835 -3900 3845 -3730
rect 3865 -3900 3875 -3730
rect 3835 -3910 3875 -3900
rect 3900 -3730 3940 -3720
rect 3900 -3900 3910 -3730
rect 3930 -3900 3940 -3730
rect 3900 -3910 3940 -3900
rect 3980 -3730 4020 -3720
rect 3980 -3900 3990 -3730
rect 4010 -3900 4020 -3730
rect 3980 -3910 4020 -3900
rect 4045 -3730 4085 -3720
rect 4045 -3900 4055 -3730
rect 4075 -3900 4085 -3730
rect 4045 -3910 4085 -3900
rect 4125 -3730 4165 -3720
rect 4125 -3900 4135 -3730
rect 4155 -3900 4165 -3730
rect 4125 -3910 4165 -3900
rect 2905 -3965 2925 -3910
rect 2985 -3965 3025 -3955
rect 2905 -3985 2995 -3965
rect 3015 -3985 3025 -3965
rect 2905 -4050 2925 -3985
rect 2985 -3995 3025 -3985
rect 3050 -3965 3070 -3910
rect 3195 -3930 3215 -3910
rect 3195 -3940 3235 -3930
rect 3130 -3965 3170 -3955
rect 3050 -3985 3140 -3965
rect 3160 -3985 3170 -3965
rect 3050 -4050 3070 -3985
rect 3130 -3995 3170 -3985
rect 3195 -3960 3205 -3940
rect 3225 -3960 3235 -3940
rect 3195 -3970 3235 -3960
rect 3195 -4050 3215 -3970
rect 3265 -4050 3285 -3910
rect 3320 -4050 3340 -3910
rect 3420 -3930 3440 -3910
rect 3555 -3930 3575 -3910
rect 3420 -3950 3575 -3930
rect 3420 -4050 3440 -3950
rect 3485 -4000 3525 -3990
rect 3485 -4020 3495 -4000
rect 3515 -4020 3525 -4000
rect 3485 -4030 3525 -4020
rect 3485 -4050 3505 -4030
rect 3555 -4050 3575 -3950
rect 3620 -3930 3640 -3910
rect 3620 -3940 3670 -3930
rect 3620 -3960 3640 -3940
rect 3660 -3960 3670 -3940
rect 3620 -3965 3670 -3960
rect 3620 -4050 3640 -3965
rect 3695 -3990 3715 -3910
rect 3670 -4000 3715 -3990
rect 3670 -4020 3680 -4000
rect 3700 -4020 3715 -4000
rect 3670 -4030 3715 -4020
rect 3775 -3995 3795 -3910
rect 3775 -4005 3815 -3995
rect 3775 -4025 3785 -4005
rect 3805 -4025 3815 -4005
rect 3775 -4035 3815 -4025
rect 3775 -4050 3795 -4035
rect 3845 -4050 3865 -3910
rect 3910 -3990 3930 -3910
rect 3910 -4010 4200 -3990
rect 3910 -4050 3930 -4010
rect 4055 -4050 4075 -4010
rect 2820 -4060 2860 -4050
rect 2820 -4130 2830 -4060
rect 2850 -4130 2860 -4060
rect 2820 -4140 2860 -4130
rect 2885 -4060 2925 -4050
rect 2885 -4130 2895 -4060
rect 2915 -4130 2925 -4060
rect 2885 -4140 2925 -4130
rect 2965 -4060 3005 -4050
rect 2965 -4130 2975 -4060
rect 2995 -4130 3005 -4060
rect 2965 -4140 3005 -4130
rect 3030 -4060 3070 -4050
rect 3030 -4130 3040 -4060
rect 3060 -4130 3070 -4060
rect 3030 -4140 3070 -4130
rect 3110 -4060 3150 -4050
rect 3110 -4130 3120 -4060
rect 3140 -4130 3150 -4060
rect 3110 -4140 3150 -4130
rect 3175 -4060 3215 -4050
rect 3175 -4130 3185 -4060
rect 3205 -4130 3215 -4060
rect 3175 -4140 3215 -4130
rect 3255 -4060 3295 -4050
rect 3255 -4130 3265 -4060
rect 3285 -4130 3295 -4060
rect 3255 -4140 3295 -4130
rect 3320 -4060 3360 -4050
rect 3320 -4130 3330 -4060
rect 3350 -4130 3360 -4060
rect 3320 -4140 3360 -4130
rect 3400 -4060 3440 -4050
rect 3400 -4130 3410 -4060
rect 3430 -4130 3440 -4060
rect 3400 -4140 3440 -4130
rect 3465 -4060 3505 -4050
rect 3465 -4130 3475 -4060
rect 3495 -4130 3505 -4060
rect 3465 -4140 3505 -4130
rect 3545 -4060 3585 -4050
rect 3545 -4130 3555 -4060
rect 3575 -4130 3585 -4060
rect 3545 -4140 3585 -4130
rect 3610 -4060 3650 -4050
rect 3610 -4130 3620 -4060
rect 3640 -4130 3650 -4060
rect 3610 -4140 3650 -4130
rect 3690 -4060 3730 -4050
rect 3690 -4130 3700 -4060
rect 3720 -4130 3730 -4060
rect 3690 -4140 3730 -4130
rect 3755 -4060 3795 -4050
rect 3755 -4130 3765 -4060
rect 3785 -4130 3795 -4060
rect 3755 -4140 3795 -4130
rect 3835 -4060 3875 -4050
rect 3835 -4130 3845 -4060
rect 3865 -4130 3875 -4060
rect 3835 -4140 3875 -4130
rect 3900 -4060 3945 -4050
rect 3900 -4130 3910 -4060
rect 3930 -4130 3945 -4060
rect 3900 -4140 3945 -4130
rect 3980 -4060 4020 -4050
rect 3980 -4130 3990 -4060
rect 4010 -4130 4020 -4060
rect 3980 -4140 4020 -4130
rect 4045 -4060 4085 -4050
rect 4045 -4130 4055 -4060
rect 4075 -4130 4085 -4060
rect 4045 -4140 4085 -4130
rect 4125 -4060 4165 -4050
rect 4125 -4130 4135 -4060
rect 4155 -4130 4165 -4060
rect 4125 -4140 4165 -4130
rect 2775 -4175 3355 -4160
rect 3845 -4175 3865 -4140
rect 3895 -4170 3935 -4160
rect 3895 -4175 3905 -4170
rect 3925 -4175 3935 -4170
rect 1450 -4930 1470 -4910
rect 1490 -4930 1520 -4910
rect 1540 -4930 1570 -4910
rect 1590 -4930 1620 -4910
rect 1640 -4930 1670 -4910
rect 1690 -4930 1720 -4910
rect 1740 -4930 1770 -4910
rect 1790 -4930 1820 -4910
rect 1840 -4930 1870 -4910
rect 1890 -4930 1920 -4910
rect 1940 -4930 1970 -4910
rect 1990 -4930 2020 -4910
rect 2040 -4930 2070 -4910
rect 2090 -4930 2120 -4910
rect 2140 -4930 2170 -4910
rect 2190 -4930 2220 -4910
rect 2240 -4930 2270 -4910
rect 1530 -5105 1550 -4930
rect 1675 -5105 1695 -4930
rect 1820 -5105 1840 -4930
rect 1520 -5115 1560 -5105
rect 1520 -5135 1530 -5115
rect 1550 -5135 1560 -5115
rect 1520 -5165 1560 -5135
rect 1520 -5185 1530 -5165
rect 1550 -5185 1560 -5165
rect 1520 -5195 1560 -5185
rect 1585 -5115 1625 -5105
rect 1585 -5135 1595 -5115
rect 1615 -5135 1625 -5115
rect 1585 -5165 1625 -5135
rect 1585 -5185 1595 -5165
rect 1615 -5185 1625 -5165
rect 1585 -5195 1625 -5185
rect 1665 -5115 1705 -5105
rect 1665 -5135 1675 -5115
rect 1695 -5135 1705 -5115
rect 1665 -5165 1705 -5135
rect 1665 -5185 1675 -5165
rect 1695 -5185 1705 -5165
rect 1665 -5195 1705 -5185
rect 1730 -5115 1770 -5105
rect 1730 -5135 1740 -5115
rect 1760 -5135 1770 -5115
rect 1730 -5165 1770 -5135
rect 1730 -5185 1740 -5165
rect 1760 -5185 1770 -5165
rect 1730 -5195 1770 -5185
rect 1810 -5115 1850 -5105
rect 1810 -5135 1820 -5115
rect 1840 -5135 1850 -5115
rect 1810 -5165 1850 -5135
rect 1810 -5185 1820 -5165
rect 1840 -5185 1850 -5165
rect 1810 -5195 1850 -5185
rect 1875 -5115 1915 -5105
rect 1875 -5135 1885 -5115
rect 1905 -5135 1915 -5115
rect 1875 -5165 1915 -5135
rect 1875 -5185 1885 -5165
rect 1905 -5185 1915 -5165
rect 1875 -5195 1915 -5185
rect 1955 -5115 1995 -5105
rect 1955 -5135 1965 -5115
rect 1985 -5135 1995 -5115
rect 1955 -5165 1995 -5135
rect 1955 -5185 1965 -5165
rect 1985 -5185 1995 -5165
rect 1955 -5195 1995 -5185
rect 2020 -5115 2060 -5105
rect 2020 -5135 2030 -5115
rect 2050 -5135 2060 -5115
rect 2020 -5165 2060 -5135
rect 2020 -5185 2030 -5165
rect 2050 -5185 2060 -5165
rect 2020 -5195 2060 -5185
rect 1605 -5260 1625 -5195
rect 1685 -5260 1725 -5250
rect 1605 -5280 1695 -5260
rect 1715 -5280 1725 -5260
rect 1605 -5335 1625 -5280
rect 1685 -5290 1725 -5280
rect 1750 -5260 1770 -5195
rect 1830 -5260 1870 -5250
rect 1750 -5280 1840 -5260
rect 1860 -5280 1870 -5260
rect 1750 -5335 1770 -5280
rect 1830 -5290 1870 -5280
rect 1895 -5275 1915 -5195
rect 1895 -5285 1935 -5275
rect 1895 -5305 1905 -5285
rect 1925 -5305 1935 -5285
rect 1895 -5315 1935 -5305
rect 1895 -5335 1915 -5315
rect 1965 -5335 1985 -5195
rect 2020 -5335 2040 -5195
rect 1520 -5345 1560 -5335
rect 1520 -5365 1530 -5345
rect 1550 -5365 1560 -5345
rect 1520 -5395 1560 -5365
rect 1520 -5415 1530 -5395
rect 1550 -5415 1560 -5395
rect 1520 -5445 1560 -5415
rect 1520 -5465 1530 -5445
rect 1550 -5465 1560 -5445
rect 1520 -5495 1560 -5465
rect 1520 -5515 1530 -5495
rect 1550 -5515 1560 -5495
rect 1520 -5525 1560 -5515
rect 1585 -5345 1625 -5335
rect 1585 -5365 1595 -5345
rect 1615 -5365 1625 -5345
rect 1585 -5395 1625 -5365
rect 1585 -5415 1595 -5395
rect 1615 -5415 1625 -5395
rect 1585 -5445 1625 -5415
rect 1585 -5465 1595 -5445
rect 1615 -5465 1625 -5445
rect 1585 -5495 1625 -5465
rect 1585 -5515 1595 -5495
rect 1615 -5515 1625 -5495
rect 1585 -5525 1625 -5515
rect 1665 -5345 1705 -5335
rect 1665 -5365 1675 -5345
rect 1695 -5365 1705 -5345
rect 1665 -5395 1705 -5365
rect 1665 -5415 1675 -5395
rect 1695 -5415 1705 -5395
rect 1665 -5445 1705 -5415
rect 1665 -5465 1675 -5445
rect 1695 -5465 1705 -5445
rect 1665 -5495 1705 -5465
rect 1665 -5515 1675 -5495
rect 1695 -5515 1705 -5495
rect 1665 -5525 1705 -5515
rect 1730 -5345 1770 -5335
rect 1730 -5365 1740 -5345
rect 1760 -5365 1770 -5345
rect 1730 -5395 1770 -5365
rect 1730 -5415 1740 -5395
rect 1760 -5415 1770 -5395
rect 1730 -5445 1770 -5415
rect 1730 -5465 1740 -5445
rect 1760 -5465 1770 -5445
rect 1730 -5495 1770 -5465
rect 1730 -5515 1740 -5495
rect 1760 -5515 1770 -5495
rect 1730 -5525 1770 -5515
rect 1810 -5345 1850 -5335
rect 1810 -5365 1820 -5345
rect 1840 -5365 1850 -5345
rect 1810 -5395 1850 -5365
rect 1810 -5415 1820 -5395
rect 1840 -5415 1850 -5395
rect 1810 -5445 1850 -5415
rect 1810 -5465 1820 -5445
rect 1840 -5465 1850 -5445
rect 1810 -5495 1850 -5465
rect 1810 -5515 1820 -5495
rect 1840 -5515 1850 -5495
rect 1810 -5525 1850 -5515
rect 1875 -5345 1915 -5335
rect 1875 -5365 1885 -5345
rect 1905 -5365 1915 -5345
rect 1875 -5395 1915 -5365
rect 1875 -5415 1885 -5395
rect 1905 -5415 1915 -5395
rect 1875 -5445 1915 -5415
rect 1875 -5465 1885 -5445
rect 1905 -5465 1915 -5445
rect 1875 -5495 1915 -5465
rect 1875 -5515 1885 -5495
rect 1905 -5515 1915 -5495
rect 1875 -5525 1915 -5515
rect 1955 -5345 1995 -5335
rect 1955 -5365 1965 -5345
rect 1985 -5365 1995 -5345
rect 1955 -5395 1995 -5365
rect 1955 -5415 1965 -5395
rect 1985 -5415 1995 -5395
rect 1955 -5445 1995 -5415
rect 1955 -5465 1965 -5445
rect 1985 -5465 1995 -5445
rect 1955 -5495 1995 -5465
rect 1955 -5515 1965 -5495
rect 1985 -5515 1995 -5495
rect 1955 -5525 1995 -5515
rect 2020 -5345 2060 -5335
rect 2020 -5365 2030 -5345
rect 2050 -5365 2060 -5345
rect 2020 -5395 2060 -5365
rect 2020 -5415 2030 -5395
rect 2050 -5415 2060 -5395
rect 2020 -5445 2060 -5415
rect 2020 -5465 2030 -5445
rect 2050 -5465 2060 -5445
rect 2020 -5495 2060 -5465
rect 2020 -5515 2030 -5495
rect 2050 -5515 2060 -5495
rect 2020 -5525 2060 -5515
rect 1530 -5610 1550 -5525
rect 1675 -5610 1695 -5525
rect 1820 -5610 1840 -5525
rect 1450 -5630 1470 -5610
rect 1490 -5630 1520 -5610
rect 1540 -5630 1570 -5610
rect 1590 -5630 1620 -5610
rect 1640 -5630 1670 -5610
rect 1690 -5630 1720 -5610
rect 1740 -5630 1770 -5610
rect 1790 -5630 1820 -5610
rect 1840 -5630 1870 -5610
rect 1890 -5630 1920 -5610
rect 1940 -5630 1970 -5610
rect 1990 -5630 2020 -5610
rect 2040 -5630 2070 -5610
rect 2090 -5630 2120 -5610
rect 2140 -5630 2170 -5610
rect 2190 -5630 2220 -5610
rect 2240 -5630 2270 -5610
rect 1595 -5725 1615 -5630
rect 1820 -5725 1840 -5630
rect 1520 -5735 1560 -5725
rect 1520 -5755 1530 -5735
rect 1550 -5755 1560 -5735
rect 1520 -5785 1560 -5755
rect 1520 -5805 1530 -5785
rect 1550 -5805 1560 -5785
rect 1520 -5835 1560 -5805
rect 1520 -5855 1530 -5835
rect 1550 -5855 1560 -5835
rect 1520 -5885 1560 -5855
rect 1520 -5905 1530 -5885
rect 1550 -5905 1560 -5885
rect 1520 -5915 1560 -5905
rect 1585 -5735 1625 -5725
rect 1585 -5755 1595 -5735
rect 1615 -5755 1625 -5735
rect 1585 -5785 1625 -5755
rect 1585 -5805 1595 -5785
rect 1615 -5805 1625 -5785
rect 1585 -5835 1625 -5805
rect 1585 -5855 1595 -5835
rect 1615 -5855 1625 -5835
rect 1585 -5885 1625 -5855
rect 1585 -5905 1595 -5885
rect 1615 -5905 1625 -5885
rect 1585 -5915 1625 -5905
rect 1665 -5735 1705 -5725
rect 1665 -5755 1675 -5735
rect 1695 -5755 1705 -5735
rect 1665 -5785 1705 -5755
rect 1665 -5805 1675 -5785
rect 1695 -5805 1705 -5785
rect 1665 -5835 1705 -5805
rect 1665 -5855 1675 -5835
rect 1695 -5855 1705 -5835
rect 1665 -5885 1705 -5855
rect 1665 -5905 1675 -5885
rect 1695 -5905 1705 -5885
rect 1665 -5915 1705 -5905
rect 1730 -5735 1770 -5725
rect 1730 -5755 1740 -5735
rect 1760 -5755 1770 -5735
rect 1730 -5785 1770 -5755
rect 1730 -5805 1740 -5785
rect 1760 -5805 1770 -5785
rect 1730 -5835 1770 -5805
rect 1730 -5855 1740 -5835
rect 1760 -5855 1770 -5835
rect 1730 -5885 1770 -5855
rect 1730 -5905 1740 -5885
rect 1760 -5905 1770 -5885
rect 1730 -5915 1770 -5905
rect 1810 -5735 1850 -5725
rect 1810 -5755 1820 -5735
rect 1840 -5755 1850 -5735
rect 1810 -5785 1850 -5755
rect 1810 -5805 1820 -5785
rect 1840 -5805 1850 -5785
rect 1810 -5835 1850 -5805
rect 1810 -5855 1820 -5835
rect 1840 -5855 1850 -5835
rect 1810 -5885 1850 -5855
rect 1810 -5905 1820 -5885
rect 1840 -5905 1850 -5885
rect 1810 -5915 1850 -5905
rect 1875 -5735 1915 -5725
rect 1875 -5755 1885 -5735
rect 1905 -5755 1915 -5735
rect 1875 -5785 1915 -5755
rect 1875 -5805 1885 -5785
rect 1905 -5805 1915 -5785
rect 1875 -5835 1915 -5805
rect 1875 -5855 1885 -5835
rect 1905 -5855 1915 -5835
rect 1875 -5885 1915 -5855
rect 1875 -5905 1885 -5885
rect 1905 -5905 1915 -5885
rect 1875 -5915 1915 -5905
rect 1955 -5735 1995 -5725
rect 1955 -5755 1965 -5735
rect 1985 -5755 1995 -5735
rect 1955 -5785 1995 -5755
rect 1955 -5805 1965 -5785
rect 1985 -5805 1995 -5785
rect 1955 -5835 1995 -5805
rect 1955 -5855 1965 -5835
rect 1985 -5855 1995 -5835
rect 1955 -5885 1995 -5855
rect 1955 -5905 1965 -5885
rect 1985 -5905 1995 -5885
rect 1955 -5915 1995 -5905
rect 2020 -5735 2060 -5725
rect 2020 -5755 2030 -5735
rect 2050 -5755 2060 -5735
rect 2020 -5785 2060 -5755
rect 2020 -5805 2030 -5785
rect 2050 -5805 2060 -5785
rect 2020 -5835 2060 -5805
rect 2020 -5855 2030 -5835
rect 2050 -5855 2060 -5835
rect 2020 -5885 2060 -5855
rect 2020 -5905 2030 -5885
rect 2050 -5905 2060 -5885
rect 2020 -5915 2060 -5905
rect 2100 -5735 2140 -5725
rect 2100 -5755 2110 -5735
rect 2130 -5755 2140 -5735
rect 2100 -5785 2140 -5755
rect 2100 -5805 2110 -5785
rect 2130 -5805 2140 -5785
rect 2100 -5835 2140 -5805
rect 2100 -5855 2110 -5835
rect 2130 -5855 2140 -5835
rect 2100 -5885 2140 -5855
rect 2100 -5905 2110 -5885
rect 2130 -5905 2140 -5885
rect 2100 -5915 2140 -5905
rect 2165 -5735 2205 -5725
rect 2165 -5755 2175 -5735
rect 2195 -5755 2205 -5735
rect 2165 -5785 2205 -5755
rect 2165 -5805 2175 -5785
rect 2195 -5805 2205 -5785
rect 2165 -5835 2205 -5805
rect 2165 -5855 2175 -5835
rect 2195 -5855 2205 -5835
rect 2165 -5885 2205 -5855
rect 2165 -5905 2175 -5885
rect 2195 -5905 2205 -5885
rect 2165 -5915 2205 -5905
rect 1540 -5935 1560 -5915
rect 1675 -5935 1695 -5915
rect 1540 -5955 1695 -5935
rect 1540 -6055 1560 -5955
rect 1605 -6005 1645 -5995
rect 1605 -6025 1615 -6005
rect 1635 -6025 1645 -6005
rect 1605 -6035 1645 -6025
rect 1605 -6055 1625 -6035
rect 1675 -6055 1695 -5955
rect 1740 -5935 1760 -5915
rect 1740 -5945 1790 -5935
rect 1740 -5965 1760 -5945
rect 1780 -5965 1790 -5945
rect 1740 -5970 1790 -5965
rect 1740 -6055 1760 -5970
rect 1815 -5995 1835 -5915
rect 1790 -6005 1835 -5995
rect 1790 -6025 1800 -6005
rect 1820 -6025 1835 -6005
rect 1790 -6035 1835 -6025
rect 1895 -6000 1915 -5915
rect 1895 -6010 1935 -6000
rect 1895 -6030 1905 -6010
rect 1925 -6030 1935 -6010
rect 1895 -6040 1935 -6030
rect 1895 -6055 1915 -6040
rect 1965 -6055 1985 -5915
rect 2030 -5995 2050 -5915
rect 2030 -6015 2225 -5995
rect 2030 -6055 2050 -6015
rect 2175 -6055 2195 -6015
rect 1520 -6065 1560 -6055
rect 1520 -6085 1530 -6065
rect 1550 -6085 1560 -6065
rect 1520 -6115 1560 -6085
rect 1520 -6135 1530 -6115
rect 1550 -6135 1560 -6115
rect 1520 -6145 1560 -6135
rect 1585 -6065 1625 -6055
rect 1585 -6085 1595 -6065
rect 1615 -6085 1625 -6065
rect 1585 -6115 1625 -6085
rect 1585 -6135 1595 -6115
rect 1615 -6135 1625 -6115
rect 1585 -6145 1625 -6135
rect 1665 -6065 1705 -6055
rect 1665 -6085 1675 -6065
rect 1695 -6085 1705 -6065
rect 1665 -6115 1705 -6085
rect 1665 -6135 1675 -6115
rect 1695 -6135 1705 -6115
rect 1665 -6145 1705 -6135
rect 1730 -6065 1770 -6055
rect 1730 -6085 1740 -6065
rect 1760 -6085 1770 -6065
rect 1730 -6115 1770 -6085
rect 1730 -6135 1740 -6115
rect 1760 -6135 1770 -6115
rect 1730 -6145 1770 -6135
rect 1810 -6065 1850 -6055
rect 1810 -6085 1820 -6065
rect 1840 -6085 1850 -6065
rect 1810 -6115 1850 -6085
rect 1810 -6135 1820 -6115
rect 1840 -6135 1850 -6115
rect 1810 -6145 1850 -6135
rect 1875 -6065 1915 -6055
rect 1875 -6085 1885 -6065
rect 1905 -6085 1915 -6065
rect 1875 -6115 1915 -6085
rect 1875 -6135 1885 -6115
rect 1905 -6135 1915 -6115
rect 1875 -6145 1915 -6135
rect 1955 -6065 1995 -6055
rect 1955 -6085 1965 -6065
rect 1985 -6085 1995 -6065
rect 1955 -6115 1995 -6085
rect 1955 -6135 1965 -6115
rect 1985 -6135 1995 -6115
rect 1955 -6145 1995 -6135
rect 2020 -6065 2065 -6055
rect 2020 -6085 2030 -6065
rect 2050 -6085 2065 -6065
rect 2020 -6115 2065 -6085
rect 2020 -6135 2030 -6115
rect 2050 -6135 2065 -6115
rect 2020 -6145 2065 -6135
rect 2100 -6065 2140 -6055
rect 2100 -6085 2110 -6065
rect 2130 -6085 2140 -6065
rect 2100 -6115 2140 -6085
rect 2100 -6135 2110 -6115
rect 2130 -6135 2140 -6115
rect 2100 -6145 2140 -6135
rect 2165 -6065 2205 -6055
rect 2165 -6085 2175 -6065
rect 2195 -6085 2205 -6065
rect 2165 -6115 2205 -6085
rect 2165 -6135 2175 -6115
rect 2195 -6135 2205 -6115
rect 2165 -6145 2205 -6135
rect 1595 -6215 1615 -6145
rect 1820 -6215 1840 -6145
rect 2110 -6215 2130 -6145
rect 1450 -6235 1470 -6215
rect 1490 -6235 1520 -6215
rect 1540 -6235 1570 -6215
rect 1590 -6235 1620 -6215
rect 1640 -6235 1670 -6215
rect 1690 -6235 1720 -6215
rect 1740 -6235 1770 -6215
rect 1790 -6235 1820 -6215
rect 1840 -6235 1870 -6215
rect 1890 -6235 1920 -6215
rect 1940 -6235 1970 -6215
rect 1990 -6235 2020 -6215
rect 2040 -6235 2070 -6215
rect 2090 -6235 2120 -6215
rect 2140 -6235 2170 -6215
rect 2190 -6235 2220 -6215
rect 2240 -6235 2270 -6215
<< viali >>
rect -30 175 -10 245
rect 340 175 360 245
rect 410 175 430 245
rect 780 175 800 245
rect 850 175 870 245
rect 1220 175 1240 245
rect 1260 175 1280 245
rect 1300 175 1320 245
rect 1670 175 1690 245
rect 1795 175 1815 245
rect 1920 175 1940 245
rect 2045 175 2065 245
rect 2170 175 2190 245
rect 2295 175 2315 245
rect 2420 175 2440 245
rect -30 15 -10 35
rect 80 15 100 35
rect 230 15 250 35
rect 340 15 360 35
rect 410 15 430 35
rect 520 15 540 35
rect 670 15 690 35
rect 780 15 800 35
rect 850 15 870 35
rect 960 15 980 35
rect 1110 15 1130 35
rect 1220 15 1240 35
rect 1260 15 1280 35
rect 1300 15 1320 35
rect 1410 15 1430 35
rect 1560 15 1580 35
rect 1670 15 1690 35
rect 1740 15 1760 35
rect 1920 15 1940 35
rect 2045 15 2065 35
rect 2170 15 2190 35
rect 2295 15 2315 35
rect 2420 15 2440 35
rect -30 -1235 -10 -1215
rect 80 -1235 100 -1215
rect 230 -1235 250 -1215
rect 340 -1235 360 -1215
rect 410 -1235 430 -1215
rect 520 -1235 540 -1215
rect 670 -1235 690 -1215
rect 780 -1235 800 -1215
rect 910 -1235 930 -1215
rect 1090 -1235 1110 -1215
rect 1215 -1235 1235 -1215
rect -30 -1445 -10 -1375
rect 340 -1445 360 -1375
rect 410 -1445 430 -1375
rect 780 -1445 800 -1375
rect 965 -1445 985 -1375
rect 1090 -1445 1110 -1375
rect 1215 -1445 1235 -1375
rect -30 -1825 -10 -1755
rect 340 -1825 360 -1755
rect 410 -1825 430 -1755
rect 780 -1825 800 -1755
rect 1015 -1825 1035 -1755
rect 1140 -1825 1160 -1755
rect 1265 -1825 1285 -1755
rect -30 -1985 -10 -1965
rect 80 -1985 100 -1965
rect 230 -1985 250 -1965
rect 340 -1985 360 -1965
rect 410 -1985 430 -1965
rect 520 -1985 540 -1965
rect 670 -1985 690 -1965
rect 780 -1985 800 -1965
rect 1015 -1985 1035 -1965
rect 1140 -1985 1160 -1965
rect 1265 -1985 1285 -1965
rect -170 -2570 -150 -2550
rect -120 -2570 -100 -2550
rect -70 -2570 -50 -2550
rect -20 -2570 0 -2550
rect 30 -2570 50 -2550
rect 80 -2570 100 -2550
rect 130 -2570 150 -2550
rect 180 -2570 200 -2550
rect 230 -2570 250 -2550
rect 280 -2570 300 -2550
rect 340 -2570 360 -2550
rect 390 -2570 410 -2550
rect 440 -2570 460 -2550
rect 490 -2570 510 -2550
rect 540 -2570 560 -2550
rect 590 -2570 610 -2550
rect 640 -2570 660 -2550
rect 690 -2570 710 -2550
rect 740 -2570 760 -2550
rect 790 -2570 810 -2550
rect 840 -2570 860 -2550
rect 890 -2570 910 -2550
rect 980 -2570 1000 -2550
rect 1030 -2570 1050 -2550
rect 1080 -2570 1100 -2550
rect 1170 -2570 1190 -2550
rect 1220 -2570 1240 -2550
rect 1270 -2570 1290 -2550
rect 1470 -2570 1490 -2550
rect 1520 -2570 1540 -2550
rect 1570 -2570 1590 -2550
rect 1620 -2570 1640 -2550
rect 1670 -2570 1690 -2550
rect 1720 -2570 1740 -2550
rect 1770 -2570 1790 -2550
rect 1820 -2570 1840 -2550
rect 1870 -2570 1890 -2550
rect 1920 -2570 1940 -2550
rect 1970 -2570 1990 -2550
rect 2020 -2570 2040 -2550
rect 2070 -2570 2090 -2550
rect 2120 -2570 2140 -2550
rect 2170 -2570 2190 -2550
rect 2220 -2570 2240 -2550
rect 85 -2625 105 -2605
rect 890 -2625 910 -2605
rect 730 -2800 750 -2780
rect 1260 -2820 1280 -2800
rect 805 -3105 825 -3085
rect -170 -3160 -150 -3140
rect -120 -3160 -100 -3140
rect -70 -3160 -50 -3140
rect -20 -3160 0 -3140
rect 30 -3160 50 -3140
rect 80 -3160 100 -3140
rect 130 -3160 150 -3140
rect 180 -3160 200 -3140
rect 230 -3160 250 -3140
rect 280 -3160 300 -3140
rect 340 -3160 360 -3140
rect 390 -3160 410 -3140
rect 440 -3160 460 -3140
rect 490 -3160 510 -3140
rect 540 -3160 560 -3140
rect 590 -3160 610 -3140
rect 640 -3160 660 -3140
rect 690 -3160 710 -3140
rect 740 -3160 760 -3140
rect 790 -3160 810 -3140
rect 840 -3160 860 -3140
rect 890 -3160 910 -3140
rect 980 -3160 1000 -3140
rect 1030 -3160 1050 -3140
rect 1080 -3160 1100 -3140
rect 1170 -3160 1190 -3140
rect 1220 -3160 1240 -3140
rect 1270 -3160 1290 -3140
rect 1470 -3160 1490 -3140
rect 1520 -3160 1540 -3140
rect 1570 -3160 1590 -3140
rect 1620 -3160 1640 -3140
rect 1670 -3160 1690 -3140
rect 1720 -3160 1740 -3140
rect 1770 -3160 1790 -3140
rect 1820 -3160 1840 -3140
rect 1870 -3160 1890 -3140
rect 1920 -3160 1940 -3140
rect 1970 -3160 1990 -3140
rect 2020 -3160 2040 -3140
rect 2070 -3160 2090 -3140
rect 2120 -3160 2140 -3140
rect 2170 -3160 2190 -3140
rect 2220 -3160 2240 -3140
rect 105 -3215 125 -3195
rect 1695 -3215 1715 -3195
rect 1985 -3215 2005 -3195
rect 740 -3500 760 -3480
rect 1280 -3500 1300 -3480
rect 1735 -3695 1755 -3675
rect 2025 -3695 2045 -3675
rect -170 -3750 -150 -3730
rect -120 -3750 -100 -3730
rect -70 -3750 -50 -3730
rect -20 -3750 0 -3730
rect 30 -3750 50 -3730
rect 80 -3750 100 -3730
rect 130 -3750 150 -3730
rect 180 -3750 200 -3730
rect 230 -3750 250 -3730
rect 280 -3750 300 -3730
rect 340 -3750 360 -3730
rect 390 -3750 410 -3730
rect 440 -3750 460 -3730
rect 490 -3750 510 -3730
rect 540 -3750 560 -3730
rect 590 -3750 610 -3730
rect 640 -3750 660 -3730
rect 690 -3750 710 -3730
rect 740 -3750 760 -3730
rect 790 -3750 810 -3730
rect 840 -3750 860 -3730
rect 890 -3750 910 -3730
rect 980 -3750 1000 -3730
rect 1030 -3750 1050 -3730
rect 1080 -3750 1100 -3730
rect 1170 -3750 1190 -3730
rect 1220 -3750 1240 -3730
rect 1270 -3750 1290 -3730
rect 1470 -3750 1490 -3730
rect 1520 -3750 1540 -3730
rect 1570 -3750 1590 -3730
rect 1620 -3750 1640 -3730
rect 1670 -3750 1690 -3730
rect 1720 -3750 1740 -3730
rect 1770 -3750 1790 -3730
rect 1820 -3750 1840 -3730
rect 1870 -3750 1890 -3730
rect 1920 -3750 1940 -3730
rect 1970 -3750 1990 -3730
rect 2020 -3750 2040 -3730
rect 2070 -3750 2090 -3730
rect 2120 -3750 2140 -3730
rect 2170 -3750 2190 -3730
rect 2220 -3750 2240 -3730
rect 1470 -4930 1490 -4910
rect 1520 -4930 1540 -4910
rect 1570 -4930 1590 -4910
rect 1620 -4930 1640 -4910
rect 1670 -4930 1690 -4910
rect 1720 -4930 1740 -4910
rect 1770 -4930 1790 -4910
rect 1820 -4930 1840 -4910
rect 1870 -4930 1890 -4910
rect 1920 -4930 1940 -4910
rect 1970 -4930 1990 -4910
rect 2020 -4930 2040 -4910
rect 2070 -4930 2090 -4910
rect 2120 -4930 2140 -4910
rect 2170 -4930 2190 -4910
rect 2220 -4930 2240 -4910
rect 1470 -5630 1490 -5610
rect 1520 -5630 1540 -5610
rect 1570 -5630 1590 -5610
rect 1620 -5630 1640 -5610
rect 1670 -5630 1690 -5610
rect 1720 -5630 1740 -5610
rect 1770 -5630 1790 -5610
rect 1820 -5630 1840 -5610
rect 1870 -5630 1890 -5610
rect 1920 -5630 1940 -5610
rect 1970 -5630 1990 -5610
rect 2020 -5630 2040 -5610
rect 2070 -5630 2090 -5610
rect 2120 -5630 2140 -5610
rect 2170 -5630 2190 -5610
rect 2220 -5630 2240 -5610
rect 1470 -6235 1490 -6215
rect 1520 -6235 1540 -6215
rect 1570 -6235 1590 -6215
rect 1620 -6235 1640 -6215
rect 1670 -6235 1690 -6215
rect 1720 -6235 1740 -6215
rect 1770 -6235 1790 -6215
rect 1820 -6235 1840 -6215
rect 1870 -6235 1890 -6215
rect 1920 -6235 1940 -6215
rect 1970 -6235 1990 -6215
rect 2020 -6235 2040 -6215
rect 2070 -6235 2090 -6215
rect 2120 -6235 2140 -6215
rect 2170 -6235 2190 -6215
rect 2220 -6235 2240 -6215
<< metal1 >>
rect -40 245 2505 260
rect -40 175 -30 245
rect -10 175 340 245
rect 360 175 410 245
rect 430 175 780 245
rect 800 175 850 245
rect 870 175 1220 245
rect 1240 175 1260 245
rect 1280 175 1300 245
rect 1320 175 1670 245
rect 1690 175 1795 245
rect 1815 175 1920 245
rect 1940 175 2045 245
rect 2065 175 2170 245
rect 2190 175 2295 245
rect 2315 175 2420 245
rect 2440 175 2505 245
rect -40 160 2505 175
rect -40 35 2505 50
rect -40 15 -30 35
rect -10 15 80 35
rect 100 15 230 35
rect 250 15 340 35
rect 360 15 410 35
rect 430 15 520 35
rect 540 15 670 35
rect 690 15 780 35
rect 800 15 850 35
rect 870 15 960 35
rect 980 15 1110 35
rect 1130 15 1220 35
rect 1240 15 1260 35
rect 1280 15 1300 35
rect 1320 15 1410 35
rect 1430 15 1560 35
rect 1580 15 1670 35
rect 1690 15 1740 35
rect 1760 15 1920 35
rect 1940 15 2045 35
rect 2065 15 2170 35
rect 2190 15 2295 35
rect 2315 15 2420 35
rect 2440 15 2505 35
rect -40 1 2505 15
rect -40 0 0 1
rect 1 0 2505 1
rect -40 -1215 830 -1200
rect -40 -1235 -30 -1215
rect -10 -1235 80 -1215
rect 100 -1235 230 -1215
rect 250 -1235 340 -1215
rect 360 -1235 410 -1215
rect 430 -1235 520 -1215
rect 540 -1235 670 -1215
rect 690 -1235 780 -1215
rect 800 -1235 830 -1215
rect -40 -1250 830 -1235
rect 890 -1215 1325 -1200
rect 890 -1235 910 -1215
rect 930 -1235 1090 -1215
rect 1110 -1235 1215 -1215
rect 1235 -1235 1325 -1215
rect 890 -1250 1325 -1235
rect -40 -1375 830 -1360
rect -40 -1445 -30 -1375
rect -10 -1445 340 -1375
rect 360 -1445 410 -1375
rect 430 -1445 780 -1375
rect 800 -1445 830 -1375
rect -40 -1460 830 -1445
rect 890 -1375 1325 -1360
rect 890 -1445 965 -1375
rect 985 -1445 1090 -1375
rect 1110 -1445 1215 -1375
rect 1235 -1445 1325 -1375
rect 890 -1460 1325 -1445
rect -40 -1755 830 -1740
rect -40 -1825 -30 -1755
rect -10 -1825 340 -1755
rect 360 -1825 410 -1755
rect 430 -1825 780 -1755
rect 800 -1825 830 -1755
rect -40 -1840 830 -1825
rect 950 -1755 1300 -1740
rect 950 -1825 1015 -1755
rect 1035 -1825 1140 -1755
rect 1160 -1825 1265 -1755
rect 1285 -1825 1300 -1755
rect 950 -1840 1300 -1825
rect -40 -1965 830 -1950
rect -40 -1985 -30 -1965
rect -10 -1985 80 -1965
rect 100 -1985 230 -1965
rect 250 -1985 340 -1965
rect 360 -1985 410 -1965
rect 430 -1985 520 -1965
rect 540 -1985 670 -1965
rect 690 -1985 780 -1965
rect 800 -1985 830 -1965
rect -40 -2000 830 -1985
rect 950 -1965 1300 -1950
rect 950 -1985 1015 -1965
rect 1035 -1985 1140 -1965
rect 1160 -1985 1265 -1965
rect 1285 -1985 1300 -1965
rect 950 -2000 1300 -1985
rect -190 -2550 1350 -2540
rect -190 -2570 -170 -2550
rect -150 -2570 -120 -2550
rect -100 -2570 -70 -2550
rect -50 -2570 -20 -2550
rect 0 -2570 30 -2550
rect 50 -2570 80 -2550
rect 100 -2570 130 -2550
rect 150 -2570 180 -2550
rect 200 -2570 230 -2550
rect 250 -2570 280 -2550
rect 300 -2570 340 -2550
rect 360 -2570 390 -2550
rect 410 -2570 440 -2550
rect 460 -2570 490 -2550
rect 510 -2570 540 -2550
rect 560 -2570 590 -2550
rect 610 -2570 640 -2550
rect 660 -2570 690 -2550
rect 710 -2570 740 -2550
rect 760 -2570 790 -2550
rect 810 -2570 840 -2550
rect 860 -2570 890 -2550
rect 910 -2570 980 -2550
rect 1000 -2570 1030 -2550
rect 1050 -2570 1080 -2550
rect 1100 -2570 1170 -2550
rect 1190 -2570 1220 -2550
rect 1240 -2570 1270 -2550
rect 1290 -2570 1350 -2550
rect -190 -2580 1350 -2570
rect 1450 -2550 2270 -2540
rect 1450 -2570 1470 -2550
rect 1490 -2570 1520 -2550
rect 1540 -2570 1570 -2550
rect 1590 -2570 1620 -2550
rect 1640 -2570 1670 -2550
rect 1690 -2570 1720 -2550
rect 1740 -2570 1770 -2550
rect 1790 -2570 1820 -2550
rect 1840 -2570 1870 -2550
rect 1890 -2570 1920 -2550
rect 1940 -2570 1970 -2550
rect 1990 -2570 2020 -2550
rect 2040 -2570 2070 -2550
rect 2090 -2570 2120 -2550
rect 2140 -2570 2170 -2550
rect 2190 -2570 2220 -2550
rect 2240 -2570 2270 -2550
rect 1450 -2580 2270 -2570
rect 75 -2605 115 -2595
rect 75 -2625 85 -2605
rect 105 -2615 115 -2605
rect 880 -2605 920 -2595
rect 880 -2615 890 -2605
rect 105 -2625 890 -2615
rect 910 -2615 920 -2605
rect 910 -2625 1325 -2615
rect 75 -2635 1325 -2625
rect 720 -2775 760 -2770
rect 720 -2805 725 -2775
rect 755 -2805 760 -2775
rect 720 -2810 760 -2805
rect 1250 -2795 1290 -2790
rect 1250 -2825 1255 -2795
rect 1285 -2825 1290 -2795
rect 1250 -2830 1290 -2825
rect 795 -3080 835 -3075
rect 795 -3110 800 -3080
rect 830 -3110 835 -3080
rect 795 -3115 835 -3110
rect -190 -3140 1345 -3130
rect -190 -3160 -170 -3140
rect -150 -3160 -120 -3140
rect -100 -3160 -70 -3140
rect -50 -3160 -20 -3140
rect 0 -3160 30 -3140
rect 50 -3160 80 -3140
rect 100 -3160 130 -3140
rect 150 -3160 180 -3140
rect 200 -3160 230 -3140
rect 250 -3160 280 -3140
rect 300 -3160 340 -3140
rect 360 -3160 390 -3140
rect 410 -3160 440 -3140
rect 460 -3160 490 -3140
rect 510 -3160 540 -3140
rect 560 -3160 590 -3140
rect 610 -3160 640 -3140
rect 660 -3160 690 -3140
rect 710 -3160 740 -3140
rect 760 -3160 790 -3140
rect 810 -3160 840 -3140
rect 860 -3160 890 -3140
rect 910 -3160 980 -3140
rect 1000 -3160 1030 -3140
rect 1050 -3160 1080 -3140
rect 1100 -3160 1170 -3140
rect 1190 -3160 1220 -3140
rect 1240 -3160 1270 -3140
rect 1290 -3160 1345 -3140
rect -190 -3170 1345 -3160
rect 1450 -3140 2270 -3130
rect 1450 -3160 1470 -3140
rect 1490 -3160 1520 -3140
rect 1540 -3160 1570 -3140
rect 1590 -3160 1620 -3140
rect 1640 -3160 1670 -3140
rect 1690 -3160 1720 -3140
rect 1740 -3160 1770 -3140
rect 1790 -3160 1820 -3140
rect 1840 -3160 1870 -3140
rect 1890 -3160 1920 -3140
rect 1940 -3160 1970 -3140
rect 1990 -3160 2020 -3140
rect 2040 -3160 2070 -3140
rect 2090 -3160 2120 -3140
rect 2140 -3160 2170 -3140
rect 2190 -3160 2220 -3140
rect 2240 -3160 2270 -3140
rect 1450 -3170 2270 -3160
rect 1745 -3175 1785 -3170
rect 95 -3195 135 -3185
rect 95 -3215 105 -3195
rect 125 -3200 135 -3195
rect 1685 -3190 1725 -3185
rect 125 -3205 1350 -3200
rect 125 -3215 785 -3205
rect 95 -3220 785 -3215
rect 95 -3225 135 -3220
rect 780 -3235 785 -3220
rect 815 -3220 1350 -3205
rect 1685 -3220 1690 -3190
rect 1720 -3220 1725 -3190
rect 1745 -3205 1750 -3175
rect 1780 -3205 1785 -3175
rect 2035 -3175 2075 -3170
rect 1745 -3210 1785 -3205
rect 1975 -3190 2015 -3185
rect 815 -3235 820 -3220
rect 1685 -3225 1725 -3220
rect 1975 -3220 1980 -3190
rect 2010 -3220 2015 -3190
rect 2035 -3205 2040 -3175
rect 2070 -3205 2075 -3175
rect 2035 -3210 2075 -3205
rect 1975 -3225 2015 -3220
rect 780 -3240 820 -3235
rect 730 -3475 770 -3470
rect 730 -3505 735 -3475
rect 765 -3505 770 -3475
rect 730 -3510 770 -3505
rect 1270 -3475 1310 -3470
rect 1270 -3505 1275 -3475
rect 1305 -3505 1310 -3475
rect 1270 -3510 1310 -3505
rect 1685 -3680 1705 -3645
rect 1665 -3685 1705 -3680
rect 1665 -3715 1670 -3685
rect 1700 -3715 1705 -3685
rect 1725 -3670 1765 -3665
rect 1725 -3700 1730 -3670
rect 1760 -3700 1765 -3670
rect 1975 -3680 1995 -3645
rect 1725 -3705 1765 -3700
rect 1955 -3685 1995 -3680
rect 1665 -3720 1705 -3715
rect 1955 -3715 1960 -3685
rect 1990 -3715 1995 -3685
rect 2015 -3670 2055 -3665
rect 2015 -3700 2020 -3670
rect 2050 -3700 2055 -3670
rect 2015 -3705 2055 -3700
rect 1955 -3720 1995 -3715
rect -190 -3730 1320 -3720
rect -190 -3750 -170 -3730
rect -150 -3750 -120 -3730
rect -100 -3750 -70 -3730
rect -50 -3750 -20 -3730
rect 0 -3750 30 -3730
rect 50 -3750 80 -3730
rect 100 -3750 130 -3730
rect 150 -3750 180 -3730
rect 200 -3750 230 -3730
rect 250 -3750 280 -3730
rect 300 -3750 340 -3730
rect 360 -3750 390 -3730
rect 410 -3750 440 -3730
rect 460 -3750 490 -3730
rect 510 -3750 540 -3730
rect 560 -3750 590 -3730
rect 610 -3750 640 -3730
rect 660 -3750 690 -3730
rect 710 -3750 740 -3730
rect 760 -3750 790 -3730
rect 810 -3750 840 -3730
rect 860 -3750 890 -3730
rect 910 -3750 980 -3730
rect 1000 -3750 1030 -3730
rect 1050 -3750 1080 -3730
rect 1100 -3750 1170 -3730
rect 1190 -3750 1220 -3730
rect 1240 -3750 1270 -3730
rect 1290 -3750 1320 -3730
rect -190 -3760 1320 -3750
rect 1450 -3730 2270 -3720
rect 1450 -3750 1470 -3730
rect 1490 -3750 1520 -3730
rect 1540 -3750 1570 -3730
rect 1590 -3750 1620 -3730
rect 1640 -3750 1670 -3730
rect 1690 -3750 1720 -3730
rect 1740 -3750 1770 -3730
rect 1790 -3750 1820 -3730
rect 1840 -3750 1870 -3730
rect 1890 -3750 1920 -3730
rect 1940 -3750 1970 -3730
rect 1990 -3750 2020 -3730
rect 2040 -3750 2070 -3730
rect 2090 -3750 2120 -3730
rect 2140 -3750 2170 -3730
rect 2190 -3750 2220 -3730
rect 2240 -3750 2270 -3730
rect 1450 -3760 2270 -3750
rect 1450 -4910 2270 -4900
rect 1450 -4930 1470 -4910
rect 1490 -4930 1520 -4910
rect 1540 -4930 1570 -4910
rect 1590 -4930 1620 -4910
rect 1640 -4930 1670 -4910
rect 1690 -4930 1720 -4910
rect 1740 -4930 1770 -4910
rect 1790 -4930 1820 -4910
rect 1840 -4930 1870 -4910
rect 1890 -4930 1920 -4910
rect 1940 -4930 1970 -4910
rect 1990 -4930 2020 -4910
rect 2040 -4930 2070 -4910
rect 2090 -4930 2120 -4910
rect 2140 -4930 2170 -4910
rect 2190 -4930 2220 -4910
rect 2240 -4930 2270 -4910
rect 1450 -4940 2270 -4930
rect 1450 -5610 2270 -5600
rect 1450 -5630 1470 -5610
rect 1490 -5630 1520 -5610
rect 1540 -5630 1570 -5610
rect 1590 -5630 1620 -5610
rect 1640 -5630 1670 -5610
rect 1690 -5630 1720 -5610
rect 1740 -5630 1770 -5610
rect 1790 -5630 1820 -5610
rect 1840 -5630 1870 -5610
rect 1890 -5630 1920 -5610
rect 1940 -5630 1970 -5610
rect 1990 -5630 2020 -5610
rect 2040 -5630 2070 -5610
rect 2090 -5630 2120 -5610
rect 2140 -5630 2170 -5610
rect 2190 -5630 2220 -5610
rect 2240 -5630 2270 -5610
rect 1450 -5640 2270 -5630
rect 1450 -6215 2270 -6205
rect 1450 -6235 1470 -6215
rect 1490 -6235 1520 -6215
rect 1540 -6235 1570 -6215
rect 1590 -6235 1620 -6215
rect 1640 -6235 1670 -6215
rect 1690 -6235 1720 -6215
rect 1740 -6235 1770 -6215
rect 1790 -6235 1820 -6215
rect 1840 -6235 1870 -6215
rect 1890 -6235 1920 -6215
rect 1940 -6235 1970 -6215
rect 1990 -6235 2020 -6215
rect 2040 -6235 2070 -6215
rect 2090 -6235 2120 -6215
rect 2140 -6235 2170 -6215
rect 2190 -6235 2220 -6215
rect 2240 -6235 2270 -6215
rect 1450 -6245 2270 -6235
<< via1 >>
rect 725 -2780 755 -2775
rect 725 -2800 730 -2780
rect 730 -2800 750 -2780
rect 750 -2800 755 -2780
rect 725 -2805 755 -2800
rect 1255 -2800 1285 -2795
rect 1255 -2820 1260 -2800
rect 1260 -2820 1280 -2800
rect 1280 -2820 1285 -2800
rect 1255 -2825 1285 -2820
rect 800 -3085 830 -3080
rect 800 -3105 805 -3085
rect 805 -3105 825 -3085
rect 825 -3105 830 -3085
rect 800 -3110 830 -3105
rect 785 -3235 815 -3205
rect 1690 -3195 1720 -3190
rect 1690 -3215 1695 -3195
rect 1695 -3215 1715 -3195
rect 1715 -3215 1720 -3195
rect 1690 -3220 1720 -3215
rect 1750 -3205 1780 -3175
rect 1980 -3195 2010 -3190
rect 1980 -3215 1985 -3195
rect 1985 -3215 2005 -3195
rect 2005 -3215 2010 -3195
rect 1980 -3220 2010 -3215
rect 2040 -3205 2070 -3175
rect 735 -3480 765 -3475
rect 735 -3500 740 -3480
rect 740 -3500 760 -3480
rect 760 -3500 765 -3480
rect 735 -3505 765 -3500
rect 1275 -3480 1305 -3475
rect 1275 -3500 1280 -3480
rect 1280 -3500 1300 -3480
rect 1300 -3500 1305 -3480
rect 1275 -3505 1305 -3500
rect 1670 -3715 1700 -3685
rect 1730 -3675 1760 -3670
rect 1730 -3695 1735 -3675
rect 1735 -3695 1755 -3675
rect 1755 -3695 1760 -3675
rect 1730 -3700 1760 -3695
rect 1960 -3715 1990 -3685
rect 2020 -3675 2050 -3670
rect 2020 -3695 2025 -3675
rect 2025 -3695 2045 -3675
rect 2045 -3695 2050 -3675
rect 2020 -3700 2050 -3695
<< metal2 >>
rect 720 -2775 760 -2770
rect 720 -2805 725 -2775
rect 755 -2805 760 -2775
rect 720 -2810 760 -2805
rect 740 -3470 760 -2810
rect 1250 -2795 1310 -2790
rect 1250 -2825 1255 -2795
rect 1285 -2825 1310 -2795
rect 1250 -2830 1310 -2825
rect 795 -3080 835 -3075
rect 795 -3110 800 -3080
rect 830 -3110 835 -3080
rect 795 -3115 835 -3110
rect 795 -3200 815 -3115
rect 780 -3205 820 -3200
rect 780 -3235 785 -3205
rect 815 -3235 820 -3205
rect 780 -3240 820 -3235
rect 1290 -3470 1310 -2830
rect 1745 -3175 1785 -3170
rect 730 -3475 770 -3470
rect 730 -3505 735 -3475
rect 765 -3505 770 -3475
rect 730 -3510 770 -3505
rect 1270 -3475 1310 -3470
rect 1270 -3505 1275 -3475
rect 1305 -3505 1310 -3475
rect 1270 -3510 1310 -3505
rect 1685 -3190 1725 -3185
rect 1685 -3220 1690 -3190
rect 1720 -3220 1725 -3190
rect 1685 -3225 1725 -3220
rect 1745 -3205 1750 -3175
rect 1780 -3205 1785 -3175
rect 2035 -3175 2075 -3170
rect 1745 -3210 1785 -3205
rect 1975 -3190 2015 -3185
rect 1685 -3680 1705 -3225
rect 1745 -3665 1765 -3210
rect 1665 -3685 1705 -3680
rect 1665 -3715 1670 -3685
rect 1700 -3715 1705 -3685
rect 1725 -3670 1765 -3665
rect 1725 -3700 1730 -3670
rect 1760 -3700 1765 -3670
rect 1975 -3220 1980 -3190
rect 2010 -3220 2015 -3190
rect 1975 -3225 2015 -3220
rect 2035 -3205 2040 -3175
rect 2070 -3205 2075 -3175
rect 2035 -3210 2075 -3205
rect 1975 -3680 1995 -3225
rect 2035 -3665 2055 -3210
rect 1725 -3705 1765 -3700
rect 1955 -3685 1995 -3680
rect 1665 -3720 1705 -3715
rect 1955 -3715 1960 -3685
rect 1990 -3715 1995 -3685
rect 2015 -3670 2055 -3665
rect 2015 -3700 2020 -3670
rect 2050 -3700 2055 -3670
rect 2015 -3705 2055 -3700
rect 1955 -3720 1995 -3715
<< labels >>
flabel poly -60 95 -60 95 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel poly 150 125 150 125 7 FreeSans 160 0 -80 0 QA_b
flabel locali 540 125 540 125 3 FreeSans 160 0 80 0 E
flabel locali 745 125 745 125 3 FreeSans 160 0 80 0 E_b
flabel poly 770 325 770 325 3 FreeSans 160 0 80 0 Reset
flabel locali 1905 130 1905 130 3 FreeSans 160 0 80 0 before_Reset
flabel poly -60 -85 -60 -85 7 FreeSans 160 0 -80 0 F_VCO
port 2 w
flabel poly 1030 135 1030 135 7 FreeSans 160 0 -80 0 QB_b
flabel locali 1430 125 1430 125 3 FreeSans 160 0 80 0 F
flabel locali 1635 110 1635 110 3 FreeSans 160 0 80 0 F_b
flabel metal1 -40 25 -40 25 7 FreeSans 160 0 -80 0 GNDA
port 6 w
flabel metal1 -40 210 -40 210 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel locali 2530 285 2530 285 3 FreeSans 160 0 80 0 QA
port 4 e
flabel locali 2530 -25 2530 -25 3 FreeSans 160 0 80 0 QB
port 5 e
flabel poly -60 -1295 -60 -1295 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel poly 150 -1325 150 -1325 7 FreeSans 160 0 -80 0 QA_b
flabel locali 540 -1325 540 -1325 3 FreeSans 160 0 80 0 E
flabel locali 745 -1325 745 -1325 3 FreeSans 160 0 80 0 E_b
flabel metal1 -40 -1225 -40 -1225 7 FreeSans 160 0 -80 0 GNDA
port 6 w
flabel metal1 -40 -1410 -40 -1410 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel locali 1075 -1330 1075 -1330 3 FreeSans 160 0 80 0 before_Reset
flabel poly 60 -2825 60 -2825 7 FreeSans 160 0 -80 0 QA_b
flabel poly -150 -2795 -150 -2795 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel locali 665 -2825 665 -2825 3 FreeSans 160 0 80 0 E_b
flabel locali 460 -2825 460 -2825 3 FreeSans 160 0 80 0 E
<< end >>
