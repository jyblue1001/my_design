magic
tech sky130A
timestamp 1723040051
<< nwell >>
rect -75 630 460 985
<< nmos >>
rect -5 425 10 525
rect 35 425 50 525
rect 100 425 115 525
rect 245 425 260 525
rect 310 425 325 525
rect 375 425 390 525
rect -5 210 10 310
rect 35 210 50 310
rect 100 210 115 310
rect 245 210 260 310
rect 310 210 325 310
rect 375 210 390 310
<< pmos >>
rect -5 865 10 965
rect 60 865 75 965
rect 125 865 140 965
rect 270 865 285 965
rect 310 865 325 965
rect 375 865 390 965
rect -5 650 10 750
rect 60 650 75 750
rect 125 650 140 750
rect 270 650 285 750
rect 310 650 325 750
rect 375 650 390 750
<< ndiff >>
rect -55 510 -5 525
rect -55 440 -40 510
rect -20 440 -5 510
rect -55 425 -5 440
rect 10 425 35 525
rect 50 510 100 525
rect 50 440 65 510
rect 85 440 100 510
rect 50 425 100 440
rect 115 510 165 525
rect 115 440 130 510
rect 150 440 165 510
rect 115 425 165 440
rect 195 510 245 525
rect 195 440 210 510
rect 230 440 245 510
rect 195 425 245 440
rect 260 510 310 525
rect 260 440 275 510
rect 295 440 310 510
rect 260 425 310 440
rect 325 510 375 525
rect 325 440 340 510
rect 360 440 375 510
rect 325 425 375 440
rect 390 510 440 525
rect 390 440 405 510
rect 425 440 440 510
rect 390 425 440 440
rect -55 295 -5 310
rect -55 225 -40 295
rect -20 225 -5 295
rect -55 210 -5 225
rect 10 210 35 310
rect 50 295 100 310
rect 50 225 65 295
rect 85 225 100 295
rect 50 210 100 225
rect 115 295 165 310
rect 115 225 130 295
rect 150 225 165 295
rect 115 210 165 225
rect 195 295 245 310
rect 195 225 210 295
rect 230 225 245 295
rect 195 210 245 225
rect 260 295 310 310
rect 260 225 275 295
rect 295 225 310 295
rect 260 210 310 225
rect 325 295 375 310
rect 325 225 340 295
rect 360 225 375 295
rect 325 210 375 225
rect 390 295 440 310
rect 390 225 405 295
rect 425 225 440 295
rect 390 210 440 225
<< pdiff >>
rect -55 950 -5 965
rect -55 880 -40 950
rect -20 880 -5 950
rect -55 865 -5 880
rect 10 950 60 965
rect 10 880 25 950
rect 45 880 60 950
rect 10 865 60 880
rect 75 950 125 965
rect 75 880 90 950
rect 110 880 125 950
rect 75 865 125 880
rect 140 950 190 965
rect 140 880 155 950
rect 175 880 190 950
rect 140 865 190 880
rect 220 950 270 965
rect 220 880 235 950
rect 255 880 270 950
rect 220 865 270 880
rect 285 865 310 965
rect 325 950 375 965
rect 325 880 340 950
rect 360 880 375 950
rect 325 865 375 880
rect 390 950 440 965
rect 390 880 405 950
rect 425 880 440 950
rect 390 865 440 880
rect -55 735 -5 750
rect -55 665 -40 735
rect -20 665 -5 735
rect -55 650 -5 665
rect 10 735 60 750
rect 10 665 25 735
rect 45 665 60 735
rect 10 650 60 665
rect 75 735 125 750
rect 75 665 90 735
rect 110 665 125 735
rect 75 650 125 665
rect 140 735 190 750
rect 140 665 155 735
rect 175 665 190 735
rect 140 650 190 665
rect 220 735 270 750
rect 220 665 235 735
rect 255 665 270 735
rect 220 650 270 665
rect 285 650 310 750
rect 325 735 375 750
rect 325 665 340 735
rect 360 665 375 735
rect 325 650 375 665
rect 390 735 440 750
rect 390 665 405 735
rect 425 665 440 735
rect 390 650 440 665
<< ndiffc >>
rect -40 440 -20 510
rect 65 440 85 510
rect 130 440 150 510
rect 210 440 230 510
rect 275 440 295 510
rect 340 440 360 510
rect 405 440 425 510
rect -40 225 -20 295
rect 65 225 85 295
rect 130 225 150 295
rect 210 225 230 295
rect 275 225 295 295
rect 340 225 360 295
rect 405 225 425 295
<< pdiffc >>
rect -40 880 -20 950
rect 25 880 45 950
rect 90 880 110 950
rect 155 880 175 950
rect 235 880 255 950
rect 340 880 360 950
rect 405 880 425 950
rect -40 665 -20 735
rect 25 665 45 735
rect 90 665 110 735
rect 155 665 175 735
rect 235 665 255 735
rect 340 665 360 735
rect 405 665 425 735
<< psubdiff >>
rect 195 380 295 395
rect 195 360 210 380
rect 280 360 295 380
rect 195 345 295 360
<< nsubdiff >>
rect -55 815 45 830
rect -55 795 -40 815
rect 30 795 45 815
rect -55 780 45 795
<< psubdiffcont >>
rect 210 360 280 380
<< nsubdiffcont >>
rect -40 795 30 815
<< poly >>
rect 350 1010 390 1020
rect 350 990 360 1010
rect 380 990 390 1010
rect 350 980 390 990
rect -5 965 10 980
rect 60 965 75 980
rect 125 965 140 980
rect 270 965 285 980
rect 310 965 325 980
rect 375 965 390 980
rect -5 855 10 865
rect -65 840 10 855
rect -5 750 10 765
rect 60 750 75 865
rect 125 850 140 865
rect 270 850 285 865
rect 100 840 140 850
rect 100 820 110 840
rect 130 820 140 840
rect 100 810 140 820
rect 165 840 285 850
rect 165 820 175 840
rect 195 835 285 840
rect 195 820 205 835
rect 165 810 205 820
rect 165 780 180 810
rect 125 765 180 780
rect 125 750 140 765
rect 270 750 285 765
rect 310 750 325 865
rect 375 850 390 865
rect 415 840 460 855
rect 415 805 430 840
rect 350 795 430 805
rect 350 775 360 795
rect 380 790 430 795
rect 380 775 390 790
rect 350 765 390 775
rect 375 750 390 765
rect -5 585 10 650
rect 60 640 75 650
rect 125 640 140 650
rect -30 575 10 585
rect -30 555 -20 575
rect 0 555 10 575
rect -30 545 10 555
rect -5 525 10 545
rect 35 625 75 640
rect 100 625 140 640
rect 270 635 285 650
rect 245 625 285 635
rect 35 525 50 625
rect 100 525 115 625
rect 245 605 255 625
rect 275 605 285 625
rect 245 595 285 605
rect 245 525 260 595
rect 310 525 325 650
rect 375 525 390 650
rect -5 410 10 425
rect -65 320 10 335
rect -5 310 10 320
rect 35 310 50 425
rect 100 405 115 425
rect 245 410 260 425
rect 75 395 115 405
rect 75 375 85 395
rect 105 380 115 395
rect 105 375 155 380
rect 75 365 155 375
rect 140 335 155 365
rect 100 310 115 325
rect 140 320 260 335
rect 245 310 260 320
rect 310 310 325 425
rect 375 415 390 425
rect 375 400 430 415
rect 350 355 390 365
rect 350 335 360 355
rect 380 335 390 355
rect 350 325 390 335
rect 375 310 390 325
rect 415 360 430 400
rect 415 350 455 360
rect 415 330 425 350
rect 445 335 455 350
rect 445 330 460 335
rect 415 320 460 330
rect -5 195 10 210
rect 35 155 50 210
rect 100 195 115 210
rect 245 195 260 210
rect 75 185 115 195
rect 75 165 85 185
rect 105 165 115 185
rect 75 155 115 165
rect 310 155 325 210
rect 375 195 390 210
rect 10 145 50 155
rect 10 125 20 145
rect 40 125 50 145
rect 10 115 50 125
rect 285 145 325 155
rect 285 125 295 145
rect 315 125 325 145
rect 285 115 325 125
<< polycont >>
rect 360 990 380 1010
rect 110 820 130 840
rect 175 820 195 840
rect 360 775 380 795
rect -20 555 0 575
rect 255 605 275 625
rect 85 375 105 395
rect 360 335 380 355
rect 425 330 445 350
rect 85 165 105 185
rect 20 125 40 145
rect 295 125 315 145
<< locali >>
rect 350 1010 390 1020
rect 350 1000 360 1010
rect -30 980 100 1000
rect -30 960 -10 980
rect 80 960 100 980
rect 285 990 360 1000
rect 380 990 390 1010
rect 285 980 390 990
rect -50 950 -10 960
rect -50 880 -40 950
rect -20 880 -10 950
rect -50 870 -10 880
rect 15 950 55 960
rect 15 880 25 950
rect 45 880 55 950
rect 15 870 55 880
rect 80 950 120 960
rect 80 880 90 950
rect 110 880 120 950
rect 80 870 120 880
rect 145 950 185 960
rect 145 880 155 950
rect 175 880 185 950
rect 145 870 185 880
rect 15 825 35 870
rect 165 850 185 870
rect 225 950 265 960
rect 225 880 235 950
rect 255 880 265 950
rect 225 870 265 880
rect 100 840 140 850
rect -50 815 40 825
rect -50 795 -40 815
rect 30 795 40 815
rect 100 820 110 840
rect 130 820 140 840
rect 100 810 140 820
rect 165 840 205 850
rect 165 820 175 840
rect 195 820 205 840
rect 165 810 205 820
rect -50 785 40 795
rect 120 790 140 810
rect 15 745 35 785
rect 120 770 165 790
rect 145 745 165 770
rect 225 745 245 870
rect 285 745 305 980
rect 330 950 370 960
rect 330 880 340 950
rect 360 880 370 950
rect 330 870 370 880
rect 395 950 435 960
rect 395 880 405 950
rect 425 880 435 950
rect 395 870 435 880
rect 350 805 370 870
rect 350 795 390 805
rect 350 775 360 795
rect 380 775 390 795
rect 350 765 390 775
rect 415 745 435 870
rect -50 735 -10 745
rect -50 665 -40 735
rect -20 665 -10 735
rect -50 655 -10 665
rect 15 735 55 745
rect 15 665 25 735
rect 45 665 55 735
rect 15 655 55 665
rect 80 735 120 745
rect 80 665 90 735
rect 110 665 120 735
rect 80 655 120 665
rect 145 735 185 745
rect 145 665 155 735
rect 175 665 185 735
rect 145 655 185 665
rect 225 735 265 745
rect 225 665 235 735
rect 255 665 265 735
rect 285 735 370 745
rect 285 725 340 735
rect 225 655 265 665
rect 330 665 340 725
rect 360 665 370 735
rect 330 655 370 665
rect 395 735 435 745
rect 395 665 405 735
rect 425 665 435 735
rect 395 655 435 665
rect -30 635 -10 655
rect 80 635 100 655
rect -30 615 100 635
rect 145 635 165 655
rect 145 625 285 635
rect 145 615 255 625
rect -70 575 10 585
rect -70 565 -20 575
rect -30 555 -20 565
rect 0 555 10 575
rect 145 565 165 615
rect 245 605 255 615
rect 275 605 285 625
rect 245 595 285 605
rect 350 620 370 655
rect 350 600 435 620
rect -30 545 10 555
rect 75 545 165 565
rect 415 585 435 600
rect 415 565 460 585
rect 75 520 95 545
rect 220 540 350 560
rect 220 520 240 540
rect 330 520 350 540
rect 415 520 435 565
rect -50 510 -10 520
rect -50 440 -40 510
rect -20 440 -10 510
rect 55 510 95 520
rect 55 450 65 510
rect -50 430 -10 440
rect 15 440 65 450
rect 85 440 95 510
rect 15 430 95 440
rect 120 510 160 520
rect 120 440 130 510
rect 150 440 160 510
rect 120 430 160 440
rect 200 510 240 520
rect 200 440 210 510
rect 230 440 240 510
rect 200 430 240 440
rect 265 510 305 520
rect 265 440 275 510
rect 295 440 305 510
rect 265 430 305 440
rect 330 510 370 520
rect 330 440 340 510
rect 360 440 370 510
rect 330 430 370 440
rect 395 510 435 520
rect 395 440 405 510
rect 425 440 435 510
rect 395 430 435 440
rect -50 305 -30 430
rect -50 295 -10 305
rect -50 225 -40 295
rect -20 225 -10 295
rect -50 215 -10 225
rect 15 195 35 430
rect 75 395 115 405
rect 75 375 85 395
rect 105 375 115 395
rect 75 365 115 375
rect 140 380 160 430
rect 265 390 285 430
rect 395 410 415 430
rect 370 390 415 410
rect 200 380 290 390
rect 75 305 95 365
rect 140 360 210 380
rect 280 360 290 380
rect 370 365 390 390
rect 140 305 160 360
rect 200 350 290 360
rect 350 355 390 365
rect 265 305 285 350
rect 350 335 360 355
rect 380 335 390 355
rect 350 325 390 335
rect 415 350 455 360
rect 415 330 425 350
rect 445 330 455 350
rect 415 320 455 330
rect 415 305 435 320
rect 55 295 95 305
rect 55 225 65 295
rect 85 225 95 295
rect 55 215 95 225
rect 120 295 160 305
rect 120 225 130 295
rect 150 225 160 295
rect 120 215 160 225
rect 200 295 240 305
rect 200 225 210 295
rect 230 225 240 295
rect 200 215 240 225
rect 265 295 305 305
rect 265 225 275 295
rect 295 225 305 295
rect 265 215 305 225
rect 330 295 370 305
rect 330 225 340 295
rect 360 225 370 295
rect 330 215 370 225
rect 395 295 435 305
rect 395 225 405 295
rect 425 225 435 295
rect 395 215 435 225
rect 220 195 240 215
rect 330 195 350 215
rect 15 185 115 195
rect 15 175 85 185
rect 75 165 85 175
rect 105 165 115 185
rect 220 175 350 195
rect 75 155 115 165
rect 10 145 50 155
rect 10 125 20 145
rect 40 125 50 145
rect 10 115 50 125
rect 285 145 325 155
rect 285 125 295 145
rect 315 125 325 145
rect 285 115 325 125
<< viali >>
rect 25 880 45 950
rect 235 880 255 950
rect -40 795 30 815
rect 405 880 425 950
rect 25 665 45 735
rect 235 665 255 735
rect 405 665 425 735
rect -40 440 -20 510
rect 130 440 150 510
rect 275 440 295 510
rect -40 225 -20 295
rect 210 360 280 380
rect 130 225 150 295
rect 275 225 295 295
rect 20 125 40 145
rect 295 125 315 145
<< metal1 >>
rect -65 950 460 965
rect -65 880 25 950
rect 45 880 235 950
rect 255 880 405 950
rect 425 880 460 950
rect -65 815 460 880
rect -65 795 -40 815
rect 30 795 460 815
rect -65 735 460 795
rect -65 665 25 735
rect 45 665 235 735
rect 255 665 405 735
rect 425 665 460 735
rect -65 650 460 665
rect -65 510 460 525
rect -65 440 -40 510
rect -20 440 130 510
rect 150 440 275 510
rect 295 440 460 510
rect -65 380 460 440
rect -65 360 210 380
rect 280 360 460 380
rect -65 295 460 360
rect -65 225 -40 295
rect -20 225 130 295
rect 150 225 275 295
rect 295 225 460 295
rect -65 210 460 225
rect -65 145 460 155
rect -65 125 20 145
rect 40 125 295 145
rect 315 125 460 145
rect -65 115 460 125
<< labels >>
flabel poly -65 845 -65 845 7 FreeSans 80 0 -40 0 Db1
port 2 w
flabel metal1 -65 805 -65 805 7 FreeSans 80 0 -40 0 VP
port 7 w
flabel metal1 -65 370 -65 370 7 FreeSans 80 0 -40 0 VN
port 8 w
flabel poly -65 325 -65 325 7 FreeSans 80 0 -40 0 Db2
port 3 w
flabel space -65 135 -65 135 7 FreeSans 80 0 -40 0 CLK
port 6 w
flabel poly 460 845 460 845 3 FreeSans 80 0 40 0 Qb1
port 5 e
flabel locali -70 575 -70 575 7 FreeSans 80 0 -40 0 D
port 1 w
flabel locali 460 575 460 575 3 FreeSans 80 0 40 0 Q
port 4 e
<< end >>
