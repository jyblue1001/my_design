magic
tech sky130A
timestamp 1752827747
<< error_s >>
rect 7380 1785 7400 1805
<< metal1 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6655 2990 6685
rect 2950 6650 2990 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6655 6085 6685
rect 3030 6650 3070 6655
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6550 2945 6580
rect 2905 6545 2945 6550
rect 2915 2710 2935 6545
rect 2960 2505 2980 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 3955 6645 3995 6650
rect 3955 6615 3960 6645
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3965 3360 3985 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 4005 6475 4045 6480
rect 4005 6445 4010 6475
rect 4040 6445 4045 6475
rect 4005 6440 4045 6445
rect 3955 3355 3995 3360
rect 3955 3325 3960 3355
rect 3990 3325 3995 3355
rect 3955 3320 3995 3325
rect 4015 2790 4035 6440
rect 5085 5465 5105 6655
rect 5730 6585 5750 6655
rect 6045 6650 6085 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5430 5115 5460
rect 5075 5425 5115 5430
rect 5385 5420 5405 6485
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5385 5415 5415
rect 5375 5380 5415 5385
rect 5495 5415 5535 5420
rect 5495 5385 5500 5415
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 5505 4805 5525 5380
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6055 3640 6075 6650
rect 6100 5460 6140 5465
rect 6100 5430 6105 5460
rect 6135 5430 6140 5460
rect 6785 5440 6805 6655
rect 7020 6650 7060 6655
rect 7100 6685 7140 6690
rect 7100 6655 7105 6685
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 6100 5425 6140 5430
rect 6425 5435 6465 5440
rect 6045 3635 6085 3640
rect 4970 3630 5010 3635
rect 4970 3600 4975 3630
rect 5005 3600 5010 3630
rect 6045 3605 6050 3635
rect 6080 3605 6085 3635
rect 6045 3600 6085 3605
rect 4970 3595 5010 3600
rect 6110 2880 6130 5425
rect 6425 5405 6430 5435
rect 6460 5405 6465 5435
rect 6425 5400 6465 5405
rect 6775 5435 6815 5440
rect 6775 5405 6780 5435
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 6435 4870 6455 5400
rect 6425 4865 6465 4870
rect 6425 4835 6430 4865
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 5085 2875 5125 2880
rect 5085 2845 5090 2875
rect 5120 2845 5125 2875
rect 5085 2840 5125 2845
rect 6100 2875 6140 2880
rect 6100 2845 6105 2875
rect 6135 2845 6140 2875
rect 6100 2840 6140 2845
rect 5095 2410 5115 2840
rect 7110 2505 7130 6650
rect 7145 6580 7185 6585
rect 7145 6550 7150 6580
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 7155 2710 7175 6545
rect 2440 1800 2480 1830
<< via1 >>
rect 2955 6655 2985 6685
rect 3035 6655 3065 6685
rect 6050 6655 6080 6685
rect 2910 6550 2940 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 3960 6615 3990 6645
rect 3550 6445 3580 6475
rect 4335 6550 4365 6580
rect 4010 6445 4040 6475
rect 3960 3325 3990 3355
rect 6705 6655 6735 6685
rect 7025 6655 7055 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 5080 5430 5110 5460
rect 5380 5385 5410 5415
rect 5500 5385 5530 5415
rect 5500 4770 5530 4800
rect 6105 5430 6135 5460
rect 7105 6655 7135 6685
rect 4975 3600 5005 3630
rect 6050 3605 6080 3635
rect 6430 5405 6460 5435
rect 6780 5405 6810 5435
rect 6430 4835 6460 4865
rect 5090 2845 5120 2875
rect 6105 2845 6135 2875
rect 7150 6550 7180 6580
<< metal2 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6680 2990 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2985 6660 3035 6680
rect 2985 6655 2990 6660
rect 2950 6650 2990 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6680 6085 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6080 6660 6705 6680
rect 6080 6655 6085 6660
rect 6045 6650 6085 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6680 7025 6685
rect 7010 6660 7025 6680
rect 6700 6650 6740 6655
rect 7020 6655 7025 6660
rect 7055 6680 7060 6685
rect 7100 6685 7140 6690
rect 7100 6680 7105 6685
rect 7055 6660 7105 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7100 6655 7105 6660
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 3955 6645 3995 6650
rect 3955 6640 3960 6645
rect 3435 6620 3960 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 3955 6615 3960 6620
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6575 2945 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2940 6555 4335 6575
rect 2940 6550 2945 6555
rect 2905 6545 2945 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7145 6580 7185 6585
rect 7145 6575 7150 6580
rect 5755 6555 7150 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7145 6550 7150 6555
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 4005 6475 4045 6480
rect 4005 6470 4010 6475
rect 3580 6450 4010 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 4005 6445 4010 6450
rect 4040 6445 4045 6475
rect 4005 6440 4045 6445
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5455 5115 5460
rect 6100 5460 6140 5465
rect 6100 5455 6105 5460
rect 5110 5435 6105 5455
rect 5110 5430 5115 5435
rect 5075 5425 5115 5430
rect 6100 5430 6105 5435
rect 6135 5430 6140 5460
rect 6100 5425 6140 5430
rect 6425 5435 6465 5440
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5410 5415 5415
rect 5495 5415 5535 5420
rect 5495 5410 5500 5415
rect 5410 5390 5500 5410
rect 5410 5385 5415 5390
rect 5375 5380 5415 5385
rect 5495 5385 5500 5390
rect 5530 5385 5535 5415
rect 6425 5405 6430 5435
rect 6460 5430 6465 5435
rect 6775 5435 6815 5440
rect 6775 5430 6780 5435
rect 6460 5410 6780 5430
rect 6460 5405 6465 5410
rect 6425 5400 6465 5405
rect 6775 5405 6780 5410
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 5495 5380 5535 5385
rect 6425 4865 6465 4870
rect 6425 4860 6430 4865
rect 5750 4840 6430 4860
rect 6425 4835 6430 4840
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6045 3635 6085 3640
rect 4970 3630 5010 3635
rect 4970 3600 4975 3630
rect 5005 3625 5010 3630
rect 6045 3625 6050 3635
rect 5005 3605 6050 3625
rect 6080 3605 6085 3635
rect 5005 3600 5010 3605
rect 6045 3600 6085 3605
rect 4970 3595 5010 3600
rect 3955 3355 3995 3360
rect 3955 3325 3960 3355
rect 3990 3340 3995 3355
rect 3990 3325 4115 3340
rect 3955 3320 4115 3325
rect 5085 2875 5125 2880
rect 5085 2845 5090 2875
rect 5120 2870 5125 2875
rect 6100 2875 6140 2880
rect 6100 2870 6105 2875
rect 5120 2850 6105 2870
rect 5120 2845 5125 2850
rect 5085 2840 5125 2845
rect 6100 2845 6105 2850
rect 6135 2845 6140 2875
rect 6100 2840 6140 2845
rect 4160 2315 4180 2335
rect 5910 2315 5930 2335
rect 2440 1800 2480 1830
rect 2645 1785 2665 1805
rect 7380 1785 7400 1805
<< metal3 >>
rect 9685 14460 9735 14465
rect 9685 14420 9690 14460
rect 9730 14420 9735 14460
rect 9685 14415 9735 14420
rect 9690 50 9730 14415
rect 9685 45 9735 50
rect 9685 5 9690 45
rect 9730 5 9735 45
rect 9685 0 9735 5
<< via3 >>
rect 9690 14420 9730 14460
rect 9690 5 9730 45
<< metal4 >>
rect 7255 14460 9735 14465
rect 7255 14420 9690 14460
rect 9730 14420 9735 14460
rect 7255 14415 9735 14420
rect 540 6700 590 6750
rect 540 0 590 50
rect 9685 45 9735 50
rect 9685 5 9690 45
rect 9730 5 9735 45
rect 9685 0 9735 5
use bgr  bgr_0
timestamp 1752419158
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic_21  two_stage_opamp_dummy_magic_21_0
timestamp 1752827590
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 565 0 565 0 5 FreeSans 800 0 0 -320 GNDA
port 2 s
flabel metal4 565 6750 565 6750 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 4160 2325 4160 2325 7 FreeSans 800 0 -320 0 VIN+
port 5 w
flabel metal2 5930 2325 5930 2325 3 FreeSans 800 0 320 0 VIN-
port 6 e
flabel metal2 2655 1785 2655 1785 5 FreeSans 800 0 0 -320 VOUT+
port 3 s
flabel metal2 7390 1785 7390 1785 5 FreeSans 800 0 0 -320 VOUT-
port 4 s
<< end >>
