magic
tech sky130A
timestamp 1738417841
<< nwell >>
rect 585 105 1945 210
<< nmos >>
rect 645 -35 660 15
rect 700 -35 715 15
rect 755 -35 770 15
rect 920 -35 935 15
rect 975 -35 990 15
rect 1030 -35 1045 15
rect 1085 -35 1100 15
rect 1250 -35 1265 15
rect 1305 -35 1320 15
rect 1360 -35 1375 15
rect 1525 -35 1540 15
rect 1580 -35 1595 15
rect 1635 -35 1650 15
rect 1690 -35 1705 15
rect 1815 -35 1830 15
<< pmos >>
rect 645 125 660 175
rect 700 125 715 175
rect 825 125 840 175
rect 880 125 895 175
rect 1050 125 1065 175
rect 1305 125 1320 175
rect 1360 125 1375 175
rect 1525 125 1540 175
rect 1580 125 1595 175
rect 1815 125 1830 175
rect 1870 125 1885 175
<< ndiff >>
rect 605 0 645 15
rect 605 -20 615 0
rect 635 -20 645 0
rect 605 -35 645 -20
rect 660 0 700 15
rect 660 -20 670 0
rect 690 -20 700 0
rect 660 -35 700 -20
rect 715 0 755 15
rect 715 -20 725 0
rect 745 -20 755 0
rect 715 -35 755 -20
rect 770 0 810 15
rect 770 -20 780 0
rect 800 -20 810 0
rect 770 -35 810 -20
rect 880 0 920 15
rect 880 -20 890 0
rect 910 -20 920 0
rect 880 -35 920 -20
rect 935 0 975 15
rect 935 -20 945 0
rect 965 -20 975 0
rect 935 -35 975 -20
rect 990 0 1030 15
rect 990 -20 1000 0
rect 1020 -20 1030 0
rect 990 -35 1030 -20
rect 1045 0 1085 15
rect 1045 -20 1055 0
rect 1075 -20 1085 0
rect 1045 -35 1085 -20
rect 1100 0 1140 15
rect 1100 -20 1110 0
rect 1130 -20 1140 0
rect 1100 -35 1140 -20
rect 1210 0 1250 15
rect 1210 -20 1220 0
rect 1240 -20 1250 0
rect 1210 -35 1250 -20
rect 1265 0 1305 15
rect 1265 -20 1275 0
rect 1295 -20 1305 0
rect 1265 -35 1305 -20
rect 1320 0 1360 15
rect 1320 -20 1330 0
rect 1350 -20 1360 0
rect 1320 -35 1360 -20
rect 1375 0 1415 15
rect 1375 -20 1385 0
rect 1405 -20 1415 0
rect 1375 -35 1415 -20
rect 1485 0 1525 15
rect 1485 -20 1495 0
rect 1515 -20 1525 0
rect 1485 -35 1525 -20
rect 1540 0 1580 15
rect 1540 -20 1550 0
rect 1570 -20 1580 0
rect 1540 -35 1580 -20
rect 1595 0 1635 15
rect 1595 -20 1605 0
rect 1625 -20 1635 0
rect 1595 -35 1635 -20
rect 1650 0 1690 15
rect 1650 -20 1660 0
rect 1680 -20 1690 0
rect 1650 -35 1690 -20
rect 1705 0 1745 15
rect 1705 -20 1715 0
rect 1735 -20 1745 0
rect 1705 -35 1745 -20
rect 1775 0 1815 15
rect 1775 -20 1785 0
rect 1805 -20 1815 0
rect 1775 -35 1815 -20
rect 1830 0 1870 15
rect 1830 -20 1840 0
rect 1860 -20 1870 0
rect 1830 -35 1870 -20
<< pdiff >>
rect 605 160 645 175
rect 605 140 615 160
rect 635 140 645 160
rect 605 125 645 140
rect 660 160 700 175
rect 660 140 670 160
rect 690 140 700 160
rect 660 125 700 140
rect 715 160 755 175
rect 715 140 725 160
rect 745 140 755 160
rect 715 125 755 140
rect 785 160 825 175
rect 785 140 795 160
rect 815 140 825 160
rect 785 125 825 140
rect 840 160 880 175
rect 840 140 850 160
rect 870 140 880 160
rect 840 125 880 140
rect 895 160 935 175
rect 895 140 905 160
rect 925 140 935 160
rect 895 125 935 140
rect 1010 160 1050 175
rect 1010 140 1020 160
rect 1040 140 1050 160
rect 1010 125 1050 140
rect 1065 160 1105 175
rect 1065 140 1075 160
rect 1095 140 1105 160
rect 1065 125 1105 140
rect 1265 160 1305 175
rect 1265 140 1275 160
rect 1295 140 1305 160
rect 1265 125 1305 140
rect 1320 160 1360 175
rect 1320 140 1330 160
rect 1350 140 1360 160
rect 1320 125 1360 140
rect 1375 160 1415 175
rect 1375 140 1385 160
rect 1405 140 1415 160
rect 1375 125 1415 140
rect 1485 160 1525 175
rect 1485 140 1495 160
rect 1515 140 1525 160
rect 1485 125 1525 140
rect 1540 160 1580 175
rect 1540 140 1550 160
rect 1570 140 1580 160
rect 1540 125 1580 140
rect 1595 160 1635 175
rect 1595 140 1605 160
rect 1625 140 1635 160
rect 1595 125 1635 140
rect 1775 160 1815 175
rect 1775 140 1785 160
rect 1805 140 1815 160
rect 1775 125 1815 140
rect 1830 160 1870 175
rect 1830 140 1840 160
rect 1860 140 1870 160
rect 1830 125 1870 140
rect 1885 160 1925 175
rect 1885 140 1895 160
rect 1915 140 1925 160
rect 1885 125 1925 140
<< ndiffc >>
rect 615 -20 635 0
rect 670 -20 690 0
rect 725 -20 745 0
rect 780 -20 800 0
rect 890 -20 910 0
rect 945 -20 965 0
rect 1000 -20 1020 0
rect 1055 -20 1075 0
rect 1110 -20 1130 0
rect 1220 -20 1240 0
rect 1275 -20 1295 0
rect 1330 -20 1350 0
rect 1385 -20 1405 0
rect 1495 -20 1515 0
rect 1550 -20 1570 0
rect 1605 -20 1625 0
rect 1660 -20 1680 0
rect 1715 -20 1735 0
rect 1785 -20 1805 0
rect 1840 -20 1860 0
<< pdiffc >>
rect 615 140 635 160
rect 670 140 690 160
rect 725 140 745 160
rect 795 140 815 160
rect 850 140 870 160
rect 905 140 925 160
rect 1020 140 1040 160
rect 1075 140 1095 160
rect 1275 140 1295 160
rect 1330 140 1350 160
rect 1385 140 1405 160
rect 1495 140 1515 160
rect 1550 140 1570 160
rect 1605 140 1625 160
rect 1785 140 1805 160
rect 1840 140 1860 160
rect 1895 140 1915 160
<< psubdiff >>
rect 1415 0 1455 15
rect 1415 -20 1425 0
rect 1445 -20 1455 0
rect 1415 -35 1455 -20
<< nsubdiff >>
rect 970 160 1010 175
rect 970 140 980 160
rect 1000 140 1010 160
rect 970 125 1010 140
<< psubdiffcont >>
rect 1425 -20 1445 0
<< nsubdiffcont >>
rect 980 140 1000 160
<< poly >>
rect 1400 225 1440 235
rect 1400 210 1410 225
rect 1360 205 1410 210
rect 1430 205 1440 225
rect 645 185 715 200
rect 1360 195 1440 205
rect 645 175 660 185
rect 700 175 715 185
rect 825 175 840 190
rect 880 175 895 190
rect 1050 175 1065 190
rect 1305 175 1320 190
rect 1360 175 1375 195
rect 1525 175 1540 190
rect 1580 175 1595 190
rect 1815 175 1830 190
rect 1870 175 1885 190
rect 1135 160 1175 170
rect 1135 140 1145 160
rect 1165 145 1175 160
rect 1165 140 1255 145
rect 1135 130 1255 140
rect 645 70 660 125
rect 700 110 715 125
rect 825 115 840 125
rect 740 100 840 115
rect 880 110 895 125
rect 865 100 905 110
rect 1050 105 1065 125
rect 1240 105 1255 130
rect 1305 105 1320 125
rect 740 85 755 100
rect 585 55 660 70
rect 645 15 660 55
rect 700 70 755 85
rect 865 80 875 100
rect 895 80 905 100
rect 865 70 905 80
rect 1030 90 1185 105
rect 1240 90 1320 105
rect 700 15 715 70
rect 780 60 820 70
rect 780 40 790 60
rect 810 40 820 60
rect 1030 40 1045 90
rect 755 25 1045 40
rect 1070 60 1110 65
rect 1070 40 1080 60
rect 1100 40 1110 60
rect 1070 30 1110 40
rect 1170 45 1185 90
rect 1235 60 1275 65
rect 1235 45 1245 60
rect 1170 40 1245 45
rect 1265 40 1275 60
rect 1170 30 1275 40
rect 755 15 770 25
rect 920 15 935 25
rect 975 15 990 25
rect 1030 15 1045 25
rect 1085 15 1100 30
rect 1250 15 1265 30
rect 1305 15 1320 90
rect 1360 15 1375 125
rect 1430 120 1470 130
rect 1430 100 1440 120
rect 1460 110 1470 120
rect 1525 110 1540 125
rect 1460 100 1540 110
rect 1430 95 1540 100
rect 1430 90 1470 95
rect 1415 60 1455 65
rect 1415 40 1425 60
rect 1445 45 1455 60
rect 1580 45 1595 125
rect 1815 115 1830 125
rect 1870 115 1885 125
rect 1630 100 1670 110
rect 1630 80 1640 100
rect 1660 85 1670 100
rect 1815 100 1885 115
rect 1730 85 1770 95
rect 1660 80 1705 85
rect 1630 70 1705 80
rect 1445 40 1650 45
rect 1415 30 1650 40
rect 1525 15 1540 30
rect 1580 15 1595 30
rect 1635 15 1650 30
rect 1690 15 1705 70
rect 1730 65 1740 85
rect 1760 80 1770 85
rect 1815 80 1830 100
rect 1760 65 1830 80
rect 1730 55 1770 65
rect 1815 15 1830 65
rect 1860 65 1900 75
rect 1860 45 1870 65
rect 1890 45 1900 65
rect 1860 35 1900 45
rect 645 -50 660 -35
rect 700 -75 715 -35
rect 755 -50 770 -35
rect 920 -50 935 -35
rect 975 -50 990 -35
rect 1030 -50 1045 -35
rect 1085 -50 1100 -35
rect 1250 -50 1265 -35
rect 1305 -50 1320 -35
rect 1360 -50 1375 -35
rect 1525 -50 1540 -35
rect 1580 -50 1595 -35
rect 1635 -50 1650 -35
rect 1690 -50 1705 -35
rect 1815 -50 1830 -35
rect 1885 -75 1900 35
rect 700 -90 1900 -75
<< polycont >>
rect 1410 205 1430 225
rect 1145 140 1165 160
rect 875 80 895 100
rect 790 40 810 60
rect 1080 40 1100 60
rect 1245 40 1265 60
rect 1440 100 1460 120
rect 1425 40 1445 60
rect 1640 80 1660 100
rect 1740 65 1760 85
rect 1870 45 1890 65
<< locali >>
rect 1400 225 1440 235
rect 1400 205 1410 225
rect 1430 215 1440 225
rect 1430 205 1625 215
rect 1400 195 1625 205
rect 1605 170 1625 195
rect 610 160 640 170
rect 610 140 615 160
rect 635 140 640 160
rect 610 130 640 140
rect 665 160 695 170
rect 665 140 670 160
rect 690 140 695 160
rect 665 130 695 140
rect 720 160 750 170
rect 720 140 725 160
rect 745 140 750 160
rect 720 130 750 140
rect 790 160 820 170
rect 790 140 795 160
rect 815 140 820 160
rect 790 130 820 140
rect 845 160 875 170
rect 845 140 850 160
rect 870 140 875 160
rect 845 130 875 140
rect 900 160 945 170
rect 900 140 905 160
rect 925 140 945 160
rect 900 130 945 140
rect 975 160 1045 170
rect 975 140 980 160
rect 1000 140 1020 160
rect 1040 140 1045 160
rect 975 130 1045 140
rect 1070 160 1100 170
rect 1135 160 1175 170
rect 1270 160 1300 170
rect 1070 140 1075 160
rect 1095 140 1145 160
rect 1165 140 1175 160
rect 1070 130 1100 140
rect 1135 130 1175 140
rect 1195 140 1275 160
rect 1295 140 1300 160
rect 615 50 635 130
rect 725 50 745 130
rect 795 110 815 130
rect 795 100 905 110
rect 795 90 875 100
rect 845 80 875 90
rect 895 80 905 100
rect 845 70 905 80
rect 780 60 820 70
rect 780 50 790 60
rect 615 40 790 50
rect 810 40 820 60
rect 615 30 820 40
rect 615 10 635 30
rect 845 10 865 70
rect 925 50 945 130
rect 1070 60 1110 65
rect 1070 50 1080 60
rect 890 40 1080 50
rect 1100 40 1110 60
rect 890 30 1110 40
rect 890 10 910 30
rect 1000 10 1020 30
rect 1135 10 1155 130
rect 610 0 640 10
rect 610 -20 615 0
rect 635 -20 640 0
rect 610 -30 640 -20
rect 665 0 695 10
rect 665 -20 670 0
rect 690 -20 695 0
rect 665 -30 695 -20
rect 720 0 750 10
rect 720 -20 725 0
rect 745 -20 750 0
rect 720 -30 750 -20
rect 775 0 865 10
rect 775 -20 780 0
rect 800 -10 865 0
rect 885 0 915 10
rect 800 -20 805 -10
rect 775 -30 805 -20
rect 885 -20 890 0
rect 910 -20 915 0
rect 885 -30 915 -20
rect 940 0 970 10
rect 940 -20 945 0
rect 965 -20 970 0
rect 940 -30 970 -20
rect 995 0 1025 10
rect 995 -20 1000 0
rect 1020 -20 1025 0
rect 995 -30 1025 -20
rect 1050 0 1080 10
rect 1050 -20 1055 0
rect 1075 -20 1080 0
rect 1050 -30 1080 -20
rect 1105 0 1155 10
rect 1105 -20 1110 0
rect 1130 -20 1155 0
rect 1195 10 1215 140
rect 1270 130 1300 140
rect 1325 160 1355 170
rect 1325 140 1330 160
rect 1350 140 1355 160
rect 1325 130 1355 140
rect 1380 160 1410 170
rect 1380 140 1385 160
rect 1405 140 1410 160
rect 1380 130 1410 140
rect 1490 160 1520 170
rect 1490 140 1495 160
rect 1515 140 1520 160
rect 1490 130 1520 140
rect 1545 160 1575 170
rect 1545 140 1550 160
rect 1570 140 1575 160
rect 1545 130 1575 140
rect 1600 160 1630 170
rect 1780 160 1810 170
rect 1600 140 1605 160
rect 1625 140 1740 160
rect 1600 130 1630 140
rect 1275 110 1295 130
rect 1385 110 1405 130
rect 1430 120 1470 130
rect 1430 110 1440 120
rect 1275 100 1440 110
rect 1460 100 1470 120
rect 1275 90 1470 100
rect 1235 60 1275 65
rect 1415 60 1455 65
rect 1235 40 1245 60
rect 1265 40 1425 60
rect 1445 40 1455 60
rect 1235 30 1275 40
rect 1415 30 1455 40
rect 1500 50 1520 130
rect 1630 100 1670 110
rect 1630 80 1640 100
rect 1660 80 1670 100
rect 1630 70 1670 80
rect 1720 95 1740 140
rect 1780 140 1785 160
rect 1805 140 1810 160
rect 1780 130 1810 140
rect 1835 160 1865 170
rect 1835 140 1840 160
rect 1860 140 1865 160
rect 1835 130 1865 140
rect 1890 160 1920 170
rect 1890 140 1895 160
rect 1915 140 1920 160
rect 1890 130 1920 140
rect 1720 85 1770 95
rect 1630 50 1650 70
rect 1500 30 1650 50
rect 1720 65 1740 85
rect 1760 65 1770 85
rect 1720 55 1770 65
rect 1840 75 1860 130
rect 1840 70 1900 75
rect 1840 65 1945 70
rect 1500 10 1520 30
rect 1610 10 1630 30
rect 1720 10 1740 55
rect 1840 45 1870 65
rect 1890 50 1945 65
rect 1890 45 1900 50
rect 1840 35 1900 45
rect 1840 10 1860 35
rect 1195 0 1245 10
rect 1195 -20 1220 0
rect 1240 -20 1245 0
rect 1105 -30 1135 -20
rect 1215 -30 1245 -20
rect 1270 0 1300 10
rect 1270 -20 1275 0
rect 1295 -20 1300 0
rect 1270 -30 1300 -20
rect 1325 0 1355 10
rect 1325 -20 1330 0
rect 1350 -20 1355 0
rect 1325 -30 1355 -20
rect 1380 0 1450 10
rect 1380 -20 1385 0
rect 1405 -20 1425 0
rect 1445 -20 1450 0
rect 1380 -30 1450 -20
rect 1490 0 1520 10
rect 1490 -20 1495 0
rect 1515 -20 1520 0
rect 1490 -30 1520 -20
rect 1545 0 1575 10
rect 1545 -20 1550 0
rect 1570 -20 1575 0
rect 1545 -30 1575 -20
rect 1600 0 1630 10
rect 1600 -20 1605 0
rect 1625 -20 1630 0
rect 1600 -30 1630 -20
rect 1655 0 1685 10
rect 1655 -20 1660 0
rect 1680 -20 1685 0
rect 1655 -30 1685 -20
rect 1710 0 1740 10
rect 1710 -20 1715 0
rect 1735 -20 1740 0
rect 1710 -30 1740 -20
rect 1780 0 1810 10
rect 1780 -20 1785 0
rect 1805 -20 1810 0
rect 1780 -30 1810 -20
rect 1835 0 1865 10
rect 1835 -20 1840 0
rect 1860 -20 1865 0
rect 1835 -30 1865 -20
<< viali >>
rect 670 140 690 160
rect 850 140 870 160
rect 980 140 1000 160
rect 1020 140 1040 160
rect 670 -20 690 0
rect 945 -20 965 0
rect 1055 -20 1075 0
rect 1330 140 1350 160
rect 1550 140 1570 160
rect 1785 140 1805 160
rect 1895 140 1915 160
rect 1385 -20 1405 0
rect 1425 -20 1445 0
rect 1550 -20 1570 0
rect 1660 -20 1680 0
rect 1785 -20 1805 0
<< metal1 >>
rect 585 160 1945 175
rect 585 140 670 160
rect 690 140 850 160
rect 870 140 980 160
rect 1000 140 1020 160
rect 1040 140 1330 160
rect 1350 140 1550 160
rect 1570 140 1785 160
rect 1805 140 1895 160
rect 1915 140 1945 160
rect 585 125 1945 140
rect 585 0 1945 15
rect 585 -20 670 0
rect 690 -20 945 0
rect 965 -20 1055 0
rect 1075 -20 1385 0
rect 1405 -20 1425 0
rect 1445 -20 1550 0
rect 1570 -20 1660 0
rect 1680 -20 1785 0
rect 1805 -20 1945 0
rect 585 -35 1945 -20
<< labels >>
flabel metal1 585 150 585 150 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel metal1 585 -10 585 -10 7 FreeSans 160 0 -80 0 GNDA
port 4 w
flabel poly 585 60 585 60 7 FreeSans 160 0 -80 0 VIN
port 2 w
flabel locali 680 50 680 50 1 FreeSans 160 0 0 80 CLK
flabel locali 795 90 795 90 7 FreeSans 160 0 -80 0 A
flabel locali 735 -30 735 -30 5 FreeSans 160 0 0 -80 B
flabel locali 945 80 945 80 3 FreeSans 160 0 80 0 C
flabel locali 1155 45 1155 45 3 FreeSans 160 0 0 0 D
flabel locali 1740 160 1740 160 3 FreeSans 160 0 80 0 I
flabel locali 1195 160 1195 160 7 FreeSans 160 0 -80 0 E
flabel locali 1285 -30 1285 -30 5 FreeSans 160 0 0 -80 F
flabel locali 1340 -30 1340 -30 5 FreeSans 160 0 0 -80 G
flabel locali 1520 70 1520 70 3 FreeSans 160 0 80 0 H
flabel locali 1945 60 1945 60 3 FreeSans 160 0 80 0 VOUT
<< end >>
