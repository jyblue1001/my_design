magic
tech sky130A
timestamp 1738175887
<< nwell >>
rect -170 190 295 430
rect 445 330 885 430
rect 445 190 955 330
rect 820 185 955 190
rect 860 165 955 185
<< nmos >>
rect 0 0 15 100
rect 700 0 715 100
<< pmos >>
rect 0 210 15 410
rect 700 210 715 410
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 650 85 700 100
rect 650 15 665 85
rect 685 15 700 85
rect 650 0 700 15
rect 715 85 765 100
rect 715 15 730 85
rect 750 15 765 85
rect 715 0 765 15
<< pdiff >>
rect -50 395 0 410
rect -50 225 -35 395
rect -15 225 0 395
rect -50 210 0 225
rect 15 395 65 410
rect 15 225 30 395
rect 50 225 65 395
rect 15 210 65 225
rect 650 395 700 410
rect 650 225 665 395
rect 685 225 700 395
rect 650 210 700 225
rect 715 395 765 410
rect 715 225 730 395
rect 750 225 765 395
rect 715 210 765 225
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 665 15 685 85
rect 730 15 750 85
<< pdiffc >>
rect -35 225 -15 395
rect 30 225 50 395
rect 665 225 685 395
rect 730 225 750 395
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 395 -50 410
rect -100 225 -85 395
rect -65 225 -50 395
rect -100 210 -50 225
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 225 -65 395
<< poly >>
rect 0 410 15 475
rect 585 440 625 450
rect 585 420 595 440
rect 615 420 625 440
rect 585 410 625 420
rect 700 410 715 425
rect 0 165 15 210
rect -185 150 15 165
rect 0 100 15 150
rect 600 125 615 410
rect 700 200 715 210
rect 700 185 835 200
rect 600 110 715 125
rect 700 100 715 110
rect 820 10 835 185
rect 805 0 845 10
rect 0 -65 15 0
rect 700 -15 715 0
rect 805 -20 815 0
rect 835 -20 845 0
rect 805 -30 845 -20
<< polycont >>
rect 595 420 615 440
rect 815 -20 835 0
<< locali >>
rect -175 500 935 510
rect -175 480 -85 500
rect -65 480 -40 500
rect -20 480 5 500
rect 25 480 50 500
rect 70 480 95 500
rect 115 480 140 500
rect 160 480 185 500
rect 205 480 230 500
rect 250 480 275 500
rect 295 480 320 500
rect 340 480 365 500
rect 385 480 410 500
rect 430 480 455 500
rect 475 480 500 500
rect 520 480 545 500
rect 565 480 620 500
rect 640 480 820 500
rect 840 480 865 500
rect 885 480 910 500
rect 930 480 935 500
rect -175 470 935 480
rect -85 405 -65 470
rect -40 405 -20 470
rect 595 450 615 470
rect 585 440 625 450
rect 585 420 595 440
rect 615 420 625 440
rect 585 410 625 420
rect -95 395 -5 405
rect -95 225 -85 395
rect -65 225 -35 395
rect -15 225 -5 395
rect -95 215 -5 225
rect 20 395 65 405
rect 20 225 30 395
rect 50 225 65 395
rect 20 215 65 225
rect 655 395 695 405
rect 655 225 665 395
rect 685 225 695 395
rect 655 215 695 225
rect 720 395 765 405
rect 720 225 730 395
rect 750 225 765 395
rect 720 215 765 225
rect 30 165 50 215
rect 665 195 685 215
rect 555 175 685 195
rect 30 145 145 165
rect 30 95 50 145
rect 665 95 685 175
rect 730 135 750 215
rect 730 115 880 135
rect 730 95 750 115
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 650 85 695 95
rect 650 15 665 85
rect 685 15 695 85
rect 650 5 695 15
rect 720 85 760 95
rect 720 15 730 85
rect 750 15 760 85
rect 720 5 760 15
rect -85 -50 -65 5
rect -40 -50 -20 5
rect 805 0 845 10
rect 805 -20 815 0
rect 835 -20 845 0
rect 805 -30 845 -20
rect 815 -50 835 -30
rect -180 -70 885 -50
rect -180 -90 -85 -70
rect -65 -90 -40 -70
rect -20 -90 5 -70
rect 25 -90 50 -70
rect 70 -90 95 -70
rect 115 -90 140 -70
rect 160 -90 185 -70
rect 205 -90 230 -70
rect 250 -90 275 -70
rect 295 -90 320 -70
rect 340 -90 365 -70
rect 385 -90 410 -70
rect 430 -90 455 -70
rect 475 -90 500 -70
rect 520 -90 540 -70
rect 560 -90 585 -70
rect 605 -90 770 -70
rect 790 -90 815 -70
rect 835 -90 860 -70
rect 880 -90 885 -70
rect -180 -110 885 -90
<< viali >>
rect -85 480 -65 500
rect -40 480 -20 500
rect 5 480 25 500
rect 50 480 70 500
rect 95 480 115 500
rect 140 480 160 500
rect 185 480 205 500
rect 230 480 250 500
rect 275 480 295 500
rect 320 480 340 500
rect 365 480 385 500
rect 410 480 430 500
rect 455 480 475 500
rect 500 480 520 500
rect 545 480 565 500
rect 620 480 640 500
rect 820 480 840 500
rect 865 480 885 500
rect 910 480 930 500
rect -85 -90 -65 -70
rect -40 -90 -20 -70
rect 5 -90 25 -70
rect 50 -90 70 -70
rect 95 -90 115 -70
rect 140 -90 160 -70
rect 185 -90 205 -70
rect 230 -90 250 -70
rect 275 -90 295 -70
rect 320 -90 340 -70
rect 365 -90 385 -70
rect 410 -90 430 -70
rect 455 -90 475 -70
rect 500 -90 520 -70
rect 540 -90 560 -70
rect 585 -90 605 -70
rect 770 -90 790 -70
rect 815 -90 835 -70
rect 860 -90 880 -70
<< metal1 >>
rect -175 500 935 520
rect -175 480 -85 500
rect -65 480 -40 500
rect -20 480 5 500
rect 25 480 50 500
rect 70 480 95 500
rect 115 480 140 500
rect 160 480 185 500
rect 205 480 230 500
rect 250 480 275 500
rect 295 480 320 500
rect 340 480 365 500
rect 385 480 410 500
rect 430 480 455 500
rect 475 480 500 500
rect 520 480 545 500
rect 565 480 620 500
rect 640 480 820 500
rect 840 480 865 500
rect 885 480 910 500
rect 930 480 935 500
rect -175 470 935 480
rect -175 460 830 470
rect 850 460 935 470
rect -180 -70 885 -40
rect -180 -90 -85 -70
rect -65 -90 -40 -70
rect -20 -90 5 -70
rect 25 -90 50 -70
rect 70 -90 95 -70
rect 115 -90 140 -70
rect 160 -90 185 -70
rect 205 -90 230 -70
rect 250 -90 275 -70
rect 295 -90 320 -70
rect 340 -90 365 -70
rect 385 -90 410 -70
rect 430 -90 455 -70
rect 475 -90 500 -70
rect 520 -90 540 -70
rect 560 -90 585 -70
rect 605 -90 770 -70
rect 790 -90 815 -70
rect 835 -90 860 -70
rect 880 -90 885 -70
rect -180 -120 885 -90
<< labels >>
flabel locali 880 125 880 125 3 FreeSans 400 0 80 0 D
flabel locali 145 155 145 155 3 FreeSans 400 0 80 0 B
flabel poly -185 155 -185 155 7 FreeSans 400 0 -80 0 A
flabel metal1 -180 -80 -180 -80 7 FreeSans 400 0 -80 0 GNDA
flabel metal1 -175 490 -175 490 7 FreeSans 400 0 -80 0 VDDA
flabel locali 555 185 555 185 7 FreeSans 400 0 -200 0 C
<< end >>
