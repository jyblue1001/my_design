magic
tech sky130A
timestamp 1740284794
<< nwell >>
rect 1175 -5 2315 580
<< nmos >>
rect 1640 -90 1655 -40
rect 1940 -90 1955 -40
rect 2240 -90 2255 -40
rect 1640 -210 1655 -160
rect 1940 -210 1955 -160
rect 2240 -210 2255 -160
rect 1505 -375 1520 -275
rect 1640 -375 1655 -275
rect 1940 -375 1955 -275
rect 2240 -375 2255 -275
<< pmos >>
rect 1235 360 1385 560
rect 1505 360 1655 560
rect 1805 360 1955 560
rect 2105 360 2255 560
rect 1640 185 1655 285
rect 1940 185 1955 285
rect 2240 185 2255 285
rect 1640 15 1655 115
rect 1940 15 1955 115
rect 2240 15 2255 115
<< ndiff >>
rect 1600 -55 1640 -40
rect 1600 -75 1610 -55
rect 1630 -75 1640 -55
rect 1600 -90 1640 -75
rect 1655 -55 1695 -40
rect 1655 -75 1665 -55
rect 1685 -75 1695 -55
rect 1655 -90 1695 -75
rect 1900 -55 1940 -40
rect 1900 -75 1910 -55
rect 1930 -75 1940 -55
rect 1900 -90 1940 -75
rect 1955 -55 1995 -40
rect 1955 -75 1965 -55
rect 1985 -75 1995 -55
rect 1955 -90 1995 -75
rect 2200 -55 2240 -40
rect 2200 -75 2210 -55
rect 2230 -75 2240 -55
rect 2200 -90 2240 -75
rect 2255 -55 2295 -40
rect 2255 -75 2265 -55
rect 2285 -75 2295 -55
rect 2255 -90 2295 -75
rect 1600 -175 1640 -160
rect 1600 -195 1610 -175
rect 1630 -195 1640 -175
rect 1600 -210 1640 -195
rect 1655 -175 1695 -160
rect 1655 -195 1665 -175
rect 1685 -195 1695 -175
rect 1655 -210 1695 -195
rect 1900 -175 1940 -160
rect 1900 -195 1910 -175
rect 1930 -195 1940 -175
rect 1900 -210 1940 -195
rect 1955 -175 1995 -160
rect 1955 -195 1965 -175
rect 1985 -195 1995 -175
rect 1955 -210 1995 -195
rect 2200 -175 2240 -160
rect 2200 -195 2210 -175
rect 2230 -195 2240 -175
rect 2200 -210 2240 -195
rect 2255 -175 2295 -160
rect 2255 -195 2265 -175
rect 2285 -195 2295 -175
rect 2255 -210 2295 -195
rect 1465 -290 1505 -275
rect 1465 -310 1475 -290
rect 1495 -310 1505 -290
rect 1465 -340 1505 -310
rect 1465 -360 1475 -340
rect 1495 -360 1505 -340
rect 1465 -375 1505 -360
rect 1520 -290 1560 -275
rect 1600 -290 1640 -275
rect 1520 -310 1530 -290
rect 1550 -310 1560 -290
rect 1600 -310 1610 -290
rect 1630 -310 1640 -290
rect 1520 -340 1560 -310
rect 1600 -340 1640 -310
rect 1520 -360 1530 -340
rect 1550 -360 1560 -340
rect 1600 -360 1610 -340
rect 1630 -360 1640 -340
rect 1520 -375 1560 -360
rect 1600 -375 1640 -360
rect 1655 -290 1695 -275
rect 1655 -310 1665 -290
rect 1685 -310 1695 -290
rect 1655 -340 1695 -310
rect 1655 -360 1665 -340
rect 1685 -360 1695 -340
rect 1655 -375 1695 -360
rect 1900 -290 1940 -275
rect 1900 -310 1910 -290
rect 1930 -310 1940 -290
rect 1900 -340 1940 -310
rect 1900 -360 1910 -340
rect 1930 -360 1940 -340
rect 1900 -375 1940 -360
rect 1955 -290 1995 -275
rect 1955 -310 1965 -290
rect 1985 -310 1995 -290
rect 1955 -340 1995 -310
rect 1955 -360 1965 -340
rect 1985 -360 1995 -340
rect 1955 -375 1995 -360
rect 2200 -290 2240 -275
rect 2200 -310 2210 -290
rect 2230 -310 2240 -290
rect 2200 -340 2240 -310
rect 2200 -360 2210 -340
rect 2230 -360 2240 -340
rect 2200 -375 2240 -360
rect 2255 -290 2295 -275
rect 2255 -310 2265 -290
rect 2285 -310 2295 -290
rect 2255 -340 2295 -310
rect 2255 -360 2265 -340
rect 2285 -360 2295 -340
rect 2255 -375 2295 -360
<< pdiff >>
rect 1195 545 1235 560
rect 1195 525 1205 545
rect 1225 525 1235 545
rect 1195 495 1235 525
rect 1195 475 1205 495
rect 1225 475 1235 495
rect 1195 445 1235 475
rect 1195 425 1205 445
rect 1225 425 1235 445
rect 1195 395 1235 425
rect 1195 375 1205 395
rect 1225 375 1235 395
rect 1195 360 1235 375
rect 1385 545 1425 560
rect 1465 545 1505 560
rect 1385 525 1395 545
rect 1415 525 1425 545
rect 1465 525 1475 545
rect 1495 525 1505 545
rect 1385 495 1425 525
rect 1465 495 1505 525
rect 1385 475 1395 495
rect 1415 475 1425 495
rect 1465 475 1475 495
rect 1495 475 1505 495
rect 1385 445 1425 475
rect 1465 445 1505 475
rect 1385 425 1395 445
rect 1415 425 1425 445
rect 1465 425 1475 445
rect 1495 425 1505 445
rect 1385 395 1425 425
rect 1465 395 1505 425
rect 1385 375 1395 395
rect 1415 375 1425 395
rect 1465 375 1475 395
rect 1495 375 1505 395
rect 1385 360 1425 375
rect 1465 360 1505 375
rect 1655 545 1695 560
rect 1655 525 1665 545
rect 1685 525 1695 545
rect 1655 495 1695 525
rect 1655 475 1665 495
rect 1685 475 1695 495
rect 1655 445 1695 475
rect 1655 425 1665 445
rect 1685 425 1695 445
rect 1655 395 1695 425
rect 1655 375 1665 395
rect 1685 375 1695 395
rect 1655 360 1695 375
rect 1765 545 1805 560
rect 1765 525 1775 545
rect 1795 525 1805 545
rect 1765 495 1805 525
rect 1765 475 1775 495
rect 1795 475 1805 495
rect 1765 445 1805 475
rect 1765 425 1775 445
rect 1795 425 1805 445
rect 1765 395 1805 425
rect 1765 375 1775 395
rect 1795 375 1805 395
rect 1765 360 1805 375
rect 1955 545 1995 560
rect 1955 525 1965 545
rect 1985 525 1995 545
rect 1955 495 1995 525
rect 1955 475 1965 495
rect 1985 475 1995 495
rect 1955 445 1995 475
rect 1955 425 1965 445
rect 1985 425 1995 445
rect 1955 395 1995 425
rect 1955 375 1965 395
rect 1985 375 1995 395
rect 1955 360 1995 375
rect 2065 545 2105 560
rect 2065 525 2075 545
rect 2095 525 2105 545
rect 2065 495 2105 525
rect 2065 475 2075 495
rect 2095 475 2105 495
rect 2065 445 2105 475
rect 2065 425 2075 445
rect 2095 425 2105 445
rect 2065 395 2105 425
rect 2065 375 2075 395
rect 2095 375 2105 395
rect 2065 360 2105 375
rect 2255 545 2295 560
rect 2255 525 2265 545
rect 2285 525 2295 545
rect 2255 495 2295 525
rect 2255 475 2265 495
rect 2285 475 2295 495
rect 2255 445 2295 475
rect 2255 425 2265 445
rect 2285 425 2295 445
rect 2255 395 2295 425
rect 2255 375 2265 395
rect 2285 375 2295 395
rect 2255 360 2295 375
rect 1600 270 1640 285
rect 1600 250 1610 270
rect 1630 250 1640 270
rect 1600 220 1640 250
rect 1600 200 1610 220
rect 1630 200 1640 220
rect 1600 185 1640 200
rect 1655 270 1695 285
rect 1655 250 1665 270
rect 1685 250 1695 270
rect 1655 220 1695 250
rect 1655 200 1665 220
rect 1685 200 1695 220
rect 1655 185 1695 200
rect 1900 270 1940 285
rect 1900 250 1910 270
rect 1930 250 1940 270
rect 1900 220 1940 250
rect 1900 200 1910 220
rect 1930 200 1940 220
rect 1900 185 1940 200
rect 1955 270 1995 285
rect 1955 250 1965 270
rect 1985 250 1995 270
rect 1955 220 1995 250
rect 1955 200 1965 220
rect 1985 200 1995 220
rect 1955 185 1995 200
rect 2200 270 2240 285
rect 2200 250 2210 270
rect 2230 250 2240 270
rect 2200 220 2240 250
rect 2200 200 2210 220
rect 2230 200 2240 220
rect 2200 185 2240 200
rect 2255 270 2295 285
rect 2255 250 2265 270
rect 2285 250 2295 270
rect 2255 220 2295 250
rect 2255 200 2265 220
rect 2285 200 2295 220
rect 2255 185 2295 200
rect 1600 100 1640 115
rect 1600 80 1610 100
rect 1630 80 1640 100
rect 1600 50 1640 80
rect 1600 30 1610 50
rect 1630 30 1640 50
rect 1600 15 1640 30
rect 1655 100 1695 115
rect 1655 80 1665 100
rect 1685 80 1695 100
rect 1655 50 1695 80
rect 1655 30 1665 50
rect 1685 30 1695 50
rect 1655 15 1695 30
rect 1900 100 1940 115
rect 1900 80 1910 100
rect 1930 80 1940 100
rect 1900 50 1940 80
rect 1900 30 1910 50
rect 1930 30 1940 50
rect 1900 15 1940 30
rect 1955 100 1995 115
rect 1955 80 1965 100
rect 1985 80 1995 100
rect 1955 50 1995 80
rect 1955 30 1965 50
rect 1985 30 1995 50
rect 1955 15 1995 30
rect 2200 100 2240 115
rect 2200 80 2210 100
rect 2230 80 2240 100
rect 2200 50 2240 80
rect 2200 30 2210 50
rect 2230 30 2240 50
rect 2200 15 2240 30
rect 2255 100 2295 115
rect 2255 80 2265 100
rect 2285 80 2295 100
rect 2255 50 2295 80
rect 2255 30 2265 50
rect 2285 30 2295 50
rect 2255 15 2295 30
<< ndiffc >>
rect 1610 -75 1630 -55
rect 1665 -75 1685 -55
rect 1910 -75 1930 -55
rect 1965 -75 1985 -55
rect 2210 -75 2230 -55
rect 2265 -75 2285 -55
rect 1610 -195 1630 -175
rect 1665 -195 1685 -175
rect 1910 -195 1930 -175
rect 1965 -195 1985 -175
rect 2210 -195 2230 -175
rect 2265 -195 2285 -175
rect 1475 -310 1495 -290
rect 1475 -360 1495 -340
rect 1530 -310 1550 -290
rect 1610 -310 1630 -290
rect 1530 -360 1550 -340
rect 1610 -360 1630 -340
rect 1665 -310 1685 -290
rect 1665 -360 1685 -340
rect 1910 -310 1930 -290
rect 1910 -360 1930 -340
rect 1965 -310 1985 -290
rect 1965 -360 1985 -340
rect 2210 -310 2230 -290
rect 2210 -360 2230 -340
rect 2265 -310 2285 -290
rect 2265 -360 2285 -340
<< pdiffc >>
rect 1205 525 1225 545
rect 1205 475 1225 495
rect 1205 425 1225 445
rect 1205 375 1225 395
rect 1395 525 1415 545
rect 1475 525 1495 545
rect 1395 475 1415 495
rect 1475 475 1495 495
rect 1395 425 1415 445
rect 1475 425 1495 445
rect 1395 375 1415 395
rect 1475 375 1495 395
rect 1665 525 1685 545
rect 1665 475 1685 495
rect 1665 425 1685 445
rect 1665 375 1685 395
rect 1775 525 1795 545
rect 1775 475 1795 495
rect 1775 425 1795 445
rect 1775 375 1795 395
rect 1965 525 1985 545
rect 1965 475 1985 495
rect 1965 425 1985 445
rect 1965 375 1985 395
rect 2075 525 2095 545
rect 2075 475 2095 495
rect 2075 425 2095 445
rect 2075 375 2095 395
rect 2265 525 2285 545
rect 2265 475 2285 495
rect 2265 425 2285 445
rect 2265 375 2285 395
rect 1610 250 1630 270
rect 1610 200 1630 220
rect 1665 250 1685 270
rect 1665 200 1685 220
rect 1910 250 1930 270
rect 1910 200 1930 220
rect 1965 250 1985 270
rect 1965 200 1985 220
rect 2210 250 2230 270
rect 2210 200 2230 220
rect 2265 250 2285 270
rect 2265 200 2285 220
rect 1610 80 1630 100
rect 1610 30 1630 50
rect 1665 80 1685 100
rect 1665 30 1685 50
rect 1910 80 1930 100
rect 1910 30 1930 50
rect 1965 80 1985 100
rect 1965 30 1985 50
rect 2210 80 2230 100
rect 2210 30 2230 50
rect 2265 80 2285 100
rect 2265 30 2285 50
<< psubdiff >>
rect 1560 -175 1600 -160
rect 1560 -195 1570 -175
rect 1590 -195 1600 -175
rect 1560 -210 1600 -195
rect 1860 -175 1900 -160
rect 1860 -195 1870 -175
rect 1890 -195 1900 -175
rect 1860 -210 1900 -195
rect 2160 -175 2200 -160
rect 2160 -195 2170 -175
rect 2190 -195 2200 -175
rect 2160 -210 2200 -195
rect 1560 -290 1600 -275
rect 1560 -310 1570 -290
rect 1590 -310 1600 -290
rect 1560 -340 1600 -310
rect 1560 -360 1570 -340
rect 1590 -360 1600 -340
rect 1560 -375 1600 -360
rect 1860 -290 1900 -275
rect 1860 -310 1870 -290
rect 1890 -310 1900 -290
rect 1860 -340 1900 -310
rect 1860 -360 1870 -340
rect 1890 -360 1900 -340
rect 1860 -375 1900 -360
rect 2160 -290 2200 -275
rect 2160 -310 2170 -290
rect 2190 -310 2200 -290
rect 2160 -340 2200 -310
rect 2160 -360 2170 -340
rect 2190 -360 2200 -340
rect 2160 -375 2200 -360
<< nsubdiff >>
rect 1425 545 1465 560
rect 1425 525 1435 545
rect 1455 525 1465 545
rect 1425 495 1465 525
rect 1425 475 1435 495
rect 1455 475 1465 495
rect 1425 445 1465 475
rect 1425 425 1435 445
rect 1455 425 1465 445
rect 1425 395 1465 425
rect 1425 375 1435 395
rect 1455 375 1465 395
rect 1425 360 1465 375
rect 1725 545 1765 560
rect 1725 525 1735 545
rect 1755 525 1765 545
rect 1725 495 1765 525
rect 1725 475 1735 495
rect 1755 475 1765 495
rect 1725 445 1765 475
rect 1725 425 1735 445
rect 1755 425 1765 445
rect 1725 395 1765 425
rect 1725 375 1735 395
rect 1755 375 1765 395
rect 1725 360 1765 375
rect 2025 545 2065 560
rect 2025 525 2035 545
rect 2055 525 2065 545
rect 2025 495 2065 525
rect 2025 475 2035 495
rect 2055 475 2065 495
rect 2025 445 2065 475
rect 2025 425 2035 445
rect 2055 425 2065 445
rect 2025 395 2065 425
rect 2025 375 2035 395
rect 2055 375 2065 395
rect 2025 360 2065 375
rect 1560 270 1600 285
rect 1560 250 1570 270
rect 1590 250 1600 270
rect 1560 220 1600 250
rect 1560 200 1570 220
rect 1590 200 1600 220
rect 1560 185 1600 200
rect 1860 270 1900 285
rect 1860 250 1870 270
rect 1890 250 1900 270
rect 1860 220 1900 250
rect 1860 200 1870 220
rect 1890 200 1900 220
rect 1860 185 1900 200
rect 2160 270 2200 285
rect 2160 250 2170 270
rect 2190 250 2200 270
rect 2160 220 2200 250
rect 2160 200 2170 220
rect 2190 200 2200 220
rect 2160 185 2200 200
<< psubdiffcont >>
rect 1570 -195 1590 -175
rect 1870 -195 1890 -175
rect 2170 -195 2190 -175
rect 1570 -310 1590 -290
rect 1570 -360 1590 -340
rect 1870 -310 1890 -290
rect 1870 -360 1890 -340
rect 2170 -310 2190 -290
rect 2170 -360 2190 -340
<< nsubdiffcont >>
rect 1435 525 1455 545
rect 1435 475 1455 495
rect 1435 425 1455 445
rect 1435 375 1455 395
rect 1735 525 1755 545
rect 1735 475 1755 495
rect 1735 425 1755 445
rect 1735 375 1755 395
rect 2035 525 2055 545
rect 2035 475 2055 495
rect 2035 425 2055 445
rect 2035 375 2055 395
rect 1570 250 1590 270
rect 1570 200 1590 220
rect 1870 250 1890 270
rect 1870 200 1890 220
rect 2170 250 2190 270
rect 2170 200 2190 220
<< poly >>
rect 1235 560 1385 575
rect 1505 560 1655 575
rect 1805 560 1955 575
rect 2105 560 2255 575
rect 1235 345 1385 360
rect 1505 345 1655 360
rect 1805 345 1955 360
rect 2105 345 2255 360
rect 1235 335 1265 345
rect 1235 315 1240 335
rect 1260 315 1265 335
rect 1235 305 1265 315
rect 1295 335 1325 345
rect 1295 315 1300 335
rect 1320 315 1325 335
rect 1295 305 1325 315
rect 1355 335 2255 345
rect 1355 315 1360 335
rect 1380 325 2255 335
rect 1380 315 1385 325
rect 1355 305 1385 315
rect 1640 285 1655 300
rect 1940 285 1955 300
rect 2240 285 2255 300
rect 1640 170 1655 185
rect 1940 170 1955 185
rect 2240 170 2255 185
rect 1505 160 1655 170
rect 1505 140 1515 160
rect 1535 155 1655 160
rect 1805 160 1955 170
rect 1535 140 1545 155
rect 1505 130 1545 140
rect 1805 140 1815 160
rect 1835 155 1955 160
rect 2105 160 2255 170
rect 1835 140 1845 155
rect 1805 130 1845 140
rect 2105 140 2115 160
rect 2135 155 2255 160
rect 2135 140 2145 155
rect 2105 130 2145 140
rect 1640 115 1655 130
rect 1940 115 1955 130
rect 2240 115 2255 130
rect 1640 -5 1655 15
rect 1710 0 1750 10
rect 1710 -5 1720 0
rect 1640 -20 1720 -5
rect 1740 -20 1750 0
rect 1640 -40 1655 -20
rect 1710 -30 1750 -20
rect 1940 -5 1955 15
rect 2010 0 2050 10
rect 2010 -5 2020 0
rect 1940 -20 2020 -5
rect 2040 -20 2050 0
rect 1940 -40 1955 -20
rect 2010 -30 2050 -20
rect 2240 -5 2255 15
rect 2310 0 2350 10
rect 2310 -5 2320 0
rect 2240 -20 2320 -5
rect 2340 -20 2350 0
rect 2240 -40 2255 -20
rect 2310 -30 2350 -20
rect 1640 -105 1655 -90
rect 1940 -105 1955 -90
rect 2240 -105 2255 -90
rect 1540 -115 1580 -105
rect 1540 -135 1550 -115
rect 1570 -130 1580 -115
rect 1840 -115 1880 -105
rect 1570 -135 1655 -130
rect 1540 -145 1655 -135
rect 1840 -135 1850 -115
rect 1870 -130 1880 -115
rect 2140 -115 2180 -105
rect 1870 -135 1955 -130
rect 1840 -145 1955 -135
rect 2140 -135 2150 -115
rect 2170 -130 2180 -115
rect 2170 -135 2255 -130
rect 2140 -145 2255 -135
rect 1640 -160 1655 -145
rect 1940 -160 1955 -145
rect 2240 -160 2255 -145
rect 1640 -225 1655 -210
rect 1940 -225 1955 -210
rect 2240 -225 2255 -210
rect 1345 -265 2255 -250
rect 1505 -275 1520 -265
rect 1640 -275 1655 -265
rect 1940 -275 1955 -265
rect 2240 -275 2255 -265
rect 1505 -390 1520 -375
rect 1640 -390 1655 -375
rect 1940 -390 1955 -375
rect 2240 -390 2255 -375
<< polycont >>
rect 1240 315 1260 335
rect 1300 315 1320 335
rect 1360 315 1380 335
rect 1515 140 1535 160
rect 1815 140 1835 160
rect 2115 140 2135 160
rect 1720 -20 1740 0
rect 2020 -20 2040 0
rect 2320 -20 2340 0
rect 1550 -135 1570 -115
rect 1850 -135 1870 -115
rect 2150 -135 2170 -115
<< locali >>
rect 1195 595 1225 615
rect 1245 595 1275 615
rect 1295 595 1325 615
rect 1345 595 1375 615
rect 1395 595 1425 615
rect 1445 595 1475 615
rect 1495 595 1525 615
rect 1545 595 1575 615
rect 1595 595 1625 615
rect 1645 595 1675 615
rect 1695 595 1725 615
rect 1745 595 1775 615
rect 1795 595 1825 615
rect 1845 595 1875 615
rect 1895 595 1925 615
rect 1945 595 1975 615
rect 1995 595 2025 615
rect 2045 595 2075 615
rect 2095 595 2125 615
rect 2145 595 2175 615
rect 2195 595 2225 615
rect 2245 595 2275 615
rect 2295 595 2325 615
rect 2345 595 2350 615
rect 1430 555 1460 595
rect 1770 555 1800 595
rect 2070 555 2100 595
rect 1200 545 1230 555
rect 1200 525 1205 545
rect 1225 525 1230 545
rect 1200 495 1230 525
rect 1200 475 1205 495
rect 1225 475 1230 495
rect 1200 445 1230 475
rect 1200 425 1205 445
rect 1225 425 1230 445
rect 1200 395 1230 425
rect 1200 375 1205 395
rect 1225 375 1230 395
rect 1200 345 1230 375
rect 1390 545 1500 555
rect 1390 525 1395 545
rect 1415 525 1435 545
rect 1455 525 1475 545
rect 1495 525 1500 545
rect 1390 495 1500 525
rect 1390 475 1395 495
rect 1415 475 1435 495
rect 1455 475 1475 495
rect 1495 475 1500 495
rect 1390 445 1500 475
rect 1390 425 1395 445
rect 1415 425 1435 445
rect 1455 425 1475 445
rect 1495 425 1500 445
rect 1390 395 1500 425
rect 1390 375 1395 395
rect 1415 375 1435 395
rect 1455 375 1475 395
rect 1495 375 1500 395
rect 1390 365 1500 375
rect 1660 545 1690 555
rect 1660 525 1665 545
rect 1685 525 1690 545
rect 1660 495 1690 525
rect 1660 475 1665 495
rect 1685 475 1690 495
rect 1660 445 1690 475
rect 1660 425 1665 445
rect 1685 425 1690 445
rect 1660 395 1690 425
rect 1660 375 1665 395
rect 1685 375 1690 395
rect 1200 335 1385 345
rect 1200 315 1240 335
rect 1260 315 1300 335
rect 1320 315 1360 335
rect 1380 315 1385 335
rect 1200 305 1385 315
rect 1365 -280 1385 305
rect 1430 280 1460 365
rect 1430 270 1635 280
rect 1430 250 1570 270
rect 1590 250 1610 270
rect 1630 250 1635 270
rect 1560 220 1635 250
rect 1560 200 1570 220
rect 1590 200 1610 220
rect 1630 200 1635 220
rect 1560 190 1635 200
rect 1660 270 1690 375
rect 1730 545 1800 555
rect 1730 525 1735 545
rect 1755 525 1775 545
rect 1795 525 1800 545
rect 1730 495 1800 525
rect 1730 475 1735 495
rect 1755 475 1775 495
rect 1795 475 1800 495
rect 1730 445 1800 475
rect 1730 425 1735 445
rect 1755 425 1775 445
rect 1795 425 1800 445
rect 1730 395 1800 425
rect 1730 375 1735 395
rect 1755 375 1775 395
rect 1795 375 1800 395
rect 1730 365 1800 375
rect 1660 250 1665 270
rect 1685 250 1690 270
rect 1770 280 1800 365
rect 1960 545 1990 555
rect 1960 525 1965 545
rect 1985 525 1990 545
rect 1960 495 1990 525
rect 1960 475 1965 495
rect 1985 475 1990 495
rect 1960 445 1990 475
rect 1960 425 1965 445
rect 1985 425 1990 445
rect 1960 395 1990 425
rect 1960 375 1965 395
rect 1985 375 1990 395
rect 1770 270 1935 280
rect 1770 250 1870 270
rect 1890 250 1910 270
rect 1930 250 1935 270
rect 1660 220 1690 250
rect 1660 200 1665 220
rect 1685 200 1690 220
rect 1505 160 1545 170
rect 1505 140 1515 160
rect 1535 140 1545 160
rect 1505 130 1545 140
rect 1605 100 1635 110
rect 1605 80 1610 100
rect 1630 80 1635 100
rect 1605 50 1635 80
rect 1605 30 1610 50
rect 1630 30 1635 50
rect 1605 10 1635 30
rect 1660 100 1690 200
rect 1860 220 1935 250
rect 1860 200 1870 220
rect 1890 200 1910 220
rect 1930 200 1935 220
rect 1860 190 1935 200
rect 1960 270 1990 375
rect 2030 545 2100 555
rect 2030 525 2035 545
rect 2055 525 2075 545
rect 2095 525 2100 545
rect 2030 495 2100 525
rect 2030 475 2035 495
rect 2055 475 2075 495
rect 2095 475 2100 495
rect 2030 445 2100 475
rect 2030 425 2035 445
rect 2055 425 2075 445
rect 2095 425 2100 445
rect 2030 395 2100 425
rect 2030 375 2035 395
rect 2055 375 2075 395
rect 2095 375 2100 395
rect 2030 365 2100 375
rect 1960 250 1965 270
rect 1985 250 1990 270
rect 2070 280 2100 365
rect 2260 545 2290 555
rect 2260 525 2265 545
rect 2285 525 2290 545
rect 2260 495 2290 525
rect 2260 475 2265 495
rect 2285 475 2290 495
rect 2260 445 2290 475
rect 2260 425 2265 445
rect 2285 425 2290 445
rect 2260 395 2290 425
rect 2260 375 2265 395
rect 2285 375 2290 395
rect 2070 270 2235 280
rect 2070 250 2170 270
rect 2190 250 2210 270
rect 2230 250 2235 270
rect 1960 220 1990 250
rect 1960 200 1965 220
rect 1985 200 1990 220
rect 1805 160 1845 170
rect 1805 140 1815 160
rect 1835 140 1845 160
rect 1805 130 1845 140
rect 1660 80 1665 100
rect 1685 80 1690 100
rect 1660 50 1690 80
rect 1660 30 1665 50
rect 1685 30 1690 50
rect 1660 20 1690 30
rect 1905 100 1935 110
rect 1905 80 1910 100
rect 1930 80 1935 100
rect 1905 50 1935 80
rect 1905 30 1910 50
rect 1930 30 1935 50
rect 1905 10 1935 30
rect 1960 100 1990 200
rect 2160 220 2235 250
rect 2160 200 2170 220
rect 2190 200 2210 220
rect 2230 200 2235 220
rect 2160 190 2235 200
rect 2260 270 2290 375
rect 2260 250 2265 270
rect 2285 250 2290 270
rect 2260 220 2290 250
rect 2260 200 2265 220
rect 2285 200 2290 220
rect 2105 160 2145 170
rect 2105 140 2115 160
rect 2135 140 2145 160
rect 2105 130 2145 140
rect 1960 80 1965 100
rect 1985 80 1990 100
rect 1960 50 1990 80
rect 1960 30 1965 50
rect 1985 30 1990 50
rect 1960 20 1990 30
rect 2205 100 2235 110
rect 2205 80 2210 100
rect 2230 80 2235 100
rect 2205 50 2235 80
rect 2205 30 2210 50
rect 2230 30 2235 50
rect 2205 10 2235 30
rect 2260 100 2290 200
rect 2260 80 2265 100
rect 2285 80 2290 100
rect 2260 50 2290 80
rect 2260 30 2265 50
rect 2285 30 2290 50
rect 2260 20 2290 30
rect 1425 0 1635 10
rect 1425 -20 1435 0
rect 1455 -20 1635 0
rect 1425 -30 1635 -20
rect 1710 0 1935 10
rect 1710 -20 1720 0
rect 1740 -20 1935 0
rect 1710 -30 1935 -20
rect 2010 0 2235 10
rect 2010 -20 2020 0
rect 2040 -20 2235 0
rect 2010 -30 2235 -20
rect 2310 0 2350 10
rect 2310 -20 2320 0
rect 2340 -20 2350 0
rect 2310 -30 2350 -20
rect 1605 -55 1635 -30
rect 1605 -75 1610 -55
rect 1630 -75 1635 -55
rect 1605 -85 1635 -75
rect 1660 -55 1690 -45
rect 1660 -75 1665 -55
rect 1685 -75 1690 -55
rect 1540 -115 1580 -105
rect 1540 -135 1550 -115
rect 1570 -135 1580 -115
rect 1540 -145 1580 -135
rect 1565 -175 1635 -165
rect 1565 -195 1570 -175
rect 1590 -195 1610 -175
rect 1630 -195 1635 -175
rect 1565 -205 1635 -195
rect 1605 -280 1635 -205
rect 1365 -290 1500 -280
rect 1365 -300 1475 -290
rect 1470 -310 1475 -300
rect 1495 -310 1500 -290
rect 1470 -340 1500 -310
rect 1470 -360 1475 -340
rect 1495 -360 1500 -340
rect 1470 -370 1500 -360
rect 1525 -290 1635 -280
rect 1525 -310 1530 -290
rect 1550 -310 1570 -290
rect 1590 -310 1610 -290
rect 1630 -310 1635 -290
rect 1525 -340 1635 -310
rect 1525 -360 1530 -340
rect 1550 -360 1570 -340
rect 1590 -360 1610 -340
rect 1630 -360 1635 -340
rect 1525 -370 1635 -360
rect 1660 -175 1690 -75
rect 1905 -55 1935 -30
rect 1905 -75 1910 -55
rect 1930 -75 1935 -55
rect 1905 -85 1935 -75
rect 1960 -55 1990 -45
rect 1960 -75 1965 -55
rect 1985 -75 1990 -55
rect 1840 -115 1880 -105
rect 1840 -135 1850 -115
rect 1870 -135 1880 -115
rect 1840 -145 1880 -135
rect 1660 -195 1665 -175
rect 1685 -195 1690 -175
rect 1660 -290 1690 -195
rect 1865 -175 1935 -165
rect 1865 -195 1870 -175
rect 1890 -195 1910 -175
rect 1930 -195 1935 -175
rect 1865 -205 1935 -195
rect 1905 -280 1935 -205
rect 1660 -310 1665 -290
rect 1685 -310 1690 -290
rect 1660 -340 1690 -310
rect 1660 -360 1665 -340
rect 1685 -360 1690 -340
rect 1660 -370 1690 -360
rect 1865 -290 1935 -280
rect 1865 -310 1870 -290
rect 1890 -310 1910 -290
rect 1930 -310 1935 -290
rect 1865 -340 1935 -310
rect 1865 -360 1870 -340
rect 1890 -360 1910 -340
rect 1930 -360 1935 -340
rect 1865 -370 1935 -360
rect 1960 -175 1990 -75
rect 2205 -55 2235 -30
rect 2205 -75 2210 -55
rect 2230 -75 2235 -55
rect 2205 -85 2235 -75
rect 2260 -55 2290 -45
rect 2260 -75 2265 -55
rect 2285 -75 2290 -55
rect 2140 -115 2180 -105
rect 2140 -135 2150 -115
rect 2170 -135 2180 -115
rect 2140 -145 2180 -135
rect 1960 -195 1965 -175
rect 1985 -195 1990 -175
rect 1960 -290 1990 -195
rect 2165 -175 2235 -165
rect 2165 -195 2170 -175
rect 2190 -195 2210 -175
rect 2230 -195 2235 -175
rect 2165 -205 2235 -195
rect 2205 -280 2235 -205
rect 1960 -310 1965 -290
rect 1985 -310 1990 -290
rect 1960 -340 1990 -310
rect 1960 -360 1965 -340
rect 1985 -360 1990 -340
rect 1960 -370 1990 -360
rect 2165 -290 2235 -280
rect 2165 -310 2170 -290
rect 2190 -310 2210 -290
rect 2230 -310 2235 -290
rect 2165 -340 2235 -310
rect 2165 -360 2170 -340
rect 2190 -360 2210 -340
rect 2230 -360 2235 -340
rect 2165 -370 2235 -360
rect 2260 -175 2290 -75
rect 2260 -195 2265 -175
rect 2285 -195 2290 -175
rect 2260 -290 2290 -195
rect 2260 -310 2265 -290
rect 2285 -310 2290 -290
rect 2260 -340 2290 -310
rect 2260 -360 2265 -340
rect 2285 -360 2290 -340
rect 2260 -370 2290 -360
rect 1565 -435 1595 -370
rect 1905 -435 1935 -370
rect 2205 -435 2235 -370
rect 1195 -455 1225 -435
rect 1245 -455 1275 -435
rect 1295 -455 1325 -435
rect 1345 -455 1375 -435
rect 1395 -455 1425 -435
rect 1445 -455 1475 -435
rect 1495 -455 1525 -435
rect 1545 -455 1575 -435
rect 1595 -455 1625 -435
rect 1645 -455 1675 -435
rect 1695 -455 1725 -435
rect 1745 -455 1775 -435
rect 1795 -455 1825 -435
rect 1845 -455 1875 -435
rect 1895 -455 1925 -435
rect 1945 -455 1975 -435
rect 1995 -455 2025 -435
rect 2045 -455 2075 -435
rect 2095 -455 2125 -435
rect 2145 -455 2175 -435
rect 2195 -455 2225 -435
rect 2245 -455 2275 -435
rect 2295 -455 2325 -435
rect 2345 -455 2350 -435
<< viali >>
rect 1225 595 1245 615
rect 1275 595 1295 615
rect 1325 595 1345 615
rect 1375 595 1395 615
rect 1425 595 1445 615
rect 1475 595 1495 615
rect 1525 595 1545 615
rect 1575 595 1595 615
rect 1625 595 1645 615
rect 1675 595 1695 615
rect 1725 595 1745 615
rect 1775 595 1795 615
rect 1825 595 1845 615
rect 1875 595 1895 615
rect 1925 595 1945 615
rect 1975 595 1995 615
rect 2025 595 2045 615
rect 2075 595 2095 615
rect 2125 595 2145 615
rect 2175 595 2195 615
rect 2225 595 2245 615
rect 2275 595 2295 615
rect 2325 595 2345 615
rect 1570 250 1590 270
rect 1570 200 1590 220
rect 1870 250 1890 270
rect 1515 140 1535 160
rect 1870 200 1890 220
rect 2170 250 2190 270
rect 1815 140 1835 160
rect 2170 200 2190 220
rect 2115 140 2135 160
rect 1435 -20 1455 0
rect 2320 -20 2340 0
rect 1550 -135 1570 -115
rect 1570 -195 1590 -175
rect 1610 -195 1630 -175
rect 1850 -135 1870 -115
rect 1870 -195 1890 -175
rect 1910 -195 1930 -175
rect 2150 -135 2170 -115
rect 2170 -195 2190 -175
rect 2210 -195 2230 -175
rect 1225 -455 1245 -435
rect 1275 -455 1295 -435
rect 1325 -455 1345 -435
rect 1375 -455 1395 -435
rect 1425 -455 1445 -435
rect 1475 -455 1495 -435
rect 1525 -455 1545 -435
rect 1575 -455 1595 -435
rect 1625 -455 1645 -435
rect 1675 -455 1695 -435
rect 1725 -455 1745 -435
rect 1775 -455 1795 -435
rect 1825 -455 1845 -435
rect 1875 -455 1895 -435
rect 1925 -455 1945 -435
rect 1975 -455 1995 -435
rect 2025 -455 2045 -435
rect 2075 -455 2095 -435
rect 2125 -455 2145 -435
rect 2175 -455 2195 -435
rect 2225 -455 2245 -435
rect 2275 -455 2295 -435
rect 2325 -455 2345 -435
<< metal1 >>
rect 1195 615 2350 625
rect 1195 595 1225 615
rect 1245 595 1275 615
rect 1295 595 1325 615
rect 1345 595 1375 615
rect 1395 595 1425 615
rect 1445 595 1475 615
rect 1495 595 1525 615
rect 1545 595 1575 615
rect 1595 595 1625 615
rect 1645 595 1675 615
rect 1695 595 1725 615
rect 1745 595 1775 615
rect 1795 595 1825 615
rect 1845 595 1875 615
rect 1895 595 1925 615
rect 1945 595 1975 615
rect 1995 595 2025 615
rect 2045 595 2075 615
rect 2095 595 2125 615
rect 2145 595 2175 615
rect 2195 595 2225 615
rect 2245 595 2275 615
rect 2295 595 2325 615
rect 2345 595 2350 615
rect 1195 585 2350 595
rect 1560 270 1600 280
rect 1560 250 1570 270
rect 1590 250 1600 270
rect 1560 220 1600 250
rect 1560 200 1570 220
rect 1590 200 1600 220
rect 1560 190 1600 200
rect 1860 270 1900 280
rect 1860 250 1870 270
rect 1890 250 1900 270
rect 1860 220 1900 250
rect 1860 200 1870 220
rect 1890 200 1900 220
rect 1860 190 1900 200
rect 2160 270 2200 280
rect 2160 250 2170 270
rect 2190 250 2200 270
rect 2160 220 2200 250
rect 2160 200 2170 220
rect 2190 200 2200 220
rect 2160 190 2200 200
rect 1505 160 1545 170
rect 1505 140 1515 160
rect 1535 140 1545 160
rect 1505 130 1545 140
rect 1425 0 1465 10
rect 1425 -20 1435 0
rect 1455 -20 1465 0
rect 1425 -30 1465 -20
rect 1425 -390 1445 -30
rect 1505 -165 1525 130
rect 1560 -105 1580 190
rect 1540 -115 1580 -105
rect 1540 -135 1550 -115
rect 1570 -135 1580 -115
rect 1540 -145 1580 -135
rect 1805 160 1845 170
rect 1805 140 1815 160
rect 1835 140 1845 160
rect 1805 130 1845 140
rect 1805 -165 1825 130
rect 1860 -105 1880 190
rect 1840 -115 1880 -105
rect 1840 -135 1850 -115
rect 1870 -135 1880 -115
rect 1840 -145 1880 -135
rect 2105 160 2145 170
rect 2105 140 2115 160
rect 2135 140 2145 160
rect 2105 130 2145 140
rect 2105 -165 2125 130
rect 2160 -105 2180 190
rect 2140 -115 2180 -105
rect 2140 -135 2150 -115
rect 2170 -135 2180 -115
rect 2140 -145 2180 -135
rect 2310 0 2350 10
rect 2310 -20 2320 0
rect 2340 -20 2350 0
rect 2310 -30 2350 -20
rect 1505 -175 1635 -165
rect 1505 -195 1570 -175
rect 1590 -195 1610 -175
rect 1630 -195 1635 -175
rect 1505 -205 1635 -195
rect 1805 -175 1935 -165
rect 1805 -195 1870 -175
rect 1890 -195 1910 -175
rect 1930 -195 1935 -175
rect 1805 -205 1935 -195
rect 2105 -175 2235 -165
rect 2105 -195 2170 -175
rect 2190 -195 2210 -175
rect 2230 -195 2235 -175
rect 2105 -205 2235 -195
rect 2310 -390 2330 -30
rect 1425 -410 2330 -390
rect 1195 -435 2350 -425
rect 1195 -455 1225 -435
rect 1245 -455 1275 -435
rect 1295 -455 1325 -435
rect 1345 -455 1375 -435
rect 1395 -455 1425 -435
rect 1445 -455 1475 -435
rect 1495 -455 1525 -435
rect 1545 -455 1575 -435
rect 1595 -455 1625 -435
rect 1645 -455 1675 -435
rect 1695 -455 1725 -435
rect 1745 -455 1775 -435
rect 1795 -455 1825 -435
rect 1845 -455 1875 -435
rect 1895 -455 1925 -435
rect 1945 -455 1975 -435
rect 1995 -455 2025 -435
rect 2045 -455 2075 -435
rect 2095 -455 2125 -435
rect 2145 -455 2175 -435
rect 2195 -455 2225 -435
rect 2245 -455 2275 -435
rect 2295 -455 2325 -435
rect 2345 -455 2350 -435
rect 1195 -465 2350 -455
<< labels >>
flabel locali 1770 10 1770 10 1 FreeSans 400 0 0 200 V8
flabel locali 2080 10 2080 10 1 FreeSans 400 0 0 200 V9
flabel locali 1690 310 1690 310 3 FreeSans 400 0 200 0 V2
flabel locali 1690 -235 1690 -235 3 FreeSans 400 0 200 0 V3
flabel locali 1990 320 1990 320 3 FreeSans 400 0 200 0 V4
flabel locali 1990 -235 1990 -235 3 FreeSans 400 0 200 0 V5
flabel locali 2290 320 2290 320 3 FreeSans 400 0 200 0 V6
flabel locali 2290 -235 2290 -235 3 FreeSans 400 0 200 0 V7
flabel locali 1365 -85 1365 -85 7 FreeSans 400 0 -200 0 V1
<< end >>
