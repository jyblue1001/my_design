magic
tech sky130A
magscale 1 2
timestamp 1746453344
<< nwell >>
rect 4300 3700 9310 5490
<< pwell >>
rect 1500 1320 2550 1340
rect 2630 1320 2670 1340
rect 1370 1187 2670 1320
rect 1370 153 1503 1187
rect 2537 153 2670 1187
rect 40 50 80 90
rect 1370 20 2670 153
rect 2710 1320 2770 1340
rect 2850 1320 4050 1340
rect 2710 1187 4050 1320
rect 2710 153 2863 1187
rect 3897 153 4050 1187
rect 2710 20 4050 153
rect 4070 1187 5390 1340
rect 4070 153 4223 1187
rect 5257 153 5390 1187
rect 4070 20 5390 153
rect 5430 1187 6750 1340
rect 5430 153 5583 1187
rect 6617 153 6750 1187
rect 5430 20 6750 153
rect 6790 1187 8110 1340
rect 6790 153 6943 1187
rect 7977 153 8110 1187
rect 6790 20 8110 153
rect 8150 1187 9470 1340
rect 8150 153 8303 1187
rect 9337 153 9470 1187
rect 8150 20 9470 153
<< nbase >>
rect 1503 153 2537 1187
rect 2863 153 3897 1187
rect 4223 153 5257 1187
rect 5583 153 6617 1187
rect 6943 153 7977 1187
rect 8303 153 9337 1187
<< nmos >>
rect 5220 3130 5340 3330
rect 5420 3130 5540 3330
rect 5620 3130 5740 3330
rect 5820 3130 5940 3330
rect 6020 3130 6140 3330
rect 6220 3130 6340 3330
rect 6580 3130 6700 3330
rect 6780 3130 6900 3330
rect 6980 3130 7100 3330
rect 7180 3130 7300 3330
rect 7380 3130 7500 3330
rect 7580 3130 7700 3330
rect 4740 1980 5540 2780
rect 5620 1980 6420 2780
rect 6500 1980 7300 2780
rect 7380 1980 8180 2780
rect 5440 1510 7440 1710
<< pmos >>
rect 4500 4650 4620 5450
rect 4700 4650 4820 5450
rect 4900 4650 5020 5450
rect 5100 4650 5220 5450
rect 5300 4650 5420 5450
rect 5500 4650 5620 5450
rect 5700 4650 5820 5450
rect 5900 4650 6020 5450
rect 6100 4650 6220 5450
rect 6300 4650 6420 5450
rect 6500 4650 6620 5450
rect 6700 4650 6820 5450
rect 6900 4650 7020 5450
rect 7100 4650 7220 5450
rect 7300 4650 7420 5450
rect 7500 4650 7620 5450
rect 7700 4650 7820 5450
rect 7900 4650 8020 5450
rect 8100 4650 8220 5450
rect 8300 4650 8420 5450
rect 4540 3740 4660 4140
rect 4740 3740 4860 4140
rect 4940 3740 5060 4140
rect 5140 3740 5260 4140
rect 5340 3740 5460 4140
rect 5540 3740 5660 4140
rect 5900 3740 6020 4140
rect 6100 3740 6220 4140
rect 6300 3740 6420 4140
rect 6500 3740 6620 4140
rect 6700 3740 6820 4140
rect 6900 3740 7020 4140
rect 7260 3740 7380 4140
rect 7460 3740 7580 4140
rect 7660 3740 7780 4140
rect 7860 3740 7980 4140
rect 8060 3740 8180 4140
rect 8260 3740 8380 4140
rect 8830 3740 8860 4140
rect 9080 3740 9110 4140
<< ndiff >>
rect 5140 3300 5220 3330
rect 5140 3260 5160 3300
rect 5200 3260 5220 3300
rect 5140 3200 5220 3260
rect 5140 3160 5160 3200
rect 5200 3160 5220 3200
rect 5140 3130 5220 3160
rect 5340 3300 5420 3330
rect 5340 3260 5360 3300
rect 5400 3260 5420 3300
rect 5340 3200 5420 3260
rect 5340 3160 5360 3200
rect 5400 3160 5420 3200
rect 5340 3130 5420 3160
rect 5540 3300 5620 3330
rect 5540 3260 5560 3300
rect 5600 3260 5620 3300
rect 5540 3200 5620 3260
rect 5540 3160 5560 3200
rect 5600 3160 5620 3200
rect 5540 3130 5620 3160
rect 5740 3300 5820 3330
rect 5740 3260 5760 3300
rect 5800 3260 5820 3300
rect 5740 3200 5820 3260
rect 5740 3160 5760 3200
rect 5800 3160 5820 3200
rect 5740 3130 5820 3160
rect 5940 3300 6020 3330
rect 5940 3260 5960 3300
rect 6000 3260 6020 3300
rect 5940 3200 6020 3260
rect 5940 3160 5960 3200
rect 6000 3160 6020 3200
rect 5940 3130 6020 3160
rect 6140 3300 6220 3330
rect 6140 3260 6160 3300
rect 6200 3260 6220 3300
rect 6140 3200 6220 3260
rect 6140 3160 6160 3200
rect 6200 3160 6220 3200
rect 6140 3130 6220 3160
rect 6340 3300 6420 3330
rect 6500 3300 6580 3330
rect 6340 3260 6360 3300
rect 6400 3260 6420 3300
rect 6500 3260 6520 3300
rect 6560 3260 6580 3300
rect 6340 3200 6420 3260
rect 6500 3200 6580 3260
rect 6340 3160 6360 3200
rect 6400 3160 6420 3200
rect 6500 3160 6520 3200
rect 6560 3160 6580 3200
rect 6340 3130 6420 3160
rect 6500 3130 6580 3160
rect 6700 3300 6780 3330
rect 6700 3260 6720 3300
rect 6760 3260 6780 3300
rect 6700 3200 6780 3260
rect 6700 3160 6720 3200
rect 6760 3160 6780 3200
rect 6700 3130 6780 3160
rect 6900 3300 6980 3330
rect 6900 3260 6920 3300
rect 6960 3260 6980 3300
rect 6900 3200 6980 3260
rect 6900 3160 6920 3200
rect 6960 3160 6980 3200
rect 6900 3130 6980 3160
rect 7100 3300 7180 3330
rect 7100 3260 7120 3300
rect 7160 3260 7180 3300
rect 7100 3200 7180 3260
rect 7100 3160 7120 3200
rect 7160 3160 7180 3200
rect 7100 3130 7180 3160
rect 7300 3300 7380 3330
rect 7300 3260 7320 3300
rect 7360 3260 7380 3300
rect 7300 3200 7380 3260
rect 7300 3160 7320 3200
rect 7360 3160 7380 3200
rect 7300 3130 7380 3160
rect 7500 3300 7580 3330
rect 7500 3260 7520 3300
rect 7560 3260 7580 3300
rect 7500 3200 7580 3260
rect 7500 3160 7520 3200
rect 7560 3160 7580 3200
rect 7500 3130 7580 3160
rect 7700 3300 7780 3330
rect 7700 3260 7720 3300
rect 7760 3260 7780 3300
rect 7700 3200 7780 3260
rect 7700 3160 7720 3200
rect 7760 3160 7780 3200
rect 7700 3130 7780 3160
rect 4660 2750 4740 2780
rect 4660 2710 4680 2750
rect 4720 2710 4740 2750
rect 4660 2650 4740 2710
rect 4660 2610 4680 2650
rect 4720 2610 4740 2650
rect 4660 2550 4740 2610
rect 4660 2510 4680 2550
rect 4720 2510 4740 2550
rect 4660 2450 4740 2510
rect 4660 2410 4680 2450
rect 4720 2410 4740 2450
rect 4660 2350 4740 2410
rect 4660 2310 4680 2350
rect 4720 2310 4740 2350
rect 4660 2250 4740 2310
rect 4660 2210 4680 2250
rect 4720 2210 4740 2250
rect 4660 2150 4740 2210
rect 4660 2110 4680 2150
rect 4720 2110 4740 2150
rect 4660 2050 4740 2110
rect 4660 2010 4680 2050
rect 4720 2010 4740 2050
rect 4660 1980 4740 2010
rect 5540 2750 5620 2780
rect 5540 2710 5560 2750
rect 5600 2710 5620 2750
rect 5540 2650 5620 2710
rect 5540 2610 5560 2650
rect 5600 2610 5620 2650
rect 5540 2550 5620 2610
rect 5540 2510 5560 2550
rect 5600 2510 5620 2550
rect 5540 2450 5620 2510
rect 5540 2410 5560 2450
rect 5600 2410 5620 2450
rect 5540 2350 5620 2410
rect 5540 2310 5560 2350
rect 5600 2310 5620 2350
rect 5540 2250 5620 2310
rect 5540 2210 5560 2250
rect 5600 2210 5620 2250
rect 5540 2150 5620 2210
rect 5540 2110 5560 2150
rect 5600 2110 5620 2150
rect 5540 2050 5620 2110
rect 5540 2010 5560 2050
rect 5600 2010 5620 2050
rect 5540 1980 5620 2010
rect 6420 2750 6500 2780
rect 6420 2710 6440 2750
rect 6480 2710 6500 2750
rect 6420 2650 6500 2710
rect 6420 2610 6440 2650
rect 6480 2610 6500 2650
rect 6420 2550 6500 2610
rect 6420 2510 6440 2550
rect 6480 2510 6500 2550
rect 6420 2450 6500 2510
rect 6420 2410 6440 2450
rect 6480 2410 6500 2450
rect 6420 2350 6500 2410
rect 6420 2310 6440 2350
rect 6480 2310 6500 2350
rect 6420 2250 6500 2310
rect 6420 2210 6440 2250
rect 6480 2210 6500 2250
rect 6420 2150 6500 2210
rect 6420 2110 6440 2150
rect 6480 2110 6500 2150
rect 6420 2050 6500 2110
rect 6420 2010 6440 2050
rect 6480 2010 6500 2050
rect 6420 1980 6500 2010
rect 7300 2750 7380 2780
rect 7300 2710 7320 2750
rect 7360 2710 7380 2750
rect 7300 2650 7380 2710
rect 7300 2610 7320 2650
rect 7360 2610 7380 2650
rect 7300 2550 7380 2610
rect 7300 2510 7320 2550
rect 7360 2510 7380 2550
rect 7300 2450 7380 2510
rect 7300 2410 7320 2450
rect 7360 2410 7380 2450
rect 7300 2350 7380 2410
rect 7300 2310 7320 2350
rect 7360 2310 7380 2350
rect 7300 2250 7380 2310
rect 7300 2210 7320 2250
rect 7360 2210 7380 2250
rect 7300 2150 7380 2210
rect 7300 2110 7320 2150
rect 7360 2110 7380 2150
rect 7300 2050 7380 2110
rect 7300 2010 7320 2050
rect 7360 2010 7380 2050
rect 7300 1980 7380 2010
rect 8180 2750 8260 2780
rect 8180 2710 8200 2750
rect 8240 2710 8260 2750
rect 8180 2650 8260 2710
rect 8180 2610 8200 2650
rect 8240 2610 8260 2650
rect 8180 2550 8260 2610
rect 8180 2510 8200 2550
rect 8240 2510 8260 2550
rect 8180 2450 8260 2510
rect 8180 2410 8200 2450
rect 8240 2410 8260 2450
rect 8180 2350 8260 2410
rect 8180 2310 8200 2350
rect 8240 2310 8260 2350
rect 8180 2250 8260 2310
rect 8180 2210 8200 2250
rect 8240 2210 8260 2250
rect 8180 2150 8260 2210
rect 8180 2110 8200 2150
rect 8240 2110 8260 2150
rect 8180 2050 8260 2110
rect 8180 2010 8200 2050
rect 8240 2010 8260 2050
rect 8180 1980 8260 2010
rect 5360 1680 5440 1710
rect 5360 1640 5380 1680
rect 5420 1640 5440 1680
rect 5360 1580 5440 1640
rect 5360 1540 5380 1580
rect 5420 1540 5440 1580
rect 5360 1510 5440 1540
rect 7440 1680 7520 1710
rect 7440 1640 7460 1680
rect 7500 1640 7520 1680
rect 7440 1580 7520 1640
rect 7440 1540 7460 1580
rect 7500 1540 7520 1580
rect 7440 1510 7520 1540
<< pdiff >>
rect 4420 5420 4500 5450
rect 4420 5380 4440 5420
rect 4480 5380 4500 5420
rect 4420 5320 4500 5380
rect 4420 5280 4440 5320
rect 4480 5280 4500 5320
rect 4420 5220 4500 5280
rect 4420 5180 4440 5220
rect 4480 5180 4500 5220
rect 4420 5120 4500 5180
rect 4420 5080 4440 5120
rect 4480 5080 4500 5120
rect 4420 5020 4500 5080
rect 4420 4980 4440 5020
rect 4480 4980 4500 5020
rect 4420 4920 4500 4980
rect 4420 4880 4440 4920
rect 4480 4880 4500 4920
rect 4420 4820 4500 4880
rect 4420 4780 4440 4820
rect 4480 4780 4500 4820
rect 4420 4720 4500 4780
rect 4420 4680 4440 4720
rect 4480 4680 4500 4720
rect 4420 4650 4500 4680
rect 4620 5420 4700 5450
rect 4620 5380 4640 5420
rect 4680 5380 4700 5420
rect 4620 5320 4700 5380
rect 4620 5280 4640 5320
rect 4680 5280 4700 5320
rect 4620 5220 4700 5280
rect 4620 5180 4640 5220
rect 4680 5180 4700 5220
rect 4620 5120 4700 5180
rect 4620 5080 4640 5120
rect 4680 5080 4700 5120
rect 4620 5020 4700 5080
rect 4620 4980 4640 5020
rect 4680 4980 4700 5020
rect 4620 4920 4700 4980
rect 4620 4880 4640 4920
rect 4680 4880 4700 4920
rect 4620 4820 4700 4880
rect 4620 4780 4640 4820
rect 4680 4780 4700 4820
rect 4620 4720 4700 4780
rect 4620 4680 4640 4720
rect 4680 4680 4700 4720
rect 4620 4650 4700 4680
rect 4820 5420 4900 5450
rect 4820 5380 4840 5420
rect 4880 5380 4900 5420
rect 4820 5320 4900 5380
rect 4820 5280 4840 5320
rect 4880 5280 4900 5320
rect 4820 5220 4900 5280
rect 4820 5180 4840 5220
rect 4880 5180 4900 5220
rect 4820 5120 4900 5180
rect 4820 5080 4840 5120
rect 4880 5080 4900 5120
rect 4820 5020 4900 5080
rect 4820 4980 4840 5020
rect 4880 4980 4900 5020
rect 4820 4920 4900 4980
rect 4820 4880 4840 4920
rect 4880 4880 4900 4920
rect 4820 4820 4900 4880
rect 4820 4780 4840 4820
rect 4880 4780 4900 4820
rect 4820 4720 4900 4780
rect 4820 4680 4840 4720
rect 4880 4680 4900 4720
rect 4820 4650 4900 4680
rect 5020 5420 5100 5450
rect 5020 5380 5040 5420
rect 5080 5380 5100 5420
rect 5020 5320 5100 5380
rect 5020 5280 5040 5320
rect 5080 5280 5100 5320
rect 5020 5220 5100 5280
rect 5020 5180 5040 5220
rect 5080 5180 5100 5220
rect 5020 5120 5100 5180
rect 5020 5080 5040 5120
rect 5080 5080 5100 5120
rect 5020 5020 5100 5080
rect 5020 4980 5040 5020
rect 5080 4980 5100 5020
rect 5020 4920 5100 4980
rect 5020 4880 5040 4920
rect 5080 4880 5100 4920
rect 5020 4820 5100 4880
rect 5020 4780 5040 4820
rect 5080 4780 5100 4820
rect 5020 4720 5100 4780
rect 5020 4680 5040 4720
rect 5080 4680 5100 4720
rect 5020 4650 5100 4680
rect 5220 5420 5300 5450
rect 5220 5380 5240 5420
rect 5280 5380 5300 5420
rect 5220 5320 5300 5380
rect 5220 5280 5240 5320
rect 5280 5280 5300 5320
rect 5220 5220 5300 5280
rect 5220 5180 5240 5220
rect 5280 5180 5300 5220
rect 5220 5120 5300 5180
rect 5220 5080 5240 5120
rect 5280 5080 5300 5120
rect 5220 5020 5300 5080
rect 5220 4980 5240 5020
rect 5280 4980 5300 5020
rect 5220 4920 5300 4980
rect 5220 4880 5240 4920
rect 5280 4880 5300 4920
rect 5220 4820 5300 4880
rect 5220 4780 5240 4820
rect 5280 4780 5300 4820
rect 5220 4720 5300 4780
rect 5220 4680 5240 4720
rect 5280 4680 5300 4720
rect 5220 4650 5300 4680
rect 5420 5420 5500 5450
rect 5420 5380 5440 5420
rect 5480 5380 5500 5420
rect 5420 5320 5500 5380
rect 5420 5280 5440 5320
rect 5480 5280 5500 5320
rect 5420 5220 5500 5280
rect 5420 5180 5440 5220
rect 5480 5180 5500 5220
rect 5420 5120 5500 5180
rect 5420 5080 5440 5120
rect 5480 5080 5500 5120
rect 5420 5020 5500 5080
rect 5420 4980 5440 5020
rect 5480 4980 5500 5020
rect 5420 4920 5500 4980
rect 5420 4880 5440 4920
rect 5480 4880 5500 4920
rect 5420 4820 5500 4880
rect 5420 4780 5440 4820
rect 5480 4780 5500 4820
rect 5420 4720 5500 4780
rect 5420 4680 5440 4720
rect 5480 4680 5500 4720
rect 5420 4650 5500 4680
rect 5620 5420 5700 5450
rect 5620 5380 5640 5420
rect 5680 5380 5700 5420
rect 5620 5320 5700 5380
rect 5620 5280 5640 5320
rect 5680 5280 5700 5320
rect 5620 5220 5700 5280
rect 5620 5180 5640 5220
rect 5680 5180 5700 5220
rect 5620 5120 5700 5180
rect 5620 5080 5640 5120
rect 5680 5080 5700 5120
rect 5620 5020 5700 5080
rect 5620 4980 5640 5020
rect 5680 4980 5700 5020
rect 5620 4920 5700 4980
rect 5620 4880 5640 4920
rect 5680 4880 5700 4920
rect 5620 4820 5700 4880
rect 5620 4780 5640 4820
rect 5680 4780 5700 4820
rect 5620 4720 5700 4780
rect 5620 4680 5640 4720
rect 5680 4680 5700 4720
rect 5620 4650 5700 4680
rect 5820 5420 5900 5450
rect 5820 5380 5840 5420
rect 5880 5380 5900 5420
rect 5820 5320 5900 5380
rect 5820 5280 5840 5320
rect 5880 5280 5900 5320
rect 5820 5220 5900 5280
rect 5820 5180 5840 5220
rect 5880 5180 5900 5220
rect 5820 5120 5900 5180
rect 5820 5080 5840 5120
rect 5880 5080 5900 5120
rect 5820 5020 5900 5080
rect 5820 4980 5840 5020
rect 5880 4980 5900 5020
rect 5820 4920 5900 4980
rect 5820 4880 5840 4920
rect 5880 4880 5900 4920
rect 5820 4820 5900 4880
rect 5820 4780 5840 4820
rect 5880 4780 5900 4820
rect 5820 4720 5900 4780
rect 5820 4680 5840 4720
rect 5880 4680 5900 4720
rect 5820 4650 5900 4680
rect 6020 5420 6100 5450
rect 6020 5380 6040 5420
rect 6080 5380 6100 5420
rect 6020 5320 6100 5380
rect 6020 5280 6040 5320
rect 6080 5280 6100 5320
rect 6020 5220 6100 5280
rect 6020 5180 6040 5220
rect 6080 5180 6100 5220
rect 6020 5120 6100 5180
rect 6020 5080 6040 5120
rect 6080 5080 6100 5120
rect 6020 5020 6100 5080
rect 6020 4980 6040 5020
rect 6080 4980 6100 5020
rect 6020 4920 6100 4980
rect 6020 4880 6040 4920
rect 6080 4880 6100 4920
rect 6020 4820 6100 4880
rect 6020 4780 6040 4820
rect 6080 4780 6100 4820
rect 6020 4720 6100 4780
rect 6020 4680 6040 4720
rect 6080 4680 6100 4720
rect 6020 4650 6100 4680
rect 6220 5420 6300 5450
rect 6220 5380 6240 5420
rect 6280 5380 6300 5420
rect 6220 5320 6300 5380
rect 6220 5280 6240 5320
rect 6280 5280 6300 5320
rect 6220 5220 6300 5280
rect 6220 5180 6240 5220
rect 6280 5180 6300 5220
rect 6220 5120 6300 5180
rect 6220 5080 6240 5120
rect 6280 5080 6300 5120
rect 6220 5020 6300 5080
rect 6220 4980 6240 5020
rect 6280 4980 6300 5020
rect 6220 4920 6300 4980
rect 6220 4880 6240 4920
rect 6280 4880 6300 4920
rect 6220 4820 6300 4880
rect 6220 4780 6240 4820
rect 6280 4780 6300 4820
rect 6220 4720 6300 4780
rect 6220 4680 6240 4720
rect 6280 4680 6300 4720
rect 6220 4650 6300 4680
rect 6420 5420 6500 5450
rect 6420 5380 6440 5420
rect 6480 5380 6500 5420
rect 6420 5320 6500 5380
rect 6420 5280 6440 5320
rect 6480 5280 6500 5320
rect 6420 5220 6500 5280
rect 6420 5180 6440 5220
rect 6480 5180 6500 5220
rect 6420 5120 6500 5180
rect 6420 5080 6440 5120
rect 6480 5080 6500 5120
rect 6420 5020 6500 5080
rect 6420 4980 6440 5020
rect 6480 4980 6500 5020
rect 6420 4920 6500 4980
rect 6420 4880 6440 4920
rect 6480 4880 6500 4920
rect 6420 4820 6500 4880
rect 6420 4780 6440 4820
rect 6480 4780 6500 4820
rect 6420 4720 6500 4780
rect 6420 4680 6440 4720
rect 6480 4680 6500 4720
rect 6420 4650 6500 4680
rect 6620 5420 6700 5450
rect 6620 5380 6640 5420
rect 6680 5380 6700 5420
rect 6620 5320 6700 5380
rect 6620 5280 6640 5320
rect 6680 5280 6700 5320
rect 6620 5220 6700 5280
rect 6620 5180 6640 5220
rect 6680 5180 6700 5220
rect 6620 5120 6700 5180
rect 6620 5080 6640 5120
rect 6680 5080 6700 5120
rect 6620 5020 6700 5080
rect 6620 4980 6640 5020
rect 6680 4980 6700 5020
rect 6620 4920 6700 4980
rect 6620 4880 6640 4920
rect 6680 4880 6700 4920
rect 6620 4820 6700 4880
rect 6620 4780 6640 4820
rect 6680 4780 6700 4820
rect 6620 4720 6700 4780
rect 6620 4680 6640 4720
rect 6680 4680 6700 4720
rect 6620 4650 6700 4680
rect 6820 5420 6900 5450
rect 6820 5380 6840 5420
rect 6880 5380 6900 5420
rect 6820 5320 6900 5380
rect 6820 5280 6840 5320
rect 6880 5280 6900 5320
rect 6820 5220 6900 5280
rect 6820 5180 6840 5220
rect 6880 5180 6900 5220
rect 6820 5120 6900 5180
rect 6820 5080 6840 5120
rect 6880 5080 6900 5120
rect 6820 5020 6900 5080
rect 6820 4980 6840 5020
rect 6880 4980 6900 5020
rect 6820 4920 6900 4980
rect 6820 4880 6840 4920
rect 6880 4880 6900 4920
rect 6820 4820 6900 4880
rect 6820 4780 6840 4820
rect 6880 4780 6900 4820
rect 6820 4720 6900 4780
rect 6820 4680 6840 4720
rect 6880 4680 6900 4720
rect 6820 4650 6900 4680
rect 7020 5420 7100 5450
rect 7020 5380 7040 5420
rect 7080 5380 7100 5420
rect 7020 5320 7100 5380
rect 7020 5280 7040 5320
rect 7080 5280 7100 5320
rect 7020 5220 7100 5280
rect 7020 5180 7040 5220
rect 7080 5180 7100 5220
rect 7020 5120 7100 5180
rect 7020 5080 7040 5120
rect 7080 5080 7100 5120
rect 7020 5020 7100 5080
rect 7020 4980 7040 5020
rect 7080 4980 7100 5020
rect 7020 4920 7100 4980
rect 7020 4880 7040 4920
rect 7080 4880 7100 4920
rect 7020 4820 7100 4880
rect 7020 4780 7040 4820
rect 7080 4780 7100 4820
rect 7020 4720 7100 4780
rect 7020 4680 7040 4720
rect 7080 4680 7100 4720
rect 7020 4650 7100 4680
rect 7220 5420 7300 5450
rect 7220 5380 7240 5420
rect 7280 5380 7300 5420
rect 7220 5320 7300 5380
rect 7220 5280 7240 5320
rect 7280 5280 7300 5320
rect 7220 5220 7300 5280
rect 7220 5180 7240 5220
rect 7280 5180 7300 5220
rect 7220 5120 7300 5180
rect 7220 5080 7240 5120
rect 7280 5080 7300 5120
rect 7220 5020 7300 5080
rect 7220 4980 7240 5020
rect 7280 4980 7300 5020
rect 7220 4920 7300 4980
rect 7220 4880 7240 4920
rect 7280 4880 7300 4920
rect 7220 4820 7300 4880
rect 7220 4780 7240 4820
rect 7280 4780 7300 4820
rect 7220 4720 7300 4780
rect 7220 4680 7240 4720
rect 7280 4680 7300 4720
rect 7220 4650 7300 4680
rect 7420 5420 7500 5450
rect 7420 5380 7440 5420
rect 7480 5380 7500 5420
rect 7420 5320 7500 5380
rect 7420 5280 7440 5320
rect 7480 5280 7500 5320
rect 7420 5220 7500 5280
rect 7420 5180 7440 5220
rect 7480 5180 7500 5220
rect 7420 5120 7500 5180
rect 7420 5080 7440 5120
rect 7480 5080 7500 5120
rect 7420 5020 7500 5080
rect 7420 4980 7440 5020
rect 7480 4980 7500 5020
rect 7420 4920 7500 4980
rect 7420 4880 7440 4920
rect 7480 4880 7500 4920
rect 7420 4820 7500 4880
rect 7420 4780 7440 4820
rect 7480 4780 7500 4820
rect 7420 4720 7500 4780
rect 7420 4680 7440 4720
rect 7480 4680 7500 4720
rect 7420 4650 7500 4680
rect 7620 5420 7700 5450
rect 7620 5380 7640 5420
rect 7680 5380 7700 5420
rect 7620 5320 7700 5380
rect 7620 5280 7640 5320
rect 7680 5280 7700 5320
rect 7620 5220 7700 5280
rect 7620 5180 7640 5220
rect 7680 5180 7700 5220
rect 7620 5120 7700 5180
rect 7620 5080 7640 5120
rect 7680 5080 7700 5120
rect 7620 5020 7700 5080
rect 7620 4980 7640 5020
rect 7680 4980 7700 5020
rect 7620 4920 7700 4980
rect 7620 4880 7640 4920
rect 7680 4880 7700 4920
rect 7620 4820 7700 4880
rect 7620 4780 7640 4820
rect 7680 4780 7700 4820
rect 7620 4720 7700 4780
rect 7620 4680 7640 4720
rect 7680 4680 7700 4720
rect 7620 4650 7700 4680
rect 7820 5420 7900 5450
rect 7820 5380 7840 5420
rect 7880 5380 7900 5420
rect 7820 5320 7900 5380
rect 7820 5280 7840 5320
rect 7880 5280 7900 5320
rect 7820 5220 7900 5280
rect 7820 5180 7840 5220
rect 7880 5180 7900 5220
rect 7820 5120 7900 5180
rect 7820 5080 7840 5120
rect 7880 5080 7900 5120
rect 7820 5020 7900 5080
rect 7820 4980 7840 5020
rect 7880 4980 7900 5020
rect 7820 4920 7900 4980
rect 7820 4880 7840 4920
rect 7880 4880 7900 4920
rect 7820 4820 7900 4880
rect 7820 4780 7840 4820
rect 7880 4780 7900 4820
rect 7820 4720 7900 4780
rect 7820 4680 7840 4720
rect 7880 4680 7900 4720
rect 7820 4650 7900 4680
rect 8020 5420 8100 5450
rect 8020 5380 8040 5420
rect 8080 5380 8100 5420
rect 8020 5320 8100 5380
rect 8020 5280 8040 5320
rect 8080 5280 8100 5320
rect 8020 5220 8100 5280
rect 8020 5180 8040 5220
rect 8080 5180 8100 5220
rect 8020 5120 8100 5180
rect 8020 5080 8040 5120
rect 8080 5080 8100 5120
rect 8020 5020 8100 5080
rect 8020 4980 8040 5020
rect 8080 4980 8100 5020
rect 8020 4920 8100 4980
rect 8020 4880 8040 4920
rect 8080 4880 8100 4920
rect 8020 4820 8100 4880
rect 8020 4780 8040 4820
rect 8080 4780 8100 4820
rect 8020 4720 8100 4780
rect 8020 4680 8040 4720
rect 8080 4680 8100 4720
rect 8020 4650 8100 4680
rect 8220 5420 8300 5450
rect 8220 5380 8240 5420
rect 8280 5380 8300 5420
rect 8220 5320 8300 5380
rect 8220 5280 8240 5320
rect 8280 5280 8300 5320
rect 8220 5220 8300 5280
rect 8220 5180 8240 5220
rect 8280 5180 8300 5220
rect 8220 5120 8300 5180
rect 8220 5080 8240 5120
rect 8280 5080 8300 5120
rect 8220 5020 8300 5080
rect 8220 4980 8240 5020
rect 8280 4980 8300 5020
rect 8220 4920 8300 4980
rect 8220 4880 8240 4920
rect 8280 4880 8300 4920
rect 8220 4820 8300 4880
rect 8220 4780 8240 4820
rect 8280 4780 8300 4820
rect 8220 4720 8300 4780
rect 8220 4680 8240 4720
rect 8280 4680 8300 4720
rect 8220 4650 8300 4680
rect 8420 5420 8500 5450
rect 8420 5380 8440 5420
rect 8480 5380 8500 5420
rect 8420 5320 8500 5380
rect 8420 5280 8440 5320
rect 8480 5280 8500 5320
rect 8420 5220 8500 5280
rect 8420 5180 8440 5220
rect 8480 5180 8500 5220
rect 8420 5120 8500 5180
rect 8420 5080 8440 5120
rect 8480 5080 8500 5120
rect 8420 5020 8500 5080
rect 8420 4980 8440 5020
rect 8480 4980 8500 5020
rect 8420 4920 8500 4980
rect 8420 4880 8440 4920
rect 8480 4880 8500 4920
rect 8420 4820 8500 4880
rect 8420 4780 8440 4820
rect 8480 4780 8500 4820
rect 8420 4720 8500 4780
rect 8420 4680 8440 4720
rect 8480 4680 8500 4720
rect 8420 4650 8500 4680
rect 4460 4110 4540 4140
rect 4460 4070 4480 4110
rect 4520 4070 4540 4110
rect 4460 4010 4540 4070
rect 4460 3970 4480 4010
rect 4520 3970 4540 4010
rect 4460 3910 4540 3970
rect 4460 3870 4480 3910
rect 4520 3870 4540 3910
rect 4460 3810 4540 3870
rect 4460 3770 4480 3810
rect 4520 3770 4540 3810
rect 4460 3740 4540 3770
rect 4660 4110 4740 4140
rect 4660 4070 4680 4110
rect 4720 4070 4740 4110
rect 4660 4010 4740 4070
rect 4660 3970 4680 4010
rect 4720 3970 4740 4010
rect 4660 3910 4740 3970
rect 4660 3870 4680 3910
rect 4720 3870 4740 3910
rect 4660 3810 4740 3870
rect 4660 3770 4680 3810
rect 4720 3770 4740 3810
rect 4660 3740 4740 3770
rect 4860 4110 4940 4140
rect 4860 4070 4880 4110
rect 4920 4070 4940 4110
rect 4860 4010 4940 4070
rect 4860 3970 4880 4010
rect 4920 3970 4940 4010
rect 4860 3910 4940 3970
rect 4860 3870 4880 3910
rect 4920 3870 4940 3910
rect 4860 3810 4940 3870
rect 4860 3770 4880 3810
rect 4920 3770 4940 3810
rect 4860 3740 4940 3770
rect 5060 4110 5140 4140
rect 5060 4070 5080 4110
rect 5120 4070 5140 4110
rect 5060 4010 5140 4070
rect 5060 3970 5080 4010
rect 5120 3970 5140 4010
rect 5060 3910 5140 3970
rect 5060 3870 5080 3910
rect 5120 3870 5140 3910
rect 5060 3810 5140 3870
rect 5060 3770 5080 3810
rect 5120 3770 5140 3810
rect 5060 3740 5140 3770
rect 5260 4110 5340 4140
rect 5260 4070 5280 4110
rect 5320 4070 5340 4110
rect 5260 4010 5340 4070
rect 5260 3970 5280 4010
rect 5320 3970 5340 4010
rect 5260 3910 5340 3970
rect 5260 3870 5280 3910
rect 5320 3870 5340 3910
rect 5260 3810 5340 3870
rect 5260 3770 5280 3810
rect 5320 3770 5340 3810
rect 5260 3740 5340 3770
rect 5460 4110 5540 4140
rect 5460 4070 5480 4110
rect 5520 4070 5540 4110
rect 5460 4010 5540 4070
rect 5460 3970 5480 4010
rect 5520 3970 5540 4010
rect 5460 3910 5540 3970
rect 5460 3870 5480 3910
rect 5520 3870 5540 3910
rect 5460 3810 5540 3870
rect 5460 3770 5480 3810
rect 5520 3770 5540 3810
rect 5460 3740 5540 3770
rect 5660 4110 5740 4140
rect 5820 4110 5900 4140
rect 5660 4070 5680 4110
rect 5720 4070 5740 4110
rect 5820 4070 5840 4110
rect 5880 4070 5900 4110
rect 5660 4010 5740 4070
rect 5820 4010 5900 4070
rect 5660 3970 5680 4010
rect 5720 3970 5740 4010
rect 5820 3970 5840 4010
rect 5880 3970 5900 4010
rect 5660 3910 5740 3970
rect 5820 3910 5900 3970
rect 5660 3870 5680 3910
rect 5720 3870 5740 3910
rect 5820 3870 5840 3910
rect 5880 3870 5900 3910
rect 5660 3810 5740 3870
rect 5820 3810 5900 3870
rect 5660 3770 5680 3810
rect 5720 3770 5740 3810
rect 5820 3770 5840 3810
rect 5880 3770 5900 3810
rect 5660 3740 5740 3770
rect 5820 3740 5900 3770
rect 6020 4110 6100 4140
rect 6020 4070 6040 4110
rect 6080 4070 6100 4110
rect 6020 4010 6100 4070
rect 6020 3970 6040 4010
rect 6080 3970 6100 4010
rect 6020 3910 6100 3970
rect 6020 3870 6040 3910
rect 6080 3870 6100 3910
rect 6020 3810 6100 3870
rect 6020 3770 6040 3810
rect 6080 3770 6100 3810
rect 6020 3740 6100 3770
rect 6220 4110 6300 4140
rect 6220 4070 6240 4110
rect 6280 4070 6300 4110
rect 6220 4010 6300 4070
rect 6220 3970 6240 4010
rect 6280 3970 6300 4010
rect 6220 3910 6300 3970
rect 6220 3870 6240 3910
rect 6280 3870 6300 3910
rect 6220 3810 6300 3870
rect 6220 3770 6240 3810
rect 6280 3770 6300 3810
rect 6220 3740 6300 3770
rect 6420 4110 6500 4140
rect 6420 4070 6440 4110
rect 6480 4070 6500 4110
rect 6420 4010 6500 4070
rect 6420 3970 6440 4010
rect 6480 3970 6500 4010
rect 6420 3910 6500 3970
rect 6420 3870 6440 3910
rect 6480 3870 6500 3910
rect 6420 3810 6500 3870
rect 6420 3770 6440 3810
rect 6480 3770 6500 3810
rect 6420 3740 6500 3770
rect 6620 4110 6700 4140
rect 6620 4070 6640 4110
rect 6680 4070 6700 4110
rect 6620 4010 6700 4070
rect 6620 3970 6640 4010
rect 6680 3970 6700 4010
rect 6620 3910 6700 3970
rect 6620 3870 6640 3910
rect 6680 3870 6700 3910
rect 6620 3810 6700 3870
rect 6620 3770 6640 3810
rect 6680 3770 6700 3810
rect 6620 3740 6700 3770
rect 6820 4110 6900 4140
rect 6820 4070 6840 4110
rect 6880 4070 6900 4110
rect 6820 4010 6900 4070
rect 6820 3970 6840 4010
rect 6880 3970 6900 4010
rect 6820 3910 6900 3970
rect 6820 3870 6840 3910
rect 6880 3870 6900 3910
rect 6820 3810 6900 3870
rect 6820 3770 6840 3810
rect 6880 3770 6900 3810
rect 6820 3740 6900 3770
rect 7020 4110 7100 4140
rect 7180 4110 7260 4140
rect 7020 4070 7040 4110
rect 7080 4070 7100 4110
rect 7180 4070 7200 4110
rect 7240 4070 7260 4110
rect 7020 4010 7100 4070
rect 7180 4010 7260 4070
rect 7020 3970 7040 4010
rect 7080 3970 7100 4010
rect 7180 3970 7200 4010
rect 7240 3970 7260 4010
rect 7020 3910 7100 3970
rect 7180 3910 7260 3970
rect 7020 3870 7040 3910
rect 7080 3870 7100 3910
rect 7180 3870 7200 3910
rect 7240 3870 7260 3910
rect 7020 3810 7100 3870
rect 7180 3810 7260 3870
rect 7020 3770 7040 3810
rect 7080 3770 7100 3810
rect 7180 3770 7200 3810
rect 7240 3770 7260 3810
rect 7020 3740 7100 3770
rect 7180 3740 7260 3770
rect 7380 4110 7460 4140
rect 7380 4070 7400 4110
rect 7440 4070 7460 4110
rect 7380 4010 7460 4070
rect 7380 3970 7400 4010
rect 7440 3970 7460 4010
rect 7380 3910 7460 3970
rect 7380 3870 7400 3910
rect 7440 3870 7460 3910
rect 7380 3810 7460 3870
rect 7380 3770 7400 3810
rect 7440 3770 7460 3810
rect 7380 3740 7460 3770
rect 7580 4110 7660 4140
rect 7580 4070 7600 4110
rect 7640 4070 7660 4110
rect 7580 4010 7660 4070
rect 7580 3970 7600 4010
rect 7640 3970 7660 4010
rect 7580 3910 7660 3970
rect 7580 3870 7600 3910
rect 7640 3870 7660 3910
rect 7580 3810 7660 3870
rect 7580 3770 7600 3810
rect 7640 3770 7660 3810
rect 7580 3740 7660 3770
rect 7780 4110 7860 4140
rect 7780 4070 7800 4110
rect 7840 4070 7860 4110
rect 7780 4010 7860 4070
rect 7780 3970 7800 4010
rect 7840 3970 7860 4010
rect 7780 3910 7860 3970
rect 7780 3870 7800 3910
rect 7840 3870 7860 3910
rect 7780 3810 7860 3870
rect 7780 3770 7800 3810
rect 7840 3770 7860 3810
rect 7780 3740 7860 3770
rect 7980 4110 8060 4140
rect 7980 4070 8000 4110
rect 8040 4070 8060 4110
rect 7980 4010 8060 4070
rect 7980 3970 8000 4010
rect 8040 3970 8060 4010
rect 7980 3910 8060 3970
rect 7980 3870 8000 3910
rect 8040 3870 8060 3910
rect 7980 3810 8060 3870
rect 7980 3770 8000 3810
rect 8040 3770 8060 3810
rect 7980 3740 8060 3770
rect 8180 4110 8260 4140
rect 8180 4070 8200 4110
rect 8240 4070 8260 4110
rect 8180 4010 8260 4070
rect 8180 3970 8200 4010
rect 8240 3970 8260 4010
rect 8180 3910 8260 3970
rect 8180 3870 8200 3910
rect 8240 3870 8260 3910
rect 8180 3810 8260 3870
rect 8180 3770 8200 3810
rect 8240 3770 8260 3810
rect 8180 3740 8260 3770
rect 8380 4110 8460 4140
rect 8380 4070 8400 4110
rect 8440 4070 8460 4110
rect 8380 4010 8460 4070
rect 8380 3970 8400 4010
rect 8440 3970 8460 4010
rect 8380 3910 8460 3970
rect 8380 3870 8400 3910
rect 8440 3870 8460 3910
rect 8380 3810 8460 3870
rect 8380 3770 8400 3810
rect 8440 3770 8460 3810
rect 8380 3740 8460 3770
rect 8750 4110 8830 4140
rect 8750 4070 8770 4110
rect 8810 4070 8830 4110
rect 8750 4010 8830 4070
rect 8750 3970 8770 4010
rect 8810 3970 8830 4010
rect 8750 3910 8830 3970
rect 8750 3870 8770 3910
rect 8810 3870 8830 3910
rect 8750 3810 8830 3870
rect 8750 3770 8770 3810
rect 8810 3770 8830 3810
rect 8750 3740 8830 3770
rect 8860 4110 8940 4140
rect 8860 4070 8880 4110
rect 8920 4070 8940 4110
rect 8860 4010 8940 4070
rect 8860 3970 8880 4010
rect 8920 3970 8940 4010
rect 8860 3910 8940 3970
rect 8860 3870 8880 3910
rect 8920 3870 8940 3910
rect 8860 3810 8940 3870
rect 8860 3770 8880 3810
rect 8920 3770 8940 3810
rect 8860 3740 8940 3770
rect 9000 4110 9080 4140
rect 9000 4070 9020 4110
rect 9060 4070 9080 4110
rect 9000 4010 9080 4070
rect 9000 3970 9020 4010
rect 9060 3970 9080 4010
rect 9000 3910 9080 3970
rect 9000 3870 9020 3910
rect 9060 3870 9080 3910
rect 9000 3810 9080 3870
rect 9000 3770 9020 3810
rect 9060 3770 9080 3810
rect 9000 3740 9080 3770
rect 9110 4110 9190 4140
rect 9110 4070 9130 4110
rect 9170 4070 9190 4110
rect 9110 4010 9190 4070
rect 9110 3970 9130 4010
rect 9170 3970 9190 4010
rect 9110 3910 9190 3970
rect 9110 3870 9130 3910
rect 9170 3870 9190 3910
rect 9110 3810 9190 3870
rect 9110 3770 9130 3810
rect 9170 3770 9190 3810
rect 9110 3740 9190 3770
rect 1680 958 2360 1010
rect 1680 924 1734 958
rect 1768 924 1824 958
rect 1858 924 1914 958
rect 1948 924 2004 958
rect 2038 924 2094 958
rect 2128 924 2184 958
rect 2218 924 2274 958
rect 2308 924 2360 958
rect 1680 868 2360 924
rect 1680 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2360 868
rect 1680 778 2360 834
rect 1680 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2360 778
rect 1680 688 2360 744
rect 1680 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2360 688
rect 1680 598 2360 654
rect 1680 564 1734 598
rect 1768 564 1824 598
rect 1858 564 1914 598
rect 1948 564 2004 598
rect 2038 564 2094 598
rect 2128 564 2184 598
rect 2218 564 2274 598
rect 2308 564 2360 598
rect 1680 508 2360 564
rect 1680 474 1734 508
rect 1768 474 1824 508
rect 1858 474 1914 508
rect 1948 474 2004 508
rect 2038 474 2094 508
rect 2128 474 2184 508
rect 2218 474 2274 508
rect 2308 474 2360 508
rect 1680 418 2360 474
rect 1680 384 1734 418
rect 1768 384 1824 418
rect 1858 384 1914 418
rect 1948 384 2004 418
rect 2038 384 2094 418
rect 2128 384 2184 418
rect 2218 384 2274 418
rect 2308 384 2360 418
rect 1680 330 2360 384
rect 3040 958 3720 1010
rect 3040 924 3094 958
rect 3128 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3720 958
rect 3040 868 3720 924
rect 3040 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3720 868
rect 3040 778 3720 834
rect 3040 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3720 778
rect 3040 688 3720 744
rect 3040 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3720 688
rect 3040 598 3720 654
rect 3040 564 3094 598
rect 3128 564 3184 598
rect 3218 564 3274 598
rect 3308 564 3364 598
rect 3398 564 3454 598
rect 3488 564 3544 598
rect 3578 564 3634 598
rect 3668 564 3720 598
rect 3040 508 3720 564
rect 3040 474 3094 508
rect 3128 474 3184 508
rect 3218 474 3274 508
rect 3308 474 3364 508
rect 3398 474 3454 508
rect 3488 474 3544 508
rect 3578 474 3634 508
rect 3668 474 3720 508
rect 3040 418 3720 474
rect 3040 384 3094 418
rect 3128 384 3184 418
rect 3218 384 3274 418
rect 3308 384 3364 418
rect 3398 384 3454 418
rect 3488 384 3544 418
rect 3578 384 3634 418
rect 3668 384 3720 418
rect 3040 330 3720 384
rect 4400 958 5080 1010
rect 4400 924 4454 958
rect 4488 924 4544 958
rect 4578 924 4634 958
rect 4668 924 4724 958
rect 4758 924 4814 958
rect 4848 924 4904 958
rect 4938 924 4994 958
rect 5028 924 5080 958
rect 4400 868 5080 924
rect 4400 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5080 868
rect 4400 778 5080 834
rect 4400 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5080 778
rect 4400 688 5080 744
rect 4400 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5080 688
rect 4400 598 5080 654
rect 4400 564 4454 598
rect 4488 564 4544 598
rect 4578 564 4634 598
rect 4668 564 4724 598
rect 4758 564 4814 598
rect 4848 564 4904 598
rect 4938 564 4994 598
rect 5028 564 5080 598
rect 4400 508 5080 564
rect 4400 474 4454 508
rect 4488 474 4544 508
rect 4578 474 4634 508
rect 4668 474 4724 508
rect 4758 474 4814 508
rect 4848 474 4904 508
rect 4938 474 4994 508
rect 5028 474 5080 508
rect 4400 418 5080 474
rect 4400 384 4454 418
rect 4488 384 4544 418
rect 4578 384 4634 418
rect 4668 384 4724 418
rect 4758 384 4814 418
rect 4848 384 4904 418
rect 4938 384 4994 418
rect 5028 384 5080 418
rect 4400 330 5080 384
rect 5760 958 6440 1010
rect 5760 924 5814 958
rect 5848 924 5904 958
rect 5938 924 5994 958
rect 6028 924 6084 958
rect 6118 924 6174 958
rect 6208 924 6264 958
rect 6298 924 6354 958
rect 6388 924 6440 958
rect 5760 868 6440 924
rect 5760 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6440 868
rect 5760 778 6440 834
rect 5760 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6440 778
rect 5760 688 6440 744
rect 5760 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6440 688
rect 5760 598 6440 654
rect 5760 564 5814 598
rect 5848 564 5904 598
rect 5938 564 5994 598
rect 6028 564 6084 598
rect 6118 564 6174 598
rect 6208 564 6264 598
rect 6298 564 6354 598
rect 6388 564 6440 598
rect 5760 508 6440 564
rect 5760 474 5814 508
rect 5848 474 5904 508
rect 5938 474 5994 508
rect 6028 474 6084 508
rect 6118 474 6174 508
rect 6208 474 6264 508
rect 6298 474 6354 508
rect 6388 474 6440 508
rect 5760 418 6440 474
rect 5760 384 5814 418
rect 5848 384 5904 418
rect 5938 384 5994 418
rect 6028 384 6084 418
rect 6118 384 6174 418
rect 6208 384 6264 418
rect 6298 384 6354 418
rect 6388 384 6440 418
rect 5760 330 6440 384
rect 7120 958 7800 1010
rect 7120 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7800 958
rect 7120 868 7800 924
rect 7120 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7800 868
rect 7120 778 7800 834
rect 7120 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7800 778
rect 7120 688 7800 744
rect 7120 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7800 688
rect 7120 598 7800 654
rect 7120 564 7174 598
rect 7208 564 7264 598
rect 7298 564 7354 598
rect 7388 564 7444 598
rect 7478 564 7534 598
rect 7568 564 7624 598
rect 7658 564 7714 598
rect 7748 564 7800 598
rect 7120 508 7800 564
rect 7120 474 7174 508
rect 7208 474 7264 508
rect 7298 474 7354 508
rect 7388 474 7444 508
rect 7478 474 7534 508
rect 7568 474 7624 508
rect 7658 474 7714 508
rect 7748 474 7800 508
rect 7120 418 7800 474
rect 7120 384 7174 418
rect 7208 384 7264 418
rect 7298 384 7354 418
rect 7388 384 7444 418
rect 7478 384 7534 418
rect 7568 384 7624 418
rect 7658 384 7714 418
rect 7748 384 7800 418
rect 7120 330 7800 384
rect 8480 958 9160 1010
rect 8480 924 8534 958
rect 8568 924 8624 958
rect 8658 924 8714 958
rect 8748 924 8804 958
rect 8838 924 8894 958
rect 8928 924 8984 958
rect 9018 924 9074 958
rect 9108 924 9160 958
rect 8480 868 9160 924
rect 8480 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9160 868
rect 8480 778 9160 834
rect 8480 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9160 778
rect 8480 688 9160 744
rect 8480 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9160 688
rect 8480 598 9160 654
rect 8480 564 8534 598
rect 8568 564 8624 598
rect 8658 564 8714 598
rect 8748 564 8804 598
rect 8838 564 8894 598
rect 8928 564 8984 598
rect 9018 564 9074 598
rect 9108 564 9160 598
rect 8480 508 9160 564
rect 8480 474 8534 508
rect 8568 474 8624 508
rect 8658 474 8714 508
rect 8748 474 8804 508
rect 8838 474 8894 508
rect 8928 474 8984 508
rect 9018 474 9074 508
rect 9108 474 9160 508
rect 8480 418 9160 474
rect 8480 384 8534 418
rect 8568 384 8624 418
rect 8658 384 8714 418
rect 8748 384 8804 418
rect 8838 384 8894 418
rect 8928 384 8984 418
rect 9018 384 9074 418
rect 9108 384 9160 418
rect 8480 330 9160 384
<< ndiffc >>
rect 5160 3260 5200 3300
rect 5160 3160 5200 3200
rect 5360 3260 5400 3300
rect 5360 3160 5400 3200
rect 5560 3260 5600 3300
rect 5560 3160 5600 3200
rect 5760 3260 5800 3300
rect 5760 3160 5800 3200
rect 5960 3260 6000 3300
rect 5960 3160 6000 3200
rect 6160 3260 6200 3300
rect 6160 3160 6200 3200
rect 6360 3260 6400 3300
rect 6520 3260 6560 3300
rect 6360 3160 6400 3200
rect 6520 3160 6560 3200
rect 6720 3260 6760 3300
rect 6720 3160 6760 3200
rect 6920 3260 6960 3300
rect 6920 3160 6960 3200
rect 7120 3260 7160 3300
rect 7120 3160 7160 3200
rect 7320 3260 7360 3300
rect 7320 3160 7360 3200
rect 7520 3260 7560 3300
rect 7520 3160 7560 3200
rect 7720 3260 7760 3300
rect 7720 3160 7760 3200
rect 4680 2710 4720 2750
rect 4680 2610 4720 2650
rect 4680 2510 4720 2550
rect 4680 2410 4720 2450
rect 4680 2310 4720 2350
rect 4680 2210 4720 2250
rect 4680 2110 4720 2150
rect 4680 2010 4720 2050
rect 5560 2710 5600 2750
rect 5560 2610 5600 2650
rect 5560 2510 5600 2550
rect 5560 2410 5600 2450
rect 5560 2310 5600 2350
rect 5560 2210 5600 2250
rect 5560 2110 5600 2150
rect 5560 2010 5600 2050
rect 6440 2710 6480 2750
rect 6440 2610 6480 2650
rect 6440 2510 6480 2550
rect 6440 2410 6480 2450
rect 6440 2310 6480 2350
rect 6440 2210 6480 2250
rect 6440 2110 6480 2150
rect 6440 2010 6480 2050
rect 7320 2710 7360 2750
rect 7320 2610 7360 2650
rect 7320 2510 7360 2550
rect 7320 2410 7360 2450
rect 7320 2310 7360 2350
rect 7320 2210 7360 2250
rect 7320 2110 7360 2150
rect 7320 2010 7360 2050
rect 8200 2710 8240 2750
rect 8200 2610 8240 2650
rect 8200 2510 8240 2550
rect 8200 2410 8240 2450
rect 8200 2310 8240 2350
rect 8200 2210 8240 2250
rect 8200 2110 8240 2150
rect 8200 2010 8240 2050
rect 5380 1640 5420 1680
rect 5380 1540 5420 1580
rect 7460 1640 7500 1680
rect 7460 1540 7500 1580
<< pdiffc >>
rect 4440 5380 4480 5420
rect 4440 5280 4480 5320
rect 4440 5180 4480 5220
rect 4440 5080 4480 5120
rect 4440 4980 4480 5020
rect 4440 4880 4480 4920
rect 4440 4780 4480 4820
rect 4440 4680 4480 4720
rect 4640 5380 4680 5420
rect 4640 5280 4680 5320
rect 4640 5180 4680 5220
rect 4640 5080 4680 5120
rect 4640 4980 4680 5020
rect 4640 4880 4680 4920
rect 4640 4780 4680 4820
rect 4640 4680 4680 4720
rect 4840 5380 4880 5420
rect 4840 5280 4880 5320
rect 4840 5180 4880 5220
rect 4840 5080 4880 5120
rect 4840 4980 4880 5020
rect 4840 4880 4880 4920
rect 4840 4780 4880 4820
rect 4840 4680 4880 4720
rect 5040 5380 5080 5420
rect 5040 5280 5080 5320
rect 5040 5180 5080 5220
rect 5040 5080 5080 5120
rect 5040 4980 5080 5020
rect 5040 4880 5080 4920
rect 5040 4780 5080 4820
rect 5040 4680 5080 4720
rect 5240 5380 5280 5420
rect 5240 5280 5280 5320
rect 5240 5180 5280 5220
rect 5240 5080 5280 5120
rect 5240 4980 5280 5020
rect 5240 4880 5280 4920
rect 5240 4780 5280 4820
rect 5240 4680 5280 4720
rect 5440 5380 5480 5420
rect 5440 5280 5480 5320
rect 5440 5180 5480 5220
rect 5440 5080 5480 5120
rect 5440 4980 5480 5020
rect 5440 4880 5480 4920
rect 5440 4780 5480 4820
rect 5440 4680 5480 4720
rect 5640 5380 5680 5420
rect 5640 5280 5680 5320
rect 5640 5180 5680 5220
rect 5640 5080 5680 5120
rect 5640 4980 5680 5020
rect 5640 4880 5680 4920
rect 5640 4780 5680 4820
rect 5640 4680 5680 4720
rect 5840 5380 5880 5420
rect 5840 5280 5880 5320
rect 5840 5180 5880 5220
rect 5840 5080 5880 5120
rect 5840 4980 5880 5020
rect 5840 4880 5880 4920
rect 5840 4780 5880 4820
rect 5840 4680 5880 4720
rect 6040 5380 6080 5420
rect 6040 5280 6080 5320
rect 6040 5180 6080 5220
rect 6040 5080 6080 5120
rect 6040 4980 6080 5020
rect 6040 4880 6080 4920
rect 6040 4780 6080 4820
rect 6040 4680 6080 4720
rect 6240 5380 6280 5420
rect 6240 5280 6280 5320
rect 6240 5180 6280 5220
rect 6240 5080 6280 5120
rect 6240 4980 6280 5020
rect 6240 4880 6280 4920
rect 6240 4780 6280 4820
rect 6240 4680 6280 4720
rect 6440 5380 6480 5420
rect 6440 5280 6480 5320
rect 6440 5180 6480 5220
rect 6440 5080 6480 5120
rect 6440 4980 6480 5020
rect 6440 4880 6480 4920
rect 6440 4780 6480 4820
rect 6440 4680 6480 4720
rect 6640 5380 6680 5420
rect 6640 5280 6680 5320
rect 6640 5180 6680 5220
rect 6640 5080 6680 5120
rect 6640 4980 6680 5020
rect 6640 4880 6680 4920
rect 6640 4780 6680 4820
rect 6640 4680 6680 4720
rect 6840 5380 6880 5420
rect 6840 5280 6880 5320
rect 6840 5180 6880 5220
rect 6840 5080 6880 5120
rect 6840 4980 6880 5020
rect 6840 4880 6880 4920
rect 6840 4780 6880 4820
rect 6840 4680 6880 4720
rect 7040 5380 7080 5420
rect 7040 5280 7080 5320
rect 7040 5180 7080 5220
rect 7040 5080 7080 5120
rect 7040 4980 7080 5020
rect 7040 4880 7080 4920
rect 7040 4780 7080 4820
rect 7040 4680 7080 4720
rect 7240 5380 7280 5420
rect 7240 5280 7280 5320
rect 7240 5180 7280 5220
rect 7240 5080 7280 5120
rect 7240 4980 7280 5020
rect 7240 4880 7280 4920
rect 7240 4780 7280 4820
rect 7240 4680 7280 4720
rect 7440 5380 7480 5420
rect 7440 5280 7480 5320
rect 7440 5180 7480 5220
rect 7440 5080 7480 5120
rect 7440 4980 7480 5020
rect 7440 4880 7480 4920
rect 7440 4780 7480 4820
rect 7440 4680 7480 4720
rect 7640 5380 7680 5420
rect 7640 5280 7680 5320
rect 7640 5180 7680 5220
rect 7640 5080 7680 5120
rect 7640 4980 7680 5020
rect 7640 4880 7680 4920
rect 7640 4780 7680 4820
rect 7640 4680 7680 4720
rect 7840 5380 7880 5420
rect 7840 5280 7880 5320
rect 7840 5180 7880 5220
rect 7840 5080 7880 5120
rect 7840 4980 7880 5020
rect 7840 4880 7880 4920
rect 7840 4780 7880 4820
rect 7840 4680 7880 4720
rect 8040 5380 8080 5420
rect 8040 5280 8080 5320
rect 8040 5180 8080 5220
rect 8040 5080 8080 5120
rect 8040 4980 8080 5020
rect 8040 4880 8080 4920
rect 8040 4780 8080 4820
rect 8040 4680 8080 4720
rect 8240 5380 8280 5420
rect 8240 5280 8280 5320
rect 8240 5180 8280 5220
rect 8240 5080 8280 5120
rect 8240 4980 8280 5020
rect 8240 4880 8280 4920
rect 8240 4780 8280 4820
rect 8240 4680 8280 4720
rect 8440 5380 8480 5420
rect 8440 5280 8480 5320
rect 8440 5180 8480 5220
rect 8440 5080 8480 5120
rect 8440 4980 8480 5020
rect 8440 4880 8480 4920
rect 8440 4780 8480 4820
rect 8440 4680 8480 4720
rect 4480 4070 4520 4110
rect 4480 3970 4520 4010
rect 4480 3870 4520 3910
rect 4480 3770 4520 3810
rect 4680 4070 4720 4110
rect 4680 3970 4720 4010
rect 4680 3870 4720 3910
rect 4680 3770 4720 3810
rect 4880 4070 4920 4110
rect 4880 3970 4920 4010
rect 4880 3870 4920 3910
rect 4880 3770 4920 3810
rect 5080 4070 5120 4110
rect 5080 3970 5120 4010
rect 5080 3870 5120 3910
rect 5080 3770 5120 3810
rect 5280 4070 5320 4110
rect 5280 3970 5320 4010
rect 5280 3870 5320 3910
rect 5280 3770 5320 3810
rect 5480 4070 5520 4110
rect 5480 3970 5520 4010
rect 5480 3870 5520 3910
rect 5480 3770 5520 3810
rect 5680 4070 5720 4110
rect 5840 4070 5880 4110
rect 5680 3970 5720 4010
rect 5840 3970 5880 4010
rect 5680 3870 5720 3910
rect 5840 3870 5880 3910
rect 5680 3770 5720 3810
rect 5840 3770 5880 3810
rect 6040 4070 6080 4110
rect 6040 3970 6080 4010
rect 6040 3870 6080 3910
rect 6040 3770 6080 3810
rect 6240 4070 6280 4110
rect 6240 3970 6280 4010
rect 6240 3870 6280 3910
rect 6240 3770 6280 3810
rect 6440 4070 6480 4110
rect 6440 3970 6480 4010
rect 6440 3870 6480 3910
rect 6440 3770 6480 3810
rect 6640 4070 6680 4110
rect 6640 3970 6680 4010
rect 6640 3870 6680 3910
rect 6640 3770 6680 3810
rect 6840 4070 6880 4110
rect 6840 3970 6880 4010
rect 6840 3870 6880 3910
rect 6840 3770 6880 3810
rect 7040 4070 7080 4110
rect 7200 4070 7240 4110
rect 7040 3970 7080 4010
rect 7200 3970 7240 4010
rect 7040 3870 7080 3910
rect 7200 3870 7240 3910
rect 7040 3770 7080 3810
rect 7200 3770 7240 3810
rect 7400 4070 7440 4110
rect 7400 3970 7440 4010
rect 7400 3870 7440 3910
rect 7400 3770 7440 3810
rect 7600 4070 7640 4110
rect 7600 3970 7640 4010
rect 7600 3870 7640 3910
rect 7600 3770 7640 3810
rect 7800 4070 7840 4110
rect 7800 3970 7840 4010
rect 7800 3870 7840 3910
rect 7800 3770 7840 3810
rect 8000 4070 8040 4110
rect 8000 3970 8040 4010
rect 8000 3870 8040 3910
rect 8000 3770 8040 3810
rect 8200 4070 8240 4110
rect 8200 3970 8240 4010
rect 8200 3870 8240 3910
rect 8200 3770 8240 3810
rect 8400 4070 8440 4110
rect 8400 3970 8440 4010
rect 8400 3870 8440 3910
rect 8400 3770 8440 3810
rect 8770 4070 8810 4110
rect 8770 3970 8810 4010
rect 8770 3870 8810 3910
rect 8770 3770 8810 3810
rect 8880 4070 8920 4110
rect 8880 3970 8920 4010
rect 8880 3870 8920 3910
rect 8880 3770 8920 3810
rect 9020 4070 9060 4110
rect 9020 3970 9060 4010
rect 9020 3870 9060 3910
rect 9020 3770 9060 3810
rect 9130 4070 9170 4110
rect 9130 3970 9170 4010
rect 9130 3870 9170 3910
rect 9130 3770 9170 3810
rect 1734 924 1768 958
rect 1824 924 1858 958
rect 1914 924 1948 958
rect 2004 924 2038 958
rect 2094 924 2128 958
rect 2184 924 2218 958
rect 2274 924 2308 958
rect 1734 834 1768 868
rect 1824 834 1858 868
rect 1914 834 1948 868
rect 2004 834 2038 868
rect 2094 834 2128 868
rect 2184 834 2218 868
rect 2274 834 2308 868
rect 1734 744 1768 778
rect 1824 744 1858 778
rect 1914 744 1948 778
rect 2004 744 2038 778
rect 2094 744 2128 778
rect 2184 744 2218 778
rect 2274 744 2308 778
rect 1734 654 1768 688
rect 1824 654 1858 688
rect 1914 654 1948 688
rect 2004 654 2038 688
rect 2094 654 2128 688
rect 2184 654 2218 688
rect 2274 654 2308 688
rect 1734 564 1768 598
rect 1824 564 1858 598
rect 1914 564 1948 598
rect 2004 564 2038 598
rect 2094 564 2128 598
rect 2184 564 2218 598
rect 2274 564 2308 598
rect 1734 474 1768 508
rect 1824 474 1858 508
rect 1914 474 1948 508
rect 2004 474 2038 508
rect 2094 474 2128 508
rect 2184 474 2218 508
rect 2274 474 2308 508
rect 1734 384 1768 418
rect 1824 384 1858 418
rect 1914 384 1948 418
rect 2004 384 2038 418
rect 2094 384 2128 418
rect 2184 384 2218 418
rect 2274 384 2308 418
rect 3094 924 3128 958
rect 3184 924 3218 958
rect 3274 924 3308 958
rect 3364 924 3398 958
rect 3454 924 3488 958
rect 3544 924 3578 958
rect 3634 924 3668 958
rect 3094 834 3128 868
rect 3184 834 3218 868
rect 3274 834 3308 868
rect 3364 834 3398 868
rect 3454 834 3488 868
rect 3544 834 3578 868
rect 3634 834 3668 868
rect 3094 744 3128 778
rect 3184 744 3218 778
rect 3274 744 3308 778
rect 3364 744 3398 778
rect 3454 744 3488 778
rect 3544 744 3578 778
rect 3634 744 3668 778
rect 3094 654 3128 688
rect 3184 654 3218 688
rect 3274 654 3308 688
rect 3364 654 3398 688
rect 3454 654 3488 688
rect 3544 654 3578 688
rect 3634 654 3668 688
rect 3094 564 3128 598
rect 3184 564 3218 598
rect 3274 564 3308 598
rect 3364 564 3398 598
rect 3454 564 3488 598
rect 3544 564 3578 598
rect 3634 564 3668 598
rect 3094 474 3128 508
rect 3184 474 3218 508
rect 3274 474 3308 508
rect 3364 474 3398 508
rect 3454 474 3488 508
rect 3544 474 3578 508
rect 3634 474 3668 508
rect 3094 384 3128 418
rect 3184 384 3218 418
rect 3274 384 3308 418
rect 3364 384 3398 418
rect 3454 384 3488 418
rect 3544 384 3578 418
rect 3634 384 3668 418
rect 4454 924 4488 958
rect 4544 924 4578 958
rect 4634 924 4668 958
rect 4724 924 4758 958
rect 4814 924 4848 958
rect 4904 924 4938 958
rect 4994 924 5028 958
rect 4454 834 4488 868
rect 4544 834 4578 868
rect 4634 834 4668 868
rect 4724 834 4758 868
rect 4814 834 4848 868
rect 4904 834 4938 868
rect 4994 834 5028 868
rect 4454 744 4488 778
rect 4544 744 4578 778
rect 4634 744 4668 778
rect 4724 744 4758 778
rect 4814 744 4848 778
rect 4904 744 4938 778
rect 4994 744 5028 778
rect 4454 654 4488 688
rect 4544 654 4578 688
rect 4634 654 4668 688
rect 4724 654 4758 688
rect 4814 654 4848 688
rect 4904 654 4938 688
rect 4994 654 5028 688
rect 4454 564 4488 598
rect 4544 564 4578 598
rect 4634 564 4668 598
rect 4724 564 4758 598
rect 4814 564 4848 598
rect 4904 564 4938 598
rect 4994 564 5028 598
rect 4454 474 4488 508
rect 4544 474 4578 508
rect 4634 474 4668 508
rect 4724 474 4758 508
rect 4814 474 4848 508
rect 4904 474 4938 508
rect 4994 474 5028 508
rect 4454 384 4488 418
rect 4544 384 4578 418
rect 4634 384 4668 418
rect 4724 384 4758 418
rect 4814 384 4848 418
rect 4904 384 4938 418
rect 4994 384 5028 418
rect 5814 924 5848 958
rect 5904 924 5938 958
rect 5994 924 6028 958
rect 6084 924 6118 958
rect 6174 924 6208 958
rect 6264 924 6298 958
rect 6354 924 6388 958
rect 5814 834 5848 868
rect 5904 834 5938 868
rect 5994 834 6028 868
rect 6084 834 6118 868
rect 6174 834 6208 868
rect 6264 834 6298 868
rect 6354 834 6388 868
rect 5814 744 5848 778
rect 5904 744 5938 778
rect 5994 744 6028 778
rect 6084 744 6118 778
rect 6174 744 6208 778
rect 6264 744 6298 778
rect 6354 744 6388 778
rect 5814 654 5848 688
rect 5904 654 5938 688
rect 5994 654 6028 688
rect 6084 654 6118 688
rect 6174 654 6208 688
rect 6264 654 6298 688
rect 6354 654 6388 688
rect 5814 564 5848 598
rect 5904 564 5938 598
rect 5994 564 6028 598
rect 6084 564 6118 598
rect 6174 564 6208 598
rect 6264 564 6298 598
rect 6354 564 6388 598
rect 5814 474 5848 508
rect 5904 474 5938 508
rect 5994 474 6028 508
rect 6084 474 6118 508
rect 6174 474 6208 508
rect 6264 474 6298 508
rect 6354 474 6388 508
rect 5814 384 5848 418
rect 5904 384 5938 418
rect 5994 384 6028 418
rect 6084 384 6118 418
rect 6174 384 6208 418
rect 6264 384 6298 418
rect 6354 384 6388 418
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7714 924 7748 958
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7714 834 7748 868
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7714 744 7748 778
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 7714 654 7748 688
rect 7174 564 7208 598
rect 7264 564 7298 598
rect 7354 564 7388 598
rect 7444 564 7478 598
rect 7534 564 7568 598
rect 7624 564 7658 598
rect 7714 564 7748 598
rect 7174 474 7208 508
rect 7264 474 7298 508
rect 7354 474 7388 508
rect 7444 474 7478 508
rect 7534 474 7568 508
rect 7624 474 7658 508
rect 7714 474 7748 508
rect 7174 384 7208 418
rect 7264 384 7298 418
rect 7354 384 7388 418
rect 7444 384 7478 418
rect 7534 384 7568 418
rect 7624 384 7658 418
rect 7714 384 7748 418
rect 8534 924 8568 958
rect 8624 924 8658 958
rect 8714 924 8748 958
rect 8804 924 8838 958
rect 8894 924 8928 958
rect 8984 924 9018 958
rect 9074 924 9108 958
rect 8534 834 8568 868
rect 8624 834 8658 868
rect 8714 834 8748 868
rect 8804 834 8838 868
rect 8894 834 8928 868
rect 8984 834 9018 868
rect 9074 834 9108 868
rect 8534 744 8568 778
rect 8624 744 8658 778
rect 8714 744 8748 778
rect 8804 744 8838 778
rect 8894 744 8928 778
rect 8984 744 9018 778
rect 9074 744 9108 778
rect 8534 654 8568 688
rect 8624 654 8658 688
rect 8714 654 8748 688
rect 8804 654 8838 688
rect 8894 654 8928 688
rect 8984 654 9018 688
rect 9074 654 9108 688
rect 8534 564 8568 598
rect 8624 564 8658 598
rect 8714 564 8748 598
rect 8804 564 8838 598
rect 8894 564 8928 598
rect 8984 564 9018 598
rect 9074 564 9108 598
rect 8534 474 8568 508
rect 8624 474 8658 508
rect 8714 474 8748 508
rect 8804 474 8838 508
rect 8894 474 8928 508
rect 8984 474 9018 508
rect 9074 474 9108 508
rect 8534 384 8568 418
rect 8624 384 8658 418
rect 8714 384 8748 418
rect 8804 384 8838 418
rect 8894 384 8928 418
rect 8984 384 9018 418
rect 9074 384 9108 418
<< psubdiff >>
rect 5060 3300 5140 3330
rect 5060 3260 5080 3300
rect 5120 3260 5140 3300
rect 5060 3200 5140 3260
rect 5060 3160 5080 3200
rect 5120 3160 5140 3200
rect 5060 3130 5140 3160
rect 6420 3300 6500 3330
rect 6420 3260 6440 3300
rect 6480 3260 6500 3300
rect 6420 3200 6500 3260
rect 6420 3160 6440 3200
rect 6480 3160 6500 3200
rect 6420 3130 6500 3160
rect 7780 3300 7860 3330
rect 7780 3260 7800 3300
rect 7840 3260 7860 3300
rect 7780 3200 7860 3260
rect 7780 3160 7800 3200
rect 7840 3160 7860 3200
rect 7780 3130 7860 3160
rect 4580 2750 4660 2780
rect 4580 2710 4600 2750
rect 4640 2710 4660 2750
rect 4580 2650 4660 2710
rect 4580 2610 4600 2650
rect 4640 2610 4660 2650
rect 4580 2550 4660 2610
rect 4580 2510 4600 2550
rect 4640 2510 4660 2550
rect 4580 2450 4660 2510
rect 4580 2410 4600 2450
rect 4640 2410 4660 2450
rect 4580 2350 4660 2410
rect 4580 2310 4600 2350
rect 4640 2310 4660 2350
rect 4580 2250 4660 2310
rect 4580 2210 4600 2250
rect 4640 2210 4660 2250
rect 4580 2150 4660 2210
rect 4580 2110 4600 2150
rect 4640 2110 4660 2150
rect 4580 2050 4660 2110
rect 4580 2010 4600 2050
rect 4640 2010 4660 2050
rect 4580 1980 4660 2010
rect 8260 2750 8340 2780
rect 8260 2710 8280 2750
rect 8320 2710 8340 2750
rect 8260 2650 8340 2710
rect 8260 2610 8280 2650
rect 8320 2610 8340 2650
rect 8260 2550 8340 2610
rect 8260 2510 8280 2550
rect 8320 2510 8340 2550
rect 8260 2450 8340 2510
rect 8260 2410 8280 2450
rect 8320 2410 8340 2450
rect 8260 2350 8340 2410
rect 8260 2310 8280 2350
rect 8320 2310 8340 2350
rect 8260 2250 8340 2310
rect 8260 2210 8280 2250
rect 8320 2210 8340 2250
rect 8260 2150 8340 2210
rect 8260 2110 8280 2150
rect 8320 2110 8340 2150
rect 8260 2050 8340 2110
rect 8260 2010 8280 2050
rect 8320 2010 8340 2050
rect 8260 1980 8340 2010
rect 7520 1680 7600 1710
rect 7520 1640 7540 1680
rect 7580 1640 7600 1680
rect 7520 1580 7600 1640
rect 7520 1540 7540 1580
rect 7580 1540 7600 1580
rect 7520 1510 7600 1540
rect 1376 1279 2664 1314
rect 1376 1256 1506 1279
rect 1376 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2664 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2664 1256
rect 1376 1213 2664 1222
rect 1376 1166 1477 1213
rect 1376 1132 1410 1166
rect 1444 1132 1477 1166
rect 2563 1166 2664 1213
rect 1376 1076 1477 1132
rect 1376 1042 1410 1076
rect 1444 1042 1477 1076
rect 1376 986 1477 1042
rect 1376 952 1410 986
rect 1444 952 1477 986
rect 1376 896 1477 952
rect 1376 862 1410 896
rect 1444 862 1477 896
rect 1376 806 1477 862
rect 1376 772 1410 806
rect 1444 772 1477 806
rect 1376 716 1477 772
rect 1376 682 1410 716
rect 1444 682 1477 716
rect 1376 626 1477 682
rect 1376 592 1410 626
rect 1444 592 1477 626
rect 1376 536 1477 592
rect 1376 502 1410 536
rect 1444 502 1477 536
rect 1376 446 1477 502
rect 1376 412 1410 446
rect 1444 412 1477 446
rect 1376 356 1477 412
rect 1376 322 1410 356
rect 1444 322 1477 356
rect 1376 266 1477 322
rect 1376 232 1410 266
rect 1444 232 1477 266
rect 1376 176 1477 232
rect 2563 1132 2597 1166
rect 2631 1132 2664 1166
rect 2563 1076 2664 1132
rect 2563 1042 2597 1076
rect 2631 1042 2664 1076
rect 2563 986 2664 1042
rect 2563 952 2597 986
rect 2631 952 2664 986
rect 2563 896 2664 952
rect 2563 862 2597 896
rect 2631 862 2664 896
rect 2563 806 2664 862
rect 2563 772 2597 806
rect 2631 772 2664 806
rect 2563 716 2664 772
rect 2563 682 2597 716
rect 2631 682 2664 716
rect 2563 626 2664 682
rect 2563 592 2597 626
rect 2631 592 2664 626
rect 2563 536 2664 592
rect 2563 502 2597 536
rect 2631 502 2664 536
rect 2563 446 2664 502
rect 2563 412 2597 446
rect 2631 412 2664 446
rect 2563 356 2664 412
rect 2563 322 2597 356
rect 2631 322 2664 356
rect 2563 266 2664 322
rect 2563 232 2597 266
rect 2631 232 2664 266
rect 1376 142 1410 176
rect 1444 142 1477 176
rect 1376 127 1477 142
rect 2563 176 2664 232
rect 2563 142 2597 176
rect 2631 142 2664 176
rect 2563 127 2664 142
rect 1376 92 2664 127
rect 40 50 80 90
rect 1376 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2664 92
rect 1376 26 2664 58
rect 2736 1279 4024 1314
rect 2736 1256 2866 1279
rect 2736 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4024 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4024 1256
rect 2736 1213 4024 1222
rect 2736 1166 2837 1213
rect 2736 1132 2770 1166
rect 2804 1132 2837 1166
rect 3923 1166 4024 1213
rect 2736 1076 2837 1132
rect 2736 1042 2770 1076
rect 2804 1042 2837 1076
rect 2736 986 2837 1042
rect 2736 952 2770 986
rect 2804 952 2837 986
rect 2736 896 2837 952
rect 2736 862 2770 896
rect 2804 862 2837 896
rect 2736 806 2837 862
rect 2736 772 2770 806
rect 2804 772 2837 806
rect 2736 716 2837 772
rect 2736 682 2770 716
rect 2804 682 2837 716
rect 2736 626 2837 682
rect 2736 592 2770 626
rect 2804 592 2837 626
rect 2736 536 2837 592
rect 2736 502 2770 536
rect 2804 502 2837 536
rect 2736 446 2837 502
rect 2736 412 2770 446
rect 2804 412 2837 446
rect 2736 356 2837 412
rect 2736 322 2770 356
rect 2804 322 2837 356
rect 2736 266 2837 322
rect 2736 232 2770 266
rect 2804 232 2837 266
rect 2736 176 2837 232
rect 3923 1132 3957 1166
rect 3991 1132 4024 1166
rect 3923 1076 4024 1132
rect 3923 1042 3957 1076
rect 3991 1042 4024 1076
rect 3923 986 4024 1042
rect 3923 952 3957 986
rect 3991 952 4024 986
rect 3923 896 4024 952
rect 3923 862 3957 896
rect 3991 862 4024 896
rect 3923 806 4024 862
rect 3923 772 3957 806
rect 3991 772 4024 806
rect 3923 716 4024 772
rect 3923 682 3957 716
rect 3991 682 4024 716
rect 3923 626 4024 682
rect 3923 592 3957 626
rect 3991 592 4024 626
rect 3923 536 4024 592
rect 3923 502 3957 536
rect 3991 502 4024 536
rect 3923 446 4024 502
rect 3923 412 3957 446
rect 3991 412 4024 446
rect 3923 356 4024 412
rect 3923 322 3957 356
rect 3991 322 4024 356
rect 3923 266 4024 322
rect 3923 232 3957 266
rect 3991 232 4024 266
rect 2736 142 2770 176
rect 2804 142 2837 176
rect 2736 127 2837 142
rect 3923 176 4024 232
rect 3923 142 3957 176
rect 3991 142 4024 176
rect 3923 127 4024 142
rect 2736 92 4024 127
rect 2736 58 2866 92
rect 2900 58 2956 92
rect 2990 58 3046 92
rect 3080 58 3136 92
rect 3170 58 3226 92
rect 3260 58 3316 92
rect 3350 58 3406 92
rect 3440 58 3496 92
rect 3530 58 3586 92
rect 3620 58 3676 92
rect 3710 58 3766 92
rect 3800 58 3856 92
rect 3890 58 4024 92
rect 2736 26 4024 58
rect 4096 1279 5384 1314
rect 4096 1256 4226 1279
rect 4096 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5384 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5384 1256
rect 4096 1213 5384 1222
rect 4096 1166 4197 1213
rect 4096 1132 4130 1166
rect 4164 1132 4197 1166
rect 5283 1166 5384 1213
rect 4096 1076 4197 1132
rect 4096 1042 4130 1076
rect 4164 1042 4197 1076
rect 4096 986 4197 1042
rect 4096 952 4130 986
rect 4164 952 4197 986
rect 4096 896 4197 952
rect 4096 862 4130 896
rect 4164 862 4197 896
rect 4096 806 4197 862
rect 4096 772 4130 806
rect 4164 772 4197 806
rect 4096 716 4197 772
rect 4096 682 4130 716
rect 4164 682 4197 716
rect 4096 626 4197 682
rect 4096 592 4130 626
rect 4164 592 4197 626
rect 4096 536 4197 592
rect 4096 502 4130 536
rect 4164 502 4197 536
rect 4096 446 4197 502
rect 4096 412 4130 446
rect 4164 412 4197 446
rect 4096 356 4197 412
rect 4096 322 4130 356
rect 4164 322 4197 356
rect 4096 266 4197 322
rect 4096 232 4130 266
rect 4164 232 4197 266
rect 4096 176 4197 232
rect 5283 1132 5317 1166
rect 5351 1132 5384 1166
rect 5283 1076 5384 1132
rect 5283 1042 5317 1076
rect 5351 1042 5384 1076
rect 5283 986 5384 1042
rect 5283 952 5317 986
rect 5351 952 5384 986
rect 5283 896 5384 952
rect 5283 862 5317 896
rect 5351 862 5384 896
rect 5283 806 5384 862
rect 5283 772 5317 806
rect 5351 772 5384 806
rect 5283 716 5384 772
rect 5283 682 5317 716
rect 5351 682 5384 716
rect 5283 626 5384 682
rect 5283 592 5317 626
rect 5351 592 5384 626
rect 5283 536 5384 592
rect 5283 502 5317 536
rect 5351 502 5384 536
rect 5283 446 5384 502
rect 5283 412 5317 446
rect 5351 412 5384 446
rect 5283 356 5384 412
rect 5283 322 5317 356
rect 5351 322 5384 356
rect 5283 266 5384 322
rect 5283 232 5317 266
rect 5351 232 5384 266
rect 4096 142 4130 176
rect 4164 142 4197 176
rect 4096 127 4197 142
rect 5283 176 5384 232
rect 5283 142 5317 176
rect 5351 142 5384 176
rect 5283 127 5384 142
rect 4096 92 5384 127
rect 4096 58 4226 92
rect 4260 58 4316 92
rect 4350 58 4406 92
rect 4440 58 4496 92
rect 4530 58 4586 92
rect 4620 58 4676 92
rect 4710 58 4766 92
rect 4800 58 4856 92
rect 4890 58 4946 92
rect 4980 58 5036 92
rect 5070 58 5126 92
rect 5160 58 5216 92
rect 5250 58 5384 92
rect 4096 26 5384 58
rect 5456 1279 6744 1314
rect 5456 1256 5586 1279
rect 5456 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6744 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6744 1256
rect 5456 1213 6744 1222
rect 5456 1166 5557 1213
rect 5456 1132 5490 1166
rect 5524 1132 5557 1166
rect 6643 1166 6744 1213
rect 5456 1076 5557 1132
rect 5456 1042 5490 1076
rect 5524 1042 5557 1076
rect 5456 986 5557 1042
rect 5456 952 5490 986
rect 5524 952 5557 986
rect 5456 896 5557 952
rect 5456 862 5490 896
rect 5524 862 5557 896
rect 5456 806 5557 862
rect 5456 772 5490 806
rect 5524 772 5557 806
rect 5456 716 5557 772
rect 5456 682 5490 716
rect 5524 682 5557 716
rect 5456 626 5557 682
rect 5456 592 5490 626
rect 5524 592 5557 626
rect 5456 536 5557 592
rect 5456 502 5490 536
rect 5524 502 5557 536
rect 5456 446 5557 502
rect 5456 412 5490 446
rect 5524 412 5557 446
rect 5456 356 5557 412
rect 5456 322 5490 356
rect 5524 322 5557 356
rect 5456 266 5557 322
rect 5456 232 5490 266
rect 5524 232 5557 266
rect 5456 176 5557 232
rect 6643 1132 6677 1166
rect 6711 1132 6744 1166
rect 6643 1076 6744 1132
rect 6643 1042 6677 1076
rect 6711 1042 6744 1076
rect 6643 986 6744 1042
rect 6643 952 6677 986
rect 6711 952 6744 986
rect 6643 896 6744 952
rect 6643 862 6677 896
rect 6711 862 6744 896
rect 6643 806 6744 862
rect 6643 772 6677 806
rect 6711 772 6744 806
rect 6643 716 6744 772
rect 6643 682 6677 716
rect 6711 682 6744 716
rect 6643 626 6744 682
rect 6643 592 6677 626
rect 6711 592 6744 626
rect 6643 536 6744 592
rect 6643 502 6677 536
rect 6711 502 6744 536
rect 6643 446 6744 502
rect 6643 412 6677 446
rect 6711 412 6744 446
rect 6643 356 6744 412
rect 6643 322 6677 356
rect 6711 322 6744 356
rect 6643 266 6744 322
rect 6643 232 6677 266
rect 6711 232 6744 266
rect 5456 142 5490 176
rect 5524 142 5557 176
rect 5456 127 5557 142
rect 6643 176 6744 232
rect 6643 142 6677 176
rect 6711 142 6744 176
rect 6643 127 6744 142
rect 5456 92 6744 127
rect 5456 58 5586 92
rect 5620 58 5676 92
rect 5710 58 5766 92
rect 5800 58 5856 92
rect 5890 58 5946 92
rect 5980 58 6036 92
rect 6070 58 6126 92
rect 6160 58 6216 92
rect 6250 58 6306 92
rect 6340 58 6396 92
rect 6430 58 6486 92
rect 6520 58 6576 92
rect 6610 58 6744 92
rect 5456 26 6744 58
rect 6816 1279 8104 1314
rect 6816 1256 6946 1279
rect 6816 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8104 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8104 1256
rect 6816 1213 8104 1222
rect 6816 1166 6917 1213
rect 6816 1132 6850 1166
rect 6884 1132 6917 1166
rect 8003 1166 8104 1213
rect 6816 1076 6917 1132
rect 6816 1042 6850 1076
rect 6884 1042 6917 1076
rect 6816 986 6917 1042
rect 6816 952 6850 986
rect 6884 952 6917 986
rect 6816 896 6917 952
rect 6816 862 6850 896
rect 6884 862 6917 896
rect 6816 806 6917 862
rect 6816 772 6850 806
rect 6884 772 6917 806
rect 6816 716 6917 772
rect 6816 682 6850 716
rect 6884 682 6917 716
rect 6816 626 6917 682
rect 6816 592 6850 626
rect 6884 592 6917 626
rect 6816 536 6917 592
rect 6816 502 6850 536
rect 6884 502 6917 536
rect 6816 446 6917 502
rect 6816 412 6850 446
rect 6884 412 6917 446
rect 6816 356 6917 412
rect 6816 322 6850 356
rect 6884 322 6917 356
rect 6816 266 6917 322
rect 6816 232 6850 266
rect 6884 232 6917 266
rect 6816 176 6917 232
rect 8003 1132 8037 1166
rect 8071 1132 8104 1166
rect 8003 1076 8104 1132
rect 8003 1042 8037 1076
rect 8071 1042 8104 1076
rect 8003 986 8104 1042
rect 8003 952 8037 986
rect 8071 952 8104 986
rect 8003 896 8104 952
rect 8003 862 8037 896
rect 8071 862 8104 896
rect 8003 806 8104 862
rect 8003 772 8037 806
rect 8071 772 8104 806
rect 8003 716 8104 772
rect 8003 682 8037 716
rect 8071 682 8104 716
rect 8003 626 8104 682
rect 8003 592 8037 626
rect 8071 592 8104 626
rect 8003 536 8104 592
rect 8003 502 8037 536
rect 8071 502 8104 536
rect 8003 446 8104 502
rect 8003 412 8037 446
rect 8071 412 8104 446
rect 8003 356 8104 412
rect 8003 322 8037 356
rect 8071 322 8104 356
rect 8003 266 8104 322
rect 8003 232 8037 266
rect 8071 232 8104 266
rect 6816 142 6850 176
rect 6884 142 6917 176
rect 6816 127 6917 142
rect 8003 176 8104 232
rect 8003 142 8037 176
rect 8071 142 8104 176
rect 8003 127 8104 142
rect 6816 92 8104 127
rect 6816 58 6946 92
rect 6980 58 7036 92
rect 7070 58 7126 92
rect 7160 58 7216 92
rect 7250 58 7306 92
rect 7340 58 7396 92
rect 7430 58 7486 92
rect 7520 58 7576 92
rect 7610 58 7666 92
rect 7700 58 7756 92
rect 7790 58 7846 92
rect 7880 58 7936 92
rect 7970 58 8104 92
rect 6816 26 8104 58
rect 8176 1279 9464 1314
rect 8176 1256 8306 1279
rect 8176 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9464 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9464 1256
rect 8176 1213 9464 1222
rect 8176 1166 8277 1213
rect 8176 1132 8210 1166
rect 8244 1132 8277 1166
rect 9363 1166 9464 1213
rect 8176 1076 8277 1132
rect 8176 1042 8210 1076
rect 8244 1042 8277 1076
rect 8176 986 8277 1042
rect 8176 952 8210 986
rect 8244 952 8277 986
rect 8176 896 8277 952
rect 8176 862 8210 896
rect 8244 862 8277 896
rect 8176 806 8277 862
rect 8176 772 8210 806
rect 8244 772 8277 806
rect 8176 716 8277 772
rect 8176 682 8210 716
rect 8244 682 8277 716
rect 8176 626 8277 682
rect 8176 592 8210 626
rect 8244 592 8277 626
rect 8176 536 8277 592
rect 8176 502 8210 536
rect 8244 502 8277 536
rect 8176 446 8277 502
rect 8176 412 8210 446
rect 8244 412 8277 446
rect 8176 356 8277 412
rect 8176 322 8210 356
rect 8244 322 8277 356
rect 8176 266 8277 322
rect 8176 232 8210 266
rect 8244 232 8277 266
rect 8176 176 8277 232
rect 9363 1132 9397 1166
rect 9431 1132 9464 1166
rect 9363 1076 9464 1132
rect 9363 1042 9397 1076
rect 9431 1042 9464 1076
rect 9363 986 9464 1042
rect 9363 952 9397 986
rect 9431 952 9464 986
rect 9363 896 9464 952
rect 9363 862 9397 896
rect 9431 862 9464 896
rect 9363 806 9464 862
rect 9363 772 9397 806
rect 9431 772 9464 806
rect 9363 716 9464 772
rect 9363 682 9397 716
rect 9431 682 9464 716
rect 9363 626 9464 682
rect 9363 592 9397 626
rect 9431 592 9464 626
rect 9363 536 9464 592
rect 9363 502 9397 536
rect 9431 502 9464 536
rect 9363 446 9464 502
rect 9363 412 9397 446
rect 9431 412 9464 446
rect 9363 356 9464 412
rect 9363 322 9397 356
rect 9431 322 9464 356
rect 9363 266 9464 322
rect 9363 232 9397 266
rect 9431 232 9464 266
rect 8176 142 8210 176
rect 8244 142 8277 176
rect 8176 127 8277 142
rect 9363 176 9464 232
rect 9363 142 9397 176
rect 9431 142 9464 176
rect 9363 127 9464 142
rect 8176 92 9464 127
rect 8176 58 8306 92
rect 8340 58 8396 92
rect 8430 58 8486 92
rect 8520 58 8576 92
rect 8610 58 8666 92
rect 8700 58 8756 92
rect 8790 58 8846 92
rect 8880 58 8936 92
rect 8970 58 9026 92
rect 9060 58 9116 92
rect 9150 58 9206 92
rect 9240 58 9296 92
rect 9330 58 9464 92
rect 8176 26 9464 58
<< nsubdiff >>
rect 4340 5420 4420 5450
rect 4340 5380 4360 5420
rect 4400 5380 4420 5420
rect 4340 5320 4420 5380
rect 4340 5280 4360 5320
rect 4400 5280 4420 5320
rect 4340 5220 4420 5280
rect 4340 5180 4360 5220
rect 4400 5180 4420 5220
rect 4340 5120 4420 5180
rect 4340 5080 4360 5120
rect 4400 5080 4420 5120
rect 4340 5020 4420 5080
rect 4340 4980 4360 5020
rect 4400 4980 4420 5020
rect 4340 4920 4420 4980
rect 4340 4880 4360 4920
rect 4400 4880 4420 4920
rect 4340 4820 4420 4880
rect 4340 4780 4360 4820
rect 4400 4780 4420 4820
rect 4340 4720 4420 4780
rect 4340 4680 4360 4720
rect 4400 4680 4420 4720
rect 4340 4650 4420 4680
rect 8500 5420 8580 5450
rect 8500 5380 8520 5420
rect 8560 5380 8580 5420
rect 8500 5320 8580 5380
rect 8500 5280 8520 5320
rect 8560 5280 8580 5320
rect 8500 5220 8580 5280
rect 8500 5180 8520 5220
rect 8560 5180 8580 5220
rect 8500 5120 8580 5180
rect 8500 5080 8520 5120
rect 8560 5080 8580 5120
rect 8500 5020 8580 5080
rect 8500 4980 8520 5020
rect 8560 4980 8580 5020
rect 8500 4920 8580 4980
rect 8500 4880 8520 4920
rect 8560 4880 8580 4920
rect 8500 4820 8580 4880
rect 8500 4780 8520 4820
rect 8560 4780 8580 4820
rect 8500 4720 8580 4780
rect 8500 4680 8520 4720
rect 8560 4680 8580 4720
rect 8500 4650 8580 4680
rect 4380 4110 4460 4140
rect 4380 4070 4400 4110
rect 4440 4070 4460 4110
rect 4380 4010 4460 4070
rect 4380 3970 4400 4010
rect 4440 3970 4460 4010
rect 4380 3910 4460 3970
rect 4380 3870 4400 3910
rect 4440 3870 4460 3910
rect 4380 3810 4460 3870
rect 4380 3770 4400 3810
rect 4440 3770 4460 3810
rect 4380 3740 4460 3770
rect 5740 4110 5820 4140
rect 5740 4070 5760 4110
rect 5800 4070 5820 4110
rect 5740 4010 5820 4070
rect 5740 3970 5760 4010
rect 5800 3970 5820 4010
rect 5740 3910 5820 3970
rect 5740 3870 5760 3910
rect 5800 3870 5820 3910
rect 5740 3810 5820 3870
rect 5740 3770 5760 3810
rect 5800 3770 5820 3810
rect 5740 3740 5820 3770
rect 7100 4110 7180 4140
rect 7100 4070 7120 4110
rect 7160 4070 7180 4110
rect 7100 4010 7180 4070
rect 7100 3970 7120 4010
rect 7160 3970 7180 4010
rect 7100 3910 7180 3970
rect 7100 3870 7120 3910
rect 7160 3870 7180 3910
rect 7100 3810 7180 3870
rect 7100 3770 7120 3810
rect 7160 3770 7180 3810
rect 7100 3740 7180 3770
rect 8460 4110 8540 4140
rect 8460 4070 8480 4110
rect 8520 4070 8540 4110
rect 8460 4010 8540 4070
rect 8460 3970 8480 4010
rect 8520 3970 8540 4010
rect 8460 3910 8540 3970
rect 8460 3870 8480 3910
rect 8520 3870 8540 3910
rect 8460 3810 8540 3870
rect 8460 3770 8480 3810
rect 8520 3770 8540 3810
rect 8460 3740 8540 3770
rect 9190 4110 9270 4140
rect 9190 4070 9210 4110
rect 9250 4070 9270 4110
rect 9190 4010 9270 4070
rect 9190 3970 9210 4010
rect 9250 3970 9270 4010
rect 9190 3910 9270 3970
rect 9190 3870 9210 3910
rect 9250 3870 9270 3910
rect 9190 3810 9270 3870
rect 9190 3770 9210 3810
rect 9250 3770 9270 3810
rect 9190 3740 9270 3770
rect 1539 1132 2501 1151
rect 1539 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 2501 1132
rect 1539 1079 2501 1098
rect 1539 1075 1611 1079
rect 1539 1041 1558 1075
rect 1592 1041 1611 1075
rect 1539 985 1611 1041
rect 2429 1056 2501 1079
rect 2429 1022 2448 1056
rect 2482 1022 2501 1056
rect 1539 951 1558 985
rect 1592 951 1611 985
rect 1539 895 1611 951
rect 1539 861 1558 895
rect 1592 861 1611 895
rect 1539 805 1611 861
rect 1539 771 1558 805
rect 1592 771 1611 805
rect 1539 715 1611 771
rect 1539 681 1558 715
rect 1592 681 1611 715
rect 1539 625 1611 681
rect 1539 591 1558 625
rect 1592 591 1611 625
rect 1539 535 1611 591
rect 1539 501 1558 535
rect 1592 501 1611 535
rect 1539 445 1611 501
rect 1539 411 1558 445
rect 1592 411 1611 445
rect 1539 355 1611 411
rect 1539 321 1558 355
rect 1592 321 1611 355
rect 2429 966 2501 1022
rect 2429 932 2448 966
rect 2482 932 2501 966
rect 2429 876 2501 932
rect 2429 842 2448 876
rect 2482 842 2501 876
rect 2429 786 2501 842
rect 2429 752 2448 786
rect 2482 752 2501 786
rect 2429 696 2501 752
rect 2429 662 2448 696
rect 2482 662 2501 696
rect 2429 606 2501 662
rect 2429 572 2448 606
rect 2482 572 2501 606
rect 2429 516 2501 572
rect 2429 482 2448 516
rect 2482 482 2501 516
rect 2429 426 2501 482
rect 2429 392 2448 426
rect 2482 392 2501 426
rect 2429 336 2501 392
rect 1539 261 1611 321
rect 2429 302 2448 336
rect 2482 302 2501 336
rect 2429 261 2501 302
rect 1539 242 2501 261
rect 1539 208 1636 242
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 208 2501 242
rect 1539 189 2501 208
rect 2899 1132 3861 1151
rect 2899 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 3861 1132
rect 2899 1079 3861 1098
rect 2899 1075 2971 1079
rect 2899 1041 2918 1075
rect 2952 1041 2971 1075
rect 2899 985 2971 1041
rect 3789 1056 3861 1079
rect 3789 1022 3808 1056
rect 3842 1022 3861 1056
rect 2899 951 2918 985
rect 2952 951 2971 985
rect 2899 895 2971 951
rect 2899 861 2918 895
rect 2952 861 2971 895
rect 2899 805 2971 861
rect 2899 771 2918 805
rect 2952 771 2971 805
rect 2899 715 2971 771
rect 2899 681 2918 715
rect 2952 681 2971 715
rect 2899 625 2971 681
rect 2899 591 2918 625
rect 2952 591 2971 625
rect 2899 535 2971 591
rect 2899 501 2918 535
rect 2952 501 2971 535
rect 2899 445 2971 501
rect 2899 411 2918 445
rect 2952 411 2971 445
rect 2899 355 2971 411
rect 2899 321 2918 355
rect 2952 321 2971 355
rect 3789 966 3861 1022
rect 3789 932 3808 966
rect 3842 932 3861 966
rect 3789 876 3861 932
rect 3789 842 3808 876
rect 3842 842 3861 876
rect 3789 786 3861 842
rect 3789 752 3808 786
rect 3842 752 3861 786
rect 3789 696 3861 752
rect 3789 662 3808 696
rect 3842 662 3861 696
rect 3789 606 3861 662
rect 3789 572 3808 606
rect 3842 572 3861 606
rect 3789 516 3861 572
rect 3789 482 3808 516
rect 3842 482 3861 516
rect 3789 426 3861 482
rect 3789 392 3808 426
rect 3842 392 3861 426
rect 3789 336 3861 392
rect 2899 261 2971 321
rect 3789 302 3808 336
rect 3842 302 3861 336
rect 3789 261 3861 302
rect 2899 242 3861 261
rect 2899 208 2996 242
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 208 3861 242
rect 2899 189 3861 208
rect 4259 1132 5221 1151
rect 4259 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5221 1132
rect 4259 1079 5221 1098
rect 4259 1075 4331 1079
rect 4259 1041 4278 1075
rect 4312 1041 4331 1075
rect 4259 985 4331 1041
rect 5149 1056 5221 1079
rect 5149 1022 5168 1056
rect 5202 1022 5221 1056
rect 4259 951 4278 985
rect 4312 951 4331 985
rect 4259 895 4331 951
rect 4259 861 4278 895
rect 4312 861 4331 895
rect 4259 805 4331 861
rect 4259 771 4278 805
rect 4312 771 4331 805
rect 4259 715 4331 771
rect 4259 681 4278 715
rect 4312 681 4331 715
rect 4259 625 4331 681
rect 4259 591 4278 625
rect 4312 591 4331 625
rect 4259 535 4331 591
rect 4259 501 4278 535
rect 4312 501 4331 535
rect 4259 445 4331 501
rect 4259 411 4278 445
rect 4312 411 4331 445
rect 4259 355 4331 411
rect 4259 321 4278 355
rect 4312 321 4331 355
rect 5149 966 5221 1022
rect 5149 932 5168 966
rect 5202 932 5221 966
rect 5149 876 5221 932
rect 5149 842 5168 876
rect 5202 842 5221 876
rect 5149 786 5221 842
rect 5149 752 5168 786
rect 5202 752 5221 786
rect 5149 696 5221 752
rect 5149 662 5168 696
rect 5202 662 5221 696
rect 5149 606 5221 662
rect 5149 572 5168 606
rect 5202 572 5221 606
rect 5149 516 5221 572
rect 5149 482 5168 516
rect 5202 482 5221 516
rect 5149 426 5221 482
rect 5149 392 5168 426
rect 5202 392 5221 426
rect 5149 336 5221 392
rect 4259 261 4331 321
rect 5149 302 5168 336
rect 5202 302 5221 336
rect 5149 261 5221 302
rect 4259 242 5221 261
rect 4259 208 4356 242
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 208 5221 242
rect 4259 189 5221 208
rect 5619 1132 6581 1151
rect 5619 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 6581 1132
rect 5619 1079 6581 1098
rect 5619 1075 5691 1079
rect 5619 1041 5638 1075
rect 5672 1041 5691 1075
rect 5619 985 5691 1041
rect 6509 1056 6581 1079
rect 6509 1022 6528 1056
rect 6562 1022 6581 1056
rect 5619 951 5638 985
rect 5672 951 5691 985
rect 5619 895 5691 951
rect 5619 861 5638 895
rect 5672 861 5691 895
rect 5619 805 5691 861
rect 5619 771 5638 805
rect 5672 771 5691 805
rect 5619 715 5691 771
rect 5619 681 5638 715
rect 5672 681 5691 715
rect 5619 625 5691 681
rect 5619 591 5638 625
rect 5672 591 5691 625
rect 5619 535 5691 591
rect 5619 501 5638 535
rect 5672 501 5691 535
rect 5619 445 5691 501
rect 5619 411 5638 445
rect 5672 411 5691 445
rect 5619 355 5691 411
rect 5619 321 5638 355
rect 5672 321 5691 355
rect 6509 966 6581 1022
rect 6509 932 6528 966
rect 6562 932 6581 966
rect 6509 876 6581 932
rect 6509 842 6528 876
rect 6562 842 6581 876
rect 6509 786 6581 842
rect 6509 752 6528 786
rect 6562 752 6581 786
rect 6509 696 6581 752
rect 6509 662 6528 696
rect 6562 662 6581 696
rect 6509 606 6581 662
rect 6509 572 6528 606
rect 6562 572 6581 606
rect 6509 516 6581 572
rect 6509 482 6528 516
rect 6562 482 6581 516
rect 6509 426 6581 482
rect 6509 392 6528 426
rect 6562 392 6581 426
rect 6509 336 6581 392
rect 5619 261 5691 321
rect 6509 302 6528 336
rect 6562 302 6581 336
rect 6509 261 6581 302
rect 5619 242 6581 261
rect 5619 208 5716 242
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 208 6581 242
rect 5619 189 6581 208
rect 6979 1132 7941 1151
rect 6979 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 7941 1132
rect 6979 1079 7941 1098
rect 6979 1075 7051 1079
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 7869 1056 7941 1079
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 6979 535 7051 591
rect 6979 501 6998 535
rect 7032 501 7051 535
rect 6979 445 7051 501
rect 6979 411 6998 445
rect 7032 411 7051 445
rect 6979 355 7051 411
rect 6979 321 6998 355
rect 7032 321 7051 355
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 516 7941 572
rect 7869 482 7888 516
rect 7922 482 7941 516
rect 7869 426 7941 482
rect 7869 392 7888 426
rect 7922 392 7941 426
rect 7869 336 7941 392
rect 6979 261 7051 321
rect 7869 302 7888 336
rect 7922 302 7941 336
rect 7869 261 7941 302
rect 6979 242 7941 261
rect 6979 208 7076 242
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 208 7941 242
rect 6979 189 7941 208
rect 8339 1132 9301 1151
rect 8339 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9301 1132
rect 8339 1079 9301 1098
rect 8339 1075 8411 1079
rect 8339 1041 8358 1075
rect 8392 1041 8411 1075
rect 8339 985 8411 1041
rect 9229 1056 9301 1079
rect 9229 1022 9248 1056
rect 9282 1022 9301 1056
rect 8339 951 8358 985
rect 8392 951 8411 985
rect 8339 895 8411 951
rect 8339 861 8358 895
rect 8392 861 8411 895
rect 8339 805 8411 861
rect 8339 771 8358 805
rect 8392 771 8411 805
rect 8339 715 8411 771
rect 8339 681 8358 715
rect 8392 681 8411 715
rect 8339 625 8411 681
rect 8339 591 8358 625
rect 8392 591 8411 625
rect 8339 535 8411 591
rect 8339 501 8358 535
rect 8392 501 8411 535
rect 8339 445 8411 501
rect 8339 411 8358 445
rect 8392 411 8411 445
rect 8339 355 8411 411
rect 8339 321 8358 355
rect 8392 321 8411 355
rect 9229 966 9301 1022
rect 9229 932 9248 966
rect 9282 932 9301 966
rect 9229 876 9301 932
rect 9229 842 9248 876
rect 9282 842 9301 876
rect 9229 786 9301 842
rect 9229 752 9248 786
rect 9282 752 9301 786
rect 9229 696 9301 752
rect 9229 662 9248 696
rect 9282 662 9301 696
rect 9229 606 9301 662
rect 9229 572 9248 606
rect 9282 572 9301 606
rect 9229 516 9301 572
rect 9229 482 9248 516
rect 9282 482 9301 516
rect 9229 426 9301 482
rect 9229 392 9248 426
rect 9282 392 9301 426
rect 9229 336 9301 392
rect 8339 261 8411 321
rect 9229 302 9248 336
rect 9282 302 9301 336
rect 9229 261 9301 302
rect 8339 242 9301 261
rect 8339 208 8436 242
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 208 9301 242
rect 8339 189 9301 208
<< psubdiffcont >>
rect 5080 3260 5120 3300
rect 5080 3160 5120 3200
rect 6440 3260 6480 3300
rect 6440 3160 6480 3200
rect 7800 3260 7840 3300
rect 7800 3160 7840 3200
rect 4600 2710 4640 2750
rect 4600 2610 4640 2650
rect 4600 2510 4640 2550
rect 4600 2410 4640 2450
rect 4600 2310 4640 2350
rect 4600 2210 4640 2250
rect 4600 2110 4640 2150
rect 4600 2010 4640 2050
rect 8280 2710 8320 2750
rect 8280 2610 8320 2650
rect 8280 2510 8320 2550
rect 8280 2410 8320 2450
rect 8280 2310 8320 2350
rect 8280 2210 8320 2250
rect 8280 2110 8320 2150
rect 8280 2010 8320 2050
rect 7540 1640 7580 1680
rect 7540 1540 7580 1580
rect 1410 1222 1444 1256
rect 1506 1245 1540 1279
rect 1596 1245 1630 1279
rect 1686 1245 1720 1279
rect 1776 1245 1810 1279
rect 1866 1245 1900 1279
rect 1956 1245 1990 1279
rect 2046 1245 2080 1279
rect 2136 1245 2170 1279
rect 2226 1245 2260 1279
rect 2316 1245 2350 1279
rect 2406 1245 2440 1279
rect 2496 1245 2530 1279
rect 2597 1222 2631 1256
rect 1410 1132 1444 1166
rect 1410 1042 1444 1076
rect 1410 952 1444 986
rect 1410 862 1444 896
rect 1410 772 1444 806
rect 1410 682 1444 716
rect 1410 592 1444 626
rect 1410 502 1444 536
rect 1410 412 1444 446
rect 1410 322 1444 356
rect 1410 232 1444 266
rect 2597 1132 2631 1166
rect 2597 1042 2631 1076
rect 2597 952 2631 986
rect 2597 862 2631 896
rect 2597 772 2631 806
rect 2597 682 2631 716
rect 2597 592 2631 626
rect 2597 502 2631 536
rect 2597 412 2631 446
rect 2597 322 2631 356
rect 2597 232 2631 266
rect 1410 142 1444 176
rect 2597 142 2631 176
rect 1506 58 1540 92
rect 1596 58 1630 92
rect 1686 58 1720 92
rect 1776 58 1810 92
rect 1866 58 1900 92
rect 1956 58 1990 92
rect 2046 58 2080 92
rect 2136 58 2170 92
rect 2226 58 2260 92
rect 2316 58 2350 92
rect 2406 58 2440 92
rect 2496 58 2530 92
rect 2770 1222 2804 1256
rect 2866 1245 2900 1279
rect 2956 1245 2990 1279
rect 3046 1245 3080 1279
rect 3136 1245 3170 1279
rect 3226 1245 3260 1279
rect 3316 1245 3350 1279
rect 3406 1245 3440 1279
rect 3496 1245 3530 1279
rect 3586 1245 3620 1279
rect 3676 1245 3710 1279
rect 3766 1245 3800 1279
rect 3856 1245 3890 1279
rect 3957 1222 3991 1256
rect 2770 1132 2804 1166
rect 2770 1042 2804 1076
rect 2770 952 2804 986
rect 2770 862 2804 896
rect 2770 772 2804 806
rect 2770 682 2804 716
rect 2770 592 2804 626
rect 2770 502 2804 536
rect 2770 412 2804 446
rect 2770 322 2804 356
rect 2770 232 2804 266
rect 3957 1132 3991 1166
rect 3957 1042 3991 1076
rect 3957 952 3991 986
rect 3957 862 3991 896
rect 3957 772 3991 806
rect 3957 682 3991 716
rect 3957 592 3991 626
rect 3957 502 3991 536
rect 3957 412 3991 446
rect 3957 322 3991 356
rect 3957 232 3991 266
rect 2770 142 2804 176
rect 3957 142 3991 176
rect 2866 58 2900 92
rect 2956 58 2990 92
rect 3046 58 3080 92
rect 3136 58 3170 92
rect 3226 58 3260 92
rect 3316 58 3350 92
rect 3406 58 3440 92
rect 3496 58 3530 92
rect 3586 58 3620 92
rect 3676 58 3710 92
rect 3766 58 3800 92
rect 3856 58 3890 92
rect 4130 1222 4164 1256
rect 4226 1245 4260 1279
rect 4316 1245 4350 1279
rect 4406 1245 4440 1279
rect 4496 1245 4530 1279
rect 4586 1245 4620 1279
rect 4676 1245 4710 1279
rect 4766 1245 4800 1279
rect 4856 1245 4890 1279
rect 4946 1245 4980 1279
rect 5036 1245 5070 1279
rect 5126 1245 5160 1279
rect 5216 1245 5250 1279
rect 5317 1222 5351 1256
rect 4130 1132 4164 1166
rect 4130 1042 4164 1076
rect 4130 952 4164 986
rect 4130 862 4164 896
rect 4130 772 4164 806
rect 4130 682 4164 716
rect 4130 592 4164 626
rect 4130 502 4164 536
rect 4130 412 4164 446
rect 4130 322 4164 356
rect 4130 232 4164 266
rect 5317 1132 5351 1166
rect 5317 1042 5351 1076
rect 5317 952 5351 986
rect 5317 862 5351 896
rect 5317 772 5351 806
rect 5317 682 5351 716
rect 5317 592 5351 626
rect 5317 502 5351 536
rect 5317 412 5351 446
rect 5317 322 5351 356
rect 5317 232 5351 266
rect 4130 142 4164 176
rect 5317 142 5351 176
rect 4226 58 4260 92
rect 4316 58 4350 92
rect 4406 58 4440 92
rect 4496 58 4530 92
rect 4586 58 4620 92
rect 4676 58 4710 92
rect 4766 58 4800 92
rect 4856 58 4890 92
rect 4946 58 4980 92
rect 5036 58 5070 92
rect 5126 58 5160 92
rect 5216 58 5250 92
rect 5490 1222 5524 1256
rect 5586 1245 5620 1279
rect 5676 1245 5710 1279
rect 5766 1245 5800 1279
rect 5856 1245 5890 1279
rect 5946 1245 5980 1279
rect 6036 1245 6070 1279
rect 6126 1245 6160 1279
rect 6216 1245 6250 1279
rect 6306 1245 6340 1279
rect 6396 1245 6430 1279
rect 6486 1245 6520 1279
rect 6576 1245 6610 1279
rect 6677 1222 6711 1256
rect 5490 1132 5524 1166
rect 5490 1042 5524 1076
rect 5490 952 5524 986
rect 5490 862 5524 896
rect 5490 772 5524 806
rect 5490 682 5524 716
rect 5490 592 5524 626
rect 5490 502 5524 536
rect 5490 412 5524 446
rect 5490 322 5524 356
rect 5490 232 5524 266
rect 6677 1132 6711 1166
rect 6677 1042 6711 1076
rect 6677 952 6711 986
rect 6677 862 6711 896
rect 6677 772 6711 806
rect 6677 682 6711 716
rect 6677 592 6711 626
rect 6677 502 6711 536
rect 6677 412 6711 446
rect 6677 322 6711 356
rect 6677 232 6711 266
rect 5490 142 5524 176
rect 6677 142 6711 176
rect 5586 58 5620 92
rect 5676 58 5710 92
rect 5766 58 5800 92
rect 5856 58 5890 92
rect 5946 58 5980 92
rect 6036 58 6070 92
rect 6126 58 6160 92
rect 6216 58 6250 92
rect 6306 58 6340 92
rect 6396 58 6430 92
rect 6486 58 6520 92
rect 6576 58 6610 92
rect 6850 1222 6884 1256
rect 6946 1245 6980 1279
rect 7036 1245 7070 1279
rect 7126 1245 7160 1279
rect 7216 1245 7250 1279
rect 7306 1245 7340 1279
rect 7396 1245 7430 1279
rect 7486 1245 7520 1279
rect 7576 1245 7610 1279
rect 7666 1245 7700 1279
rect 7756 1245 7790 1279
rect 7846 1245 7880 1279
rect 7936 1245 7970 1279
rect 8037 1222 8071 1256
rect 6850 1132 6884 1166
rect 6850 1042 6884 1076
rect 6850 952 6884 986
rect 6850 862 6884 896
rect 6850 772 6884 806
rect 6850 682 6884 716
rect 6850 592 6884 626
rect 6850 502 6884 536
rect 6850 412 6884 446
rect 6850 322 6884 356
rect 6850 232 6884 266
rect 8037 1132 8071 1166
rect 8037 1042 8071 1076
rect 8037 952 8071 986
rect 8037 862 8071 896
rect 8037 772 8071 806
rect 8037 682 8071 716
rect 8037 592 8071 626
rect 8037 502 8071 536
rect 8037 412 8071 446
rect 8037 322 8071 356
rect 8037 232 8071 266
rect 6850 142 6884 176
rect 8037 142 8071 176
rect 6946 58 6980 92
rect 7036 58 7070 92
rect 7126 58 7160 92
rect 7216 58 7250 92
rect 7306 58 7340 92
rect 7396 58 7430 92
rect 7486 58 7520 92
rect 7576 58 7610 92
rect 7666 58 7700 92
rect 7756 58 7790 92
rect 7846 58 7880 92
rect 7936 58 7970 92
rect 8210 1222 8244 1256
rect 8306 1245 8340 1279
rect 8396 1245 8430 1279
rect 8486 1245 8520 1279
rect 8576 1245 8610 1279
rect 8666 1245 8700 1279
rect 8756 1245 8790 1279
rect 8846 1245 8880 1279
rect 8936 1245 8970 1279
rect 9026 1245 9060 1279
rect 9116 1245 9150 1279
rect 9206 1245 9240 1279
rect 9296 1245 9330 1279
rect 9397 1222 9431 1256
rect 8210 1132 8244 1166
rect 8210 1042 8244 1076
rect 8210 952 8244 986
rect 8210 862 8244 896
rect 8210 772 8244 806
rect 8210 682 8244 716
rect 8210 592 8244 626
rect 8210 502 8244 536
rect 8210 412 8244 446
rect 8210 322 8244 356
rect 8210 232 8244 266
rect 9397 1132 9431 1166
rect 9397 1042 9431 1076
rect 9397 952 9431 986
rect 9397 862 9431 896
rect 9397 772 9431 806
rect 9397 682 9431 716
rect 9397 592 9431 626
rect 9397 502 9431 536
rect 9397 412 9431 446
rect 9397 322 9431 356
rect 9397 232 9431 266
rect 8210 142 8244 176
rect 9397 142 9431 176
rect 8306 58 8340 92
rect 8396 58 8430 92
rect 8486 58 8520 92
rect 8576 58 8610 92
rect 8666 58 8700 92
rect 8756 58 8790 92
rect 8846 58 8880 92
rect 8936 58 8970 92
rect 9026 58 9060 92
rect 9116 58 9150 92
rect 9206 58 9240 92
rect 9296 58 9330 92
<< nsubdiffcont >>
rect 4360 5380 4400 5420
rect 4360 5280 4400 5320
rect 4360 5180 4400 5220
rect 4360 5080 4400 5120
rect 4360 4980 4400 5020
rect 4360 4880 4400 4920
rect 4360 4780 4400 4820
rect 4360 4680 4400 4720
rect 8520 5380 8560 5420
rect 8520 5280 8560 5320
rect 8520 5180 8560 5220
rect 8520 5080 8560 5120
rect 8520 4980 8560 5020
rect 8520 4880 8560 4920
rect 8520 4780 8560 4820
rect 8520 4680 8560 4720
rect 4400 4070 4440 4110
rect 4400 3970 4440 4010
rect 4400 3870 4440 3910
rect 4400 3770 4440 3810
rect 5760 4070 5800 4110
rect 5760 3970 5800 4010
rect 5760 3870 5800 3910
rect 5760 3770 5800 3810
rect 7120 4070 7160 4110
rect 7120 3970 7160 4010
rect 7120 3870 7160 3910
rect 7120 3770 7160 3810
rect 8480 4070 8520 4110
rect 8480 3970 8520 4010
rect 8480 3870 8520 3910
rect 8480 3770 8520 3810
rect 9210 4070 9250 4110
rect 9210 3970 9250 4010
rect 9210 3870 9250 3910
rect 9210 3770 9250 3810
rect 1670 1098 1704 1132
rect 1760 1098 1794 1132
rect 1850 1098 1884 1132
rect 1940 1098 1974 1132
rect 2030 1098 2064 1132
rect 2120 1098 2154 1132
rect 2210 1098 2244 1132
rect 2300 1098 2334 1132
rect 2390 1098 2424 1132
rect 1558 1041 1592 1075
rect 2448 1022 2482 1056
rect 1558 951 1592 985
rect 1558 861 1592 895
rect 1558 771 1592 805
rect 1558 681 1592 715
rect 1558 591 1592 625
rect 1558 501 1592 535
rect 1558 411 1592 445
rect 1558 321 1592 355
rect 2448 932 2482 966
rect 2448 842 2482 876
rect 2448 752 2482 786
rect 2448 662 2482 696
rect 2448 572 2482 606
rect 2448 482 2482 516
rect 2448 392 2482 426
rect 2448 302 2482 336
rect 1636 208 1670 242
rect 1726 208 1760 242
rect 1816 208 1850 242
rect 1906 208 1940 242
rect 1996 208 2030 242
rect 2086 208 2120 242
rect 2176 208 2210 242
rect 2266 208 2300 242
rect 2356 208 2390 242
rect 3030 1098 3064 1132
rect 3120 1098 3154 1132
rect 3210 1098 3244 1132
rect 3300 1098 3334 1132
rect 3390 1098 3424 1132
rect 3480 1098 3514 1132
rect 3570 1098 3604 1132
rect 3660 1098 3694 1132
rect 3750 1098 3784 1132
rect 2918 1041 2952 1075
rect 3808 1022 3842 1056
rect 2918 951 2952 985
rect 2918 861 2952 895
rect 2918 771 2952 805
rect 2918 681 2952 715
rect 2918 591 2952 625
rect 2918 501 2952 535
rect 2918 411 2952 445
rect 2918 321 2952 355
rect 3808 932 3842 966
rect 3808 842 3842 876
rect 3808 752 3842 786
rect 3808 662 3842 696
rect 3808 572 3842 606
rect 3808 482 3842 516
rect 3808 392 3842 426
rect 3808 302 3842 336
rect 2996 208 3030 242
rect 3086 208 3120 242
rect 3176 208 3210 242
rect 3266 208 3300 242
rect 3356 208 3390 242
rect 3446 208 3480 242
rect 3536 208 3570 242
rect 3626 208 3660 242
rect 3716 208 3750 242
rect 4390 1098 4424 1132
rect 4480 1098 4514 1132
rect 4570 1098 4604 1132
rect 4660 1098 4694 1132
rect 4750 1098 4784 1132
rect 4840 1098 4874 1132
rect 4930 1098 4964 1132
rect 5020 1098 5054 1132
rect 5110 1098 5144 1132
rect 4278 1041 4312 1075
rect 5168 1022 5202 1056
rect 4278 951 4312 985
rect 4278 861 4312 895
rect 4278 771 4312 805
rect 4278 681 4312 715
rect 4278 591 4312 625
rect 4278 501 4312 535
rect 4278 411 4312 445
rect 4278 321 4312 355
rect 5168 932 5202 966
rect 5168 842 5202 876
rect 5168 752 5202 786
rect 5168 662 5202 696
rect 5168 572 5202 606
rect 5168 482 5202 516
rect 5168 392 5202 426
rect 5168 302 5202 336
rect 4356 208 4390 242
rect 4446 208 4480 242
rect 4536 208 4570 242
rect 4626 208 4660 242
rect 4716 208 4750 242
rect 4806 208 4840 242
rect 4896 208 4930 242
rect 4986 208 5020 242
rect 5076 208 5110 242
rect 5750 1098 5784 1132
rect 5840 1098 5874 1132
rect 5930 1098 5964 1132
rect 6020 1098 6054 1132
rect 6110 1098 6144 1132
rect 6200 1098 6234 1132
rect 6290 1098 6324 1132
rect 6380 1098 6414 1132
rect 6470 1098 6504 1132
rect 5638 1041 5672 1075
rect 6528 1022 6562 1056
rect 5638 951 5672 985
rect 5638 861 5672 895
rect 5638 771 5672 805
rect 5638 681 5672 715
rect 5638 591 5672 625
rect 5638 501 5672 535
rect 5638 411 5672 445
rect 5638 321 5672 355
rect 6528 932 6562 966
rect 6528 842 6562 876
rect 6528 752 6562 786
rect 6528 662 6562 696
rect 6528 572 6562 606
rect 6528 482 6562 516
rect 6528 392 6562 426
rect 6528 302 6562 336
rect 5716 208 5750 242
rect 5806 208 5840 242
rect 5896 208 5930 242
rect 5986 208 6020 242
rect 6076 208 6110 242
rect 6166 208 6200 242
rect 6256 208 6290 242
rect 6346 208 6380 242
rect 6436 208 6470 242
rect 7110 1098 7144 1132
rect 7200 1098 7234 1132
rect 7290 1098 7324 1132
rect 7380 1098 7414 1132
rect 7470 1098 7504 1132
rect 7560 1098 7594 1132
rect 7650 1098 7684 1132
rect 7740 1098 7774 1132
rect 7830 1098 7864 1132
rect 6998 1041 7032 1075
rect 7888 1022 7922 1056
rect 6998 951 7032 985
rect 6998 861 7032 895
rect 6998 771 7032 805
rect 6998 681 7032 715
rect 6998 591 7032 625
rect 6998 501 7032 535
rect 6998 411 7032 445
rect 6998 321 7032 355
rect 7888 932 7922 966
rect 7888 842 7922 876
rect 7888 752 7922 786
rect 7888 662 7922 696
rect 7888 572 7922 606
rect 7888 482 7922 516
rect 7888 392 7922 426
rect 7888 302 7922 336
rect 7076 208 7110 242
rect 7166 208 7200 242
rect 7256 208 7290 242
rect 7346 208 7380 242
rect 7436 208 7470 242
rect 7526 208 7560 242
rect 7616 208 7650 242
rect 7706 208 7740 242
rect 7796 208 7830 242
rect 8470 1098 8504 1132
rect 8560 1098 8594 1132
rect 8650 1098 8684 1132
rect 8740 1098 8774 1132
rect 8830 1098 8864 1132
rect 8920 1098 8954 1132
rect 9010 1098 9044 1132
rect 9100 1098 9134 1132
rect 9190 1098 9224 1132
rect 8358 1041 8392 1075
rect 9248 1022 9282 1056
rect 8358 951 8392 985
rect 8358 861 8392 895
rect 8358 771 8392 805
rect 8358 681 8392 715
rect 8358 591 8392 625
rect 8358 501 8392 535
rect 8358 411 8392 445
rect 8358 321 8392 355
rect 9248 932 9282 966
rect 9248 842 9282 876
rect 9248 752 9282 786
rect 9248 662 9282 696
rect 9248 572 9282 606
rect 9248 482 9282 516
rect 9248 392 9282 426
rect 9248 302 9282 336
rect 8436 208 8470 242
rect 8526 208 8560 242
rect 8616 208 8650 242
rect 8706 208 8740 242
rect 8796 208 8830 242
rect 8886 208 8920 242
rect 8976 208 9010 242
rect 9066 208 9100 242
rect 9156 208 9190 242
<< poly >>
rect 4500 5450 4620 5480
rect 4700 5450 4820 5480
rect 4900 5450 5020 5480
rect 5100 5450 5220 5480
rect 5300 5450 5420 5480
rect 5500 5450 5620 5480
rect 5700 5450 5820 5480
rect 5900 5450 6020 5480
rect 6100 5450 6220 5480
rect 6300 5450 6420 5480
rect 6500 5450 6620 5480
rect 6700 5450 6820 5480
rect 6900 5450 7020 5480
rect 7100 5450 7220 5480
rect 7300 5450 7420 5480
rect 7500 5450 7620 5480
rect 7700 5450 7820 5480
rect 7900 5450 8020 5480
rect 8100 5450 8220 5480
rect 8300 5450 8420 5480
rect 4500 4620 4620 4650
rect 4700 4630 4820 4650
rect 4900 4630 5020 4650
rect 5100 4630 5220 4650
rect 5300 4630 5420 4650
rect 5500 4630 5620 4650
rect 5700 4630 5820 4650
rect 5900 4630 6020 4650
rect 6100 4630 6220 4650
rect 6300 4630 6420 4650
rect 6500 4630 6620 4650
rect 6700 4630 6820 4650
rect 6900 4630 7020 4650
rect 7100 4630 7220 4650
rect 7300 4630 7420 4650
rect 7500 4630 7620 4650
rect 7700 4630 7820 4650
rect 7900 4630 8020 4650
rect 8100 4630 8220 4650
rect 4700 4600 8220 4630
rect 8300 4620 8420 4650
rect 6220 4560 6240 4600
rect 6280 4560 6300 4600
rect 6220 4540 6300 4560
rect 6620 4560 6640 4600
rect 6680 4560 6700 4600
rect 6620 4540 6700 4560
rect 8140 4560 8160 4600
rect 8200 4560 8220 4600
rect 8140 4540 8220 4560
rect 9030 4310 9110 4330
rect 9030 4270 9050 4310
rect 9090 4270 9110 4310
rect 9030 4250 9110 4270
rect 4540 4140 4660 4170
rect 4740 4140 4860 4170
rect 4940 4140 5060 4170
rect 5140 4140 5260 4170
rect 5340 4140 5460 4170
rect 5540 4140 5660 4170
rect 5900 4140 6020 4170
rect 6100 4140 6220 4170
rect 6300 4140 6420 4170
rect 6500 4140 6620 4170
rect 6700 4140 6820 4170
rect 6900 4140 7020 4170
rect 7260 4140 7380 4170
rect 7460 4140 7580 4170
rect 7660 4140 7780 4170
rect 7860 4140 7980 4170
rect 8060 4140 8180 4170
rect 8260 4140 8380 4170
rect 8830 4140 8860 4170
rect 9080 4140 9110 4250
rect 4540 3710 4660 3740
rect 4740 3720 4860 3740
rect 4940 3720 5060 3740
rect 5140 3720 5260 3740
rect 5340 3720 5460 3740
rect 4740 3690 5460 3720
rect 5540 3710 5660 3740
rect 5900 3710 6020 3740
rect 6100 3720 6220 3740
rect 6300 3720 6420 3740
rect 6500 3720 6620 3740
rect 6700 3720 6820 3740
rect 6100 3690 6820 3720
rect 6900 3710 7020 3740
rect 7260 3710 7380 3740
rect 7460 3720 7580 3740
rect 7660 3720 7780 3740
rect 7860 3720 7980 3740
rect 8060 3720 8180 3740
rect 7460 3690 8180 3720
rect 8260 3710 8380 3740
rect 5260 3650 5280 3690
rect 5320 3650 5340 3690
rect 5260 3630 5340 3650
rect 6140 3620 6180 3690
rect 6740 3620 6780 3690
rect 7580 3650 7600 3690
rect 7640 3650 7660 3690
rect 7580 3630 7660 3650
rect 8830 3660 8860 3740
rect 9080 3710 9110 3740
rect 8970 3660 9050 3680
rect 8830 3620 8990 3660
rect 9030 3620 9050 3660
rect 6120 3600 6200 3620
rect 6120 3560 6140 3600
rect 6180 3560 6200 3600
rect 6120 3540 6200 3560
rect 6720 3600 6800 3620
rect 8970 3600 9050 3620
rect 6720 3560 6740 3600
rect 6780 3560 6800 3600
rect 6720 3540 6800 3560
rect 6060 3420 6140 3440
rect 6060 3380 6080 3420
rect 6120 3380 6140 3420
rect 5220 3330 5340 3360
rect 5420 3330 5540 3360
rect 5620 3330 5740 3360
rect 5820 3350 6140 3380
rect 6780 3420 6860 3440
rect 6780 3380 6800 3420
rect 6840 3380 6860 3420
rect 5820 3330 5940 3350
rect 6020 3330 6140 3350
rect 6220 3330 6340 3360
rect 6580 3330 6700 3360
rect 6780 3350 7100 3380
rect 6780 3330 6900 3350
rect 6980 3330 7100 3350
rect 7180 3330 7300 3360
rect 7380 3330 7500 3360
rect 7580 3330 7700 3360
rect 5220 3100 5340 3130
rect 5420 3110 5540 3130
rect 5620 3110 5740 3130
rect 5420 3080 5740 3110
rect 5820 3100 5940 3130
rect 6020 3100 6140 3130
rect 6220 3100 6340 3130
rect 6580 3100 6700 3130
rect 6780 3100 6900 3130
rect 6980 3100 7100 3130
rect 7180 3110 7300 3130
rect 7380 3110 7500 3130
rect 7180 3080 7500 3110
rect 7580 3100 7700 3130
rect 5540 3040 5560 3080
rect 5600 3040 5620 3080
rect 5540 3020 5620 3040
rect 7300 3040 7320 3080
rect 7360 3040 7380 3080
rect 7300 3020 7380 3040
rect 5620 2870 7300 2890
rect 5620 2830 5640 2870
rect 5680 2830 5720 2870
rect 5760 2830 5800 2870
rect 5840 2830 5880 2870
rect 5920 2830 5960 2870
rect 6000 2830 6040 2870
rect 6080 2830 6120 2870
rect 6160 2830 6200 2870
rect 6240 2830 6280 2870
rect 6320 2830 6360 2870
rect 6400 2830 6440 2870
rect 6480 2830 6520 2870
rect 6560 2830 6600 2870
rect 6640 2830 6680 2870
rect 6720 2830 6760 2870
rect 6800 2830 6840 2870
rect 6880 2830 6920 2870
rect 6960 2830 7000 2870
rect 7040 2830 7080 2870
rect 7120 2830 7160 2870
rect 7200 2830 7240 2870
rect 7280 2830 7300 2870
rect 5620 2810 7300 2830
rect 4740 2780 5540 2810
rect 5620 2780 6420 2810
rect 6500 2780 7300 2810
rect 7380 2780 8180 2810
rect 4740 1930 5540 1980
rect 5620 1950 6420 1980
rect 6500 1950 7300 1980
rect 4740 1890 4760 1930
rect 4800 1890 4840 1930
rect 4880 1890 4920 1930
rect 4960 1890 5000 1930
rect 5040 1890 5080 1930
rect 5120 1890 5160 1930
rect 5200 1890 5240 1930
rect 5280 1890 5320 1930
rect 5360 1890 5400 1930
rect 5440 1890 5480 1930
rect 5520 1890 5540 1930
rect 4740 1870 5540 1890
rect 7380 1930 8180 1980
rect 7380 1890 7400 1930
rect 7440 1890 7480 1930
rect 7520 1890 7560 1930
rect 7600 1890 7640 1930
rect 7680 1890 7720 1930
rect 7760 1890 7800 1930
rect 7840 1890 7880 1930
rect 7920 1890 7960 1930
rect 8000 1890 8040 1930
rect 8080 1890 8120 1930
rect 8160 1890 8180 1930
rect 7380 1870 8180 1890
rect 5440 1800 5520 1820
rect 5440 1760 5460 1800
rect 5500 1760 5520 1800
rect 5440 1740 5520 1760
rect 5600 1800 5680 1820
rect 5600 1760 5620 1800
rect 5660 1760 5680 1800
rect 5600 1740 5680 1760
rect 5760 1800 5840 1820
rect 5760 1760 5780 1800
rect 5820 1760 5840 1800
rect 5760 1740 5840 1760
rect 5920 1800 6000 1820
rect 5920 1760 5940 1800
rect 5980 1760 6000 1800
rect 5920 1740 6000 1760
rect 6080 1800 6160 1820
rect 6080 1760 6100 1800
rect 6140 1760 6160 1800
rect 6080 1740 6160 1760
rect 6240 1800 6320 1820
rect 6240 1760 6260 1800
rect 6300 1760 6320 1800
rect 6240 1740 6320 1760
rect 6400 1800 6480 1820
rect 6400 1760 6420 1800
rect 6460 1760 6480 1800
rect 6400 1740 6480 1760
rect 6560 1800 6640 1820
rect 6560 1760 6580 1800
rect 6620 1760 6640 1800
rect 6560 1740 6640 1760
rect 6720 1800 6800 1820
rect 6720 1760 6740 1800
rect 6780 1760 6800 1800
rect 6720 1740 6800 1760
rect 6880 1800 6960 1820
rect 6880 1760 6900 1800
rect 6940 1760 6960 1800
rect 6880 1740 6960 1760
rect 7040 1800 7120 1820
rect 7040 1760 7060 1800
rect 7100 1760 7120 1800
rect 7040 1740 7120 1760
rect 7200 1800 7280 1820
rect 7200 1760 7220 1800
rect 7260 1760 7280 1800
rect 7200 1740 7280 1760
rect 7360 1800 7440 1820
rect 7360 1760 7380 1800
rect 7420 1760 7440 1800
rect 7360 1740 7440 1760
rect 5440 1710 7440 1740
rect 5440 1480 7440 1510
<< polycont >>
rect 6240 4560 6280 4600
rect 6640 4560 6680 4600
rect 8160 4560 8200 4600
rect 9050 4270 9090 4310
rect 5280 3650 5320 3690
rect 7600 3650 7640 3690
rect 8990 3620 9030 3660
rect 6140 3560 6180 3600
rect 6740 3560 6780 3600
rect 6080 3380 6120 3420
rect 6800 3380 6840 3420
rect 5560 3040 5600 3080
rect 7320 3040 7360 3080
rect 5640 2830 5680 2870
rect 5720 2830 5760 2870
rect 5800 2830 5840 2870
rect 5880 2830 5920 2870
rect 5960 2830 6000 2870
rect 6040 2830 6080 2870
rect 6120 2830 6160 2870
rect 6200 2830 6240 2870
rect 6280 2830 6320 2870
rect 6360 2830 6400 2870
rect 6440 2830 6480 2870
rect 6520 2830 6560 2870
rect 6600 2830 6640 2870
rect 6680 2830 6720 2870
rect 6760 2830 6800 2870
rect 6840 2830 6880 2870
rect 6920 2830 6960 2870
rect 7000 2830 7040 2870
rect 7080 2830 7120 2870
rect 7160 2830 7200 2870
rect 7240 2830 7280 2870
rect 4760 1890 4800 1930
rect 4840 1890 4880 1930
rect 4920 1890 4960 1930
rect 5000 1890 5040 1930
rect 5080 1890 5120 1930
rect 5160 1890 5200 1930
rect 5240 1890 5280 1930
rect 5320 1890 5360 1930
rect 5400 1890 5440 1930
rect 5480 1890 5520 1930
rect 7400 1890 7440 1930
rect 7480 1890 7520 1930
rect 7560 1890 7600 1930
rect 7640 1890 7680 1930
rect 7720 1890 7760 1930
rect 7800 1890 7840 1930
rect 7880 1890 7920 1930
rect 7960 1890 8000 1930
rect 8040 1890 8080 1930
rect 8120 1890 8160 1930
rect 5460 1760 5500 1800
rect 5620 1760 5660 1800
rect 5780 1760 5820 1800
rect 5940 1760 5980 1800
rect 6100 1760 6140 1800
rect 6260 1760 6300 1800
rect 6420 1760 6460 1800
rect 6580 1760 6620 1800
rect 6740 1760 6780 1800
rect 6900 1760 6940 1800
rect 7060 1760 7100 1800
rect 7220 1760 7260 1800
rect 7380 1760 7420 1800
<< xpolycontact >>
rect 2010 4970 2450 5040
rect 3790 4970 4230 5040
rect 2010 4850 2450 4920
rect 3790 4850 4230 4920
rect 2010 4730 2450 4800
rect 3790 4730 4230 4800
rect 2010 4610 2450 4680
rect 3790 4610 4230 4680
rect 2010 4490 2450 4560
rect 3790 4490 4230 4560
rect 2010 3970 2450 4040
rect 3790 3970 4230 4040
rect 2010 3850 2450 3920
rect 3790 3850 4230 3920
rect 2010 3730 2450 3800
rect 3790 3730 4230 3800
rect 2010 3610 2450 3680
rect 3790 3610 4230 3680
rect 2010 3490 2450 3560
rect 3790 3490 4230 3560
rect 2010 3020 2450 3090
rect 3150 3020 3590 3090
rect 2010 2900 2450 2970
rect 3790 2900 4230 2970
rect 2010 2780 2450 2850
rect 3790 2780 4230 2850
rect 2010 2660 2450 2730
rect 3790 2660 4230 2730
rect 2010 2540 2450 2610
rect 3790 2540 4230 2610
rect 2010 2420 2450 2490
rect 3790 2420 4230 2490
<< xpolyres >>
rect 2450 4970 3790 5040
rect 2450 4850 3790 4920
rect 2450 4730 3790 4800
rect 2450 4610 3790 4680
rect 2450 4490 3790 4560
rect 2450 3970 3790 4040
rect 2450 3850 3790 3920
rect 2450 3730 3790 3800
rect 2450 3610 3790 3680
rect 2450 3490 3790 3560
rect 2450 3020 3150 3090
rect 2450 2900 3790 2970
rect 2450 2780 3790 2850
rect 2450 2660 3790 2730
rect 2450 2540 3790 2610
rect 2450 2420 3790 2490
<< locali >>
rect 4620 5540 4700 5560
rect 4620 5500 4640 5540
rect 4680 5500 4700 5540
rect 4620 5480 4700 5500
rect 5020 5540 5100 5560
rect 5020 5500 5040 5540
rect 5080 5500 5100 5540
rect 5020 5480 5100 5500
rect 5420 5540 5500 5560
rect 5420 5500 5440 5540
rect 5480 5500 5500 5540
rect 5420 5480 5500 5500
rect 5820 5540 5900 5560
rect 5820 5500 5840 5540
rect 5880 5500 5900 5540
rect 5820 5480 5900 5500
rect 6220 5540 6300 5560
rect 6220 5500 6240 5540
rect 6280 5500 6300 5540
rect 6220 5480 6300 5500
rect 6420 5540 6500 5560
rect 6420 5500 6440 5540
rect 6480 5500 6500 5540
rect 6420 5480 6500 5500
rect 6620 5540 6700 5560
rect 6620 5500 6640 5540
rect 6680 5500 6700 5540
rect 6620 5480 6700 5500
rect 7020 5540 7100 5560
rect 7020 5500 7040 5540
rect 7080 5500 7100 5540
rect 7020 5480 7100 5500
rect 7420 5540 7500 5560
rect 7420 5500 7440 5540
rect 7480 5500 7500 5540
rect 7420 5480 7500 5500
rect 7820 5540 7900 5560
rect 7820 5500 7840 5540
rect 7880 5500 7900 5540
rect 7820 5480 7900 5500
rect 8220 5540 8300 5560
rect 8220 5500 8240 5540
rect 8280 5500 8300 5540
rect 8220 5480 8300 5500
rect 4640 5440 4680 5480
rect 5040 5440 5080 5480
rect 5440 5440 5480 5480
rect 5840 5440 5880 5480
rect 6240 5440 6280 5480
rect 4350 5420 4490 5440
rect 4350 5380 4360 5420
rect 4400 5380 4440 5420
rect 4480 5380 4490 5420
rect 4350 5320 4490 5380
rect 4350 5280 4360 5320
rect 4400 5280 4440 5320
rect 4480 5280 4490 5320
rect 4350 5220 4490 5280
rect 4350 5180 4360 5220
rect 4400 5180 4440 5220
rect 4480 5180 4490 5220
rect 4350 5120 4490 5180
rect 4350 5080 4360 5120
rect 4400 5080 4440 5120
rect 4480 5080 4490 5120
rect 1890 5020 2010 5040
rect 1890 4980 1910 5020
rect 1950 4980 2010 5020
rect 1890 4970 2010 4980
rect 1890 4960 1970 4970
rect 3790 4920 4230 4970
rect 4350 5020 4490 5080
rect 4350 4980 4360 5020
rect 4400 4980 4440 5020
rect 4480 4980 4490 5020
rect 4350 4920 4490 4980
rect 4350 4880 4360 4920
rect 4400 4880 4440 4920
rect 4480 4880 4490 4920
rect 2010 4800 2450 4850
rect 4350 4820 4490 4880
rect 3790 4680 4230 4730
rect 4350 4780 4360 4820
rect 4400 4780 4440 4820
rect 4480 4780 4490 4820
rect 4350 4720 4490 4780
rect 4350 4680 4360 4720
rect 4400 4680 4440 4720
rect 4480 4680 4490 4720
rect 4350 4660 4490 4680
rect 4630 5420 4690 5440
rect 4630 5380 4640 5420
rect 4680 5380 4690 5420
rect 4630 5320 4690 5380
rect 4630 5280 4640 5320
rect 4680 5280 4690 5320
rect 4630 5220 4690 5280
rect 4630 5180 4640 5220
rect 4680 5180 4690 5220
rect 4630 5120 4690 5180
rect 4630 5080 4640 5120
rect 4680 5080 4690 5120
rect 4630 5020 4690 5080
rect 4630 4980 4640 5020
rect 4680 4980 4690 5020
rect 4630 4920 4690 4980
rect 4630 4880 4640 4920
rect 4680 4880 4690 4920
rect 4630 4820 4690 4880
rect 4630 4780 4640 4820
rect 4680 4780 4690 4820
rect 4630 4720 4690 4780
rect 4630 4680 4640 4720
rect 4680 4680 4690 4720
rect 4630 4660 4690 4680
rect 4830 5420 4890 5440
rect 4830 5380 4840 5420
rect 4880 5380 4890 5420
rect 4830 5320 4890 5380
rect 4830 5280 4840 5320
rect 4880 5280 4890 5320
rect 4830 5220 4890 5280
rect 4830 5180 4840 5220
rect 4880 5180 4890 5220
rect 4830 5120 4890 5180
rect 4830 5080 4840 5120
rect 4880 5080 4890 5120
rect 4830 5020 4890 5080
rect 4830 4980 4840 5020
rect 4880 4980 4890 5020
rect 4830 4920 4890 4980
rect 4830 4880 4840 4920
rect 4880 4880 4890 4920
rect 4830 4820 4890 4880
rect 4830 4780 4840 4820
rect 4880 4780 4890 4820
rect 4830 4720 4890 4780
rect 4830 4680 4840 4720
rect 4880 4680 4890 4720
rect 4830 4660 4890 4680
rect 5030 5420 5090 5440
rect 5030 5380 5040 5420
rect 5080 5380 5090 5420
rect 5030 5320 5090 5380
rect 5030 5280 5040 5320
rect 5080 5280 5090 5320
rect 5030 5220 5090 5280
rect 5030 5180 5040 5220
rect 5080 5180 5090 5220
rect 5030 5120 5090 5180
rect 5030 5080 5040 5120
rect 5080 5080 5090 5120
rect 5030 5020 5090 5080
rect 5030 4980 5040 5020
rect 5080 4980 5090 5020
rect 5030 4920 5090 4980
rect 5030 4880 5040 4920
rect 5080 4880 5090 4920
rect 5030 4820 5090 4880
rect 5030 4780 5040 4820
rect 5080 4780 5090 4820
rect 5030 4720 5090 4780
rect 5030 4680 5040 4720
rect 5080 4680 5090 4720
rect 5030 4660 5090 4680
rect 5230 5420 5290 5440
rect 5230 5380 5240 5420
rect 5280 5380 5290 5420
rect 5230 5320 5290 5380
rect 5230 5280 5240 5320
rect 5280 5280 5290 5320
rect 5230 5220 5290 5280
rect 5230 5180 5240 5220
rect 5280 5180 5290 5220
rect 5230 5120 5290 5180
rect 5230 5080 5240 5120
rect 5280 5080 5290 5120
rect 5230 5020 5290 5080
rect 5230 4980 5240 5020
rect 5280 4980 5290 5020
rect 5230 4920 5290 4980
rect 5230 4880 5240 4920
rect 5280 4880 5290 4920
rect 5230 4820 5290 4880
rect 5230 4780 5240 4820
rect 5280 4780 5290 4820
rect 5230 4720 5290 4780
rect 5230 4680 5240 4720
rect 5280 4680 5290 4720
rect 5230 4660 5290 4680
rect 5430 5420 5490 5440
rect 5430 5380 5440 5420
rect 5480 5380 5490 5420
rect 5430 5320 5490 5380
rect 5430 5280 5440 5320
rect 5480 5280 5490 5320
rect 5430 5220 5490 5280
rect 5430 5180 5440 5220
rect 5480 5180 5490 5220
rect 5430 5120 5490 5180
rect 5430 5080 5440 5120
rect 5480 5080 5490 5120
rect 5430 5020 5490 5080
rect 5430 4980 5440 5020
rect 5480 4980 5490 5020
rect 5430 4920 5490 4980
rect 5430 4880 5440 4920
rect 5480 4880 5490 4920
rect 5430 4820 5490 4880
rect 5430 4780 5440 4820
rect 5480 4780 5490 4820
rect 5430 4720 5490 4780
rect 5430 4680 5440 4720
rect 5480 4680 5490 4720
rect 5430 4660 5490 4680
rect 5630 5420 5690 5440
rect 5630 5380 5640 5420
rect 5680 5380 5690 5420
rect 5630 5320 5690 5380
rect 5630 5280 5640 5320
rect 5680 5280 5690 5320
rect 5630 5220 5690 5280
rect 5630 5180 5640 5220
rect 5680 5180 5690 5220
rect 5630 5120 5690 5180
rect 5630 5080 5640 5120
rect 5680 5080 5690 5120
rect 5630 5020 5690 5080
rect 5630 4980 5640 5020
rect 5680 4980 5690 5020
rect 5630 4920 5690 4980
rect 5630 4880 5640 4920
rect 5680 4880 5690 4920
rect 5630 4820 5690 4880
rect 5630 4780 5640 4820
rect 5680 4780 5690 4820
rect 5630 4720 5690 4780
rect 5630 4680 5640 4720
rect 5680 4680 5690 4720
rect 5630 4660 5690 4680
rect 5830 5420 5890 5440
rect 5830 5380 5840 5420
rect 5880 5380 5890 5420
rect 5830 5320 5890 5380
rect 5830 5280 5840 5320
rect 5880 5280 5890 5320
rect 5830 5220 5890 5280
rect 5830 5180 5840 5220
rect 5880 5180 5890 5220
rect 5830 5120 5890 5180
rect 5830 5080 5840 5120
rect 5880 5080 5890 5120
rect 5830 5020 5890 5080
rect 5830 4980 5840 5020
rect 5880 4980 5890 5020
rect 5830 4920 5890 4980
rect 5830 4880 5840 4920
rect 5880 4880 5890 4920
rect 5830 4820 5890 4880
rect 5830 4780 5840 4820
rect 5880 4780 5890 4820
rect 5830 4720 5890 4780
rect 5830 4680 5840 4720
rect 5880 4680 5890 4720
rect 5830 4660 5890 4680
rect 6030 5420 6090 5440
rect 6030 5380 6040 5420
rect 6080 5380 6090 5420
rect 6030 5320 6090 5380
rect 6030 5280 6040 5320
rect 6080 5280 6090 5320
rect 6030 5220 6090 5280
rect 6030 5180 6040 5220
rect 6080 5180 6090 5220
rect 6030 5120 6090 5180
rect 6030 5080 6040 5120
rect 6080 5080 6090 5120
rect 6030 5020 6090 5080
rect 6030 4980 6040 5020
rect 6080 4980 6090 5020
rect 6030 4920 6090 4980
rect 6030 4880 6040 4920
rect 6080 4880 6090 4920
rect 6030 4820 6090 4880
rect 6030 4780 6040 4820
rect 6080 4780 6090 4820
rect 6030 4720 6090 4780
rect 6030 4680 6040 4720
rect 6080 4680 6090 4720
rect 6030 4660 6090 4680
rect 6230 5420 6290 5440
rect 6230 5380 6240 5420
rect 6280 5380 6290 5420
rect 6230 5320 6290 5380
rect 6230 5280 6240 5320
rect 6280 5280 6290 5320
rect 6230 5220 6290 5280
rect 6230 5180 6240 5220
rect 6280 5180 6290 5220
rect 6230 5120 6290 5180
rect 6230 5080 6240 5120
rect 6280 5080 6290 5120
rect 6230 5020 6290 5080
rect 6230 4980 6240 5020
rect 6280 4980 6290 5020
rect 6230 4920 6290 4980
rect 6230 4880 6240 4920
rect 6280 4880 6290 4920
rect 6230 4820 6290 4880
rect 6230 4780 6240 4820
rect 6280 4780 6290 4820
rect 6230 4720 6290 4780
rect 6230 4680 6240 4720
rect 6280 4680 6290 4720
rect 6230 4660 6290 4680
rect 6430 5420 6490 5480
rect 6640 5440 6680 5480
rect 7040 5440 7080 5480
rect 7440 5440 7480 5480
rect 7840 5440 7880 5480
rect 8240 5440 8280 5480
rect 6430 5380 6440 5420
rect 6480 5380 6490 5420
rect 6430 5320 6490 5380
rect 6430 5280 6440 5320
rect 6480 5280 6490 5320
rect 6430 5220 6490 5280
rect 6430 5180 6440 5220
rect 6480 5180 6490 5220
rect 6430 5120 6490 5180
rect 6430 5080 6440 5120
rect 6480 5080 6490 5120
rect 6430 5020 6490 5080
rect 6430 4980 6440 5020
rect 6480 4980 6490 5020
rect 6430 4920 6490 4980
rect 6430 4880 6440 4920
rect 6480 4880 6490 4920
rect 6430 4820 6490 4880
rect 6430 4780 6440 4820
rect 6480 4780 6490 4820
rect 6430 4720 6490 4780
rect 6430 4680 6440 4720
rect 6480 4680 6490 4720
rect 6430 4660 6490 4680
rect 6630 5420 6690 5440
rect 6630 5380 6640 5420
rect 6680 5380 6690 5420
rect 6630 5320 6690 5380
rect 6630 5280 6640 5320
rect 6680 5280 6690 5320
rect 6630 5220 6690 5280
rect 6630 5180 6640 5220
rect 6680 5180 6690 5220
rect 6630 5120 6690 5180
rect 6630 5080 6640 5120
rect 6680 5080 6690 5120
rect 6630 5020 6690 5080
rect 6630 4980 6640 5020
rect 6680 4980 6690 5020
rect 6630 4920 6690 4980
rect 6630 4880 6640 4920
rect 6680 4880 6690 4920
rect 6630 4820 6690 4880
rect 6630 4780 6640 4820
rect 6680 4780 6690 4820
rect 6630 4720 6690 4780
rect 6630 4680 6640 4720
rect 6680 4680 6690 4720
rect 6630 4660 6690 4680
rect 6830 5420 6890 5440
rect 6830 5380 6840 5420
rect 6880 5380 6890 5420
rect 6830 5320 6890 5380
rect 6830 5280 6840 5320
rect 6880 5280 6890 5320
rect 6830 5220 6890 5280
rect 6830 5180 6840 5220
rect 6880 5180 6890 5220
rect 6830 5120 6890 5180
rect 6830 5080 6840 5120
rect 6880 5080 6890 5120
rect 6830 5020 6890 5080
rect 6830 4980 6840 5020
rect 6880 4980 6890 5020
rect 6830 4920 6890 4980
rect 6830 4880 6840 4920
rect 6880 4880 6890 4920
rect 6830 4820 6890 4880
rect 6830 4780 6840 4820
rect 6880 4780 6890 4820
rect 6830 4720 6890 4780
rect 6830 4680 6840 4720
rect 6880 4680 6890 4720
rect 6830 4660 6890 4680
rect 7030 5420 7090 5440
rect 7030 5380 7040 5420
rect 7080 5380 7090 5420
rect 7030 5320 7090 5380
rect 7030 5280 7040 5320
rect 7080 5280 7090 5320
rect 7030 5220 7090 5280
rect 7030 5180 7040 5220
rect 7080 5180 7090 5220
rect 7030 5120 7090 5180
rect 7030 5080 7040 5120
rect 7080 5080 7090 5120
rect 7030 5020 7090 5080
rect 7030 4980 7040 5020
rect 7080 4980 7090 5020
rect 7030 4920 7090 4980
rect 7030 4880 7040 4920
rect 7080 4880 7090 4920
rect 7030 4820 7090 4880
rect 7030 4780 7040 4820
rect 7080 4780 7090 4820
rect 7030 4720 7090 4780
rect 7030 4680 7040 4720
rect 7080 4680 7090 4720
rect 7030 4660 7090 4680
rect 7230 5420 7290 5440
rect 7230 5380 7240 5420
rect 7280 5380 7290 5420
rect 7230 5320 7290 5380
rect 7230 5280 7240 5320
rect 7280 5280 7290 5320
rect 7230 5220 7290 5280
rect 7230 5180 7240 5220
rect 7280 5180 7290 5220
rect 7230 5120 7290 5180
rect 7230 5080 7240 5120
rect 7280 5080 7290 5120
rect 7230 5020 7290 5080
rect 7230 4980 7240 5020
rect 7280 4980 7290 5020
rect 7230 4920 7290 4980
rect 7230 4880 7240 4920
rect 7280 4880 7290 4920
rect 7230 4820 7290 4880
rect 7230 4780 7240 4820
rect 7280 4780 7290 4820
rect 7230 4720 7290 4780
rect 7230 4680 7240 4720
rect 7280 4680 7290 4720
rect 7230 4660 7290 4680
rect 7430 5420 7490 5440
rect 7430 5380 7440 5420
rect 7480 5380 7490 5420
rect 7430 5320 7490 5380
rect 7430 5280 7440 5320
rect 7480 5280 7490 5320
rect 7430 5220 7490 5280
rect 7430 5180 7440 5220
rect 7480 5180 7490 5220
rect 7430 5120 7490 5180
rect 7430 5080 7440 5120
rect 7480 5080 7490 5120
rect 7430 5020 7490 5080
rect 7430 4980 7440 5020
rect 7480 4980 7490 5020
rect 7430 4920 7490 4980
rect 7430 4880 7440 4920
rect 7480 4880 7490 4920
rect 7430 4820 7490 4880
rect 7430 4780 7440 4820
rect 7480 4780 7490 4820
rect 7430 4720 7490 4780
rect 7430 4680 7440 4720
rect 7480 4680 7490 4720
rect 7430 4660 7490 4680
rect 7630 5420 7690 5440
rect 7630 5380 7640 5420
rect 7680 5380 7690 5420
rect 7630 5320 7690 5380
rect 7630 5280 7640 5320
rect 7680 5280 7690 5320
rect 7630 5220 7690 5280
rect 7630 5180 7640 5220
rect 7680 5180 7690 5220
rect 7630 5120 7690 5180
rect 7630 5080 7640 5120
rect 7680 5080 7690 5120
rect 7630 5020 7690 5080
rect 7630 4980 7640 5020
rect 7680 4980 7690 5020
rect 7630 4920 7690 4980
rect 7630 4880 7640 4920
rect 7680 4880 7690 4920
rect 7630 4820 7690 4880
rect 7630 4780 7640 4820
rect 7680 4780 7690 4820
rect 7630 4720 7690 4780
rect 7630 4680 7640 4720
rect 7680 4680 7690 4720
rect 7630 4660 7690 4680
rect 7830 5420 7890 5440
rect 7830 5380 7840 5420
rect 7880 5380 7890 5420
rect 7830 5320 7890 5380
rect 7830 5280 7840 5320
rect 7880 5280 7890 5320
rect 7830 5220 7890 5280
rect 7830 5180 7840 5220
rect 7880 5180 7890 5220
rect 7830 5120 7890 5180
rect 7830 5080 7840 5120
rect 7880 5080 7890 5120
rect 7830 5020 7890 5080
rect 7830 4980 7840 5020
rect 7880 4980 7890 5020
rect 7830 4920 7890 4980
rect 7830 4880 7840 4920
rect 7880 4880 7890 4920
rect 7830 4820 7890 4880
rect 7830 4780 7840 4820
rect 7880 4780 7890 4820
rect 7830 4720 7890 4780
rect 7830 4680 7840 4720
rect 7880 4680 7890 4720
rect 7830 4660 7890 4680
rect 8030 5420 8090 5440
rect 8030 5380 8040 5420
rect 8080 5380 8090 5420
rect 8030 5320 8090 5380
rect 8030 5280 8040 5320
rect 8080 5280 8090 5320
rect 8030 5220 8090 5280
rect 8030 5180 8040 5220
rect 8080 5180 8090 5220
rect 8030 5120 8090 5180
rect 8030 5080 8040 5120
rect 8080 5080 8090 5120
rect 8030 5020 8090 5080
rect 8030 4980 8040 5020
rect 8080 4980 8090 5020
rect 8030 4920 8090 4980
rect 8030 4880 8040 4920
rect 8080 4880 8090 4920
rect 8030 4820 8090 4880
rect 8030 4780 8040 4820
rect 8080 4780 8090 4820
rect 8030 4720 8090 4780
rect 8030 4680 8040 4720
rect 8080 4680 8090 4720
rect 8030 4660 8090 4680
rect 8230 5420 8290 5440
rect 8230 5380 8240 5420
rect 8280 5380 8290 5420
rect 8230 5320 8290 5380
rect 8230 5280 8240 5320
rect 8280 5280 8290 5320
rect 8230 5220 8290 5280
rect 8230 5180 8240 5220
rect 8280 5180 8290 5220
rect 8230 5120 8290 5180
rect 8230 5080 8240 5120
rect 8280 5080 8290 5120
rect 8230 5020 8290 5080
rect 8230 4980 8240 5020
rect 8280 4980 8290 5020
rect 8230 4920 8290 4980
rect 8230 4880 8240 4920
rect 8280 4880 8290 4920
rect 8230 4820 8290 4880
rect 8230 4780 8240 4820
rect 8280 4780 8290 4820
rect 8230 4720 8290 4780
rect 8230 4680 8240 4720
rect 8280 4680 8290 4720
rect 8230 4660 8290 4680
rect 8430 5420 8570 5440
rect 8430 5380 8440 5420
rect 8480 5380 8520 5420
rect 8560 5380 8570 5420
rect 8430 5320 8570 5380
rect 8430 5280 8440 5320
rect 8480 5280 8520 5320
rect 8560 5280 8570 5320
rect 8430 5220 8570 5280
rect 8430 5180 8440 5220
rect 8480 5180 8520 5220
rect 8560 5180 8570 5220
rect 8430 5120 8570 5180
rect 8430 5080 8440 5120
rect 8480 5080 8520 5120
rect 8560 5080 8570 5120
rect 8430 5020 8570 5080
rect 8430 4980 8440 5020
rect 8480 4980 8520 5020
rect 8560 4980 8570 5020
rect 8430 4920 8570 4980
rect 8430 4880 8440 4920
rect 8480 4880 8520 4920
rect 8560 4880 8570 4920
rect 8430 4820 8570 4880
rect 8430 4780 8440 4820
rect 8480 4780 8520 4820
rect 8560 4780 8570 4820
rect 8430 4720 8570 4780
rect 8430 4680 8440 4720
rect 8480 4680 8520 4720
rect 8560 4680 8570 4720
rect 8430 4660 8570 4680
rect 4840 4620 4880 4660
rect 2010 4560 2450 4610
rect 4820 4600 4900 4620
rect 4820 4560 4840 4600
rect 4880 4560 4900 4600
rect 4820 4540 4900 4560
rect 5240 4530 5280 4660
rect 3790 4430 4230 4490
rect 5220 4510 5300 4530
rect 5220 4470 5240 4510
rect 5280 4470 5300 4510
rect 5220 4450 5300 4470
rect 5640 4440 5680 4660
rect 6040 4530 6080 4660
rect 6220 4600 6300 4620
rect 6220 4560 6240 4600
rect 6280 4560 6300 4600
rect 6220 4540 6300 4560
rect 6020 4510 6100 4530
rect 6020 4470 6040 4510
rect 6080 4470 6100 4510
rect 6020 4450 6100 4470
rect 6440 4440 6480 4660
rect 6840 4620 6880 4660
rect 6620 4600 6700 4620
rect 6620 4560 6640 4600
rect 6680 4560 6700 4600
rect 6620 4540 6700 4560
rect 6820 4600 6900 4620
rect 6820 4560 6840 4600
rect 6880 4560 6900 4600
rect 6820 4540 6900 4560
rect 7240 4440 7280 4660
rect 7640 4620 7680 4660
rect 7620 4600 7700 4620
rect 7620 4560 7640 4600
rect 7680 4560 7700 4600
rect 7620 4540 7700 4560
rect 8040 4530 8080 4660
rect 8140 4600 8220 4620
rect 8140 4560 8160 4600
rect 8200 4560 8220 4600
rect 8140 4540 8220 4560
rect 8020 4510 8100 4530
rect 8020 4470 8040 4510
rect 8080 4470 8100 4510
rect 8020 4450 8100 4470
rect 3790 4390 3810 4430
rect 3850 4390 3900 4430
rect 3940 4390 3990 4430
rect 4030 4390 4080 4430
rect 4120 4390 4170 4430
rect 4210 4390 4230 4430
rect 3790 4370 4230 4390
rect 5620 4420 5700 4440
rect 5620 4380 5640 4420
rect 5680 4380 5700 4420
rect 5620 4360 5700 4380
rect 6420 4420 6500 4440
rect 6420 4380 6440 4420
rect 6480 4380 6500 4420
rect 6420 4360 6500 4380
rect 7220 4420 7300 4440
rect 7220 4380 7240 4420
rect 7280 4380 7300 4420
rect 7220 4360 7300 4380
rect 8750 4330 8830 4350
rect 8750 4290 8770 4330
rect 8810 4310 9110 4330
rect 8810 4290 9050 4310
rect 8750 4270 8830 4290
rect 9030 4270 9050 4290
rect 9090 4270 9110 4310
rect 4460 4230 4540 4250
rect 4460 4190 4480 4230
rect 4520 4190 4540 4230
rect 4460 4170 4540 4190
rect 4660 4230 4740 4250
rect 4660 4190 4680 4230
rect 4720 4190 4740 4230
rect 4660 4170 4740 4190
rect 5060 4230 5140 4250
rect 5060 4190 5080 4230
rect 5120 4190 5140 4230
rect 5060 4170 5140 4190
rect 5460 4230 5540 4250
rect 5460 4190 5480 4230
rect 5520 4190 5540 4230
rect 5460 4170 5540 4190
rect 5660 4230 5740 4250
rect 5660 4190 5680 4230
rect 5720 4190 5740 4230
rect 5660 4170 5740 4190
rect 5820 4230 5900 4250
rect 5820 4190 5840 4230
rect 5880 4190 5900 4230
rect 5820 4170 5900 4190
rect 6020 4230 6100 4250
rect 6020 4190 6040 4230
rect 6080 4190 6100 4230
rect 6020 4170 6100 4190
rect 6220 4230 6300 4250
rect 6220 4190 6240 4230
rect 6280 4190 6300 4230
rect 6220 4170 6300 4190
rect 6420 4230 6500 4250
rect 6420 4190 6440 4230
rect 6480 4190 6500 4230
rect 6420 4170 6500 4190
rect 6620 4230 6700 4250
rect 6620 4190 6640 4230
rect 6680 4190 6700 4230
rect 6620 4170 6700 4190
rect 6820 4230 6900 4250
rect 6820 4190 6840 4230
rect 6880 4190 6900 4230
rect 6820 4170 6900 4190
rect 7020 4230 7100 4250
rect 7020 4190 7040 4230
rect 7080 4190 7100 4230
rect 7020 4170 7100 4190
rect 7180 4230 7260 4250
rect 7180 4190 7200 4230
rect 7240 4190 7260 4230
rect 7180 4170 7260 4190
rect 7380 4230 7460 4250
rect 7380 4190 7400 4230
rect 7440 4190 7460 4230
rect 7380 4170 7460 4190
rect 7780 4230 7860 4250
rect 7780 4190 7800 4230
rect 7840 4190 7860 4230
rect 7780 4170 7860 4190
rect 8180 4230 8260 4250
rect 8180 4190 8200 4230
rect 8240 4190 8260 4230
rect 8180 4170 8260 4190
rect 8380 4230 8460 4250
rect 8380 4190 8400 4230
rect 8440 4190 8460 4230
rect 8380 4170 8460 4190
rect 4480 4130 4520 4170
rect 4680 4130 4720 4170
rect 5080 4130 5120 4170
rect 5480 4130 5520 4170
rect 5680 4130 5720 4170
rect 5840 4130 5880 4170
rect 6040 4130 6080 4170
rect 6240 4130 6280 4170
rect 6440 4130 6480 4170
rect 6640 4130 6680 4170
rect 6840 4130 6880 4170
rect 7040 4130 7080 4170
rect 7200 4130 7240 4170
rect 7400 4130 7440 4170
rect 7800 4130 7840 4170
rect 8200 4130 8240 4170
rect 8400 4130 8440 4170
rect 8770 4130 8810 4270
rect 9030 4250 9110 4270
rect 9150 4230 9230 4250
rect 9150 4190 9170 4230
rect 9210 4190 9230 4230
rect 9150 4170 9230 4190
rect 9170 4130 9210 4170
rect 4390 4110 4530 4130
rect 4390 4070 4400 4110
rect 4440 4070 4480 4110
rect 4520 4070 4530 4110
rect 1890 4020 2010 4040
rect 1890 3980 1910 4020
rect 1950 3980 2010 4020
rect 1890 3970 2010 3980
rect 1890 3960 1970 3970
rect 3790 3920 4230 3970
rect 4390 4010 4530 4070
rect 4390 3970 4400 4010
rect 4440 3970 4480 4010
rect 4520 3970 4530 4010
rect 4390 3910 4530 3970
rect 4390 3870 4400 3910
rect 4440 3870 4480 3910
rect 4520 3870 4530 3910
rect 2010 3800 2450 3850
rect 4390 3810 4530 3870
rect 4390 3770 4400 3810
rect 4440 3770 4480 3810
rect 4520 3770 4530 3810
rect 4390 3750 4530 3770
rect 4670 4110 4730 4130
rect 4670 4070 4680 4110
rect 4720 4070 4730 4110
rect 4670 4010 4730 4070
rect 4670 3970 4680 4010
rect 4720 3970 4730 4010
rect 4670 3910 4730 3970
rect 4670 3870 4680 3910
rect 4720 3870 4730 3910
rect 4670 3810 4730 3870
rect 4670 3770 4680 3810
rect 4720 3770 4730 3810
rect 4670 3750 4730 3770
rect 4870 4110 4930 4130
rect 4870 4070 4880 4110
rect 4920 4070 4930 4110
rect 4870 4010 4930 4070
rect 4870 3970 4880 4010
rect 4920 3970 4930 4010
rect 4870 3910 4930 3970
rect 4870 3870 4880 3910
rect 4920 3870 4930 3910
rect 4870 3810 4930 3870
rect 4870 3770 4880 3810
rect 4920 3770 4930 3810
rect 4870 3750 4930 3770
rect 5070 4110 5130 4130
rect 5070 4070 5080 4110
rect 5120 4070 5130 4110
rect 5070 4010 5130 4070
rect 5070 3970 5080 4010
rect 5120 3970 5130 4010
rect 5070 3910 5130 3970
rect 5070 3870 5080 3910
rect 5120 3870 5130 3910
rect 5070 3810 5130 3870
rect 5070 3770 5080 3810
rect 5120 3770 5130 3810
rect 5070 3750 5130 3770
rect 5270 4110 5330 4130
rect 5270 4070 5280 4110
rect 5320 4070 5330 4110
rect 5270 4010 5330 4070
rect 5270 3970 5280 4010
rect 5320 3970 5330 4010
rect 5270 3910 5330 3970
rect 5270 3870 5280 3910
rect 5320 3870 5330 3910
rect 5270 3810 5330 3870
rect 5270 3770 5280 3810
rect 5320 3770 5330 3810
rect 5270 3750 5330 3770
rect 5470 4110 5530 4130
rect 5470 4070 5480 4110
rect 5520 4070 5530 4110
rect 5470 4010 5530 4070
rect 5470 3970 5480 4010
rect 5520 3970 5530 4010
rect 5470 3910 5530 3970
rect 5470 3870 5480 3910
rect 5520 3870 5530 3910
rect 5470 3810 5530 3870
rect 5470 3770 5480 3810
rect 5520 3770 5530 3810
rect 5470 3750 5530 3770
rect 5670 4110 5890 4130
rect 5670 4070 5680 4110
rect 5720 4070 5760 4110
rect 5800 4070 5840 4110
rect 5880 4070 5890 4110
rect 5670 4010 5890 4070
rect 5670 3970 5680 4010
rect 5720 3970 5760 4010
rect 5800 3970 5840 4010
rect 5880 3970 5890 4010
rect 5670 3910 5890 3970
rect 5670 3870 5680 3910
rect 5720 3870 5760 3910
rect 5800 3870 5840 3910
rect 5880 3870 5890 3910
rect 5670 3810 5890 3870
rect 5670 3770 5680 3810
rect 5720 3770 5760 3810
rect 5800 3770 5840 3810
rect 5880 3770 5890 3810
rect 5670 3750 5890 3770
rect 6030 4110 6090 4130
rect 6030 4070 6040 4110
rect 6080 4070 6090 4110
rect 6030 4010 6090 4070
rect 6030 3970 6040 4010
rect 6080 3970 6090 4010
rect 6030 3910 6090 3970
rect 6030 3870 6040 3910
rect 6080 3870 6090 3910
rect 6030 3810 6090 3870
rect 6030 3770 6040 3810
rect 6080 3770 6090 3810
rect 6030 3750 6090 3770
rect 6230 4110 6290 4130
rect 6230 4070 6240 4110
rect 6280 4070 6290 4110
rect 6230 4010 6290 4070
rect 6230 3970 6240 4010
rect 6280 3970 6290 4010
rect 6230 3910 6290 3970
rect 6230 3870 6240 3910
rect 6280 3870 6290 3910
rect 6230 3810 6290 3870
rect 6230 3770 6240 3810
rect 6280 3770 6290 3810
rect 6230 3750 6290 3770
rect 6430 4110 6490 4130
rect 6430 4070 6440 4110
rect 6480 4070 6490 4110
rect 6430 4010 6490 4070
rect 6430 3970 6440 4010
rect 6480 3970 6490 4010
rect 6430 3910 6490 3970
rect 6430 3870 6440 3910
rect 6480 3870 6490 3910
rect 6430 3810 6490 3870
rect 6430 3770 6440 3810
rect 6480 3770 6490 3810
rect 6430 3750 6490 3770
rect 6630 4110 6690 4130
rect 6630 4070 6640 4110
rect 6680 4070 6690 4110
rect 6630 4010 6690 4070
rect 6630 3970 6640 4010
rect 6680 3970 6690 4010
rect 6630 3910 6690 3970
rect 6630 3870 6640 3910
rect 6680 3870 6690 3910
rect 6630 3810 6690 3870
rect 6630 3770 6640 3810
rect 6680 3770 6690 3810
rect 6630 3750 6690 3770
rect 6830 4110 6890 4130
rect 6830 4070 6840 4110
rect 6880 4070 6890 4110
rect 6830 4010 6890 4070
rect 6830 3970 6840 4010
rect 6880 3970 6890 4010
rect 6830 3910 6890 3970
rect 6830 3870 6840 3910
rect 6880 3870 6890 3910
rect 6830 3810 6890 3870
rect 6830 3770 6840 3810
rect 6880 3770 6890 3810
rect 6830 3750 6890 3770
rect 7030 4110 7250 4130
rect 7030 4070 7040 4110
rect 7080 4070 7120 4110
rect 7160 4070 7200 4110
rect 7240 4070 7250 4110
rect 7030 4010 7250 4070
rect 7030 3970 7040 4010
rect 7080 3970 7120 4010
rect 7160 3970 7200 4010
rect 7240 3970 7250 4010
rect 7030 3910 7250 3970
rect 7030 3870 7040 3910
rect 7080 3870 7120 3910
rect 7160 3870 7200 3910
rect 7240 3870 7250 3910
rect 7030 3810 7250 3870
rect 7030 3770 7040 3810
rect 7080 3770 7120 3810
rect 7160 3770 7200 3810
rect 7240 3770 7250 3810
rect 7030 3750 7250 3770
rect 7390 4110 7450 4130
rect 7390 4070 7400 4110
rect 7440 4070 7450 4110
rect 7390 4010 7450 4070
rect 7390 3970 7400 4010
rect 7440 3970 7450 4010
rect 7390 3910 7450 3970
rect 7390 3870 7400 3910
rect 7440 3870 7450 3910
rect 7390 3810 7450 3870
rect 7390 3770 7400 3810
rect 7440 3770 7450 3810
rect 7390 3750 7450 3770
rect 7590 4110 7650 4130
rect 7590 4070 7600 4110
rect 7640 4070 7650 4110
rect 7590 4010 7650 4070
rect 7590 3970 7600 4010
rect 7640 3970 7650 4010
rect 7590 3910 7650 3970
rect 7590 3870 7600 3910
rect 7640 3870 7650 3910
rect 7590 3810 7650 3870
rect 7590 3770 7600 3810
rect 7640 3770 7650 3810
rect 7590 3750 7650 3770
rect 7790 4110 7850 4130
rect 7790 4070 7800 4110
rect 7840 4070 7850 4110
rect 7790 4010 7850 4070
rect 7790 3970 7800 4010
rect 7840 3970 7850 4010
rect 7790 3910 7850 3970
rect 7790 3870 7800 3910
rect 7840 3870 7850 3910
rect 7790 3810 7850 3870
rect 7790 3770 7800 3810
rect 7840 3770 7850 3810
rect 7790 3750 7850 3770
rect 7990 4110 8050 4130
rect 7990 4070 8000 4110
rect 8040 4070 8050 4110
rect 7990 4010 8050 4070
rect 7990 3970 8000 4010
rect 8040 3970 8050 4010
rect 7990 3910 8050 3970
rect 7990 3870 8000 3910
rect 8040 3870 8050 3910
rect 7990 3810 8050 3870
rect 7990 3770 8000 3810
rect 8040 3770 8050 3810
rect 7990 3750 8050 3770
rect 8190 4110 8250 4130
rect 8190 4070 8200 4110
rect 8240 4070 8250 4110
rect 8190 4010 8250 4070
rect 8190 3970 8200 4010
rect 8240 3970 8250 4010
rect 8190 3910 8250 3970
rect 8190 3870 8200 3910
rect 8240 3870 8250 3910
rect 8190 3810 8250 3870
rect 8190 3770 8200 3810
rect 8240 3770 8250 3810
rect 8190 3750 8250 3770
rect 8390 4110 8530 4130
rect 8390 4070 8400 4110
rect 8440 4070 8480 4110
rect 8520 4070 8530 4110
rect 8390 4010 8530 4070
rect 8390 3970 8400 4010
rect 8440 3970 8480 4010
rect 8520 3970 8530 4010
rect 8390 3910 8530 3970
rect 8390 3870 8400 3910
rect 8440 3870 8480 3910
rect 8520 3870 8530 3910
rect 8390 3810 8530 3870
rect 8390 3770 8400 3810
rect 8440 3770 8480 3810
rect 8520 3770 8530 3810
rect 8390 3750 8530 3770
rect 8760 4110 8820 4130
rect 8760 4070 8770 4110
rect 8810 4070 8820 4110
rect 8760 4010 8820 4070
rect 8760 3970 8770 4010
rect 8810 3970 8820 4010
rect 8760 3910 8820 3970
rect 8760 3870 8770 3910
rect 8810 3870 8820 3910
rect 8760 3810 8820 3870
rect 8760 3770 8770 3810
rect 8810 3770 8820 3810
rect 8760 3750 8820 3770
rect 8870 4110 8930 4130
rect 8870 4070 8880 4110
rect 8920 4070 8930 4110
rect 8870 4010 8930 4070
rect 8870 3970 8880 4010
rect 8920 3970 8930 4010
rect 8870 3910 8930 3970
rect 8870 3870 8880 3910
rect 8920 3870 8930 3910
rect 8870 3810 8930 3870
rect 8870 3770 8880 3810
rect 8920 3770 8930 3810
rect 8870 3750 8930 3770
rect 9010 4110 9070 4130
rect 9010 4070 9020 4110
rect 9060 4070 9070 4110
rect 9010 4010 9070 4070
rect 9010 3970 9020 4010
rect 9060 3970 9070 4010
rect 9010 3910 9070 3970
rect 9010 3870 9020 3910
rect 9060 3870 9070 3910
rect 9010 3810 9070 3870
rect 9010 3770 9020 3810
rect 9060 3770 9070 3810
rect 9010 3750 9070 3770
rect 9120 4110 9260 4130
rect 9120 4070 9130 4110
rect 9170 4070 9210 4110
rect 9250 4070 9260 4110
rect 9120 4010 9260 4070
rect 9120 3970 9130 4010
rect 9170 3970 9210 4010
rect 9250 3970 9260 4010
rect 9120 3910 9260 3970
rect 9120 3870 9130 3910
rect 9170 3870 9210 3910
rect 9250 3870 9260 3910
rect 9120 3810 9260 3870
rect 9120 3770 9130 3810
rect 9170 3770 9210 3810
rect 9250 3770 9260 3810
rect 9120 3750 9260 3770
rect 3790 3680 4230 3730
rect 4880 3620 4920 3750
rect 5280 3710 5320 3750
rect 6240 3710 6280 3750
rect 6640 3710 6680 3750
rect 7600 3710 7640 3750
rect 5260 3690 5340 3710
rect 5260 3650 5280 3690
rect 5320 3650 5340 3690
rect 6240 3690 6680 3710
rect 6240 3670 6440 3690
rect 5260 3630 5340 3650
rect 6420 3650 6440 3670
rect 6480 3670 6680 3690
rect 7580 3690 7660 3710
rect 6480 3650 6500 3670
rect 6420 3630 6500 3650
rect 7580 3650 7600 3690
rect 7640 3650 7660 3690
rect 7580 3630 7660 3650
rect 8000 3620 8040 3750
rect 2010 3560 2450 3610
rect 4860 3600 4940 3620
rect 4860 3560 4880 3600
rect 4920 3560 4940 3600
rect 4860 3540 4940 3560
rect 5540 3540 5620 3620
rect 6120 3600 6200 3620
rect 6120 3560 6140 3600
rect 6180 3560 6200 3600
rect 6120 3540 6200 3560
rect 6720 3600 6800 3620
rect 6720 3560 6740 3600
rect 6780 3560 6800 3600
rect 6720 3540 6800 3560
rect 7300 3540 7380 3620
rect 7980 3600 8060 3620
rect 7980 3560 8000 3600
rect 8040 3560 8060 3600
rect 7980 3540 8060 3560
rect 3790 3430 4230 3490
rect 6420 3510 6500 3530
rect 6420 3470 6440 3510
rect 6480 3470 6500 3510
rect 6420 3450 6500 3470
rect 8880 3440 8920 3750
rect 9010 3680 9050 3750
rect 8970 3660 9050 3680
rect 8970 3620 8990 3660
rect 9030 3620 9050 3660
rect 8970 3600 9050 3620
rect 3790 3390 3810 3430
rect 3850 3390 3900 3430
rect 3940 3390 3990 3430
rect 4030 3390 4080 3430
rect 4120 3390 4170 3430
rect 4210 3390 4230 3430
rect 3790 3370 4230 3390
rect 5540 3420 5620 3440
rect 5540 3380 5560 3420
rect 5600 3380 5620 3420
rect 5540 3360 5620 3380
rect 5940 3420 6020 3440
rect 5940 3380 5960 3420
rect 6000 3380 6020 3420
rect 5940 3360 6020 3380
rect 6060 3420 6140 3440
rect 6060 3380 6080 3420
rect 6120 3380 6140 3420
rect 6060 3360 6140 3380
rect 6780 3420 6860 3440
rect 6780 3380 6800 3420
rect 6840 3380 6860 3420
rect 6780 3360 6860 3380
rect 6900 3420 6980 3440
rect 6900 3380 6920 3420
rect 6960 3380 6980 3420
rect 6900 3360 6980 3380
rect 7300 3420 7380 3440
rect 7300 3380 7320 3420
rect 7360 3380 7380 3420
rect 7300 3360 7380 3380
rect 8860 3420 8940 3440
rect 8860 3380 8880 3420
rect 8920 3380 8940 3420
rect 8860 3360 8940 3380
rect 5560 3320 5600 3360
rect 5960 3320 6000 3360
rect 6920 3320 6960 3360
rect 7320 3320 7360 3360
rect 5060 3300 5210 3320
rect 5060 3260 5080 3300
rect 5120 3260 5160 3300
rect 5200 3260 5210 3300
rect 5060 3200 5210 3260
rect 5060 3160 5080 3200
rect 5120 3160 5160 3200
rect 5200 3160 5210 3200
rect 5060 3140 5210 3160
rect 5350 3300 5410 3320
rect 5350 3260 5360 3300
rect 5400 3260 5410 3300
rect 5350 3200 5410 3260
rect 5350 3160 5360 3200
rect 5400 3160 5410 3200
rect 5350 3140 5410 3160
rect 5550 3300 5610 3320
rect 5550 3260 5560 3300
rect 5600 3260 5610 3300
rect 5550 3200 5610 3260
rect 5550 3160 5560 3200
rect 5600 3160 5610 3200
rect 5550 3140 5610 3160
rect 5750 3300 5810 3320
rect 5750 3260 5760 3300
rect 5800 3260 5810 3300
rect 5750 3200 5810 3260
rect 5750 3160 5760 3200
rect 5800 3160 5810 3200
rect 5750 3140 5810 3160
rect 5950 3300 6010 3320
rect 5950 3260 5960 3300
rect 6000 3260 6010 3300
rect 5950 3200 6010 3260
rect 5950 3160 5960 3200
rect 6000 3160 6010 3200
rect 5950 3140 6010 3160
rect 6150 3300 6210 3320
rect 6150 3260 6160 3300
rect 6200 3260 6210 3300
rect 6150 3200 6210 3260
rect 6150 3160 6160 3200
rect 6200 3160 6210 3200
rect 6150 3140 6210 3160
rect 6350 3300 6570 3320
rect 6350 3260 6360 3300
rect 6400 3260 6440 3300
rect 6480 3260 6520 3300
rect 6560 3260 6570 3300
rect 6350 3200 6570 3260
rect 6350 3160 6360 3200
rect 6400 3160 6440 3200
rect 6480 3160 6520 3200
rect 6560 3160 6570 3200
rect 6350 3140 6570 3160
rect 6710 3300 6770 3320
rect 6710 3260 6720 3300
rect 6760 3260 6770 3300
rect 6710 3200 6770 3260
rect 6710 3160 6720 3200
rect 6760 3160 6770 3200
rect 6710 3140 6770 3160
rect 6910 3300 6970 3320
rect 6910 3260 6920 3300
rect 6960 3260 6970 3300
rect 6910 3200 6970 3260
rect 6910 3160 6920 3200
rect 6960 3160 6970 3200
rect 6910 3140 6970 3160
rect 7110 3300 7170 3320
rect 7110 3260 7120 3300
rect 7160 3260 7170 3300
rect 7110 3200 7170 3260
rect 7110 3160 7120 3200
rect 7160 3160 7170 3200
rect 7110 3140 7170 3160
rect 7310 3300 7370 3320
rect 7310 3260 7320 3300
rect 7360 3260 7370 3300
rect 7310 3200 7370 3260
rect 7310 3160 7320 3200
rect 7360 3160 7370 3200
rect 7310 3140 7370 3160
rect 7510 3300 7570 3320
rect 7510 3260 7520 3300
rect 7560 3260 7570 3300
rect 7510 3200 7570 3260
rect 7510 3160 7520 3200
rect 7560 3160 7570 3200
rect 7510 3140 7570 3160
rect 7710 3300 7850 3320
rect 7710 3260 7720 3300
rect 7760 3260 7800 3300
rect 7840 3260 7850 3300
rect 7710 3200 7850 3260
rect 7710 3160 7720 3200
rect 7760 3160 7800 3200
rect 7840 3160 7850 3200
rect 7710 3140 7850 3160
rect 1890 3070 2010 3090
rect 1890 3030 1910 3070
rect 1950 3030 2010 3070
rect 1890 3020 2010 3030
rect 3590 3070 4230 3090
rect 3590 3030 3810 3070
rect 3850 3030 3900 3070
rect 3940 3030 3990 3070
rect 4030 3030 4080 3070
rect 4120 3030 4170 3070
rect 4210 3030 4230 3070
rect 3590 3020 4230 3030
rect 1890 3010 1970 3020
rect 3790 2970 4230 3020
rect 5160 3010 5200 3140
rect 5360 3010 5400 3140
rect 5540 3080 5620 3100
rect 5540 3040 5560 3080
rect 5600 3040 5620 3080
rect 5540 3020 5620 3040
rect 5760 3010 5800 3140
rect 6160 3010 6200 3140
rect 6360 3010 6400 3140
rect 6520 3010 6560 3140
rect 6720 3010 6760 3140
rect 7120 3010 7160 3140
rect 7300 3080 7380 3100
rect 7300 3040 7320 3080
rect 7360 3040 7380 3080
rect 7300 3020 7380 3040
rect 7520 3010 7560 3140
rect 7720 3010 7760 3140
rect 5140 2990 5220 3010
rect 5140 2950 5160 2990
rect 5200 2950 5220 2990
rect 5140 2930 5220 2950
rect 5340 2990 5420 3010
rect 5340 2950 5360 2990
rect 5400 2950 5420 2990
rect 5340 2930 5420 2950
rect 5740 2990 5820 3010
rect 5740 2950 5760 2990
rect 5800 2950 5820 2990
rect 5740 2930 5820 2950
rect 6140 2990 6220 3010
rect 6140 2950 6160 2990
rect 6200 2950 6220 2990
rect 6140 2930 6220 2950
rect 6340 2990 6420 3010
rect 6340 2950 6360 2990
rect 6400 2950 6420 2990
rect 6340 2930 6420 2950
rect 6500 2990 6580 3010
rect 6500 2950 6520 2990
rect 6560 2950 6580 2990
rect 6500 2930 6580 2950
rect 6700 2990 6780 3010
rect 6700 2950 6720 2990
rect 6760 2950 6780 2990
rect 6700 2930 6780 2950
rect 7100 2990 7180 3010
rect 7100 2950 7120 2990
rect 7160 2950 7180 2990
rect 7100 2930 7180 2950
rect 7500 2990 7580 3010
rect 7500 2950 7520 2990
rect 7560 2950 7580 2990
rect 7500 2930 7580 2950
rect 7700 2990 7780 3010
rect 7700 2950 7720 2990
rect 7760 2950 7780 2990
rect 7700 2930 7780 2950
rect 2010 2850 2450 2900
rect 5760 2890 5800 2930
rect 6160 2890 6200 2930
rect 5620 2870 7380 2890
rect 5620 2830 5640 2870
rect 5680 2830 5720 2870
rect 5760 2830 5800 2870
rect 5840 2830 5880 2870
rect 5920 2830 5960 2870
rect 6000 2830 6040 2870
rect 6080 2830 6120 2870
rect 6160 2830 6200 2870
rect 6240 2830 6280 2870
rect 6320 2830 6360 2870
rect 6400 2830 6440 2870
rect 6480 2830 6520 2870
rect 6560 2830 6600 2870
rect 6640 2830 6680 2870
rect 6720 2830 6760 2870
rect 6800 2830 6840 2870
rect 6880 2830 6920 2870
rect 6960 2830 7000 2870
rect 7040 2830 7080 2870
rect 7120 2830 7160 2870
rect 7200 2830 7240 2870
rect 7280 2830 7320 2870
rect 7360 2830 7380 2870
rect 5620 2810 7380 2830
rect 3790 2730 4230 2780
rect 4590 2750 4730 2770
rect 4590 2710 4600 2750
rect 4640 2710 4680 2750
rect 4720 2710 4730 2750
rect 2010 2610 2450 2660
rect 4590 2650 4730 2710
rect 4590 2610 4600 2650
rect 4640 2610 4680 2650
rect 4720 2610 4730 2650
rect 1890 2490 1970 2500
rect 3790 2490 4230 2540
rect 1890 2480 2010 2490
rect 1890 2440 1910 2480
rect 1950 2440 2010 2480
rect 1890 2420 2010 2440
rect 4590 2550 4730 2610
rect 4590 2510 4600 2550
rect 4640 2510 4680 2550
rect 4720 2510 4730 2550
rect 4590 2450 4730 2510
rect 4590 2410 4600 2450
rect 4640 2410 4680 2450
rect 4720 2410 4730 2450
rect 4590 2350 4730 2410
rect 4590 2310 4600 2350
rect 4640 2310 4680 2350
rect 4720 2310 4730 2350
rect 4590 2250 4730 2310
rect 4590 2210 4600 2250
rect 4640 2210 4680 2250
rect 4720 2210 4730 2250
rect 4590 2150 4730 2210
rect 4590 2110 4600 2150
rect 4640 2110 4680 2150
rect 4720 2110 4730 2150
rect 4590 2050 4730 2110
rect 4590 2010 4600 2050
rect 4640 2010 4680 2050
rect 4720 2010 4730 2050
rect 4590 1990 4730 2010
rect 5550 2750 5610 2770
rect 5550 2710 5560 2750
rect 5600 2710 5610 2750
rect 5550 2650 5610 2710
rect 5550 2610 5560 2650
rect 5600 2610 5610 2650
rect 5550 2550 5610 2610
rect 5550 2510 5560 2550
rect 5600 2510 5610 2550
rect 5550 2450 5610 2510
rect 5550 2410 5560 2450
rect 5600 2410 5610 2450
rect 5550 2350 5610 2410
rect 5550 2310 5560 2350
rect 5600 2310 5610 2350
rect 5550 2250 5610 2310
rect 5550 2210 5560 2250
rect 5600 2210 5610 2250
rect 5550 2150 5610 2210
rect 5550 2110 5560 2150
rect 5600 2110 5610 2150
rect 5550 2050 5610 2110
rect 5550 2010 5560 2050
rect 5600 2010 5610 2050
rect 5550 1990 5610 2010
rect 6430 2750 6490 2810
rect 6430 2710 6440 2750
rect 6480 2710 6490 2750
rect 6430 2650 6490 2710
rect 6430 2610 6440 2650
rect 6480 2610 6490 2650
rect 6430 2550 6490 2610
rect 6430 2510 6440 2550
rect 6480 2510 6490 2550
rect 6430 2450 6490 2510
rect 6430 2410 6440 2450
rect 6480 2410 6490 2450
rect 6430 2350 6490 2410
rect 6430 2310 6440 2350
rect 6480 2310 6490 2350
rect 6430 2250 6490 2310
rect 6430 2210 6440 2250
rect 6480 2210 6490 2250
rect 6430 2150 6490 2210
rect 6430 2110 6440 2150
rect 6480 2110 6490 2150
rect 6430 2050 6490 2110
rect 6430 2010 6440 2050
rect 6480 2010 6490 2050
rect 6430 1990 6490 2010
rect 7310 2750 7370 2770
rect 7310 2710 7320 2750
rect 7360 2710 7370 2750
rect 7310 2650 7370 2710
rect 7310 2610 7320 2650
rect 7360 2610 7370 2650
rect 7310 2550 7370 2610
rect 7310 2510 7320 2550
rect 7360 2510 7370 2550
rect 7310 2450 7370 2510
rect 7310 2410 7320 2450
rect 7360 2410 7370 2450
rect 7310 2350 7370 2410
rect 7310 2310 7320 2350
rect 7360 2310 7370 2350
rect 7310 2250 7370 2310
rect 7310 2210 7320 2250
rect 7360 2210 7370 2250
rect 7310 2150 7370 2210
rect 7310 2110 7320 2150
rect 7360 2110 7370 2150
rect 7310 2050 7370 2110
rect 7310 2010 7320 2050
rect 7360 2010 7370 2050
rect 7310 1990 7370 2010
rect 8190 2750 8330 2770
rect 8190 2710 8200 2750
rect 8240 2710 8280 2750
rect 8320 2710 8330 2750
rect 8190 2650 8330 2710
rect 8190 2610 8200 2650
rect 8240 2610 8280 2650
rect 8320 2610 8330 2650
rect 8190 2550 8330 2610
rect 8190 2510 8200 2550
rect 8240 2510 8280 2550
rect 8320 2510 8330 2550
rect 8190 2450 8330 2510
rect 8190 2410 8200 2450
rect 8240 2410 8280 2450
rect 8320 2410 8330 2450
rect 8190 2350 8330 2410
rect 8190 2310 8200 2350
rect 8240 2310 8280 2350
rect 8320 2310 8330 2350
rect 8190 2250 8330 2310
rect 8190 2210 8200 2250
rect 8240 2210 8280 2250
rect 8320 2210 8330 2250
rect 8190 2150 8330 2210
rect 8190 2110 8200 2150
rect 8240 2110 8280 2150
rect 8320 2110 8330 2150
rect 8190 2050 8330 2110
rect 8190 2010 8200 2050
rect 8240 2010 8280 2050
rect 8320 2010 8330 2050
rect 8190 1990 8330 2010
rect 4680 1950 4720 1990
rect 5560 1950 5600 1990
rect 7320 1950 7360 1990
rect 8190 1950 8260 1990
rect 4660 1930 5620 1950
rect 4660 1890 4680 1930
rect 4720 1890 4760 1930
rect 4800 1890 4840 1930
rect 4880 1890 4920 1930
rect 4960 1890 5000 1930
rect 5040 1890 5080 1930
rect 5120 1890 5160 1930
rect 5200 1890 5240 1930
rect 5280 1890 5320 1930
rect 5360 1890 5400 1930
rect 5440 1890 5480 1930
rect 5520 1890 5560 1930
rect 5600 1890 5620 1930
rect 4660 1870 5620 1890
rect 7300 1930 8260 1950
rect 7300 1890 7320 1930
rect 7360 1890 7400 1930
rect 7440 1890 7480 1930
rect 7520 1890 7560 1930
rect 7600 1890 7640 1930
rect 7680 1890 7720 1930
rect 7760 1890 7800 1930
rect 7840 1890 7880 1930
rect 7920 1890 7960 1930
rect 8000 1890 8040 1930
rect 8080 1890 8120 1930
rect 8160 1890 8200 1930
rect 8240 1890 8260 1930
rect 7300 1870 8260 1890
rect 5380 1800 7520 1820
rect 5380 1760 5460 1800
rect 5500 1760 5620 1800
rect 5660 1760 5780 1800
rect 5820 1760 5940 1800
rect 5980 1760 6100 1800
rect 6140 1760 6260 1800
rect 6300 1760 6420 1800
rect 6460 1760 6580 1800
rect 6620 1760 6740 1800
rect 6780 1760 6900 1800
rect 6940 1760 7060 1800
rect 7100 1760 7220 1800
rect 7260 1760 7380 1800
rect 7420 1760 7460 1800
rect 7500 1760 7520 1800
rect 5380 1740 7520 1760
rect 5380 1700 5420 1740
rect 5370 1680 5430 1700
rect 5370 1640 5380 1680
rect 5420 1640 5430 1680
rect 5370 1580 5430 1640
rect 5370 1540 5380 1580
rect 5420 1540 5430 1580
rect 5370 1520 5430 1540
rect 7450 1680 7590 1700
rect 7450 1640 7460 1680
rect 7500 1640 7540 1680
rect 7580 1650 7590 1680
rect 7580 1640 7670 1650
rect 7450 1630 7670 1640
rect 7450 1590 7610 1630
rect 7650 1590 7670 1630
rect 7450 1580 7670 1590
rect 7450 1540 7460 1580
rect 7500 1540 7540 1580
rect 7580 1570 7670 1580
rect 7580 1540 7590 1570
rect 7450 1520 7590 1540
rect 10 1279 9470 1320
rect 10 1256 1506 1279
rect 10 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2866 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4226 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5586 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6946 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8306 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9470 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9470 1256
rect 10 1166 9470 1222
rect 10 1132 1410 1166
rect 1444 1132 2597 1166
rect 2631 1132 2770 1166
rect 2804 1132 3957 1166
rect 3991 1132 4130 1166
rect 4164 1132 5317 1166
rect 5351 1132 5490 1166
rect 5524 1132 6677 1166
rect 6711 1132 6850 1166
rect 6884 1132 8037 1166
rect 8071 1132 8210 1166
rect 8244 1132 9397 1166
rect 9431 1132 9470 1166
rect 10 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9470 1132
rect 10 1076 9470 1098
rect 10 1070 1410 1076
rect 10 270 260 1070
rect 1060 1042 1410 1070
rect 1444 1075 2597 1076
rect 1444 1042 1558 1075
rect 1060 1041 1558 1042
rect 1592 1070 2597 1075
rect 1592 1041 1620 1070
rect 1060 986 1620 1041
rect 2420 1056 2597 1070
rect 2420 1022 2448 1056
rect 2482 1042 2597 1056
rect 2631 1042 2770 1076
rect 2804 1075 3957 1076
rect 2804 1042 2918 1075
rect 2482 1041 2918 1042
rect 2952 1070 3957 1075
rect 2952 1041 2980 1070
rect 2482 1022 2980 1041
rect 1060 952 1410 986
rect 1444 985 1620 986
rect 1444 952 1558 985
rect 1060 951 1558 952
rect 1592 951 1620 985
rect 1060 896 1620 951
rect 1060 862 1410 896
rect 1444 895 1620 896
rect 1444 862 1558 895
rect 1060 861 1558 862
rect 1592 861 1620 895
rect 1060 806 1620 861
rect 1060 772 1410 806
rect 1444 805 1620 806
rect 1444 772 1558 805
rect 1060 771 1558 772
rect 1592 771 1620 805
rect 1060 716 1620 771
rect 1060 682 1410 716
rect 1444 715 1620 716
rect 1444 682 1558 715
rect 1060 681 1558 682
rect 1592 681 1620 715
rect 1060 626 1620 681
rect 1060 592 1410 626
rect 1444 625 1620 626
rect 1444 592 1558 625
rect 1060 591 1558 592
rect 1592 591 1620 625
rect 1060 536 1620 591
rect 1060 502 1410 536
rect 1444 535 1620 536
rect 1444 502 1558 535
rect 1060 501 1558 502
rect 1592 501 1620 535
rect 1060 446 1620 501
rect 1060 412 1410 446
rect 1444 445 1620 446
rect 1444 412 1558 445
rect 1060 411 1558 412
rect 1592 411 1620 445
rect 1060 356 1620 411
rect 1060 322 1410 356
rect 1444 355 1620 356
rect 1444 322 1558 355
rect 1060 321 1558 322
rect 1592 321 1620 355
rect 1673 958 2367 1017
rect 1673 924 1734 958
rect 1768 930 1824 958
rect 1858 930 1914 958
rect 1948 930 2004 958
rect 1780 924 1824 930
rect 1880 924 1914 930
rect 1980 924 2004 930
rect 2038 930 2094 958
rect 2038 924 2046 930
rect 1673 896 1746 924
rect 1780 896 1846 924
rect 1880 896 1946 924
rect 1980 896 2046 924
rect 2080 924 2094 930
rect 2128 930 2184 958
rect 2128 924 2146 930
rect 2080 896 2146 924
rect 2180 924 2184 930
rect 2218 930 2274 958
rect 2218 924 2246 930
rect 2308 924 2367 958
rect 2180 896 2246 924
rect 2280 896 2367 924
rect 1673 868 2367 896
rect 1673 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2367 868
rect 1673 830 2367 834
rect 1673 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2367 830
rect 1673 778 2367 796
rect 1673 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2367 778
rect 1673 730 2367 744
rect 1673 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2367 730
rect 1673 688 2367 696
rect 1673 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2367 688
rect 1673 630 2367 654
rect 1673 598 1746 630
rect 1780 598 1846 630
rect 1880 598 1946 630
rect 1980 598 2046 630
rect 1673 564 1734 598
rect 1780 596 1824 598
rect 1880 596 1914 598
rect 1980 596 2004 598
rect 1768 564 1824 596
rect 1858 564 1914 596
rect 1948 564 2004 596
rect 2038 596 2046 598
rect 2080 598 2146 630
rect 2080 596 2094 598
rect 2038 564 2094 596
rect 2128 596 2146 598
rect 2180 598 2246 630
rect 2280 598 2367 630
rect 2180 596 2184 598
rect 2128 564 2184 596
rect 2218 596 2246 598
rect 2218 564 2274 596
rect 2308 564 2367 598
rect 1673 530 2367 564
rect 1673 508 1746 530
rect 1780 508 1846 530
rect 1880 508 1946 530
rect 1980 508 2046 530
rect 1673 474 1734 508
rect 1780 496 1824 508
rect 1880 496 1914 508
rect 1980 496 2004 508
rect 1768 474 1824 496
rect 1858 474 1914 496
rect 1948 474 2004 496
rect 2038 496 2046 508
rect 2080 508 2146 530
rect 2080 496 2094 508
rect 2038 474 2094 496
rect 2128 496 2146 508
rect 2180 508 2246 530
rect 2280 508 2367 530
rect 2180 496 2184 508
rect 2128 474 2184 496
rect 2218 496 2246 508
rect 2218 474 2274 496
rect 2308 474 2367 508
rect 1673 430 2367 474
rect 1673 418 1746 430
rect 1780 418 1846 430
rect 1880 418 1946 430
rect 1980 418 2046 430
rect 1673 384 1734 418
rect 1780 396 1824 418
rect 1880 396 1914 418
rect 1980 396 2004 418
rect 1768 384 1824 396
rect 1858 384 1914 396
rect 1948 384 2004 396
rect 2038 396 2046 418
rect 2080 418 2146 430
rect 2080 396 2094 418
rect 2038 384 2094 396
rect 2128 396 2146 418
rect 2180 418 2246 430
rect 2280 418 2367 430
rect 2180 396 2184 418
rect 2128 384 2184 396
rect 2218 396 2246 418
rect 2218 384 2274 396
rect 2308 384 2367 418
rect 1673 323 2367 384
rect 2420 986 2980 1022
rect 3780 1056 3957 1070
rect 3780 1022 3808 1056
rect 3842 1042 3957 1056
rect 3991 1042 4130 1076
rect 4164 1075 5317 1076
rect 4164 1042 4278 1075
rect 3842 1041 4278 1042
rect 4312 1070 5317 1075
rect 4312 1041 4340 1070
rect 3842 1022 4340 1041
rect 2420 966 2597 986
rect 2420 932 2448 966
rect 2482 952 2597 966
rect 2631 952 2770 986
rect 2804 985 2980 986
rect 2804 952 2918 985
rect 2482 951 2918 952
rect 2952 951 2980 985
rect 2482 932 2980 951
rect 2420 896 2980 932
rect 2420 876 2597 896
rect 2420 842 2448 876
rect 2482 862 2597 876
rect 2631 862 2770 896
rect 2804 895 2980 896
rect 2804 862 2918 895
rect 2482 861 2918 862
rect 2952 861 2980 895
rect 2482 842 2980 861
rect 2420 806 2980 842
rect 2420 786 2597 806
rect 2420 752 2448 786
rect 2482 772 2597 786
rect 2631 772 2770 806
rect 2804 805 2980 806
rect 2804 772 2918 805
rect 2482 771 2918 772
rect 2952 771 2980 805
rect 2482 752 2980 771
rect 2420 716 2980 752
rect 2420 696 2597 716
rect 2420 662 2448 696
rect 2482 682 2597 696
rect 2631 682 2770 716
rect 2804 715 2980 716
rect 2804 682 2918 715
rect 2482 681 2918 682
rect 2952 681 2980 715
rect 2482 662 2980 681
rect 2420 626 2980 662
rect 2420 606 2597 626
rect 2420 572 2448 606
rect 2482 592 2597 606
rect 2631 592 2770 626
rect 2804 625 2980 626
rect 2804 592 2918 625
rect 2482 591 2918 592
rect 2952 591 2980 625
rect 2482 572 2980 591
rect 2420 536 2980 572
rect 2420 516 2597 536
rect 2420 482 2448 516
rect 2482 502 2597 516
rect 2631 502 2770 536
rect 2804 535 2980 536
rect 2804 502 2918 535
rect 2482 501 2918 502
rect 2952 501 2980 535
rect 2482 482 2980 501
rect 2420 446 2980 482
rect 2420 426 2597 446
rect 2420 392 2448 426
rect 2482 412 2597 426
rect 2631 412 2770 446
rect 2804 445 2980 446
rect 2804 412 2918 445
rect 2482 411 2918 412
rect 2952 411 2980 445
rect 2482 392 2980 411
rect 2420 356 2980 392
rect 2420 336 2597 356
rect 1060 270 1620 321
rect 2420 302 2448 336
rect 2482 322 2597 336
rect 2631 322 2770 356
rect 2804 355 2980 356
rect 2804 322 2918 355
rect 2482 321 2918 322
rect 2952 321 2980 355
rect 3033 958 3727 1017
rect 3033 924 3094 958
rect 3128 930 3184 958
rect 3218 930 3274 958
rect 3308 930 3364 958
rect 3140 924 3184 930
rect 3240 924 3274 930
rect 3340 924 3364 930
rect 3398 930 3454 958
rect 3398 924 3406 930
rect 3033 896 3106 924
rect 3140 896 3206 924
rect 3240 896 3306 924
rect 3340 896 3406 924
rect 3440 924 3454 930
rect 3488 930 3544 958
rect 3488 924 3506 930
rect 3440 896 3506 924
rect 3540 924 3544 930
rect 3578 930 3634 958
rect 3578 924 3606 930
rect 3668 924 3727 958
rect 3540 896 3606 924
rect 3640 896 3727 924
rect 3033 868 3727 896
rect 3033 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3727 868
rect 3033 830 3727 834
rect 3033 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3727 830
rect 3033 778 3727 796
rect 3033 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3727 778
rect 3033 730 3727 744
rect 3033 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3727 730
rect 3033 688 3727 696
rect 3033 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3727 688
rect 3033 630 3727 654
rect 3033 598 3106 630
rect 3140 598 3206 630
rect 3240 598 3306 630
rect 3340 598 3406 630
rect 3033 564 3094 598
rect 3140 596 3184 598
rect 3240 596 3274 598
rect 3340 596 3364 598
rect 3128 564 3184 596
rect 3218 564 3274 596
rect 3308 564 3364 596
rect 3398 596 3406 598
rect 3440 598 3506 630
rect 3440 596 3454 598
rect 3398 564 3454 596
rect 3488 596 3506 598
rect 3540 598 3606 630
rect 3640 598 3727 630
rect 3540 596 3544 598
rect 3488 564 3544 596
rect 3578 596 3606 598
rect 3578 564 3634 596
rect 3668 564 3727 598
rect 3033 530 3727 564
rect 3033 508 3106 530
rect 3140 508 3206 530
rect 3240 508 3306 530
rect 3340 508 3406 530
rect 3033 474 3094 508
rect 3140 496 3184 508
rect 3240 496 3274 508
rect 3340 496 3364 508
rect 3128 474 3184 496
rect 3218 474 3274 496
rect 3308 474 3364 496
rect 3398 496 3406 508
rect 3440 508 3506 530
rect 3440 496 3454 508
rect 3398 474 3454 496
rect 3488 496 3506 508
rect 3540 508 3606 530
rect 3640 508 3727 530
rect 3540 496 3544 508
rect 3488 474 3544 496
rect 3578 496 3606 508
rect 3578 474 3634 496
rect 3668 474 3727 508
rect 3033 430 3727 474
rect 3033 418 3106 430
rect 3140 418 3206 430
rect 3240 418 3306 430
rect 3340 418 3406 430
rect 3033 384 3094 418
rect 3140 396 3184 418
rect 3240 396 3274 418
rect 3340 396 3364 418
rect 3128 384 3184 396
rect 3218 384 3274 396
rect 3308 384 3364 396
rect 3398 396 3406 418
rect 3440 418 3506 430
rect 3440 396 3454 418
rect 3398 384 3454 396
rect 3488 396 3506 418
rect 3540 418 3606 430
rect 3640 418 3727 430
rect 3540 396 3544 418
rect 3488 384 3544 396
rect 3578 396 3606 418
rect 3578 384 3634 396
rect 3668 384 3727 418
rect 3033 323 3727 384
rect 3780 986 4340 1022
rect 5140 1056 5317 1070
rect 5140 1022 5168 1056
rect 5202 1042 5317 1056
rect 5351 1042 5490 1076
rect 5524 1075 6677 1076
rect 5524 1042 5638 1075
rect 5202 1041 5638 1042
rect 5672 1070 6677 1075
rect 5672 1041 5700 1070
rect 5202 1022 5700 1041
rect 3780 966 3957 986
rect 3780 932 3808 966
rect 3842 952 3957 966
rect 3991 952 4130 986
rect 4164 985 4340 986
rect 4164 952 4278 985
rect 3842 951 4278 952
rect 4312 951 4340 985
rect 3842 932 4340 951
rect 3780 896 4340 932
rect 3780 876 3957 896
rect 3780 842 3808 876
rect 3842 862 3957 876
rect 3991 862 4130 896
rect 4164 895 4340 896
rect 4164 862 4278 895
rect 3842 861 4278 862
rect 4312 861 4340 895
rect 3842 842 4340 861
rect 3780 806 4340 842
rect 3780 786 3957 806
rect 3780 752 3808 786
rect 3842 772 3957 786
rect 3991 772 4130 806
rect 4164 805 4340 806
rect 4164 772 4278 805
rect 3842 771 4278 772
rect 4312 771 4340 805
rect 3842 752 4340 771
rect 3780 716 4340 752
rect 3780 696 3957 716
rect 3780 662 3808 696
rect 3842 682 3957 696
rect 3991 682 4130 716
rect 4164 715 4340 716
rect 4164 682 4278 715
rect 3842 681 4278 682
rect 4312 681 4340 715
rect 3842 662 4340 681
rect 3780 626 4340 662
rect 3780 606 3957 626
rect 3780 572 3808 606
rect 3842 592 3957 606
rect 3991 592 4130 626
rect 4164 625 4340 626
rect 4164 592 4278 625
rect 3842 591 4278 592
rect 4312 591 4340 625
rect 3842 572 4340 591
rect 3780 536 4340 572
rect 3780 516 3957 536
rect 3780 482 3808 516
rect 3842 502 3957 516
rect 3991 502 4130 536
rect 4164 535 4340 536
rect 4164 502 4278 535
rect 3842 501 4278 502
rect 4312 501 4340 535
rect 3842 482 4340 501
rect 3780 446 4340 482
rect 3780 426 3957 446
rect 3780 392 3808 426
rect 3842 412 3957 426
rect 3991 412 4130 446
rect 4164 445 4340 446
rect 4164 412 4278 445
rect 3842 411 4278 412
rect 4312 411 4340 445
rect 3842 392 4340 411
rect 3780 356 4340 392
rect 3780 336 3957 356
rect 2482 302 2980 321
rect 2420 270 2980 302
rect 3780 302 3808 336
rect 3842 322 3957 336
rect 3991 322 4130 356
rect 4164 355 4340 356
rect 4164 322 4278 355
rect 3842 321 4278 322
rect 4312 321 4340 355
rect 4393 958 5087 1017
rect 4393 924 4454 958
rect 4488 930 4544 958
rect 4578 930 4634 958
rect 4668 930 4724 958
rect 4500 924 4544 930
rect 4600 924 4634 930
rect 4700 924 4724 930
rect 4758 930 4814 958
rect 4758 924 4766 930
rect 4393 896 4466 924
rect 4500 896 4566 924
rect 4600 896 4666 924
rect 4700 896 4766 924
rect 4800 924 4814 930
rect 4848 930 4904 958
rect 4848 924 4866 930
rect 4800 896 4866 924
rect 4900 924 4904 930
rect 4938 930 4994 958
rect 4938 924 4966 930
rect 5028 924 5087 958
rect 4900 896 4966 924
rect 5000 896 5087 924
rect 4393 868 5087 896
rect 4393 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5087 868
rect 4393 830 5087 834
rect 4393 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5087 830
rect 4393 778 5087 796
rect 4393 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5087 778
rect 4393 730 5087 744
rect 4393 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5087 730
rect 4393 688 5087 696
rect 4393 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5087 688
rect 4393 630 5087 654
rect 4393 598 4466 630
rect 4500 598 4566 630
rect 4600 598 4666 630
rect 4700 598 4766 630
rect 4393 564 4454 598
rect 4500 596 4544 598
rect 4600 596 4634 598
rect 4700 596 4724 598
rect 4488 564 4544 596
rect 4578 564 4634 596
rect 4668 564 4724 596
rect 4758 596 4766 598
rect 4800 598 4866 630
rect 4800 596 4814 598
rect 4758 564 4814 596
rect 4848 596 4866 598
rect 4900 598 4966 630
rect 5000 598 5087 630
rect 4900 596 4904 598
rect 4848 564 4904 596
rect 4938 596 4966 598
rect 4938 564 4994 596
rect 5028 564 5087 598
rect 4393 530 5087 564
rect 4393 508 4466 530
rect 4500 508 4566 530
rect 4600 508 4666 530
rect 4700 508 4766 530
rect 4393 474 4454 508
rect 4500 496 4544 508
rect 4600 496 4634 508
rect 4700 496 4724 508
rect 4488 474 4544 496
rect 4578 474 4634 496
rect 4668 474 4724 496
rect 4758 496 4766 508
rect 4800 508 4866 530
rect 4800 496 4814 508
rect 4758 474 4814 496
rect 4848 496 4866 508
rect 4900 508 4966 530
rect 5000 508 5087 530
rect 4900 496 4904 508
rect 4848 474 4904 496
rect 4938 496 4966 508
rect 4938 474 4994 496
rect 5028 474 5087 508
rect 4393 430 5087 474
rect 4393 418 4466 430
rect 4500 418 4566 430
rect 4600 418 4666 430
rect 4700 418 4766 430
rect 4393 384 4454 418
rect 4500 396 4544 418
rect 4600 396 4634 418
rect 4700 396 4724 418
rect 4488 384 4544 396
rect 4578 384 4634 396
rect 4668 384 4724 396
rect 4758 396 4766 418
rect 4800 418 4866 430
rect 4800 396 4814 418
rect 4758 384 4814 396
rect 4848 396 4866 418
rect 4900 418 4966 430
rect 5000 418 5087 430
rect 4900 396 4904 418
rect 4848 384 4904 396
rect 4938 396 4966 418
rect 4938 384 4994 396
rect 5028 384 5087 418
rect 4393 323 5087 384
rect 5140 986 5700 1022
rect 6500 1056 6677 1070
rect 6500 1022 6528 1056
rect 6562 1042 6677 1056
rect 6711 1042 6850 1076
rect 6884 1075 8037 1076
rect 6884 1042 6998 1075
rect 6562 1041 6998 1042
rect 7032 1070 8037 1075
rect 7032 1041 7060 1070
rect 6562 1022 7060 1041
rect 5140 966 5317 986
rect 5140 932 5168 966
rect 5202 952 5317 966
rect 5351 952 5490 986
rect 5524 985 5700 986
rect 5524 952 5638 985
rect 5202 951 5638 952
rect 5672 951 5700 985
rect 5202 932 5700 951
rect 5140 896 5700 932
rect 5140 876 5317 896
rect 5140 842 5168 876
rect 5202 862 5317 876
rect 5351 862 5490 896
rect 5524 895 5700 896
rect 5524 862 5638 895
rect 5202 861 5638 862
rect 5672 861 5700 895
rect 5202 842 5700 861
rect 5140 806 5700 842
rect 5140 786 5317 806
rect 5140 752 5168 786
rect 5202 772 5317 786
rect 5351 772 5490 806
rect 5524 805 5700 806
rect 5524 772 5638 805
rect 5202 771 5638 772
rect 5672 771 5700 805
rect 5202 752 5700 771
rect 5140 716 5700 752
rect 5140 696 5317 716
rect 5140 662 5168 696
rect 5202 682 5317 696
rect 5351 682 5490 716
rect 5524 715 5700 716
rect 5524 682 5638 715
rect 5202 681 5638 682
rect 5672 681 5700 715
rect 5202 662 5700 681
rect 5140 626 5700 662
rect 5140 606 5317 626
rect 5140 572 5168 606
rect 5202 592 5317 606
rect 5351 592 5490 626
rect 5524 625 5700 626
rect 5524 592 5638 625
rect 5202 591 5638 592
rect 5672 591 5700 625
rect 5202 572 5700 591
rect 5140 536 5700 572
rect 5140 516 5317 536
rect 5140 482 5168 516
rect 5202 502 5317 516
rect 5351 502 5490 536
rect 5524 535 5700 536
rect 5524 502 5638 535
rect 5202 501 5638 502
rect 5672 501 5700 535
rect 5202 482 5700 501
rect 5140 446 5700 482
rect 5140 426 5317 446
rect 5140 392 5168 426
rect 5202 412 5317 426
rect 5351 412 5490 446
rect 5524 445 5700 446
rect 5524 412 5638 445
rect 5202 411 5638 412
rect 5672 411 5700 445
rect 5202 392 5700 411
rect 5140 356 5700 392
rect 5140 336 5317 356
rect 3842 302 4340 321
rect 3780 270 4340 302
rect 5140 302 5168 336
rect 5202 322 5317 336
rect 5351 322 5490 356
rect 5524 355 5700 356
rect 5524 322 5638 355
rect 5202 321 5638 322
rect 5672 321 5700 355
rect 5753 958 6447 1017
rect 5753 924 5814 958
rect 5848 930 5904 958
rect 5938 930 5994 958
rect 6028 930 6084 958
rect 5860 924 5904 930
rect 5960 924 5994 930
rect 6060 924 6084 930
rect 6118 930 6174 958
rect 6118 924 6126 930
rect 5753 896 5826 924
rect 5860 896 5926 924
rect 5960 896 6026 924
rect 6060 896 6126 924
rect 6160 924 6174 930
rect 6208 930 6264 958
rect 6208 924 6226 930
rect 6160 896 6226 924
rect 6260 924 6264 930
rect 6298 930 6354 958
rect 6298 924 6326 930
rect 6388 924 6447 958
rect 6260 896 6326 924
rect 6360 896 6447 924
rect 5753 868 6447 896
rect 5753 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6447 868
rect 5753 830 6447 834
rect 5753 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6447 830
rect 5753 778 6447 796
rect 5753 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6447 778
rect 5753 730 6447 744
rect 5753 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6447 730
rect 5753 688 6447 696
rect 5753 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6447 688
rect 5753 630 6447 654
rect 5753 598 5826 630
rect 5860 598 5926 630
rect 5960 598 6026 630
rect 6060 598 6126 630
rect 5753 564 5814 598
rect 5860 596 5904 598
rect 5960 596 5994 598
rect 6060 596 6084 598
rect 5848 564 5904 596
rect 5938 564 5994 596
rect 6028 564 6084 596
rect 6118 596 6126 598
rect 6160 598 6226 630
rect 6160 596 6174 598
rect 6118 564 6174 596
rect 6208 596 6226 598
rect 6260 598 6326 630
rect 6360 598 6447 630
rect 6260 596 6264 598
rect 6208 564 6264 596
rect 6298 596 6326 598
rect 6298 564 6354 596
rect 6388 564 6447 598
rect 5753 530 6447 564
rect 5753 508 5826 530
rect 5860 508 5926 530
rect 5960 508 6026 530
rect 6060 508 6126 530
rect 5753 474 5814 508
rect 5860 496 5904 508
rect 5960 496 5994 508
rect 6060 496 6084 508
rect 5848 474 5904 496
rect 5938 474 5994 496
rect 6028 474 6084 496
rect 6118 496 6126 508
rect 6160 508 6226 530
rect 6160 496 6174 508
rect 6118 474 6174 496
rect 6208 496 6226 508
rect 6260 508 6326 530
rect 6360 508 6447 530
rect 6260 496 6264 508
rect 6208 474 6264 496
rect 6298 496 6326 508
rect 6298 474 6354 496
rect 6388 474 6447 508
rect 5753 430 6447 474
rect 5753 418 5826 430
rect 5860 418 5926 430
rect 5960 418 6026 430
rect 6060 418 6126 430
rect 5753 384 5814 418
rect 5860 396 5904 418
rect 5960 396 5994 418
rect 6060 396 6084 418
rect 5848 384 5904 396
rect 5938 384 5994 396
rect 6028 384 6084 396
rect 6118 396 6126 418
rect 6160 418 6226 430
rect 6160 396 6174 418
rect 6118 384 6174 396
rect 6208 396 6226 418
rect 6260 418 6326 430
rect 6360 418 6447 430
rect 6260 396 6264 418
rect 6208 384 6264 396
rect 6298 396 6326 418
rect 6298 384 6354 396
rect 6388 384 6447 418
rect 5753 323 6447 384
rect 6500 986 7060 1022
rect 7860 1056 8037 1070
rect 7860 1022 7888 1056
rect 7922 1042 8037 1056
rect 8071 1042 8210 1076
rect 8244 1075 9397 1076
rect 8244 1042 8358 1075
rect 7922 1041 8358 1042
rect 8392 1070 9397 1075
rect 8392 1041 8420 1070
rect 7922 1022 8420 1041
rect 6500 966 6677 986
rect 6500 932 6528 966
rect 6562 952 6677 966
rect 6711 952 6850 986
rect 6884 985 7060 986
rect 6884 952 6998 985
rect 6562 951 6998 952
rect 7032 951 7060 985
rect 6562 932 7060 951
rect 6500 896 7060 932
rect 6500 876 6677 896
rect 6500 842 6528 876
rect 6562 862 6677 876
rect 6711 862 6850 896
rect 6884 895 7060 896
rect 6884 862 6998 895
rect 6562 861 6998 862
rect 7032 861 7060 895
rect 6562 842 7060 861
rect 6500 806 7060 842
rect 6500 786 6677 806
rect 6500 752 6528 786
rect 6562 772 6677 786
rect 6711 772 6850 806
rect 6884 805 7060 806
rect 6884 772 6998 805
rect 6562 771 6998 772
rect 7032 771 7060 805
rect 6562 752 7060 771
rect 6500 716 7060 752
rect 6500 696 6677 716
rect 6500 662 6528 696
rect 6562 682 6677 696
rect 6711 682 6850 716
rect 6884 715 7060 716
rect 6884 682 6998 715
rect 6562 681 6998 682
rect 7032 681 7060 715
rect 6562 662 7060 681
rect 6500 626 7060 662
rect 6500 606 6677 626
rect 6500 572 6528 606
rect 6562 592 6677 606
rect 6711 592 6850 626
rect 6884 625 7060 626
rect 6884 592 6998 625
rect 6562 591 6998 592
rect 7032 591 7060 625
rect 6562 572 7060 591
rect 6500 536 7060 572
rect 6500 516 6677 536
rect 6500 482 6528 516
rect 6562 502 6677 516
rect 6711 502 6850 536
rect 6884 535 7060 536
rect 6884 502 6998 535
rect 6562 501 6998 502
rect 7032 501 7060 535
rect 6562 482 7060 501
rect 6500 446 7060 482
rect 6500 426 6677 446
rect 6500 392 6528 426
rect 6562 412 6677 426
rect 6711 412 6850 446
rect 6884 445 7060 446
rect 6884 412 6998 445
rect 6562 411 6998 412
rect 7032 411 7060 445
rect 6562 392 7060 411
rect 6500 356 7060 392
rect 6500 336 6677 356
rect 5202 302 5700 321
rect 5140 270 5700 302
rect 6500 302 6528 336
rect 6562 322 6677 336
rect 6711 322 6850 356
rect 6884 355 7060 356
rect 6884 322 6998 355
rect 6562 321 6998 322
rect 7032 321 7060 355
rect 7113 958 7807 1017
rect 7113 924 7174 958
rect 7208 930 7264 958
rect 7298 930 7354 958
rect 7388 930 7444 958
rect 7220 924 7264 930
rect 7320 924 7354 930
rect 7420 924 7444 930
rect 7478 930 7534 958
rect 7478 924 7486 930
rect 7113 896 7186 924
rect 7220 896 7286 924
rect 7320 896 7386 924
rect 7420 896 7486 924
rect 7520 924 7534 930
rect 7568 930 7624 958
rect 7568 924 7586 930
rect 7520 896 7586 924
rect 7620 924 7624 930
rect 7658 930 7714 958
rect 7658 924 7686 930
rect 7748 924 7807 958
rect 7620 896 7686 924
rect 7720 896 7807 924
rect 7113 868 7807 896
rect 7113 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7807 868
rect 7113 830 7807 834
rect 7113 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7807 830
rect 7113 778 7807 796
rect 7113 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7807 778
rect 7113 730 7807 744
rect 7113 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7807 730
rect 7113 688 7807 696
rect 7113 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7807 688
rect 7113 630 7807 654
rect 7113 598 7186 630
rect 7220 598 7286 630
rect 7320 598 7386 630
rect 7420 598 7486 630
rect 7113 564 7174 598
rect 7220 596 7264 598
rect 7320 596 7354 598
rect 7420 596 7444 598
rect 7208 564 7264 596
rect 7298 564 7354 596
rect 7388 564 7444 596
rect 7478 596 7486 598
rect 7520 598 7586 630
rect 7520 596 7534 598
rect 7478 564 7534 596
rect 7568 596 7586 598
rect 7620 598 7686 630
rect 7720 598 7807 630
rect 7620 596 7624 598
rect 7568 564 7624 596
rect 7658 596 7686 598
rect 7658 564 7714 596
rect 7748 564 7807 598
rect 7113 530 7807 564
rect 7113 508 7186 530
rect 7220 508 7286 530
rect 7320 508 7386 530
rect 7420 508 7486 530
rect 7113 474 7174 508
rect 7220 496 7264 508
rect 7320 496 7354 508
rect 7420 496 7444 508
rect 7208 474 7264 496
rect 7298 474 7354 496
rect 7388 474 7444 496
rect 7478 496 7486 508
rect 7520 508 7586 530
rect 7520 496 7534 508
rect 7478 474 7534 496
rect 7568 496 7586 508
rect 7620 508 7686 530
rect 7720 508 7807 530
rect 7620 496 7624 508
rect 7568 474 7624 496
rect 7658 496 7686 508
rect 7658 474 7714 496
rect 7748 474 7807 508
rect 7113 430 7807 474
rect 7113 418 7186 430
rect 7220 418 7286 430
rect 7320 418 7386 430
rect 7420 418 7486 430
rect 7113 384 7174 418
rect 7220 396 7264 418
rect 7320 396 7354 418
rect 7420 396 7444 418
rect 7208 384 7264 396
rect 7298 384 7354 396
rect 7388 384 7444 396
rect 7478 396 7486 418
rect 7520 418 7586 430
rect 7520 396 7534 418
rect 7478 384 7534 396
rect 7568 396 7586 418
rect 7620 418 7686 430
rect 7720 418 7807 430
rect 7620 396 7624 418
rect 7568 384 7624 396
rect 7658 396 7686 418
rect 7658 384 7714 396
rect 7748 384 7807 418
rect 7113 323 7807 384
rect 7860 986 8420 1022
rect 9220 1056 9397 1070
rect 9220 1022 9248 1056
rect 9282 1042 9397 1056
rect 9431 1042 9470 1076
rect 9282 1022 9470 1042
rect 7860 966 8037 986
rect 7860 932 7888 966
rect 7922 952 8037 966
rect 8071 952 8210 986
rect 8244 985 8420 986
rect 8244 952 8358 985
rect 7922 951 8358 952
rect 8392 951 8420 985
rect 7922 932 8420 951
rect 7860 896 8420 932
rect 7860 876 8037 896
rect 7860 842 7888 876
rect 7922 862 8037 876
rect 8071 862 8210 896
rect 8244 895 8420 896
rect 8244 862 8358 895
rect 7922 861 8358 862
rect 8392 861 8420 895
rect 7922 842 8420 861
rect 7860 806 8420 842
rect 7860 786 8037 806
rect 7860 752 7888 786
rect 7922 772 8037 786
rect 8071 772 8210 806
rect 8244 805 8420 806
rect 8244 772 8358 805
rect 7922 771 8358 772
rect 8392 771 8420 805
rect 7922 752 8420 771
rect 7860 716 8420 752
rect 7860 696 8037 716
rect 7860 662 7888 696
rect 7922 682 8037 696
rect 8071 682 8210 716
rect 8244 715 8420 716
rect 8244 682 8358 715
rect 7922 681 8358 682
rect 8392 681 8420 715
rect 7922 662 8420 681
rect 7860 626 8420 662
rect 7860 606 8037 626
rect 7860 572 7888 606
rect 7922 592 8037 606
rect 8071 592 8210 626
rect 8244 625 8420 626
rect 8244 592 8358 625
rect 7922 591 8358 592
rect 8392 591 8420 625
rect 7922 572 8420 591
rect 7860 536 8420 572
rect 7860 516 8037 536
rect 7860 482 7888 516
rect 7922 502 8037 516
rect 8071 502 8210 536
rect 8244 535 8420 536
rect 8244 502 8358 535
rect 7922 501 8358 502
rect 8392 501 8420 535
rect 7922 482 8420 501
rect 7860 446 8420 482
rect 7860 426 8037 446
rect 7860 392 7888 426
rect 7922 412 8037 426
rect 8071 412 8210 446
rect 8244 445 8420 446
rect 8244 412 8358 445
rect 7922 411 8358 412
rect 8392 411 8420 445
rect 7922 392 8420 411
rect 7860 356 8420 392
rect 7860 336 8037 356
rect 6562 302 7060 321
rect 6500 270 7060 302
rect 7860 302 7888 336
rect 7922 322 8037 336
rect 8071 322 8210 356
rect 8244 355 8420 356
rect 8244 322 8358 355
rect 7922 321 8358 322
rect 8392 321 8420 355
rect 8473 958 9167 1017
rect 8473 924 8534 958
rect 8568 930 8624 958
rect 8658 930 8714 958
rect 8748 930 8804 958
rect 8580 924 8624 930
rect 8680 924 8714 930
rect 8780 924 8804 930
rect 8838 930 8894 958
rect 8838 924 8846 930
rect 8473 896 8546 924
rect 8580 896 8646 924
rect 8680 896 8746 924
rect 8780 896 8846 924
rect 8880 924 8894 930
rect 8928 930 8984 958
rect 8928 924 8946 930
rect 8880 896 8946 924
rect 8980 924 8984 930
rect 9018 930 9074 958
rect 9018 924 9046 930
rect 9108 924 9167 958
rect 8980 896 9046 924
rect 9080 896 9167 924
rect 8473 868 9167 896
rect 8473 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9167 868
rect 8473 830 9167 834
rect 8473 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9167 830
rect 8473 778 9167 796
rect 8473 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9167 778
rect 8473 730 9167 744
rect 8473 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9167 730
rect 8473 688 9167 696
rect 8473 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9167 688
rect 8473 630 9167 654
rect 8473 598 8546 630
rect 8580 598 8646 630
rect 8680 598 8746 630
rect 8780 598 8846 630
rect 8473 564 8534 598
rect 8580 596 8624 598
rect 8680 596 8714 598
rect 8780 596 8804 598
rect 8568 564 8624 596
rect 8658 564 8714 596
rect 8748 564 8804 596
rect 8838 596 8846 598
rect 8880 598 8946 630
rect 8880 596 8894 598
rect 8838 564 8894 596
rect 8928 596 8946 598
rect 8980 598 9046 630
rect 9080 598 9167 630
rect 8980 596 8984 598
rect 8928 564 8984 596
rect 9018 596 9046 598
rect 9018 564 9074 596
rect 9108 564 9167 598
rect 8473 530 9167 564
rect 8473 508 8546 530
rect 8580 508 8646 530
rect 8680 508 8746 530
rect 8780 508 8846 530
rect 8473 474 8534 508
rect 8580 496 8624 508
rect 8680 496 8714 508
rect 8780 496 8804 508
rect 8568 474 8624 496
rect 8658 474 8714 496
rect 8748 474 8804 496
rect 8838 496 8846 508
rect 8880 508 8946 530
rect 8880 496 8894 508
rect 8838 474 8894 496
rect 8928 496 8946 508
rect 8980 508 9046 530
rect 9080 508 9167 530
rect 8980 496 8984 508
rect 8928 474 8984 496
rect 9018 496 9046 508
rect 9018 474 9074 496
rect 9108 474 9167 508
rect 8473 430 9167 474
rect 8473 418 8546 430
rect 8580 418 8646 430
rect 8680 418 8746 430
rect 8780 418 8846 430
rect 8473 384 8534 418
rect 8580 396 8624 418
rect 8680 396 8714 418
rect 8780 396 8804 418
rect 8568 384 8624 396
rect 8658 384 8714 396
rect 8748 384 8804 396
rect 8838 396 8846 418
rect 8880 418 8946 430
rect 8880 396 8894 418
rect 8838 384 8894 396
rect 8928 396 8946 418
rect 8980 418 9046 430
rect 9080 418 9167 430
rect 8980 396 8984 418
rect 8928 384 8984 396
rect 9018 396 9046 418
rect 9018 384 9074 396
rect 9108 384 9167 418
rect 8473 323 9167 384
rect 9220 986 9470 1022
rect 9220 966 9397 986
rect 9220 932 9248 966
rect 9282 952 9397 966
rect 9431 952 9470 986
rect 9282 932 9470 952
rect 9220 896 9470 932
rect 9220 876 9397 896
rect 9220 842 9248 876
rect 9282 862 9397 876
rect 9431 862 9470 896
rect 9282 842 9470 862
rect 9220 806 9470 842
rect 9220 786 9397 806
rect 9220 752 9248 786
rect 9282 772 9397 786
rect 9431 772 9470 806
rect 9282 752 9470 772
rect 9220 716 9470 752
rect 9220 696 9397 716
rect 9220 662 9248 696
rect 9282 682 9397 696
rect 9431 682 9470 716
rect 9282 662 9470 682
rect 9220 626 9470 662
rect 9220 606 9397 626
rect 9220 572 9248 606
rect 9282 592 9397 606
rect 9431 592 9470 626
rect 9282 572 9470 592
rect 9220 536 9470 572
rect 9220 516 9397 536
rect 9220 482 9248 516
rect 9282 502 9397 516
rect 9431 502 9470 536
rect 9282 482 9470 502
rect 9220 446 9470 482
rect 9220 426 9397 446
rect 9220 392 9248 426
rect 9282 412 9397 426
rect 9431 412 9470 446
rect 9282 392 9470 412
rect 9220 356 9470 392
rect 9220 336 9397 356
rect 7922 302 8420 321
rect 7860 270 8420 302
rect 9220 302 9248 336
rect 9282 322 9397 336
rect 9431 322 9470 356
rect 9282 302 9470 322
rect 9220 270 9470 302
rect 10 266 9470 270
rect 10 232 1410 266
rect 1444 242 2597 266
rect 1444 232 1636 242
rect 10 208 1636 232
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 232 2597 242
rect 2631 232 2770 266
rect 2804 242 3957 266
rect 2804 232 2996 242
rect 2390 208 2996 232
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 232 3957 242
rect 3991 232 4130 266
rect 4164 242 5317 266
rect 4164 232 4356 242
rect 3750 208 4356 232
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 232 5317 242
rect 5351 232 5490 266
rect 5524 242 6677 266
rect 5524 232 5716 242
rect 5110 208 5716 232
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 232 6677 242
rect 6711 232 6850 266
rect 6884 242 8037 266
rect 6884 232 7076 242
rect 6470 208 7076 232
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 232 8037 242
rect 8071 232 8210 266
rect 8244 242 9397 266
rect 8244 232 8436 242
rect 7830 208 8436 232
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 232 9397 242
rect 9431 232 9470 266
rect 9190 208 9470 232
rect 10 176 9470 208
rect 10 142 1410 176
rect 1444 142 2597 176
rect 2631 142 2770 176
rect 2804 142 3957 176
rect 3991 142 4130 176
rect 4164 142 5317 176
rect 5351 142 5490 176
rect 5524 142 6677 176
rect 6711 142 6850 176
rect 6884 142 8037 176
rect 8071 142 8210 176
rect 8244 142 9397 176
rect 9431 142 9470 176
rect 10 92 9470 142
rect 10 90 1506 92
rect 1540 90 1596 92
rect 1630 90 1686 92
rect 1720 90 1776 92
rect 1810 90 1866 92
rect 1900 90 1956 92
rect 1990 90 2046 92
rect 2080 90 2136 92
rect 2170 90 2226 92
rect 2260 90 2316 92
rect 2350 90 2406 92
rect 2440 90 2496 92
rect 2530 90 2866 92
rect 2900 90 2956 92
rect 2990 90 3046 92
rect 3080 90 3136 92
rect 3170 90 3226 92
rect 3260 90 3316 92
rect 3350 90 3406 92
rect 3440 90 3496 92
rect 3530 90 3586 92
rect 3620 90 3676 92
rect 3710 90 3766 92
rect 3800 90 3856 92
rect 3890 90 4226 92
rect 4260 90 4316 92
rect 4350 90 4406 92
rect 4440 90 4496 92
rect 4530 90 4586 92
rect 4620 90 4676 92
rect 4710 90 4766 92
rect 4800 90 4856 92
rect 4890 90 4946 92
rect 4980 90 5036 92
rect 5070 90 5126 92
rect 5160 90 5216 92
rect 5250 90 5586 92
rect 5620 90 5676 92
rect 5710 90 5766 92
rect 5800 90 5856 92
rect 5890 90 5946 92
rect 5980 90 6036 92
rect 6070 90 6126 92
rect 6160 90 6216 92
rect 6250 90 6306 92
rect 6340 90 6396 92
rect 6430 90 6486 92
rect 6520 90 6576 92
rect 6610 90 6946 92
rect 6980 90 7036 92
rect 7070 90 7126 92
rect 7160 90 7216 92
rect 7250 90 7306 92
rect 7340 90 7396 92
rect 7430 90 7486 92
rect 7520 90 7576 92
rect 7610 90 7666 92
rect 7700 90 7756 92
rect 7790 90 7846 92
rect 7880 90 7936 92
rect 7970 90 8306 92
rect 8340 90 8396 92
rect 8430 90 8486 92
rect 8520 90 8576 92
rect 8610 90 8666 92
rect 8700 90 8756 92
rect 8790 90 8846 92
rect 8880 90 8936 92
rect 8970 90 9026 92
rect 9060 90 9116 92
rect 9150 90 9206 92
rect 9240 90 9296 92
rect 9330 90 9470 92
rect 10 50 40 90
rect 80 50 140 90
rect 180 50 240 90
rect 280 50 330 90
rect 370 50 410 90
rect 450 50 500 90
rect 540 50 590 90
rect 630 50 680 90
rect 720 50 770 90
rect 810 50 860 90
rect 900 50 950 90
rect 990 50 1040 90
rect 1080 50 1130 90
rect 1170 50 1230 90
rect 1270 50 1320 90
rect 1360 50 1420 90
rect 1460 50 1500 90
rect 1540 50 1590 90
rect 1630 50 1680 90
rect 1720 50 1770 90
rect 1810 50 1860 90
rect 1900 50 1950 90
rect 1990 50 2040 90
rect 2080 50 2130 90
rect 2170 50 2220 90
rect 2260 50 2310 90
rect 2350 50 2400 90
rect 2440 50 2490 90
rect 2530 50 2590 90
rect 2630 50 2680 90
rect 2720 50 2770 90
rect 2810 50 2860 90
rect 2900 50 2950 90
rect 2990 50 3040 90
rect 3080 50 3130 90
rect 3170 50 3220 90
rect 3260 50 3310 90
rect 3350 50 3400 90
rect 3440 50 3490 90
rect 3530 50 3580 90
rect 3620 50 3670 90
rect 3710 50 3760 90
rect 3800 50 3850 90
rect 3890 50 3950 90
rect 3990 50 4040 90
rect 4080 50 4130 90
rect 4170 50 4220 90
rect 4260 50 4310 90
rect 4350 50 4400 90
rect 4440 50 4490 90
rect 4530 50 4580 90
rect 4620 50 4670 90
rect 4710 50 4760 90
rect 4800 50 4850 90
rect 4890 50 4940 90
rect 4980 50 5030 90
rect 5070 50 5120 90
rect 5160 50 5210 90
rect 5250 50 5310 90
rect 5350 50 5400 90
rect 5440 50 5490 90
rect 5530 50 5580 90
rect 5620 50 5670 90
rect 5710 50 5760 90
rect 5800 50 5850 90
rect 5890 50 5940 90
rect 5980 50 6030 90
rect 6070 50 6120 90
rect 6160 50 6210 90
rect 6250 50 6300 90
rect 6340 50 6390 90
rect 6430 50 6480 90
rect 6520 50 6570 90
rect 6610 50 6660 90
rect 6700 50 6760 90
rect 6800 50 6850 90
rect 6890 50 6940 90
rect 6980 50 7030 90
rect 7070 50 7120 90
rect 7160 50 7210 90
rect 7250 50 7300 90
rect 7340 50 7390 90
rect 7430 50 7480 90
rect 7520 50 7570 90
rect 7610 50 7660 90
rect 7700 50 7750 90
rect 7790 50 7840 90
rect 7880 50 7930 90
rect 7970 50 8020 90
rect 8060 50 8120 90
rect 8160 50 8210 90
rect 8250 50 8300 90
rect 8340 50 8390 90
rect 8430 50 8480 90
rect 8520 50 8570 90
rect 8610 50 8660 90
rect 8700 50 8750 90
rect 8790 50 8840 90
rect 8880 50 8930 90
rect 8970 50 9020 90
rect 9060 50 9110 90
rect 9150 50 9200 90
rect 9240 50 9290 90
rect 9330 50 9390 90
rect 9430 50 9470 90
rect 10 20 9470 50
<< viali >>
rect 4640 5500 4680 5540
rect 5040 5500 5080 5540
rect 5440 5500 5480 5540
rect 5840 5500 5880 5540
rect 6240 5500 6280 5540
rect 6440 5500 6480 5540
rect 6640 5500 6680 5540
rect 7040 5500 7080 5540
rect 7440 5500 7480 5540
rect 7840 5500 7880 5540
rect 8240 5500 8280 5540
rect 1910 4980 1950 5020
rect 4840 4560 4880 4600
rect 5240 4470 5280 4510
rect 6240 4560 6280 4600
rect 6040 4470 6080 4510
rect 6640 4560 6680 4600
rect 6840 4560 6880 4600
rect 7640 4560 7680 4600
rect 8160 4560 8200 4600
rect 8040 4470 8080 4510
rect 3810 4390 3850 4430
rect 3900 4390 3940 4430
rect 3990 4390 4030 4430
rect 4080 4390 4120 4430
rect 4170 4390 4210 4430
rect 5640 4380 5680 4420
rect 6440 4380 6480 4420
rect 7240 4380 7280 4420
rect 8770 4290 8810 4330
rect 4480 4190 4520 4230
rect 4680 4190 4720 4230
rect 5080 4190 5120 4230
rect 5480 4190 5520 4230
rect 5680 4190 5720 4230
rect 5840 4190 5880 4230
rect 6040 4190 6080 4230
rect 6240 4190 6280 4230
rect 6440 4190 6480 4230
rect 6640 4190 6680 4230
rect 6840 4190 6880 4230
rect 7040 4190 7080 4230
rect 7200 4190 7240 4230
rect 7400 4190 7440 4230
rect 7800 4190 7840 4230
rect 8200 4190 8240 4230
rect 8400 4190 8440 4230
rect 9170 4190 9210 4230
rect 1910 3980 1950 4020
rect 5280 3650 5320 3690
rect 6440 3650 6480 3690
rect 7600 3650 7640 3690
rect 4880 3560 4920 3600
rect 6140 3560 6180 3600
rect 6740 3560 6780 3600
rect 8000 3560 8040 3600
rect 6440 3470 6480 3510
rect 8990 3620 9030 3660
rect 3810 3390 3850 3430
rect 3900 3390 3940 3430
rect 3990 3390 4030 3430
rect 4080 3390 4120 3430
rect 4170 3390 4210 3430
rect 5560 3380 5600 3420
rect 5960 3380 6000 3420
rect 6080 3380 6120 3420
rect 6800 3380 6840 3420
rect 6920 3380 6960 3420
rect 7320 3380 7360 3420
rect 8880 3380 8920 3420
rect 1910 3030 1950 3070
rect 3810 3030 3850 3070
rect 3900 3030 3940 3070
rect 3990 3030 4030 3070
rect 4080 3030 4120 3070
rect 4170 3030 4210 3070
rect 5560 3040 5600 3080
rect 7320 3040 7360 3080
rect 5160 2950 5200 2990
rect 5360 2950 5400 2990
rect 5760 2950 5800 2990
rect 6160 2950 6200 2990
rect 6360 2950 6400 2990
rect 6520 2950 6560 2990
rect 6720 2950 6760 2990
rect 7120 2950 7160 2990
rect 7520 2950 7560 2990
rect 7720 2950 7760 2990
rect 7320 2830 7360 2870
rect 1910 2440 1950 2480
rect 4680 1890 4720 1930
rect 4760 1890 4800 1930
rect 4840 1890 4880 1930
rect 4920 1890 4960 1930
rect 5000 1890 5040 1930
rect 5080 1890 5120 1930
rect 5160 1890 5200 1930
rect 5240 1890 5280 1930
rect 5320 1890 5360 1930
rect 5400 1890 5440 1930
rect 5480 1890 5520 1930
rect 5560 1890 5600 1930
rect 7320 1890 7360 1930
rect 7400 1890 7440 1930
rect 7480 1890 7520 1930
rect 7560 1890 7600 1930
rect 7640 1890 7680 1930
rect 7720 1890 7760 1930
rect 7800 1890 7840 1930
rect 7880 1890 7920 1930
rect 7960 1890 8000 1930
rect 8040 1890 8080 1930
rect 8120 1890 8160 1930
rect 8200 1890 8240 1930
rect 7460 1760 7500 1800
rect 7610 1590 7650 1630
rect 1746 924 1768 930
rect 1768 924 1780 930
rect 1846 924 1858 930
rect 1858 924 1880 930
rect 1946 924 1948 930
rect 1948 924 1980 930
rect 1746 896 1780 924
rect 1846 896 1880 924
rect 1946 896 1980 924
rect 2046 896 2080 930
rect 2146 896 2180 930
rect 2246 924 2274 930
rect 2274 924 2280 930
rect 2246 896 2280 924
rect 1746 796 1780 830
rect 1846 796 1880 830
rect 1946 796 1980 830
rect 2046 796 2080 830
rect 2146 796 2180 830
rect 2246 796 2280 830
rect 1746 696 1780 730
rect 1846 696 1880 730
rect 1946 696 1980 730
rect 2046 696 2080 730
rect 2146 696 2180 730
rect 2246 696 2280 730
rect 1746 598 1780 630
rect 1846 598 1880 630
rect 1946 598 1980 630
rect 1746 596 1768 598
rect 1768 596 1780 598
rect 1846 596 1858 598
rect 1858 596 1880 598
rect 1946 596 1948 598
rect 1948 596 1980 598
rect 2046 596 2080 630
rect 2146 596 2180 630
rect 2246 598 2280 630
rect 2246 596 2274 598
rect 2274 596 2280 598
rect 1746 508 1780 530
rect 1846 508 1880 530
rect 1946 508 1980 530
rect 1746 496 1768 508
rect 1768 496 1780 508
rect 1846 496 1858 508
rect 1858 496 1880 508
rect 1946 496 1948 508
rect 1948 496 1980 508
rect 2046 496 2080 530
rect 2146 496 2180 530
rect 2246 508 2280 530
rect 2246 496 2274 508
rect 2274 496 2280 508
rect 1746 418 1780 430
rect 1846 418 1880 430
rect 1946 418 1980 430
rect 1746 396 1768 418
rect 1768 396 1780 418
rect 1846 396 1858 418
rect 1858 396 1880 418
rect 1946 396 1948 418
rect 1948 396 1980 418
rect 2046 396 2080 430
rect 2146 396 2180 430
rect 2246 418 2280 430
rect 2246 396 2274 418
rect 2274 396 2280 418
rect 3106 924 3128 930
rect 3128 924 3140 930
rect 3206 924 3218 930
rect 3218 924 3240 930
rect 3306 924 3308 930
rect 3308 924 3340 930
rect 3106 896 3140 924
rect 3206 896 3240 924
rect 3306 896 3340 924
rect 3406 896 3440 930
rect 3506 896 3540 930
rect 3606 924 3634 930
rect 3634 924 3640 930
rect 3606 896 3640 924
rect 3106 796 3140 830
rect 3206 796 3240 830
rect 3306 796 3340 830
rect 3406 796 3440 830
rect 3506 796 3540 830
rect 3606 796 3640 830
rect 3106 696 3140 730
rect 3206 696 3240 730
rect 3306 696 3340 730
rect 3406 696 3440 730
rect 3506 696 3540 730
rect 3606 696 3640 730
rect 3106 598 3140 630
rect 3206 598 3240 630
rect 3306 598 3340 630
rect 3106 596 3128 598
rect 3128 596 3140 598
rect 3206 596 3218 598
rect 3218 596 3240 598
rect 3306 596 3308 598
rect 3308 596 3340 598
rect 3406 596 3440 630
rect 3506 596 3540 630
rect 3606 598 3640 630
rect 3606 596 3634 598
rect 3634 596 3640 598
rect 3106 508 3140 530
rect 3206 508 3240 530
rect 3306 508 3340 530
rect 3106 496 3128 508
rect 3128 496 3140 508
rect 3206 496 3218 508
rect 3218 496 3240 508
rect 3306 496 3308 508
rect 3308 496 3340 508
rect 3406 496 3440 530
rect 3506 496 3540 530
rect 3606 508 3640 530
rect 3606 496 3634 508
rect 3634 496 3640 508
rect 3106 418 3140 430
rect 3206 418 3240 430
rect 3306 418 3340 430
rect 3106 396 3128 418
rect 3128 396 3140 418
rect 3206 396 3218 418
rect 3218 396 3240 418
rect 3306 396 3308 418
rect 3308 396 3340 418
rect 3406 396 3440 430
rect 3506 396 3540 430
rect 3606 418 3640 430
rect 3606 396 3634 418
rect 3634 396 3640 418
rect 4466 924 4488 930
rect 4488 924 4500 930
rect 4566 924 4578 930
rect 4578 924 4600 930
rect 4666 924 4668 930
rect 4668 924 4700 930
rect 4466 896 4500 924
rect 4566 896 4600 924
rect 4666 896 4700 924
rect 4766 896 4800 930
rect 4866 896 4900 930
rect 4966 924 4994 930
rect 4994 924 5000 930
rect 4966 896 5000 924
rect 4466 796 4500 830
rect 4566 796 4600 830
rect 4666 796 4700 830
rect 4766 796 4800 830
rect 4866 796 4900 830
rect 4966 796 5000 830
rect 4466 696 4500 730
rect 4566 696 4600 730
rect 4666 696 4700 730
rect 4766 696 4800 730
rect 4866 696 4900 730
rect 4966 696 5000 730
rect 4466 598 4500 630
rect 4566 598 4600 630
rect 4666 598 4700 630
rect 4466 596 4488 598
rect 4488 596 4500 598
rect 4566 596 4578 598
rect 4578 596 4600 598
rect 4666 596 4668 598
rect 4668 596 4700 598
rect 4766 596 4800 630
rect 4866 596 4900 630
rect 4966 598 5000 630
rect 4966 596 4994 598
rect 4994 596 5000 598
rect 4466 508 4500 530
rect 4566 508 4600 530
rect 4666 508 4700 530
rect 4466 496 4488 508
rect 4488 496 4500 508
rect 4566 496 4578 508
rect 4578 496 4600 508
rect 4666 496 4668 508
rect 4668 496 4700 508
rect 4766 496 4800 530
rect 4866 496 4900 530
rect 4966 508 5000 530
rect 4966 496 4994 508
rect 4994 496 5000 508
rect 4466 418 4500 430
rect 4566 418 4600 430
rect 4666 418 4700 430
rect 4466 396 4488 418
rect 4488 396 4500 418
rect 4566 396 4578 418
rect 4578 396 4600 418
rect 4666 396 4668 418
rect 4668 396 4700 418
rect 4766 396 4800 430
rect 4866 396 4900 430
rect 4966 418 5000 430
rect 4966 396 4994 418
rect 4994 396 5000 418
rect 5826 924 5848 930
rect 5848 924 5860 930
rect 5926 924 5938 930
rect 5938 924 5960 930
rect 6026 924 6028 930
rect 6028 924 6060 930
rect 5826 896 5860 924
rect 5926 896 5960 924
rect 6026 896 6060 924
rect 6126 896 6160 930
rect 6226 896 6260 930
rect 6326 924 6354 930
rect 6354 924 6360 930
rect 6326 896 6360 924
rect 5826 796 5860 830
rect 5926 796 5960 830
rect 6026 796 6060 830
rect 6126 796 6160 830
rect 6226 796 6260 830
rect 6326 796 6360 830
rect 5826 696 5860 730
rect 5926 696 5960 730
rect 6026 696 6060 730
rect 6126 696 6160 730
rect 6226 696 6260 730
rect 6326 696 6360 730
rect 5826 598 5860 630
rect 5926 598 5960 630
rect 6026 598 6060 630
rect 5826 596 5848 598
rect 5848 596 5860 598
rect 5926 596 5938 598
rect 5938 596 5960 598
rect 6026 596 6028 598
rect 6028 596 6060 598
rect 6126 596 6160 630
rect 6226 596 6260 630
rect 6326 598 6360 630
rect 6326 596 6354 598
rect 6354 596 6360 598
rect 5826 508 5860 530
rect 5926 508 5960 530
rect 6026 508 6060 530
rect 5826 496 5848 508
rect 5848 496 5860 508
rect 5926 496 5938 508
rect 5938 496 5960 508
rect 6026 496 6028 508
rect 6028 496 6060 508
rect 6126 496 6160 530
rect 6226 496 6260 530
rect 6326 508 6360 530
rect 6326 496 6354 508
rect 6354 496 6360 508
rect 5826 418 5860 430
rect 5926 418 5960 430
rect 6026 418 6060 430
rect 5826 396 5848 418
rect 5848 396 5860 418
rect 5926 396 5938 418
rect 5938 396 5960 418
rect 6026 396 6028 418
rect 6028 396 6060 418
rect 6126 396 6160 430
rect 6226 396 6260 430
rect 6326 418 6360 430
rect 6326 396 6354 418
rect 6354 396 6360 418
rect 7186 924 7208 930
rect 7208 924 7220 930
rect 7286 924 7298 930
rect 7298 924 7320 930
rect 7386 924 7388 930
rect 7388 924 7420 930
rect 7186 896 7220 924
rect 7286 896 7320 924
rect 7386 896 7420 924
rect 7486 896 7520 930
rect 7586 896 7620 930
rect 7686 924 7714 930
rect 7714 924 7720 930
rect 7686 896 7720 924
rect 7186 796 7220 830
rect 7286 796 7320 830
rect 7386 796 7420 830
rect 7486 796 7520 830
rect 7586 796 7620 830
rect 7686 796 7720 830
rect 7186 696 7220 730
rect 7286 696 7320 730
rect 7386 696 7420 730
rect 7486 696 7520 730
rect 7586 696 7620 730
rect 7686 696 7720 730
rect 7186 598 7220 630
rect 7286 598 7320 630
rect 7386 598 7420 630
rect 7186 596 7208 598
rect 7208 596 7220 598
rect 7286 596 7298 598
rect 7298 596 7320 598
rect 7386 596 7388 598
rect 7388 596 7420 598
rect 7486 596 7520 630
rect 7586 596 7620 630
rect 7686 598 7720 630
rect 7686 596 7714 598
rect 7714 596 7720 598
rect 7186 508 7220 530
rect 7286 508 7320 530
rect 7386 508 7420 530
rect 7186 496 7208 508
rect 7208 496 7220 508
rect 7286 496 7298 508
rect 7298 496 7320 508
rect 7386 496 7388 508
rect 7388 496 7420 508
rect 7486 496 7520 530
rect 7586 496 7620 530
rect 7686 508 7720 530
rect 7686 496 7714 508
rect 7714 496 7720 508
rect 7186 418 7220 430
rect 7286 418 7320 430
rect 7386 418 7420 430
rect 7186 396 7208 418
rect 7208 396 7220 418
rect 7286 396 7298 418
rect 7298 396 7320 418
rect 7386 396 7388 418
rect 7388 396 7420 418
rect 7486 396 7520 430
rect 7586 396 7620 430
rect 7686 418 7720 430
rect 7686 396 7714 418
rect 7714 396 7720 418
rect 8546 924 8568 930
rect 8568 924 8580 930
rect 8646 924 8658 930
rect 8658 924 8680 930
rect 8746 924 8748 930
rect 8748 924 8780 930
rect 8546 896 8580 924
rect 8646 896 8680 924
rect 8746 896 8780 924
rect 8846 896 8880 930
rect 8946 896 8980 930
rect 9046 924 9074 930
rect 9074 924 9080 930
rect 9046 896 9080 924
rect 8546 796 8580 830
rect 8646 796 8680 830
rect 8746 796 8780 830
rect 8846 796 8880 830
rect 8946 796 8980 830
rect 9046 796 9080 830
rect 8546 696 8580 730
rect 8646 696 8680 730
rect 8746 696 8780 730
rect 8846 696 8880 730
rect 8946 696 8980 730
rect 9046 696 9080 730
rect 8546 598 8580 630
rect 8646 598 8680 630
rect 8746 598 8780 630
rect 8546 596 8568 598
rect 8568 596 8580 598
rect 8646 596 8658 598
rect 8658 596 8680 598
rect 8746 596 8748 598
rect 8748 596 8780 598
rect 8846 596 8880 630
rect 8946 596 8980 630
rect 9046 598 9080 630
rect 9046 596 9074 598
rect 9074 596 9080 598
rect 8546 508 8580 530
rect 8646 508 8680 530
rect 8746 508 8780 530
rect 8546 496 8568 508
rect 8568 496 8580 508
rect 8646 496 8658 508
rect 8658 496 8680 508
rect 8746 496 8748 508
rect 8748 496 8780 508
rect 8846 496 8880 530
rect 8946 496 8980 530
rect 9046 508 9080 530
rect 9046 496 9074 508
rect 9074 496 9080 508
rect 8546 418 8580 430
rect 8646 418 8680 430
rect 8746 418 8780 430
rect 8546 396 8568 418
rect 8568 396 8580 418
rect 8646 396 8658 418
rect 8658 396 8680 418
rect 8746 396 8748 418
rect 8748 396 8780 418
rect 8846 396 8880 430
rect 8946 396 8980 430
rect 9046 418 9080 430
rect 9046 396 9074 418
rect 9074 396 9080 418
rect 40 50 80 90
rect 140 50 180 90
rect 240 50 280 90
rect 330 50 370 90
rect 410 50 450 90
rect 500 50 540 90
rect 590 50 630 90
rect 680 50 720 90
rect 770 50 810 90
rect 860 50 900 90
rect 950 50 990 90
rect 1040 50 1080 90
rect 1130 50 1170 90
rect 1230 50 1270 90
rect 1320 50 1360 90
rect 1420 50 1460 90
rect 1500 58 1506 90
rect 1506 58 1540 90
rect 1500 50 1540 58
rect 1590 58 1596 90
rect 1596 58 1630 90
rect 1590 50 1630 58
rect 1680 58 1686 90
rect 1686 58 1720 90
rect 1680 50 1720 58
rect 1770 58 1776 90
rect 1776 58 1810 90
rect 1770 50 1810 58
rect 1860 58 1866 90
rect 1866 58 1900 90
rect 1860 50 1900 58
rect 1950 58 1956 90
rect 1956 58 1990 90
rect 1950 50 1990 58
rect 2040 58 2046 90
rect 2046 58 2080 90
rect 2040 50 2080 58
rect 2130 58 2136 90
rect 2136 58 2170 90
rect 2130 50 2170 58
rect 2220 58 2226 90
rect 2226 58 2260 90
rect 2220 50 2260 58
rect 2310 58 2316 90
rect 2316 58 2350 90
rect 2310 50 2350 58
rect 2400 58 2406 90
rect 2406 58 2440 90
rect 2400 50 2440 58
rect 2490 58 2496 90
rect 2496 58 2530 90
rect 2490 50 2530 58
rect 2590 50 2630 90
rect 2680 50 2720 90
rect 2770 50 2810 90
rect 2860 58 2866 90
rect 2866 58 2900 90
rect 2860 50 2900 58
rect 2950 58 2956 90
rect 2956 58 2990 90
rect 2950 50 2990 58
rect 3040 58 3046 90
rect 3046 58 3080 90
rect 3040 50 3080 58
rect 3130 58 3136 90
rect 3136 58 3170 90
rect 3130 50 3170 58
rect 3220 58 3226 90
rect 3226 58 3260 90
rect 3220 50 3260 58
rect 3310 58 3316 90
rect 3316 58 3350 90
rect 3310 50 3350 58
rect 3400 58 3406 90
rect 3406 58 3440 90
rect 3400 50 3440 58
rect 3490 58 3496 90
rect 3496 58 3530 90
rect 3490 50 3530 58
rect 3580 58 3586 90
rect 3586 58 3620 90
rect 3580 50 3620 58
rect 3670 58 3676 90
rect 3676 58 3710 90
rect 3670 50 3710 58
rect 3760 58 3766 90
rect 3766 58 3800 90
rect 3760 50 3800 58
rect 3850 58 3856 90
rect 3856 58 3890 90
rect 3850 50 3890 58
rect 3950 50 3990 90
rect 4040 50 4080 90
rect 4130 50 4170 90
rect 4220 58 4226 90
rect 4226 58 4260 90
rect 4220 50 4260 58
rect 4310 58 4316 90
rect 4316 58 4350 90
rect 4310 50 4350 58
rect 4400 58 4406 90
rect 4406 58 4440 90
rect 4400 50 4440 58
rect 4490 58 4496 90
rect 4496 58 4530 90
rect 4490 50 4530 58
rect 4580 58 4586 90
rect 4586 58 4620 90
rect 4580 50 4620 58
rect 4670 58 4676 90
rect 4676 58 4710 90
rect 4670 50 4710 58
rect 4760 58 4766 90
rect 4766 58 4800 90
rect 4760 50 4800 58
rect 4850 58 4856 90
rect 4856 58 4890 90
rect 4850 50 4890 58
rect 4940 58 4946 90
rect 4946 58 4980 90
rect 4940 50 4980 58
rect 5030 58 5036 90
rect 5036 58 5070 90
rect 5030 50 5070 58
rect 5120 58 5126 90
rect 5126 58 5160 90
rect 5120 50 5160 58
rect 5210 58 5216 90
rect 5216 58 5250 90
rect 5210 50 5250 58
rect 5310 50 5350 90
rect 5400 50 5440 90
rect 5490 50 5530 90
rect 5580 58 5586 90
rect 5586 58 5620 90
rect 5580 50 5620 58
rect 5670 58 5676 90
rect 5676 58 5710 90
rect 5670 50 5710 58
rect 5760 58 5766 90
rect 5766 58 5800 90
rect 5760 50 5800 58
rect 5850 58 5856 90
rect 5856 58 5890 90
rect 5850 50 5890 58
rect 5940 58 5946 90
rect 5946 58 5980 90
rect 5940 50 5980 58
rect 6030 58 6036 90
rect 6036 58 6070 90
rect 6030 50 6070 58
rect 6120 58 6126 90
rect 6126 58 6160 90
rect 6120 50 6160 58
rect 6210 58 6216 90
rect 6216 58 6250 90
rect 6210 50 6250 58
rect 6300 58 6306 90
rect 6306 58 6340 90
rect 6300 50 6340 58
rect 6390 58 6396 90
rect 6396 58 6430 90
rect 6390 50 6430 58
rect 6480 58 6486 90
rect 6486 58 6520 90
rect 6480 50 6520 58
rect 6570 58 6576 90
rect 6576 58 6610 90
rect 6570 50 6610 58
rect 6660 50 6700 90
rect 6760 50 6800 90
rect 6850 50 6890 90
rect 6940 58 6946 90
rect 6946 58 6980 90
rect 6940 50 6980 58
rect 7030 58 7036 90
rect 7036 58 7070 90
rect 7030 50 7070 58
rect 7120 58 7126 90
rect 7126 58 7160 90
rect 7120 50 7160 58
rect 7210 58 7216 90
rect 7216 58 7250 90
rect 7210 50 7250 58
rect 7300 58 7306 90
rect 7306 58 7340 90
rect 7300 50 7340 58
rect 7390 58 7396 90
rect 7396 58 7430 90
rect 7390 50 7430 58
rect 7480 58 7486 90
rect 7486 58 7520 90
rect 7480 50 7520 58
rect 7570 58 7576 90
rect 7576 58 7610 90
rect 7570 50 7610 58
rect 7660 58 7666 90
rect 7666 58 7700 90
rect 7660 50 7700 58
rect 7750 58 7756 90
rect 7756 58 7790 90
rect 7750 50 7790 58
rect 7840 58 7846 90
rect 7846 58 7880 90
rect 7840 50 7880 58
rect 7930 58 7936 90
rect 7936 58 7970 90
rect 7930 50 7970 58
rect 8020 50 8060 90
rect 8120 50 8160 90
rect 8210 50 8250 90
rect 8300 58 8306 90
rect 8306 58 8340 90
rect 8300 50 8340 58
rect 8390 58 8396 90
rect 8396 58 8430 90
rect 8390 50 8430 58
rect 8480 58 8486 90
rect 8486 58 8520 90
rect 8480 50 8520 58
rect 8570 58 8576 90
rect 8576 58 8610 90
rect 8570 50 8610 58
rect 8660 58 8666 90
rect 8666 58 8700 90
rect 8660 50 8700 58
rect 8750 58 8756 90
rect 8756 58 8790 90
rect 8750 50 8790 58
rect 8840 58 8846 90
rect 8846 58 8880 90
rect 8840 50 8880 58
rect 8930 58 8936 90
rect 8936 58 8970 90
rect 8930 50 8970 58
rect 9020 58 9026 90
rect 9026 58 9060 90
rect 9020 50 9060 58
rect 9110 58 9116 90
rect 9116 58 9150 90
rect 9110 50 9150 58
rect 9200 58 9206 90
rect 9206 58 9240 90
rect 9200 50 9240 58
rect 9290 58 9296 90
rect 9296 58 9330 90
rect 9290 50 9330 58
rect 9390 50 9430 90
<< metal1 >>
rect 6440 5560 6480 6300
rect 4620 5550 4700 5560
rect 4620 5490 4630 5550
rect 4690 5490 4700 5550
rect 4620 5480 4700 5490
rect 5020 5550 5100 5560
rect 5020 5490 5030 5550
rect 5090 5490 5100 5550
rect 5020 5480 5100 5490
rect 5420 5550 5500 5560
rect 5420 5490 5430 5550
rect 5490 5490 5500 5550
rect 5420 5480 5500 5490
rect 5820 5550 5900 5560
rect 5820 5490 5830 5550
rect 5890 5490 5900 5550
rect 5820 5480 5900 5490
rect 6220 5550 6300 5560
rect 6220 5490 6230 5550
rect 6290 5490 6300 5550
rect 6220 5480 6300 5490
rect 6420 5540 6500 5560
rect 6420 5500 6440 5540
rect 6480 5500 6500 5540
rect 6420 5480 6500 5500
rect 6620 5550 6700 5560
rect 6620 5490 6630 5550
rect 6690 5490 6700 5550
rect 6620 5480 6700 5490
rect 7020 5550 7100 5560
rect 7020 5490 7030 5550
rect 7090 5490 7100 5550
rect 7020 5480 7100 5490
rect 7420 5550 7500 5560
rect 7420 5490 7430 5550
rect 7490 5490 7500 5550
rect 7420 5480 7500 5490
rect 7820 5550 7900 5560
rect 7820 5490 7830 5550
rect 7890 5490 7900 5550
rect 7820 5480 7900 5490
rect 8220 5550 8300 5560
rect 8220 5490 8230 5550
rect 8290 5490 8300 5550
rect 8220 5480 8300 5490
rect 1890 5030 1970 5040
rect 1890 4970 1900 5030
rect 1960 4970 1970 5030
rect 1890 4960 1970 4970
rect 4300 4610 4380 4620
rect 4300 4550 4310 4610
rect 4370 4550 4380 4610
rect 4300 4540 4380 4550
rect 4820 4610 4900 4620
rect 4820 4550 4830 4610
rect 4890 4550 4900 4610
rect 4820 4540 4900 4550
rect 6220 4600 6300 4620
rect 6220 4560 6240 4600
rect 6280 4560 6300 4600
rect 6220 4540 6300 4560
rect 6620 4600 6700 4620
rect 6620 4560 6640 4600
rect 6680 4560 6700 4600
rect 6620 4540 6700 4560
rect 6820 4610 6900 4620
rect 6820 4550 6830 4610
rect 6890 4550 6900 4610
rect 6820 4540 6900 4550
rect 7620 4610 7700 4620
rect 7620 4550 7630 4610
rect 7690 4550 7700 4610
rect 7620 4540 7700 4550
rect 8140 4610 8220 4620
rect 8140 4550 8150 4610
rect 8210 4550 8220 4610
rect 8140 4540 8220 4550
rect 8750 4610 8830 4620
rect 8750 4550 8760 4610
rect 8820 4550 8830 4610
rect 8750 4540 8830 4550
rect 3790 4440 4230 4450
rect 3790 4380 3800 4440
rect 4220 4380 4230 4440
rect 3790 4370 4230 4380
rect 1890 4030 1970 4040
rect 1890 3970 1900 4030
rect 1960 3970 1970 4030
rect 1890 3960 1970 3970
rect 880 3440 960 3450
rect 880 3380 890 3440
rect 950 3380 960 3440
rect 880 1450 960 3380
rect 3790 3440 4230 3450
rect 4320 3440 4360 4540
rect 5220 4520 5300 4530
rect 5220 4460 5230 4520
rect 5290 4460 5300 4520
rect 5220 4450 5300 4460
rect 6020 4520 6100 4530
rect 6020 4460 6030 4520
rect 6090 4460 6100 4520
rect 6020 4450 6100 4460
rect 5620 4430 5700 4440
rect 5620 4370 5630 4430
rect 5690 4370 5700 4430
rect 5620 4360 5700 4370
rect 6240 4250 6280 4540
rect 6420 4430 6500 4440
rect 6420 4370 6430 4430
rect 6490 4370 6500 4430
rect 6420 4360 6500 4370
rect 6640 4250 6680 4540
rect 8020 4520 8100 4530
rect 8020 4460 8030 4520
rect 8090 4460 8100 4520
rect 8020 4450 8100 4460
rect 8630 4520 8710 4530
rect 8630 4460 8640 4520
rect 8700 4460 8710 4520
rect 8630 4450 8710 4460
rect 7220 4430 7300 4440
rect 7220 4370 7230 4430
rect 7290 4370 7300 4430
rect 7220 4360 7300 4370
rect 4460 4240 4540 4250
rect 4460 4180 4470 4240
rect 4530 4180 4540 4240
rect 4460 4170 4540 4180
rect 4660 4240 4740 4250
rect 4660 4180 4670 4240
rect 4730 4180 4740 4240
rect 4660 4170 4740 4180
rect 5060 4240 5140 4250
rect 5060 4180 5070 4240
rect 5130 4180 5140 4240
rect 5060 4170 5140 4180
rect 5460 4240 5540 4250
rect 5460 4180 5470 4240
rect 5530 4180 5540 4240
rect 5460 4170 5540 4180
rect 5660 4240 5740 4250
rect 5660 4180 5670 4240
rect 5730 4180 5740 4240
rect 5660 4170 5740 4180
rect 5820 4240 5900 4250
rect 5820 4180 5830 4240
rect 5890 4180 5900 4240
rect 5820 4170 5900 4180
rect 6020 4240 6100 4250
rect 6020 4180 6030 4240
rect 6090 4180 6100 4240
rect 6020 4170 6100 4180
rect 6220 4230 6300 4250
rect 6220 4190 6240 4230
rect 6280 4190 6300 4230
rect 6220 4170 6300 4190
rect 6420 4240 6500 4250
rect 6420 4180 6430 4240
rect 6490 4180 6500 4240
rect 6420 4170 6500 4180
rect 6620 4230 6700 4250
rect 6620 4190 6640 4230
rect 6680 4190 6700 4230
rect 6620 4170 6700 4190
rect 6820 4240 6900 4250
rect 6820 4180 6830 4240
rect 6890 4180 6900 4240
rect 6820 4170 6900 4180
rect 7020 4240 7100 4250
rect 7020 4180 7030 4240
rect 7090 4180 7100 4240
rect 7020 4170 7100 4180
rect 7180 4240 7260 4250
rect 7180 4180 7190 4240
rect 7250 4180 7260 4240
rect 7180 4170 7260 4180
rect 7380 4240 7460 4250
rect 7380 4180 7390 4240
rect 7450 4180 7460 4240
rect 7380 4170 7460 4180
rect 7780 4240 7860 4250
rect 7780 4180 7790 4240
rect 7850 4180 7860 4240
rect 7780 4170 7860 4180
rect 8180 4240 8260 4250
rect 8180 4180 8190 4240
rect 8250 4180 8260 4240
rect 8180 4170 8260 4180
rect 8380 4240 8460 4250
rect 8380 4180 8390 4240
rect 8450 4180 8460 4240
rect 8380 4170 8460 4180
rect 5260 3700 5340 3710
rect 5260 3640 5270 3700
rect 5330 3640 5340 3700
rect 5260 3630 5340 3640
rect 5940 3700 6020 3710
rect 5940 3640 5950 3700
rect 6010 3640 6020 3700
rect 5940 3630 6020 3640
rect 6420 3690 6500 3710
rect 6420 3650 6440 3690
rect 6480 3650 6500 3690
rect 6420 3630 6500 3650
rect 6900 3700 6980 3710
rect 6900 3640 6910 3700
rect 6970 3640 6980 3700
rect 6900 3630 6980 3640
rect 7580 3700 7660 3710
rect 7580 3640 7590 3700
rect 7650 3640 7660 3700
rect 7580 3630 7660 3640
rect 4860 3610 4940 3620
rect 4860 3550 4870 3610
rect 4930 3550 4940 3610
rect 4860 3540 4940 3550
rect 5540 3610 5620 3620
rect 5540 3550 5550 3610
rect 5610 3550 5620 3610
rect 5540 3540 5620 3550
rect 5560 3440 5600 3540
rect 5960 3440 6000 3630
rect 6120 3610 6200 3620
rect 6120 3550 6130 3610
rect 6190 3550 6200 3610
rect 6120 3540 6200 3550
rect 6440 3530 6480 3630
rect 6720 3610 6800 3620
rect 6720 3550 6730 3610
rect 6790 3550 6800 3610
rect 6720 3540 6800 3550
rect 6420 3520 6500 3530
rect 6420 3460 6430 3520
rect 6490 3460 6500 3520
rect 6420 3450 6500 3460
rect 6920 3440 6960 3630
rect 7300 3610 7380 3620
rect 7300 3550 7310 3610
rect 7370 3550 7380 3610
rect 7300 3540 7380 3550
rect 7980 3610 8060 3620
rect 7980 3550 7990 3610
rect 8050 3550 8060 3610
rect 7980 3540 8060 3550
rect 7320 3440 7360 3540
rect 8440 3520 8520 3530
rect 8440 3460 8450 3520
rect 8510 3460 8520 3520
rect 8440 3450 8520 3460
rect 3790 3380 3800 3440
rect 4220 3380 4230 3440
rect 3790 3370 4230 3380
rect 4300 3430 4380 3440
rect 4300 3370 4310 3430
rect 4370 3370 4380 3430
rect 4300 3360 4380 3370
rect 5540 3420 5620 3440
rect 5540 3380 5560 3420
rect 5600 3380 5620 3420
rect 5540 3360 5620 3380
rect 5940 3420 6020 3440
rect 5940 3380 5960 3420
rect 6000 3380 6020 3420
rect 5940 3360 6020 3380
rect 6060 3430 6140 3440
rect 6060 3370 6070 3430
rect 6130 3370 6140 3430
rect 6060 3360 6140 3370
rect 6780 3430 6860 3440
rect 6780 3370 6790 3430
rect 6850 3370 6860 3430
rect 6780 3360 6860 3370
rect 6900 3420 6980 3440
rect 6900 3380 6920 3420
rect 6960 3380 6980 3420
rect 6900 3360 6980 3380
rect 7300 3420 7380 3440
rect 7300 3380 7320 3420
rect 7360 3380 7380 3420
rect 7300 3360 7380 3380
rect 5540 3090 5620 3100
rect 360 370 960 1450
rect 1720 3080 1800 3090
rect 1720 3020 1730 3080
rect 1790 3020 1800 3080
rect 1720 1460 1800 3020
rect 1890 3080 1970 3090
rect 1890 3020 1900 3080
rect 1960 3020 1970 3080
rect 1890 3010 1970 3020
rect 3790 3080 4230 3090
rect 3790 3020 3800 3080
rect 4220 3020 4230 3080
rect 5540 3030 5550 3090
rect 5610 3030 5620 3090
rect 5540 3020 5620 3030
rect 7300 3090 7380 3100
rect 7300 3030 7310 3090
rect 7370 3030 7380 3090
rect 7300 3020 7380 3030
rect 3790 3010 4230 3020
rect 5140 3000 5220 3010
rect 5140 2940 5150 3000
rect 5210 2940 5220 3000
rect 5140 2930 5220 2940
rect 5340 3000 5420 3010
rect 5340 2940 5350 3000
rect 5410 2940 5420 3000
rect 5340 2930 5420 2940
rect 5740 3000 5820 3010
rect 5740 2940 5750 3000
rect 5810 2940 5820 3000
rect 5740 2930 5820 2940
rect 6140 3000 6220 3010
rect 6140 2940 6150 3000
rect 6210 2940 6220 3000
rect 6140 2930 6220 2940
rect 6340 3000 6420 3010
rect 6340 2940 6350 3000
rect 6410 2940 6420 3000
rect 6340 2930 6420 2940
rect 6500 3000 6580 3010
rect 6500 2940 6510 3000
rect 6570 2940 6580 3000
rect 6500 2930 6580 2940
rect 6700 3000 6780 3010
rect 6700 2940 6710 3000
rect 6770 2940 6780 3000
rect 6700 2930 6780 2940
rect 7100 3000 7180 3010
rect 7100 2940 7110 3000
rect 7170 2940 7180 3000
rect 7100 2930 7180 2940
rect 7500 3000 7580 3010
rect 7500 2940 7510 3000
rect 7570 2940 7580 3000
rect 7500 2930 7580 2940
rect 7700 3000 7780 3010
rect 7700 2940 7710 3000
rect 7770 2940 7780 3000
rect 7700 2930 7780 2940
rect 8460 2890 8500 3450
rect 8650 3100 8690 4450
rect 8770 4350 8810 4540
rect 8750 4330 8830 4350
rect 8750 4290 8770 4330
rect 8810 4290 8830 4330
rect 8750 4270 8830 4290
rect 9150 4240 9230 4250
rect 9150 4180 9160 4240
rect 9220 4180 9230 4240
rect 9150 4170 9230 4180
rect 8970 3660 9050 3680
rect 8970 3620 8990 3660
rect 9030 3620 9050 3660
rect 8970 3600 9050 3620
rect 8860 3430 8940 3440
rect 8860 3370 8870 3430
rect 8930 3370 8940 3430
rect 8860 3360 8940 3370
rect 8630 3090 8710 3100
rect 8630 3030 8640 3090
rect 8700 3030 8710 3090
rect 8630 3020 8710 3030
rect 7300 2880 7380 2890
rect 7300 2820 7310 2880
rect 7370 2820 7380 2880
rect 7300 2810 7380 2820
rect 8440 2880 8520 2890
rect 8440 2820 8450 2880
rect 8510 2820 8520 2880
rect 8440 2810 8520 2820
rect 1890 2490 1970 2500
rect 1890 2430 1900 2490
rect 1960 2430 1970 2490
rect 1890 2420 1970 2430
rect 4660 1940 5620 1950
rect 4660 1880 4670 1940
rect 4730 1880 4750 1940
rect 4810 1880 4830 1940
rect 4890 1880 4910 1940
rect 4970 1880 4990 1940
rect 5050 1880 5070 1940
rect 5130 1880 5150 1940
rect 5210 1880 5230 1940
rect 5290 1880 5310 1940
rect 5370 1880 5390 1940
rect 5450 1880 5470 1940
rect 5530 1880 5550 1940
rect 5610 1880 5620 1940
rect 4660 1870 5620 1880
rect 7300 1940 8260 1950
rect 7300 1880 7310 1940
rect 7370 1880 7390 1940
rect 7450 1880 7470 1940
rect 7530 1880 7550 1940
rect 7610 1880 7630 1940
rect 7690 1880 7710 1940
rect 7770 1880 7790 1940
rect 7850 1880 7870 1940
rect 7930 1880 7950 1940
rect 8010 1880 8030 1940
rect 8090 1880 8110 1940
rect 8170 1880 8190 1940
rect 8250 1880 8260 1940
rect 7300 1870 8260 1880
rect 9010 1820 9050 3600
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1750 7520 1810
rect 7440 1740 7520 1750
rect 8990 1810 9070 1820
rect 8990 1750 9000 1810
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect 7590 1640 7670 1650
rect 7590 1580 7600 1640
rect 7660 1580 7670 1640
rect 7590 1570 7670 1580
rect 1720 1380 9120 1460
rect 1720 975 2320 1380
rect 3080 975 3680 1380
rect 4440 975 5040 1380
rect 5800 975 6400 1380
rect 7160 975 7760 1380
rect 8520 975 9120 1380
rect 1715 930 2325 975
rect 1715 896 1746 930
rect 1780 896 1846 930
rect 1880 896 1946 930
rect 1980 896 2046 930
rect 2080 896 2146 930
rect 2180 896 2246 930
rect 2280 896 2325 930
rect 1715 830 2325 896
rect 1715 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2325 830
rect 1715 730 2325 796
rect 1715 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2325 730
rect 1715 630 2325 696
rect 1715 596 1746 630
rect 1780 596 1846 630
rect 1880 596 1946 630
rect 1980 596 2046 630
rect 2080 596 2146 630
rect 2180 596 2246 630
rect 2280 596 2325 630
rect 1715 530 2325 596
rect 1715 496 1746 530
rect 1780 496 1846 530
rect 1880 496 1946 530
rect 1980 496 2046 530
rect 2080 496 2146 530
rect 2180 496 2246 530
rect 2280 496 2325 530
rect 1715 430 2325 496
rect 1715 396 1746 430
rect 1780 396 1846 430
rect 1880 396 1946 430
rect 1980 396 2046 430
rect 2080 396 2146 430
rect 2180 396 2246 430
rect 2280 396 2325 430
rect 1715 365 2325 396
rect 3075 930 3685 975
rect 3075 896 3106 930
rect 3140 896 3206 930
rect 3240 896 3306 930
rect 3340 896 3406 930
rect 3440 896 3506 930
rect 3540 896 3606 930
rect 3640 896 3685 930
rect 3075 830 3685 896
rect 3075 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3685 830
rect 3075 730 3685 796
rect 3075 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3685 730
rect 3075 630 3685 696
rect 3075 596 3106 630
rect 3140 596 3206 630
rect 3240 596 3306 630
rect 3340 596 3406 630
rect 3440 596 3506 630
rect 3540 596 3606 630
rect 3640 596 3685 630
rect 3075 530 3685 596
rect 3075 496 3106 530
rect 3140 496 3206 530
rect 3240 496 3306 530
rect 3340 496 3406 530
rect 3440 496 3506 530
rect 3540 496 3606 530
rect 3640 496 3685 530
rect 3075 430 3685 496
rect 3075 396 3106 430
rect 3140 396 3206 430
rect 3240 396 3306 430
rect 3340 396 3406 430
rect 3440 396 3506 430
rect 3540 396 3606 430
rect 3640 396 3685 430
rect 3075 365 3685 396
rect 4435 930 5045 975
rect 4435 896 4466 930
rect 4500 896 4566 930
rect 4600 896 4666 930
rect 4700 896 4766 930
rect 4800 896 4866 930
rect 4900 896 4966 930
rect 5000 896 5045 930
rect 4435 830 5045 896
rect 4435 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5045 830
rect 4435 730 5045 796
rect 4435 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5045 730
rect 4435 630 5045 696
rect 4435 596 4466 630
rect 4500 596 4566 630
rect 4600 596 4666 630
rect 4700 596 4766 630
rect 4800 596 4866 630
rect 4900 596 4966 630
rect 5000 596 5045 630
rect 4435 530 5045 596
rect 4435 496 4466 530
rect 4500 496 4566 530
rect 4600 496 4666 530
rect 4700 496 4766 530
rect 4800 496 4866 530
rect 4900 496 4966 530
rect 5000 496 5045 530
rect 4435 430 5045 496
rect 4435 396 4466 430
rect 4500 396 4566 430
rect 4600 396 4666 430
rect 4700 396 4766 430
rect 4800 396 4866 430
rect 4900 396 4966 430
rect 5000 396 5045 430
rect 4435 365 5045 396
rect 5795 930 6405 975
rect 5795 896 5826 930
rect 5860 896 5926 930
rect 5960 896 6026 930
rect 6060 896 6126 930
rect 6160 896 6226 930
rect 6260 896 6326 930
rect 6360 896 6405 930
rect 5795 830 6405 896
rect 5795 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6405 830
rect 5795 730 6405 796
rect 5795 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6405 730
rect 5795 630 6405 696
rect 5795 596 5826 630
rect 5860 596 5926 630
rect 5960 596 6026 630
rect 6060 596 6126 630
rect 6160 596 6226 630
rect 6260 596 6326 630
rect 6360 596 6405 630
rect 5795 530 6405 596
rect 5795 496 5826 530
rect 5860 496 5926 530
rect 5960 496 6026 530
rect 6060 496 6126 530
rect 6160 496 6226 530
rect 6260 496 6326 530
rect 6360 496 6405 530
rect 5795 430 6405 496
rect 5795 396 5826 430
rect 5860 396 5926 430
rect 5960 396 6026 430
rect 6060 396 6126 430
rect 6160 396 6226 430
rect 6260 396 6326 430
rect 6360 396 6405 430
rect 5795 365 6405 396
rect 7155 930 7765 975
rect 7155 896 7186 930
rect 7220 896 7286 930
rect 7320 896 7386 930
rect 7420 896 7486 930
rect 7520 896 7586 930
rect 7620 896 7686 930
rect 7720 896 7765 930
rect 7155 830 7765 896
rect 7155 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7765 830
rect 7155 730 7765 796
rect 7155 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7765 730
rect 7155 630 7765 696
rect 7155 596 7186 630
rect 7220 596 7286 630
rect 7320 596 7386 630
rect 7420 596 7486 630
rect 7520 596 7586 630
rect 7620 596 7686 630
rect 7720 596 7765 630
rect 7155 530 7765 596
rect 7155 496 7186 530
rect 7220 496 7286 530
rect 7320 496 7386 530
rect 7420 496 7486 530
rect 7520 496 7586 530
rect 7620 496 7686 530
rect 7720 496 7765 530
rect 7155 430 7765 496
rect 7155 396 7186 430
rect 7220 396 7286 430
rect 7320 396 7386 430
rect 7420 396 7486 430
rect 7520 396 7586 430
rect 7620 396 7686 430
rect 7720 396 7765 430
rect 7155 365 7765 396
rect 8515 930 9125 975
rect 8515 896 8546 930
rect 8580 896 8646 930
rect 8680 896 8746 930
rect 8780 896 8846 930
rect 8880 896 8946 930
rect 8980 896 9046 930
rect 9080 896 9125 930
rect 8515 830 9125 896
rect 8515 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9125 830
rect 8515 730 9125 796
rect 8515 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9125 730
rect 8515 630 9125 696
rect 8515 596 8546 630
rect 8580 596 8646 630
rect 8680 596 8746 630
rect 8780 596 8846 630
rect 8880 596 8946 630
rect 8980 596 9046 630
rect 9080 596 9125 630
rect 8515 530 9125 596
rect 8515 496 8546 530
rect 8580 496 8646 530
rect 8680 496 8746 530
rect 8780 496 8846 530
rect 8880 496 8946 530
rect 8980 496 9046 530
rect 9080 496 9125 530
rect 8515 430 9125 496
rect 8515 396 8546 430
rect 8580 396 8646 430
rect 8680 396 8746 430
rect 8780 396 8846 430
rect 8880 396 8946 430
rect 8980 396 9046 430
rect 9080 396 9125 430
rect 8515 365 9125 396
rect 10 100 9460 120
rect 10 40 30 100
rect 90 40 130 100
rect 190 40 230 100
rect 290 40 320 100
rect 380 40 400 100
rect 460 40 490 100
rect 550 40 580 100
rect 640 40 670 100
rect 730 40 760 100
rect 820 40 850 100
rect 910 40 940 100
rect 1000 40 1030 100
rect 1090 40 1120 100
rect 1180 40 1220 100
rect 1280 40 1310 100
rect 1370 40 1410 100
rect 1470 40 1490 100
rect 1550 40 1580 100
rect 1640 40 1670 100
rect 1730 40 1760 100
rect 1820 40 1850 100
rect 1910 40 1940 100
rect 2000 40 2030 100
rect 2090 40 2120 100
rect 2180 40 2210 100
rect 2270 40 2300 100
rect 2360 40 2390 100
rect 2450 40 2480 100
rect 2540 40 2580 100
rect 2640 40 2670 100
rect 2730 40 2760 100
rect 2820 40 2850 100
rect 2910 40 2940 100
rect 3000 40 3030 100
rect 3090 40 3120 100
rect 3180 40 3210 100
rect 3270 40 3300 100
rect 3360 40 3390 100
rect 3450 40 3480 100
rect 3540 40 3570 100
rect 3630 40 3660 100
rect 3720 40 3750 100
rect 3810 40 3840 100
rect 3900 40 3940 100
rect 4000 40 4030 100
rect 4090 40 4120 100
rect 4180 40 4210 100
rect 4270 40 4300 100
rect 4360 40 4390 100
rect 4450 40 4480 100
rect 4540 40 4570 100
rect 4630 40 4660 100
rect 4720 40 4750 100
rect 4810 40 4840 100
rect 4900 40 4930 100
rect 4990 40 5020 100
rect 5080 40 5110 100
rect 5170 40 5200 100
rect 5260 40 5300 100
rect 5360 40 5390 100
rect 5450 40 5480 100
rect 5540 40 5570 100
rect 5630 40 5660 100
rect 5720 40 5750 100
rect 5810 40 5840 100
rect 5900 40 5930 100
rect 5990 40 6020 100
rect 6080 40 6110 100
rect 6170 40 6200 100
rect 6260 40 6290 100
rect 6350 40 6380 100
rect 6440 40 6470 100
rect 6530 40 6560 100
rect 6620 40 6650 100
rect 6710 40 6750 100
rect 6810 40 6840 100
rect 6900 40 6930 100
rect 6990 40 7020 100
rect 7080 40 7110 100
rect 7170 40 7200 100
rect 7260 40 7290 100
rect 7350 40 7380 100
rect 7440 40 7470 100
rect 7530 40 7560 100
rect 7620 40 7650 100
rect 7710 40 7740 100
rect 7800 40 7830 100
rect 7890 40 7920 100
rect 7980 40 8010 100
rect 8070 40 8110 100
rect 8170 40 8200 100
rect 8260 40 8290 100
rect 8350 40 8380 100
rect 8440 40 8470 100
rect 8530 40 8560 100
rect 8620 40 8650 100
rect 8710 40 8740 100
rect 8800 40 8830 100
rect 8890 40 8920 100
rect 8980 40 9010 100
rect 9070 40 9100 100
rect 9160 40 9190 100
rect 9250 40 9280 100
rect 9340 40 9380 100
rect 9440 40 9460 100
rect 10 20 9460 40
<< via1 >>
rect 4630 5540 4690 5550
rect 4630 5500 4640 5540
rect 4640 5500 4680 5540
rect 4680 5500 4690 5540
rect 4630 5490 4690 5500
rect 5030 5540 5090 5550
rect 5030 5500 5040 5540
rect 5040 5500 5080 5540
rect 5080 5500 5090 5540
rect 5030 5490 5090 5500
rect 5430 5540 5490 5550
rect 5430 5500 5440 5540
rect 5440 5500 5480 5540
rect 5480 5500 5490 5540
rect 5430 5490 5490 5500
rect 5830 5540 5890 5550
rect 5830 5500 5840 5540
rect 5840 5500 5880 5540
rect 5880 5500 5890 5540
rect 5830 5490 5890 5500
rect 6230 5540 6290 5550
rect 6230 5500 6240 5540
rect 6240 5500 6280 5540
rect 6280 5500 6290 5540
rect 6230 5490 6290 5500
rect 6630 5540 6690 5550
rect 6630 5500 6640 5540
rect 6640 5500 6680 5540
rect 6680 5500 6690 5540
rect 6630 5490 6690 5500
rect 7030 5540 7090 5550
rect 7030 5500 7040 5540
rect 7040 5500 7080 5540
rect 7080 5500 7090 5540
rect 7030 5490 7090 5500
rect 7430 5540 7490 5550
rect 7430 5500 7440 5540
rect 7440 5500 7480 5540
rect 7480 5500 7490 5540
rect 7430 5490 7490 5500
rect 7830 5540 7890 5550
rect 7830 5500 7840 5540
rect 7840 5500 7880 5540
rect 7880 5500 7890 5540
rect 7830 5490 7890 5500
rect 8230 5540 8290 5550
rect 8230 5500 8240 5540
rect 8240 5500 8280 5540
rect 8280 5500 8290 5540
rect 8230 5490 8290 5500
rect 1900 5020 1960 5030
rect 1900 4980 1910 5020
rect 1910 4980 1950 5020
rect 1950 4980 1960 5020
rect 1900 4970 1960 4980
rect 4310 4550 4370 4610
rect 4830 4600 4890 4610
rect 4830 4560 4840 4600
rect 4840 4560 4880 4600
rect 4880 4560 4890 4600
rect 4830 4550 4890 4560
rect 6830 4600 6890 4610
rect 6830 4560 6840 4600
rect 6840 4560 6880 4600
rect 6880 4560 6890 4600
rect 6830 4550 6890 4560
rect 7630 4600 7690 4610
rect 7630 4560 7640 4600
rect 7640 4560 7680 4600
rect 7680 4560 7690 4600
rect 7630 4550 7690 4560
rect 8150 4600 8210 4610
rect 8150 4560 8160 4600
rect 8160 4560 8200 4600
rect 8200 4560 8210 4600
rect 8150 4550 8210 4560
rect 8760 4550 8820 4610
rect 3800 4430 4220 4440
rect 3800 4390 3810 4430
rect 3810 4390 3850 4430
rect 3850 4390 3900 4430
rect 3900 4390 3940 4430
rect 3940 4390 3990 4430
rect 3990 4390 4030 4430
rect 4030 4390 4080 4430
rect 4080 4390 4120 4430
rect 4120 4390 4170 4430
rect 4170 4390 4210 4430
rect 4210 4390 4220 4430
rect 3800 4380 4220 4390
rect 1900 4020 1960 4030
rect 1900 3980 1910 4020
rect 1910 3980 1950 4020
rect 1950 3980 1960 4020
rect 1900 3970 1960 3980
rect 890 3380 950 3440
rect 5230 4510 5290 4520
rect 5230 4470 5240 4510
rect 5240 4470 5280 4510
rect 5280 4470 5290 4510
rect 5230 4460 5290 4470
rect 6030 4510 6090 4520
rect 6030 4470 6040 4510
rect 6040 4470 6080 4510
rect 6080 4470 6090 4510
rect 6030 4460 6090 4470
rect 5630 4420 5690 4430
rect 5630 4380 5640 4420
rect 5640 4380 5680 4420
rect 5680 4380 5690 4420
rect 5630 4370 5690 4380
rect 6430 4420 6490 4430
rect 6430 4380 6440 4420
rect 6440 4380 6480 4420
rect 6480 4380 6490 4420
rect 6430 4370 6490 4380
rect 8030 4510 8090 4520
rect 8030 4470 8040 4510
rect 8040 4470 8080 4510
rect 8080 4470 8090 4510
rect 8030 4460 8090 4470
rect 8640 4460 8700 4520
rect 7230 4420 7290 4430
rect 7230 4380 7240 4420
rect 7240 4380 7280 4420
rect 7280 4380 7290 4420
rect 7230 4370 7290 4380
rect 4470 4230 4530 4240
rect 4470 4190 4480 4230
rect 4480 4190 4520 4230
rect 4520 4190 4530 4230
rect 4470 4180 4530 4190
rect 4670 4230 4730 4240
rect 4670 4190 4680 4230
rect 4680 4190 4720 4230
rect 4720 4190 4730 4230
rect 4670 4180 4730 4190
rect 5070 4230 5130 4240
rect 5070 4190 5080 4230
rect 5080 4190 5120 4230
rect 5120 4190 5130 4230
rect 5070 4180 5130 4190
rect 5470 4230 5530 4240
rect 5470 4190 5480 4230
rect 5480 4190 5520 4230
rect 5520 4190 5530 4230
rect 5470 4180 5530 4190
rect 5670 4230 5730 4240
rect 5670 4190 5680 4230
rect 5680 4190 5720 4230
rect 5720 4190 5730 4230
rect 5670 4180 5730 4190
rect 5830 4230 5890 4240
rect 5830 4190 5840 4230
rect 5840 4190 5880 4230
rect 5880 4190 5890 4230
rect 5830 4180 5890 4190
rect 6030 4230 6090 4240
rect 6030 4190 6040 4230
rect 6040 4190 6080 4230
rect 6080 4190 6090 4230
rect 6030 4180 6090 4190
rect 6430 4230 6490 4240
rect 6430 4190 6440 4230
rect 6440 4190 6480 4230
rect 6480 4190 6490 4230
rect 6430 4180 6490 4190
rect 6830 4230 6890 4240
rect 6830 4190 6840 4230
rect 6840 4190 6880 4230
rect 6880 4190 6890 4230
rect 6830 4180 6890 4190
rect 7030 4230 7090 4240
rect 7030 4190 7040 4230
rect 7040 4190 7080 4230
rect 7080 4190 7090 4230
rect 7030 4180 7090 4190
rect 7190 4230 7250 4240
rect 7190 4190 7200 4230
rect 7200 4190 7240 4230
rect 7240 4190 7250 4230
rect 7190 4180 7250 4190
rect 7390 4230 7450 4240
rect 7390 4190 7400 4230
rect 7400 4190 7440 4230
rect 7440 4190 7450 4230
rect 7390 4180 7450 4190
rect 7790 4230 7850 4240
rect 7790 4190 7800 4230
rect 7800 4190 7840 4230
rect 7840 4190 7850 4230
rect 7790 4180 7850 4190
rect 8190 4230 8250 4240
rect 8190 4190 8200 4230
rect 8200 4190 8240 4230
rect 8240 4190 8250 4230
rect 8190 4180 8250 4190
rect 8390 4230 8450 4240
rect 8390 4190 8400 4230
rect 8400 4190 8440 4230
rect 8440 4190 8450 4230
rect 8390 4180 8450 4190
rect 5270 3690 5330 3700
rect 5270 3650 5280 3690
rect 5280 3650 5320 3690
rect 5320 3650 5330 3690
rect 5270 3640 5330 3650
rect 5950 3640 6010 3700
rect 6910 3640 6970 3700
rect 7590 3690 7650 3700
rect 7590 3650 7600 3690
rect 7600 3650 7640 3690
rect 7640 3650 7650 3690
rect 7590 3640 7650 3650
rect 4870 3600 4930 3610
rect 4870 3560 4880 3600
rect 4880 3560 4920 3600
rect 4920 3560 4930 3600
rect 4870 3550 4930 3560
rect 5550 3550 5610 3610
rect 6130 3600 6190 3610
rect 6130 3560 6140 3600
rect 6140 3560 6180 3600
rect 6180 3560 6190 3600
rect 6130 3550 6190 3560
rect 6730 3600 6790 3610
rect 6730 3560 6740 3600
rect 6740 3560 6780 3600
rect 6780 3560 6790 3600
rect 6730 3550 6790 3560
rect 6430 3510 6490 3520
rect 6430 3470 6440 3510
rect 6440 3470 6480 3510
rect 6480 3470 6490 3510
rect 6430 3460 6490 3470
rect 7310 3550 7370 3610
rect 7990 3600 8050 3610
rect 7990 3560 8000 3600
rect 8000 3560 8040 3600
rect 8040 3560 8050 3600
rect 7990 3550 8050 3560
rect 8450 3460 8510 3520
rect 3800 3430 4220 3440
rect 3800 3390 3810 3430
rect 3810 3390 3850 3430
rect 3850 3390 3900 3430
rect 3900 3390 3940 3430
rect 3940 3390 3990 3430
rect 3990 3390 4030 3430
rect 4030 3390 4080 3430
rect 4080 3390 4120 3430
rect 4120 3390 4170 3430
rect 4170 3390 4210 3430
rect 4210 3390 4220 3430
rect 3800 3380 4220 3390
rect 4310 3370 4370 3430
rect 6070 3420 6130 3430
rect 6070 3380 6080 3420
rect 6080 3380 6120 3420
rect 6120 3380 6130 3420
rect 6070 3370 6130 3380
rect 6790 3420 6850 3430
rect 6790 3380 6800 3420
rect 6800 3380 6840 3420
rect 6840 3380 6850 3420
rect 6790 3370 6850 3380
rect 1730 3020 1790 3080
rect 1900 3070 1960 3080
rect 1900 3030 1910 3070
rect 1910 3030 1950 3070
rect 1950 3030 1960 3070
rect 1900 3020 1960 3030
rect 3800 3070 4220 3080
rect 3800 3030 3810 3070
rect 3810 3030 3850 3070
rect 3850 3030 3900 3070
rect 3900 3030 3940 3070
rect 3940 3030 3990 3070
rect 3990 3030 4030 3070
rect 4030 3030 4080 3070
rect 4080 3030 4120 3070
rect 4120 3030 4170 3070
rect 4170 3030 4210 3070
rect 4210 3030 4220 3070
rect 3800 3020 4220 3030
rect 5550 3080 5610 3090
rect 5550 3040 5560 3080
rect 5560 3040 5600 3080
rect 5600 3040 5610 3080
rect 5550 3030 5610 3040
rect 7310 3080 7370 3090
rect 7310 3040 7320 3080
rect 7320 3040 7360 3080
rect 7360 3040 7370 3080
rect 7310 3030 7370 3040
rect 5150 2990 5210 3000
rect 5150 2950 5160 2990
rect 5160 2950 5200 2990
rect 5200 2950 5210 2990
rect 5150 2940 5210 2950
rect 5350 2990 5410 3000
rect 5350 2950 5360 2990
rect 5360 2950 5400 2990
rect 5400 2950 5410 2990
rect 5350 2940 5410 2950
rect 5750 2990 5810 3000
rect 5750 2950 5760 2990
rect 5760 2950 5800 2990
rect 5800 2950 5810 2990
rect 5750 2940 5810 2950
rect 6150 2990 6210 3000
rect 6150 2950 6160 2990
rect 6160 2950 6200 2990
rect 6200 2950 6210 2990
rect 6150 2940 6210 2950
rect 6350 2990 6410 3000
rect 6350 2950 6360 2990
rect 6360 2950 6400 2990
rect 6400 2950 6410 2990
rect 6350 2940 6410 2950
rect 6510 2990 6570 3000
rect 6510 2950 6520 2990
rect 6520 2950 6560 2990
rect 6560 2950 6570 2990
rect 6510 2940 6570 2950
rect 6710 2990 6770 3000
rect 6710 2950 6720 2990
rect 6720 2950 6760 2990
rect 6760 2950 6770 2990
rect 6710 2940 6770 2950
rect 7110 2990 7170 3000
rect 7110 2950 7120 2990
rect 7120 2950 7160 2990
rect 7160 2950 7170 2990
rect 7110 2940 7170 2950
rect 7510 2990 7570 3000
rect 7510 2950 7520 2990
rect 7520 2950 7560 2990
rect 7560 2950 7570 2990
rect 7510 2940 7570 2950
rect 7710 2990 7770 3000
rect 7710 2950 7720 2990
rect 7720 2950 7760 2990
rect 7760 2950 7770 2990
rect 7710 2940 7770 2950
rect 9160 4230 9220 4240
rect 9160 4190 9170 4230
rect 9170 4190 9210 4230
rect 9210 4190 9220 4230
rect 9160 4180 9220 4190
rect 8870 3420 8930 3430
rect 8870 3380 8880 3420
rect 8880 3380 8920 3420
rect 8920 3380 8930 3420
rect 8870 3370 8930 3380
rect 8640 3030 8700 3090
rect 7310 2870 7370 2880
rect 7310 2830 7320 2870
rect 7320 2830 7360 2870
rect 7360 2830 7370 2870
rect 7310 2820 7370 2830
rect 8450 2820 8510 2880
rect 1900 2480 1960 2490
rect 1900 2440 1910 2480
rect 1910 2440 1950 2480
rect 1950 2440 1960 2480
rect 1900 2430 1960 2440
rect 4670 1930 4730 1940
rect 4670 1890 4680 1930
rect 4680 1890 4720 1930
rect 4720 1890 4730 1930
rect 4670 1880 4730 1890
rect 4750 1930 4810 1940
rect 4750 1890 4760 1930
rect 4760 1890 4800 1930
rect 4800 1890 4810 1930
rect 4750 1880 4810 1890
rect 4830 1930 4890 1940
rect 4830 1890 4840 1930
rect 4840 1890 4880 1930
rect 4880 1890 4890 1930
rect 4830 1880 4890 1890
rect 4910 1930 4970 1940
rect 4910 1890 4920 1930
rect 4920 1890 4960 1930
rect 4960 1890 4970 1930
rect 4910 1880 4970 1890
rect 4990 1930 5050 1940
rect 4990 1890 5000 1930
rect 5000 1890 5040 1930
rect 5040 1890 5050 1930
rect 4990 1880 5050 1890
rect 5070 1930 5130 1940
rect 5070 1890 5080 1930
rect 5080 1890 5120 1930
rect 5120 1890 5130 1930
rect 5070 1880 5130 1890
rect 5150 1930 5210 1940
rect 5150 1890 5160 1930
rect 5160 1890 5200 1930
rect 5200 1890 5210 1930
rect 5150 1880 5210 1890
rect 5230 1930 5290 1940
rect 5230 1890 5240 1930
rect 5240 1890 5280 1930
rect 5280 1890 5290 1930
rect 5230 1880 5290 1890
rect 5310 1930 5370 1940
rect 5310 1890 5320 1930
rect 5320 1890 5360 1930
rect 5360 1890 5370 1930
rect 5310 1880 5370 1890
rect 5390 1930 5450 1940
rect 5390 1890 5400 1930
rect 5400 1890 5440 1930
rect 5440 1890 5450 1930
rect 5390 1880 5450 1890
rect 5470 1930 5530 1940
rect 5470 1890 5480 1930
rect 5480 1890 5520 1930
rect 5520 1890 5530 1930
rect 5470 1880 5530 1890
rect 5550 1930 5610 1940
rect 5550 1890 5560 1930
rect 5560 1890 5600 1930
rect 5600 1890 5610 1930
rect 5550 1880 5610 1890
rect 7310 1930 7370 1940
rect 7310 1890 7320 1930
rect 7320 1890 7360 1930
rect 7360 1890 7370 1930
rect 7310 1880 7370 1890
rect 7390 1930 7450 1940
rect 7390 1890 7400 1930
rect 7400 1890 7440 1930
rect 7440 1890 7450 1930
rect 7390 1880 7450 1890
rect 7470 1930 7530 1940
rect 7470 1890 7480 1930
rect 7480 1890 7520 1930
rect 7520 1890 7530 1930
rect 7470 1880 7530 1890
rect 7550 1930 7610 1940
rect 7550 1890 7560 1930
rect 7560 1890 7600 1930
rect 7600 1890 7610 1930
rect 7550 1880 7610 1890
rect 7630 1930 7690 1940
rect 7630 1890 7640 1930
rect 7640 1890 7680 1930
rect 7680 1890 7690 1930
rect 7630 1880 7690 1890
rect 7710 1930 7770 1940
rect 7710 1890 7720 1930
rect 7720 1890 7760 1930
rect 7760 1890 7770 1930
rect 7710 1880 7770 1890
rect 7790 1930 7850 1940
rect 7790 1890 7800 1930
rect 7800 1890 7840 1930
rect 7840 1890 7850 1930
rect 7790 1880 7850 1890
rect 7870 1930 7930 1940
rect 7870 1890 7880 1930
rect 7880 1890 7920 1930
rect 7920 1890 7930 1930
rect 7870 1880 7930 1890
rect 7950 1930 8010 1940
rect 7950 1890 7960 1930
rect 7960 1890 8000 1930
rect 8000 1890 8010 1930
rect 7950 1880 8010 1890
rect 8030 1930 8090 1940
rect 8030 1890 8040 1930
rect 8040 1890 8080 1930
rect 8080 1890 8090 1930
rect 8030 1880 8090 1890
rect 8110 1930 8170 1940
rect 8110 1890 8120 1930
rect 8120 1890 8160 1930
rect 8160 1890 8170 1930
rect 8110 1880 8170 1890
rect 8190 1930 8250 1940
rect 8190 1890 8200 1930
rect 8200 1890 8240 1930
rect 8240 1890 8250 1930
rect 8190 1880 8250 1890
rect 7450 1800 7510 1810
rect 7450 1760 7460 1800
rect 7460 1760 7500 1800
rect 7500 1760 7510 1800
rect 7450 1750 7510 1760
rect 9000 1750 9060 1810
rect 7600 1630 7660 1640
rect 7600 1590 7610 1630
rect 7610 1590 7650 1630
rect 7650 1590 7660 1630
rect 7600 1580 7660 1590
rect 30 90 90 100
rect 30 50 40 90
rect 40 50 80 90
rect 80 50 90 90
rect 30 40 90 50
rect 130 90 190 100
rect 130 50 140 90
rect 140 50 180 90
rect 180 50 190 90
rect 130 40 190 50
rect 230 90 290 100
rect 230 50 240 90
rect 240 50 280 90
rect 280 50 290 90
rect 230 40 290 50
rect 320 90 380 100
rect 320 50 330 90
rect 330 50 370 90
rect 370 50 380 90
rect 320 40 380 50
rect 400 90 460 100
rect 400 50 410 90
rect 410 50 450 90
rect 450 50 460 90
rect 400 40 460 50
rect 490 90 550 100
rect 490 50 500 90
rect 500 50 540 90
rect 540 50 550 90
rect 490 40 550 50
rect 580 90 640 100
rect 580 50 590 90
rect 590 50 630 90
rect 630 50 640 90
rect 580 40 640 50
rect 670 90 730 100
rect 670 50 680 90
rect 680 50 720 90
rect 720 50 730 90
rect 670 40 730 50
rect 760 90 820 100
rect 760 50 770 90
rect 770 50 810 90
rect 810 50 820 90
rect 760 40 820 50
rect 850 90 910 100
rect 850 50 860 90
rect 860 50 900 90
rect 900 50 910 90
rect 850 40 910 50
rect 940 90 1000 100
rect 940 50 950 90
rect 950 50 990 90
rect 990 50 1000 90
rect 940 40 1000 50
rect 1030 90 1090 100
rect 1030 50 1040 90
rect 1040 50 1080 90
rect 1080 50 1090 90
rect 1030 40 1090 50
rect 1120 90 1180 100
rect 1120 50 1130 90
rect 1130 50 1170 90
rect 1170 50 1180 90
rect 1120 40 1180 50
rect 1220 90 1280 100
rect 1220 50 1230 90
rect 1230 50 1270 90
rect 1270 50 1280 90
rect 1220 40 1280 50
rect 1310 90 1370 100
rect 1310 50 1320 90
rect 1320 50 1360 90
rect 1360 50 1370 90
rect 1310 40 1370 50
rect 1410 90 1470 100
rect 1410 50 1420 90
rect 1420 50 1460 90
rect 1460 50 1470 90
rect 1410 40 1470 50
rect 1490 90 1550 100
rect 1490 50 1500 90
rect 1500 50 1540 90
rect 1540 50 1550 90
rect 1490 40 1550 50
rect 1580 90 1640 100
rect 1580 50 1590 90
rect 1590 50 1630 90
rect 1630 50 1640 90
rect 1580 40 1640 50
rect 1670 90 1730 100
rect 1670 50 1680 90
rect 1680 50 1720 90
rect 1720 50 1730 90
rect 1670 40 1730 50
rect 1760 90 1820 100
rect 1760 50 1770 90
rect 1770 50 1810 90
rect 1810 50 1820 90
rect 1760 40 1820 50
rect 1850 90 1910 100
rect 1850 50 1860 90
rect 1860 50 1900 90
rect 1900 50 1910 90
rect 1850 40 1910 50
rect 1940 90 2000 100
rect 1940 50 1950 90
rect 1950 50 1990 90
rect 1990 50 2000 90
rect 1940 40 2000 50
rect 2030 90 2090 100
rect 2030 50 2040 90
rect 2040 50 2080 90
rect 2080 50 2090 90
rect 2030 40 2090 50
rect 2120 90 2180 100
rect 2120 50 2130 90
rect 2130 50 2170 90
rect 2170 50 2180 90
rect 2120 40 2180 50
rect 2210 90 2270 100
rect 2210 50 2220 90
rect 2220 50 2260 90
rect 2260 50 2270 90
rect 2210 40 2270 50
rect 2300 90 2360 100
rect 2300 50 2310 90
rect 2310 50 2350 90
rect 2350 50 2360 90
rect 2300 40 2360 50
rect 2390 90 2450 100
rect 2390 50 2400 90
rect 2400 50 2440 90
rect 2440 50 2450 90
rect 2390 40 2450 50
rect 2480 90 2540 100
rect 2480 50 2490 90
rect 2490 50 2530 90
rect 2530 50 2540 90
rect 2480 40 2540 50
rect 2580 90 2640 100
rect 2580 50 2590 90
rect 2590 50 2630 90
rect 2630 50 2640 90
rect 2580 40 2640 50
rect 2670 90 2730 100
rect 2670 50 2680 90
rect 2680 50 2720 90
rect 2720 50 2730 90
rect 2670 40 2730 50
rect 2760 90 2820 100
rect 2760 50 2770 90
rect 2770 50 2810 90
rect 2810 50 2820 90
rect 2760 40 2820 50
rect 2850 90 2910 100
rect 2850 50 2860 90
rect 2860 50 2900 90
rect 2900 50 2910 90
rect 2850 40 2910 50
rect 2940 90 3000 100
rect 2940 50 2950 90
rect 2950 50 2990 90
rect 2990 50 3000 90
rect 2940 40 3000 50
rect 3030 90 3090 100
rect 3030 50 3040 90
rect 3040 50 3080 90
rect 3080 50 3090 90
rect 3030 40 3090 50
rect 3120 90 3180 100
rect 3120 50 3130 90
rect 3130 50 3170 90
rect 3170 50 3180 90
rect 3120 40 3180 50
rect 3210 90 3270 100
rect 3210 50 3220 90
rect 3220 50 3260 90
rect 3260 50 3270 90
rect 3210 40 3270 50
rect 3300 90 3360 100
rect 3300 50 3310 90
rect 3310 50 3350 90
rect 3350 50 3360 90
rect 3300 40 3360 50
rect 3390 90 3450 100
rect 3390 50 3400 90
rect 3400 50 3440 90
rect 3440 50 3450 90
rect 3390 40 3450 50
rect 3480 90 3540 100
rect 3480 50 3490 90
rect 3490 50 3530 90
rect 3530 50 3540 90
rect 3480 40 3540 50
rect 3570 90 3630 100
rect 3570 50 3580 90
rect 3580 50 3620 90
rect 3620 50 3630 90
rect 3570 40 3630 50
rect 3660 90 3720 100
rect 3660 50 3670 90
rect 3670 50 3710 90
rect 3710 50 3720 90
rect 3660 40 3720 50
rect 3750 90 3810 100
rect 3750 50 3760 90
rect 3760 50 3800 90
rect 3800 50 3810 90
rect 3750 40 3810 50
rect 3840 90 3900 100
rect 3840 50 3850 90
rect 3850 50 3890 90
rect 3890 50 3900 90
rect 3840 40 3900 50
rect 3940 90 4000 100
rect 3940 50 3950 90
rect 3950 50 3990 90
rect 3990 50 4000 90
rect 3940 40 4000 50
rect 4030 90 4090 100
rect 4030 50 4040 90
rect 4040 50 4080 90
rect 4080 50 4090 90
rect 4030 40 4090 50
rect 4120 90 4180 100
rect 4120 50 4130 90
rect 4130 50 4170 90
rect 4170 50 4180 90
rect 4120 40 4180 50
rect 4210 90 4270 100
rect 4210 50 4220 90
rect 4220 50 4260 90
rect 4260 50 4270 90
rect 4210 40 4270 50
rect 4300 90 4360 100
rect 4300 50 4310 90
rect 4310 50 4350 90
rect 4350 50 4360 90
rect 4300 40 4360 50
rect 4390 90 4450 100
rect 4390 50 4400 90
rect 4400 50 4440 90
rect 4440 50 4450 90
rect 4390 40 4450 50
rect 4480 90 4540 100
rect 4480 50 4490 90
rect 4490 50 4530 90
rect 4530 50 4540 90
rect 4480 40 4540 50
rect 4570 90 4630 100
rect 4570 50 4580 90
rect 4580 50 4620 90
rect 4620 50 4630 90
rect 4570 40 4630 50
rect 4660 90 4720 100
rect 4660 50 4670 90
rect 4670 50 4710 90
rect 4710 50 4720 90
rect 4660 40 4720 50
rect 4750 90 4810 100
rect 4750 50 4760 90
rect 4760 50 4800 90
rect 4800 50 4810 90
rect 4750 40 4810 50
rect 4840 90 4900 100
rect 4840 50 4850 90
rect 4850 50 4890 90
rect 4890 50 4900 90
rect 4840 40 4900 50
rect 4930 90 4990 100
rect 4930 50 4940 90
rect 4940 50 4980 90
rect 4980 50 4990 90
rect 4930 40 4990 50
rect 5020 90 5080 100
rect 5020 50 5030 90
rect 5030 50 5070 90
rect 5070 50 5080 90
rect 5020 40 5080 50
rect 5110 90 5170 100
rect 5110 50 5120 90
rect 5120 50 5160 90
rect 5160 50 5170 90
rect 5110 40 5170 50
rect 5200 90 5260 100
rect 5200 50 5210 90
rect 5210 50 5250 90
rect 5250 50 5260 90
rect 5200 40 5260 50
rect 5300 90 5360 100
rect 5300 50 5310 90
rect 5310 50 5350 90
rect 5350 50 5360 90
rect 5300 40 5360 50
rect 5390 90 5450 100
rect 5390 50 5400 90
rect 5400 50 5440 90
rect 5440 50 5450 90
rect 5390 40 5450 50
rect 5480 90 5540 100
rect 5480 50 5490 90
rect 5490 50 5530 90
rect 5530 50 5540 90
rect 5480 40 5540 50
rect 5570 90 5630 100
rect 5570 50 5580 90
rect 5580 50 5620 90
rect 5620 50 5630 90
rect 5570 40 5630 50
rect 5660 90 5720 100
rect 5660 50 5670 90
rect 5670 50 5710 90
rect 5710 50 5720 90
rect 5660 40 5720 50
rect 5750 90 5810 100
rect 5750 50 5760 90
rect 5760 50 5800 90
rect 5800 50 5810 90
rect 5750 40 5810 50
rect 5840 90 5900 100
rect 5840 50 5850 90
rect 5850 50 5890 90
rect 5890 50 5900 90
rect 5840 40 5900 50
rect 5930 90 5990 100
rect 5930 50 5940 90
rect 5940 50 5980 90
rect 5980 50 5990 90
rect 5930 40 5990 50
rect 6020 90 6080 100
rect 6020 50 6030 90
rect 6030 50 6070 90
rect 6070 50 6080 90
rect 6020 40 6080 50
rect 6110 90 6170 100
rect 6110 50 6120 90
rect 6120 50 6160 90
rect 6160 50 6170 90
rect 6110 40 6170 50
rect 6200 90 6260 100
rect 6200 50 6210 90
rect 6210 50 6250 90
rect 6250 50 6260 90
rect 6200 40 6260 50
rect 6290 90 6350 100
rect 6290 50 6300 90
rect 6300 50 6340 90
rect 6340 50 6350 90
rect 6290 40 6350 50
rect 6380 90 6440 100
rect 6380 50 6390 90
rect 6390 50 6430 90
rect 6430 50 6440 90
rect 6380 40 6440 50
rect 6470 90 6530 100
rect 6470 50 6480 90
rect 6480 50 6520 90
rect 6520 50 6530 90
rect 6470 40 6530 50
rect 6560 90 6620 100
rect 6560 50 6570 90
rect 6570 50 6610 90
rect 6610 50 6620 90
rect 6560 40 6620 50
rect 6650 90 6710 100
rect 6650 50 6660 90
rect 6660 50 6700 90
rect 6700 50 6710 90
rect 6650 40 6710 50
rect 6750 90 6810 100
rect 6750 50 6760 90
rect 6760 50 6800 90
rect 6800 50 6810 90
rect 6750 40 6810 50
rect 6840 90 6900 100
rect 6840 50 6850 90
rect 6850 50 6890 90
rect 6890 50 6900 90
rect 6840 40 6900 50
rect 6930 90 6990 100
rect 6930 50 6940 90
rect 6940 50 6980 90
rect 6980 50 6990 90
rect 6930 40 6990 50
rect 7020 90 7080 100
rect 7020 50 7030 90
rect 7030 50 7070 90
rect 7070 50 7080 90
rect 7020 40 7080 50
rect 7110 90 7170 100
rect 7110 50 7120 90
rect 7120 50 7160 90
rect 7160 50 7170 90
rect 7110 40 7170 50
rect 7200 90 7260 100
rect 7200 50 7210 90
rect 7210 50 7250 90
rect 7250 50 7260 90
rect 7200 40 7260 50
rect 7290 90 7350 100
rect 7290 50 7300 90
rect 7300 50 7340 90
rect 7340 50 7350 90
rect 7290 40 7350 50
rect 7380 90 7440 100
rect 7380 50 7390 90
rect 7390 50 7430 90
rect 7430 50 7440 90
rect 7380 40 7440 50
rect 7470 90 7530 100
rect 7470 50 7480 90
rect 7480 50 7520 90
rect 7520 50 7530 90
rect 7470 40 7530 50
rect 7560 90 7620 100
rect 7560 50 7570 90
rect 7570 50 7610 90
rect 7610 50 7620 90
rect 7560 40 7620 50
rect 7650 90 7710 100
rect 7650 50 7660 90
rect 7660 50 7700 90
rect 7700 50 7710 90
rect 7650 40 7710 50
rect 7740 90 7800 100
rect 7740 50 7750 90
rect 7750 50 7790 90
rect 7790 50 7800 90
rect 7740 40 7800 50
rect 7830 90 7890 100
rect 7830 50 7840 90
rect 7840 50 7880 90
rect 7880 50 7890 90
rect 7830 40 7890 50
rect 7920 90 7980 100
rect 7920 50 7930 90
rect 7930 50 7970 90
rect 7970 50 7980 90
rect 7920 40 7980 50
rect 8010 90 8070 100
rect 8010 50 8020 90
rect 8020 50 8060 90
rect 8060 50 8070 90
rect 8010 40 8070 50
rect 8110 90 8170 100
rect 8110 50 8120 90
rect 8120 50 8160 90
rect 8160 50 8170 90
rect 8110 40 8170 50
rect 8200 90 8260 100
rect 8200 50 8210 90
rect 8210 50 8250 90
rect 8250 50 8260 90
rect 8200 40 8260 50
rect 8290 90 8350 100
rect 8290 50 8300 90
rect 8300 50 8340 90
rect 8340 50 8350 90
rect 8290 40 8350 50
rect 8380 90 8440 100
rect 8380 50 8390 90
rect 8390 50 8430 90
rect 8430 50 8440 90
rect 8380 40 8440 50
rect 8470 90 8530 100
rect 8470 50 8480 90
rect 8480 50 8520 90
rect 8520 50 8530 90
rect 8470 40 8530 50
rect 8560 90 8620 100
rect 8560 50 8570 90
rect 8570 50 8610 90
rect 8610 50 8620 90
rect 8560 40 8620 50
rect 8650 90 8710 100
rect 8650 50 8660 90
rect 8660 50 8700 90
rect 8700 50 8710 90
rect 8650 40 8710 50
rect 8740 90 8800 100
rect 8740 50 8750 90
rect 8750 50 8790 90
rect 8790 50 8800 90
rect 8740 40 8800 50
rect 8830 90 8890 100
rect 8830 50 8840 90
rect 8840 50 8880 90
rect 8880 50 8890 90
rect 8830 40 8890 50
rect 8920 90 8980 100
rect 8920 50 8930 90
rect 8930 50 8970 90
rect 8970 50 8980 90
rect 8920 40 8980 50
rect 9010 90 9070 100
rect 9010 50 9020 90
rect 9020 50 9060 90
rect 9060 50 9070 90
rect 9010 40 9070 50
rect 9100 90 9160 100
rect 9100 50 9110 90
rect 9110 50 9150 90
rect 9150 50 9160 90
rect 9100 40 9160 50
rect 9190 90 9250 100
rect 9190 50 9200 90
rect 9200 50 9240 90
rect 9240 50 9250 90
rect 9190 40 9250 50
rect 9280 90 9340 100
rect 9280 50 9290 90
rect 9290 50 9330 90
rect 9330 50 9340 90
rect 9280 40 9340 50
rect 9380 90 9440 100
rect 9380 50 9390 90
rect 9390 50 9430 90
rect 9430 50 9440 90
rect 9380 40 9440 50
<< metal2 >>
rect -260 5800 -180 5810
rect -260 5740 -250 5800
rect -190 5740 -180 5800
rect -260 5730 -180 5740
rect 9660 5800 9740 5810
rect 9660 5740 9670 5800
rect 9730 5740 9740 5800
rect 9660 5730 9740 5740
rect -260 5550 -180 5560
rect -260 5490 -250 5550
rect -190 5540 -180 5550
rect 4620 5550 4700 5560
rect 4620 5540 4630 5550
rect -190 5500 4630 5540
rect -190 5490 -180 5500
rect -260 5480 -180 5490
rect 4620 5490 4630 5500
rect 4690 5540 4700 5550
rect 5020 5550 5100 5560
rect 5020 5540 5030 5550
rect 4690 5500 5030 5540
rect 4690 5490 4700 5500
rect 4620 5480 4700 5490
rect 5020 5490 5030 5500
rect 5090 5540 5100 5550
rect 5420 5550 5500 5560
rect 5420 5540 5430 5550
rect 5090 5500 5430 5540
rect 5090 5490 5100 5500
rect 5020 5480 5100 5490
rect 5420 5490 5430 5500
rect 5490 5540 5500 5550
rect 5820 5550 5900 5560
rect 5820 5540 5830 5550
rect 5490 5500 5830 5540
rect 5490 5490 5500 5500
rect 5420 5480 5500 5490
rect 5820 5490 5830 5500
rect 5890 5540 5900 5550
rect 6220 5550 6300 5560
rect 6220 5540 6230 5550
rect 5890 5500 6230 5540
rect 5890 5490 5900 5500
rect 5820 5480 5900 5490
rect 6220 5490 6230 5500
rect 6290 5540 6300 5550
rect 6620 5550 6700 5560
rect 6620 5540 6630 5550
rect 6290 5500 6630 5540
rect 6290 5490 6300 5500
rect 6220 5480 6300 5490
rect 6620 5490 6630 5500
rect 6690 5540 6700 5550
rect 7020 5550 7100 5560
rect 7020 5540 7030 5550
rect 6690 5500 7030 5540
rect 6690 5490 6700 5500
rect 6620 5480 6700 5490
rect 7020 5490 7030 5500
rect 7090 5540 7100 5550
rect 7420 5550 7500 5560
rect 7420 5540 7430 5550
rect 7090 5500 7430 5540
rect 7090 5490 7100 5500
rect 7020 5480 7100 5490
rect 7420 5490 7430 5500
rect 7490 5540 7500 5550
rect 7820 5550 7900 5560
rect 7820 5540 7830 5550
rect 7490 5500 7830 5540
rect 7490 5490 7500 5500
rect 7420 5480 7500 5490
rect 7820 5490 7830 5500
rect 7890 5540 7900 5550
rect 8220 5550 8300 5560
rect 8220 5540 8230 5550
rect 7890 5500 8230 5540
rect 7890 5490 7900 5500
rect 7820 5480 7900 5490
rect 8220 5490 8230 5500
rect 8290 5540 8300 5550
rect 9660 5550 9740 5560
rect 9660 5540 9670 5550
rect 8290 5500 9670 5540
rect 8290 5490 8300 5500
rect 8220 5480 8300 5490
rect 9660 5490 9670 5500
rect 9730 5490 9740 5550
rect 9660 5480 9740 5490
rect -110 5030 1970 5040
rect -110 4970 -100 5030
rect -40 4970 1900 5030
rect 1960 4970 1970 5030
rect -110 4960 1970 4970
rect 4300 4610 4380 4620
rect 4300 4550 4310 4610
rect 4370 4600 4380 4610
rect 4820 4610 4900 4620
rect 4820 4600 4830 4610
rect 4370 4560 4830 4600
rect 4370 4550 4380 4560
rect 4300 4540 4380 4550
rect 4820 4550 4830 4560
rect 4890 4600 4900 4610
rect 6820 4610 6900 4620
rect 6820 4600 6830 4610
rect 4890 4560 6830 4600
rect 4890 4550 4900 4560
rect 4820 4540 4900 4550
rect 6820 4550 6830 4560
rect 6890 4600 6900 4610
rect 7620 4610 7700 4620
rect 7620 4600 7630 4610
rect 6890 4560 7630 4600
rect 6890 4550 6900 4560
rect 6820 4540 6900 4550
rect 7620 4550 7630 4560
rect 7690 4550 7700 4610
rect 7620 4540 7700 4550
rect 8140 4610 8220 4620
rect 8140 4550 8150 4610
rect 8210 4600 8220 4610
rect 8750 4610 8830 4620
rect 8750 4600 8760 4610
rect 8210 4560 8760 4600
rect 8210 4550 8220 4560
rect 8140 4540 8220 4550
rect 8750 4550 8760 4560
rect 8820 4550 8830 4610
rect 8750 4540 8830 4550
rect 5220 4520 5300 4530
rect 5220 4460 5230 4520
rect 5290 4510 5300 4520
rect 6020 4520 6100 4530
rect 6020 4510 6030 4520
rect 5290 4470 6030 4510
rect 5290 4460 5300 4470
rect 5220 4450 5300 4460
rect 6020 4460 6030 4470
rect 6090 4510 6100 4520
rect 8020 4520 8100 4530
rect 8020 4510 8030 4520
rect 6090 4470 8030 4510
rect 6090 4460 6100 4470
rect 6020 4450 6100 4460
rect 8020 4460 8030 4470
rect 8090 4510 8100 4520
rect 8630 4520 8710 4530
rect 8630 4510 8640 4520
rect 8090 4470 8640 4510
rect 8090 4460 8100 4470
rect 8020 4450 8100 4460
rect 8630 4460 8640 4470
rect 8700 4460 8710 4520
rect 8630 4450 8710 4460
rect 3790 4440 4230 4450
rect 3790 4380 3800 4440
rect 4220 4420 4230 4440
rect 5620 4430 5700 4440
rect 5620 4420 5630 4430
rect 4220 4380 5630 4420
rect 3790 4370 4230 4380
rect 5620 4370 5630 4380
rect 5690 4420 5700 4430
rect 6420 4430 6500 4440
rect 6420 4420 6430 4430
rect 5690 4380 6430 4420
rect 5690 4370 5700 4380
rect 5620 4360 5700 4370
rect 6420 4370 6430 4380
rect 6490 4420 6500 4430
rect 7220 4430 7300 4440
rect 7220 4420 7230 4430
rect 6490 4380 7230 4420
rect 6490 4370 6500 4380
rect 6420 4360 6500 4370
rect 7220 4370 7230 4380
rect 7290 4370 7300 4430
rect 7220 4360 7300 4370
rect -260 4240 -180 4250
rect -260 4180 -250 4240
rect -190 4230 -180 4240
rect 4460 4240 4540 4250
rect 4460 4230 4470 4240
rect -190 4190 4470 4230
rect -190 4180 -180 4190
rect -260 4170 -180 4180
rect 4460 4180 4470 4190
rect 4530 4230 4540 4240
rect 4660 4240 4740 4250
rect 4660 4230 4670 4240
rect 4530 4190 4670 4230
rect 4530 4180 4540 4190
rect 4460 4170 4540 4180
rect 4660 4180 4670 4190
rect 4730 4230 4740 4240
rect 5060 4240 5140 4250
rect 5060 4230 5070 4240
rect 4730 4190 5070 4230
rect 4730 4180 4740 4190
rect 4660 4170 4740 4180
rect 5060 4180 5070 4190
rect 5130 4230 5140 4240
rect 5460 4240 5540 4250
rect 5460 4230 5470 4240
rect 5130 4190 5470 4230
rect 5130 4180 5140 4190
rect 5060 4170 5140 4180
rect 5460 4180 5470 4190
rect 5530 4230 5540 4240
rect 5660 4240 5740 4250
rect 5660 4230 5670 4240
rect 5530 4190 5670 4230
rect 5530 4180 5540 4190
rect 5460 4170 5540 4180
rect 5660 4180 5670 4190
rect 5730 4230 5740 4240
rect 5820 4240 5900 4250
rect 5820 4230 5830 4240
rect 5730 4190 5830 4230
rect 5730 4180 5740 4190
rect 5660 4170 5740 4180
rect 5820 4180 5830 4190
rect 5890 4230 5900 4240
rect 6020 4240 6100 4250
rect 6020 4230 6030 4240
rect 5890 4190 6030 4230
rect 5890 4180 5900 4190
rect 5820 4170 5900 4180
rect 6020 4180 6030 4190
rect 6090 4230 6100 4240
rect 6420 4240 6500 4250
rect 6420 4230 6430 4240
rect 6090 4190 6430 4230
rect 6090 4180 6100 4190
rect 6020 4170 6100 4180
rect 6420 4180 6430 4190
rect 6490 4230 6500 4240
rect 6820 4240 6900 4250
rect 6820 4230 6830 4240
rect 6490 4190 6830 4230
rect 6490 4180 6500 4190
rect 6420 4170 6500 4180
rect 6820 4180 6830 4190
rect 6890 4230 6900 4240
rect 7020 4240 7100 4250
rect 7020 4230 7030 4240
rect 6890 4190 7030 4230
rect 6890 4180 6900 4190
rect 6820 4170 6900 4180
rect 7020 4180 7030 4190
rect 7090 4230 7100 4240
rect 7180 4240 7260 4250
rect 7180 4230 7190 4240
rect 7090 4190 7190 4230
rect 7090 4180 7100 4190
rect 7020 4170 7100 4180
rect 7180 4180 7190 4190
rect 7250 4230 7260 4240
rect 7380 4240 7460 4250
rect 7380 4230 7390 4240
rect 7250 4190 7390 4230
rect 7250 4180 7260 4190
rect 7180 4170 7260 4180
rect 7380 4180 7390 4190
rect 7450 4230 7460 4240
rect 7780 4240 7860 4250
rect 7780 4230 7790 4240
rect 7450 4190 7790 4230
rect 7450 4180 7460 4190
rect 7380 4170 7460 4180
rect 7780 4180 7790 4190
rect 7850 4230 7860 4240
rect 8180 4240 8260 4250
rect 8180 4230 8190 4240
rect 7850 4190 8190 4230
rect 7850 4180 7860 4190
rect 7780 4170 7860 4180
rect 8180 4180 8190 4190
rect 8250 4230 8260 4240
rect 8380 4240 8460 4250
rect 8380 4230 8390 4240
rect 8250 4190 8390 4230
rect 8250 4180 8260 4190
rect 8180 4170 8260 4180
rect 8380 4180 8390 4190
rect 8450 4230 8460 4240
rect 9150 4240 9230 4250
rect 9150 4230 9160 4240
rect 8450 4190 9160 4230
rect 8450 4180 8460 4190
rect 8380 4170 8460 4180
rect 9150 4180 9160 4190
rect 9220 4230 9230 4240
rect 9660 4240 9740 4250
rect 9660 4230 9670 4240
rect 9220 4190 9670 4230
rect 9220 4180 9230 4190
rect 9150 4170 9230 4180
rect 9660 4180 9670 4190
rect 9730 4180 9740 4240
rect 9660 4170 9740 4180
rect -110 4030 1970 4040
rect -110 3970 -100 4030
rect -40 3970 1900 4030
rect 1960 3970 1970 4030
rect -110 3960 1970 3970
rect 5260 3700 5340 3710
rect 5260 3640 5270 3700
rect 5330 3690 5340 3700
rect 5940 3700 6020 3710
rect 5940 3690 5950 3700
rect 5330 3650 5950 3690
rect 5330 3640 5340 3650
rect 5260 3630 5340 3640
rect 5940 3640 5950 3650
rect 6010 3690 6020 3700
rect 6900 3700 6980 3710
rect 6900 3690 6910 3700
rect 6010 3650 6910 3690
rect 6010 3640 6020 3650
rect 5940 3630 6020 3640
rect 6900 3640 6910 3650
rect 6970 3690 6980 3700
rect 7580 3700 7660 3710
rect 7580 3690 7590 3700
rect 6970 3650 7590 3690
rect 6970 3640 6980 3650
rect 6900 3630 6980 3640
rect 7580 3640 7590 3650
rect 7650 3640 7660 3700
rect 7580 3630 7660 3640
rect 4860 3610 4940 3620
rect 4860 3550 4870 3610
rect 4930 3600 4940 3610
rect 5540 3610 5620 3620
rect 5540 3600 5550 3610
rect 4930 3560 5550 3600
rect 4930 3550 4940 3560
rect 4860 3540 4940 3550
rect 5540 3550 5550 3560
rect 5610 3600 5620 3610
rect 6120 3610 6200 3620
rect 6120 3600 6130 3610
rect 5610 3560 6130 3600
rect 5610 3550 5620 3560
rect 5540 3540 5620 3550
rect 6120 3550 6130 3560
rect 6190 3600 6200 3610
rect 6720 3610 6800 3620
rect 6720 3600 6730 3610
rect 6190 3560 6730 3600
rect 6190 3550 6200 3560
rect 6120 3540 6200 3550
rect 6720 3550 6730 3560
rect 6790 3600 6800 3610
rect 7300 3610 7380 3620
rect 7300 3600 7310 3610
rect 6790 3560 7310 3600
rect 6790 3550 6800 3560
rect 6720 3540 6800 3550
rect 7300 3550 7310 3560
rect 7370 3600 7380 3610
rect 7980 3610 8060 3620
rect 7980 3600 7990 3610
rect 7370 3560 7990 3600
rect 7370 3550 7380 3560
rect 7300 3540 7380 3550
rect 7980 3550 7990 3560
rect 8050 3550 8060 3610
rect 7980 3540 8060 3550
rect 6420 3520 6500 3530
rect 6420 3460 6430 3520
rect 6490 3510 6500 3520
rect 8440 3520 8520 3530
rect 8440 3510 8450 3520
rect 6490 3470 8450 3510
rect 6490 3460 6500 3470
rect 6420 3450 6500 3460
rect 8440 3460 8450 3470
rect 8510 3460 8520 3520
rect 8440 3450 8520 3460
rect 880 3440 4230 3450
rect 880 3380 890 3440
rect 950 3380 3800 3440
rect 4220 3420 4230 3440
rect 4300 3430 4380 3440
rect 4300 3420 4310 3430
rect 4220 3380 4310 3420
rect 880 3370 4230 3380
rect 4300 3370 4310 3380
rect 4370 3420 4380 3430
rect 6060 3430 6140 3440
rect 6060 3420 6070 3430
rect 4370 3380 6070 3420
rect 4370 3370 4380 3380
rect 4300 3360 4380 3370
rect 6060 3370 6070 3380
rect 6130 3420 6140 3430
rect 6780 3430 6860 3440
rect 6780 3420 6790 3430
rect 6130 3380 6790 3420
rect 6130 3370 6140 3380
rect 6060 3360 6140 3370
rect 6780 3370 6790 3380
rect 6850 3420 6860 3430
rect 8860 3430 8940 3440
rect 8860 3420 8870 3430
rect 6850 3380 8870 3420
rect 6850 3370 6860 3380
rect 6780 3360 6860 3370
rect 8860 3370 8870 3380
rect 8930 3370 8940 3430
rect 8860 3360 8940 3370
rect 5540 3090 5620 3100
rect 1720 3080 1970 3090
rect 1720 3020 1730 3080
rect 1790 3020 1900 3080
rect 1960 3020 1970 3080
rect 1720 3010 1970 3020
rect 3790 3080 4230 3090
rect 5540 3080 5550 3090
rect 3790 3020 3800 3080
rect 4220 3040 5550 3080
rect 4220 3020 4230 3040
rect 5540 3030 5550 3040
rect 5610 3080 5620 3090
rect 7300 3090 7380 3100
rect 7300 3080 7310 3090
rect 5610 3040 7310 3080
rect 5610 3030 5620 3040
rect 5540 3020 5620 3030
rect 7300 3030 7310 3040
rect 7370 3080 7380 3090
rect 8630 3090 8710 3100
rect 8630 3080 8640 3090
rect 7370 3040 8640 3080
rect 7370 3030 7380 3040
rect 7300 3020 7380 3030
rect 8630 3030 8640 3040
rect 8700 3030 8710 3090
rect 8630 3020 8710 3030
rect 3790 3010 4230 3020
rect 5140 3000 5220 3010
rect 5140 2940 5150 3000
rect 5210 2990 5220 3000
rect 5340 3000 5420 3010
rect 5340 2990 5350 3000
rect 5210 2950 5350 2990
rect 5210 2940 5220 2950
rect 5140 2930 5220 2940
rect 5340 2940 5350 2950
rect 5410 2990 5420 3000
rect 5740 3000 5820 3010
rect 5740 2990 5750 3000
rect 5410 2950 5750 2990
rect 5410 2940 5420 2950
rect 5340 2930 5420 2940
rect 5740 2940 5750 2950
rect 5810 2990 5820 3000
rect 6140 3000 6220 3010
rect 6140 2990 6150 3000
rect 5810 2950 6150 2990
rect 5810 2940 5820 2950
rect 5740 2930 5820 2940
rect 6140 2940 6150 2950
rect 6210 2990 6220 3000
rect 6340 3000 6420 3010
rect 6340 2990 6350 3000
rect 6210 2950 6350 2990
rect 6210 2940 6220 2950
rect 6140 2930 6220 2940
rect 6340 2940 6350 2950
rect 6410 2990 6420 3000
rect 6500 3000 6580 3010
rect 6500 2990 6510 3000
rect 6410 2950 6510 2990
rect 6410 2940 6420 2950
rect 6340 2930 6420 2940
rect 6500 2940 6510 2950
rect 6570 2990 6580 3000
rect 6700 3000 6780 3010
rect 6700 2990 6710 3000
rect 6570 2950 6710 2990
rect 6570 2940 6580 2950
rect 6500 2930 6580 2940
rect 6700 2940 6710 2950
rect 6770 2990 6780 3000
rect 7100 3000 7180 3010
rect 7100 2990 7110 3000
rect 6770 2950 7110 2990
rect 6770 2940 6780 2950
rect 6700 2930 6780 2940
rect 7100 2940 7110 2950
rect 7170 2990 7180 3000
rect 7500 3000 7580 3010
rect 7500 2990 7510 3000
rect 7170 2950 7510 2990
rect 7170 2940 7180 2950
rect 7100 2930 7180 2940
rect 7500 2940 7510 2950
rect 7570 2990 7580 3000
rect 7700 3000 7780 3010
rect 7700 2990 7710 3000
rect 7570 2950 7710 2990
rect 7570 2940 7580 2950
rect 7500 2930 7580 2940
rect 7700 2940 7710 2950
rect 7770 2940 7780 3000
rect 7700 2930 7780 2940
rect 7300 2880 7380 2890
rect 7300 2820 7310 2880
rect 7370 2870 7380 2880
rect 8440 2880 8520 2890
rect 8440 2870 8450 2880
rect 7370 2830 8450 2870
rect 7370 2820 7380 2830
rect 7300 2810 7380 2820
rect 8440 2820 8450 2830
rect 8510 2820 8520 2880
rect 8440 2810 8520 2820
rect -110 2490 1970 2500
rect -110 2430 -100 2490
rect -40 2430 1900 2490
rect 1960 2430 1970 2490
rect -110 2420 1970 2430
rect 4660 1940 5620 1950
rect 4660 1880 4670 1940
rect 4730 1880 4750 1940
rect 4810 1880 4830 1940
rect 4890 1880 4910 1940
rect 4970 1880 4990 1940
rect 5050 1880 5070 1940
rect 5130 1880 5150 1940
rect 5210 1880 5230 1940
rect 5290 1880 5310 1940
rect 5370 1880 5390 1940
rect 5450 1880 5470 1940
rect 5530 1880 5550 1940
rect 5610 1930 5620 1940
rect 7300 1940 8260 1950
rect 7300 1930 7310 1940
rect 5610 1890 7310 1930
rect 5610 1880 5620 1890
rect 4660 1870 5620 1880
rect 7300 1880 7310 1890
rect 7370 1880 7390 1940
rect 7450 1880 7470 1940
rect 7530 1880 7550 1940
rect 7610 1880 7630 1940
rect 7690 1880 7710 1940
rect 7770 1880 7790 1940
rect 7850 1880 7870 1940
rect 7930 1880 7950 1940
rect 8010 1880 8030 1940
rect 8090 1880 8110 1940
rect 8170 1880 8190 1940
rect 8250 1930 8260 1940
rect 9510 1940 9590 1950
rect 9510 1930 9520 1940
rect 8250 1890 9520 1930
rect 8250 1880 8260 1890
rect 7300 1870 8260 1880
rect 9510 1880 9520 1890
rect 9580 1880 9590 1940
rect 9510 1870 9590 1880
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1800 7520 1810
rect 8990 1810 9070 1820
rect 8990 1800 9000 1810
rect 7510 1760 9000 1800
rect 7510 1750 7520 1760
rect 7440 1740 7520 1750
rect 8990 1750 9000 1760
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect 7590 1640 7670 1650
rect 7590 1580 7600 1640
rect 7660 1630 7670 1640
rect 9510 1640 9590 1650
rect 9510 1630 9520 1640
rect 7660 1590 9520 1630
rect 7660 1580 7670 1590
rect 7590 1570 7670 1580
rect 9510 1580 9520 1590
rect 9580 1580 9590 1640
rect 9510 1570 9590 1580
rect -110 100 9590 110
rect -110 40 -100 100
rect -40 40 30 100
rect 90 40 130 100
rect 190 40 230 100
rect 290 40 320 100
rect 380 40 400 100
rect 460 40 490 100
rect 550 40 580 100
rect 640 40 670 100
rect 730 40 760 100
rect 820 40 850 100
rect 910 40 940 100
rect 1000 40 1030 100
rect 1090 40 1120 100
rect 1180 40 1220 100
rect 1280 40 1310 100
rect 1370 40 1410 100
rect 1470 40 1490 100
rect 1550 40 1580 100
rect 1640 40 1670 100
rect 1730 40 1760 100
rect 1820 40 1850 100
rect 1910 40 1940 100
rect 2000 40 2030 100
rect 2090 40 2120 100
rect 2180 40 2210 100
rect 2270 40 2300 100
rect 2360 40 2390 100
rect 2450 40 2480 100
rect 2540 40 2580 100
rect 2640 40 2670 100
rect 2730 40 2760 100
rect 2820 40 2850 100
rect 2910 40 2940 100
rect 3000 40 3030 100
rect 3090 40 3120 100
rect 3180 40 3210 100
rect 3270 40 3300 100
rect 3360 40 3390 100
rect 3450 40 3480 100
rect 3540 40 3570 100
rect 3630 40 3660 100
rect 3720 40 3750 100
rect 3810 40 3840 100
rect 3900 40 3940 100
rect 4000 40 4030 100
rect 4090 40 4120 100
rect 4180 40 4210 100
rect 4270 40 4300 100
rect 4360 40 4390 100
rect 4450 40 4480 100
rect 4540 40 4570 100
rect 4630 40 4660 100
rect 4720 40 4750 100
rect 4810 40 4840 100
rect 4900 40 4930 100
rect 4990 40 5020 100
rect 5080 40 5110 100
rect 5170 40 5200 100
rect 5260 40 5300 100
rect 5360 40 5390 100
rect 5450 40 5480 100
rect 5540 40 5570 100
rect 5630 40 5660 100
rect 5720 40 5750 100
rect 5810 40 5840 100
rect 5900 40 5930 100
rect 5990 40 6020 100
rect 6080 40 6110 100
rect 6170 40 6200 100
rect 6260 40 6290 100
rect 6350 40 6380 100
rect 6440 40 6470 100
rect 6530 40 6560 100
rect 6620 40 6650 100
rect 6710 40 6750 100
rect 6810 40 6840 100
rect 6900 40 6930 100
rect 6990 40 7020 100
rect 7080 40 7110 100
rect 7170 40 7200 100
rect 7260 40 7290 100
rect 7350 40 7380 100
rect 7440 40 7470 100
rect 7530 40 7560 100
rect 7620 40 7650 100
rect 7710 40 7740 100
rect 7800 40 7830 100
rect 7890 40 7920 100
rect 7980 40 8010 100
rect 8070 40 8110 100
rect 8170 40 8200 100
rect 8260 40 8290 100
rect 8350 40 8380 100
rect 8440 40 8470 100
rect 8530 40 8560 100
rect 8620 40 8650 100
rect 8710 40 8740 100
rect 8800 40 8830 100
rect 8890 40 8920 100
rect 8980 40 9010 100
rect 9070 40 9100 100
rect 9160 40 9190 100
rect 9250 40 9280 100
rect 9340 40 9380 100
rect 9440 40 9520 100
rect 9580 40 9590 100
rect -110 30 9590 40
rect -260 -180 -180 -170
rect -260 -240 -250 -180
rect -190 -240 -180 -180
rect -260 -250 -180 -240
<< via2 >>
rect -250 5740 -190 5800
rect 9670 5740 9730 5800
rect -250 5490 -190 5550
rect 9670 5490 9730 5550
rect -100 4970 -40 5030
rect -250 4180 -190 4240
rect 9670 4180 9730 4240
rect -100 3970 -40 4030
rect -100 2430 -40 2490
rect 9520 1880 9580 1940
rect 9520 1580 9580 1640
rect -100 40 -40 100
rect 9520 40 9580 100
rect -250 -240 -190 -180
<< metal3 >>
rect -270 5810 -170 5820
rect -270 5730 -260 5810
rect -180 5730 -170 5810
rect -270 5720 -170 5730
rect 9650 5810 9750 5820
rect 9650 5730 9660 5810
rect 9740 5730 9750 5810
rect 9650 5720 9750 5730
rect -260 5550 -180 5720
rect -120 5660 -20 5670
rect -120 5580 -110 5660
rect -30 5580 -20 5660
rect -120 5570 -20 5580
rect 9500 5660 9600 5670
rect 9500 5580 9510 5660
rect 9590 5580 9600 5660
rect 9500 5570 9600 5580
rect -260 5490 -250 5550
rect -190 5490 -180 5550
rect -260 4240 -180 5490
rect -260 4180 -250 4240
rect -190 4180 -180 4240
rect -260 -160 -180 4180
rect -110 5030 -30 5570
rect -110 4970 -100 5030
rect -40 4970 -30 5030
rect -110 4030 -30 4970
rect -110 3970 -100 4030
rect -40 3970 -30 4030
rect -110 2490 -30 3970
rect -110 2430 -100 2490
rect -40 2430 -30 2490
rect -110 100 -30 2430
rect -110 40 -100 100
rect -40 40 -30 100
rect -110 -10 -30 40
rect 9510 1940 9590 5570
rect 9510 1880 9520 1940
rect 9580 1880 9590 1940
rect 9510 1640 9590 1880
rect 9510 1580 9520 1640
rect 9580 1580 9590 1640
rect 9510 100 9590 1580
rect 9510 40 9520 100
rect 9580 40 9590 100
rect 9510 -10 9590 40
rect 9660 5550 9740 5720
rect 9660 5490 9670 5550
rect 9730 5490 9740 5550
rect 9660 4240 9740 5490
rect 9660 4180 9670 4240
rect 9730 4180 9740 4240
rect -120 -20 -20 -10
rect -120 -100 -110 -20
rect -30 -100 -20 -20
rect -120 -110 -20 -100
rect 9500 -20 9600 -10
rect 9500 -100 9510 -20
rect 9590 -100 9600 -20
rect 9500 -110 9600 -100
rect 9660 -160 9740 4180
rect -270 -170 -170 -160
rect -270 -250 -260 -170
rect -180 -250 -170 -170
rect -270 -260 -170 -250
rect 9650 -170 9750 -160
rect 9650 -250 9660 -170
rect 9740 -250 9750 -170
rect 9650 -260 9750 -250
<< via3 >>
rect -260 5800 -180 5810
rect -260 5740 -250 5800
rect -250 5740 -190 5800
rect -190 5740 -180 5800
rect -260 5730 -180 5740
rect 9660 5800 9740 5810
rect 9660 5740 9670 5800
rect 9670 5740 9730 5800
rect 9730 5740 9740 5800
rect 9660 5730 9740 5740
rect -110 5580 -30 5660
rect 9510 5580 9590 5660
rect -110 -100 -30 -20
rect 9510 -100 9590 -20
rect -260 -180 -180 -170
rect -260 -240 -250 -180
rect -250 -240 -190 -180
rect -190 -240 -180 -180
rect -260 -250 -180 -240
rect 9660 -250 9740 -170
<< metal4 >>
rect -270 5810 -170 5820
rect 9650 5810 9750 5820
rect -270 5730 -260 5810
rect -180 5730 9660 5810
rect 9740 5730 9750 5810
rect -270 5720 -170 5730
rect 9650 5720 9750 5730
rect -120 5660 -20 5670
rect 9500 5660 9600 5670
rect -120 5580 -110 5660
rect -30 5580 9510 5660
rect 9590 5580 9600 5660
rect -120 5570 -20 5580
rect 9500 5570 9600 5580
rect -120 -20 -20 -10
rect 9500 -20 9600 -10
rect -120 -100 -110 -20
rect -30 -100 9510 -20
rect 9590 -100 9600 -20
rect -120 -110 -20 -100
rect 9500 -110 9600 -100
rect -270 -170 -170 -160
rect 9650 -170 9750 -160
rect -270 -250 -260 -170
rect -180 -250 9660 -170
rect 9740 -250 9750 -170
rect -270 -260 -170 -250
rect 9650 -260 9750 -250
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 2710 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 -10 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 1350 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 2710 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 4070 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 5430 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 6790 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 4070 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 5430 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1723858470
transform 1 0 6790 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1723858470
transform 1 0 8150 0 1 0
box 0 0 1340 1340
<< labels >>
flabel locali s 8740 1102 8858 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 8763 1252 8864 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 8704 626 8952 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 7380 1102 7498 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 7403 1252 7504 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 7344 626 7592 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 6020 1102 6138 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 6043 1252 6144 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 5984 626 6232 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 4660 1102 4778 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 4683 1252 4784 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 4624 626 4872 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3300 1102 3418 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 3323 1252 3424 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 3264 626 3512 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 1940 1102 2058 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1963 1252 2064 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 1904 626 2152 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel metal3 9740 2800 9740 2800 3 FreeSans 1600 0 160 0 VDDA
port 1 e
flabel metal3 9590 2350 9590 2350 3 FreeSans 1600 0 160 0 GNDA
port 6 e
flabel metal2 4570 3040 4570 3040 5 FreeSans 800 0 0 -160 Vin+
flabel metal2 4570 3380 4570 3380 5 FreeSans 800 0 0 -160 Vin-
flabel metal1 6460 6300 6460 6300 1 FreeSans 1600 0 0 800 V_out
port 5 n
flabel metal1 8830 4580 8830 4580 3 FreeSans 800 0 160 0 V_TOP
flabel metal1 1800 2080 1800 2080 3 FreeSans 800 0 160 0 Vbe2
flabel metal1 9050 3230 9050 3230 3 FreeSans 800 0 160 0 start_up
flabel metal1 5960 3510 5960 3510 7 FreeSans 400 0 -160 0 V_mirror
flabel locali 5760 2910 5760 2910 7 FreeSans 400 0 -160 0 V_p
flabel metal2 8060 3580 8060 3580 3 FreeSans 400 0 160 0 1st_Vout
<< end >>
