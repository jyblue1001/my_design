magic
tech sky130A
timestamp 1752584700
<< nwell >>
rect -30 2305 310 2695
rect 440 2305 780 2525
rect 910 2305 1250 2695
rect 1378 2305 1718 2695
rect -1225 1730 -345 2120
rect -100 1730 780 2120
rect 910 1730 1790 2120
rect 2035 1730 2915 2120
rect -1195 815 -375 1455
rect 395 1215 1295 1505
rect 2065 815 2885 1455
rect -1195 400 -375 640
rect 2065 400 2885 640
<< nmos >>
rect -65 700 -50 850
rect -10 700 5 850
rect 45 700 60 850
rect 100 700 115 850
rect 155 700 170 850
rect 210 700 225 850
rect 265 700 280 850
rect 320 700 335 850
rect 375 700 390 850
rect 430 700 445 850
rect 485 700 500 850
rect 540 700 555 850
rect 755 625 770 875
rect 810 625 825 875
rect 865 625 880 875
rect 920 625 935 875
rect 1135 700 1150 850
rect 1190 700 1205 850
rect 1245 700 1260 850
rect 1300 700 1315 850
rect 1355 700 1370 850
rect 1410 700 1425 850
rect 1465 700 1480 850
rect 1520 700 1535 850
rect 1575 700 1590 850
rect 1630 700 1645 850
rect 1685 700 1700 850
rect 1740 700 1755 850
rect -65 305 -50 455
rect -10 305 5 455
rect 45 305 60 455
rect 100 305 115 455
rect 155 305 170 455
rect 210 305 225 455
rect 265 305 280 455
rect 320 305 335 455
rect 375 305 390 455
rect 430 305 445 455
rect 485 305 500 455
rect 540 305 555 455
rect 755 305 770 455
rect 810 305 825 455
rect 865 305 880 455
rect 920 305 935 455
rect 1135 305 1150 455
rect 1190 305 1205 455
rect 1245 305 1260 455
rect 1300 305 1315 455
rect 1355 305 1370 455
rect 1410 305 1425 455
rect 1465 305 1480 455
rect 1520 305 1535 455
rect 1575 305 1590 455
rect 1630 305 1645 455
rect 1685 305 1700 455
rect 1740 305 1755 455
rect -1095 -70 -1080 230
rect -1040 -70 -1025 230
rect -985 -70 -970 230
rect -930 -70 -915 230
rect -875 -70 -860 230
rect -820 -70 -805 230
rect -765 -70 -750 230
rect -710 -70 -695 230
rect -655 -70 -640 230
rect -600 -70 -585 230
rect -545 -70 -530 230
rect -490 -70 -475 230
rect 755 -290 770 -40
rect 810 -290 825 -40
rect 865 -290 880 -40
rect 920 -290 935 -40
rect 2165 -70 2180 230
rect 2220 -70 2235 230
rect 2275 -70 2290 230
rect 2330 -70 2345 230
rect 2385 -70 2400 230
rect 2440 -70 2455 230
rect 2495 -70 2510 230
rect 2550 -70 2565 230
rect 2605 -70 2620 230
rect 2660 -70 2675 230
rect 2715 -70 2730 230
rect 2770 -70 2785 230
rect -985 -1055 -925 -355
rect -885 -1055 -825 -355
rect -785 -1055 -725 -355
rect -685 -1055 -625 -355
rect -585 -1055 -525 -355
rect -485 -1055 -425 -355
rect 315 -785 330 -535
rect 370 -785 385 -535
rect 425 -785 440 -535
rect 480 -785 495 -535
rect 535 -785 550 -535
rect 590 -785 605 -535
rect 645 -785 660 -535
rect 700 -785 715 -535
rect 755 -785 770 -535
rect 810 -785 825 -535
rect 865 -785 880 -535
rect 920 -785 935 -535
rect 975 -785 990 -535
rect 1030 -785 1045 -535
rect 1085 -785 1100 -535
rect 1140 -785 1155 -535
rect 1195 -785 1210 -535
rect 1250 -785 1265 -535
rect 1305 -785 1320 -535
rect 1360 -785 1375 -535
rect 1415 -785 1430 -535
rect 535 -1100 550 -950
rect 590 -1100 605 -950
rect 645 -1100 660 -950
rect 700 -1100 715 -950
rect 755 -1100 770 -950
rect 810 -1100 825 -950
rect 1000 -1100 1300 -950
rect 2115 -1055 2175 -355
rect 2215 -1055 2275 -355
rect 2315 -1055 2375 -355
rect 2415 -1055 2475 -355
rect 2515 -1055 2575 -355
rect 2615 -1055 2675 -355
<< pmos >>
rect 70 2325 90 2675
rect 130 2325 150 2675
rect 190 2325 210 2675
rect 540 2325 560 2505
rect 600 2325 620 2505
rect 660 2325 680 2505
rect 1010 2325 1030 2675
rect 1070 2325 1090 2675
rect 1130 2325 1150 2675
rect 1478 2325 1498 2675
rect 1538 2325 1558 2675
rect 1598 2325 1618 2675
rect -1125 1750 -1105 2100
rect -1065 1750 -1045 2100
rect -1005 1750 -985 2100
rect -945 1750 -925 2100
rect -885 1750 -865 2100
rect -825 1750 -805 2100
rect -765 1750 -745 2100
rect -705 1750 -685 2100
rect -645 1750 -625 2100
rect -585 1750 -565 2100
rect -525 1750 -505 2100
rect -465 1750 -445 2100
rect 0 1750 20 2100
rect 60 1750 80 2100
rect 120 1750 140 2100
rect 180 1750 200 2100
rect 240 1750 260 2100
rect 300 1750 320 2100
rect 360 1750 380 2100
rect 420 1750 440 2100
rect 480 1750 500 2100
rect 540 1750 560 2100
rect 600 1750 620 2100
rect 660 1750 680 2100
rect 1010 1750 1030 2100
rect 1070 1750 1090 2100
rect 1130 1750 1150 2100
rect 1190 1750 1210 2100
rect 1250 1750 1270 2100
rect 1310 1750 1330 2100
rect 1370 1750 1390 2100
rect 1430 1750 1450 2100
rect 1490 1750 1510 2100
rect 1550 1750 1570 2100
rect 1610 1750 1630 2100
rect 1670 1750 1690 2100
rect 2135 1750 2155 2100
rect 2195 1750 2215 2100
rect 2255 1750 2275 2100
rect 2315 1750 2335 2100
rect 2375 1750 2395 2100
rect 2435 1750 2455 2100
rect 2495 1750 2515 2100
rect 2555 1750 2575 2100
rect 2615 1750 2635 2100
rect 2675 1750 2695 2100
rect 2735 1750 2755 2100
rect 2795 1750 2815 2100
rect -1095 835 -1080 1435
rect -1040 835 -1025 1435
rect -985 835 -970 1435
rect -930 835 -915 1435
rect -875 835 -860 1435
rect -820 835 -805 1435
rect -765 835 -750 1435
rect -710 835 -695 1435
rect -655 835 -640 1435
rect -600 835 -585 1435
rect -545 835 -530 1435
rect -490 835 -475 1435
rect 495 1235 510 1485
rect 550 1235 565 1485
rect 605 1235 620 1485
rect 660 1235 675 1485
rect 715 1235 730 1485
rect 770 1235 785 1485
rect 905 1235 920 1485
rect 960 1235 975 1485
rect 1015 1235 1030 1485
rect 1070 1235 1085 1485
rect 1125 1235 1140 1485
rect 1180 1235 1195 1485
rect 2165 835 2180 1435
rect 2220 835 2235 1435
rect 2275 835 2290 1435
rect 2330 835 2345 1435
rect 2385 835 2400 1435
rect 2440 835 2455 1435
rect 2495 835 2510 1435
rect 2550 835 2565 1435
rect 2605 835 2620 1435
rect 2660 835 2675 1435
rect 2715 835 2730 1435
rect 2770 835 2785 1435
rect -1095 420 -1080 620
rect -1040 420 -1025 620
rect -985 420 -970 620
rect -930 420 -915 620
rect -875 420 -860 620
rect -820 420 -805 620
rect -765 420 -750 620
rect -710 420 -695 620
rect -655 420 -640 620
rect -600 420 -585 620
rect -545 420 -530 620
rect -490 420 -475 620
rect 2165 420 2180 620
rect 2220 420 2235 620
rect 2275 420 2290 620
rect 2330 420 2345 620
rect 2385 420 2400 620
rect 2440 420 2455 620
rect 2495 420 2510 620
rect 2550 420 2565 620
rect 2605 420 2620 620
rect 2660 420 2675 620
rect 2715 420 2730 620
rect 2770 420 2785 620
<< ndiff >>
rect 715 860 755 875
rect -105 835 -65 850
rect -105 815 -95 835
rect -75 815 -65 835
rect -105 785 -65 815
rect -105 765 -95 785
rect -75 765 -65 785
rect -105 735 -65 765
rect -105 715 -95 735
rect -75 715 -65 735
rect -105 700 -65 715
rect -50 835 -10 850
rect -50 815 -40 835
rect -20 815 -10 835
rect -50 785 -10 815
rect -50 765 -40 785
rect -20 765 -10 785
rect -50 735 -10 765
rect -50 715 -40 735
rect -20 715 -10 735
rect -50 700 -10 715
rect 5 835 45 850
rect 5 815 15 835
rect 35 815 45 835
rect 5 785 45 815
rect 5 765 15 785
rect 35 765 45 785
rect 5 735 45 765
rect 5 715 15 735
rect 35 715 45 735
rect 5 700 45 715
rect 60 835 100 850
rect 60 815 70 835
rect 90 815 100 835
rect 60 785 100 815
rect 60 765 70 785
rect 90 765 100 785
rect 60 735 100 765
rect 60 715 70 735
rect 90 715 100 735
rect 60 700 100 715
rect 115 835 155 850
rect 115 815 125 835
rect 145 815 155 835
rect 115 785 155 815
rect 115 765 125 785
rect 145 765 155 785
rect 115 735 155 765
rect 115 715 125 735
rect 145 715 155 735
rect 115 700 155 715
rect 170 835 210 850
rect 170 815 180 835
rect 200 815 210 835
rect 170 785 210 815
rect 170 765 180 785
rect 200 765 210 785
rect 170 735 210 765
rect 170 715 180 735
rect 200 715 210 735
rect 170 700 210 715
rect 225 835 265 850
rect 225 815 235 835
rect 255 815 265 835
rect 225 785 265 815
rect 225 765 235 785
rect 255 765 265 785
rect 225 735 265 765
rect 225 715 235 735
rect 255 715 265 735
rect 225 700 265 715
rect 280 835 320 850
rect 280 815 290 835
rect 310 815 320 835
rect 280 785 320 815
rect 280 765 290 785
rect 310 765 320 785
rect 280 735 320 765
rect 280 715 290 735
rect 310 715 320 735
rect 280 700 320 715
rect 335 835 375 850
rect 335 815 345 835
rect 365 815 375 835
rect 335 785 375 815
rect 335 765 345 785
rect 365 765 375 785
rect 335 735 375 765
rect 335 715 345 735
rect 365 715 375 735
rect 335 700 375 715
rect 390 835 430 850
rect 390 815 400 835
rect 420 815 430 835
rect 390 785 430 815
rect 390 765 400 785
rect 420 765 430 785
rect 390 735 430 765
rect 390 715 400 735
rect 420 715 430 735
rect 390 700 430 715
rect 445 835 485 850
rect 445 815 455 835
rect 475 815 485 835
rect 445 785 485 815
rect 445 765 455 785
rect 475 765 485 785
rect 445 735 485 765
rect 445 715 455 735
rect 475 715 485 735
rect 445 700 485 715
rect 500 835 540 850
rect 500 815 510 835
rect 530 815 540 835
rect 500 785 540 815
rect 500 765 510 785
rect 530 765 540 785
rect 500 735 540 765
rect 500 715 510 735
rect 530 715 540 735
rect 500 700 540 715
rect 555 835 595 850
rect 555 815 565 835
rect 585 815 595 835
rect 555 785 595 815
rect 555 765 565 785
rect 585 765 595 785
rect 555 735 595 765
rect 555 715 565 735
rect 585 715 595 735
rect 555 700 595 715
rect 715 840 725 860
rect 745 840 755 860
rect 715 810 755 840
rect 715 790 725 810
rect 745 790 755 810
rect 715 760 755 790
rect 715 740 725 760
rect 745 740 755 760
rect 715 710 755 740
rect 715 690 725 710
rect 745 690 755 710
rect 715 660 755 690
rect 715 640 725 660
rect 745 640 755 660
rect 715 625 755 640
rect 770 860 810 875
rect 770 840 780 860
rect 800 840 810 860
rect 770 810 810 840
rect 770 790 780 810
rect 800 790 810 810
rect 770 760 810 790
rect 770 740 780 760
rect 800 740 810 760
rect 770 710 810 740
rect 770 690 780 710
rect 800 690 810 710
rect 770 660 810 690
rect 770 640 780 660
rect 800 640 810 660
rect 770 625 810 640
rect 825 860 865 875
rect 825 840 835 860
rect 855 840 865 860
rect 825 810 865 840
rect 825 790 835 810
rect 855 790 865 810
rect 825 760 865 790
rect 825 740 835 760
rect 855 740 865 760
rect 825 710 865 740
rect 825 690 835 710
rect 855 690 865 710
rect 825 660 865 690
rect 825 640 835 660
rect 855 640 865 660
rect 825 625 865 640
rect 880 860 920 875
rect 880 840 890 860
rect 910 840 920 860
rect 880 810 920 840
rect 880 790 890 810
rect 910 790 920 810
rect 880 760 920 790
rect 880 740 890 760
rect 910 740 920 760
rect 880 710 920 740
rect 880 690 890 710
rect 910 690 920 710
rect 880 660 920 690
rect 880 640 890 660
rect 910 640 920 660
rect 880 625 920 640
rect 935 860 975 875
rect 935 840 945 860
rect 965 840 975 860
rect 935 810 975 840
rect 935 790 945 810
rect 965 790 975 810
rect 935 760 975 790
rect 935 740 945 760
rect 965 740 975 760
rect 935 710 975 740
rect 935 690 945 710
rect 965 690 975 710
rect 1095 835 1135 850
rect 1095 815 1105 835
rect 1125 815 1135 835
rect 1095 785 1135 815
rect 1095 765 1105 785
rect 1125 765 1135 785
rect 1095 735 1135 765
rect 1095 715 1105 735
rect 1125 715 1135 735
rect 1095 700 1135 715
rect 1150 835 1190 850
rect 1150 815 1160 835
rect 1180 815 1190 835
rect 1150 785 1190 815
rect 1150 765 1160 785
rect 1180 765 1190 785
rect 1150 735 1190 765
rect 1150 715 1160 735
rect 1180 715 1190 735
rect 1150 700 1190 715
rect 1205 835 1245 850
rect 1205 815 1215 835
rect 1235 815 1245 835
rect 1205 785 1245 815
rect 1205 765 1215 785
rect 1235 765 1245 785
rect 1205 735 1245 765
rect 1205 715 1215 735
rect 1235 715 1245 735
rect 1205 700 1245 715
rect 1260 835 1300 850
rect 1260 815 1270 835
rect 1290 815 1300 835
rect 1260 785 1300 815
rect 1260 765 1270 785
rect 1290 765 1300 785
rect 1260 735 1300 765
rect 1260 715 1270 735
rect 1290 715 1300 735
rect 1260 700 1300 715
rect 1315 835 1355 850
rect 1315 815 1325 835
rect 1345 815 1355 835
rect 1315 785 1355 815
rect 1315 765 1325 785
rect 1345 765 1355 785
rect 1315 735 1355 765
rect 1315 715 1325 735
rect 1345 715 1355 735
rect 1315 700 1355 715
rect 1370 835 1410 850
rect 1370 815 1380 835
rect 1400 815 1410 835
rect 1370 785 1410 815
rect 1370 765 1380 785
rect 1400 765 1410 785
rect 1370 735 1410 765
rect 1370 715 1380 735
rect 1400 715 1410 735
rect 1370 700 1410 715
rect 1425 835 1465 850
rect 1425 815 1435 835
rect 1455 815 1465 835
rect 1425 785 1465 815
rect 1425 765 1435 785
rect 1455 765 1465 785
rect 1425 735 1465 765
rect 1425 715 1435 735
rect 1455 715 1465 735
rect 1425 700 1465 715
rect 1480 835 1520 850
rect 1480 815 1490 835
rect 1510 815 1520 835
rect 1480 785 1520 815
rect 1480 765 1490 785
rect 1510 765 1520 785
rect 1480 735 1520 765
rect 1480 715 1490 735
rect 1510 715 1520 735
rect 1480 700 1520 715
rect 1535 835 1575 850
rect 1535 815 1545 835
rect 1565 815 1575 835
rect 1535 785 1575 815
rect 1535 765 1545 785
rect 1565 765 1575 785
rect 1535 735 1575 765
rect 1535 715 1545 735
rect 1565 715 1575 735
rect 1535 700 1575 715
rect 1590 835 1630 850
rect 1590 815 1600 835
rect 1620 815 1630 835
rect 1590 785 1630 815
rect 1590 765 1600 785
rect 1620 765 1630 785
rect 1590 735 1630 765
rect 1590 715 1600 735
rect 1620 715 1630 735
rect 1590 700 1630 715
rect 1645 835 1685 850
rect 1645 815 1655 835
rect 1675 815 1685 835
rect 1645 785 1685 815
rect 1645 765 1655 785
rect 1675 765 1685 785
rect 1645 735 1685 765
rect 1645 715 1655 735
rect 1675 715 1685 735
rect 1645 700 1685 715
rect 1700 835 1740 850
rect 1700 815 1710 835
rect 1730 815 1740 835
rect 1700 785 1740 815
rect 1700 765 1710 785
rect 1730 765 1740 785
rect 1700 735 1740 765
rect 1700 715 1710 735
rect 1730 715 1740 735
rect 1700 700 1740 715
rect 1755 835 1795 850
rect 1755 815 1765 835
rect 1785 815 1795 835
rect 1755 785 1795 815
rect 1755 765 1765 785
rect 1785 765 1795 785
rect 1755 735 1795 765
rect 1755 715 1765 735
rect 1785 715 1795 735
rect 1755 700 1795 715
rect 935 660 975 690
rect 935 640 945 660
rect 965 640 975 660
rect 935 625 975 640
rect -105 440 -65 455
rect -105 420 -95 440
rect -75 420 -65 440
rect -105 390 -65 420
rect -105 370 -95 390
rect -75 370 -65 390
rect -105 340 -65 370
rect -105 320 -95 340
rect -75 320 -65 340
rect -105 305 -65 320
rect -50 440 -10 455
rect -50 420 -40 440
rect -20 420 -10 440
rect -50 390 -10 420
rect -50 370 -40 390
rect -20 370 -10 390
rect -50 340 -10 370
rect -50 320 -40 340
rect -20 320 -10 340
rect -50 305 -10 320
rect 5 440 45 455
rect 5 420 15 440
rect 35 420 45 440
rect 5 390 45 420
rect 5 370 15 390
rect 35 370 45 390
rect 5 340 45 370
rect 5 320 15 340
rect 35 320 45 340
rect 5 305 45 320
rect 60 440 100 455
rect 60 420 70 440
rect 90 420 100 440
rect 60 390 100 420
rect 60 370 70 390
rect 90 370 100 390
rect 60 340 100 370
rect 60 320 70 340
rect 90 320 100 340
rect 60 305 100 320
rect 115 440 155 455
rect 115 420 125 440
rect 145 420 155 440
rect 115 390 155 420
rect 115 370 125 390
rect 145 370 155 390
rect 115 340 155 370
rect 115 320 125 340
rect 145 320 155 340
rect 115 305 155 320
rect 170 440 210 455
rect 170 420 180 440
rect 200 420 210 440
rect 170 390 210 420
rect 170 370 180 390
rect 200 370 210 390
rect 170 340 210 370
rect 170 320 180 340
rect 200 320 210 340
rect 170 305 210 320
rect 225 440 265 455
rect 225 420 235 440
rect 255 420 265 440
rect 225 390 265 420
rect 225 370 235 390
rect 255 370 265 390
rect 225 340 265 370
rect 225 320 235 340
rect 255 320 265 340
rect 225 305 265 320
rect 280 440 320 455
rect 280 420 290 440
rect 310 420 320 440
rect 280 390 320 420
rect 280 370 290 390
rect 310 370 320 390
rect 280 340 320 370
rect 280 320 290 340
rect 310 320 320 340
rect 280 305 320 320
rect 335 440 375 455
rect 335 420 345 440
rect 365 420 375 440
rect 335 390 375 420
rect 335 370 345 390
rect 365 370 375 390
rect 335 340 375 370
rect 335 320 345 340
rect 365 320 375 340
rect 335 305 375 320
rect 390 440 430 455
rect 390 420 400 440
rect 420 420 430 440
rect 390 390 430 420
rect 390 370 400 390
rect 420 370 430 390
rect 390 340 430 370
rect 390 320 400 340
rect 420 320 430 340
rect 390 305 430 320
rect 445 440 485 455
rect 445 420 455 440
rect 475 420 485 440
rect 445 390 485 420
rect 445 370 455 390
rect 475 370 485 390
rect 445 340 485 370
rect 445 320 455 340
rect 475 320 485 340
rect 445 305 485 320
rect 500 440 540 455
rect 500 420 510 440
rect 530 420 540 440
rect 500 390 540 420
rect 500 370 510 390
rect 530 370 540 390
rect 500 340 540 370
rect 500 320 510 340
rect 530 320 540 340
rect 500 305 540 320
rect 555 440 595 455
rect 555 420 565 440
rect 585 420 595 440
rect 555 390 595 420
rect 555 370 565 390
rect 585 370 595 390
rect 555 340 595 370
rect 555 320 565 340
rect 585 320 595 340
rect 555 305 595 320
rect 715 440 755 455
rect 715 420 725 440
rect 745 420 755 440
rect 715 390 755 420
rect 715 370 725 390
rect 745 370 755 390
rect 715 340 755 370
rect 715 320 725 340
rect 745 320 755 340
rect 715 305 755 320
rect 770 440 810 455
rect 770 420 780 440
rect 800 420 810 440
rect 770 390 810 420
rect 770 370 780 390
rect 800 370 810 390
rect 770 340 810 370
rect 770 320 780 340
rect 800 320 810 340
rect 770 305 810 320
rect 825 440 865 455
rect 825 420 835 440
rect 855 420 865 440
rect 825 390 865 420
rect 825 370 835 390
rect 855 370 865 390
rect 825 340 865 370
rect 825 320 835 340
rect 855 320 865 340
rect 825 305 865 320
rect 880 440 920 455
rect 880 420 890 440
rect 910 420 920 440
rect 880 390 920 420
rect 880 370 890 390
rect 910 370 920 390
rect 880 340 920 370
rect 880 320 890 340
rect 910 320 920 340
rect 880 305 920 320
rect 935 440 975 455
rect 935 420 945 440
rect 965 420 975 440
rect 935 390 975 420
rect 935 370 945 390
rect 965 370 975 390
rect 935 340 975 370
rect 935 320 945 340
rect 965 320 975 340
rect 935 305 975 320
rect 1095 440 1135 455
rect 1095 420 1105 440
rect 1125 420 1135 440
rect 1095 390 1135 420
rect 1095 370 1105 390
rect 1125 370 1135 390
rect 1095 340 1135 370
rect 1095 320 1105 340
rect 1125 320 1135 340
rect 1095 305 1135 320
rect 1150 440 1190 455
rect 1150 420 1160 440
rect 1180 420 1190 440
rect 1150 390 1190 420
rect 1150 370 1160 390
rect 1180 370 1190 390
rect 1150 340 1190 370
rect 1150 320 1160 340
rect 1180 320 1190 340
rect 1150 305 1190 320
rect 1205 440 1245 455
rect 1205 420 1215 440
rect 1235 420 1245 440
rect 1205 390 1245 420
rect 1205 370 1215 390
rect 1235 370 1245 390
rect 1205 340 1245 370
rect 1205 320 1215 340
rect 1235 320 1245 340
rect 1205 305 1245 320
rect 1260 440 1300 455
rect 1260 420 1270 440
rect 1290 420 1300 440
rect 1260 390 1300 420
rect 1260 370 1270 390
rect 1290 370 1300 390
rect 1260 340 1300 370
rect 1260 320 1270 340
rect 1290 320 1300 340
rect 1260 305 1300 320
rect 1315 440 1355 455
rect 1315 420 1325 440
rect 1345 420 1355 440
rect 1315 390 1355 420
rect 1315 370 1325 390
rect 1345 370 1355 390
rect 1315 340 1355 370
rect 1315 320 1325 340
rect 1345 320 1355 340
rect 1315 305 1355 320
rect 1370 440 1410 455
rect 1370 420 1380 440
rect 1400 420 1410 440
rect 1370 390 1410 420
rect 1370 370 1380 390
rect 1400 370 1410 390
rect 1370 340 1410 370
rect 1370 320 1380 340
rect 1400 320 1410 340
rect 1370 305 1410 320
rect 1425 440 1465 455
rect 1425 420 1435 440
rect 1455 420 1465 440
rect 1425 390 1465 420
rect 1425 370 1435 390
rect 1455 370 1465 390
rect 1425 340 1465 370
rect 1425 320 1435 340
rect 1455 320 1465 340
rect 1425 305 1465 320
rect 1480 440 1520 455
rect 1480 420 1490 440
rect 1510 420 1520 440
rect 1480 390 1520 420
rect 1480 370 1490 390
rect 1510 370 1520 390
rect 1480 340 1520 370
rect 1480 320 1490 340
rect 1510 320 1520 340
rect 1480 305 1520 320
rect 1535 440 1575 455
rect 1535 420 1545 440
rect 1565 420 1575 440
rect 1535 390 1575 420
rect 1535 370 1545 390
rect 1565 370 1575 390
rect 1535 340 1575 370
rect 1535 320 1545 340
rect 1565 320 1575 340
rect 1535 305 1575 320
rect 1590 440 1630 455
rect 1590 420 1600 440
rect 1620 420 1630 440
rect 1590 390 1630 420
rect 1590 370 1600 390
rect 1620 370 1630 390
rect 1590 340 1630 370
rect 1590 320 1600 340
rect 1620 320 1630 340
rect 1590 305 1630 320
rect 1645 440 1685 455
rect 1645 420 1655 440
rect 1675 420 1685 440
rect 1645 390 1685 420
rect 1645 370 1655 390
rect 1675 370 1685 390
rect 1645 340 1685 370
rect 1645 320 1655 340
rect 1675 320 1685 340
rect 1645 305 1685 320
rect 1700 440 1740 455
rect 1700 420 1710 440
rect 1730 420 1740 440
rect 1700 390 1740 420
rect 1700 370 1710 390
rect 1730 370 1740 390
rect 1700 340 1740 370
rect 1700 320 1710 340
rect 1730 320 1740 340
rect 1700 305 1740 320
rect 1755 440 1795 455
rect 1755 420 1765 440
rect 1785 420 1795 440
rect 1755 390 1795 420
rect 1755 370 1765 390
rect 1785 370 1795 390
rect 1755 340 1795 370
rect 1755 320 1765 340
rect 1785 320 1795 340
rect 1755 305 1795 320
rect -1135 215 -1095 230
rect -1135 195 -1125 215
rect -1105 195 -1095 215
rect -1135 165 -1095 195
rect -1135 145 -1125 165
rect -1105 145 -1095 165
rect -1135 115 -1095 145
rect -1135 95 -1125 115
rect -1105 95 -1095 115
rect -1135 65 -1095 95
rect -1135 45 -1125 65
rect -1105 45 -1095 65
rect -1135 15 -1095 45
rect -1135 -5 -1125 15
rect -1105 -5 -1095 15
rect -1135 -35 -1095 -5
rect -1135 -55 -1125 -35
rect -1105 -55 -1095 -35
rect -1135 -70 -1095 -55
rect -1080 215 -1040 230
rect -1080 195 -1070 215
rect -1050 195 -1040 215
rect -1080 165 -1040 195
rect -1080 145 -1070 165
rect -1050 145 -1040 165
rect -1080 115 -1040 145
rect -1080 95 -1070 115
rect -1050 95 -1040 115
rect -1080 65 -1040 95
rect -1080 45 -1070 65
rect -1050 45 -1040 65
rect -1080 15 -1040 45
rect -1080 -5 -1070 15
rect -1050 -5 -1040 15
rect -1080 -35 -1040 -5
rect -1080 -55 -1070 -35
rect -1050 -55 -1040 -35
rect -1080 -70 -1040 -55
rect -1025 215 -985 230
rect -1025 195 -1015 215
rect -995 195 -985 215
rect -1025 165 -985 195
rect -1025 145 -1015 165
rect -995 145 -985 165
rect -1025 115 -985 145
rect -1025 95 -1015 115
rect -995 95 -985 115
rect -1025 65 -985 95
rect -1025 45 -1015 65
rect -995 45 -985 65
rect -1025 15 -985 45
rect -1025 -5 -1015 15
rect -995 -5 -985 15
rect -1025 -35 -985 -5
rect -1025 -55 -1015 -35
rect -995 -55 -985 -35
rect -1025 -70 -985 -55
rect -970 215 -930 230
rect -970 195 -960 215
rect -940 195 -930 215
rect -970 165 -930 195
rect -970 145 -960 165
rect -940 145 -930 165
rect -970 115 -930 145
rect -970 95 -960 115
rect -940 95 -930 115
rect -970 65 -930 95
rect -970 45 -960 65
rect -940 45 -930 65
rect -970 15 -930 45
rect -970 -5 -960 15
rect -940 -5 -930 15
rect -970 -35 -930 -5
rect -970 -55 -960 -35
rect -940 -55 -930 -35
rect -970 -70 -930 -55
rect -915 215 -875 230
rect -915 195 -905 215
rect -885 195 -875 215
rect -915 165 -875 195
rect -915 145 -905 165
rect -885 145 -875 165
rect -915 115 -875 145
rect -915 95 -905 115
rect -885 95 -875 115
rect -915 65 -875 95
rect -915 45 -905 65
rect -885 45 -875 65
rect -915 15 -875 45
rect -915 -5 -905 15
rect -885 -5 -875 15
rect -915 -35 -875 -5
rect -915 -55 -905 -35
rect -885 -55 -875 -35
rect -915 -70 -875 -55
rect -860 215 -820 230
rect -860 195 -850 215
rect -830 195 -820 215
rect -860 165 -820 195
rect -860 145 -850 165
rect -830 145 -820 165
rect -860 115 -820 145
rect -860 95 -850 115
rect -830 95 -820 115
rect -860 65 -820 95
rect -860 45 -850 65
rect -830 45 -820 65
rect -860 15 -820 45
rect -860 -5 -850 15
rect -830 -5 -820 15
rect -860 -35 -820 -5
rect -860 -55 -850 -35
rect -830 -55 -820 -35
rect -860 -70 -820 -55
rect -805 215 -765 230
rect -805 195 -795 215
rect -775 195 -765 215
rect -805 165 -765 195
rect -805 145 -795 165
rect -775 145 -765 165
rect -805 115 -765 145
rect -805 95 -795 115
rect -775 95 -765 115
rect -805 65 -765 95
rect -805 45 -795 65
rect -775 45 -765 65
rect -805 15 -765 45
rect -805 -5 -795 15
rect -775 -5 -765 15
rect -805 -35 -765 -5
rect -805 -55 -795 -35
rect -775 -55 -765 -35
rect -805 -70 -765 -55
rect -750 215 -710 230
rect -750 195 -740 215
rect -720 195 -710 215
rect -750 165 -710 195
rect -750 145 -740 165
rect -720 145 -710 165
rect -750 115 -710 145
rect -750 95 -740 115
rect -720 95 -710 115
rect -750 65 -710 95
rect -750 45 -740 65
rect -720 45 -710 65
rect -750 15 -710 45
rect -750 -5 -740 15
rect -720 -5 -710 15
rect -750 -35 -710 -5
rect -750 -55 -740 -35
rect -720 -55 -710 -35
rect -750 -70 -710 -55
rect -695 215 -655 230
rect -695 195 -685 215
rect -665 195 -655 215
rect -695 165 -655 195
rect -695 145 -685 165
rect -665 145 -655 165
rect -695 115 -655 145
rect -695 95 -685 115
rect -665 95 -655 115
rect -695 65 -655 95
rect -695 45 -685 65
rect -665 45 -655 65
rect -695 15 -655 45
rect -695 -5 -685 15
rect -665 -5 -655 15
rect -695 -35 -655 -5
rect -695 -55 -685 -35
rect -665 -55 -655 -35
rect -695 -70 -655 -55
rect -640 215 -600 230
rect -640 195 -630 215
rect -610 195 -600 215
rect -640 165 -600 195
rect -640 145 -630 165
rect -610 145 -600 165
rect -640 115 -600 145
rect -640 95 -630 115
rect -610 95 -600 115
rect -640 65 -600 95
rect -640 45 -630 65
rect -610 45 -600 65
rect -640 15 -600 45
rect -640 -5 -630 15
rect -610 -5 -600 15
rect -640 -35 -600 -5
rect -640 -55 -630 -35
rect -610 -55 -600 -35
rect -640 -70 -600 -55
rect -585 215 -545 230
rect -585 195 -575 215
rect -555 195 -545 215
rect -585 165 -545 195
rect -585 145 -575 165
rect -555 145 -545 165
rect -585 115 -545 145
rect -585 95 -575 115
rect -555 95 -545 115
rect -585 65 -545 95
rect -585 45 -575 65
rect -555 45 -545 65
rect -585 15 -545 45
rect -585 -5 -575 15
rect -555 -5 -545 15
rect -585 -35 -545 -5
rect -585 -55 -575 -35
rect -555 -55 -545 -35
rect -585 -70 -545 -55
rect -530 215 -490 230
rect -530 195 -520 215
rect -500 195 -490 215
rect -530 165 -490 195
rect -530 145 -520 165
rect -500 145 -490 165
rect -530 115 -490 145
rect -530 95 -520 115
rect -500 95 -490 115
rect -530 65 -490 95
rect -530 45 -520 65
rect -500 45 -490 65
rect -530 15 -490 45
rect -530 -5 -520 15
rect -500 -5 -490 15
rect -530 -35 -490 -5
rect -530 -55 -520 -35
rect -500 -55 -490 -35
rect -530 -70 -490 -55
rect -475 215 -435 230
rect -475 195 -465 215
rect -445 195 -435 215
rect -475 165 -435 195
rect -475 145 -465 165
rect -445 145 -435 165
rect -475 115 -435 145
rect -475 95 -465 115
rect -445 95 -435 115
rect -475 65 -435 95
rect -475 45 -465 65
rect -445 45 -435 65
rect -475 15 -435 45
rect 2125 215 2165 230
rect 2125 195 2135 215
rect 2155 195 2165 215
rect 2125 165 2165 195
rect 2125 145 2135 165
rect 2155 145 2165 165
rect 2125 115 2165 145
rect 2125 95 2135 115
rect 2155 95 2165 115
rect 2125 65 2165 95
rect 2125 45 2135 65
rect 2155 45 2165 65
rect -475 -5 -465 15
rect -445 -5 -435 15
rect -475 -35 -435 -5
rect 2125 15 2165 45
rect 2125 -5 2135 15
rect 2155 -5 2165 15
rect -475 -55 -465 -35
rect -445 -55 -435 -35
rect 2125 -35 2165 -5
rect -475 -70 -435 -55
rect 715 -55 755 -40
rect 715 -75 725 -55
rect 745 -75 755 -55
rect 715 -105 755 -75
rect 715 -125 725 -105
rect 745 -125 755 -105
rect 715 -155 755 -125
rect 715 -175 725 -155
rect 745 -175 755 -155
rect 715 -205 755 -175
rect 715 -225 725 -205
rect 745 -225 755 -205
rect 715 -255 755 -225
rect 715 -275 725 -255
rect 745 -275 755 -255
rect 715 -290 755 -275
rect 770 -55 810 -40
rect 770 -75 780 -55
rect 800 -75 810 -55
rect 770 -105 810 -75
rect 770 -125 780 -105
rect 800 -125 810 -105
rect 770 -155 810 -125
rect 770 -175 780 -155
rect 800 -175 810 -155
rect 770 -205 810 -175
rect 770 -225 780 -205
rect 800 -225 810 -205
rect 770 -255 810 -225
rect 770 -275 780 -255
rect 800 -275 810 -255
rect 770 -290 810 -275
rect 825 -55 865 -40
rect 825 -75 835 -55
rect 855 -75 865 -55
rect 825 -105 865 -75
rect 825 -125 835 -105
rect 855 -125 865 -105
rect 825 -155 865 -125
rect 825 -175 835 -155
rect 855 -175 865 -155
rect 825 -205 865 -175
rect 825 -225 835 -205
rect 855 -225 865 -205
rect 825 -255 865 -225
rect 825 -275 835 -255
rect 855 -275 865 -255
rect 825 -290 865 -275
rect 880 -55 920 -40
rect 880 -75 890 -55
rect 910 -75 920 -55
rect 880 -105 920 -75
rect 880 -125 890 -105
rect 910 -125 920 -105
rect 880 -155 920 -125
rect 880 -175 890 -155
rect 910 -175 920 -155
rect 880 -205 920 -175
rect 880 -225 890 -205
rect 910 -225 920 -205
rect 880 -255 920 -225
rect 880 -275 890 -255
rect 910 -275 920 -255
rect 880 -290 920 -275
rect 935 -55 975 -40
rect 935 -75 945 -55
rect 965 -75 975 -55
rect 2125 -55 2135 -35
rect 2155 -55 2165 -35
rect 2125 -70 2165 -55
rect 2180 215 2220 230
rect 2180 195 2190 215
rect 2210 195 2220 215
rect 2180 165 2220 195
rect 2180 145 2190 165
rect 2210 145 2220 165
rect 2180 115 2220 145
rect 2180 95 2190 115
rect 2210 95 2220 115
rect 2180 65 2220 95
rect 2180 45 2190 65
rect 2210 45 2220 65
rect 2180 15 2220 45
rect 2180 -5 2190 15
rect 2210 -5 2220 15
rect 2180 -35 2220 -5
rect 2180 -55 2190 -35
rect 2210 -55 2220 -35
rect 2180 -70 2220 -55
rect 2235 215 2275 230
rect 2235 195 2245 215
rect 2265 195 2275 215
rect 2235 165 2275 195
rect 2235 145 2245 165
rect 2265 145 2275 165
rect 2235 115 2275 145
rect 2235 95 2245 115
rect 2265 95 2275 115
rect 2235 65 2275 95
rect 2235 45 2245 65
rect 2265 45 2275 65
rect 2235 15 2275 45
rect 2235 -5 2245 15
rect 2265 -5 2275 15
rect 2235 -35 2275 -5
rect 2235 -55 2245 -35
rect 2265 -55 2275 -35
rect 2235 -70 2275 -55
rect 2290 215 2330 230
rect 2290 195 2300 215
rect 2320 195 2330 215
rect 2290 165 2330 195
rect 2290 145 2300 165
rect 2320 145 2330 165
rect 2290 115 2330 145
rect 2290 95 2300 115
rect 2320 95 2330 115
rect 2290 65 2330 95
rect 2290 45 2300 65
rect 2320 45 2330 65
rect 2290 15 2330 45
rect 2290 -5 2300 15
rect 2320 -5 2330 15
rect 2290 -35 2330 -5
rect 2290 -55 2300 -35
rect 2320 -55 2330 -35
rect 2290 -70 2330 -55
rect 2345 215 2385 230
rect 2345 195 2355 215
rect 2375 195 2385 215
rect 2345 165 2385 195
rect 2345 145 2355 165
rect 2375 145 2385 165
rect 2345 115 2385 145
rect 2345 95 2355 115
rect 2375 95 2385 115
rect 2345 65 2385 95
rect 2345 45 2355 65
rect 2375 45 2385 65
rect 2345 15 2385 45
rect 2345 -5 2355 15
rect 2375 -5 2385 15
rect 2345 -35 2385 -5
rect 2345 -55 2355 -35
rect 2375 -55 2385 -35
rect 2345 -70 2385 -55
rect 2400 215 2440 230
rect 2400 195 2410 215
rect 2430 195 2440 215
rect 2400 165 2440 195
rect 2400 145 2410 165
rect 2430 145 2440 165
rect 2400 115 2440 145
rect 2400 95 2410 115
rect 2430 95 2440 115
rect 2400 65 2440 95
rect 2400 45 2410 65
rect 2430 45 2440 65
rect 2400 15 2440 45
rect 2400 -5 2410 15
rect 2430 -5 2440 15
rect 2400 -35 2440 -5
rect 2400 -55 2410 -35
rect 2430 -55 2440 -35
rect 2400 -70 2440 -55
rect 2455 215 2495 230
rect 2455 195 2465 215
rect 2485 195 2495 215
rect 2455 165 2495 195
rect 2455 145 2465 165
rect 2485 145 2495 165
rect 2455 115 2495 145
rect 2455 95 2465 115
rect 2485 95 2495 115
rect 2455 65 2495 95
rect 2455 45 2465 65
rect 2485 45 2495 65
rect 2455 15 2495 45
rect 2455 -5 2465 15
rect 2485 -5 2495 15
rect 2455 -35 2495 -5
rect 2455 -55 2465 -35
rect 2485 -55 2495 -35
rect 2455 -70 2495 -55
rect 2510 215 2550 230
rect 2510 195 2520 215
rect 2540 195 2550 215
rect 2510 165 2550 195
rect 2510 145 2520 165
rect 2540 145 2550 165
rect 2510 115 2550 145
rect 2510 95 2520 115
rect 2540 95 2550 115
rect 2510 65 2550 95
rect 2510 45 2520 65
rect 2540 45 2550 65
rect 2510 15 2550 45
rect 2510 -5 2520 15
rect 2540 -5 2550 15
rect 2510 -35 2550 -5
rect 2510 -55 2520 -35
rect 2540 -55 2550 -35
rect 2510 -70 2550 -55
rect 2565 215 2605 230
rect 2565 195 2575 215
rect 2595 195 2605 215
rect 2565 165 2605 195
rect 2565 145 2575 165
rect 2595 145 2605 165
rect 2565 115 2605 145
rect 2565 95 2575 115
rect 2595 95 2605 115
rect 2565 65 2605 95
rect 2565 45 2575 65
rect 2595 45 2605 65
rect 2565 15 2605 45
rect 2565 -5 2575 15
rect 2595 -5 2605 15
rect 2565 -35 2605 -5
rect 2565 -55 2575 -35
rect 2595 -55 2605 -35
rect 2565 -70 2605 -55
rect 2620 215 2660 230
rect 2620 195 2630 215
rect 2650 195 2660 215
rect 2620 165 2660 195
rect 2620 145 2630 165
rect 2650 145 2660 165
rect 2620 115 2660 145
rect 2620 95 2630 115
rect 2650 95 2660 115
rect 2620 65 2660 95
rect 2620 45 2630 65
rect 2650 45 2660 65
rect 2620 15 2660 45
rect 2620 -5 2630 15
rect 2650 -5 2660 15
rect 2620 -35 2660 -5
rect 2620 -55 2630 -35
rect 2650 -55 2660 -35
rect 2620 -70 2660 -55
rect 2675 215 2715 230
rect 2675 195 2685 215
rect 2705 195 2715 215
rect 2675 165 2715 195
rect 2675 145 2685 165
rect 2705 145 2715 165
rect 2675 115 2715 145
rect 2675 95 2685 115
rect 2705 95 2715 115
rect 2675 65 2715 95
rect 2675 45 2685 65
rect 2705 45 2715 65
rect 2675 15 2715 45
rect 2675 -5 2685 15
rect 2705 -5 2715 15
rect 2675 -35 2715 -5
rect 2675 -55 2685 -35
rect 2705 -55 2715 -35
rect 2675 -70 2715 -55
rect 2730 215 2770 230
rect 2730 195 2740 215
rect 2760 195 2770 215
rect 2730 165 2770 195
rect 2730 145 2740 165
rect 2760 145 2770 165
rect 2730 115 2770 145
rect 2730 95 2740 115
rect 2760 95 2770 115
rect 2730 65 2770 95
rect 2730 45 2740 65
rect 2760 45 2770 65
rect 2730 15 2770 45
rect 2730 -5 2740 15
rect 2760 -5 2770 15
rect 2730 -35 2770 -5
rect 2730 -55 2740 -35
rect 2760 -55 2770 -35
rect 2730 -70 2770 -55
rect 2785 215 2825 230
rect 2785 195 2795 215
rect 2815 195 2825 215
rect 2785 165 2825 195
rect 2785 145 2795 165
rect 2815 145 2825 165
rect 2785 115 2825 145
rect 2785 95 2795 115
rect 2815 95 2825 115
rect 2785 65 2825 95
rect 2785 45 2795 65
rect 2815 45 2825 65
rect 2785 15 2825 45
rect 2785 -5 2795 15
rect 2815 -5 2825 15
rect 2785 -35 2825 -5
rect 2785 -55 2795 -35
rect 2815 -55 2825 -35
rect 2785 -70 2825 -55
rect 935 -105 975 -75
rect 935 -125 945 -105
rect 965 -125 975 -105
rect 935 -155 975 -125
rect 935 -175 945 -155
rect 965 -175 975 -155
rect 935 -205 975 -175
rect 935 -225 945 -205
rect 965 -225 975 -205
rect 935 -255 975 -225
rect 935 -275 945 -255
rect 965 -275 975 -255
rect 935 -290 975 -275
rect -1025 -370 -985 -355
rect -1025 -390 -1015 -370
rect -995 -390 -985 -370
rect -1025 -420 -985 -390
rect -1025 -440 -1015 -420
rect -995 -440 -985 -420
rect -1025 -470 -985 -440
rect -1025 -490 -1015 -470
rect -995 -490 -985 -470
rect -1025 -520 -985 -490
rect -1025 -540 -1015 -520
rect -995 -540 -985 -520
rect -1025 -570 -985 -540
rect -1025 -590 -1015 -570
rect -995 -590 -985 -570
rect -1025 -620 -985 -590
rect -1025 -640 -1015 -620
rect -995 -640 -985 -620
rect -1025 -670 -985 -640
rect -1025 -690 -1015 -670
rect -995 -690 -985 -670
rect -1025 -720 -985 -690
rect -1025 -740 -1015 -720
rect -995 -740 -985 -720
rect -1025 -770 -985 -740
rect -1025 -790 -1015 -770
rect -995 -790 -985 -770
rect -1025 -820 -985 -790
rect -1025 -840 -1015 -820
rect -995 -840 -985 -820
rect -1025 -870 -985 -840
rect -1025 -890 -1015 -870
rect -995 -890 -985 -870
rect -1025 -920 -985 -890
rect -1025 -940 -1015 -920
rect -995 -940 -985 -920
rect -1025 -970 -985 -940
rect -1025 -990 -1015 -970
rect -995 -990 -985 -970
rect -1025 -1020 -985 -990
rect -1025 -1040 -1015 -1020
rect -995 -1040 -985 -1020
rect -1025 -1055 -985 -1040
rect -925 -370 -885 -355
rect -925 -390 -915 -370
rect -895 -390 -885 -370
rect -925 -420 -885 -390
rect -925 -440 -915 -420
rect -895 -440 -885 -420
rect -925 -470 -885 -440
rect -925 -490 -915 -470
rect -895 -490 -885 -470
rect -925 -520 -885 -490
rect -925 -540 -915 -520
rect -895 -540 -885 -520
rect -925 -570 -885 -540
rect -925 -590 -915 -570
rect -895 -590 -885 -570
rect -925 -620 -885 -590
rect -925 -640 -915 -620
rect -895 -640 -885 -620
rect -925 -670 -885 -640
rect -925 -690 -915 -670
rect -895 -690 -885 -670
rect -925 -720 -885 -690
rect -925 -740 -915 -720
rect -895 -740 -885 -720
rect -925 -770 -885 -740
rect -925 -790 -915 -770
rect -895 -790 -885 -770
rect -925 -820 -885 -790
rect -925 -840 -915 -820
rect -895 -840 -885 -820
rect -925 -870 -885 -840
rect -925 -890 -915 -870
rect -895 -890 -885 -870
rect -925 -920 -885 -890
rect -925 -940 -915 -920
rect -895 -940 -885 -920
rect -925 -970 -885 -940
rect -925 -990 -915 -970
rect -895 -990 -885 -970
rect -925 -1020 -885 -990
rect -925 -1040 -915 -1020
rect -895 -1040 -885 -1020
rect -925 -1055 -885 -1040
rect -825 -370 -785 -355
rect -825 -390 -815 -370
rect -795 -390 -785 -370
rect -825 -420 -785 -390
rect -825 -440 -815 -420
rect -795 -440 -785 -420
rect -825 -470 -785 -440
rect -825 -490 -815 -470
rect -795 -490 -785 -470
rect -825 -520 -785 -490
rect -825 -540 -815 -520
rect -795 -540 -785 -520
rect -825 -570 -785 -540
rect -825 -590 -815 -570
rect -795 -590 -785 -570
rect -825 -620 -785 -590
rect -825 -640 -815 -620
rect -795 -640 -785 -620
rect -825 -670 -785 -640
rect -825 -690 -815 -670
rect -795 -690 -785 -670
rect -825 -720 -785 -690
rect -825 -740 -815 -720
rect -795 -740 -785 -720
rect -825 -770 -785 -740
rect -825 -790 -815 -770
rect -795 -790 -785 -770
rect -825 -820 -785 -790
rect -825 -840 -815 -820
rect -795 -840 -785 -820
rect -825 -870 -785 -840
rect -825 -890 -815 -870
rect -795 -890 -785 -870
rect -825 -920 -785 -890
rect -825 -940 -815 -920
rect -795 -940 -785 -920
rect -825 -970 -785 -940
rect -825 -990 -815 -970
rect -795 -990 -785 -970
rect -825 -1020 -785 -990
rect -825 -1040 -815 -1020
rect -795 -1040 -785 -1020
rect -825 -1055 -785 -1040
rect -725 -370 -685 -355
rect -725 -390 -715 -370
rect -695 -390 -685 -370
rect -725 -420 -685 -390
rect -725 -440 -715 -420
rect -695 -440 -685 -420
rect -725 -470 -685 -440
rect -725 -490 -715 -470
rect -695 -490 -685 -470
rect -725 -520 -685 -490
rect -725 -540 -715 -520
rect -695 -540 -685 -520
rect -725 -570 -685 -540
rect -725 -590 -715 -570
rect -695 -590 -685 -570
rect -725 -620 -685 -590
rect -725 -640 -715 -620
rect -695 -640 -685 -620
rect -725 -670 -685 -640
rect -725 -690 -715 -670
rect -695 -690 -685 -670
rect -725 -720 -685 -690
rect -725 -740 -715 -720
rect -695 -740 -685 -720
rect -725 -770 -685 -740
rect -725 -790 -715 -770
rect -695 -790 -685 -770
rect -725 -820 -685 -790
rect -725 -840 -715 -820
rect -695 -840 -685 -820
rect -725 -870 -685 -840
rect -725 -890 -715 -870
rect -695 -890 -685 -870
rect -725 -920 -685 -890
rect -725 -940 -715 -920
rect -695 -940 -685 -920
rect -725 -970 -685 -940
rect -725 -990 -715 -970
rect -695 -990 -685 -970
rect -725 -1020 -685 -990
rect -725 -1040 -715 -1020
rect -695 -1040 -685 -1020
rect -725 -1055 -685 -1040
rect -625 -370 -585 -355
rect -625 -390 -615 -370
rect -595 -390 -585 -370
rect -625 -420 -585 -390
rect -625 -440 -615 -420
rect -595 -440 -585 -420
rect -625 -470 -585 -440
rect -625 -490 -615 -470
rect -595 -490 -585 -470
rect -625 -520 -585 -490
rect -625 -540 -615 -520
rect -595 -540 -585 -520
rect -625 -570 -585 -540
rect -625 -590 -615 -570
rect -595 -590 -585 -570
rect -625 -620 -585 -590
rect -625 -640 -615 -620
rect -595 -640 -585 -620
rect -625 -670 -585 -640
rect -625 -690 -615 -670
rect -595 -690 -585 -670
rect -625 -720 -585 -690
rect -625 -740 -615 -720
rect -595 -740 -585 -720
rect -625 -770 -585 -740
rect -625 -790 -615 -770
rect -595 -790 -585 -770
rect -625 -820 -585 -790
rect -625 -840 -615 -820
rect -595 -840 -585 -820
rect -625 -870 -585 -840
rect -625 -890 -615 -870
rect -595 -890 -585 -870
rect -625 -920 -585 -890
rect -625 -940 -615 -920
rect -595 -940 -585 -920
rect -625 -970 -585 -940
rect -625 -990 -615 -970
rect -595 -990 -585 -970
rect -625 -1020 -585 -990
rect -625 -1040 -615 -1020
rect -595 -1040 -585 -1020
rect -625 -1055 -585 -1040
rect -525 -370 -485 -355
rect -525 -390 -515 -370
rect -495 -390 -485 -370
rect -525 -420 -485 -390
rect -525 -440 -515 -420
rect -495 -440 -485 -420
rect -525 -470 -485 -440
rect -525 -490 -515 -470
rect -495 -490 -485 -470
rect -525 -520 -485 -490
rect -525 -540 -515 -520
rect -495 -540 -485 -520
rect -525 -570 -485 -540
rect -525 -590 -515 -570
rect -495 -590 -485 -570
rect -525 -620 -485 -590
rect -525 -640 -515 -620
rect -495 -640 -485 -620
rect -525 -670 -485 -640
rect -525 -690 -515 -670
rect -495 -690 -485 -670
rect -525 -720 -485 -690
rect -525 -740 -515 -720
rect -495 -740 -485 -720
rect -525 -770 -485 -740
rect -525 -790 -515 -770
rect -495 -790 -485 -770
rect -525 -820 -485 -790
rect -525 -840 -515 -820
rect -495 -840 -485 -820
rect -525 -870 -485 -840
rect -525 -890 -515 -870
rect -495 -890 -485 -870
rect -525 -920 -485 -890
rect -525 -940 -515 -920
rect -495 -940 -485 -920
rect -525 -970 -485 -940
rect -525 -990 -515 -970
rect -495 -990 -485 -970
rect -525 -1020 -485 -990
rect -525 -1040 -515 -1020
rect -495 -1040 -485 -1020
rect -525 -1055 -485 -1040
rect -425 -370 -385 -355
rect -425 -390 -415 -370
rect -395 -390 -385 -370
rect -425 -420 -385 -390
rect -425 -440 -415 -420
rect -395 -440 -385 -420
rect -425 -470 -385 -440
rect -425 -490 -415 -470
rect -395 -490 -385 -470
rect 2075 -370 2115 -355
rect 2075 -390 2085 -370
rect 2105 -390 2115 -370
rect 2075 -420 2115 -390
rect 2075 -440 2085 -420
rect 2105 -440 2115 -420
rect 2075 -470 2115 -440
rect -425 -520 -385 -490
rect 2075 -490 2085 -470
rect 2105 -490 2115 -470
rect -425 -540 -415 -520
rect -395 -540 -385 -520
rect 2075 -520 2115 -490
rect -425 -570 -385 -540
rect -425 -590 -415 -570
rect -395 -590 -385 -570
rect -425 -620 -385 -590
rect -425 -640 -415 -620
rect -395 -640 -385 -620
rect -425 -670 -385 -640
rect -425 -690 -415 -670
rect -395 -690 -385 -670
rect -425 -720 -385 -690
rect -425 -740 -415 -720
rect -395 -740 -385 -720
rect -425 -770 -385 -740
rect -425 -790 -415 -770
rect -395 -790 -385 -770
rect 275 -550 315 -535
rect 275 -570 285 -550
rect 305 -570 315 -550
rect 275 -600 315 -570
rect 275 -620 285 -600
rect 305 -620 315 -600
rect 275 -650 315 -620
rect 275 -670 285 -650
rect 305 -670 315 -650
rect 275 -700 315 -670
rect 275 -720 285 -700
rect 305 -720 315 -700
rect 275 -750 315 -720
rect 275 -770 285 -750
rect 305 -770 315 -750
rect 275 -785 315 -770
rect 330 -550 370 -535
rect 330 -570 340 -550
rect 360 -570 370 -550
rect 330 -600 370 -570
rect 330 -620 340 -600
rect 360 -620 370 -600
rect 330 -650 370 -620
rect 330 -670 340 -650
rect 360 -670 370 -650
rect 330 -700 370 -670
rect 330 -720 340 -700
rect 360 -720 370 -700
rect 330 -750 370 -720
rect 330 -770 340 -750
rect 360 -770 370 -750
rect 330 -785 370 -770
rect 385 -550 425 -535
rect 385 -570 395 -550
rect 415 -570 425 -550
rect 385 -600 425 -570
rect 385 -620 395 -600
rect 415 -620 425 -600
rect 385 -650 425 -620
rect 385 -670 395 -650
rect 415 -670 425 -650
rect 385 -700 425 -670
rect 385 -720 395 -700
rect 415 -720 425 -700
rect 385 -750 425 -720
rect 385 -770 395 -750
rect 415 -770 425 -750
rect 385 -785 425 -770
rect 440 -550 480 -535
rect 440 -570 450 -550
rect 470 -570 480 -550
rect 440 -600 480 -570
rect 440 -620 450 -600
rect 470 -620 480 -600
rect 440 -650 480 -620
rect 440 -670 450 -650
rect 470 -670 480 -650
rect 440 -700 480 -670
rect 440 -720 450 -700
rect 470 -720 480 -700
rect 440 -750 480 -720
rect 440 -770 450 -750
rect 470 -770 480 -750
rect 440 -785 480 -770
rect 495 -550 535 -535
rect 495 -570 505 -550
rect 525 -570 535 -550
rect 495 -600 535 -570
rect 495 -620 505 -600
rect 525 -620 535 -600
rect 495 -650 535 -620
rect 495 -670 505 -650
rect 525 -670 535 -650
rect 495 -700 535 -670
rect 495 -720 505 -700
rect 525 -720 535 -700
rect 495 -750 535 -720
rect 495 -770 505 -750
rect 525 -770 535 -750
rect 495 -785 535 -770
rect 550 -550 590 -535
rect 550 -570 560 -550
rect 580 -570 590 -550
rect 550 -600 590 -570
rect 550 -620 560 -600
rect 580 -620 590 -600
rect 550 -650 590 -620
rect 550 -670 560 -650
rect 580 -670 590 -650
rect 550 -700 590 -670
rect 550 -720 560 -700
rect 580 -720 590 -700
rect 550 -750 590 -720
rect 550 -770 560 -750
rect 580 -770 590 -750
rect 550 -785 590 -770
rect 605 -550 645 -535
rect 605 -570 615 -550
rect 635 -570 645 -550
rect 605 -600 645 -570
rect 605 -620 615 -600
rect 635 -620 645 -600
rect 605 -650 645 -620
rect 605 -670 615 -650
rect 635 -670 645 -650
rect 605 -700 645 -670
rect 605 -720 615 -700
rect 635 -720 645 -700
rect 605 -750 645 -720
rect 605 -770 615 -750
rect 635 -770 645 -750
rect 605 -785 645 -770
rect 660 -550 700 -535
rect 660 -570 670 -550
rect 690 -570 700 -550
rect 660 -600 700 -570
rect 660 -620 670 -600
rect 690 -620 700 -600
rect 660 -650 700 -620
rect 660 -670 670 -650
rect 690 -670 700 -650
rect 660 -700 700 -670
rect 660 -720 670 -700
rect 690 -720 700 -700
rect 660 -750 700 -720
rect 660 -770 670 -750
rect 690 -770 700 -750
rect 660 -785 700 -770
rect 715 -550 755 -535
rect 715 -570 725 -550
rect 745 -570 755 -550
rect 715 -600 755 -570
rect 715 -620 725 -600
rect 745 -620 755 -600
rect 715 -650 755 -620
rect 715 -670 725 -650
rect 745 -670 755 -650
rect 715 -700 755 -670
rect 715 -720 725 -700
rect 745 -720 755 -700
rect 715 -750 755 -720
rect 715 -770 725 -750
rect 745 -770 755 -750
rect 715 -785 755 -770
rect 770 -550 810 -535
rect 770 -570 780 -550
rect 800 -570 810 -550
rect 770 -600 810 -570
rect 770 -620 780 -600
rect 800 -620 810 -600
rect 770 -650 810 -620
rect 770 -670 780 -650
rect 800 -670 810 -650
rect 770 -700 810 -670
rect 770 -720 780 -700
rect 800 -720 810 -700
rect 770 -750 810 -720
rect 770 -770 780 -750
rect 800 -770 810 -750
rect 770 -785 810 -770
rect 825 -550 865 -535
rect 825 -570 835 -550
rect 855 -570 865 -550
rect 825 -600 865 -570
rect 825 -620 835 -600
rect 855 -620 865 -600
rect 825 -650 865 -620
rect 825 -670 835 -650
rect 855 -670 865 -650
rect 825 -700 865 -670
rect 825 -720 835 -700
rect 855 -720 865 -700
rect 825 -750 865 -720
rect 825 -770 835 -750
rect 855 -770 865 -750
rect 825 -785 865 -770
rect 880 -550 920 -535
rect 880 -570 890 -550
rect 910 -570 920 -550
rect 880 -600 920 -570
rect 880 -620 890 -600
rect 910 -620 920 -600
rect 880 -650 920 -620
rect 880 -670 890 -650
rect 910 -670 920 -650
rect 880 -700 920 -670
rect 880 -720 890 -700
rect 910 -720 920 -700
rect 880 -750 920 -720
rect 880 -770 890 -750
rect 910 -770 920 -750
rect 880 -785 920 -770
rect 935 -550 975 -535
rect 935 -570 945 -550
rect 965 -570 975 -550
rect 935 -600 975 -570
rect 935 -620 945 -600
rect 965 -620 975 -600
rect 935 -650 975 -620
rect 935 -670 945 -650
rect 965 -670 975 -650
rect 935 -700 975 -670
rect 935 -720 945 -700
rect 965 -720 975 -700
rect 935 -750 975 -720
rect 935 -770 945 -750
rect 965 -770 975 -750
rect 935 -785 975 -770
rect 990 -550 1030 -535
rect 990 -570 1000 -550
rect 1020 -570 1030 -550
rect 990 -600 1030 -570
rect 990 -620 1000 -600
rect 1020 -620 1030 -600
rect 990 -650 1030 -620
rect 990 -670 1000 -650
rect 1020 -670 1030 -650
rect 990 -700 1030 -670
rect 990 -720 1000 -700
rect 1020 -720 1030 -700
rect 990 -750 1030 -720
rect 990 -770 1000 -750
rect 1020 -770 1030 -750
rect 990 -785 1030 -770
rect 1045 -550 1085 -535
rect 1045 -570 1055 -550
rect 1075 -570 1085 -550
rect 1045 -600 1085 -570
rect 1045 -620 1055 -600
rect 1075 -620 1085 -600
rect 1045 -650 1085 -620
rect 1045 -670 1055 -650
rect 1075 -670 1085 -650
rect 1045 -700 1085 -670
rect 1045 -720 1055 -700
rect 1075 -720 1085 -700
rect 1045 -750 1085 -720
rect 1045 -770 1055 -750
rect 1075 -770 1085 -750
rect 1045 -785 1085 -770
rect 1100 -550 1140 -535
rect 1100 -570 1110 -550
rect 1130 -570 1140 -550
rect 1100 -600 1140 -570
rect 1100 -620 1110 -600
rect 1130 -620 1140 -600
rect 1100 -650 1140 -620
rect 1100 -670 1110 -650
rect 1130 -670 1140 -650
rect 1100 -700 1140 -670
rect 1100 -720 1110 -700
rect 1130 -720 1140 -700
rect 1100 -750 1140 -720
rect 1100 -770 1110 -750
rect 1130 -770 1140 -750
rect 1100 -785 1140 -770
rect 1155 -550 1195 -535
rect 1155 -570 1165 -550
rect 1185 -570 1195 -550
rect 1155 -600 1195 -570
rect 1155 -620 1165 -600
rect 1185 -620 1195 -600
rect 1155 -650 1195 -620
rect 1155 -670 1165 -650
rect 1185 -670 1195 -650
rect 1155 -700 1195 -670
rect 1155 -720 1165 -700
rect 1185 -720 1195 -700
rect 1155 -750 1195 -720
rect 1155 -770 1165 -750
rect 1185 -770 1195 -750
rect 1155 -785 1195 -770
rect 1210 -550 1250 -535
rect 1210 -570 1220 -550
rect 1240 -570 1250 -550
rect 1210 -600 1250 -570
rect 1210 -620 1220 -600
rect 1240 -620 1250 -600
rect 1210 -650 1250 -620
rect 1210 -670 1220 -650
rect 1240 -670 1250 -650
rect 1210 -700 1250 -670
rect 1210 -720 1220 -700
rect 1240 -720 1250 -700
rect 1210 -750 1250 -720
rect 1210 -770 1220 -750
rect 1240 -770 1250 -750
rect 1210 -785 1250 -770
rect 1265 -550 1305 -535
rect 1265 -570 1275 -550
rect 1295 -570 1305 -550
rect 1265 -600 1305 -570
rect 1265 -620 1275 -600
rect 1295 -620 1305 -600
rect 1265 -650 1305 -620
rect 1265 -670 1275 -650
rect 1295 -670 1305 -650
rect 1265 -700 1305 -670
rect 1265 -720 1275 -700
rect 1295 -720 1305 -700
rect 1265 -750 1305 -720
rect 1265 -770 1275 -750
rect 1295 -770 1305 -750
rect 1265 -785 1305 -770
rect 1320 -550 1360 -535
rect 1320 -570 1330 -550
rect 1350 -570 1360 -550
rect 1320 -600 1360 -570
rect 1320 -620 1330 -600
rect 1350 -620 1360 -600
rect 1320 -650 1360 -620
rect 1320 -670 1330 -650
rect 1350 -670 1360 -650
rect 1320 -700 1360 -670
rect 1320 -720 1330 -700
rect 1350 -720 1360 -700
rect 1320 -750 1360 -720
rect 1320 -770 1330 -750
rect 1350 -770 1360 -750
rect 1320 -785 1360 -770
rect 1375 -550 1415 -535
rect 1375 -570 1385 -550
rect 1405 -570 1415 -550
rect 1375 -600 1415 -570
rect 1375 -620 1385 -600
rect 1405 -620 1415 -600
rect 1375 -650 1415 -620
rect 1375 -670 1385 -650
rect 1405 -670 1415 -650
rect 1375 -700 1415 -670
rect 1375 -720 1385 -700
rect 1405 -720 1415 -700
rect 1375 -750 1415 -720
rect 1375 -770 1385 -750
rect 1405 -770 1415 -750
rect 1375 -785 1415 -770
rect 1430 -550 1470 -535
rect 1430 -570 1440 -550
rect 1460 -570 1470 -550
rect 1430 -600 1470 -570
rect 1430 -620 1440 -600
rect 1460 -620 1470 -600
rect 1430 -650 1470 -620
rect 1430 -670 1440 -650
rect 1460 -670 1470 -650
rect 1430 -700 1470 -670
rect 1430 -720 1440 -700
rect 1460 -720 1470 -700
rect 1430 -750 1470 -720
rect 1430 -770 1440 -750
rect 1460 -770 1470 -750
rect 1430 -785 1470 -770
rect 2075 -540 2085 -520
rect 2105 -540 2115 -520
rect 2075 -570 2115 -540
rect 2075 -590 2085 -570
rect 2105 -590 2115 -570
rect 2075 -620 2115 -590
rect 2075 -640 2085 -620
rect 2105 -640 2115 -620
rect 2075 -670 2115 -640
rect 2075 -690 2085 -670
rect 2105 -690 2115 -670
rect 2075 -720 2115 -690
rect 2075 -740 2085 -720
rect 2105 -740 2115 -720
rect 2075 -770 2115 -740
rect -425 -820 -385 -790
rect 2075 -790 2085 -770
rect 2105 -790 2115 -770
rect -425 -840 -415 -820
rect -395 -840 -385 -820
rect 2075 -820 2115 -790
rect 2075 -840 2085 -820
rect 2105 -840 2115 -820
rect -425 -870 -385 -840
rect -425 -890 -415 -870
rect -395 -890 -385 -870
rect -425 -920 -385 -890
rect 2075 -870 2115 -840
rect 2075 -890 2085 -870
rect 2105 -890 2115 -870
rect -425 -940 -415 -920
rect -395 -940 -385 -920
rect -425 -970 -385 -940
rect 2075 -920 2115 -890
rect 2075 -940 2085 -920
rect 2105 -940 2115 -920
rect -425 -990 -415 -970
rect -395 -990 -385 -970
rect -425 -1020 -385 -990
rect -425 -1040 -415 -1020
rect -395 -1040 -385 -1020
rect -425 -1055 -385 -1040
rect 495 -965 535 -950
rect 495 -985 505 -965
rect 525 -985 535 -965
rect 495 -1015 535 -985
rect 495 -1035 505 -1015
rect 525 -1035 535 -1015
rect 495 -1065 535 -1035
rect 495 -1085 505 -1065
rect 525 -1085 535 -1065
rect 495 -1100 535 -1085
rect 550 -965 590 -950
rect 550 -985 560 -965
rect 580 -985 590 -965
rect 550 -1015 590 -985
rect 550 -1035 560 -1015
rect 580 -1035 590 -1015
rect 550 -1065 590 -1035
rect 550 -1085 560 -1065
rect 580 -1085 590 -1065
rect 550 -1100 590 -1085
rect 605 -965 645 -950
rect 605 -985 615 -965
rect 635 -985 645 -965
rect 605 -1015 645 -985
rect 605 -1035 615 -1015
rect 635 -1035 645 -1015
rect 605 -1065 645 -1035
rect 605 -1085 615 -1065
rect 635 -1085 645 -1065
rect 605 -1100 645 -1085
rect 660 -965 700 -950
rect 660 -985 670 -965
rect 690 -985 700 -965
rect 660 -1015 700 -985
rect 660 -1035 670 -1015
rect 690 -1035 700 -1015
rect 660 -1065 700 -1035
rect 660 -1085 670 -1065
rect 690 -1085 700 -1065
rect 660 -1100 700 -1085
rect 715 -965 755 -950
rect 715 -985 725 -965
rect 745 -985 755 -965
rect 715 -1015 755 -985
rect 715 -1035 725 -1015
rect 745 -1035 755 -1015
rect 715 -1065 755 -1035
rect 715 -1085 725 -1065
rect 745 -1085 755 -1065
rect 715 -1100 755 -1085
rect 770 -965 810 -950
rect 770 -985 780 -965
rect 800 -985 810 -965
rect 770 -1015 810 -985
rect 770 -1035 780 -1015
rect 800 -1035 810 -1015
rect 770 -1065 810 -1035
rect 770 -1085 780 -1065
rect 800 -1085 810 -1065
rect 770 -1100 810 -1085
rect 825 -965 865 -950
rect 825 -985 835 -965
rect 855 -985 865 -965
rect 825 -1015 865 -985
rect 825 -1035 835 -1015
rect 855 -1035 865 -1015
rect 825 -1065 865 -1035
rect 825 -1085 835 -1065
rect 855 -1085 865 -1065
rect 825 -1100 865 -1085
rect 960 -965 1000 -950
rect 960 -985 970 -965
rect 990 -985 1000 -965
rect 960 -1015 1000 -985
rect 960 -1035 970 -1015
rect 990 -1035 1000 -1015
rect 960 -1065 1000 -1035
rect 960 -1085 970 -1065
rect 990 -1085 1000 -1065
rect 960 -1100 1000 -1085
rect 1300 -965 1340 -950
rect 1300 -985 1310 -965
rect 1330 -985 1340 -965
rect 1300 -1015 1340 -985
rect 1300 -1035 1310 -1015
rect 1330 -1035 1340 -1015
rect 1300 -1065 1340 -1035
rect 2075 -970 2115 -940
rect 2075 -990 2085 -970
rect 2105 -990 2115 -970
rect 2075 -1020 2115 -990
rect 2075 -1040 2085 -1020
rect 2105 -1040 2115 -1020
rect 2075 -1055 2115 -1040
rect 2175 -370 2215 -355
rect 2175 -390 2185 -370
rect 2205 -390 2215 -370
rect 2175 -420 2215 -390
rect 2175 -440 2185 -420
rect 2205 -440 2215 -420
rect 2175 -470 2215 -440
rect 2175 -490 2185 -470
rect 2205 -490 2215 -470
rect 2175 -520 2215 -490
rect 2175 -540 2185 -520
rect 2205 -540 2215 -520
rect 2175 -570 2215 -540
rect 2175 -590 2185 -570
rect 2205 -590 2215 -570
rect 2175 -620 2215 -590
rect 2175 -640 2185 -620
rect 2205 -640 2215 -620
rect 2175 -670 2215 -640
rect 2175 -690 2185 -670
rect 2205 -690 2215 -670
rect 2175 -720 2215 -690
rect 2175 -740 2185 -720
rect 2205 -740 2215 -720
rect 2175 -770 2215 -740
rect 2175 -790 2185 -770
rect 2205 -790 2215 -770
rect 2175 -820 2215 -790
rect 2175 -840 2185 -820
rect 2205 -840 2215 -820
rect 2175 -870 2215 -840
rect 2175 -890 2185 -870
rect 2205 -890 2215 -870
rect 2175 -920 2215 -890
rect 2175 -940 2185 -920
rect 2205 -940 2215 -920
rect 2175 -970 2215 -940
rect 2175 -990 2185 -970
rect 2205 -990 2215 -970
rect 2175 -1020 2215 -990
rect 2175 -1040 2185 -1020
rect 2205 -1040 2215 -1020
rect 2175 -1055 2215 -1040
rect 2275 -370 2315 -355
rect 2275 -390 2285 -370
rect 2305 -390 2315 -370
rect 2275 -420 2315 -390
rect 2275 -440 2285 -420
rect 2305 -440 2315 -420
rect 2275 -470 2315 -440
rect 2275 -490 2285 -470
rect 2305 -490 2315 -470
rect 2275 -520 2315 -490
rect 2275 -540 2285 -520
rect 2305 -540 2315 -520
rect 2275 -570 2315 -540
rect 2275 -590 2285 -570
rect 2305 -590 2315 -570
rect 2275 -620 2315 -590
rect 2275 -640 2285 -620
rect 2305 -640 2315 -620
rect 2275 -670 2315 -640
rect 2275 -690 2285 -670
rect 2305 -690 2315 -670
rect 2275 -720 2315 -690
rect 2275 -740 2285 -720
rect 2305 -740 2315 -720
rect 2275 -770 2315 -740
rect 2275 -790 2285 -770
rect 2305 -790 2315 -770
rect 2275 -820 2315 -790
rect 2275 -840 2285 -820
rect 2305 -840 2315 -820
rect 2275 -870 2315 -840
rect 2275 -890 2285 -870
rect 2305 -890 2315 -870
rect 2275 -920 2315 -890
rect 2275 -940 2285 -920
rect 2305 -940 2315 -920
rect 2275 -970 2315 -940
rect 2275 -990 2285 -970
rect 2305 -990 2315 -970
rect 2275 -1020 2315 -990
rect 2275 -1040 2285 -1020
rect 2305 -1040 2315 -1020
rect 2275 -1055 2315 -1040
rect 2375 -370 2415 -355
rect 2375 -390 2385 -370
rect 2405 -390 2415 -370
rect 2375 -420 2415 -390
rect 2375 -440 2385 -420
rect 2405 -440 2415 -420
rect 2375 -470 2415 -440
rect 2375 -490 2385 -470
rect 2405 -490 2415 -470
rect 2375 -520 2415 -490
rect 2375 -540 2385 -520
rect 2405 -540 2415 -520
rect 2375 -570 2415 -540
rect 2375 -590 2385 -570
rect 2405 -590 2415 -570
rect 2375 -620 2415 -590
rect 2375 -640 2385 -620
rect 2405 -640 2415 -620
rect 2375 -670 2415 -640
rect 2375 -690 2385 -670
rect 2405 -690 2415 -670
rect 2375 -720 2415 -690
rect 2375 -740 2385 -720
rect 2405 -740 2415 -720
rect 2375 -770 2415 -740
rect 2375 -790 2385 -770
rect 2405 -790 2415 -770
rect 2375 -820 2415 -790
rect 2375 -840 2385 -820
rect 2405 -840 2415 -820
rect 2375 -870 2415 -840
rect 2375 -890 2385 -870
rect 2405 -890 2415 -870
rect 2375 -920 2415 -890
rect 2375 -940 2385 -920
rect 2405 -940 2415 -920
rect 2375 -970 2415 -940
rect 2375 -990 2385 -970
rect 2405 -990 2415 -970
rect 2375 -1020 2415 -990
rect 2375 -1040 2385 -1020
rect 2405 -1040 2415 -1020
rect 2375 -1055 2415 -1040
rect 2475 -370 2515 -355
rect 2475 -390 2485 -370
rect 2505 -390 2515 -370
rect 2475 -420 2515 -390
rect 2475 -440 2485 -420
rect 2505 -440 2515 -420
rect 2475 -470 2515 -440
rect 2475 -490 2485 -470
rect 2505 -490 2515 -470
rect 2475 -520 2515 -490
rect 2475 -540 2485 -520
rect 2505 -540 2515 -520
rect 2475 -570 2515 -540
rect 2475 -590 2485 -570
rect 2505 -590 2515 -570
rect 2475 -620 2515 -590
rect 2475 -640 2485 -620
rect 2505 -640 2515 -620
rect 2475 -670 2515 -640
rect 2475 -690 2485 -670
rect 2505 -690 2515 -670
rect 2475 -720 2515 -690
rect 2475 -740 2485 -720
rect 2505 -740 2515 -720
rect 2475 -770 2515 -740
rect 2475 -790 2485 -770
rect 2505 -790 2515 -770
rect 2475 -820 2515 -790
rect 2475 -840 2485 -820
rect 2505 -840 2515 -820
rect 2475 -870 2515 -840
rect 2475 -890 2485 -870
rect 2505 -890 2515 -870
rect 2475 -920 2515 -890
rect 2475 -940 2485 -920
rect 2505 -940 2515 -920
rect 2475 -970 2515 -940
rect 2475 -990 2485 -970
rect 2505 -990 2515 -970
rect 2475 -1020 2515 -990
rect 2475 -1040 2485 -1020
rect 2505 -1040 2515 -1020
rect 2475 -1055 2515 -1040
rect 2575 -370 2615 -355
rect 2575 -390 2585 -370
rect 2605 -390 2615 -370
rect 2575 -420 2615 -390
rect 2575 -440 2585 -420
rect 2605 -440 2615 -420
rect 2575 -470 2615 -440
rect 2575 -490 2585 -470
rect 2605 -490 2615 -470
rect 2575 -520 2615 -490
rect 2575 -540 2585 -520
rect 2605 -540 2615 -520
rect 2575 -570 2615 -540
rect 2575 -590 2585 -570
rect 2605 -590 2615 -570
rect 2575 -620 2615 -590
rect 2575 -640 2585 -620
rect 2605 -640 2615 -620
rect 2575 -670 2615 -640
rect 2575 -690 2585 -670
rect 2605 -690 2615 -670
rect 2575 -720 2615 -690
rect 2575 -740 2585 -720
rect 2605 -740 2615 -720
rect 2575 -770 2615 -740
rect 2575 -790 2585 -770
rect 2605 -790 2615 -770
rect 2575 -820 2615 -790
rect 2575 -840 2585 -820
rect 2605 -840 2615 -820
rect 2575 -870 2615 -840
rect 2575 -890 2585 -870
rect 2605 -890 2615 -870
rect 2575 -920 2615 -890
rect 2575 -940 2585 -920
rect 2605 -940 2615 -920
rect 2575 -970 2615 -940
rect 2575 -990 2585 -970
rect 2605 -990 2615 -970
rect 2575 -1020 2615 -990
rect 2575 -1040 2585 -1020
rect 2605 -1040 2615 -1020
rect 2575 -1055 2615 -1040
rect 2675 -370 2715 -355
rect 2675 -390 2685 -370
rect 2705 -390 2715 -370
rect 2675 -420 2715 -390
rect 2675 -440 2685 -420
rect 2705 -440 2715 -420
rect 2675 -470 2715 -440
rect 2675 -490 2685 -470
rect 2705 -490 2715 -470
rect 2675 -520 2715 -490
rect 2675 -540 2685 -520
rect 2705 -540 2715 -520
rect 2675 -570 2715 -540
rect 2675 -590 2685 -570
rect 2705 -590 2715 -570
rect 2675 -620 2715 -590
rect 2675 -640 2685 -620
rect 2705 -640 2715 -620
rect 2675 -670 2715 -640
rect 2675 -690 2685 -670
rect 2705 -690 2715 -670
rect 2675 -720 2715 -690
rect 2675 -740 2685 -720
rect 2705 -740 2715 -720
rect 2675 -770 2715 -740
rect 2675 -790 2685 -770
rect 2705 -790 2715 -770
rect 2675 -820 2715 -790
rect 2675 -840 2685 -820
rect 2705 -840 2715 -820
rect 2675 -870 2715 -840
rect 2675 -890 2685 -870
rect 2705 -890 2715 -870
rect 2675 -920 2715 -890
rect 2675 -940 2685 -920
rect 2705 -940 2715 -920
rect 2675 -970 2715 -940
rect 2675 -990 2685 -970
rect 2705 -990 2715 -970
rect 2675 -1020 2715 -990
rect 2675 -1040 2685 -1020
rect 2705 -1040 2715 -1020
rect 2675 -1055 2715 -1040
rect 1300 -1085 1310 -1065
rect 1330 -1085 1340 -1065
rect 1300 -1100 1340 -1085
<< pdiff >>
rect 30 2660 70 2675
rect 30 2640 40 2660
rect 60 2640 70 2660
rect 30 2610 70 2640
rect 30 2590 40 2610
rect 60 2590 70 2610
rect 30 2560 70 2590
rect 30 2540 40 2560
rect 60 2540 70 2560
rect 30 2510 70 2540
rect 30 2490 40 2510
rect 60 2490 70 2510
rect 30 2460 70 2490
rect 30 2440 40 2460
rect 60 2440 70 2460
rect 30 2410 70 2440
rect 30 2390 40 2410
rect 60 2390 70 2410
rect 30 2360 70 2390
rect 30 2340 40 2360
rect 60 2340 70 2360
rect 30 2325 70 2340
rect 90 2660 130 2675
rect 90 2640 100 2660
rect 120 2640 130 2660
rect 90 2610 130 2640
rect 90 2590 100 2610
rect 120 2590 130 2610
rect 90 2560 130 2590
rect 90 2540 100 2560
rect 120 2540 130 2560
rect 90 2510 130 2540
rect 90 2490 100 2510
rect 120 2490 130 2510
rect 90 2460 130 2490
rect 90 2440 100 2460
rect 120 2440 130 2460
rect 90 2410 130 2440
rect 90 2390 100 2410
rect 120 2390 130 2410
rect 90 2360 130 2390
rect 90 2340 100 2360
rect 120 2340 130 2360
rect 90 2325 130 2340
rect 150 2660 190 2675
rect 150 2640 160 2660
rect 180 2640 190 2660
rect 150 2610 190 2640
rect 150 2590 160 2610
rect 180 2590 190 2610
rect 150 2560 190 2590
rect 150 2540 160 2560
rect 180 2540 190 2560
rect 150 2510 190 2540
rect 150 2490 160 2510
rect 180 2490 190 2510
rect 150 2460 190 2490
rect 150 2440 160 2460
rect 180 2440 190 2460
rect 150 2410 190 2440
rect 150 2390 160 2410
rect 180 2390 190 2410
rect 150 2360 190 2390
rect 150 2340 160 2360
rect 180 2340 190 2360
rect 150 2325 190 2340
rect 210 2660 250 2675
rect 210 2640 220 2660
rect 240 2640 250 2660
rect 210 2610 250 2640
rect 210 2590 220 2610
rect 240 2590 250 2610
rect 210 2560 250 2590
rect 970 2660 1010 2675
rect 970 2640 980 2660
rect 1000 2640 1010 2660
rect 970 2610 1010 2640
rect 970 2590 980 2610
rect 1000 2590 1010 2610
rect 970 2560 1010 2590
rect 210 2540 220 2560
rect 240 2540 250 2560
rect 210 2510 250 2540
rect 970 2540 980 2560
rect 1000 2540 1010 2560
rect 210 2490 220 2510
rect 240 2490 250 2510
rect 970 2510 1010 2540
rect 210 2460 250 2490
rect 210 2440 220 2460
rect 240 2440 250 2460
rect 210 2410 250 2440
rect 210 2390 220 2410
rect 240 2390 250 2410
rect 210 2360 250 2390
rect 210 2340 220 2360
rect 240 2340 250 2360
rect 210 2325 250 2340
rect 500 2360 540 2505
rect 500 2340 510 2360
rect 530 2340 540 2360
rect 500 2325 540 2340
rect 560 2360 600 2505
rect 560 2340 570 2360
rect 590 2340 600 2360
rect 560 2325 600 2340
rect 620 2360 660 2505
rect 620 2340 630 2360
rect 650 2340 660 2360
rect 620 2325 660 2340
rect 680 2360 720 2505
rect 680 2340 690 2360
rect 710 2340 720 2360
rect 680 2325 720 2340
rect 970 2490 980 2510
rect 1000 2490 1010 2510
rect 970 2460 1010 2490
rect 970 2440 980 2460
rect 1000 2440 1010 2460
rect 970 2410 1010 2440
rect 970 2390 980 2410
rect 1000 2390 1010 2410
rect 970 2360 1010 2390
rect 970 2340 980 2360
rect 1000 2340 1010 2360
rect 970 2325 1010 2340
rect 1030 2660 1070 2675
rect 1030 2640 1040 2660
rect 1060 2640 1070 2660
rect 1030 2610 1070 2640
rect 1030 2590 1040 2610
rect 1060 2590 1070 2610
rect 1030 2560 1070 2590
rect 1030 2540 1040 2560
rect 1060 2540 1070 2560
rect 1030 2510 1070 2540
rect 1030 2490 1040 2510
rect 1060 2490 1070 2510
rect 1030 2460 1070 2490
rect 1030 2440 1040 2460
rect 1060 2440 1070 2460
rect 1030 2410 1070 2440
rect 1030 2390 1040 2410
rect 1060 2390 1070 2410
rect 1030 2360 1070 2390
rect 1030 2340 1040 2360
rect 1060 2340 1070 2360
rect 1030 2325 1070 2340
rect 1090 2660 1130 2675
rect 1090 2640 1100 2660
rect 1120 2640 1130 2660
rect 1090 2610 1130 2640
rect 1090 2590 1100 2610
rect 1120 2590 1130 2610
rect 1090 2560 1130 2590
rect 1090 2540 1100 2560
rect 1120 2540 1130 2560
rect 1090 2510 1130 2540
rect 1090 2490 1100 2510
rect 1120 2490 1130 2510
rect 1090 2460 1130 2490
rect 1090 2440 1100 2460
rect 1120 2440 1130 2460
rect 1090 2410 1130 2440
rect 1090 2390 1100 2410
rect 1120 2390 1130 2410
rect 1090 2360 1130 2390
rect 1090 2340 1100 2360
rect 1120 2340 1130 2360
rect 1090 2325 1130 2340
rect 1150 2660 1190 2675
rect 1150 2640 1160 2660
rect 1180 2640 1190 2660
rect 1150 2610 1190 2640
rect 1150 2590 1160 2610
rect 1180 2590 1190 2610
rect 1150 2560 1190 2590
rect 1150 2540 1160 2560
rect 1180 2540 1190 2560
rect 1150 2510 1190 2540
rect 1150 2490 1160 2510
rect 1180 2490 1190 2510
rect 1150 2460 1190 2490
rect 1150 2440 1160 2460
rect 1180 2440 1190 2460
rect 1150 2410 1190 2440
rect 1150 2390 1160 2410
rect 1180 2390 1190 2410
rect 1150 2360 1190 2390
rect 1150 2340 1160 2360
rect 1180 2340 1190 2360
rect 1150 2325 1190 2340
rect 1438 2660 1478 2675
rect 1438 2640 1448 2660
rect 1468 2640 1478 2660
rect 1438 2610 1478 2640
rect 1438 2590 1448 2610
rect 1468 2590 1478 2610
rect 1438 2560 1478 2590
rect 1438 2540 1448 2560
rect 1468 2540 1478 2560
rect 1438 2510 1478 2540
rect 1438 2490 1448 2510
rect 1468 2490 1478 2510
rect 1438 2460 1478 2490
rect 1438 2440 1448 2460
rect 1468 2440 1478 2460
rect 1438 2410 1478 2440
rect 1438 2390 1448 2410
rect 1468 2390 1478 2410
rect 1438 2360 1478 2390
rect 1438 2340 1448 2360
rect 1468 2340 1478 2360
rect 1438 2325 1478 2340
rect 1498 2660 1538 2675
rect 1498 2640 1508 2660
rect 1528 2640 1538 2660
rect 1498 2610 1538 2640
rect 1498 2590 1508 2610
rect 1528 2590 1538 2610
rect 1498 2560 1538 2590
rect 1498 2540 1508 2560
rect 1528 2540 1538 2560
rect 1498 2510 1538 2540
rect 1498 2490 1508 2510
rect 1528 2490 1538 2510
rect 1498 2460 1538 2490
rect 1498 2440 1508 2460
rect 1528 2440 1538 2460
rect 1498 2410 1538 2440
rect 1498 2390 1508 2410
rect 1528 2390 1538 2410
rect 1498 2360 1538 2390
rect 1498 2340 1508 2360
rect 1528 2340 1538 2360
rect 1498 2325 1538 2340
rect 1558 2660 1598 2675
rect 1558 2640 1568 2660
rect 1588 2640 1598 2660
rect 1558 2610 1598 2640
rect 1558 2590 1568 2610
rect 1588 2590 1598 2610
rect 1558 2560 1598 2590
rect 1558 2540 1568 2560
rect 1588 2540 1598 2560
rect 1558 2510 1598 2540
rect 1558 2490 1568 2510
rect 1588 2490 1598 2510
rect 1558 2460 1598 2490
rect 1558 2440 1568 2460
rect 1588 2440 1598 2460
rect 1558 2410 1598 2440
rect 1558 2390 1568 2410
rect 1588 2390 1598 2410
rect 1558 2360 1598 2390
rect 1558 2340 1568 2360
rect 1588 2340 1598 2360
rect 1558 2325 1598 2340
rect 1618 2660 1658 2675
rect 1618 2640 1628 2660
rect 1648 2640 1658 2660
rect 1618 2610 1658 2640
rect 1618 2590 1628 2610
rect 1648 2590 1658 2610
rect 1618 2560 1658 2590
rect 1618 2540 1628 2560
rect 1648 2540 1658 2560
rect 1618 2510 1658 2540
rect 1618 2490 1628 2510
rect 1648 2490 1658 2510
rect 1618 2460 1658 2490
rect 1618 2440 1628 2460
rect 1648 2440 1658 2460
rect 1618 2410 1658 2440
rect 1618 2390 1628 2410
rect 1648 2390 1658 2410
rect 1618 2360 1658 2390
rect 1618 2340 1628 2360
rect 1648 2340 1658 2360
rect 1618 2325 1658 2340
rect -1165 2085 -1125 2100
rect -1165 2065 -1155 2085
rect -1135 2065 -1125 2085
rect -1165 2035 -1125 2065
rect -1165 2015 -1155 2035
rect -1135 2015 -1125 2035
rect -1165 1985 -1125 2015
rect -1165 1965 -1155 1985
rect -1135 1965 -1125 1985
rect -1165 1935 -1125 1965
rect -1165 1915 -1155 1935
rect -1135 1915 -1125 1935
rect -1165 1885 -1125 1915
rect -1165 1865 -1155 1885
rect -1135 1865 -1125 1885
rect -1165 1835 -1125 1865
rect -1165 1815 -1155 1835
rect -1135 1815 -1125 1835
rect -1165 1785 -1125 1815
rect -1165 1765 -1155 1785
rect -1135 1765 -1125 1785
rect -1165 1750 -1125 1765
rect -1105 2085 -1065 2100
rect -1105 2065 -1095 2085
rect -1075 2065 -1065 2085
rect -1105 2035 -1065 2065
rect -1105 2015 -1095 2035
rect -1075 2015 -1065 2035
rect -1105 1985 -1065 2015
rect -1105 1965 -1095 1985
rect -1075 1965 -1065 1985
rect -1105 1935 -1065 1965
rect -1105 1915 -1095 1935
rect -1075 1915 -1065 1935
rect -1105 1885 -1065 1915
rect -1105 1865 -1095 1885
rect -1075 1865 -1065 1885
rect -1105 1835 -1065 1865
rect -1105 1815 -1095 1835
rect -1075 1815 -1065 1835
rect -1105 1785 -1065 1815
rect -1105 1765 -1095 1785
rect -1075 1765 -1065 1785
rect -1105 1750 -1065 1765
rect -1045 2085 -1005 2100
rect -1045 2065 -1035 2085
rect -1015 2065 -1005 2085
rect -1045 2035 -1005 2065
rect -1045 2015 -1035 2035
rect -1015 2015 -1005 2035
rect -1045 1985 -1005 2015
rect -1045 1965 -1035 1985
rect -1015 1965 -1005 1985
rect -1045 1935 -1005 1965
rect -1045 1915 -1035 1935
rect -1015 1915 -1005 1935
rect -1045 1885 -1005 1915
rect -1045 1865 -1035 1885
rect -1015 1865 -1005 1885
rect -1045 1835 -1005 1865
rect -1045 1815 -1035 1835
rect -1015 1815 -1005 1835
rect -1045 1785 -1005 1815
rect -1045 1765 -1035 1785
rect -1015 1765 -1005 1785
rect -1045 1750 -1005 1765
rect -985 2085 -945 2100
rect -985 2065 -975 2085
rect -955 2065 -945 2085
rect -985 2035 -945 2065
rect -985 2015 -975 2035
rect -955 2015 -945 2035
rect -985 1985 -945 2015
rect -985 1965 -975 1985
rect -955 1965 -945 1985
rect -985 1935 -945 1965
rect -985 1915 -975 1935
rect -955 1915 -945 1935
rect -985 1885 -945 1915
rect -985 1865 -975 1885
rect -955 1865 -945 1885
rect -985 1835 -945 1865
rect -985 1815 -975 1835
rect -955 1815 -945 1835
rect -985 1785 -945 1815
rect -985 1765 -975 1785
rect -955 1765 -945 1785
rect -985 1750 -945 1765
rect -925 2085 -885 2100
rect -925 2065 -915 2085
rect -895 2065 -885 2085
rect -925 2035 -885 2065
rect -925 2015 -915 2035
rect -895 2015 -885 2035
rect -925 1985 -885 2015
rect -925 1965 -915 1985
rect -895 1965 -885 1985
rect -925 1935 -885 1965
rect -925 1915 -915 1935
rect -895 1915 -885 1935
rect -925 1885 -885 1915
rect -925 1865 -915 1885
rect -895 1865 -885 1885
rect -925 1835 -885 1865
rect -925 1815 -915 1835
rect -895 1815 -885 1835
rect -925 1785 -885 1815
rect -925 1765 -915 1785
rect -895 1765 -885 1785
rect -925 1750 -885 1765
rect -865 2085 -825 2100
rect -865 2065 -855 2085
rect -835 2065 -825 2085
rect -865 2035 -825 2065
rect -865 2015 -855 2035
rect -835 2015 -825 2035
rect -865 1985 -825 2015
rect -865 1965 -855 1985
rect -835 1965 -825 1985
rect -865 1935 -825 1965
rect -865 1915 -855 1935
rect -835 1915 -825 1935
rect -865 1885 -825 1915
rect -865 1865 -855 1885
rect -835 1865 -825 1885
rect -865 1835 -825 1865
rect -865 1815 -855 1835
rect -835 1815 -825 1835
rect -865 1785 -825 1815
rect -865 1765 -855 1785
rect -835 1765 -825 1785
rect -865 1750 -825 1765
rect -805 2085 -765 2100
rect -805 2065 -795 2085
rect -775 2065 -765 2085
rect -805 2035 -765 2065
rect -805 2015 -795 2035
rect -775 2015 -765 2035
rect -805 1985 -765 2015
rect -805 1965 -795 1985
rect -775 1965 -765 1985
rect -805 1935 -765 1965
rect -805 1915 -795 1935
rect -775 1915 -765 1935
rect -805 1885 -765 1915
rect -805 1865 -795 1885
rect -775 1865 -765 1885
rect -805 1835 -765 1865
rect -805 1815 -795 1835
rect -775 1815 -765 1835
rect -805 1785 -765 1815
rect -805 1765 -795 1785
rect -775 1765 -765 1785
rect -805 1750 -765 1765
rect -745 2085 -705 2100
rect -745 2065 -735 2085
rect -715 2065 -705 2085
rect -745 2035 -705 2065
rect -745 2015 -735 2035
rect -715 2015 -705 2035
rect -745 1985 -705 2015
rect -745 1965 -735 1985
rect -715 1965 -705 1985
rect -745 1935 -705 1965
rect -745 1915 -735 1935
rect -715 1915 -705 1935
rect -745 1885 -705 1915
rect -745 1865 -735 1885
rect -715 1865 -705 1885
rect -745 1835 -705 1865
rect -745 1815 -735 1835
rect -715 1815 -705 1835
rect -745 1785 -705 1815
rect -745 1765 -735 1785
rect -715 1765 -705 1785
rect -745 1750 -705 1765
rect -685 2085 -645 2100
rect -685 2065 -675 2085
rect -655 2065 -645 2085
rect -685 2035 -645 2065
rect -685 2015 -675 2035
rect -655 2015 -645 2035
rect -685 1985 -645 2015
rect -685 1965 -675 1985
rect -655 1965 -645 1985
rect -685 1935 -645 1965
rect -685 1915 -675 1935
rect -655 1915 -645 1935
rect -685 1885 -645 1915
rect -685 1865 -675 1885
rect -655 1865 -645 1885
rect -685 1835 -645 1865
rect -685 1815 -675 1835
rect -655 1815 -645 1835
rect -685 1785 -645 1815
rect -685 1765 -675 1785
rect -655 1765 -645 1785
rect -685 1750 -645 1765
rect -625 2085 -585 2100
rect -625 2065 -615 2085
rect -595 2065 -585 2085
rect -625 2035 -585 2065
rect -625 2015 -615 2035
rect -595 2015 -585 2035
rect -625 1985 -585 2015
rect -625 1965 -615 1985
rect -595 1965 -585 1985
rect -625 1935 -585 1965
rect -625 1915 -615 1935
rect -595 1915 -585 1935
rect -625 1885 -585 1915
rect -625 1865 -615 1885
rect -595 1865 -585 1885
rect -625 1835 -585 1865
rect -625 1815 -615 1835
rect -595 1815 -585 1835
rect -625 1785 -585 1815
rect -625 1765 -615 1785
rect -595 1765 -585 1785
rect -625 1750 -585 1765
rect -565 2085 -525 2100
rect -565 2065 -555 2085
rect -535 2065 -525 2085
rect -565 2035 -525 2065
rect -565 2015 -555 2035
rect -535 2015 -525 2035
rect -565 1985 -525 2015
rect -565 1965 -555 1985
rect -535 1965 -525 1985
rect -565 1935 -525 1965
rect -565 1915 -555 1935
rect -535 1915 -525 1935
rect -565 1885 -525 1915
rect -565 1865 -555 1885
rect -535 1865 -525 1885
rect -565 1835 -525 1865
rect -565 1815 -555 1835
rect -535 1815 -525 1835
rect -565 1785 -525 1815
rect -565 1765 -555 1785
rect -535 1765 -525 1785
rect -565 1750 -525 1765
rect -505 2085 -465 2100
rect -505 2065 -495 2085
rect -475 2065 -465 2085
rect -505 2035 -465 2065
rect -505 2015 -495 2035
rect -475 2015 -465 2035
rect -505 1985 -465 2015
rect -505 1965 -495 1985
rect -475 1965 -465 1985
rect -505 1935 -465 1965
rect -505 1915 -495 1935
rect -475 1915 -465 1935
rect -505 1885 -465 1915
rect -505 1865 -495 1885
rect -475 1865 -465 1885
rect -505 1835 -465 1865
rect -505 1815 -495 1835
rect -475 1815 -465 1835
rect -505 1785 -465 1815
rect -505 1765 -495 1785
rect -475 1765 -465 1785
rect -505 1750 -465 1765
rect -445 2085 -405 2100
rect -445 2065 -435 2085
rect -415 2065 -405 2085
rect -445 2035 -405 2065
rect -445 2015 -435 2035
rect -415 2015 -405 2035
rect -445 1985 -405 2015
rect -445 1965 -435 1985
rect -415 1965 -405 1985
rect -445 1935 -405 1965
rect -445 1915 -435 1935
rect -415 1915 -405 1935
rect -445 1885 -405 1915
rect -445 1865 -435 1885
rect -415 1865 -405 1885
rect -445 1835 -405 1865
rect -445 1815 -435 1835
rect -415 1815 -405 1835
rect -445 1785 -405 1815
rect -445 1765 -435 1785
rect -415 1765 -405 1785
rect -445 1750 -405 1765
rect -40 2085 0 2100
rect -40 2065 -30 2085
rect -10 2065 0 2085
rect -40 2035 0 2065
rect -40 2015 -30 2035
rect -10 2015 0 2035
rect -40 1985 0 2015
rect -40 1965 -30 1985
rect -10 1965 0 1985
rect -40 1935 0 1965
rect -40 1915 -30 1935
rect -10 1915 0 1935
rect -40 1885 0 1915
rect -40 1865 -30 1885
rect -10 1865 0 1885
rect -40 1835 0 1865
rect -40 1815 -30 1835
rect -10 1815 0 1835
rect -40 1785 0 1815
rect -40 1765 -30 1785
rect -10 1765 0 1785
rect -40 1750 0 1765
rect 20 2085 60 2100
rect 20 2065 30 2085
rect 50 2065 60 2085
rect 20 2035 60 2065
rect 20 2015 30 2035
rect 50 2015 60 2035
rect 20 1985 60 2015
rect 20 1965 30 1985
rect 50 1965 60 1985
rect 20 1935 60 1965
rect 20 1915 30 1935
rect 50 1915 60 1935
rect 20 1885 60 1915
rect 20 1865 30 1885
rect 50 1865 60 1885
rect 20 1835 60 1865
rect 20 1815 30 1835
rect 50 1815 60 1835
rect 20 1785 60 1815
rect 20 1765 30 1785
rect 50 1765 60 1785
rect 20 1750 60 1765
rect 80 2085 120 2100
rect 80 2065 90 2085
rect 110 2065 120 2085
rect 80 2035 120 2065
rect 80 2015 90 2035
rect 110 2015 120 2035
rect 80 1985 120 2015
rect 80 1965 90 1985
rect 110 1965 120 1985
rect 80 1935 120 1965
rect 80 1915 90 1935
rect 110 1915 120 1935
rect 80 1885 120 1915
rect 80 1865 90 1885
rect 110 1865 120 1885
rect 80 1835 120 1865
rect 80 1815 90 1835
rect 110 1815 120 1835
rect 80 1785 120 1815
rect 80 1765 90 1785
rect 110 1765 120 1785
rect 80 1750 120 1765
rect 140 2085 180 2100
rect 140 2065 150 2085
rect 170 2065 180 2085
rect 140 2035 180 2065
rect 140 2015 150 2035
rect 170 2015 180 2035
rect 140 1985 180 2015
rect 140 1965 150 1985
rect 170 1965 180 1985
rect 140 1935 180 1965
rect 140 1915 150 1935
rect 170 1915 180 1935
rect 140 1885 180 1915
rect 140 1865 150 1885
rect 170 1865 180 1885
rect 140 1835 180 1865
rect 140 1815 150 1835
rect 170 1815 180 1835
rect 140 1785 180 1815
rect 140 1765 150 1785
rect 170 1765 180 1785
rect 140 1750 180 1765
rect 200 2085 240 2100
rect 200 2065 210 2085
rect 230 2065 240 2085
rect 200 2035 240 2065
rect 200 2015 210 2035
rect 230 2015 240 2035
rect 200 1985 240 2015
rect 200 1965 210 1985
rect 230 1965 240 1985
rect 200 1935 240 1965
rect 200 1915 210 1935
rect 230 1915 240 1935
rect 200 1885 240 1915
rect 200 1865 210 1885
rect 230 1865 240 1885
rect 200 1835 240 1865
rect 200 1815 210 1835
rect 230 1815 240 1835
rect 200 1785 240 1815
rect 200 1765 210 1785
rect 230 1765 240 1785
rect 200 1750 240 1765
rect 260 2085 300 2100
rect 260 2065 270 2085
rect 290 2065 300 2085
rect 260 2035 300 2065
rect 260 2015 270 2035
rect 290 2015 300 2035
rect 260 1985 300 2015
rect 260 1965 270 1985
rect 290 1965 300 1985
rect 260 1935 300 1965
rect 260 1915 270 1935
rect 290 1915 300 1935
rect 260 1885 300 1915
rect 260 1865 270 1885
rect 290 1865 300 1885
rect 260 1835 300 1865
rect 260 1815 270 1835
rect 290 1815 300 1835
rect 260 1785 300 1815
rect 260 1765 270 1785
rect 290 1765 300 1785
rect 260 1750 300 1765
rect 320 2085 360 2100
rect 320 2065 330 2085
rect 350 2065 360 2085
rect 320 2035 360 2065
rect 320 2015 330 2035
rect 350 2015 360 2035
rect 320 1985 360 2015
rect 320 1965 330 1985
rect 350 1965 360 1985
rect 320 1935 360 1965
rect 320 1915 330 1935
rect 350 1915 360 1935
rect 320 1885 360 1915
rect 320 1865 330 1885
rect 350 1865 360 1885
rect 320 1835 360 1865
rect 320 1815 330 1835
rect 350 1815 360 1835
rect 320 1785 360 1815
rect 320 1765 330 1785
rect 350 1765 360 1785
rect 320 1750 360 1765
rect 380 2085 420 2100
rect 380 2065 390 2085
rect 410 2065 420 2085
rect 380 2035 420 2065
rect 380 2015 390 2035
rect 410 2015 420 2035
rect 380 1985 420 2015
rect 380 1965 390 1985
rect 410 1965 420 1985
rect 380 1935 420 1965
rect 380 1915 390 1935
rect 410 1915 420 1935
rect 380 1885 420 1915
rect 380 1865 390 1885
rect 410 1865 420 1885
rect 380 1835 420 1865
rect 380 1815 390 1835
rect 410 1815 420 1835
rect 380 1785 420 1815
rect 380 1765 390 1785
rect 410 1765 420 1785
rect 380 1750 420 1765
rect 440 2085 480 2100
rect 440 2065 450 2085
rect 470 2065 480 2085
rect 440 2035 480 2065
rect 440 2015 450 2035
rect 470 2015 480 2035
rect 440 1985 480 2015
rect 440 1965 450 1985
rect 470 1965 480 1985
rect 440 1935 480 1965
rect 440 1915 450 1935
rect 470 1915 480 1935
rect 440 1885 480 1915
rect 440 1865 450 1885
rect 470 1865 480 1885
rect 440 1835 480 1865
rect 440 1815 450 1835
rect 470 1815 480 1835
rect 440 1785 480 1815
rect 440 1765 450 1785
rect 470 1765 480 1785
rect 440 1750 480 1765
rect 500 2085 540 2100
rect 500 2065 510 2085
rect 530 2065 540 2085
rect 500 2035 540 2065
rect 500 2015 510 2035
rect 530 2015 540 2035
rect 500 1985 540 2015
rect 500 1965 510 1985
rect 530 1965 540 1985
rect 500 1935 540 1965
rect 500 1915 510 1935
rect 530 1915 540 1935
rect 500 1885 540 1915
rect 500 1865 510 1885
rect 530 1865 540 1885
rect 500 1835 540 1865
rect 500 1815 510 1835
rect 530 1815 540 1835
rect 500 1785 540 1815
rect 500 1765 510 1785
rect 530 1765 540 1785
rect 500 1750 540 1765
rect 560 2085 600 2100
rect 560 2065 570 2085
rect 590 2065 600 2085
rect 560 2035 600 2065
rect 560 2015 570 2035
rect 590 2015 600 2035
rect 560 1985 600 2015
rect 560 1965 570 1985
rect 590 1965 600 1985
rect 560 1935 600 1965
rect 560 1915 570 1935
rect 590 1915 600 1935
rect 560 1885 600 1915
rect 560 1865 570 1885
rect 590 1865 600 1885
rect 560 1835 600 1865
rect 560 1815 570 1835
rect 590 1815 600 1835
rect 560 1785 600 1815
rect 560 1765 570 1785
rect 590 1765 600 1785
rect 560 1750 600 1765
rect 620 2085 660 2100
rect 620 2065 630 2085
rect 650 2065 660 2085
rect 620 2035 660 2065
rect 620 2015 630 2035
rect 650 2015 660 2035
rect 620 1985 660 2015
rect 620 1965 630 1985
rect 650 1965 660 1985
rect 620 1935 660 1965
rect 620 1915 630 1935
rect 650 1915 660 1935
rect 620 1885 660 1915
rect 620 1865 630 1885
rect 650 1865 660 1885
rect 620 1835 660 1865
rect 620 1815 630 1835
rect 650 1815 660 1835
rect 620 1785 660 1815
rect 620 1765 630 1785
rect 650 1765 660 1785
rect 620 1750 660 1765
rect 680 2085 720 2100
rect 680 2065 690 2085
rect 710 2065 720 2085
rect 680 2035 720 2065
rect 680 2015 690 2035
rect 710 2015 720 2035
rect 680 1985 720 2015
rect 680 1965 690 1985
rect 710 1965 720 1985
rect 680 1935 720 1965
rect 680 1915 690 1935
rect 710 1915 720 1935
rect 680 1885 720 1915
rect 680 1865 690 1885
rect 710 1865 720 1885
rect 680 1835 720 1865
rect 680 1815 690 1835
rect 710 1815 720 1835
rect 680 1785 720 1815
rect 680 1765 690 1785
rect 710 1765 720 1785
rect 680 1750 720 1765
rect 970 2085 1010 2100
rect 970 2065 980 2085
rect 1000 2065 1010 2085
rect 970 2035 1010 2065
rect 970 2015 980 2035
rect 1000 2015 1010 2035
rect 970 1985 1010 2015
rect 970 1965 980 1985
rect 1000 1965 1010 1985
rect 970 1935 1010 1965
rect 970 1915 980 1935
rect 1000 1915 1010 1935
rect 970 1885 1010 1915
rect 970 1865 980 1885
rect 1000 1865 1010 1885
rect 970 1835 1010 1865
rect 970 1815 980 1835
rect 1000 1815 1010 1835
rect 970 1785 1010 1815
rect 970 1765 980 1785
rect 1000 1765 1010 1785
rect 970 1750 1010 1765
rect 1030 2085 1070 2100
rect 1030 2065 1040 2085
rect 1060 2065 1070 2085
rect 1030 2035 1070 2065
rect 1030 2015 1040 2035
rect 1060 2015 1070 2035
rect 1030 1985 1070 2015
rect 1030 1965 1040 1985
rect 1060 1965 1070 1985
rect 1030 1935 1070 1965
rect 1030 1915 1040 1935
rect 1060 1915 1070 1935
rect 1030 1885 1070 1915
rect 1030 1865 1040 1885
rect 1060 1865 1070 1885
rect 1030 1835 1070 1865
rect 1030 1815 1040 1835
rect 1060 1815 1070 1835
rect 1030 1785 1070 1815
rect 1030 1765 1040 1785
rect 1060 1765 1070 1785
rect 1030 1750 1070 1765
rect 1090 2085 1130 2100
rect 1090 2065 1100 2085
rect 1120 2065 1130 2085
rect 1090 2035 1130 2065
rect 1090 2015 1100 2035
rect 1120 2015 1130 2035
rect 1090 1985 1130 2015
rect 1090 1965 1100 1985
rect 1120 1965 1130 1985
rect 1090 1935 1130 1965
rect 1090 1915 1100 1935
rect 1120 1915 1130 1935
rect 1090 1885 1130 1915
rect 1090 1865 1100 1885
rect 1120 1865 1130 1885
rect 1090 1835 1130 1865
rect 1090 1815 1100 1835
rect 1120 1815 1130 1835
rect 1090 1785 1130 1815
rect 1090 1765 1100 1785
rect 1120 1765 1130 1785
rect 1090 1750 1130 1765
rect 1150 2085 1190 2100
rect 1150 2065 1160 2085
rect 1180 2065 1190 2085
rect 1150 2035 1190 2065
rect 1150 2015 1160 2035
rect 1180 2015 1190 2035
rect 1150 1985 1190 2015
rect 1150 1965 1160 1985
rect 1180 1965 1190 1985
rect 1150 1935 1190 1965
rect 1150 1915 1160 1935
rect 1180 1915 1190 1935
rect 1150 1885 1190 1915
rect 1150 1865 1160 1885
rect 1180 1865 1190 1885
rect 1150 1835 1190 1865
rect 1150 1815 1160 1835
rect 1180 1815 1190 1835
rect 1150 1785 1190 1815
rect 1150 1765 1160 1785
rect 1180 1765 1190 1785
rect 1150 1750 1190 1765
rect 1210 2085 1250 2100
rect 1210 2065 1220 2085
rect 1240 2065 1250 2085
rect 1210 2035 1250 2065
rect 1210 2015 1220 2035
rect 1240 2015 1250 2035
rect 1210 1985 1250 2015
rect 1210 1965 1220 1985
rect 1240 1965 1250 1985
rect 1210 1935 1250 1965
rect 1210 1915 1220 1935
rect 1240 1915 1250 1935
rect 1210 1885 1250 1915
rect 1210 1865 1220 1885
rect 1240 1865 1250 1885
rect 1210 1835 1250 1865
rect 1210 1815 1220 1835
rect 1240 1815 1250 1835
rect 1210 1785 1250 1815
rect 1210 1765 1220 1785
rect 1240 1765 1250 1785
rect 1210 1750 1250 1765
rect 1270 2085 1310 2100
rect 1270 2065 1280 2085
rect 1300 2065 1310 2085
rect 1270 2035 1310 2065
rect 1270 2015 1280 2035
rect 1300 2015 1310 2035
rect 1270 1985 1310 2015
rect 1270 1965 1280 1985
rect 1300 1965 1310 1985
rect 1270 1935 1310 1965
rect 1270 1915 1280 1935
rect 1300 1915 1310 1935
rect 1270 1885 1310 1915
rect 1270 1865 1280 1885
rect 1300 1865 1310 1885
rect 1270 1835 1310 1865
rect 1270 1815 1280 1835
rect 1300 1815 1310 1835
rect 1270 1785 1310 1815
rect 1270 1765 1280 1785
rect 1300 1765 1310 1785
rect 1270 1750 1310 1765
rect 1330 2085 1370 2100
rect 1330 2065 1340 2085
rect 1360 2065 1370 2085
rect 1330 2035 1370 2065
rect 1330 2015 1340 2035
rect 1360 2015 1370 2035
rect 1330 1985 1370 2015
rect 1330 1965 1340 1985
rect 1360 1965 1370 1985
rect 1330 1935 1370 1965
rect 1330 1915 1340 1935
rect 1360 1915 1370 1935
rect 1330 1885 1370 1915
rect 1330 1865 1340 1885
rect 1360 1865 1370 1885
rect 1330 1835 1370 1865
rect 1330 1815 1340 1835
rect 1360 1815 1370 1835
rect 1330 1785 1370 1815
rect 1330 1765 1340 1785
rect 1360 1765 1370 1785
rect 1330 1750 1370 1765
rect 1390 2085 1430 2100
rect 1390 2065 1400 2085
rect 1420 2065 1430 2085
rect 1390 2035 1430 2065
rect 1390 2015 1400 2035
rect 1420 2015 1430 2035
rect 1390 1985 1430 2015
rect 1390 1965 1400 1985
rect 1420 1965 1430 1985
rect 1390 1935 1430 1965
rect 1390 1915 1400 1935
rect 1420 1915 1430 1935
rect 1390 1885 1430 1915
rect 1390 1865 1400 1885
rect 1420 1865 1430 1885
rect 1390 1835 1430 1865
rect 1390 1815 1400 1835
rect 1420 1815 1430 1835
rect 1390 1785 1430 1815
rect 1390 1765 1400 1785
rect 1420 1765 1430 1785
rect 1390 1750 1430 1765
rect 1450 2085 1490 2100
rect 1450 2065 1460 2085
rect 1480 2065 1490 2085
rect 1450 2035 1490 2065
rect 1450 2015 1460 2035
rect 1480 2015 1490 2035
rect 1450 1985 1490 2015
rect 1450 1965 1460 1985
rect 1480 1965 1490 1985
rect 1450 1935 1490 1965
rect 1450 1915 1460 1935
rect 1480 1915 1490 1935
rect 1450 1885 1490 1915
rect 1450 1865 1460 1885
rect 1480 1865 1490 1885
rect 1450 1835 1490 1865
rect 1450 1815 1460 1835
rect 1480 1815 1490 1835
rect 1450 1785 1490 1815
rect 1450 1765 1460 1785
rect 1480 1765 1490 1785
rect 1450 1750 1490 1765
rect 1510 2085 1550 2100
rect 1510 2065 1520 2085
rect 1540 2065 1550 2085
rect 1510 2035 1550 2065
rect 1510 2015 1520 2035
rect 1540 2015 1550 2035
rect 1510 1985 1550 2015
rect 1510 1965 1520 1985
rect 1540 1965 1550 1985
rect 1510 1935 1550 1965
rect 1510 1915 1520 1935
rect 1540 1915 1550 1935
rect 1510 1885 1550 1915
rect 1510 1865 1520 1885
rect 1540 1865 1550 1885
rect 1510 1835 1550 1865
rect 1510 1815 1520 1835
rect 1540 1815 1550 1835
rect 1510 1785 1550 1815
rect 1510 1765 1520 1785
rect 1540 1765 1550 1785
rect 1510 1750 1550 1765
rect 1570 2085 1610 2100
rect 1570 2065 1580 2085
rect 1600 2065 1610 2085
rect 1570 2035 1610 2065
rect 1570 2015 1580 2035
rect 1600 2015 1610 2035
rect 1570 1985 1610 2015
rect 1570 1965 1580 1985
rect 1600 1965 1610 1985
rect 1570 1935 1610 1965
rect 1570 1915 1580 1935
rect 1600 1915 1610 1935
rect 1570 1885 1610 1915
rect 1570 1865 1580 1885
rect 1600 1865 1610 1885
rect 1570 1835 1610 1865
rect 1570 1815 1580 1835
rect 1600 1815 1610 1835
rect 1570 1785 1610 1815
rect 1570 1765 1580 1785
rect 1600 1765 1610 1785
rect 1570 1750 1610 1765
rect 1630 2085 1670 2100
rect 1630 2065 1640 2085
rect 1660 2065 1670 2085
rect 1630 2035 1670 2065
rect 1630 2015 1640 2035
rect 1660 2015 1670 2035
rect 1630 1985 1670 2015
rect 1630 1965 1640 1985
rect 1660 1965 1670 1985
rect 1630 1935 1670 1965
rect 1630 1915 1640 1935
rect 1660 1915 1670 1935
rect 1630 1885 1670 1915
rect 1630 1865 1640 1885
rect 1660 1865 1670 1885
rect 1630 1835 1670 1865
rect 1630 1815 1640 1835
rect 1660 1815 1670 1835
rect 1630 1785 1670 1815
rect 1630 1765 1640 1785
rect 1660 1765 1670 1785
rect 1630 1750 1670 1765
rect 1690 2085 1730 2100
rect 1690 2065 1700 2085
rect 1720 2065 1730 2085
rect 1690 2035 1730 2065
rect 1690 2015 1700 2035
rect 1720 2015 1730 2035
rect 1690 1985 1730 2015
rect 1690 1965 1700 1985
rect 1720 1965 1730 1985
rect 1690 1935 1730 1965
rect 1690 1915 1700 1935
rect 1720 1915 1730 1935
rect 1690 1885 1730 1915
rect 1690 1865 1700 1885
rect 1720 1865 1730 1885
rect 1690 1835 1730 1865
rect 1690 1815 1700 1835
rect 1720 1815 1730 1835
rect 1690 1785 1730 1815
rect 1690 1765 1700 1785
rect 1720 1765 1730 1785
rect 1690 1750 1730 1765
rect 2095 2085 2135 2100
rect 2095 2065 2105 2085
rect 2125 2065 2135 2085
rect 2095 2035 2135 2065
rect 2095 2015 2105 2035
rect 2125 2015 2135 2035
rect 2095 1985 2135 2015
rect 2095 1965 2105 1985
rect 2125 1965 2135 1985
rect 2095 1935 2135 1965
rect 2095 1915 2105 1935
rect 2125 1915 2135 1935
rect 2095 1885 2135 1915
rect 2095 1865 2105 1885
rect 2125 1865 2135 1885
rect 2095 1835 2135 1865
rect 2095 1815 2105 1835
rect 2125 1815 2135 1835
rect 2095 1785 2135 1815
rect 2095 1765 2105 1785
rect 2125 1765 2135 1785
rect 2095 1750 2135 1765
rect 2155 2085 2195 2100
rect 2155 2065 2165 2085
rect 2185 2065 2195 2085
rect 2155 2035 2195 2065
rect 2155 2015 2165 2035
rect 2185 2015 2195 2035
rect 2155 1985 2195 2015
rect 2155 1965 2165 1985
rect 2185 1965 2195 1985
rect 2155 1935 2195 1965
rect 2155 1915 2165 1935
rect 2185 1915 2195 1935
rect 2155 1885 2195 1915
rect 2155 1865 2165 1885
rect 2185 1865 2195 1885
rect 2155 1835 2195 1865
rect 2155 1815 2165 1835
rect 2185 1815 2195 1835
rect 2155 1785 2195 1815
rect 2155 1765 2165 1785
rect 2185 1765 2195 1785
rect 2155 1750 2195 1765
rect 2215 2085 2255 2100
rect 2215 2065 2225 2085
rect 2245 2065 2255 2085
rect 2215 2035 2255 2065
rect 2215 2015 2225 2035
rect 2245 2015 2255 2035
rect 2215 1985 2255 2015
rect 2215 1965 2225 1985
rect 2245 1965 2255 1985
rect 2215 1935 2255 1965
rect 2215 1915 2225 1935
rect 2245 1915 2255 1935
rect 2215 1885 2255 1915
rect 2215 1865 2225 1885
rect 2245 1865 2255 1885
rect 2215 1835 2255 1865
rect 2215 1815 2225 1835
rect 2245 1815 2255 1835
rect 2215 1785 2255 1815
rect 2215 1765 2225 1785
rect 2245 1765 2255 1785
rect 2215 1750 2255 1765
rect 2275 2085 2315 2100
rect 2275 2065 2285 2085
rect 2305 2065 2315 2085
rect 2275 2035 2315 2065
rect 2275 2015 2285 2035
rect 2305 2015 2315 2035
rect 2275 1985 2315 2015
rect 2275 1965 2285 1985
rect 2305 1965 2315 1985
rect 2275 1935 2315 1965
rect 2275 1915 2285 1935
rect 2305 1915 2315 1935
rect 2275 1885 2315 1915
rect 2275 1865 2285 1885
rect 2305 1865 2315 1885
rect 2275 1835 2315 1865
rect 2275 1815 2285 1835
rect 2305 1815 2315 1835
rect 2275 1785 2315 1815
rect 2275 1765 2285 1785
rect 2305 1765 2315 1785
rect 2275 1750 2315 1765
rect 2335 2085 2375 2100
rect 2335 2065 2345 2085
rect 2365 2065 2375 2085
rect 2335 2035 2375 2065
rect 2335 2015 2345 2035
rect 2365 2015 2375 2035
rect 2335 1985 2375 2015
rect 2335 1965 2345 1985
rect 2365 1965 2375 1985
rect 2335 1935 2375 1965
rect 2335 1915 2345 1935
rect 2365 1915 2375 1935
rect 2335 1885 2375 1915
rect 2335 1865 2345 1885
rect 2365 1865 2375 1885
rect 2335 1835 2375 1865
rect 2335 1815 2345 1835
rect 2365 1815 2375 1835
rect 2335 1785 2375 1815
rect 2335 1765 2345 1785
rect 2365 1765 2375 1785
rect 2335 1750 2375 1765
rect 2395 2085 2435 2100
rect 2395 2065 2405 2085
rect 2425 2065 2435 2085
rect 2395 2035 2435 2065
rect 2395 2015 2405 2035
rect 2425 2015 2435 2035
rect 2395 1985 2435 2015
rect 2395 1965 2405 1985
rect 2425 1965 2435 1985
rect 2395 1935 2435 1965
rect 2395 1915 2405 1935
rect 2425 1915 2435 1935
rect 2395 1885 2435 1915
rect 2395 1865 2405 1885
rect 2425 1865 2435 1885
rect 2395 1835 2435 1865
rect 2395 1815 2405 1835
rect 2425 1815 2435 1835
rect 2395 1785 2435 1815
rect 2395 1765 2405 1785
rect 2425 1765 2435 1785
rect 2395 1750 2435 1765
rect 2455 2085 2495 2100
rect 2455 2065 2465 2085
rect 2485 2065 2495 2085
rect 2455 2035 2495 2065
rect 2455 2015 2465 2035
rect 2485 2015 2495 2035
rect 2455 1985 2495 2015
rect 2455 1965 2465 1985
rect 2485 1965 2495 1985
rect 2455 1935 2495 1965
rect 2455 1915 2465 1935
rect 2485 1915 2495 1935
rect 2455 1885 2495 1915
rect 2455 1865 2465 1885
rect 2485 1865 2495 1885
rect 2455 1835 2495 1865
rect 2455 1815 2465 1835
rect 2485 1815 2495 1835
rect 2455 1785 2495 1815
rect 2455 1765 2465 1785
rect 2485 1765 2495 1785
rect 2455 1750 2495 1765
rect 2515 2085 2555 2100
rect 2515 2065 2525 2085
rect 2545 2065 2555 2085
rect 2515 2035 2555 2065
rect 2515 2015 2525 2035
rect 2545 2015 2555 2035
rect 2515 1985 2555 2015
rect 2515 1965 2525 1985
rect 2545 1965 2555 1985
rect 2515 1935 2555 1965
rect 2515 1915 2525 1935
rect 2545 1915 2555 1935
rect 2515 1885 2555 1915
rect 2515 1865 2525 1885
rect 2545 1865 2555 1885
rect 2515 1835 2555 1865
rect 2515 1815 2525 1835
rect 2545 1815 2555 1835
rect 2515 1785 2555 1815
rect 2515 1765 2525 1785
rect 2545 1765 2555 1785
rect 2515 1750 2555 1765
rect 2575 2085 2615 2100
rect 2575 2065 2585 2085
rect 2605 2065 2615 2085
rect 2575 2035 2615 2065
rect 2575 2015 2585 2035
rect 2605 2015 2615 2035
rect 2575 1985 2615 2015
rect 2575 1965 2585 1985
rect 2605 1965 2615 1985
rect 2575 1935 2615 1965
rect 2575 1915 2585 1935
rect 2605 1915 2615 1935
rect 2575 1885 2615 1915
rect 2575 1865 2585 1885
rect 2605 1865 2615 1885
rect 2575 1835 2615 1865
rect 2575 1815 2585 1835
rect 2605 1815 2615 1835
rect 2575 1785 2615 1815
rect 2575 1765 2585 1785
rect 2605 1765 2615 1785
rect 2575 1750 2615 1765
rect 2635 2085 2675 2100
rect 2635 2065 2645 2085
rect 2665 2065 2675 2085
rect 2635 2035 2675 2065
rect 2635 2015 2645 2035
rect 2665 2015 2675 2035
rect 2635 1985 2675 2015
rect 2635 1965 2645 1985
rect 2665 1965 2675 1985
rect 2635 1935 2675 1965
rect 2635 1915 2645 1935
rect 2665 1915 2675 1935
rect 2635 1885 2675 1915
rect 2635 1865 2645 1885
rect 2665 1865 2675 1885
rect 2635 1835 2675 1865
rect 2635 1815 2645 1835
rect 2665 1815 2675 1835
rect 2635 1785 2675 1815
rect 2635 1765 2645 1785
rect 2665 1765 2675 1785
rect 2635 1750 2675 1765
rect 2695 2085 2735 2100
rect 2695 2065 2705 2085
rect 2725 2065 2735 2085
rect 2695 2035 2735 2065
rect 2695 2015 2705 2035
rect 2725 2015 2735 2035
rect 2695 1985 2735 2015
rect 2695 1965 2705 1985
rect 2725 1965 2735 1985
rect 2695 1935 2735 1965
rect 2695 1915 2705 1935
rect 2725 1915 2735 1935
rect 2695 1885 2735 1915
rect 2695 1865 2705 1885
rect 2725 1865 2735 1885
rect 2695 1835 2735 1865
rect 2695 1815 2705 1835
rect 2725 1815 2735 1835
rect 2695 1785 2735 1815
rect 2695 1765 2705 1785
rect 2725 1765 2735 1785
rect 2695 1750 2735 1765
rect 2755 2085 2795 2100
rect 2755 2065 2765 2085
rect 2785 2065 2795 2085
rect 2755 2035 2795 2065
rect 2755 2015 2765 2035
rect 2785 2015 2795 2035
rect 2755 1985 2795 2015
rect 2755 1965 2765 1985
rect 2785 1965 2795 1985
rect 2755 1935 2795 1965
rect 2755 1915 2765 1935
rect 2785 1915 2795 1935
rect 2755 1885 2795 1915
rect 2755 1865 2765 1885
rect 2785 1865 2795 1885
rect 2755 1835 2795 1865
rect 2755 1815 2765 1835
rect 2785 1815 2795 1835
rect 2755 1785 2795 1815
rect 2755 1765 2765 1785
rect 2785 1765 2795 1785
rect 2755 1750 2795 1765
rect 2815 2085 2855 2100
rect 2815 2065 2825 2085
rect 2845 2065 2855 2085
rect 2815 2035 2855 2065
rect 2815 2015 2825 2035
rect 2845 2015 2855 2035
rect 2815 1985 2855 2015
rect 2815 1965 2825 1985
rect 2845 1965 2855 1985
rect 2815 1935 2855 1965
rect 2815 1915 2825 1935
rect 2845 1915 2855 1935
rect 2815 1885 2855 1915
rect 2815 1865 2825 1885
rect 2845 1865 2855 1885
rect 2815 1835 2855 1865
rect 2815 1815 2825 1835
rect 2845 1815 2855 1835
rect 2815 1785 2855 1815
rect 2815 1765 2825 1785
rect 2845 1765 2855 1785
rect 2815 1750 2855 1765
rect 455 1470 495 1485
rect 455 1450 465 1470
rect 485 1450 495 1470
rect -1135 1420 -1095 1435
rect -1135 1400 -1125 1420
rect -1105 1400 -1095 1420
rect -1135 1370 -1095 1400
rect -1135 1350 -1125 1370
rect -1105 1350 -1095 1370
rect -1135 1320 -1095 1350
rect -1135 1300 -1125 1320
rect -1105 1300 -1095 1320
rect -1135 1270 -1095 1300
rect -1135 1250 -1125 1270
rect -1105 1250 -1095 1270
rect -1135 1220 -1095 1250
rect -1135 1200 -1125 1220
rect -1105 1200 -1095 1220
rect -1135 1170 -1095 1200
rect -1135 1150 -1125 1170
rect -1105 1150 -1095 1170
rect -1135 1120 -1095 1150
rect -1135 1100 -1125 1120
rect -1105 1100 -1095 1120
rect -1135 1070 -1095 1100
rect -1135 1050 -1125 1070
rect -1105 1050 -1095 1070
rect -1135 1020 -1095 1050
rect -1135 1000 -1125 1020
rect -1105 1000 -1095 1020
rect -1135 970 -1095 1000
rect -1135 950 -1125 970
rect -1105 950 -1095 970
rect -1135 920 -1095 950
rect -1135 900 -1125 920
rect -1105 900 -1095 920
rect -1135 870 -1095 900
rect -1135 850 -1125 870
rect -1105 850 -1095 870
rect -1135 835 -1095 850
rect -1080 1420 -1040 1435
rect -1080 1400 -1070 1420
rect -1050 1400 -1040 1420
rect -1080 1370 -1040 1400
rect -1080 1350 -1070 1370
rect -1050 1350 -1040 1370
rect -1080 1320 -1040 1350
rect -1080 1300 -1070 1320
rect -1050 1300 -1040 1320
rect -1080 1270 -1040 1300
rect -1080 1250 -1070 1270
rect -1050 1250 -1040 1270
rect -1080 1220 -1040 1250
rect -1080 1200 -1070 1220
rect -1050 1200 -1040 1220
rect -1080 1170 -1040 1200
rect -1080 1150 -1070 1170
rect -1050 1150 -1040 1170
rect -1080 1120 -1040 1150
rect -1080 1100 -1070 1120
rect -1050 1100 -1040 1120
rect -1080 1070 -1040 1100
rect -1080 1050 -1070 1070
rect -1050 1050 -1040 1070
rect -1080 1020 -1040 1050
rect -1080 1000 -1070 1020
rect -1050 1000 -1040 1020
rect -1080 970 -1040 1000
rect -1080 950 -1070 970
rect -1050 950 -1040 970
rect -1080 920 -1040 950
rect -1080 900 -1070 920
rect -1050 900 -1040 920
rect -1080 870 -1040 900
rect -1080 850 -1070 870
rect -1050 850 -1040 870
rect -1080 835 -1040 850
rect -1025 1420 -985 1435
rect -1025 1400 -1015 1420
rect -995 1400 -985 1420
rect -1025 1370 -985 1400
rect -1025 1350 -1015 1370
rect -995 1350 -985 1370
rect -1025 1320 -985 1350
rect -1025 1300 -1015 1320
rect -995 1300 -985 1320
rect -1025 1270 -985 1300
rect -1025 1250 -1015 1270
rect -995 1250 -985 1270
rect -1025 1220 -985 1250
rect -1025 1200 -1015 1220
rect -995 1200 -985 1220
rect -1025 1170 -985 1200
rect -1025 1150 -1015 1170
rect -995 1150 -985 1170
rect -1025 1120 -985 1150
rect -1025 1100 -1015 1120
rect -995 1100 -985 1120
rect -1025 1070 -985 1100
rect -1025 1050 -1015 1070
rect -995 1050 -985 1070
rect -1025 1020 -985 1050
rect -1025 1000 -1015 1020
rect -995 1000 -985 1020
rect -1025 970 -985 1000
rect -1025 950 -1015 970
rect -995 950 -985 970
rect -1025 920 -985 950
rect -1025 900 -1015 920
rect -995 900 -985 920
rect -1025 870 -985 900
rect -1025 850 -1015 870
rect -995 850 -985 870
rect -1025 835 -985 850
rect -970 1420 -930 1435
rect -970 1400 -960 1420
rect -940 1400 -930 1420
rect -970 1370 -930 1400
rect -970 1350 -960 1370
rect -940 1350 -930 1370
rect -970 1320 -930 1350
rect -970 1300 -960 1320
rect -940 1300 -930 1320
rect -970 1270 -930 1300
rect -970 1250 -960 1270
rect -940 1250 -930 1270
rect -970 1220 -930 1250
rect -970 1200 -960 1220
rect -940 1200 -930 1220
rect -970 1170 -930 1200
rect -970 1150 -960 1170
rect -940 1150 -930 1170
rect -970 1120 -930 1150
rect -970 1100 -960 1120
rect -940 1100 -930 1120
rect -970 1070 -930 1100
rect -970 1050 -960 1070
rect -940 1050 -930 1070
rect -970 1020 -930 1050
rect -970 1000 -960 1020
rect -940 1000 -930 1020
rect -970 970 -930 1000
rect -970 950 -960 970
rect -940 950 -930 970
rect -970 920 -930 950
rect -970 900 -960 920
rect -940 900 -930 920
rect -970 870 -930 900
rect -970 850 -960 870
rect -940 850 -930 870
rect -970 835 -930 850
rect -915 1420 -875 1435
rect -915 1400 -905 1420
rect -885 1400 -875 1420
rect -915 1370 -875 1400
rect -915 1350 -905 1370
rect -885 1350 -875 1370
rect -915 1320 -875 1350
rect -915 1300 -905 1320
rect -885 1300 -875 1320
rect -915 1270 -875 1300
rect -915 1250 -905 1270
rect -885 1250 -875 1270
rect -915 1220 -875 1250
rect -915 1200 -905 1220
rect -885 1200 -875 1220
rect -915 1170 -875 1200
rect -915 1150 -905 1170
rect -885 1150 -875 1170
rect -915 1120 -875 1150
rect -915 1100 -905 1120
rect -885 1100 -875 1120
rect -915 1070 -875 1100
rect -915 1050 -905 1070
rect -885 1050 -875 1070
rect -915 1020 -875 1050
rect -915 1000 -905 1020
rect -885 1000 -875 1020
rect -915 970 -875 1000
rect -915 950 -905 970
rect -885 950 -875 970
rect -915 920 -875 950
rect -915 900 -905 920
rect -885 900 -875 920
rect -915 870 -875 900
rect -915 850 -905 870
rect -885 850 -875 870
rect -915 835 -875 850
rect -860 1420 -820 1435
rect -860 1400 -850 1420
rect -830 1400 -820 1420
rect -860 1370 -820 1400
rect -860 1350 -850 1370
rect -830 1350 -820 1370
rect -860 1320 -820 1350
rect -860 1300 -850 1320
rect -830 1300 -820 1320
rect -860 1270 -820 1300
rect -860 1250 -850 1270
rect -830 1250 -820 1270
rect -860 1220 -820 1250
rect -860 1200 -850 1220
rect -830 1200 -820 1220
rect -860 1170 -820 1200
rect -860 1150 -850 1170
rect -830 1150 -820 1170
rect -860 1120 -820 1150
rect -860 1100 -850 1120
rect -830 1100 -820 1120
rect -860 1070 -820 1100
rect -860 1050 -850 1070
rect -830 1050 -820 1070
rect -860 1020 -820 1050
rect -860 1000 -850 1020
rect -830 1000 -820 1020
rect -860 970 -820 1000
rect -860 950 -850 970
rect -830 950 -820 970
rect -860 920 -820 950
rect -860 900 -850 920
rect -830 900 -820 920
rect -860 870 -820 900
rect -860 850 -850 870
rect -830 850 -820 870
rect -860 835 -820 850
rect -805 1420 -765 1435
rect -805 1400 -795 1420
rect -775 1400 -765 1420
rect -805 1370 -765 1400
rect -805 1350 -795 1370
rect -775 1350 -765 1370
rect -805 1320 -765 1350
rect -805 1300 -795 1320
rect -775 1300 -765 1320
rect -805 1270 -765 1300
rect -805 1250 -795 1270
rect -775 1250 -765 1270
rect -805 1220 -765 1250
rect -805 1200 -795 1220
rect -775 1200 -765 1220
rect -805 1170 -765 1200
rect -805 1150 -795 1170
rect -775 1150 -765 1170
rect -805 1120 -765 1150
rect -805 1100 -795 1120
rect -775 1100 -765 1120
rect -805 1070 -765 1100
rect -805 1050 -795 1070
rect -775 1050 -765 1070
rect -805 1020 -765 1050
rect -805 1000 -795 1020
rect -775 1000 -765 1020
rect -805 970 -765 1000
rect -805 950 -795 970
rect -775 950 -765 970
rect -805 920 -765 950
rect -805 900 -795 920
rect -775 900 -765 920
rect -805 870 -765 900
rect -805 850 -795 870
rect -775 850 -765 870
rect -805 835 -765 850
rect -750 1420 -710 1435
rect -750 1400 -740 1420
rect -720 1400 -710 1420
rect -750 1370 -710 1400
rect -750 1350 -740 1370
rect -720 1350 -710 1370
rect -750 1320 -710 1350
rect -750 1300 -740 1320
rect -720 1300 -710 1320
rect -750 1270 -710 1300
rect -750 1250 -740 1270
rect -720 1250 -710 1270
rect -750 1220 -710 1250
rect -750 1200 -740 1220
rect -720 1200 -710 1220
rect -750 1170 -710 1200
rect -750 1150 -740 1170
rect -720 1150 -710 1170
rect -750 1120 -710 1150
rect -750 1100 -740 1120
rect -720 1100 -710 1120
rect -750 1070 -710 1100
rect -750 1050 -740 1070
rect -720 1050 -710 1070
rect -750 1020 -710 1050
rect -750 1000 -740 1020
rect -720 1000 -710 1020
rect -750 970 -710 1000
rect -750 950 -740 970
rect -720 950 -710 970
rect -750 920 -710 950
rect -750 900 -740 920
rect -720 900 -710 920
rect -750 870 -710 900
rect -750 850 -740 870
rect -720 850 -710 870
rect -750 835 -710 850
rect -695 1420 -655 1435
rect -695 1400 -685 1420
rect -665 1400 -655 1420
rect -695 1370 -655 1400
rect -695 1350 -685 1370
rect -665 1350 -655 1370
rect -695 1320 -655 1350
rect -695 1300 -685 1320
rect -665 1300 -655 1320
rect -695 1270 -655 1300
rect -695 1250 -685 1270
rect -665 1250 -655 1270
rect -695 1220 -655 1250
rect -695 1200 -685 1220
rect -665 1200 -655 1220
rect -695 1170 -655 1200
rect -695 1150 -685 1170
rect -665 1150 -655 1170
rect -695 1120 -655 1150
rect -695 1100 -685 1120
rect -665 1100 -655 1120
rect -695 1070 -655 1100
rect -695 1050 -685 1070
rect -665 1050 -655 1070
rect -695 1020 -655 1050
rect -695 1000 -685 1020
rect -665 1000 -655 1020
rect -695 970 -655 1000
rect -695 950 -685 970
rect -665 950 -655 970
rect -695 920 -655 950
rect -695 900 -685 920
rect -665 900 -655 920
rect -695 870 -655 900
rect -695 850 -685 870
rect -665 850 -655 870
rect -695 835 -655 850
rect -640 1420 -600 1435
rect -640 1400 -630 1420
rect -610 1400 -600 1420
rect -640 1370 -600 1400
rect -640 1350 -630 1370
rect -610 1350 -600 1370
rect -640 1320 -600 1350
rect -640 1300 -630 1320
rect -610 1300 -600 1320
rect -640 1270 -600 1300
rect -640 1250 -630 1270
rect -610 1250 -600 1270
rect -640 1220 -600 1250
rect -640 1200 -630 1220
rect -610 1200 -600 1220
rect -640 1170 -600 1200
rect -640 1150 -630 1170
rect -610 1150 -600 1170
rect -640 1120 -600 1150
rect -640 1100 -630 1120
rect -610 1100 -600 1120
rect -640 1070 -600 1100
rect -640 1050 -630 1070
rect -610 1050 -600 1070
rect -640 1020 -600 1050
rect -640 1000 -630 1020
rect -610 1000 -600 1020
rect -640 970 -600 1000
rect -640 950 -630 970
rect -610 950 -600 970
rect -640 920 -600 950
rect -640 900 -630 920
rect -610 900 -600 920
rect -640 870 -600 900
rect -640 850 -630 870
rect -610 850 -600 870
rect -640 835 -600 850
rect -585 1420 -545 1435
rect -585 1400 -575 1420
rect -555 1400 -545 1420
rect -585 1370 -545 1400
rect -585 1350 -575 1370
rect -555 1350 -545 1370
rect -585 1320 -545 1350
rect -585 1300 -575 1320
rect -555 1300 -545 1320
rect -585 1270 -545 1300
rect -585 1250 -575 1270
rect -555 1250 -545 1270
rect -585 1220 -545 1250
rect -585 1200 -575 1220
rect -555 1200 -545 1220
rect -585 1170 -545 1200
rect -585 1150 -575 1170
rect -555 1150 -545 1170
rect -585 1120 -545 1150
rect -585 1100 -575 1120
rect -555 1100 -545 1120
rect -585 1070 -545 1100
rect -585 1050 -575 1070
rect -555 1050 -545 1070
rect -585 1020 -545 1050
rect -585 1000 -575 1020
rect -555 1000 -545 1020
rect -585 970 -545 1000
rect -585 950 -575 970
rect -555 950 -545 970
rect -585 920 -545 950
rect -585 900 -575 920
rect -555 900 -545 920
rect -585 870 -545 900
rect -585 850 -575 870
rect -555 850 -545 870
rect -585 835 -545 850
rect -530 1420 -490 1435
rect -530 1400 -520 1420
rect -500 1400 -490 1420
rect -530 1370 -490 1400
rect -530 1350 -520 1370
rect -500 1350 -490 1370
rect -530 1320 -490 1350
rect -530 1300 -520 1320
rect -500 1300 -490 1320
rect -530 1270 -490 1300
rect -530 1250 -520 1270
rect -500 1250 -490 1270
rect -530 1220 -490 1250
rect -530 1200 -520 1220
rect -500 1200 -490 1220
rect -530 1170 -490 1200
rect -530 1150 -520 1170
rect -500 1150 -490 1170
rect -530 1120 -490 1150
rect -530 1100 -520 1120
rect -500 1100 -490 1120
rect -530 1070 -490 1100
rect -530 1050 -520 1070
rect -500 1050 -490 1070
rect -530 1020 -490 1050
rect -530 1000 -520 1020
rect -500 1000 -490 1020
rect -530 970 -490 1000
rect -530 950 -520 970
rect -500 950 -490 970
rect -530 920 -490 950
rect -530 900 -520 920
rect -500 900 -490 920
rect -530 870 -490 900
rect -530 850 -520 870
rect -500 850 -490 870
rect -530 835 -490 850
rect -475 1420 -435 1435
rect -475 1400 -465 1420
rect -445 1400 -435 1420
rect -475 1370 -435 1400
rect -475 1350 -465 1370
rect -445 1350 -435 1370
rect -475 1320 -435 1350
rect -475 1300 -465 1320
rect -445 1300 -435 1320
rect -475 1270 -435 1300
rect -475 1250 -465 1270
rect -445 1250 -435 1270
rect -475 1220 -435 1250
rect 455 1420 495 1450
rect 455 1400 465 1420
rect 485 1400 495 1420
rect 455 1370 495 1400
rect 455 1350 465 1370
rect 485 1350 495 1370
rect 455 1320 495 1350
rect 455 1300 465 1320
rect 485 1300 495 1320
rect 455 1270 495 1300
rect 455 1250 465 1270
rect 485 1250 495 1270
rect 455 1235 495 1250
rect 510 1470 550 1485
rect 510 1450 520 1470
rect 540 1450 550 1470
rect 510 1420 550 1450
rect 510 1400 520 1420
rect 540 1400 550 1420
rect 510 1370 550 1400
rect 510 1350 520 1370
rect 540 1350 550 1370
rect 510 1320 550 1350
rect 510 1300 520 1320
rect 540 1300 550 1320
rect 510 1270 550 1300
rect 510 1250 520 1270
rect 540 1250 550 1270
rect 510 1235 550 1250
rect 565 1470 605 1485
rect 565 1450 575 1470
rect 595 1450 605 1470
rect 565 1420 605 1450
rect 565 1400 575 1420
rect 595 1400 605 1420
rect 565 1370 605 1400
rect 565 1350 575 1370
rect 595 1350 605 1370
rect 565 1320 605 1350
rect 565 1300 575 1320
rect 595 1300 605 1320
rect 565 1270 605 1300
rect 565 1250 575 1270
rect 595 1250 605 1270
rect 565 1235 605 1250
rect 620 1470 660 1485
rect 620 1450 630 1470
rect 650 1450 660 1470
rect 620 1420 660 1450
rect 620 1400 630 1420
rect 650 1400 660 1420
rect 620 1370 660 1400
rect 620 1350 630 1370
rect 650 1350 660 1370
rect 620 1320 660 1350
rect 620 1300 630 1320
rect 650 1300 660 1320
rect 620 1270 660 1300
rect 620 1250 630 1270
rect 650 1250 660 1270
rect 620 1235 660 1250
rect 675 1470 715 1485
rect 675 1450 685 1470
rect 705 1450 715 1470
rect 675 1420 715 1450
rect 675 1400 685 1420
rect 705 1400 715 1420
rect 675 1370 715 1400
rect 675 1350 685 1370
rect 705 1350 715 1370
rect 675 1320 715 1350
rect 675 1300 685 1320
rect 705 1300 715 1320
rect 675 1270 715 1300
rect 675 1250 685 1270
rect 705 1250 715 1270
rect 675 1235 715 1250
rect 730 1470 770 1485
rect 730 1450 740 1470
rect 760 1450 770 1470
rect 730 1420 770 1450
rect 730 1400 740 1420
rect 760 1400 770 1420
rect 730 1370 770 1400
rect 730 1350 740 1370
rect 760 1350 770 1370
rect 730 1320 770 1350
rect 730 1300 740 1320
rect 760 1300 770 1320
rect 730 1270 770 1300
rect 730 1250 740 1270
rect 760 1250 770 1270
rect 730 1235 770 1250
rect 785 1470 825 1485
rect 865 1470 905 1485
rect 785 1450 795 1470
rect 815 1450 825 1470
rect 865 1450 875 1470
rect 895 1450 905 1470
rect 785 1420 825 1450
rect 865 1420 905 1450
rect 785 1400 795 1420
rect 815 1400 825 1420
rect 865 1400 875 1420
rect 895 1400 905 1420
rect 785 1370 825 1400
rect 865 1370 905 1400
rect 785 1350 795 1370
rect 815 1350 825 1370
rect 865 1350 875 1370
rect 895 1350 905 1370
rect 785 1320 825 1350
rect 865 1320 905 1350
rect 785 1300 795 1320
rect 815 1300 825 1320
rect 865 1300 875 1320
rect 895 1300 905 1320
rect 785 1270 825 1300
rect 865 1270 905 1300
rect 785 1250 795 1270
rect 815 1250 825 1270
rect 865 1250 875 1270
rect 895 1250 905 1270
rect 785 1235 825 1250
rect 865 1235 905 1250
rect 920 1470 960 1485
rect 920 1450 930 1470
rect 950 1450 960 1470
rect 920 1420 960 1450
rect 920 1400 930 1420
rect 950 1400 960 1420
rect 920 1370 960 1400
rect 920 1350 930 1370
rect 950 1350 960 1370
rect 920 1320 960 1350
rect 920 1300 930 1320
rect 950 1300 960 1320
rect 920 1270 960 1300
rect 920 1250 930 1270
rect 950 1250 960 1270
rect 920 1235 960 1250
rect 975 1470 1015 1485
rect 975 1450 985 1470
rect 1005 1450 1015 1470
rect 975 1420 1015 1450
rect 975 1400 985 1420
rect 1005 1400 1015 1420
rect 975 1370 1015 1400
rect 975 1350 985 1370
rect 1005 1350 1015 1370
rect 975 1320 1015 1350
rect 975 1300 985 1320
rect 1005 1300 1015 1320
rect 975 1270 1015 1300
rect 975 1250 985 1270
rect 1005 1250 1015 1270
rect 975 1235 1015 1250
rect 1030 1470 1070 1485
rect 1030 1450 1040 1470
rect 1060 1450 1070 1470
rect 1030 1420 1070 1450
rect 1030 1400 1040 1420
rect 1060 1400 1070 1420
rect 1030 1370 1070 1400
rect 1030 1350 1040 1370
rect 1060 1350 1070 1370
rect 1030 1320 1070 1350
rect 1030 1300 1040 1320
rect 1060 1300 1070 1320
rect 1030 1270 1070 1300
rect 1030 1250 1040 1270
rect 1060 1250 1070 1270
rect 1030 1235 1070 1250
rect 1085 1470 1125 1485
rect 1085 1450 1095 1470
rect 1115 1450 1125 1470
rect 1085 1420 1125 1450
rect 1085 1400 1095 1420
rect 1115 1400 1125 1420
rect 1085 1370 1125 1400
rect 1085 1350 1095 1370
rect 1115 1350 1125 1370
rect 1085 1320 1125 1350
rect 1085 1300 1095 1320
rect 1115 1300 1125 1320
rect 1085 1270 1125 1300
rect 1085 1250 1095 1270
rect 1115 1250 1125 1270
rect 1085 1235 1125 1250
rect 1140 1470 1180 1485
rect 1140 1450 1150 1470
rect 1170 1450 1180 1470
rect 1140 1420 1180 1450
rect 1140 1400 1150 1420
rect 1170 1400 1180 1420
rect 1140 1370 1180 1400
rect 1140 1350 1150 1370
rect 1170 1350 1180 1370
rect 1140 1320 1180 1350
rect 1140 1300 1150 1320
rect 1170 1300 1180 1320
rect 1140 1270 1180 1300
rect 1140 1250 1150 1270
rect 1170 1250 1180 1270
rect 1140 1235 1180 1250
rect 1195 1470 1235 1485
rect 1195 1450 1205 1470
rect 1225 1450 1235 1470
rect 1195 1420 1235 1450
rect 1195 1400 1205 1420
rect 1225 1400 1235 1420
rect 1195 1370 1235 1400
rect 1195 1350 1205 1370
rect 1225 1350 1235 1370
rect 1195 1320 1235 1350
rect 1195 1300 1205 1320
rect 1225 1300 1235 1320
rect 1195 1270 1235 1300
rect 1195 1250 1205 1270
rect 1225 1250 1235 1270
rect 1195 1235 1235 1250
rect 2125 1420 2165 1435
rect 2125 1400 2135 1420
rect 2155 1400 2165 1420
rect 2125 1370 2165 1400
rect 2125 1350 2135 1370
rect 2155 1350 2165 1370
rect 2125 1320 2165 1350
rect 2125 1300 2135 1320
rect 2155 1300 2165 1320
rect 2125 1270 2165 1300
rect 2125 1250 2135 1270
rect 2155 1250 2165 1270
rect -475 1200 -465 1220
rect -445 1200 -435 1220
rect 2125 1220 2165 1250
rect -475 1170 -435 1200
rect 2125 1200 2135 1220
rect 2155 1200 2165 1220
rect -475 1150 -465 1170
rect -445 1150 -435 1170
rect -475 1120 -435 1150
rect -475 1100 -465 1120
rect -445 1100 -435 1120
rect -475 1070 -435 1100
rect -475 1050 -465 1070
rect -445 1050 -435 1070
rect -475 1020 -435 1050
rect -475 1000 -465 1020
rect -445 1000 -435 1020
rect -475 970 -435 1000
rect -475 950 -465 970
rect -445 950 -435 970
rect -475 920 -435 950
rect 2125 1170 2165 1200
rect 2125 1150 2135 1170
rect 2155 1150 2165 1170
rect 2125 1120 2165 1150
rect 2125 1100 2135 1120
rect 2155 1100 2165 1120
rect 2125 1070 2165 1100
rect 2125 1050 2135 1070
rect 2155 1050 2165 1070
rect 2125 1020 2165 1050
rect 2125 1000 2135 1020
rect 2155 1000 2165 1020
rect 2125 970 2165 1000
rect 2125 950 2135 970
rect 2155 950 2165 970
rect -475 900 -465 920
rect -445 900 -435 920
rect -475 870 -435 900
rect 2125 920 2165 950
rect 2125 900 2135 920
rect 2155 900 2165 920
rect -475 850 -465 870
rect -445 850 -435 870
rect -475 835 -435 850
rect 2125 870 2165 900
rect 2125 850 2135 870
rect 2155 850 2165 870
rect 2125 835 2165 850
rect 2180 1420 2220 1435
rect 2180 1400 2190 1420
rect 2210 1400 2220 1420
rect 2180 1370 2220 1400
rect 2180 1350 2190 1370
rect 2210 1350 2220 1370
rect 2180 1320 2220 1350
rect 2180 1300 2190 1320
rect 2210 1300 2220 1320
rect 2180 1270 2220 1300
rect 2180 1250 2190 1270
rect 2210 1250 2220 1270
rect 2180 1220 2220 1250
rect 2180 1200 2190 1220
rect 2210 1200 2220 1220
rect 2180 1170 2220 1200
rect 2180 1150 2190 1170
rect 2210 1150 2220 1170
rect 2180 1120 2220 1150
rect 2180 1100 2190 1120
rect 2210 1100 2220 1120
rect 2180 1070 2220 1100
rect 2180 1050 2190 1070
rect 2210 1050 2220 1070
rect 2180 1020 2220 1050
rect 2180 1000 2190 1020
rect 2210 1000 2220 1020
rect 2180 970 2220 1000
rect 2180 950 2190 970
rect 2210 950 2220 970
rect 2180 920 2220 950
rect 2180 900 2190 920
rect 2210 900 2220 920
rect 2180 870 2220 900
rect 2180 850 2190 870
rect 2210 850 2220 870
rect 2180 835 2220 850
rect 2235 1420 2275 1435
rect 2235 1400 2245 1420
rect 2265 1400 2275 1420
rect 2235 1370 2275 1400
rect 2235 1350 2245 1370
rect 2265 1350 2275 1370
rect 2235 1320 2275 1350
rect 2235 1300 2245 1320
rect 2265 1300 2275 1320
rect 2235 1270 2275 1300
rect 2235 1250 2245 1270
rect 2265 1250 2275 1270
rect 2235 1220 2275 1250
rect 2235 1200 2245 1220
rect 2265 1200 2275 1220
rect 2235 1170 2275 1200
rect 2235 1150 2245 1170
rect 2265 1150 2275 1170
rect 2235 1120 2275 1150
rect 2235 1100 2245 1120
rect 2265 1100 2275 1120
rect 2235 1070 2275 1100
rect 2235 1050 2245 1070
rect 2265 1050 2275 1070
rect 2235 1020 2275 1050
rect 2235 1000 2245 1020
rect 2265 1000 2275 1020
rect 2235 970 2275 1000
rect 2235 950 2245 970
rect 2265 950 2275 970
rect 2235 920 2275 950
rect 2235 900 2245 920
rect 2265 900 2275 920
rect 2235 870 2275 900
rect 2235 850 2245 870
rect 2265 850 2275 870
rect 2235 835 2275 850
rect 2290 1420 2330 1435
rect 2290 1400 2300 1420
rect 2320 1400 2330 1420
rect 2290 1370 2330 1400
rect 2290 1350 2300 1370
rect 2320 1350 2330 1370
rect 2290 1320 2330 1350
rect 2290 1300 2300 1320
rect 2320 1300 2330 1320
rect 2290 1270 2330 1300
rect 2290 1250 2300 1270
rect 2320 1250 2330 1270
rect 2290 1220 2330 1250
rect 2290 1200 2300 1220
rect 2320 1200 2330 1220
rect 2290 1170 2330 1200
rect 2290 1150 2300 1170
rect 2320 1150 2330 1170
rect 2290 1120 2330 1150
rect 2290 1100 2300 1120
rect 2320 1100 2330 1120
rect 2290 1070 2330 1100
rect 2290 1050 2300 1070
rect 2320 1050 2330 1070
rect 2290 1020 2330 1050
rect 2290 1000 2300 1020
rect 2320 1000 2330 1020
rect 2290 970 2330 1000
rect 2290 950 2300 970
rect 2320 950 2330 970
rect 2290 920 2330 950
rect 2290 900 2300 920
rect 2320 900 2330 920
rect 2290 870 2330 900
rect 2290 850 2300 870
rect 2320 850 2330 870
rect 2290 835 2330 850
rect 2345 1420 2385 1435
rect 2345 1400 2355 1420
rect 2375 1400 2385 1420
rect 2345 1370 2385 1400
rect 2345 1350 2355 1370
rect 2375 1350 2385 1370
rect 2345 1320 2385 1350
rect 2345 1300 2355 1320
rect 2375 1300 2385 1320
rect 2345 1270 2385 1300
rect 2345 1250 2355 1270
rect 2375 1250 2385 1270
rect 2345 1220 2385 1250
rect 2345 1200 2355 1220
rect 2375 1200 2385 1220
rect 2345 1170 2385 1200
rect 2345 1150 2355 1170
rect 2375 1150 2385 1170
rect 2345 1120 2385 1150
rect 2345 1100 2355 1120
rect 2375 1100 2385 1120
rect 2345 1070 2385 1100
rect 2345 1050 2355 1070
rect 2375 1050 2385 1070
rect 2345 1020 2385 1050
rect 2345 1000 2355 1020
rect 2375 1000 2385 1020
rect 2345 970 2385 1000
rect 2345 950 2355 970
rect 2375 950 2385 970
rect 2345 920 2385 950
rect 2345 900 2355 920
rect 2375 900 2385 920
rect 2345 870 2385 900
rect 2345 850 2355 870
rect 2375 850 2385 870
rect 2345 835 2385 850
rect 2400 1420 2440 1435
rect 2400 1400 2410 1420
rect 2430 1400 2440 1420
rect 2400 1370 2440 1400
rect 2400 1350 2410 1370
rect 2430 1350 2440 1370
rect 2400 1320 2440 1350
rect 2400 1300 2410 1320
rect 2430 1300 2440 1320
rect 2400 1270 2440 1300
rect 2400 1250 2410 1270
rect 2430 1250 2440 1270
rect 2400 1220 2440 1250
rect 2400 1200 2410 1220
rect 2430 1200 2440 1220
rect 2400 1170 2440 1200
rect 2400 1150 2410 1170
rect 2430 1150 2440 1170
rect 2400 1120 2440 1150
rect 2400 1100 2410 1120
rect 2430 1100 2440 1120
rect 2400 1070 2440 1100
rect 2400 1050 2410 1070
rect 2430 1050 2440 1070
rect 2400 1020 2440 1050
rect 2400 1000 2410 1020
rect 2430 1000 2440 1020
rect 2400 970 2440 1000
rect 2400 950 2410 970
rect 2430 950 2440 970
rect 2400 920 2440 950
rect 2400 900 2410 920
rect 2430 900 2440 920
rect 2400 870 2440 900
rect 2400 850 2410 870
rect 2430 850 2440 870
rect 2400 835 2440 850
rect 2455 1420 2495 1435
rect 2455 1400 2465 1420
rect 2485 1400 2495 1420
rect 2455 1370 2495 1400
rect 2455 1350 2465 1370
rect 2485 1350 2495 1370
rect 2455 1320 2495 1350
rect 2455 1300 2465 1320
rect 2485 1300 2495 1320
rect 2455 1270 2495 1300
rect 2455 1250 2465 1270
rect 2485 1250 2495 1270
rect 2455 1220 2495 1250
rect 2455 1200 2465 1220
rect 2485 1200 2495 1220
rect 2455 1170 2495 1200
rect 2455 1150 2465 1170
rect 2485 1150 2495 1170
rect 2455 1120 2495 1150
rect 2455 1100 2465 1120
rect 2485 1100 2495 1120
rect 2455 1070 2495 1100
rect 2455 1050 2465 1070
rect 2485 1050 2495 1070
rect 2455 1020 2495 1050
rect 2455 1000 2465 1020
rect 2485 1000 2495 1020
rect 2455 970 2495 1000
rect 2455 950 2465 970
rect 2485 950 2495 970
rect 2455 920 2495 950
rect 2455 900 2465 920
rect 2485 900 2495 920
rect 2455 870 2495 900
rect 2455 850 2465 870
rect 2485 850 2495 870
rect 2455 835 2495 850
rect 2510 1420 2550 1435
rect 2510 1400 2520 1420
rect 2540 1400 2550 1420
rect 2510 1370 2550 1400
rect 2510 1350 2520 1370
rect 2540 1350 2550 1370
rect 2510 1320 2550 1350
rect 2510 1300 2520 1320
rect 2540 1300 2550 1320
rect 2510 1270 2550 1300
rect 2510 1250 2520 1270
rect 2540 1250 2550 1270
rect 2510 1220 2550 1250
rect 2510 1200 2520 1220
rect 2540 1200 2550 1220
rect 2510 1170 2550 1200
rect 2510 1150 2520 1170
rect 2540 1150 2550 1170
rect 2510 1120 2550 1150
rect 2510 1100 2520 1120
rect 2540 1100 2550 1120
rect 2510 1070 2550 1100
rect 2510 1050 2520 1070
rect 2540 1050 2550 1070
rect 2510 1020 2550 1050
rect 2510 1000 2520 1020
rect 2540 1000 2550 1020
rect 2510 970 2550 1000
rect 2510 950 2520 970
rect 2540 950 2550 970
rect 2510 920 2550 950
rect 2510 900 2520 920
rect 2540 900 2550 920
rect 2510 870 2550 900
rect 2510 850 2520 870
rect 2540 850 2550 870
rect 2510 835 2550 850
rect 2565 1420 2605 1435
rect 2565 1400 2575 1420
rect 2595 1400 2605 1420
rect 2565 1370 2605 1400
rect 2565 1350 2575 1370
rect 2595 1350 2605 1370
rect 2565 1320 2605 1350
rect 2565 1300 2575 1320
rect 2595 1300 2605 1320
rect 2565 1270 2605 1300
rect 2565 1250 2575 1270
rect 2595 1250 2605 1270
rect 2565 1220 2605 1250
rect 2565 1200 2575 1220
rect 2595 1200 2605 1220
rect 2565 1170 2605 1200
rect 2565 1150 2575 1170
rect 2595 1150 2605 1170
rect 2565 1120 2605 1150
rect 2565 1100 2575 1120
rect 2595 1100 2605 1120
rect 2565 1070 2605 1100
rect 2565 1050 2575 1070
rect 2595 1050 2605 1070
rect 2565 1020 2605 1050
rect 2565 1000 2575 1020
rect 2595 1000 2605 1020
rect 2565 970 2605 1000
rect 2565 950 2575 970
rect 2595 950 2605 970
rect 2565 920 2605 950
rect 2565 900 2575 920
rect 2595 900 2605 920
rect 2565 870 2605 900
rect 2565 850 2575 870
rect 2595 850 2605 870
rect 2565 835 2605 850
rect 2620 1420 2660 1435
rect 2620 1400 2630 1420
rect 2650 1400 2660 1420
rect 2620 1370 2660 1400
rect 2620 1350 2630 1370
rect 2650 1350 2660 1370
rect 2620 1320 2660 1350
rect 2620 1300 2630 1320
rect 2650 1300 2660 1320
rect 2620 1270 2660 1300
rect 2620 1250 2630 1270
rect 2650 1250 2660 1270
rect 2620 1220 2660 1250
rect 2620 1200 2630 1220
rect 2650 1200 2660 1220
rect 2620 1170 2660 1200
rect 2620 1150 2630 1170
rect 2650 1150 2660 1170
rect 2620 1120 2660 1150
rect 2620 1100 2630 1120
rect 2650 1100 2660 1120
rect 2620 1070 2660 1100
rect 2620 1050 2630 1070
rect 2650 1050 2660 1070
rect 2620 1020 2660 1050
rect 2620 1000 2630 1020
rect 2650 1000 2660 1020
rect 2620 970 2660 1000
rect 2620 950 2630 970
rect 2650 950 2660 970
rect 2620 920 2660 950
rect 2620 900 2630 920
rect 2650 900 2660 920
rect 2620 870 2660 900
rect 2620 850 2630 870
rect 2650 850 2660 870
rect 2620 835 2660 850
rect 2675 1420 2715 1435
rect 2675 1400 2685 1420
rect 2705 1400 2715 1420
rect 2675 1370 2715 1400
rect 2675 1350 2685 1370
rect 2705 1350 2715 1370
rect 2675 1320 2715 1350
rect 2675 1300 2685 1320
rect 2705 1300 2715 1320
rect 2675 1270 2715 1300
rect 2675 1250 2685 1270
rect 2705 1250 2715 1270
rect 2675 1220 2715 1250
rect 2675 1200 2685 1220
rect 2705 1200 2715 1220
rect 2675 1170 2715 1200
rect 2675 1150 2685 1170
rect 2705 1150 2715 1170
rect 2675 1120 2715 1150
rect 2675 1100 2685 1120
rect 2705 1100 2715 1120
rect 2675 1070 2715 1100
rect 2675 1050 2685 1070
rect 2705 1050 2715 1070
rect 2675 1020 2715 1050
rect 2675 1000 2685 1020
rect 2705 1000 2715 1020
rect 2675 970 2715 1000
rect 2675 950 2685 970
rect 2705 950 2715 970
rect 2675 920 2715 950
rect 2675 900 2685 920
rect 2705 900 2715 920
rect 2675 870 2715 900
rect 2675 850 2685 870
rect 2705 850 2715 870
rect 2675 835 2715 850
rect 2730 1420 2770 1435
rect 2730 1400 2740 1420
rect 2760 1400 2770 1420
rect 2730 1370 2770 1400
rect 2730 1350 2740 1370
rect 2760 1350 2770 1370
rect 2730 1320 2770 1350
rect 2730 1300 2740 1320
rect 2760 1300 2770 1320
rect 2730 1270 2770 1300
rect 2730 1250 2740 1270
rect 2760 1250 2770 1270
rect 2730 1220 2770 1250
rect 2730 1200 2740 1220
rect 2760 1200 2770 1220
rect 2730 1170 2770 1200
rect 2730 1150 2740 1170
rect 2760 1150 2770 1170
rect 2730 1120 2770 1150
rect 2730 1100 2740 1120
rect 2760 1100 2770 1120
rect 2730 1070 2770 1100
rect 2730 1050 2740 1070
rect 2760 1050 2770 1070
rect 2730 1020 2770 1050
rect 2730 1000 2740 1020
rect 2760 1000 2770 1020
rect 2730 970 2770 1000
rect 2730 950 2740 970
rect 2760 950 2770 970
rect 2730 920 2770 950
rect 2730 900 2740 920
rect 2760 900 2770 920
rect 2730 870 2770 900
rect 2730 850 2740 870
rect 2760 850 2770 870
rect 2730 835 2770 850
rect 2785 1420 2825 1435
rect 2785 1400 2795 1420
rect 2815 1400 2825 1420
rect 2785 1370 2825 1400
rect 2785 1350 2795 1370
rect 2815 1350 2825 1370
rect 2785 1320 2825 1350
rect 2785 1300 2795 1320
rect 2815 1300 2825 1320
rect 2785 1270 2825 1300
rect 2785 1250 2795 1270
rect 2815 1250 2825 1270
rect 2785 1220 2825 1250
rect 2785 1200 2795 1220
rect 2815 1200 2825 1220
rect 2785 1170 2825 1200
rect 2785 1150 2795 1170
rect 2815 1150 2825 1170
rect 2785 1120 2825 1150
rect 2785 1100 2795 1120
rect 2815 1100 2825 1120
rect 2785 1070 2825 1100
rect 2785 1050 2795 1070
rect 2815 1050 2825 1070
rect 2785 1020 2825 1050
rect 2785 1000 2795 1020
rect 2815 1000 2825 1020
rect 2785 970 2825 1000
rect 2785 950 2795 970
rect 2815 950 2825 970
rect 2785 920 2825 950
rect 2785 900 2795 920
rect 2815 900 2825 920
rect 2785 870 2825 900
rect 2785 850 2795 870
rect 2815 850 2825 870
rect 2785 835 2825 850
rect -1135 605 -1095 620
rect -1135 585 -1125 605
rect -1105 585 -1095 605
rect -1135 555 -1095 585
rect -1135 535 -1125 555
rect -1105 535 -1095 555
rect -1135 505 -1095 535
rect -1135 485 -1125 505
rect -1105 485 -1095 505
rect -1135 455 -1095 485
rect -1135 435 -1125 455
rect -1105 435 -1095 455
rect -1135 420 -1095 435
rect -1080 605 -1040 620
rect -1080 585 -1070 605
rect -1050 585 -1040 605
rect -1080 555 -1040 585
rect -1080 535 -1070 555
rect -1050 535 -1040 555
rect -1080 505 -1040 535
rect -1080 485 -1070 505
rect -1050 485 -1040 505
rect -1080 455 -1040 485
rect -1080 435 -1070 455
rect -1050 435 -1040 455
rect -1080 420 -1040 435
rect -1025 605 -985 620
rect -1025 585 -1015 605
rect -995 585 -985 605
rect -1025 555 -985 585
rect -1025 535 -1015 555
rect -995 535 -985 555
rect -1025 505 -985 535
rect -1025 485 -1015 505
rect -995 485 -985 505
rect -1025 455 -985 485
rect -1025 435 -1015 455
rect -995 435 -985 455
rect -1025 420 -985 435
rect -970 605 -930 620
rect -970 585 -960 605
rect -940 585 -930 605
rect -970 555 -930 585
rect -970 535 -960 555
rect -940 535 -930 555
rect -970 505 -930 535
rect -970 485 -960 505
rect -940 485 -930 505
rect -970 455 -930 485
rect -970 435 -960 455
rect -940 435 -930 455
rect -970 420 -930 435
rect -915 605 -875 620
rect -915 585 -905 605
rect -885 585 -875 605
rect -915 555 -875 585
rect -915 535 -905 555
rect -885 535 -875 555
rect -915 505 -875 535
rect -915 485 -905 505
rect -885 485 -875 505
rect -915 455 -875 485
rect -915 435 -905 455
rect -885 435 -875 455
rect -915 420 -875 435
rect -860 605 -820 620
rect -860 585 -850 605
rect -830 585 -820 605
rect -860 555 -820 585
rect -860 535 -850 555
rect -830 535 -820 555
rect -860 505 -820 535
rect -860 485 -850 505
rect -830 485 -820 505
rect -860 455 -820 485
rect -860 435 -850 455
rect -830 435 -820 455
rect -860 420 -820 435
rect -805 605 -765 620
rect -805 585 -795 605
rect -775 585 -765 605
rect -805 555 -765 585
rect -805 535 -795 555
rect -775 535 -765 555
rect -805 505 -765 535
rect -805 485 -795 505
rect -775 485 -765 505
rect -805 455 -765 485
rect -805 435 -795 455
rect -775 435 -765 455
rect -805 420 -765 435
rect -750 605 -710 620
rect -750 585 -740 605
rect -720 585 -710 605
rect -750 555 -710 585
rect -750 535 -740 555
rect -720 535 -710 555
rect -750 505 -710 535
rect -750 485 -740 505
rect -720 485 -710 505
rect -750 455 -710 485
rect -750 435 -740 455
rect -720 435 -710 455
rect -750 420 -710 435
rect -695 605 -655 620
rect -695 585 -685 605
rect -665 585 -655 605
rect -695 555 -655 585
rect -695 535 -685 555
rect -665 535 -655 555
rect -695 505 -655 535
rect -695 485 -685 505
rect -665 485 -655 505
rect -695 455 -655 485
rect -695 435 -685 455
rect -665 435 -655 455
rect -695 420 -655 435
rect -640 605 -600 620
rect -640 585 -630 605
rect -610 585 -600 605
rect -640 555 -600 585
rect -640 535 -630 555
rect -610 535 -600 555
rect -640 505 -600 535
rect -640 485 -630 505
rect -610 485 -600 505
rect -640 455 -600 485
rect -640 435 -630 455
rect -610 435 -600 455
rect -640 420 -600 435
rect -585 605 -545 620
rect -585 585 -575 605
rect -555 585 -545 605
rect -585 555 -545 585
rect -585 535 -575 555
rect -555 535 -545 555
rect -585 505 -545 535
rect -585 485 -575 505
rect -555 485 -545 505
rect -585 455 -545 485
rect -585 435 -575 455
rect -555 435 -545 455
rect -585 420 -545 435
rect -530 605 -490 620
rect -530 585 -520 605
rect -500 585 -490 605
rect -530 555 -490 585
rect -530 535 -520 555
rect -500 535 -490 555
rect -530 505 -490 535
rect -530 485 -520 505
rect -500 485 -490 505
rect -530 455 -490 485
rect -530 435 -520 455
rect -500 435 -490 455
rect -530 420 -490 435
rect -475 605 -435 620
rect -475 585 -465 605
rect -445 585 -435 605
rect -475 555 -435 585
rect 2125 605 2165 620
rect 2125 585 2135 605
rect 2155 585 2165 605
rect -475 535 -465 555
rect -445 535 -435 555
rect -475 505 -435 535
rect 2125 555 2165 585
rect 2125 535 2135 555
rect 2155 535 2165 555
rect -475 485 -465 505
rect -445 485 -435 505
rect -475 455 -435 485
rect 2125 505 2165 535
rect 2125 485 2135 505
rect 2155 485 2165 505
rect 2125 455 2165 485
rect -475 435 -465 455
rect -445 435 -435 455
rect -475 420 -435 435
rect 2125 435 2135 455
rect 2155 435 2165 455
rect 2125 420 2165 435
rect 2180 605 2220 620
rect 2180 585 2190 605
rect 2210 585 2220 605
rect 2180 555 2220 585
rect 2180 535 2190 555
rect 2210 535 2220 555
rect 2180 505 2220 535
rect 2180 485 2190 505
rect 2210 485 2220 505
rect 2180 455 2220 485
rect 2180 435 2190 455
rect 2210 435 2220 455
rect 2180 420 2220 435
rect 2235 605 2275 620
rect 2235 585 2245 605
rect 2265 585 2275 605
rect 2235 555 2275 585
rect 2235 535 2245 555
rect 2265 535 2275 555
rect 2235 505 2275 535
rect 2235 485 2245 505
rect 2265 485 2275 505
rect 2235 455 2275 485
rect 2235 435 2245 455
rect 2265 435 2275 455
rect 2235 420 2275 435
rect 2290 605 2330 620
rect 2290 585 2300 605
rect 2320 585 2330 605
rect 2290 555 2330 585
rect 2290 535 2300 555
rect 2320 535 2330 555
rect 2290 505 2330 535
rect 2290 485 2300 505
rect 2320 485 2330 505
rect 2290 455 2330 485
rect 2290 435 2300 455
rect 2320 435 2330 455
rect 2290 420 2330 435
rect 2345 605 2385 620
rect 2345 585 2355 605
rect 2375 585 2385 605
rect 2345 555 2385 585
rect 2345 535 2355 555
rect 2375 535 2385 555
rect 2345 505 2385 535
rect 2345 485 2355 505
rect 2375 485 2385 505
rect 2345 455 2385 485
rect 2345 435 2355 455
rect 2375 435 2385 455
rect 2345 420 2385 435
rect 2400 605 2440 620
rect 2400 585 2410 605
rect 2430 585 2440 605
rect 2400 555 2440 585
rect 2400 535 2410 555
rect 2430 535 2440 555
rect 2400 505 2440 535
rect 2400 485 2410 505
rect 2430 485 2440 505
rect 2400 455 2440 485
rect 2400 435 2410 455
rect 2430 435 2440 455
rect 2400 420 2440 435
rect 2455 605 2495 620
rect 2455 585 2465 605
rect 2485 585 2495 605
rect 2455 555 2495 585
rect 2455 535 2465 555
rect 2485 535 2495 555
rect 2455 505 2495 535
rect 2455 485 2465 505
rect 2485 485 2495 505
rect 2455 455 2495 485
rect 2455 435 2465 455
rect 2485 435 2495 455
rect 2455 420 2495 435
rect 2510 605 2550 620
rect 2510 585 2520 605
rect 2540 585 2550 605
rect 2510 555 2550 585
rect 2510 535 2520 555
rect 2540 535 2550 555
rect 2510 505 2550 535
rect 2510 485 2520 505
rect 2540 485 2550 505
rect 2510 455 2550 485
rect 2510 435 2520 455
rect 2540 435 2550 455
rect 2510 420 2550 435
rect 2565 605 2605 620
rect 2565 585 2575 605
rect 2595 585 2605 605
rect 2565 555 2605 585
rect 2565 535 2575 555
rect 2595 535 2605 555
rect 2565 505 2605 535
rect 2565 485 2575 505
rect 2595 485 2605 505
rect 2565 455 2605 485
rect 2565 435 2575 455
rect 2595 435 2605 455
rect 2565 420 2605 435
rect 2620 605 2660 620
rect 2620 585 2630 605
rect 2650 585 2660 605
rect 2620 555 2660 585
rect 2620 535 2630 555
rect 2650 535 2660 555
rect 2620 505 2660 535
rect 2620 485 2630 505
rect 2650 485 2660 505
rect 2620 455 2660 485
rect 2620 435 2630 455
rect 2650 435 2660 455
rect 2620 420 2660 435
rect 2675 605 2715 620
rect 2675 585 2685 605
rect 2705 585 2715 605
rect 2675 555 2715 585
rect 2675 535 2685 555
rect 2705 535 2715 555
rect 2675 505 2715 535
rect 2675 485 2685 505
rect 2705 485 2715 505
rect 2675 455 2715 485
rect 2675 435 2685 455
rect 2705 435 2715 455
rect 2675 420 2715 435
rect 2730 605 2770 620
rect 2730 585 2740 605
rect 2760 585 2770 605
rect 2730 555 2770 585
rect 2730 535 2740 555
rect 2760 535 2770 555
rect 2730 505 2770 535
rect 2730 485 2740 505
rect 2760 485 2770 505
rect 2730 455 2770 485
rect 2730 435 2740 455
rect 2760 435 2770 455
rect 2730 420 2770 435
rect 2785 605 2825 620
rect 2785 585 2795 605
rect 2815 585 2825 605
rect 2785 555 2825 585
rect 2785 535 2795 555
rect 2815 535 2825 555
rect 2785 505 2825 535
rect 2785 485 2795 505
rect 2815 485 2825 505
rect 2785 455 2825 485
rect 2785 435 2795 455
rect 2815 435 2825 455
rect 2785 420 2825 435
<< ndiffc >>
rect -95 815 -75 835
rect -95 765 -75 785
rect -95 715 -75 735
rect -40 815 -20 835
rect -40 765 -20 785
rect -40 715 -20 735
rect 15 815 35 835
rect 15 765 35 785
rect 15 715 35 735
rect 70 815 90 835
rect 70 765 90 785
rect 70 715 90 735
rect 125 815 145 835
rect 125 765 145 785
rect 125 715 145 735
rect 180 815 200 835
rect 180 765 200 785
rect 180 715 200 735
rect 235 815 255 835
rect 235 765 255 785
rect 235 715 255 735
rect 290 815 310 835
rect 290 765 310 785
rect 290 715 310 735
rect 345 815 365 835
rect 345 765 365 785
rect 345 715 365 735
rect 400 815 420 835
rect 400 765 420 785
rect 400 715 420 735
rect 455 815 475 835
rect 455 765 475 785
rect 455 715 475 735
rect 510 815 530 835
rect 510 765 530 785
rect 510 715 530 735
rect 565 815 585 835
rect 565 765 585 785
rect 565 715 585 735
rect 725 840 745 860
rect 725 790 745 810
rect 725 740 745 760
rect 725 690 745 710
rect 725 640 745 660
rect 780 840 800 860
rect 780 790 800 810
rect 780 740 800 760
rect 780 690 800 710
rect 780 640 800 660
rect 835 840 855 860
rect 835 790 855 810
rect 835 740 855 760
rect 835 690 855 710
rect 835 640 855 660
rect 890 840 910 860
rect 890 790 910 810
rect 890 740 910 760
rect 890 690 910 710
rect 890 640 910 660
rect 945 840 965 860
rect 945 790 965 810
rect 945 740 965 760
rect 945 690 965 710
rect 1105 815 1125 835
rect 1105 765 1125 785
rect 1105 715 1125 735
rect 1160 815 1180 835
rect 1160 765 1180 785
rect 1160 715 1180 735
rect 1215 815 1235 835
rect 1215 765 1235 785
rect 1215 715 1235 735
rect 1270 815 1290 835
rect 1270 765 1290 785
rect 1270 715 1290 735
rect 1325 815 1345 835
rect 1325 765 1345 785
rect 1325 715 1345 735
rect 1380 815 1400 835
rect 1380 765 1400 785
rect 1380 715 1400 735
rect 1435 815 1455 835
rect 1435 765 1455 785
rect 1435 715 1455 735
rect 1490 815 1510 835
rect 1490 765 1510 785
rect 1490 715 1510 735
rect 1545 815 1565 835
rect 1545 765 1565 785
rect 1545 715 1565 735
rect 1600 815 1620 835
rect 1600 765 1620 785
rect 1600 715 1620 735
rect 1655 815 1675 835
rect 1655 765 1675 785
rect 1655 715 1675 735
rect 1710 815 1730 835
rect 1710 765 1730 785
rect 1710 715 1730 735
rect 1765 815 1785 835
rect 1765 765 1785 785
rect 1765 715 1785 735
rect 945 640 965 660
rect -95 420 -75 440
rect -95 370 -75 390
rect -95 320 -75 340
rect -40 420 -20 440
rect -40 370 -20 390
rect -40 320 -20 340
rect 15 420 35 440
rect 15 370 35 390
rect 15 320 35 340
rect 70 420 90 440
rect 70 370 90 390
rect 70 320 90 340
rect 125 420 145 440
rect 125 370 145 390
rect 125 320 145 340
rect 180 420 200 440
rect 180 370 200 390
rect 180 320 200 340
rect 235 420 255 440
rect 235 370 255 390
rect 235 320 255 340
rect 290 420 310 440
rect 290 370 310 390
rect 290 320 310 340
rect 345 420 365 440
rect 345 370 365 390
rect 345 320 365 340
rect 400 420 420 440
rect 400 370 420 390
rect 400 320 420 340
rect 455 420 475 440
rect 455 370 475 390
rect 455 320 475 340
rect 510 420 530 440
rect 510 370 530 390
rect 510 320 530 340
rect 565 420 585 440
rect 565 370 585 390
rect 565 320 585 340
rect 725 420 745 440
rect 725 370 745 390
rect 725 320 745 340
rect 780 420 800 440
rect 780 370 800 390
rect 780 320 800 340
rect 835 420 855 440
rect 835 370 855 390
rect 835 320 855 340
rect 890 420 910 440
rect 890 370 910 390
rect 890 320 910 340
rect 945 420 965 440
rect 945 370 965 390
rect 945 320 965 340
rect 1105 420 1125 440
rect 1105 370 1125 390
rect 1105 320 1125 340
rect 1160 420 1180 440
rect 1160 370 1180 390
rect 1160 320 1180 340
rect 1215 420 1235 440
rect 1215 370 1235 390
rect 1215 320 1235 340
rect 1270 420 1290 440
rect 1270 370 1290 390
rect 1270 320 1290 340
rect 1325 420 1345 440
rect 1325 370 1345 390
rect 1325 320 1345 340
rect 1380 420 1400 440
rect 1380 370 1400 390
rect 1380 320 1400 340
rect 1435 420 1455 440
rect 1435 370 1455 390
rect 1435 320 1455 340
rect 1490 420 1510 440
rect 1490 370 1510 390
rect 1490 320 1510 340
rect 1545 420 1565 440
rect 1545 370 1565 390
rect 1545 320 1565 340
rect 1600 420 1620 440
rect 1600 370 1620 390
rect 1600 320 1620 340
rect 1655 420 1675 440
rect 1655 370 1675 390
rect 1655 320 1675 340
rect 1710 420 1730 440
rect 1710 370 1730 390
rect 1710 320 1730 340
rect 1765 420 1785 440
rect 1765 370 1785 390
rect 1765 320 1785 340
rect -1125 195 -1105 215
rect -1125 145 -1105 165
rect -1125 95 -1105 115
rect -1125 45 -1105 65
rect -1125 -5 -1105 15
rect -1125 -55 -1105 -35
rect -1070 195 -1050 215
rect -1070 145 -1050 165
rect -1070 95 -1050 115
rect -1070 45 -1050 65
rect -1070 -5 -1050 15
rect -1070 -55 -1050 -35
rect -1015 195 -995 215
rect -1015 145 -995 165
rect -1015 95 -995 115
rect -1015 45 -995 65
rect -1015 -5 -995 15
rect -1015 -55 -995 -35
rect -960 195 -940 215
rect -960 145 -940 165
rect -960 95 -940 115
rect -960 45 -940 65
rect -960 -5 -940 15
rect -960 -55 -940 -35
rect -905 195 -885 215
rect -905 145 -885 165
rect -905 95 -885 115
rect -905 45 -885 65
rect -905 -5 -885 15
rect -905 -55 -885 -35
rect -850 195 -830 215
rect -850 145 -830 165
rect -850 95 -830 115
rect -850 45 -830 65
rect -850 -5 -830 15
rect -850 -55 -830 -35
rect -795 195 -775 215
rect -795 145 -775 165
rect -795 95 -775 115
rect -795 45 -775 65
rect -795 -5 -775 15
rect -795 -55 -775 -35
rect -740 195 -720 215
rect -740 145 -720 165
rect -740 95 -720 115
rect -740 45 -720 65
rect -740 -5 -720 15
rect -740 -55 -720 -35
rect -685 195 -665 215
rect -685 145 -665 165
rect -685 95 -665 115
rect -685 45 -665 65
rect -685 -5 -665 15
rect -685 -55 -665 -35
rect -630 195 -610 215
rect -630 145 -610 165
rect -630 95 -610 115
rect -630 45 -610 65
rect -630 -5 -610 15
rect -630 -55 -610 -35
rect -575 195 -555 215
rect -575 145 -555 165
rect -575 95 -555 115
rect -575 45 -555 65
rect -575 -5 -555 15
rect -575 -55 -555 -35
rect -520 195 -500 215
rect -520 145 -500 165
rect -520 95 -500 115
rect -520 45 -500 65
rect -520 -5 -500 15
rect -520 -55 -500 -35
rect -465 195 -445 215
rect -465 145 -445 165
rect -465 95 -445 115
rect -465 45 -445 65
rect 2135 195 2155 215
rect 2135 145 2155 165
rect 2135 95 2155 115
rect 2135 45 2155 65
rect -465 -5 -445 15
rect 2135 -5 2155 15
rect -465 -55 -445 -35
rect 725 -75 745 -55
rect 725 -125 745 -105
rect 725 -175 745 -155
rect 725 -225 745 -205
rect 725 -275 745 -255
rect 780 -75 800 -55
rect 780 -125 800 -105
rect 780 -175 800 -155
rect 780 -225 800 -205
rect 780 -275 800 -255
rect 835 -75 855 -55
rect 835 -125 855 -105
rect 835 -175 855 -155
rect 835 -225 855 -205
rect 835 -275 855 -255
rect 890 -75 910 -55
rect 890 -125 910 -105
rect 890 -175 910 -155
rect 890 -225 910 -205
rect 890 -275 910 -255
rect 945 -75 965 -55
rect 2135 -55 2155 -35
rect 2190 195 2210 215
rect 2190 145 2210 165
rect 2190 95 2210 115
rect 2190 45 2210 65
rect 2190 -5 2210 15
rect 2190 -55 2210 -35
rect 2245 195 2265 215
rect 2245 145 2265 165
rect 2245 95 2265 115
rect 2245 45 2265 65
rect 2245 -5 2265 15
rect 2245 -55 2265 -35
rect 2300 195 2320 215
rect 2300 145 2320 165
rect 2300 95 2320 115
rect 2300 45 2320 65
rect 2300 -5 2320 15
rect 2300 -55 2320 -35
rect 2355 195 2375 215
rect 2355 145 2375 165
rect 2355 95 2375 115
rect 2355 45 2375 65
rect 2355 -5 2375 15
rect 2355 -55 2375 -35
rect 2410 195 2430 215
rect 2410 145 2430 165
rect 2410 95 2430 115
rect 2410 45 2430 65
rect 2410 -5 2430 15
rect 2410 -55 2430 -35
rect 2465 195 2485 215
rect 2465 145 2485 165
rect 2465 95 2485 115
rect 2465 45 2485 65
rect 2465 -5 2485 15
rect 2465 -55 2485 -35
rect 2520 195 2540 215
rect 2520 145 2540 165
rect 2520 95 2540 115
rect 2520 45 2540 65
rect 2520 -5 2540 15
rect 2520 -55 2540 -35
rect 2575 195 2595 215
rect 2575 145 2595 165
rect 2575 95 2595 115
rect 2575 45 2595 65
rect 2575 -5 2595 15
rect 2575 -55 2595 -35
rect 2630 195 2650 215
rect 2630 145 2650 165
rect 2630 95 2650 115
rect 2630 45 2650 65
rect 2630 -5 2650 15
rect 2630 -55 2650 -35
rect 2685 195 2705 215
rect 2685 145 2705 165
rect 2685 95 2705 115
rect 2685 45 2705 65
rect 2685 -5 2705 15
rect 2685 -55 2705 -35
rect 2740 195 2760 215
rect 2740 145 2760 165
rect 2740 95 2760 115
rect 2740 45 2760 65
rect 2740 -5 2760 15
rect 2740 -55 2760 -35
rect 2795 195 2815 215
rect 2795 145 2815 165
rect 2795 95 2815 115
rect 2795 45 2815 65
rect 2795 -5 2815 15
rect 2795 -55 2815 -35
rect 945 -125 965 -105
rect 945 -175 965 -155
rect 945 -225 965 -205
rect 945 -275 965 -255
rect -1015 -390 -995 -370
rect -1015 -440 -995 -420
rect -1015 -490 -995 -470
rect -1015 -540 -995 -520
rect -1015 -590 -995 -570
rect -1015 -640 -995 -620
rect -1015 -690 -995 -670
rect -1015 -740 -995 -720
rect -1015 -790 -995 -770
rect -1015 -840 -995 -820
rect -1015 -890 -995 -870
rect -1015 -940 -995 -920
rect -1015 -990 -995 -970
rect -1015 -1040 -995 -1020
rect -915 -390 -895 -370
rect -915 -440 -895 -420
rect -915 -490 -895 -470
rect -915 -540 -895 -520
rect -915 -590 -895 -570
rect -915 -640 -895 -620
rect -915 -690 -895 -670
rect -915 -740 -895 -720
rect -915 -790 -895 -770
rect -915 -840 -895 -820
rect -915 -890 -895 -870
rect -915 -940 -895 -920
rect -915 -990 -895 -970
rect -915 -1040 -895 -1020
rect -815 -390 -795 -370
rect -815 -440 -795 -420
rect -815 -490 -795 -470
rect -815 -540 -795 -520
rect -815 -590 -795 -570
rect -815 -640 -795 -620
rect -815 -690 -795 -670
rect -815 -740 -795 -720
rect -815 -790 -795 -770
rect -815 -840 -795 -820
rect -815 -890 -795 -870
rect -815 -940 -795 -920
rect -815 -990 -795 -970
rect -815 -1040 -795 -1020
rect -715 -390 -695 -370
rect -715 -440 -695 -420
rect -715 -490 -695 -470
rect -715 -540 -695 -520
rect -715 -590 -695 -570
rect -715 -640 -695 -620
rect -715 -690 -695 -670
rect -715 -740 -695 -720
rect -715 -790 -695 -770
rect -715 -840 -695 -820
rect -715 -890 -695 -870
rect -715 -940 -695 -920
rect -715 -990 -695 -970
rect -715 -1040 -695 -1020
rect -615 -390 -595 -370
rect -615 -440 -595 -420
rect -615 -490 -595 -470
rect -615 -540 -595 -520
rect -615 -590 -595 -570
rect -615 -640 -595 -620
rect -615 -690 -595 -670
rect -615 -740 -595 -720
rect -615 -790 -595 -770
rect -615 -840 -595 -820
rect -615 -890 -595 -870
rect -615 -940 -595 -920
rect -615 -990 -595 -970
rect -615 -1040 -595 -1020
rect -515 -390 -495 -370
rect -515 -440 -495 -420
rect -515 -490 -495 -470
rect -515 -540 -495 -520
rect -515 -590 -495 -570
rect -515 -640 -495 -620
rect -515 -690 -495 -670
rect -515 -740 -495 -720
rect -515 -790 -495 -770
rect -515 -840 -495 -820
rect -515 -890 -495 -870
rect -515 -940 -495 -920
rect -515 -990 -495 -970
rect -515 -1040 -495 -1020
rect -415 -390 -395 -370
rect -415 -440 -395 -420
rect -415 -490 -395 -470
rect 2085 -390 2105 -370
rect 2085 -440 2105 -420
rect 2085 -490 2105 -470
rect -415 -540 -395 -520
rect -415 -590 -395 -570
rect -415 -640 -395 -620
rect -415 -690 -395 -670
rect -415 -740 -395 -720
rect -415 -790 -395 -770
rect 285 -570 305 -550
rect 285 -620 305 -600
rect 285 -670 305 -650
rect 285 -720 305 -700
rect 285 -770 305 -750
rect 340 -570 360 -550
rect 340 -620 360 -600
rect 340 -670 360 -650
rect 340 -720 360 -700
rect 340 -770 360 -750
rect 395 -570 415 -550
rect 395 -620 415 -600
rect 395 -670 415 -650
rect 395 -720 415 -700
rect 395 -770 415 -750
rect 450 -570 470 -550
rect 450 -620 470 -600
rect 450 -670 470 -650
rect 450 -720 470 -700
rect 450 -770 470 -750
rect 505 -570 525 -550
rect 505 -620 525 -600
rect 505 -670 525 -650
rect 505 -720 525 -700
rect 505 -770 525 -750
rect 560 -570 580 -550
rect 560 -620 580 -600
rect 560 -670 580 -650
rect 560 -720 580 -700
rect 560 -770 580 -750
rect 615 -570 635 -550
rect 615 -620 635 -600
rect 615 -670 635 -650
rect 615 -720 635 -700
rect 615 -770 635 -750
rect 670 -570 690 -550
rect 670 -620 690 -600
rect 670 -670 690 -650
rect 670 -720 690 -700
rect 670 -770 690 -750
rect 725 -570 745 -550
rect 725 -620 745 -600
rect 725 -670 745 -650
rect 725 -720 745 -700
rect 725 -770 745 -750
rect 780 -570 800 -550
rect 780 -620 800 -600
rect 780 -670 800 -650
rect 780 -720 800 -700
rect 780 -770 800 -750
rect 835 -570 855 -550
rect 835 -620 855 -600
rect 835 -670 855 -650
rect 835 -720 855 -700
rect 835 -770 855 -750
rect 890 -570 910 -550
rect 890 -620 910 -600
rect 890 -670 910 -650
rect 890 -720 910 -700
rect 890 -770 910 -750
rect 945 -570 965 -550
rect 945 -620 965 -600
rect 945 -670 965 -650
rect 945 -720 965 -700
rect 945 -770 965 -750
rect 1000 -570 1020 -550
rect 1000 -620 1020 -600
rect 1000 -670 1020 -650
rect 1000 -720 1020 -700
rect 1000 -770 1020 -750
rect 1055 -570 1075 -550
rect 1055 -620 1075 -600
rect 1055 -670 1075 -650
rect 1055 -720 1075 -700
rect 1055 -770 1075 -750
rect 1110 -570 1130 -550
rect 1110 -620 1130 -600
rect 1110 -670 1130 -650
rect 1110 -720 1130 -700
rect 1110 -770 1130 -750
rect 1165 -570 1185 -550
rect 1165 -620 1185 -600
rect 1165 -670 1185 -650
rect 1165 -720 1185 -700
rect 1165 -770 1185 -750
rect 1220 -570 1240 -550
rect 1220 -620 1240 -600
rect 1220 -670 1240 -650
rect 1220 -720 1240 -700
rect 1220 -770 1240 -750
rect 1275 -570 1295 -550
rect 1275 -620 1295 -600
rect 1275 -670 1295 -650
rect 1275 -720 1295 -700
rect 1275 -770 1295 -750
rect 1330 -570 1350 -550
rect 1330 -620 1350 -600
rect 1330 -670 1350 -650
rect 1330 -720 1350 -700
rect 1330 -770 1350 -750
rect 1385 -570 1405 -550
rect 1385 -620 1405 -600
rect 1385 -670 1405 -650
rect 1385 -720 1405 -700
rect 1385 -770 1405 -750
rect 1440 -570 1460 -550
rect 1440 -620 1460 -600
rect 1440 -670 1460 -650
rect 1440 -720 1460 -700
rect 1440 -770 1460 -750
rect 2085 -540 2105 -520
rect 2085 -590 2105 -570
rect 2085 -640 2105 -620
rect 2085 -690 2105 -670
rect 2085 -740 2105 -720
rect 2085 -790 2105 -770
rect -415 -840 -395 -820
rect 2085 -840 2105 -820
rect -415 -890 -395 -870
rect 2085 -890 2105 -870
rect -415 -940 -395 -920
rect 2085 -940 2105 -920
rect -415 -990 -395 -970
rect -415 -1040 -395 -1020
rect 505 -985 525 -965
rect 505 -1035 525 -1015
rect 505 -1085 525 -1065
rect 560 -985 580 -965
rect 560 -1035 580 -1015
rect 560 -1085 580 -1065
rect 615 -985 635 -965
rect 615 -1035 635 -1015
rect 615 -1085 635 -1065
rect 670 -985 690 -965
rect 670 -1035 690 -1015
rect 670 -1085 690 -1065
rect 725 -985 745 -965
rect 725 -1035 745 -1015
rect 725 -1085 745 -1065
rect 780 -985 800 -965
rect 780 -1035 800 -1015
rect 780 -1085 800 -1065
rect 835 -985 855 -965
rect 835 -1035 855 -1015
rect 835 -1085 855 -1065
rect 970 -985 990 -965
rect 970 -1035 990 -1015
rect 970 -1085 990 -1065
rect 1310 -985 1330 -965
rect 1310 -1035 1330 -1015
rect 2085 -990 2105 -970
rect 2085 -1040 2105 -1020
rect 2185 -390 2205 -370
rect 2185 -440 2205 -420
rect 2185 -490 2205 -470
rect 2185 -540 2205 -520
rect 2185 -590 2205 -570
rect 2185 -640 2205 -620
rect 2185 -690 2205 -670
rect 2185 -740 2205 -720
rect 2185 -790 2205 -770
rect 2185 -840 2205 -820
rect 2185 -890 2205 -870
rect 2185 -940 2205 -920
rect 2185 -990 2205 -970
rect 2185 -1040 2205 -1020
rect 2285 -390 2305 -370
rect 2285 -440 2305 -420
rect 2285 -490 2305 -470
rect 2285 -540 2305 -520
rect 2285 -590 2305 -570
rect 2285 -640 2305 -620
rect 2285 -690 2305 -670
rect 2285 -740 2305 -720
rect 2285 -790 2305 -770
rect 2285 -840 2305 -820
rect 2285 -890 2305 -870
rect 2285 -940 2305 -920
rect 2285 -990 2305 -970
rect 2285 -1040 2305 -1020
rect 2385 -390 2405 -370
rect 2385 -440 2405 -420
rect 2385 -490 2405 -470
rect 2385 -540 2405 -520
rect 2385 -590 2405 -570
rect 2385 -640 2405 -620
rect 2385 -690 2405 -670
rect 2385 -740 2405 -720
rect 2385 -790 2405 -770
rect 2385 -840 2405 -820
rect 2385 -890 2405 -870
rect 2385 -940 2405 -920
rect 2385 -990 2405 -970
rect 2385 -1040 2405 -1020
rect 2485 -390 2505 -370
rect 2485 -440 2505 -420
rect 2485 -490 2505 -470
rect 2485 -540 2505 -520
rect 2485 -590 2505 -570
rect 2485 -640 2505 -620
rect 2485 -690 2505 -670
rect 2485 -740 2505 -720
rect 2485 -790 2505 -770
rect 2485 -840 2505 -820
rect 2485 -890 2505 -870
rect 2485 -940 2505 -920
rect 2485 -990 2505 -970
rect 2485 -1040 2505 -1020
rect 2585 -390 2605 -370
rect 2585 -440 2605 -420
rect 2585 -490 2605 -470
rect 2585 -540 2605 -520
rect 2585 -590 2605 -570
rect 2585 -640 2605 -620
rect 2585 -690 2605 -670
rect 2585 -740 2605 -720
rect 2585 -790 2605 -770
rect 2585 -840 2605 -820
rect 2585 -890 2605 -870
rect 2585 -940 2605 -920
rect 2585 -990 2605 -970
rect 2585 -1040 2605 -1020
rect 2685 -390 2705 -370
rect 2685 -440 2705 -420
rect 2685 -490 2705 -470
rect 2685 -540 2705 -520
rect 2685 -590 2705 -570
rect 2685 -640 2705 -620
rect 2685 -690 2705 -670
rect 2685 -740 2705 -720
rect 2685 -790 2705 -770
rect 2685 -840 2705 -820
rect 2685 -890 2705 -870
rect 2685 -940 2705 -920
rect 2685 -990 2705 -970
rect 2685 -1040 2705 -1020
rect 1310 -1085 1330 -1065
<< pdiffc >>
rect 40 2640 60 2660
rect 40 2590 60 2610
rect 40 2540 60 2560
rect 40 2490 60 2510
rect 40 2440 60 2460
rect 40 2390 60 2410
rect 40 2340 60 2360
rect 100 2640 120 2660
rect 100 2590 120 2610
rect 100 2540 120 2560
rect 100 2490 120 2510
rect 100 2440 120 2460
rect 100 2390 120 2410
rect 100 2340 120 2360
rect 160 2640 180 2660
rect 160 2590 180 2610
rect 160 2540 180 2560
rect 160 2490 180 2510
rect 160 2440 180 2460
rect 160 2390 180 2410
rect 160 2340 180 2360
rect 220 2640 240 2660
rect 220 2590 240 2610
rect 980 2640 1000 2660
rect 980 2590 1000 2610
rect 220 2540 240 2560
rect 980 2540 1000 2560
rect 220 2490 240 2510
rect 220 2440 240 2460
rect 220 2390 240 2410
rect 220 2340 240 2360
rect 510 2340 530 2360
rect 570 2340 590 2360
rect 630 2340 650 2360
rect 690 2340 710 2360
rect 980 2490 1000 2510
rect 980 2440 1000 2460
rect 980 2390 1000 2410
rect 980 2340 1000 2360
rect 1040 2640 1060 2660
rect 1040 2590 1060 2610
rect 1040 2540 1060 2560
rect 1040 2490 1060 2510
rect 1040 2440 1060 2460
rect 1040 2390 1060 2410
rect 1040 2340 1060 2360
rect 1100 2640 1120 2660
rect 1100 2590 1120 2610
rect 1100 2540 1120 2560
rect 1100 2490 1120 2510
rect 1100 2440 1120 2460
rect 1100 2390 1120 2410
rect 1100 2340 1120 2360
rect 1160 2640 1180 2660
rect 1160 2590 1180 2610
rect 1160 2540 1180 2560
rect 1160 2490 1180 2510
rect 1160 2440 1180 2460
rect 1160 2390 1180 2410
rect 1160 2340 1180 2360
rect 1448 2640 1468 2660
rect 1448 2590 1468 2610
rect 1448 2540 1468 2560
rect 1448 2490 1468 2510
rect 1448 2440 1468 2460
rect 1448 2390 1468 2410
rect 1448 2340 1468 2360
rect 1508 2640 1528 2660
rect 1508 2590 1528 2610
rect 1508 2540 1528 2560
rect 1508 2490 1528 2510
rect 1508 2440 1528 2460
rect 1508 2390 1528 2410
rect 1508 2340 1528 2360
rect 1568 2640 1588 2660
rect 1568 2590 1588 2610
rect 1568 2540 1588 2560
rect 1568 2490 1588 2510
rect 1568 2440 1588 2460
rect 1568 2390 1588 2410
rect 1568 2340 1588 2360
rect 1628 2640 1648 2660
rect 1628 2590 1648 2610
rect 1628 2540 1648 2560
rect 1628 2490 1648 2510
rect 1628 2440 1648 2460
rect 1628 2390 1648 2410
rect 1628 2340 1648 2360
rect -1155 2065 -1135 2085
rect -1155 2015 -1135 2035
rect -1155 1965 -1135 1985
rect -1155 1915 -1135 1935
rect -1155 1865 -1135 1885
rect -1155 1815 -1135 1835
rect -1155 1765 -1135 1785
rect -1095 2065 -1075 2085
rect -1095 2015 -1075 2035
rect -1095 1965 -1075 1985
rect -1095 1915 -1075 1935
rect -1095 1865 -1075 1885
rect -1095 1815 -1075 1835
rect -1095 1765 -1075 1785
rect -1035 2065 -1015 2085
rect -1035 2015 -1015 2035
rect -1035 1965 -1015 1985
rect -1035 1915 -1015 1935
rect -1035 1865 -1015 1885
rect -1035 1815 -1015 1835
rect -1035 1765 -1015 1785
rect -975 2065 -955 2085
rect -975 2015 -955 2035
rect -975 1965 -955 1985
rect -975 1915 -955 1935
rect -975 1865 -955 1885
rect -975 1815 -955 1835
rect -975 1765 -955 1785
rect -915 2065 -895 2085
rect -915 2015 -895 2035
rect -915 1965 -895 1985
rect -915 1915 -895 1935
rect -915 1865 -895 1885
rect -915 1815 -895 1835
rect -915 1765 -895 1785
rect -855 2065 -835 2085
rect -855 2015 -835 2035
rect -855 1965 -835 1985
rect -855 1915 -835 1935
rect -855 1865 -835 1885
rect -855 1815 -835 1835
rect -855 1765 -835 1785
rect -795 2065 -775 2085
rect -795 2015 -775 2035
rect -795 1965 -775 1985
rect -795 1915 -775 1935
rect -795 1865 -775 1885
rect -795 1815 -775 1835
rect -795 1765 -775 1785
rect -735 2065 -715 2085
rect -735 2015 -715 2035
rect -735 1965 -715 1985
rect -735 1915 -715 1935
rect -735 1865 -715 1885
rect -735 1815 -715 1835
rect -735 1765 -715 1785
rect -675 2065 -655 2085
rect -675 2015 -655 2035
rect -675 1965 -655 1985
rect -675 1915 -655 1935
rect -675 1865 -655 1885
rect -675 1815 -655 1835
rect -675 1765 -655 1785
rect -615 2065 -595 2085
rect -615 2015 -595 2035
rect -615 1965 -595 1985
rect -615 1915 -595 1935
rect -615 1865 -595 1885
rect -615 1815 -595 1835
rect -615 1765 -595 1785
rect -555 2065 -535 2085
rect -555 2015 -535 2035
rect -555 1965 -535 1985
rect -555 1915 -535 1935
rect -555 1865 -535 1885
rect -555 1815 -535 1835
rect -555 1765 -535 1785
rect -495 2065 -475 2085
rect -495 2015 -475 2035
rect -495 1965 -475 1985
rect -495 1915 -475 1935
rect -495 1865 -475 1885
rect -495 1815 -475 1835
rect -495 1765 -475 1785
rect -435 2065 -415 2085
rect -435 2015 -415 2035
rect -435 1965 -415 1985
rect -435 1915 -415 1935
rect -435 1865 -415 1885
rect -435 1815 -415 1835
rect -435 1765 -415 1785
rect -30 2065 -10 2085
rect -30 2015 -10 2035
rect -30 1965 -10 1985
rect -30 1915 -10 1935
rect -30 1865 -10 1885
rect -30 1815 -10 1835
rect -30 1765 -10 1785
rect 30 2065 50 2085
rect 30 2015 50 2035
rect 30 1965 50 1985
rect 30 1915 50 1935
rect 30 1865 50 1885
rect 30 1815 50 1835
rect 30 1765 50 1785
rect 90 2065 110 2085
rect 90 2015 110 2035
rect 90 1965 110 1985
rect 90 1915 110 1935
rect 90 1865 110 1885
rect 90 1815 110 1835
rect 90 1765 110 1785
rect 150 2065 170 2085
rect 150 2015 170 2035
rect 150 1965 170 1985
rect 150 1915 170 1935
rect 150 1865 170 1885
rect 150 1815 170 1835
rect 150 1765 170 1785
rect 210 2065 230 2085
rect 210 2015 230 2035
rect 210 1965 230 1985
rect 210 1915 230 1935
rect 210 1865 230 1885
rect 210 1815 230 1835
rect 210 1765 230 1785
rect 270 2065 290 2085
rect 270 2015 290 2035
rect 270 1965 290 1985
rect 270 1915 290 1935
rect 270 1865 290 1885
rect 270 1815 290 1835
rect 270 1765 290 1785
rect 330 2065 350 2085
rect 330 2015 350 2035
rect 330 1965 350 1985
rect 330 1915 350 1935
rect 330 1865 350 1885
rect 330 1815 350 1835
rect 330 1765 350 1785
rect 390 2065 410 2085
rect 390 2015 410 2035
rect 390 1965 410 1985
rect 390 1915 410 1935
rect 390 1865 410 1885
rect 390 1815 410 1835
rect 390 1765 410 1785
rect 450 2065 470 2085
rect 450 2015 470 2035
rect 450 1965 470 1985
rect 450 1915 470 1935
rect 450 1865 470 1885
rect 450 1815 470 1835
rect 450 1765 470 1785
rect 510 2065 530 2085
rect 510 2015 530 2035
rect 510 1965 530 1985
rect 510 1915 530 1935
rect 510 1865 530 1885
rect 510 1815 530 1835
rect 510 1765 530 1785
rect 570 2065 590 2085
rect 570 2015 590 2035
rect 570 1965 590 1985
rect 570 1915 590 1935
rect 570 1865 590 1885
rect 570 1815 590 1835
rect 570 1765 590 1785
rect 630 2065 650 2085
rect 630 2015 650 2035
rect 630 1965 650 1985
rect 630 1915 650 1935
rect 630 1865 650 1885
rect 630 1815 650 1835
rect 630 1765 650 1785
rect 690 2065 710 2085
rect 690 2015 710 2035
rect 690 1965 710 1985
rect 690 1915 710 1935
rect 690 1865 710 1885
rect 690 1815 710 1835
rect 690 1765 710 1785
rect 980 2065 1000 2085
rect 980 2015 1000 2035
rect 980 1965 1000 1985
rect 980 1915 1000 1935
rect 980 1865 1000 1885
rect 980 1815 1000 1835
rect 980 1765 1000 1785
rect 1040 2065 1060 2085
rect 1040 2015 1060 2035
rect 1040 1965 1060 1985
rect 1040 1915 1060 1935
rect 1040 1865 1060 1885
rect 1040 1815 1060 1835
rect 1040 1765 1060 1785
rect 1100 2065 1120 2085
rect 1100 2015 1120 2035
rect 1100 1965 1120 1985
rect 1100 1915 1120 1935
rect 1100 1865 1120 1885
rect 1100 1815 1120 1835
rect 1100 1765 1120 1785
rect 1160 2065 1180 2085
rect 1160 2015 1180 2035
rect 1160 1965 1180 1985
rect 1160 1915 1180 1935
rect 1160 1865 1180 1885
rect 1160 1815 1180 1835
rect 1160 1765 1180 1785
rect 1220 2065 1240 2085
rect 1220 2015 1240 2035
rect 1220 1965 1240 1985
rect 1220 1915 1240 1935
rect 1220 1865 1240 1885
rect 1220 1815 1240 1835
rect 1220 1765 1240 1785
rect 1280 2065 1300 2085
rect 1280 2015 1300 2035
rect 1280 1965 1300 1985
rect 1280 1915 1300 1935
rect 1280 1865 1300 1885
rect 1280 1815 1300 1835
rect 1280 1765 1300 1785
rect 1340 2065 1360 2085
rect 1340 2015 1360 2035
rect 1340 1965 1360 1985
rect 1340 1915 1360 1935
rect 1340 1865 1360 1885
rect 1340 1815 1360 1835
rect 1340 1765 1360 1785
rect 1400 2065 1420 2085
rect 1400 2015 1420 2035
rect 1400 1965 1420 1985
rect 1400 1915 1420 1935
rect 1400 1865 1420 1885
rect 1400 1815 1420 1835
rect 1400 1765 1420 1785
rect 1460 2065 1480 2085
rect 1460 2015 1480 2035
rect 1460 1965 1480 1985
rect 1460 1915 1480 1935
rect 1460 1865 1480 1885
rect 1460 1815 1480 1835
rect 1460 1765 1480 1785
rect 1520 2065 1540 2085
rect 1520 2015 1540 2035
rect 1520 1965 1540 1985
rect 1520 1915 1540 1935
rect 1520 1865 1540 1885
rect 1520 1815 1540 1835
rect 1520 1765 1540 1785
rect 1580 2065 1600 2085
rect 1580 2015 1600 2035
rect 1580 1965 1600 1985
rect 1580 1915 1600 1935
rect 1580 1865 1600 1885
rect 1580 1815 1600 1835
rect 1580 1765 1600 1785
rect 1640 2065 1660 2085
rect 1640 2015 1660 2035
rect 1640 1965 1660 1985
rect 1640 1915 1660 1935
rect 1640 1865 1660 1885
rect 1640 1815 1660 1835
rect 1640 1765 1660 1785
rect 1700 2065 1720 2085
rect 1700 2015 1720 2035
rect 1700 1965 1720 1985
rect 1700 1915 1720 1935
rect 1700 1865 1720 1885
rect 1700 1815 1720 1835
rect 1700 1765 1720 1785
rect 2105 2065 2125 2085
rect 2105 2015 2125 2035
rect 2105 1965 2125 1985
rect 2105 1915 2125 1935
rect 2105 1865 2125 1885
rect 2105 1815 2125 1835
rect 2105 1765 2125 1785
rect 2165 2065 2185 2085
rect 2165 2015 2185 2035
rect 2165 1965 2185 1985
rect 2165 1915 2185 1935
rect 2165 1865 2185 1885
rect 2165 1815 2185 1835
rect 2165 1765 2185 1785
rect 2225 2065 2245 2085
rect 2225 2015 2245 2035
rect 2225 1965 2245 1985
rect 2225 1915 2245 1935
rect 2225 1865 2245 1885
rect 2225 1815 2245 1835
rect 2225 1765 2245 1785
rect 2285 2065 2305 2085
rect 2285 2015 2305 2035
rect 2285 1965 2305 1985
rect 2285 1915 2305 1935
rect 2285 1865 2305 1885
rect 2285 1815 2305 1835
rect 2285 1765 2305 1785
rect 2345 2065 2365 2085
rect 2345 2015 2365 2035
rect 2345 1965 2365 1985
rect 2345 1915 2365 1935
rect 2345 1865 2365 1885
rect 2345 1815 2365 1835
rect 2345 1765 2365 1785
rect 2405 2065 2425 2085
rect 2405 2015 2425 2035
rect 2405 1965 2425 1985
rect 2405 1915 2425 1935
rect 2405 1865 2425 1885
rect 2405 1815 2425 1835
rect 2405 1765 2425 1785
rect 2465 2065 2485 2085
rect 2465 2015 2485 2035
rect 2465 1965 2485 1985
rect 2465 1915 2485 1935
rect 2465 1865 2485 1885
rect 2465 1815 2485 1835
rect 2465 1765 2485 1785
rect 2525 2065 2545 2085
rect 2525 2015 2545 2035
rect 2525 1965 2545 1985
rect 2525 1915 2545 1935
rect 2525 1865 2545 1885
rect 2525 1815 2545 1835
rect 2525 1765 2545 1785
rect 2585 2065 2605 2085
rect 2585 2015 2605 2035
rect 2585 1965 2605 1985
rect 2585 1915 2605 1935
rect 2585 1865 2605 1885
rect 2585 1815 2605 1835
rect 2585 1765 2605 1785
rect 2645 2065 2665 2085
rect 2645 2015 2665 2035
rect 2645 1965 2665 1985
rect 2645 1915 2665 1935
rect 2645 1865 2665 1885
rect 2645 1815 2665 1835
rect 2645 1765 2665 1785
rect 2705 2065 2725 2085
rect 2705 2015 2725 2035
rect 2705 1965 2725 1985
rect 2705 1915 2725 1935
rect 2705 1865 2725 1885
rect 2705 1815 2725 1835
rect 2705 1765 2725 1785
rect 2765 2065 2785 2085
rect 2765 2015 2785 2035
rect 2765 1965 2785 1985
rect 2765 1915 2785 1935
rect 2765 1865 2785 1885
rect 2765 1815 2785 1835
rect 2765 1765 2785 1785
rect 2825 2065 2845 2085
rect 2825 2015 2845 2035
rect 2825 1965 2845 1985
rect 2825 1915 2845 1935
rect 2825 1865 2845 1885
rect 2825 1815 2845 1835
rect 2825 1765 2845 1785
rect 465 1450 485 1470
rect -1125 1400 -1105 1420
rect -1125 1350 -1105 1370
rect -1125 1300 -1105 1320
rect -1125 1250 -1105 1270
rect -1125 1200 -1105 1220
rect -1125 1150 -1105 1170
rect -1125 1100 -1105 1120
rect -1125 1050 -1105 1070
rect -1125 1000 -1105 1020
rect -1125 950 -1105 970
rect -1125 900 -1105 920
rect -1125 850 -1105 870
rect -1070 1400 -1050 1420
rect -1070 1350 -1050 1370
rect -1070 1300 -1050 1320
rect -1070 1250 -1050 1270
rect -1070 1200 -1050 1220
rect -1070 1150 -1050 1170
rect -1070 1100 -1050 1120
rect -1070 1050 -1050 1070
rect -1070 1000 -1050 1020
rect -1070 950 -1050 970
rect -1070 900 -1050 920
rect -1070 850 -1050 870
rect -1015 1400 -995 1420
rect -1015 1350 -995 1370
rect -1015 1300 -995 1320
rect -1015 1250 -995 1270
rect -1015 1200 -995 1220
rect -1015 1150 -995 1170
rect -1015 1100 -995 1120
rect -1015 1050 -995 1070
rect -1015 1000 -995 1020
rect -1015 950 -995 970
rect -1015 900 -995 920
rect -1015 850 -995 870
rect -960 1400 -940 1420
rect -960 1350 -940 1370
rect -960 1300 -940 1320
rect -960 1250 -940 1270
rect -960 1200 -940 1220
rect -960 1150 -940 1170
rect -960 1100 -940 1120
rect -960 1050 -940 1070
rect -960 1000 -940 1020
rect -960 950 -940 970
rect -960 900 -940 920
rect -960 850 -940 870
rect -905 1400 -885 1420
rect -905 1350 -885 1370
rect -905 1300 -885 1320
rect -905 1250 -885 1270
rect -905 1200 -885 1220
rect -905 1150 -885 1170
rect -905 1100 -885 1120
rect -905 1050 -885 1070
rect -905 1000 -885 1020
rect -905 950 -885 970
rect -905 900 -885 920
rect -905 850 -885 870
rect -850 1400 -830 1420
rect -850 1350 -830 1370
rect -850 1300 -830 1320
rect -850 1250 -830 1270
rect -850 1200 -830 1220
rect -850 1150 -830 1170
rect -850 1100 -830 1120
rect -850 1050 -830 1070
rect -850 1000 -830 1020
rect -850 950 -830 970
rect -850 900 -830 920
rect -850 850 -830 870
rect -795 1400 -775 1420
rect -795 1350 -775 1370
rect -795 1300 -775 1320
rect -795 1250 -775 1270
rect -795 1200 -775 1220
rect -795 1150 -775 1170
rect -795 1100 -775 1120
rect -795 1050 -775 1070
rect -795 1000 -775 1020
rect -795 950 -775 970
rect -795 900 -775 920
rect -795 850 -775 870
rect -740 1400 -720 1420
rect -740 1350 -720 1370
rect -740 1300 -720 1320
rect -740 1250 -720 1270
rect -740 1200 -720 1220
rect -740 1150 -720 1170
rect -740 1100 -720 1120
rect -740 1050 -720 1070
rect -740 1000 -720 1020
rect -740 950 -720 970
rect -740 900 -720 920
rect -740 850 -720 870
rect -685 1400 -665 1420
rect -685 1350 -665 1370
rect -685 1300 -665 1320
rect -685 1250 -665 1270
rect -685 1200 -665 1220
rect -685 1150 -665 1170
rect -685 1100 -665 1120
rect -685 1050 -665 1070
rect -685 1000 -665 1020
rect -685 950 -665 970
rect -685 900 -665 920
rect -685 850 -665 870
rect -630 1400 -610 1420
rect -630 1350 -610 1370
rect -630 1300 -610 1320
rect -630 1250 -610 1270
rect -630 1200 -610 1220
rect -630 1150 -610 1170
rect -630 1100 -610 1120
rect -630 1050 -610 1070
rect -630 1000 -610 1020
rect -630 950 -610 970
rect -630 900 -610 920
rect -630 850 -610 870
rect -575 1400 -555 1420
rect -575 1350 -555 1370
rect -575 1300 -555 1320
rect -575 1250 -555 1270
rect -575 1200 -555 1220
rect -575 1150 -555 1170
rect -575 1100 -555 1120
rect -575 1050 -555 1070
rect -575 1000 -555 1020
rect -575 950 -555 970
rect -575 900 -555 920
rect -575 850 -555 870
rect -520 1400 -500 1420
rect -520 1350 -500 1370
rect -520 1300 -500 1320
rect -520 1250 -500 1270
rect -520 1200 -500 1220
rect -520 1150 -500 1170
rect -520 1100 -500 1120
rect -520 1050 -500 1070
rect -520 1000 -500 1020
rect -520 950 -500 970
rect -520 900 -500 920
rect -520 850 -500 870
rect -465 1400 -445 1420
rect -465 1350 -445 1370
rect -465 1300 -445 1320
rect -465 1250 -445 1270
rect 465 1400 485 1420
rect 465 1350 485 1370
rect 465 1300 485 1320
rect 465 1250 485 1270
rect 520 1450 540 1470
rect 520 1400 540 1420
rect 520 1350 540 1370
rect 520 1300 540 1320
rect 520 1250 540 1270
rect 575 1450 595 1470
rect 575 1400 595 1420
rect 575 1350 595 1370
rect 575 1300 595 1320
rect 575 1250 595 1270
rect 630 1450 650 1470
rect 630 1400 650 1420
rect 630 1350 650 1370
rect 630 1300 650 1320
rect 630 1250 650 1270
rect 685 1450 705 1470
rect 685 1400 705 1420
rect 685 1350 705 1370
rect 685 1300 705 1320
rect 685 1250 705 1270
rect 740 1450 760 1470
rect 740 1400 760 1420
rect 740 1350 760 1370
rect 740 1300 760 1320
rect 740 1250 760 1270
rect 795 1450 815 1470
rect 875 1450 895 1470
rect 795 1400 815 1420
rect 875 1400 895 1420
rect 795 1350 815 1370
rect 875 1350 895 1370
rect 795 1300 815 1320
rect 875 1300 895 1320
rect 795 1250 815 1270
rect 875 1250 895 1270
rect 930 1450 950 1470
rect 930 1400 950 1420
rect 930 1350 950 1370
rect 930 1300 950 1320
rect 930 1250 950 1270
rect 985 1450 1005 1470
rect 985 1400 1005 1420
rect 985 1350 1005 1370
rect 985 1300 1005 1320
rect 985 1250 1005 1270
rect 1040 1450 1060 1470
rect 1040 1400 1060 1420
rect 1040 1350 1060 1370
rect 1040 1300 1060 1320
rect 1040 1250 1060 1270
rect 1095 1450 1115 1470
rect 1095 1400 1115 1420
rect 1095 1350 1115 1370
rect 1095 1300 1115 1320
rect 1095 1250 1115 1270
rect 1150 1450 1170 1470
rect 1150 1400 1170 1420
rect 1150 1350 1170 1370
rect 1150 1300 1170 1320
rect 1150 1250 1170 1270
rect 1205 1450 1225 1470
rect 1205 1400 1225 1420
rect 1205 1350 1225 1370
rect 1205 1300 1225 1320
rect 1205 1250 1225 1270
rect 2135 1400 2155 1420
rect 2135 1350 2155 1370
rect 2135 1300 2155 1320
rect 2135 1250 2155 1270
rect -465 1200 -445 1220
rect 2135 1200 2155 1220
rect -465 1150 -445 1170
rect -465 1100 -445 1120
rect -465 1050 -445 1070
rect -465 1000 -445 1020
rect -465 950 -445 970
rect 2135 1150 2155 1170
rect 2135 1100 2155 1120
rect 2135 1050 2155 1070
rect 2135 1000 2155 1020
rect 2135 950 2155 970
rect -465 900 -445 920
rect 2135 900 2155 920
rect -465 850 -445 870
rect 2135 850 2155 870
rect 2190 1400 2210 1420
rect 2190 1350 2210 1370
rect 2190 1300 2210 1320
rect 2190 1250 2210 1270
rect 2190 1200 2210 1220
rect 2190 1150 2210 1170
rect 2190 1100 2210 1120
rect 2190 1050 2210 1070
rect 2190 1000 2210 1020
rect 2190 950 2210 970
rect 2190 900 2210 920
rect 2190 850 2210 870
rect 2245 1400 2265 1420
rect 2245 1350 2265 1370
rect 2245 1300 2265 1320
rect 2245 1250 2265 1270
rect 2245 1200 2265 1220
rect 2245 1150 2265 1170
rect 2245 1100 2265 1120
rect 2245 1050 2265 1070
rect 2245 1000 2265 1020
rect 2245 950 2265 970
rect 2245 900 2265 920
rect 2245 850 2265 870
rect 2300 1400 2320 1420
rect 2300 1350 2320 1370
rect 2300 1300 2320 1320
rect 2300 1250 2320 1270
rect 2300 1200 2320 1220
rect 2300 1150 2320 1170
rect 2300 1100 2320 1120
rect 2300 1050 2320 1070
rect 2300 1000 2320 1020
rect 2300 950 2320 970
rect 2300 900 2320 920
rect 2300 850 2320 870
rect 2355 1400 2375 1420
rect 2355 1350 2375 1370
rect 2355 1300 2375 1320
rect 2355 1250 2375 1270
rect 2355 1200 2375 1220
rect 2355 1150 2375 1170
rect 2355 1100 2375 1120
rect 2355 1050 2375 1070
rect 2355 1000 2375 1020
rect 2355 950 2375 970
rect 2355 900 2375 920
rect 2355 850 2375 870
rect 2410 1400 2430 1420
rect 2410 1350 2430 1370
rect 2410 1300 2430 1320
rect 2410 1250 2430 1270
rect 2410 1200 2430 1220
rect 2410 1150 2430 1170
rect 2410 1100 2430 1120
rect 2410 1050 2430 1070
rect 2410 1000 2430 1020
rect 2410 950 2430 970
rect 2410 900 2430 920
rect 2410 850 2430 870
rect 2465 1400 2485 1420
rect 2465 1350 2485 1370
rect 2465 1300 2485 1320
rect 2465 1250 2485 1270
rect 2465 1200 2485 1220
rect 2465 1150 2485 1170
rect 2465 1100 2485 1120
rect 2465 1050 2485 1070
rect 2465 1000 2485 1020
rect 2465 950 2485 970
rect 2465 900 2485 920
rect 2465 850 2485 870
rect 2520 1400 2540 1420
rect 2520 1350 2540 1370
rect 2520 1300 2540 1320
rect 2520 1250 2540 1270
rect 2520 1200 2540 1220
rect 2520 1150 2540 1170
rect 2520 1100 2540 1120
rect 2520 1050 2540 1070
rect 2520 1000 2540 1020
rect 2520 950 2540 970
rect 2520 900 2540 920
rect 2520 850 2540 870
rect 2575 1400 2595 1420
rect 2575 1350 2595 1370
rect 2575 1300 2595 1320
rect 2575 1250 2595 1270
rect 2575 1200 2595 1220
rect 2575 1150 2595 1170
rect 2575 1100 2595 1120
rect 2575 1050 2595 1070
rect 2575 1000 2595 1020
rect 2575 950 2595 970
rect 2575 900 2595 920
rect 2575 850 2595 870
rect 2630 1400 2650 1420
rect 2630 1350 2650 1370
rect 2630 1300 2650 1320
rect 2630 1250 2650 1270
rect 2630 1200 2650 1220
rect 2630 1150 2650 1170
rect 2630 1100 2650 1120
rect 2630 1050 2650 1070
rect 2630 1000 2650 1020
rect 2630 950 2650 970
rect 2630 900 2650 920
rect 2630 850 2650 870
rect 2685 1400 2705 1420
rect 2685 1350 2705 1370
rect 2685 1300 2705 1320
rect 2685 1250 2705 1270
rect 2685 1200 2705 1220
rect 2685 1150 2705 1170
rect 2685 1100 2705 1120
rect 2685 1050 2705 1070
rect 2685 1000 2705 1020
rect 2685 950 2705 970
rect 2685 900 2705 920
rect 2685 850 2705 870
rect 2740 1400 2760 1420
rect 2740 1350 2760 1370
rect 2740 1300 2760 1320
rect 2740 1250 2760 1270
rect 2740 1200 2760 1220
rect 2740 1150 2760 1170
rect 2740 1100 2760 1120
rect 2740 1050 2760 1070
rect 2740 1000 2760 1020
rect 2740 950 2760 970
rect 2740 900 2760 920
rect 2740 850 2760 870
rect 2795 1400 2815 1420
rect 2795 1350 2815 1370
rect 2795 1300 2815 1320
rect 2795 1250 2815 1270
rect 2795 1200 2815 1220
rect 2795 1150 2815 1170
rect 2795 1100 2815 1120
rect 2795 1050 2815 1070
rect 2795 1000 2815 1020
rect 2795 950 2815 970
rect 2795 900 2815 920
rect 2795 850 2815 870
rect -1125 585 -1105 605
rect -1125 535 -1105 555
rect -1125 485 -1105 505
rect -1125 435 -1105 455
rect -1070 585 -1050 605
rect -1070 535 -1050 555
rect -1070 485 -1050 505
rect -1070 435 -1050 455
rect -1015 585 -995 605
rect -1015 535 -995 555
rect -1015 485 -995 505
rect -1015 435 -995 455
rect -960 585 -940 605
rect -960 535 -940 555
rect -960 485 -940 505
rect -960 435 -940 455
rect -905 585 -885 605
rect -905 535 -885 555
rect -905 485 -885 505
rect -905 435 -885 455
rect -850 585 -830 605
rect -850 535 -830 555
rect -850 485 -830 505
rect -850 435 -830 455
rect -795 585 -775 605
rect -795 535 -775 555
rect -795 485 -775 505
rect -795 435 -775 455
rect -740 585 -720 605
rect -740 535 -720 555
rect -740 485 -720 505
rect -740 435 -720 455
rect -685 585 -665 605
rect -685 535 -665 555
rect -685 485 -665 505
rect -685 435 -665 455
rect -630 585 -610 605
rect -630 535 -610 555
rect -630 485 -610 505
rect -630 435 -610 455
rect -575 585 -555 605
rect -575 535 -555 555
rect -575 485 -555 505
rect -575 435 -555 455
rect -520 585 -500 605
rect -520 535 -500 555
rect -520 485 -500 505
rect -520 435 -500 455
rect -465 585 -445 605
rect 2135 585 2155 605
rect -465 535 -445 555
rect 2135 535 2155 555
rect -465 485 -445 505
rect 2135 485 2155 505
rect -465 435 -445 455
rect 2135 435 2155 455
rect 2190 585 2210 605
rect 2190 535 2210 555
rect 2190 485 2210 505
rect 2190 435 2210 455
rect 2245 585 2265 605
rect 2245 535 2265 555
rect 2245 485 2265 505
rect 2245 435 2265 455
rect 2300 585 2320 605
rect 2300 535 2320 555
rect 2300 485 2320 505
rect 2300 435 2320 455
rect 2355 585 2375 605
rect 2355 535 2375 555
rect 2355 485 2375 505
rect 2355 435 2375 455
rect 2410 585 2430 605
rect 2410 535 2430 555
rect 2410 485 2430 505
rect 2410 435 2430 455
rect 2465 585 2485 605
rect 2465 535 2485 555
rect 2465 485 2485 505
rect 2465 435 2485 455
rect 2520 585 2540 605
rect 2520 535 2540 555
rect 2520 485 2540 505
rect 2520 435 2540 455
rect 2575 585 2595 605
rect 2575 535 2595 555
rect 2575 485 2595 505
rect 2575 435 2595 455
rect 2630 585 2650 605
rect 2630 535 2650 555
rect 2630 485 2650 505
rect 2630 435 2650 455
rect 2685 585 2705 605
rect 2685 535 2705 555
rect 2685 485 2705 505
rect 2685 435 2705 455
rect 2740 585 2760 605
rect 2740 535 2760 555
rect 2740 485 2760 505
rect 2740 435 2760 455
rect 2795 585 2815 605
rect 2795 535 2815 555
rect 2795 485 2815 505
rect 2795 435 2815 455
<< psubdiff >>
rect 675 860 715 875
rect -145 835 -105 850
rect -145 815 -135 835
rect -115 815 -105 835
rect -145 785 -105 815
rect -145 765 -135 785
rect -115 765 -105 785
rect -145 735 -105 765
rect -145 715 -135 735
rect -115 715 -105 735
rect -145 700 -105 715
rect 595 835 635 850
rect 595 815 605 835
rect 625 815 635 835
rect 595 785 635 815
rect 595 765 605 785
rect 625 765 635 785
rect 595 735 635 765
rect 595 715 605 735
rect 625 715 635 735
rect 595 700 635 715
rect 675 840 685 860
rect 705 840 715 860
rect 675 810 715 840
rect 675 790 685 810
rect 705 790 715 810
rect 675 760 715 790
rect 675 740 685 760
rect 705 740 715 760
rect 675 710 715 740
rect 675 690 685 710
rect 705 690 715 710
rect 675 660 715 690
rect 675 640 685 660
rect 705 640 715 660
rect 675 625 715 640
rect 975 860 1015 875
rect 975 840 985 860
rect 1005 840 1015 860
rect 975 810 1015 840
rect 975 790 985 810
rect 1005 790 1015 810
rect 975 760 1015 790
rect 975 740 985 760
rect 1005 740 1015 760
rect 975 710 1015 740
rect 975 690 985 710
rect 1005 690 1015 710
rect 1055 835 1095 850
rect 1055 815 1065 835
rect 1085 815 1095 835
rect 1055 785 1095 815
rect 1055 765 1065 785
rect 1085 765 1095 785
rect 1055 735 1095 765
rect 1055 715 1065 735
rect 1085 715 1095 735
rect 1055 700 1095 715
rect 1795 835 1835 850
rect 1795 815 1805 835
rect 1825 815 1835 835
rect 1795 785 1835 815
rect 1795 765 1805 785
rect 1825 765 1835 785
rect 1795 735 1835 765
rect 1795 715 1805 735
rect 1825 715 1835 735
rect 1795 700 1835 715
rect 975 660 1015 690
rect 975 640 985 660
rect 1005 640 1015 660
rect 975 625 1015 640
rect -145 440 -105 455
rect -145 420 -135 440
rect -115 420 -105 440
rect -145 390 -105 420
rect -145 370 -135 390
rect -115 370 -105 390
rect -145 340 -105 370
rect -145 320 -135 340
rect -115 320 -105 340
rect -145 305 -105 320
rect 595 440 635 455
rect 595 420 605 440
rect 625 420 635 440
rect 595 390 635 420
rect 595 370 605 390
rect 625 370 635 390
rect 595 340 635 370
rect 595 320 605 340
rect 625 320 635 340
rect 595 305 635 320
rect 675 440 715 455
rect 675 420 685 440
rect 705 420 715 440
rect 675 390 715 420
rect 675 370 685 390
rect 705 370 715 390
rect 675 340 715 370
rect 675 320 685 340
rect 705 320 715 340
rect 675 305 715 320
rect 975 440 1015 455
rect 975 420 985 440
rect 1005 420 1015 440
rect 975 390 1015 420
rect 975 370 985 390
rect 1005 370 1015 390
rect 975 340 1015 370
rect 975 320 985 340
rect 1005 320 1015 340
rect 975 305 1015 320
rect 1055 440 1095 455
rect 1055 420 1065 440
rect 1085 420 1095 440
rect 1055 390 1095 420
rect 1055 370 1065 390
rect 1085 370 1095 390
rect 1055 340 1095 370
rect 1055 320 1065 340
rect 1085 320 1095 340
rect 1055 305 1095 320
rect 1795 440 1835 455
rect 1795 420 1805 440
rect 1825 420 1835 440
rect 1795 390 1835 420
rect 1795 370 1805 390
rect 1825 370 1835 390
rect 1795 340 1835 370
rect 1795 320 1805 340
rect 1825 320 1835 340
rect 1795 305 1835 320
rect -1175 215 -1135 230
rect -1175 195 -1165 215
rect -1145 195 -1135 215
rect -1175 165 -1135 195
rect -1175 145 -1165 165
rect -1145 145 -1135 165
rect -1175 115 -1135 145
rect -1175 95 -1165 115
rect -1145 95 -1135 115
rect -1175 65 -1135 95
rect -1175 45 -1165 65
rect -1145 45 -1135 65
rect -1175 15 -1135 45
rect -1175 -5 -1165 15
rect -1145 -5 -1135 15
rect -1175 -35 -1135 -5
rect -1175 -55 -1165 -35
rect -1145 -55 -1135 -35
rect -1175 -70 -1135 -55
rect -435 215 -395 230
rect -435 195 -425 215
rect -405 195 -395 215
rect -435 165 -395 195
rect -435 145 -425 165
rect -405 145 -395 165
rect -435 115 -395 145
rect -435 95 -425 115
rect -405 95 -395 115
rect -435 65 -395 95
rect -435 45 -425 65
rect -405 45 -395 65
rect -435 15 -395 45
rect 2085 215 2125 230
rect 2085 195 2095 215
rect 2115 195 2125 215
rect 2085 165 2125 195
rect 2085 145 2095 165
rect 2115 145 2125 165
rect 2085 115 2125 145
rect 2085 95 2095 115
rect 2115 95 2125 115
rect 2085 65 2125 95
rect 2085 45 2095 65
rect 2115 45 2125 65
rect -435 -5 -425 15
rect -405 -5 -395 15
rect -435 -35 -395 -5
rect 2085 15 2125 45
rect 2085 -5 2095 15
rect 2115 -5 2125 15
rect -435 -55 -425 -35
rect -405 -55 -395 -35
rect 2085 -35 2125 -5
rect -435 -70 -395 -55
rect 675 -55 715 -40
rect 675 -75 685 -55
rect 705 -75 715 -55
rect 675 -105 715 -75
rect 675 -125 685 -105
rect 705 -125 715 -105
rect 675 -155 715 -125
rect 675 -175 685 -155
rect 705 -175 715 -155
rect 675 -205 715 -175
rect 675 -225 685 -205
rect 705 -225 715 -205
rect 675 -255 715 -225
rect 675 -275 685 -255
rect 705 -275 715 -255
rect 675 -290 715 -275
rect 975 -55 1015 -40
rect 975 -75 985 -55
rect 1005 -75 1015 -55
rect 2085 -55 2095 -35
rect 2115 -55 2125 -35
rect 2085 -70 2125 -55
rect 2825 215 2865 230
rect 2825 195 2835 215
rect 2855 195 2865 215
rect 2825 165 2865 195
rect 2825 145 2835 165
rect 2855 145 2865 165
rect 2825 115 2865 145
rect 2825 95 2835 115
rect 2855 95 2865 115
rect 2825 65 2865 95
rect 2825 45 2835 65
rect 2855 45 2865 65
rect 2825 15 2865 45
rect 2825 -5 2835 15
rect 2855 -5 2865 15
rect 2825 -35 2865 -5
rect 2825 -55 2835 -35
rect 2855 -55 2865 -35
rect 2825 -70 2865 -55
rect 975 -105 1015 -75
rect 975 -125 985 -105
rect 1005 -125 1015 -105
rect 975 -155 1015 -125
rect 975 -175 985 -155
rect 1005 -175 1015 -155
rect 975 -205 1015 -175
rect 975 -225 985 -205
rect 1005 -225 1015 -205
rect 975 -255 1015 -225
rect 975 -275 985 -255
rect 1005 -275 1015 -255
rect 975 -290 1015 -275
rect -1065 -370 -1025 -355
rect -1065 -390 -1055 -370
rect -1035 -390 -1025 -370
rect -1065 -420 -1025 -390
rect -1065 -440 -1055 -420
rect -1035 -440 -1025 -420
rect -1065 -470 -1025 -440
rect -1065 -490 -1055 -470
rect -1035 -490 -1025 -470
rect -1065 -520 -1025 -490
rect -1065 -540 -1055 -520
rect -1035 -540 -1025 -520
rect -1065 -570 -1025 -540
rect -1065 -590 -1055 -570
rect -1035 -590 -1025 -570
rect -1065 -620 -1025 -590
rect -1065 -640 -1055 -620
rect -1035 -640 -1025 -620
rect -1065 -670 -1025 -640
rect -1065 -690 -1055 -670
rect -1035 -690 -1025 -670
rect -1065 -720 -1025 -690
rect -1065 -740 -1055 -720
rect -1035 -740 -1025 -720
rect -1065 -770 -1025 -740
rect -1065 -790 -1055 -770
rect -1035 -790 -1025 -770
rect -1065 -820 -1025 -790
rect -1065 -840 -1055 -820
rect -1035 -840 -1025 -820
rect -1065 -870 -1025 -840
rect -1065 -890 -1055 -870
rect -1035 -890 -1025 -870
rect -1065 -920 -1025 -890
rect -1065 -940 -1055 -920
rect -1035 -940 -1025 -920
rect -1065 -970 -1025 -940
rect -1065 -990 -1055 -970
rect -1035 -990 -1025 -970
rect -1065 -1020 -1025 -990
rect -1065 -1040 -1055 -1020
rect -1035 -1040 -1025 -1020
rect -1065 -1055 -1025 -1040
rect -385 -370 -345 -355
rect -385 -390 -375 -370
rect -355 -390 -345 -370
rect -385 -420 -345 -390
rect -385 -440 -375 -420
rect -355 -440 -345 -420
rect -385 -470 -345 -440
rect -385 -490 -375 -470
rect -355 -490 -345 -470
rect 2035 -370 2075 -355
rect 2035 -390 2045 -370
rect 2065 -390 2075 -370
rect 2035 -420 2075 -390
rect 2035 -440 2045 -420
rect 2065 -440 2075 -420
rect 2035 -470 2075 -440
rect -385 -520 -345 -490
rect 2035 -490 2045 -470
rect 2065 -490 2075 -470
rect -385 -540 -375 -520
rect -355 -540 -345 -520
rect 2035 -520 2075 -490
rect -385 -570 -345 -540
rect -385 -590 -375 -570
rect -355 -590 -345 -570
rect -385 -620 -345 -590
rect -385 -640 -375 -620
rect -355 -640 -345 -620
rect -385 -670 -345 -640
rect -385 -690 -375 -670
rect -355 -690 -345 -670
rect -385 -720 -345 -690
rect -385 -740 -375 -720
rect -355 -740 -345 -720
rect -385 -770 -345 -740
rect -385 -790 -375 -770
rect -355 -790 -345 -770
rect 235 -550 275 -535
rect 235 -570 245 -550
rect 265 -570 275 -550
rect 235 -600 275 -570
rect 235 -620 245 -600
rect 265 -620 275 -600
rect 235 -650 275 -620
rect 235 -670 245 -650
rect 265 -670 275 -650
rect 235 -700 275 -670
rect 235 -720 245 -700
rect 265 -720 275 -700
rect 235 -750 275 -720
rect 235 -770 245 -750
rect 265 -770 275 -750
rect 235 -785 275 -770
rect 1470 -550 1510 -535
rect 1470 -570 1480 -550
rect 1500 -570 1510 -550
rect 1470 -600 1510 -570
rect 1470 -620 1480 -600
rect 1500 -620 1510 -600
rect 1470 -650 1510 -620
rect 1470 -670 1480 -650
rect 1500 -670 1510 -650
rect 1470 -700 1510 -670
rect 1470 -720 1480 -700
rect 1500 -720 1510 -700
rect 1470 -750 1510 -720
rect 1470 -770 1480 -750
rect 1500 -770 1510 -750
rect 1470 -785 1510 -770
rect 2035 -540 2045 -520
rect 2065 -540 2075 -520
rect 2035 -570 2075 -540
rect 2035 -590 2045 -570
rect 2065 -590 2075 -570
rect 2035 -620 2075 -590
rect 2035 -640 2045 -620
rect 2065 -640 2075 -620
rect 2035 -670 2075 -640
rect 2035 -690 2045 -670
rect 2065 -690 2075 -670
rect 2035 -720 2075 -690
rect 2035 -740 2045 -720
rect 2065 -740 2075 -720
rect 2035 -770 2075 -740
rect -385 -820 -345 -790
rect 2035 -790 2045 -770
rect 2065 -790 2075 -770
rect -385 -840 -375 -820
rect -355 -840 -345 -820
rect 2035 -820 2075 -790
rect 2035 -840 2045 -820
rect 2065 -840 2075 -820
rect -385 -870 -345 -840
rect -385 -890 -375 -870
rect -355 -890 -345 -870
rect -385 -920 -345 -890
rect 2035 -870 2075 -840
rect 2035 -890 2045 -870
rect 2065 -890 2075 -870
rect -385 -940 -375 -920
rect -355 -940 -345 -920
rect -385 -970 -345 -940
rect 2035 -920 2075 -890
rect 2035 -940 2045 -920
rect 2065 -940 2075 -920
rect -385 -990 -375 -970
rect -355 -990 -345 -970
rect -385 -1020 -345 -990
rect -385 -1040 -375 -1020
rect -355 -1040 -345 -1020
rect -385 -1055 -345 -1040
rect 455 -965 495 -950
rect 455 -985 465 -965
rect 485 -985 495 -965
rect 455 -1015 495 -985
rect 455 -1035 465 -1015
rect 485 -1035 495 -1015
rect 455 -1065 495 -1035
rect 455 -1085 465 -1065
rect 485 -1085 495 -1065
rect 455 -1100 495 -1085
rect 865 -965 905 -950
rect 865 -985 875 -965
rect 895 -985 905 -965
rect 865 -1015 905 -985
rect 865 -1035 875 -1015
rect 895 -1035 905 -1015
rect 865 -1065 905 -1035
rect 865 -1085 875 -1065
rect 895 -1085 905 -1065
rect 865 -1100 905 -1085
rect 2035 -970 2075 -940
rect 2035 -990 2045 -970
rect 2065 -990 2075 -970
rect 2035 -1020 2075 -990
rect 2035 -1040 2045 -1020
rect 2065 -1040 2075 -1020
rect 2035 -1055 2075 -1040
rect 2715 -370 2755 -355
rect 2715 -390 2725 -370
rect 2745 -390 2755 -370
rect 2715 -420 2755 -390
rect 2715 -440 2725 -420
rect 2745 -440 2755 -420
rect 2715 -470 2755 -440
rect 2715 -490 2725 -470
rect 2745 -490 2755 -470
rect 2715 -520 2755 -490
rect 2715 -540 2725 -520
rect 2745 -540 2755 -520
rect 2715 -570 2755 -540
rect 2715 -590 2725 -570
rect 2745 -590 2755 -570
rect 2715 -620 2755 -590
rect 2715 -640 2725 -620
rect 2745 -640 2755 -620
rect 2715 -670 2755 -640
rect 2715 -690 2725 -670
rect 2745 -690 2755 -670
rect 2715 -720 2755 -690
rect 2715 -740 2725 -720
rect 2745 -740 2755 -720
rect 2715 -770 2755 -740
rect 2715 -790 2725 -770
rect 2745 -790 2755 -770
rect 2715 -820 2755 -790
rect 2715 -840 2725 -820
rect 2745 -840 2755 -820
rect 2715 -870 2755 -840
rect 2715 -890 2725 -870
rect 2745 -890 2755 -870
rect 2715 -920 2755 -890
rect 2715 -940 2725 -920
rect 2745 -940 2755 -920
rect 2715 -970 2755 -940
rect 2715 -990 2725 -970
rect 2745 -990 2755 -970
rect 2715 -1020 2755 -990
rect 2715 -1040 2725 -1020
rect 2745 -1040 2755 -1020
rect 2715 -1055 2755 -1040
<< nsubdiff >>
rect -10 2660 30 2675
rect -10 2640 0 2660
rect 20 2640 30 2660
rect -10 2610 30 2640
rect -10 2590 0 2610
rect 20 2590 30 2610
rect -10 2560 30 2590
rect -10 2540 0 2560
rect 20 2540 30 2560
rect -10 2510 30 2540
rect -10 2490 0 2510
rect 20 2490 30 2510
rect -10 2460 30 2490
rect -10 2440 0 2460
rect 20 2440 30 2460
rect -10 2410 30 2440
rect -10 2390 0 2410
rect 20 2390 30 2410
rect -10 2360 30 2390
rect -10 2340 0 2360
rect 20 2340 30 2360
rect -10 2325 30 2340
rect 250 2660 290 2675
rect 250 2640 260 2660
rect 280 2640 290 2660
rect 250 2610 290 2640
rect 250 2590 260 2610
rect 280 2590 290 2610
rect 250 2560 290 2590
rect 930 2660 970 2675
rect 930 2640 940 2660
rect 960 2640 970 2660
rect 930 2610 970 2640
rect 930 2590 940 2610
rect 960 2590 970 2610
rect 930 2560 970 2590
rect 250 2540 260 2560
rect 280 2540 290 2560
rect 250 2510 290 2540
rect 930 2540 940 2560
rect 960 2540 970 2560
rect 250 2490 260 2510
rect 280 2490 290 2510
rect 930 2510 970 2540
rect 250 2460 290 2490
rect 250 2440 260 2460
rect 280 2440 290 2460
rect 250 2410 290 2440
rect 250 2390 260 2410
rect 280 2390 290 2410
rect 250 2360 290 2390
rect 250 2340 260 2360
rect 280 2340 290 2360
rect 250 2325 290 2340
rect 460 2360 500 2505
rect 460 2340 470 2360
rect 490 2340 500 2360
rect 460 2325 500 2340
rect 720 2360 760 2505
rect 720 2340 730 2360
rect 750 2340 760 2360
rect 720 2325 760 2340
rect 930 2490 940 2510
rect 960 2490 970 2510
rect 930 2460 970 2490
rect 930 2440 940 2460
rect 960 2440 970 2460
rect 930 2410 970 2440
rect 930 2390 940 2410
rect 960 2390 970 2410
rect 930 2360 970 2390
rect 930 2340 940 2360
rect 960 2340 970 2360
rect 930 2325 970 2340
rect 1190 2660 1230 2675
rect 1190 2640 1200 2660
rect 1220 2640 1230 2660
rect 1190 2610 1230 2640
rect 1190 2590 1200 2610
rect 1220 2590 1230 2610
rect 1190 2560 1230 2590
rect 1190 2540 1200 2560
rect 1220 2540 1230 2560
rect 1190 2510 1230 2540
rect 1190 2490 1200 2510
rect 1220 2490 1230 2510
rect 1190 2460 1230 2490
rect 1190 2440 1200 2460
rect 1220 2440 1230 2460
rect 1190 2410 1230 2440
rect 1190 2390 1200 2410
rect 1220 2390 1230 2410
rect 1190 2360 1230 2390
rect 1190 2340 1200 2360
rect 1220 2340 1230 2360
rect 1190 2325 1230 2340
rect 1398 2660 1438 2675
rect 1398 2640 1408 2660
rect 1428 2640 1438 2660
rect 1398 2610 1438 2640
rect 1398 2590 1408 2610
rect 1428 2590 1438 2610
rect 1398 2560 1438 2590
rect 1398 2540 1408 2560
rect 1428 2540 1438 2560
rect 1398 2510 1438 2540
rect 1398 2490 1408 2510
rect 1428 2490 1438 2510
rect 1398 2460 1438 2490
rect 1398 2440 1408 2460
rect 1428 2440 1438 2460
rect 1398 2410 1438 2440
rect 1398 2390 1408 2410
rect 1428 2390 1438 2410
rect 1398 2360 1438 2390
rect 1398 2340 1408 2360
rect 1428 2340 1438 2360
rect 1398 2325 1438 2340
rect 1658 2660 1698 2675
rect 1658 2640 1668 2660
rect 1688 2640 1698 2660
rect 1658 2610 1698 2640
rect 1658 2590 1668 2610
rect 1688 2590 1698 2610
rect 1658 2560 1698 2590
rect 1658 2540 1668 2560
rect 1688 2540 1698 2560
rect 1658 2510 1698 2540
rect 1658 2490 1668 2510
rect 1688 2490 1698 2510
rect 1658 2460 1698 2490
rect 1658 2440 1668 2460
rect 1688 2440 1698 2460
rect 1658 2410 1698 2440
rect 1658 2390 1668 2410
rect 1688 2390 1698 2410
rect 1658 2360 1698 2390
rect 1658 2340 1668 2360
rect 1688 2340 1698 2360
rect 1658 2325 1698 2340
rect -1205 2085 -1165 2100
rect -1205 2065 -1195 2085
rect -1175 2065 -1165 2085
rect -1205 2035 -1165 2065
rect -1205 2015 -1195 2035
rect -1175 2015 -1165 2035
rect -1205 1985 -1165 2015
rect -1205 1965 -1195 1985
rect -1175 1965 -1165 1985
rect -1205 1935 -1165 1965
rect -1205 1915 -1195 1935
rect -1175 1915 -1165 1935
rect -1205 1885 -1165 1915
rect -1205 1865 -1195 1885
rect -1175 1865 -1165 1885
rect -1205 1835 -1165 1865
rect -1205 1815 -1195 1835
rect -1175 1815 -1165 1835
rect -1205 1785 -1165 1815
rect -1205 1765 -1195 1785
rect -1175 1765 -1165 1785
rect -1205 1750 -1165 1765
rect -405 2085 -365 2100
rect -405 2065 -395 2085
rect -375 2065 -365 2085
rect -405 2035 -365 2065
rect -405 2015 -395 2035
rect -375 2015 -365 2035
rect -405 1985 -365 2015
rect -405 1965 -395 1985
rect -375 1965 -365 1985
rect -405 1935 -365 1965
rect -405 1915 -395 1935
rect -375 1915 -365 1935
rect -405 1885 -365 1915
rect -405 1865 -395 1885
rect -375 1865 -365 1885
rect -405 1835 -365 1865
rect -405 1815 -395 1835
rect -375 1815 -365 1835
rect -405 1785 -365 1815
rect -405 1765 -395 1785
rect -375 1765 -365 1785
rect -405 1750 -365 1765
rect -80 2085 -40 2100
rect -80 2065 -70 2085
rect -50 2065 -40 2085
rect -80 2035 -40 2065
rect -80 2015 -70 2035
rect -50 2015 -40 2035
rect -80 1985 -40 2015
rect -80 1965 -70 1985
rect -50 1965 -40 1985
rect -80 1935 -40 1965
rect -80 1915 -70 1935
rect -50 1915 -40 1935
rect -80 1885 -40 1915
rect -80 1865 -70 1885
rect -50 1865 -40 1885
rect -80 1835 -40 1865
rect -80 1815 -70 1835
rect -50 1815 -40 1835
rect -80 1785 -40 1815
rect -80 1765 -70 1785
rect -50 1765 -40 1785
rect -80 1750 -40 1765
rect 720 2085 760 2100
rect 720 2065 730 2085
rect 750 2065 760 2085
rect 720 2035 760 2065
rect 720 2015 730 2035
rect 750 2015 760 2035
rect 720 1985 760 2015
rect 720 1965 730 1985
rect 750 1965 760 1985
rect 720 1935 760 1965
rect 720 1915 730 1935
rect 750 1915 760 1935
rect 720 1885 760 1915
rect 720 1865 730 1885
rect 750 1865 760 1885
rect 720 1835 760 1865
rect 720 1815 730 1835
rect 750 1815 760 1835
rect 720 1785 760 1815
rect 720 1765 730 1785
rect 750 1765 760 1785
rect 720 1750 760 1765
rect 930 2085 970 2100
rect 930 2065 940 2085
rect 960 2065 970 2085
rect 930 2035 970 2065
rect 930 2015 940 2035
rect 960 2015 970 2035
rect 930 1985 970 2015
rect 930 1965 940 1985
rect 960 1965 970 1985
rect 930 1935 970 1965
rect 930 1915 940 1935
rect 960 1915 970 1935
rect 930 1885 970 1915
rect 930 1865 940 1885
rect 960 1865 970 1885
rect 930 1835 970 1865
rect 930 1815 940 1835
rect 960 1815 970 1835
rect 930 1785 970 1815
rect 930 1765 940 1785
rect 960 1765 970 1785
rect 930 1750 970 1765
rect 1730 2085 1770 2100
rect 1730 2065 1740 2085
rect 1760 2065 1770 2085
rect 1730 2035 1770 2065
rect 1730 2015 1740 2035
rect 1760 2015 1770 2035
rect 1730 1985 1770 2015
rect 1730 1965 1740 1985
rect 1760 1965 1770 1985
rect 1730 1935 1770 1965
rect 1730 1915 1740 1935
rect 1760 1915 1770 1935
rect 1730 1885 1770 1915
rect 1730 1865 1740 1885
rect 1760 1865 1770 1885
rect 1730 1835 1770 1865
rect 1730 1815 1740 1835
rect 1760 1815 1770 1835
rect 1730 1785 1770 1815
rect 1730 1765 1740 1785
rect 1760 1765 1770 1785
rect 1730 1750 1770 1765
rect 2055 2085 2095 2100
rect 2055 2065 2065 2085
rect 2085 2065 2095 2085
rect 2055 2035 2095 2065
rect 2055 2015 2065 2035
rect 2085 2015 2095 2035
rect 2055 1985 2095 2015
rect 2055 1965 2065 1985
rect 2085 1965 2095 1985
rect 2055 1935 2095 1965
rect 2055 1915 2065 1935
rect 2085 1915 2095 1935
rect 2055 1885 2095 1915
rect 2055 1865 2065 1885
rect 2085 1865 2095 1885
rect 2055 1835 2095 1865
rect 2055 1815 2065 1835
rect 2085 1815 2095 1835
rect 2055 1785 2095 1815
rect 2055 1765 2065 1785
rect 2085 1765 2095 1785
rect 2055 1750 2095 1765
rect 2855 2085 2895 2100
rect 2855 2065 2865 2085
rect 2885 2065 2895 2085
rect 2855 2035 2895 2065
rect 2855 2015 2865 2035
rect 2885 2015 2895 2035
rect 2855 1985 2895 2015
rect 2855 1965 2865 1985
rect 2885 1965 2895 1985
rect 2855 1935 2895 1965
rect 2855 1915 2865 1935
rect 2885 1915 2895 1935
rect 2855 1885 2895 1915
rect 2855 1865 2865 1885
rect 2885 1865 2895 1885
rect 2855 1835 2895 1865
rect 2855 1815 2865 1835
rect 2885 1815 2895 1835
rect 2855 1785 2895 1815
rect 2855 1765 2865 1785
rect 2885 1765 2895 1785
rect 2855 1750 2895 1765
rect 415 1470 455 1485
rect 415 1450 425 1470
rect 445 1450 455 1470
rect -1175 1420 -1135 1435
rect -1175 1400 -1165 1420
rect -1145 1400 -1135 1420
rect -1175 1370 -1135 1400
rect -1175 1350 -1165 1370
rect -1145 1350 -1135 1370
rect -1175 1320 -1135 1350
rect -1175 1300 -1165 1320
rect -1145 1300 -1135 1320
rect -1175 1270 -1135 1300
rect -1175 1250 -1165 1270
rect -1145 1250 -1135 1270
rect -1175 1220 -1135 1250
rect -1175 1200 -1165 1220
rect -1145 1200 -1135 1220
rect -1175 1170 -1135 1200
rect -1175 1150 -1165 1170
rect -1145 1150 -1135 1170
rect -1175 1120 -1135 1150
rect -1175 1100 -1165 1120
rect -1145 1100 -1135 1120
rect -1175 1070 -1135 1100
rect -1175 1050 -1165 1070
rect -1145 1050 -1135 1070
rect -1175 1020 -1135 1050
rect -1175 1000 -1165 1020
rect -1145 1000 -1135 1020
rect -1175 970 -1135 1000
rect -1175 950 -1165 970
rect -1145 950 -1135 970
rect -1175 920 -1135 950
rect -1175 900 -1165 920
rect -1145 900 -1135 920
rect -1175 870 -1135 900
rect -1175 850 -1165 870
rect -1145 850 -1135 870
rect -1175 835 -1135 850
rect -435 1420 -395 1435
rect -435 1400 -425 1420
rect -405 1400 -395 1420
rect -435 1370 -395 1400
rect -435 1350 -425 1370
rect -405 1350 -395 1370
rect -435 1320 -395 1350
rect -435 1300 -425 1320
rect -405 1300 -395 1320
rect -435 1270 -395 1300
rect -435 1250 -425 1270
rect -405 1250 -395 1270
rect -435 1220 -395 1250
rect 415 1420 455 1450
rect 415 1400 425 1420
rect 445 1400 455 1420
rect 415 1370 455 1400
rect 415 1350 425 1370
rect 445 1350 455 1370
rect 415 1320 455 1350
rect 415 1300 425 1320
rect 445 1300 455 1320
rect 415 1270 455 1300
rect 415 1250 425 1270
rect 445 1250 455 1270
rect 415 1235 455 1250
rect 825 1470 865 1485
rect 825 1450 835 1470
rect 855 1450 865 1470
rect 825 1420 865 1450
rect 825 1400 835 1420
rect 855 1400 865 1420
rect 825 1370 865 1400
rect 825 1350 835 1370
rect 855 1350 865 1370
rect 825 1320 865 1350
rect 825 1300 835 1320
rect 855 1300 865 1320
rect 825 1270 865 1300
rect 825 1250 835 1270
rect 855 1250 865 1270
rect 825 1235 865 1250
rect 1235 1470 1275 1485
rect 1235 1450 1245 1470
rect 1265 1450 1275 1470
rect 1235 1420 1275 1450
rect 1235 1400 1245 1420
rect 1265 1400 1275 1420
rect 1235 1370 1275 1400
rect 1235 1350 1245 1370
rect 1265 1350 1275 1370
rect 1235 1320 1275 1350
rect 1235 1300 1245 1320
rect 1265 1300 1275 1320
rect 1235 1270 1275 1300
rect 1235 1250 1245 1270
rect 1265 1250 1275 1270
rect 1235 1235 1275 1250
rect 2085 1420 2125 1435
rect 2085 1400 2095 1420
rect 2115 1400 2125 1420
rect 2085 1370 2125 1400
rect 2085 1350 2095 1370
rect 2115 1350 2125 1370
rect 2085 1320 2125 1350
rect 2085 1300 2095 1320
rect 2115 1300 2125 1320
rect 2085 1270 2125 1300
rect 2085 1250 2095 1270
rect 2115 1250 2125 1270
rect -435 1200 -425 1220
rect -405 1200 -395 1220
rect 2085 1220 2125 1250
rect -435 1170 -395 1200
rect 2085 1200 2095 1220
rect 2115 1200 2125 1220
rect -435 1150 -425 1170
rect -405 1150 -395 1170
rect -435 1120 -395 1150
rect -435 1100 -425 1120
rect -405 1100 -395 1120
rect -435 1070 -395 1100
rect -435 1050 -425 1070
rect -405 1050 -395 1070
rect -435 1020 -395 1050
rect -435 1000 -425 1020
rect -405 1000 -395 1020
rect -435 970 -395 1000
rect -435 950 -425 970
rect -405 950 -395 970
rect -435 920 -395 950
rect 2085 1170 2125 1200
rect 2085 1150 2095 1170
rect 2115 1150 2125 1170
rect 2085 1120 2125 1150
rect 2085 1100 2095 1120
rect 2115 1100 2125 1120
rect 2085 1070 2125 1100
rect 2085 1050 2095 1070
rect 2115 1050 2125 1070
rect 2085 1020 2125 1050
rect 2085 1000 2095 1020
rect 2115 1000 2125 1020
rect 2085 970 2125 1000
rect 2085 950 2095 970
rect 2115 950 2125 970
rect -435 900 -425 920
rect -405 900 -395 920
rect -435 870 -395 900
rect 2085 920 2125 950
rect 2085 900 2095 920
rect 2115 900 2125 920
rect -435 850 -425 870
rect -405 850 -395 870
rect -435 835 -395 850
rect 2085 870 2125 900
rect 2085 850 2095 870
rect 2115 850 2125 870
rect 2085 835 2125 850
rect 2825 1420 2865 1435
rect 2825 1400 2835 1420
rect 2855 1400 2865 1420
rect 2825 1370 2865 1400
rect 2825 1350 2835 1370
rect 2855 1350 2865 1370
rect 2825 1320 2865 1350
rect 2825 1300 2835 1320
rect 2855 1300 2865 1320
rect 2825 1270 2865 1300
rect 2825 1250 2835 1270
rect 2855 1250 2865 1270
rect 2825 1220 2865 1250
rect 2825 1200 2835 1220
rect 2855 1200 2865 1220
rect 2825 1170 2865 1200
rect 2825 1150 2835 1170
rect 2855 1150 2865 1170
rect 2825 1120 2865 1150
rect 2825 1100 2835 1120
rect 2855 1100 2865 1120
rect 2825 1070 2865 1100
rect 2825 1050 2835 1070
rect 2855 1050 2865 1070
rect 2825 1020 2865 1050
rect 2825 1000 2835 1020
rect 2855 1000 2865 1020
rect 2825 970 2865 1000
rect 2825 950 2835 970
rect 2855 950 2865 970
rect 2825 920 2865 950
rect 2825 900 2835 920
rect 2855 900 2865 920
rect 2825 870 2865 900
rect 2825 850 2835 870
rect 2855 850 2865 870
rect 2825 835 2865 850
rect -1175 605 -1135 620
rect -1175 585 -1165 605
rect -1145 585 -1135 605
rect -1175 555 -1135 585
rect -1175 535 -1165 555
rect -1145 535 -1135 555
rect -1175 505 -1135 535
rect -1175 485 -1165 505
rect -1145 485 -1135 505
rect -1175 455 -1135 485
rect -1175 435 -1165 455
rect -1145 435 -1135 455
rect -1175 420 -1135 435
rect -435 605 -395 620
rect -435 585 -425 605
rect -405 585 -395 605
rect -435 555 -395 585
rect 2085 605 2125 620
rect 2085 585 2095 605
rect 2115 585 2125 605
rect -435 535 -425 555
rect -405 535 -395 555
rect -435 505 -395 535
rect 2085 555 2125 585
rect 2085 535 2095 555
rect 2115 535 2125 555
rect -435 485 -425 505
rect -405 485 -395 505
rect -435 455 -395 485
rect 2085 505 2125 535
rect 2085 485 2095 505
rect 2115 485 2125 505
rect 2085 455 2125 485
rect -435 435 -425 455
rect -405 435 -395 455
rect -435 420 -395 435
rect 2085 435 2095 455
rect 2115 435 2125 455
rect 2085 420 2125 435
rect 2825 605 2865 620
rect 2825 585 2835 605
rect 2855 585 2865 605
rect 2825 555 2865 585
rect 2825 535 2835 555
rect 2855 535 2865 555
rect 2825 505 2865 535
rect 2825 485 2835 505
rect 2855 485 2865 505
rect 2825 455 2865 485
rect 2825 435 2835 455
rect 2855 435 2865 455
rect 2825 420 2865 435
<< psubdiffcont >>
rect -135 815 -115 835
rect -135 765 -115 785
rect -135 715 -115 735
rect 605 815 625 835
rect 605 765 625 785
rect 605 715 625 735
rect 685 840 705 860
rect 685 790 705 810
rect 685 740 705 760
rect 685 690 705 710
rect 685 640 705 660
rect 985 840 1005 860
rect 985 790 1005 810
rect 985 740 1005 760
rect 985 690 1005 710
rect 1065 815 1085 835
rect 1065 765 1085 785
rect 1065 715 1085 735
rect 1805 815 1825 835
rect 1805 765 1825 785
rect 1805 715 1825 735
rect 985 640 1005 660
rect -135 420 -115 440
rect -135 370 -115 390
rect -135 320 -115 340
rect 605 420 625 440
rect 605 370 625 390
rect 605 320 625 340
rect 685 420 705 440
rect 685 370 705 390
rect 685 320 705 340
rect 985 420 1005 440
rect 985 370 1005 390
rect 985 320 1005 340
rect 1065 420 1085 440
rect 1065 370 1085 390
rect 1065 320 1085 340
rect 1805 420 1825 440
rect 1805 370 1825 390
rect 1805 320 1825 340
rect -1165 195 -1145 215
rect -1165 145 -1145 165
rect -1165 95 -1145 115
rect -1165 45 -1145 65
rect -1165 -5 -1145 15
rect -1165 -55 -1145 -35
rect -425 195 -405 215
rect -425 145 -405 165
rect -425 95 -405 115
rect -425 45 -405 65
rect 2095 195 2115 215
rect 2095 145 2115 165
rect 2095 95 2115 115
rect 2095 45 2115 65
rect -425 -5 -405 15
rect 2095 -5 2115 15
rect -425 -55 -405 -35
rect 685 -75 705 -55
rect 685 -125 705 -105
rect 685 -175 705 -155
rect 685 -225 705 -205
rect 685 -275 705 -255
rect 985 -75 1005 -55
rect 2095 -55 2115 -35
rect 2835 195 2855 215
rect 2835 145 2855 165
rect 2835 95 2855 115
rect 2835 45 2855 65
rect 2835 -5 2855 15
rect 2835 -55 2855 -35
rect 985 -125 1005 -105
rect 985 -175 1005 -155
rect 985 -225 1005 -205
rect 985 -275 1005 -255
rect -1055 -390 -1035 -370
rect -1055 -440 -1035 -420
rect -1055 -490 -1035 -470
rect -1055 -540 -1035 -520
rect -1055 -590 -1035 -570
rect -1055 -640 -1035 -620
rect -1055 -690 -1035 -670
rect -1055 -740 -1035 -720
rect -1055 -790 -1035 -770
rect -1055 -840 -1035 -820
rect -1055 -890 -1035 -870
rect -1055 -940 -1035 -920
rect -1055 -990 -1035 -970
rect -1055 -1040 -1035 -1020
rect -375 -390 -355 -370
rect -375 -440 -355 -420
rect -375 -490 -355 -470
rect 2045 -390 2065 -370
rect 2045 -440 2065 -420
rect 2045 -490 2065 -470
rect -375 -540 -355 -520
rect -375 -590 -355 -570
rect -375 -640 -355 -620
rect -375 -690 -355 -670
rect -375 -740 -355 -720
rect -375 -790 -355 -770
rect 245 -570 265 -550
rect 245 -620 265 -600
rect 245 -670 265 -650
rect 245 -720 265 -700
rect 245 -770 265 -750
rect 1480 -570 1500 -550
rect 1480 -620 1500 -600
rect 1480 -670 1500 -650
rect 1480 -720 1500 -700
rect 1480 -770 1500 -750
rect 2045 -540 2065 -520
rect 2045 -590 2065 -570
rect 2045 -640 2065 -620
rect 2045 -690 2065 -670
rect 2045 -740 2065 -720
rect 2045 -790 2065 -770
rect -375 -840 -355 -820
rect 2045 -840 2065 -820
rect -375 -890 -355 -870
rect 2045 -890 2065 -870
rect -375 -940 -355 -920
rect 2045 -940 2065 -920
rect -375 -990 -355 -970
rect -375 -1040 -355 -1020
rect 465 -985 485 -965
rect 465 -1035 485 -1015
rect 465 -1085 485 -1065
rect 875 -985 895 -965
rect 875 -1035 895 -1015
rect 875 -1085 895 -1065
rect 2045 -990 2065 -970
rect 2045 -1040 2065 -1020
rect 2725 -390 2745 -370
rect 2725 -440 2745 -420
rect 2725 -490 2745 -470
rect 2725 -540 2745 -520
rect 2725 -590 2745 -570
rect 2725 -640 2745 -620
rect 2725 -690 2745 -670
rect 2725 -740 2745 -720
rect 2725 -790 2745 -770
rect 2725 -840 2745 -820
rect 2725 -890 2745 -870
rect 2725 -940 2745 -920
rect 2725 -990 2745 -970
rect 2725 -1040 2745 -1020
<< nsubdiffcont >>
rect 0 2640 20 2660
rect 0 2590 20 2610
rect 0 2540 20 2560
rect 0 2490 20 2510
rect 0 2440 20 2460
rect 0 2390 20 2410
rect 0 2340 20 2360
rect 260 2640 280 2660
rect 260 2590 280 2610
rect 940 2640 960 2660
rect 940 2590 960 2610
rect 260 2540 280 2560
rect 940 2540 960 2560
rect 260 2490 280 2510
rect 260 2440 280 2460
rect 260 2390 280 2410
rect 260 2340 280 2360
rect 470 2340 490 2360
rect 730 2340 750 2360
rect 940 2490 960 2510
rect 940 2440 960 2460
rect 940 2390 960 2410
rect 940 2340 960 2360
rect 1200 2640 1220 2660
rect 1200 2590 1220 2610
rect 1200 2540 1220 2560
rect 1200 2490 1220 2510
rect 1200 2440 1220 2460
rect 1200 2390 1220 2410
rect 1200 2340 1220 2360
rect 1408 2640 1428 2660
rect 1408 2590 1428 2610
rect 1408 2540 1428 2560
rect 1408 2490 1428 2510
rect 1408 2440 1428 2460
rect 1408 2390 1428 2410
rect 1408 2340 1428 2360
rect 1668 2640 1688 2660
rect 1668 2590 1688 2610
rect 1668 2540 1688 2560
rect 1668 2490 1688 2510
rect 1668 2440 1688 2460
rect 1668 2390 1688 2410
rect 1668 2340 1688 2360
rect -1195 2065 -1175 2085
rect -1195 2015 -1175 2035
rect -1195 1965 -1175 1985
rect -1195 1915 -1175 1935
rect -1195 1865 -1175 1885
rect -1195 1815 -1175 1835
rect -1195 1765 -1175 1785
rect -395 2065 -375 2085
rect -395 2015 -375 2035
rect -395 1965 -375 1985
rect -395 1915 -375 1935
rect -395 1865 -375 1885
rect -395 1815 -375 1835
rect -395 1765 -375 1785
rect -70 2065 -50 2085
rect -70 2015 -50 2035
rect -70 1965 -50 1985
rect -70 1915 -50 1935
rect -70 1865 -50 1885
rect -70 1815 -50 1835
rect -70 1765 -50 1785
rect 730 2065 750 2085
rect 730 2015 750 2035
rect 730 1965 750 1985
rect 730 1915 750 1935
rect 730 1865 750 1885
rect 730 1815 750 1835
rect 730 1765 750 1785
rect 940 2065 960 2085
rect 940 2015 960 2035
rect 940 1965 960 1985
rect 940 1915 960 1935
rect 940 1865 960 1885
rect 940 1815 960 1835
rect 940 1765 960 1785
rect 1740 2065 1760 2085
rect 1740 2015 1760 2035
rect 1740 1965 1760 1985
rect 1740 1915 1760 1935
rect 1740 1865 1760 1885
rect 1740 1815 1760 1835
rect 1740 1765 1760 1785
rect 2065 2065 2085 2085
rect 2065 2015 2085 2035
rect 2065 1965 2085 1985
rect 2065 1915 2085 1935
rect 2065 1865 2085 1885
rect 2065 1815 2085 1835
rect 2065 1765 2085 1785
rect 2865 2065 2885 2085
rect 2865 2015 2885 2035
rect 2865 1965 2885 1985
rect 2865 1915 2885 1935
rect 2865 1865 2885 1885
rect 2865 1815 2885 1835
rect 2865 1765 2885 1785
rect 425 1450 445 1470
rect -1165 1400 -1145 1420
rect -1165 1350 -1145 1370
rect -1165 1300 -1145 1320
rect -1165 1250 -1145 1270
rect -1165 1200 -1145 1220
rect -1165 1150 -1145 1170
rect -1165 1100 -1145 1120
rect -1165 1050 -1145 1070
rect -1165 1000 -1145 1020
rect -1165 950 -1145 970
rect -1165 900 -1145 920
rect -1165 850 -1145 870
rect -425 1400 -405 1420
rect -425 1350 -405 1370
rect -425 1300 -405 1320
rect -425 1250 -405 1270
rect 425 1400 445 1420
rect 425 1350 445 1370
rect 425 1300 445 1320
rect 425 1250 445 1270
rect 835 1450 855 1470
rect 835 1400 855 1420
rect 835 1350 855 1370
rect 835 1300 855 1320
rect 835 1250 855 1270
rect 1245 1450 1265 1470
rect 1245 1400 1265 1420
rect 1245 1350 1265 1370
rect 1245 1300 1265 1320
rect 1245 1250 1265 1270
rect 2095 1400 2115 1420
rect 2095 1350 2115 1370
rect 2095 1300 2115 1320
rect 2095 1250 2115 1270
rect -425 1200 -405 1220
rect 2095 1200 2115 1220
rect -425 1150 -405 1170
rect -425 1100 -405 1120
rect -425 1050 -405 1070
rect -425 1000 -405 1020
rect -425 950 -405 970
rect 2095 1150 2115 1170
rect 2095 1100 2115 1120
rect 2095 1050 2115 1070
rect 2095 1000 2115 1020
rect 2095 950 2115 970
rect -425 900 -405 920
rect 2095 900 2115 920
rect -425 850 -405 870
rect 2095 850 2115 870
rect 2835 1400 2855 1420
rect 2835 1350 2855 1370
rect 2835 1300 2855 1320
rect 2835 1250 2855 1270
rect 2835 1200 2855 1220
rect 2835 1150 2855 1170
rect 2835 1100 2855 1120
rect 2835 1050 2855 1070
rect 2835 1000 2855 1020
rect 2835 950 2855 970
rect 2835 900 2855 920
rect 2835 850 2855 870
rect -1165 585 -1145 605
rect -1165 535 -1145 555
rect -1165 485 -1145 505
rect -1165 435 -1145 455
rect -425 585 -405 605
rect 2095 585 2115 605
rect -425 535 -405 555
rect 2095 535 2115 555
rect -425 485 -405 505
rect 2095 485 2115 505
rect -425 435 -405 455
rect 2095 435 2115 455
rect 2835 585 2855 605
rect 2835 535 2855 555
rect 2835 485 2855 505
rect 2835 435 2855 455
<< poly >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2705 70 2720
rect 210 2720 250 2730
rect 210 2705 220 2720
rect 60 2700 90 2705
rect 30 2690 90 2700
rect 190 2700 220 2705
rect 240 2700 250 2720
rect 190 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2705 1010 2720
rect 1150 2720 1190 2730
rect 1150 2705 1160 2720
rect 1000 2700 1030 2705
rect 970 2690 1030 2700
rect 1130 2700 1160 2705
rect 1180 2700 1190 2720
rect 1130 2690 1190 2700
rect 1438 2720 1478 2730
rect 1438 2700 1448 2720
rect 1468 2705 1478 2720
rect 1618 2720 1658 2730
rect 1618 2705 1628 2720
rect 1468 2700 1498 2705
rect 1438 2690 1498 2700
rect 1598 2700 1628 2705
rect 1648 2700 1658 2720
rect 1598 2690 1658 2700
rect 70 2675 90 2690
rect 130 2675 150 2690
rect 190 2675 210 2690
rect 1010 2675 1030 2690
rect 1070 2675 1090 2690
rect 1130 2675 1150 2690
rect 1478 2675 1498 2690
rect 1538 2675 1558 2690
rect 1598 2675 1618 2690
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2535 540 2550
rect 680 2550 720 2560
rect 680 2535 690 2550
rect 530 2530 560 2535
rect 500 2520 560 2530
rect 660 2530 690 2535
rect 710 2530 720 2550
rect 660 2520 720 2530
rect 540 2505 560 2520
rect 600 2505 620 2520
rect 660 2505 680 2520
rect 70 2310 90 2325
rect 130 2310 150 2325
rect 190 2310 210 2325
rect 540 2310 560 2325
rect 600 2310 620 2325
rect 660 2310 680 2325
rect 1010 2310 1030 2325
rect 1070 2310 1090 2325
rect 1130 2310 1150 2325
rect 1478 2310 1498 2325
rect 1538 2310 1558 2325
rect 1598 2310 1618 2325
rect 130 2300 169 2310
rect 130 2295 144 2300
rect 139 2280 144 2295
rect 164 2280 169 2300
rect 600 2300 639 2310
rect 600 2295 614 2300
rect 139 2270 169 2280
rect 609 2280 614 2295
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1090 2310
rect 1051 2280 1056 2300
rect 1076 2295 1090 2300
rect 1519 2300 1558 2310
rect 1076 2280 1081 2295
rect 1051 2270 1081 2280
rect 1519 2280 1524 2300
rect 1544 2295 1558 2300
rect 1544 2280 1549 2295
rect 1519 2270 1549 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2130 -1125 2145
rect -445 2145 -405 2155
rect -445 2130 -435 2145
rect -1135 2125 -1105 2130
rect -1165 2115 -1105 2125
rect -465 2125 -435 2130
rect -415 2125 -405 2145
rect -465 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2130 0 2145
rect 680 2145 720 2155
rect 680 2130 690 2145
rect -10 2125 20 2130
rect -40 2115 20 2125
rect 660 2125 690 2130
rect 710 2125 720 2145
rect 660 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2130 1010 2145
rect 1690 2145 1730 2155
rect 1690 2130 1700 2145
rect 1000 2125 1030 2130
rect 970 2115 1030 2125
rect 1670 2125 1700 2130
rect 1720 2125 1730 2145
rect 1670 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2130 2135 2145
rect 2815 2145 2855 2155
rect 2815 2130 2825 2145
rect 2125 2125 2155 2130
rect 2095 2115 2155 2125
rect 2795 2125 2825 2130
rect 2845 2125 2855 2145
rect 2795 2115 2855 2125
rect -1125 2100 -1105 2115
rect -1065 2100 -1045 2115
rect -1005 2100 -985 2115
rect -945 2100 -925 2115
rect -885 2100 -865 2115
rect -825 2100 -805 2115
rect -765 2100 -745 2115
rect -705 2100 -685 2115
rect -645 2100 -625 2115
rect -585 2100 -565 2115
rect -525 2100 -505 2115
rect -465 2100 -445 2115
rect 0 2100 20 2115
rect 60 2100 80 2115
rect 120 2100 140 2115
rect 180 2100 200 2115
rect 240 2100 260 2115
rect 300 2100 320 2115
rect 360 2100 380 2115
rect 420 2100 440 2115
rect 480 2100 500 2115
rect 540 2100 560 2115
rect 600 2100 620 2115
rect 660 2100 680 2115
rect 1010 2100 1030 2115
rect 1070 2100 1090 2115
rect 1130 2100 1150 2115
rect 1190 2100 1210 2115
rect 1250 2100 1270 2115
rect 1310 2100 1330 2115
rect 1370 2100 1390 2115
rect 1430 2100 1450 2115
rect 1490 2100 1510 2115
rect 1550 2100 1570 2115
rect 1610 2100 1630 2115
rect 1670 2100 1690 2115
rect 2135 2100 2155 2115
rect 2195 2100 2215 2115
rect 2255 2100 2275 2115
rect 2315 2100 2335 2115
rect 2375 2100 2395 2115
rect 2435 2100 2455 2115
rect 2495 2100 2515 2115
rect 2555 2100 2575 2115
rect 2615 2100 2635 2115
rect 2675 2100 2695 2115
rect 2735 2100 2755 2115
rect 2795 2100 2815 2115
rect -1125 1735 -1105 1750
rect -1065 1740 -1045 1750
rect -1005 1740 -985 1750
rect -945 1740 -925 1750
rect -885 1740 -865 1750
rect -825 1740 -805 1750
rect -765 1740 -745 1750
rect -705 1740 -685 1750
rect -645 1740 -625 1750
rect -585 1740 -565 1750
rect -525 1740 -505 1750
rect -1065 1725 -505 1740
rect -465 1735 -445 1750
rect 0 1735 20 1750
rect 60 1740 80 1750
rect 120 1740 140 1750
rect 180 1740 200 1750
rect 240 1740 260 1750
rect 300 1740 320 1750
rect 360 1740 380 1750
rect 420 1740 440 1750
rect 480 1740 500 1750
rect 540 1740 560 1750
rect 600 1740 620 1750
rect 60 1725 620 1740
rect 660 1735 680 1750
rect 1010 1735 1030 1750
rect 1070 1740 1090 1750
rect 1130 1740 1150 1750
rect 1190 1740 1210 1750
rect 1250 1740 1270 1750
rect 1310 1740 1330 1750
rect 1370 1740 1390 1750
rect 1430 1740 1450 1750
rect 1490 1740 1510 1750
rect 1550 1740 1570 1750
rect 1610 1740 1630 1750
rect 1070 1725 1630 1740
rect 1670 1735 1690 1750
rect 2135 1735 2155 1750
rect 2195 1740 2215 1750
rect 2255 1740 2275 1750
rect 2315 1740 2335 1750
rect 2375 1740 2395 1750
rect 2435 1740 2455 1750
rect 2495 1740 2515 1750
rect 2555 1740 2575 1750
rect 2615 1740 2635 1750
rect 2675 1740 2695 1750
rect 2735 1740 2755 1750
rect 2195 1725 2755 1740
rect 2795 1735 2815 1750
rect -800 1720 -770 1725
rect -800 1700 -795 1720
rect -775 1700 -770 1720
rect -800 1690 -770 1700
rect 325 1720 355 1725
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 1335 1720 1365 1725
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 2460 1720 2490 1725
rect 2460 1700 2465 1720
rect 2485 1700 2490 1720
rect 2460 1690 2490 1700
rect 455 1575 495 1585
rect 455 1555 465 1575
rect 485 1560 495 1575
rect 785 1575 825 1585
rect 785 1560 795 1575
rect 485 1555 510 1560
rect 455 1545 510 1555
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1465 -1095 1480
rect -475 1480 -435 1490
rect 495 1485 510 1545
rect 770 1555 795 1560
rect 815 1555 825 1575
rect 770 1545 825 1555
rect 865 1575 905 1585
rect 865 1555 875 1575
rect 895 1560 905 1575
rect 1195 1575 1235 1585
rect 1195 1560 1205 1575
rect 895 1555 920 1560
rect 865 1545 920 1555
rect 550 1485 565 1500
rect 605 1485 620 1500
rect 660 1485 675 1500
rect 715 1485 730 1500
rect 770 1485 785 1545
rect 905 1485 920 1545
rect 1180 1555 1205 1560
rect 1225 1555 1235 1575
rect 1180 1545 1235 1555
rect 960 1485 975 1500
rect 1015 1485 1030 1500
rect 1070 1485 1085 1500
rect 1125 1485 1140 1500
rect 1180 1485 1195 1545
rect -475 1465 -465 1480
rect -1105 1460 -1080 1465
rect -1135 1450 -1080 1460
rect -490 1460 -465 1465
rect -445 1460 -435 1480
rect -490 1450 -435 1460
rect -1095 1435 -1080 1450
rect -1040 1435 -1025 1450
rect -985 1435 -970 1450
rect -930 1435 -915 1450
rect -875 1435 -860 1450
rect -820 1435 -805 1450
rect -765 1435 -750 1450
rect -710 1435 -695 1450
rect -655 1435 -640 1450
rect -600 1435 -585 1450
rect -545 1435 -530 1450
rect -490 1435 -475 1450
rect 2125 1480 2165 1490
rect 2125 1460 2135 1480
rect 2155 1465 2165 1480
rect 2785 1480 2825 1490
rect 2785 1465 2795 1480
rect 2155 1460 2180 1465
rect 2125 1450 2180 1460
rect 2770 1460 2795 1465
rect 2815 1460 2825 1480
rect 2770 1450 2825 1460
rect 2165 1435 2180 1450
rect 2220 1435 2235 1450
rect 2275 1435 2290 1450
rect 2330 1435 2345 1450
rect 2385 1435 2400 1450
rect 2440 1435 2455 1450
rect 2495 1435 2510 1450
rect 2550 1435 2565 1450
rect 2605 1435 2620 1450
rect 2660 1435 2675 1450
rect 2715 1435 2730 1450
rect 2770 1435 2785 1450
rect 495 1220 510 1235
rect 550 1220 565 1235
rect 605 1225 620 1235
rect 660 1225 675 1235
rect 550 1210 582 1220
rect 605 1210 675 1225
rect 715 1220 730 1235
rect 770 1220 785 1235
rect 905 1220 920 1235
rect 960 1220 975 1235
rect 1015 1225 1030 1235
rect 1070 1225 1085 1235
rect 698 1210 730 1220
rect 960 1210 992 1220
rect 1015 1210 1085 1225
rect 1125 1220 1140 1235
rect 1180 1220 1195 1235
rect 1108 1210 1140 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 698 1180 728 1190
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 962 1180 992 1190
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1108 1180 1138 1190
rect 795 920 835 930
rect 230 900 260 910
rect 230 880 235 900
rect 255 880 260 900
rect 795 900 805 920
rect 825 900 835 920
rect 1430 900 1460 910
rect 230 875 260 880
rect 755 875 770 890
rect 795 885 880 900
rect 810 875 825 885
rect 865 875 880 885
rect 920 875 935 890
rect 1430 880 1435 900
rect 1455 880 1460 900
rect 1430 875 1460 880
rect -65 850 -50 865
rect -10 860 500 875
rect -10 850 5 860
rect 45 850 60 860
rect 100 850 115 860
rect 155 850 170 860
rect 210 850 225 860
rect 265 850 280 860
rect 320 850 335 860
rect 375 850 390 860
rect 430 850 445 860
rect 485 850 500 860
rect 540 850 555 865
rect -1095 820 -1080 835
rect -1040 825 -1025 835
rect -985 825 -970 835
rect -930 825 -915 835
rect -875 825 -860 835
rect -820 825 -805 835
rect -765 825 -750 835
rect -710 825 -695 835
rect -655 825 -640 835
rect -600 825 -585 835
rect -545 825 -530 835
rect -1040 810 -530 825
rect -490 820 -475 835
rect -800 800 -770 810
rect -800 780 -795 800
rect -775 780 -770 800
rect -800 770 -770 780
rect -65 685 -50 700
rect -10 685 5 700
rect 45 685 60 700
rect 100 685 115 700
rect 155 685 170 700
rect 210 685 225 700
rect 265 685 280 700
rect 320 685 335 700
rect 375 685 390 700
rect 430 685 445 700
rect 485 685 500 700
rect 540 685 555 700
rect -100 675 -50 685
rect -1145 665 -1105 675
rect -1145 645 -1135 665
rect -1115 650 -1105 665
rect -465 665 -425 675
rect -465 650 -455 665
rect -1115 645 -1080 650
rect -1145 635 -1080 645
rect -490 645 -455 650
rect -435 645 -425 665
rect -100 655 -95 675
rect -75 670 -50 675
rect 540 675 590 685
rect 540 670 565 675
rect -75 655 -70 670
rect -100 645 -70 655
rect 560 655 565 670
rect 585 655 590 675
rect 560 645 590 655
rect -490 635 -425 645
rect -1095 620 -1080 635
rect -1040 620 -1025 635
rect -985 620 -970 635
rect -930 620 -915 635
rect -875 620 -860 635
rect -820 620 -805 635
rect -765 620 -750 635
rect -710 620 -695 635
rect -655 620 -640 635
rect -600 620 -585 635
rect -545 620 -530 635
rect -490 620 -475 635
rect 1135 850 1150 865
rect 1190 860 1700 875
rect 1190 850 1205 860
rect 1245 850 1260 860
rect 1300 850 1315 860
rect 1355 850 1370 860
rect 1410 850 1425 860
rect 1465 850 1480 860
rect 1520 850 1535 860
rect 1575 850 1590 860
rect 1630 850 1645 860
rect 1685 850 1700 860
rect 1740 850 1755 865
rect 2165 820 2180 835
rect 2220 825 2235 835
rect 2275 825 2290 835
rect 2330 825 2345 835
rect 2385 825 2400 835
rect 2440 825 2455 835
rect 2495 825 2510 835
rect 2550 825 2565 835
rect 2605 825 2620 835
rect 2660 825 2675 835
rect 2715 825 2730 835
rect 2220 810 2730 825
rect 2770 820 2785 835
rect 2460 800 2490 810
rect 2460 780 2465 800
rect 2485 780 2490 800
rect 2460 770 2490 780
rect 1135 685 1150 700
rect 1190 685 1205 700
rect 1245 685 1260 700
rect 1300 685 1315 700
rect 1355 685 1370 700
rect 1410 685 1425 700
rect 1465 685 1480 700
rect 1520 685 1535 700
rect 1575 685 1590 700
rect 1630 685 1645 700
rect 1685 685 1700 700
rect 1740 685 1755 700
rect 1100 675 1150 685
rect 1100 655 1105 675
rect 1125 670 1150 675
rect 1740 675 1790 685
rect 1740 670 1765 675
rect 1125 655 1130 670
rect 1100 645 1130 655
rect 1760 655 1765 670
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2115 665 2155 675
rect 2115 645 2125 665
rect 2145 650 2155 665
rect 2795 665 2835 675
rect 2795 650 2805 665
rect 2145 645 2180 650
rect 2115 635 2180 645
rect 2770 645 2805 650
rect 2825 645 2835 665
rect 2770 635 2835 645
rect 755 610 770 625
rect 810 610 825 625
rect 865 610 880 625
rect 920 610 935 625
rect 2165 620 2180 635
rect 2220 620 2235 635
rect 2275 620 2290 635
rect 2330 620 2345 635
rect 2385 620 2400 635
rect 2440 620 2455 635
rect 2495 620 2510 635
rect 2550 620 2565 635
rect 2605 620 2620 635
rect 2660 620 2675 635
rect 2715 620 2730 635
rect 2770 620 2785 635
rect 715 600 770 610
rect 715 580 725 600
rect 745 595 770 600
rect 920 600 975 610
rect 920 595 945 600
rect 745 580 755 595
rect 715 570 755 580
rect 935 580 945 595
rect 965 580 975 600
rect 935 570 975 580
rect 230 500 260 510
rect 230 480 235 500
rect 255 480 260 500
rect 715 500 755 510
rect 715 480 725 500
rect 745 485 755 500
rect 795 500 825 510
rect 745 480 770 485
rect -65 455 -50 470
rect -10 465 500 480
rect 715 470 770 480
rect 795 480 800 500
rect 820 480 825 500
rect 795 470 825 480
rect -10 455 5 465
rect 45 455 60 465
rect 100 455 115 465
rect 155 455 170 465
rect 210 455 225 465
rect 265 455 280 465
rect 320 455 335 465
rect 375 455 390 465
rect 430 455 445 465
rect 485 455 500 465
rect 540 455 555 470
rect 755 455 770 470
rect 810 455 825 470
rect 865 500 895 510
rect 865 480 870 500
rect 890 480 895 500
rect 935 500 975 510
rect 935 485 945 500
rect 865 470 895 480
rect 920 480 945 485
rect 965 480 975 500
rect 1430 500 1460 510
rect 1430 480 1435 500
rect 1455 480 1460 500
rect 920 470 975 480
rect 865 455 880 470
rect 920 455 935 470
rect 1135 455 1150 470
rect 1190 465 1700 480
rect 1190 455 1205 465
rect 1245 455 1260 465
rect 1300 455 1315 465
rect 1355 455 1370 465
rect 1410 455 1425 465
rect 1465 455 1480 465
rect 1520 455 1535 465
rect 1575 455 1590 465
rect 1630 455 1645 465
rect 1685 455 1700 465
rect 1740 455 1755 470
rect -1095 405 -1080 420
rect -1040 410 -1025 420
rect -985 410 -970 420
rect -930 410 -915 420
rect -875 410 -860 420
rect -820 410 -805 420
rect -765 410 -750 420
rect -710 410 -695 420
rect -655 410 -640 420
rect -600 410 -585 420
rect -545 410 -530 420
rect -1040 395 -530 410
rect -490 405 -475 420
rect -745 390 -715 395
rect -745 370 -740 390
rect -720 370 -715 390
rect -745 360 -715 370
rect 2165 405 2180 420
rect 2220 410 2235 420
rect 2275 410 2290 420
rect 2330 410 2345 420
rect 2385 410 2400 420
rect 2440 410 2455 420
rect 2495 410 2510 420
rect 2550 410 2565 420
rect 2605 410 2620 420
rect 2660 410 2675 420
rect 2715 410 2730 420
rect 2220 395 2730 410
rect 2770 405 2785 420
rect 2405 390 2435 395
rect 2405 370 2410 390
rect 2430 370 2435 390
rect 2405 360 2435 370
rect -65 290 -50 305
rect -10 290 5 305
rect 45 290 60 305
rect 100 290 115 305
rect 155 290 170 305
rect 210 290 225 305
rect 265 290 280 305
rect 320 290 335 305
rect 375 290 390 305
rect 430 290 445 305
rect 485 290 500 305
rect 540 290 555 305
rect 755 290 770 305
rect 810 290 825 305
rect 865 290 880 305
rect 920 290 935 305
rect 1135 290 1150 305
rect 1190 290 1205 305
rect 1245 290 1260 305
rect 1300 290 1315 305
rect 1355 290 1370 305
rect 1410 290 1425 305
rect 1465 290 1480 305
rect 1520 290 1535 305
rect 1575 290 1590 305
rect 1630 290 1645 305
rect 1685 290 1700 305
rect 1740 290 1755 305
rect -745 280 -715 290
rect -745 260 -740 280
rect -720 260 -715 280
rect -745 255 -715 260
rect -100 280 -50 290
rect -100 260 -95 280
rect -75 275 -50 280
rect 540 280 630 290
rect 540 275 605 280
rect -75 260 -70 275
rect -1095 230 -1080 245
rect -1040 240 -530 255
rect -100 250 -70 260
rect 600 260 605 275
rect 625 260 630 280
rect 600 250 630 260
rect 1060 280 1150 290
rect 1060 260 1065 280
rect 1085 275 1150 280
rect 1740 280 1790 290
rect 1740 275 1765 280
rect 1085 260 1090 275
rect 1060 250 1090 260
rect 1760 260 1765 275
rect 1785 260 1790 280
rect 1760 250 1790 260
rect 2405 280 2435 290
rect 2405 260 2410 280
rect 2430 260 2435 280
rect 2405 255 2435 260
rect -1040 230 -1025 240
rect -985 230 -970 240
rect -930 230 -915 240
rect -875 230 -860 240
rect -820 230 -805 240
rect -765 230 -750 240
rect -710 230 -695 240
rect -655 230 -640 240
rect -600 230 -585 240
rect -545 230 -530 240
rect -490 230 -475 245
rect 2165 230 2180 245
rect 2220 240 2730 255
rect 2220 230 2235 240
rect 2275 230 2290 240
rect 2330 230 2345 240
rect 2385 230 2400 240
rect 2440 230 2455 240
rect 2495 230 2510 240
rect 2550 230 2565 240
rect 2605 230 2620 240
rect 2660 230 2675 240
rect 2715 230 2730 240
rect 2770 230 2785 245
rect 830 10 860 20
rect 830 -10 835 10
rect 855 -10 860 10
rect 830 -15 860 -10
rect 755 -40 770 -25
rect 810 -30 880 -15
rect 810 -40 825 -30
rect 865 -40 880 -30
rect 920 -40 935 -25
rect -1095 -85 -1080 -70
rect -1040 -85 -1025 -70
rect -985 -85 -970 -70
rect -930 -85 -915 -70
rect -875 -85 -860 -70
rect -820 -85 -805 -70
rect -765 -85 -750 -70
rect -710 -85 -695 -70
rect -655 -85 -640 -70
rect -600 -85 -585 -70
rect -545 -85 -530 -70
rect -490 -85 -475 -70
rect -1145 -95 -1080 -85
rect -1145 -115 -1135 -95
rect -1115 -100 -1080 -95
rect -490 -95 -425 -85
rect -490 -100 -455 -95
rect -1115 -115 -1105 -100
rect -1145 -125 -1105 -115
rect -465 -115 -455 -100
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect 2165 -85 2180 -70
rect 2220 -85 2235 -70
rect 2275 -85 2290 -70
rect 2330 -85 2345 -70
rect 2385 -85 2400 -70
rect 2440 -85 2455 -70
rect 2495 -85 2510 -70
rect 2550 -85 2565 -70
rect 2605 -85 2620 -70
rect 2660 -85 2675 -70
rect 2715 -85 2730 -70
rect 2770 -85 2785 -70
rect 2115 -95 2180 -85
rect 2115 -115 2125 -95
rect 2145 -100 2180 -95
rect 2770 -95 2835 -85
rect 2770 -100 2805 -95
rect 2145 -115 2155 -100
rect 2115 -125 2155 -115
rect 2795 -115 2805 -100
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect -625 -305 -585 -295
rect 755 -305 770 -290
rect 810 -305 825 -290
rect 865 -305 880 -290
rect 920 -305 935 -290
rect 2275 -305 2315 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -330 -585 -325
rect 715 -315 770 -305
rect -985 -355 -925 -340
rect -885 -345 -525 -330
rect 715 -335 725 -315
rect 745 -320 770 -315
rect 920 -315 975 -305
rect 920 -320 945 -315
rect 745 -335 755 -320
rect -885 -355 -825 -345
rect -785 -355 -725 -345
rect -685 -355 -625 -345
rect -585 -355 -525 -345
rect -485 -355 -425 -340
rect 715 -345 755 -335
rect 935 -335 945 -320
rect 965 -335 975 -315
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -330 2315 -325
rect 935 -345 975 -335
rect 2115 -355 2175 -340
rect 2215 -345 2575 -330
rect 2215 -355 2275 -345
rect 2315 -355 2375 -345
rect 2415 -355 2475 -345
rect 2515 -355 2575 -345
rect 2615 -355 2675 -340
rect 445 -485 475 -475
rect 445 -505 450 -485
rect 470 -505 475 -485
rect 445 -510 475 -505
rect 1341 -485 1371 -475
rect 1341 -505 1346 -485
rect 1366 -500 1371 -485
rect 1366 -505 1375 -500
rect 315 -535 330 -520
rect 370 -525 1320 -510
rect 1341 -515 1375 -505
rect 370 -535 385 -525
rect 425 -535 440 -525
rect 480 -535 495 -525
rect 535 -535 550 -525
rect 590 -535 605 -525
rect 645 -535 660 -525
rect 700 -535 715 -525
rect 755 -535 770 -525
rect 810 -535 825 -525
rect 865 -535 880 -525
rect 920 -535 935 -525
rect 975 -535 990 -525
rect 1030 -535 1045 -525
rect 1085 -535 1100 -525
rect 1140 -535 1155 -525
rect 1195 -535 1210 -525
rect 1250 -535 1265 -525
rect 1305 -535 1320 -525
rect 1360 -535 1375 -515
rect 1415 -535 1430 -520
rect 315 -800 330 -785
rect 370 -800 385 -785
rect 425 -800 440 -785
rect 480 -800 495 -785
rect 535 -800 550 -785
rect 590 -800 605 -785
rect 645 -800 660 -785
rect 700 -800 715 -785
rect 755 -800 770 -785
rect 810 -800 825 -785
rect 865 -800 880 -785
rect 920 -800 935 -785
rect 975 -800 990 -785
rect 1030 -800 1045 -785
rect 1085 -800 1100 -785
rect 1140 -800 1155 -785
rect 1195 -800 1210 -785
rect 1250 -800 1265 -785
rect 1305 -800 1320 -785
rect 1360 -800 1375 -785
rect 1415 -800 1430 -785
rect 265 -810 330 -800
rect 265 -830 275 -810
rect 295 -815 330 -810
rect 1415 -810 1470 -800
rect 1415 -815 1440 -810
rect 295 -830 305 -815
rect 265 -840 305 -830
rect 1430 -830 1440 -815
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 660 -905 700 -895
rect 660 -925 670 -905
rect 690 -925 700 -905
rect 1005 -905 1045 -895
rect 1005 -925 1015 -905
rect 1035 -925 1045 -905
rect 535 -950 550 -935
rect 590 -940 770 -925
rect 1005 -935 1045 -925
rect 1125 -905 1165 -895
rect 1125 -925 1135 -905
rect 1155 -925 1165 -905
rect 1125 -935 1165 -925
rect 1255 -905 1295 -895
rect 1255 -925 1265 -905
rect 1285 -925 1295 -905
rect 1255 -935 1295 -925
rect 590 -950 605 -940
rect 645 -950 660 -940
rect 700 -950 715 -940
rect 755 -950 770 -940
rect 810 -950 825 -935
rect 1000 -950 1300 -935
rect -985 -1070 -925 -1055
rect -885 -1070 -825 -1055
rect -785 -1070 -725 -1055
rect -685 -1070 -625 -1055
rect -585 -1070 -525 -1055
rect -485 -1070 -425 -1055
rect -1025 -1080 -925 -1070
rect -1025 -1100 -1015 -1080
rect -995 -1085 -925 -1080
rect -485 -1080 -385 -1070
rect -485 -1085 -415 -1080
rect -995 -1100 -985 -1085
rect -1025 -1110 -985 -1100
rect -425 -1100 -415 -1085
rect -395 -1100 -385 -1080
rect 2115 -1070 2175 -1055
rect 2215 -1070 2275 -1055
rect 2315 -1070 2375 -1055
rect 2415 -1070 2475 -1055
rect 2515 -1070 2575 -1055
rect 2615 -1070 2675 -1055
rect 2075 -1080 2175 -1070
rect 2075 -1100 2085 -1080
rect 2105 -1085 2175 -1080
rect 2615 -1080 2715 -1070
rect 2615 -1085 2685 -1080
rect 2105 -1100 2115 -1085
rect -425 -1110 -385 -1100
rect 535 -1115 550 -1100
rect 590 -1115 605 -1100
rect 645 -1115 660 -1100
rect 700 -1115 715 -1100
rect 755 -1115 770 -1100
rect 810 -1115 825 -1100
rect 1000 -1115 1300 -1100
rect 2075 -1110 2115 -1100
rect 2675 -1100 2685 -1085
rect 2705 -1100 2715 -1080
rect 2675 -1110 2715 -1100
rect 500 -1125 550 -1115
rect 500 -1145 505 -1125
rect 525 -1130 550 -1125
rect 810 -1125 860 -1115
rect 810 -1130 835 -1125
rect 525 -1145 530 -1130
rect 500 -1155 530 -1145
rect 830 -1145 835 -1130
rect 855 -1145 860 -1125
rect 830 -1155 860 -1145
<< polycont >>
rect 40 2700 60 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1160 2700 1180 2720
rect 1448 2700 1468 2720
rect 1628 2700 1648 2720
rect 510 2530 530 2550
rect 690 2530 710 2550
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1524 2280 1544 2300
rect -1155 2125 -1135 2145
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect 2825 2125 2845 2145
rect -795 1700 -775 1720
rect 330 1700 350 1720
rect 1340 1700 1360 1720
rect 2465 1700 2485 1720
rect 465 1555 485 1575
rect -1125 1460 -1105 1480
rect 795 1555 815 1575
rect 875 1555 895 1575
rect 1205 1555 1225 1575
rect -465 1460 -445 1480
rect 2135 1460 2155 1480
rect 2795 1460 2815 1480
rect 557 1190 577 1210
rect 630 1190 650 1210
rect 703 1190 723 1210
rect 967 1190 987 1210
rect 1040 1190 1060 1210
rect 1113 1190 1133 1210
rect 235 880 255 900
rect 805 900 825 920
rect 1435 880 1455 900
rect -795 780 -775 800
rect -1135 645 -1115 665
rect -455 645 -435 665
rect -95 655 -75 675
rect 565 655 585 675
rect 2465 780 2485 800
rect 1105 655 1125 675
rect 1765 655 1785 675
rect 2125 645 2145 665
rect 2805 645 2825 665
rect 725 580 745 600
rect 945 580 965 600
rect 235 480 255 500
rect 725 480 745 500
rect 800 480 820 500
rect 870 480 890 500
rect 945 480 965 500
rect 1435 480 1455 500
rect -740 370 -720 390
rect 2410 370 2430 390
rect -740 260 -720 280
rect -95 260 -75 280
rect 605 260 625 280
rect 1065 260 1085 280
rect 1765 260 1785 280
rect 2410 260 2430 280
rect 835 -10 855 10
rect -1135 -115 -1115 -95
rect -455 -115 -435 -95
rect 2125 -115 2145 -95
rect 2805 -115 2825 -95
rect -615 -325 -595 -305
rect 725 -335 745 -315
rect 945 -335 965 -315
rect 2285 -325 2305 -305
rect 450 -505 470 -485
rect 1346 -505 1366 -485
rect 275 -830 295 -810
rect 1440 -830 1460 -810
rect 670 -925 690 -905
rect 1015 -925 1035 -905
rect 1135 -925 1155 -905
rect 1265 -925 1285 -905
rect -1015 -1100 -995 -1080
rect -415 -1100 -395 -1080
rect 2085 -1100 2105 -1080
rect 2685 -1100 2705 -1080
rect 505 -1145 525 -1125
rect 835 -1145 855 -1125
<< xpolycontact >>
rect -1501 1170 -1360 1390
rect -1501 825 -1360 1045
rect 3050 1170 3191 1390
rect 3050 825 3191 1045
rect -1490 297 -1455 517
rect -1490 -85 -1455 138
rect -1430 297 -1395 517
rect -1430 -85 -1395 138
rect -1370 297 -1335 517
rect -1370 -85 -1335 138
rect -1310 297 -1275 517
rect 2965 297 3000 517
rect -1310 -85 -1275 138
rect 2965 -85 3000 138
rect 3025 297 3060 517
rect 3025 -85 3060 138
rect 3085 297 3120 517
rect 3085 -85 3120 138
rect 3145 297 3180 517
rect 3145 -85 3180 138
rect -1210 -638 -1175 -415
rect -1210 -1105 -1175 -885
rect -1150 -638 -1115 -415
rect -1150 -1105 -1115 -885
rect 2805 -638 2840 -415
rect 2805 -1105 2840 -885
rect 2865 -638 2900 -415
rect 2865 -1105 2900 -885
<< ppolyres >>
rect -1501 1045 -1360 1170
rect 3050 1045 3191 1170
<< xpolyres >>
rect -1490 138 -1455 297
rect -1430 138 -1395 297
rect -1370 138 -1335 297
rect -1310 138 -1275 297
rect 2965 138 3000 297
rect 3025 138 3060 297
rect 3085 138 3120 297
rect 3145 138 3180 297
rect -1210 -885 -1175 -638
rect -1150 -885 -1115 -638
rect 2805 -885 2840 -638
rect 2865 -885 2900 -638
<< locali >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2700 70 2720
rect 30 2690 70 2700
rect 150 2720 190 2730
rect 150 2700 160 2720
rect 180 2700 190 2720
rect 150 2690 190 2700
rect 210 2720 250 2730
rect 210 2700 220 2720
rect 240 2700 250 2720
rect 210 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2700 1010 2720
rect 970 2690 1010 2700
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 1035 2690 1065 2700
rect 1090 2720 1130 2730
rect 1090 2700 1100 2720
rect 1120 2700 1130 2720
rect 1090 2690 1130 2700
rect 1150 2720 1190 2730
rect 1150 2700 1160 2720
rect 1180 2700 1190 2720
rect 1150 2690 1190 2700
rect 1438 2720 1478 2730
rect 1438 2700 1448 2720
rect 1468 2700 1478 2720
rect 1438 2690 1478 2700
rect 1498 2720 1538 2730
rect 1498 2700 1508 2720
rect 1528 2700 1538 2720
rect 1498 2690 1538 2700
rect 1618 2720 1658 2730
rect 1618 2700 1628 2720
rect 1648 2700 1658 2720
rect 1618 2690 1658 2700
rect 40 2670 60 2690
rect 160 2670 180 2690
rect 220 2670 240 2690
rect 980 2670 1000 2690
rect 1040 2670 1060 2690
rect 1100 2670 1120 2690
rect 1160 2670 1180 2690
rect 1448 2670 1468 2690
rect 1508 2670 1528 2690
rect 1628 2670 1648 2690
rect -5 2660 65 2670
rect -5 2640 0 2660
rect 20 2640 40 2660
rect 60 2640 65 2660
rect -5 2610 65 2640
rect -5 2590 0 2610
rect 20 2590 40 2610
rect 60 2590 65 2610
rect -5 2560 65 2590
rect -5 2540 0 2560
rect 20 2540 40 2560
rect 60 2540 65 2560
rect -5 2510 65 2540
rect -5 2490 0 2510
rect 20 2490 40 2510
rect 60 2490 65 2510
rect -5 2460 65 2490
rect -5 2440 0 2460
rect 20 2440 40 2460
rect 60 2440 65 2460
rect -5 2410 65 2440
rect -5 2390 0 2410
rect 20 2390 40 2410
rect 60 2390 65 2410
rect -5 2360 65 2390
rect -5 2340 0 2360
rect 20 2340 40 2360
rect 60 2340 65 2360
rect -5 2330 65 2340
rect 95 2660 125 2670
rect 95 2640 100 2660
rect 120 2640 125 2660
rect 95 2610 125 2640
rect 95 2590 100 2610
rect 120 2590 125 2610
rect 95 2560 125 2590
rect 95 2540 100 2560
rect 120 2540 125 2560
rect 95 2510 125 2540
rect 95 2490 100 2510
rect 120 2490 125 2510
rect 95 2460 125 2490
rect 95 2440 100 2460
rect 120 2440 125 2460
rect 95 2410 125 2440
rect 95 2390 100 2410
rect 120 2390 125 2410
rect 95 2360 125 2390
rect 95 2340 100 2360
rect 120 2340 125 2360
rect 95 2330 125 2340
rect 155 2660 185 2670
rect 155 2640 160 2660
rect 180 2640 185 2660
rect 155 2610 185 2640
rect 155 2590 160 2610
rect 180 2590 185 2610
rect 155 2560 185 2590
rect 155 2540 160 2560
rect 180 2540 185 2560
rect 155 2510 185 2540
rect 155 2490 160 2510
rect 180 2490 185 2510
rect 155 2460 185 2490
rect 155 2440 160 2460
rect 180 2440 185 2460
rect 155 2410 185 2440
rect 155 2390 160 2410
rect 180 2390 185 2410
rect 155 2360 185 2390
rect 155 2340 160 2360
rect 180 2340 185 2360
rect 155 2330 185 2340
rect 215 2660 285 2670
rect 215 2640 220 2660
rect 240 2640 260 2660
rect 280 2640 285 2660
rect 215 2610 285 2640
rect 215 2590 220 2610
rect 240 2590 260 2610
rect 280 2590 285 2610
rect 215 2560 285 2590
rect 935 2660 1005 2670
rect 935 2640 940 2660
rect 960 2640 980 2660
rect 1000 2640 1005 2660
rect 935 2610 1005 2640
rect 935 2590 940 2610
rect 960 2590 980 2610
rect 1000 2590 1005 2610
rect 935 2560 1005 2590
rect 215 2540 220 2560
rect 240 2540 260 2560
rect 280 2540 285 2560
rect 215 2510 285 2540
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2530 540 2550
rect 500 2520 540 2530
rect 560 2550 600 2560
rect 560 2530 570 2550
rect 590 2530 600 2550
rect 560 2520 600 2530
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 625 2520 655 2530
rect 680 2550 720 2560
rect 680 2530 690 2550
rect 710 2530 720 2550
rect 680 2520 720 2530
rect 935 2540 940 2560
rect 960 2540 980 2560
rect 1000 2540 1005 2560
rect 215 2490 220 2510
rect 240 2490 260 2510
rect 280 2490 285 2510
rect 510 2500 530 2520
rect 570 2500 590 2520
rect 630 2500 650 2520
rect 690 2500 710 2520
rect 935 2510 1005 2540
rect 215 2460 285 2490
rect 215 2440 220 2460
rect 240 2440 260 2460
rect 280 2440 285 2460
rect 215 2410 285 2440
rect 215 2390 220 2410
rect 240 2390 260 2410
rect 280 2390 285 2410
rect 215 2360 285 2390
rect 215 2340 220 2360
rect 240 2340 260 2360
rect 280 2340 285 2360
rect 215 2330 285 2340
rect 465 2360 535 2500
rect 465 2340 470 2360
rect 490 2340 510 2360
rect 530 2340 535 2360
rect 465 2330 535 2340
rect 565 2360 595 2500
rect 565 2340 570 2360
rect 590 2340 595 2360
rect 565 2330 595 2340
rect 625 2360 655 2500
rect 625 2340 630 2360
rect 650 2340 655 2360
rect 625 2330 655 2340
rect 685 2360 755 2500
rect 685 2340 690 2360
rect 710 2340 730 2360
rect 750 2340 755 2360
rect 685 2330 755 2340
rect 935 2490 940 2510
rect 960 2490 980 2510
rect 1000 2490 1005 2510
rect 935 2460 1005 2490
rect 935 2440 940 2460
rect 960 2440 980 2460
rect 1000 2440 1005 2460
rect 935 2410 1005 2440
rect 935 2390 940 2410
rect 960 2390 980 2410
rect 1000 2390 1005 2410
rect 935 2360 1005 2390
rect 935 2340 940 2360
rect 960 2340 980 2360
rect 1000 2340 1005 2360
rect 935 2330 1005 2340
rect 1035 2660 1065 2670
rect 1035 2640 1040 2660
rect 1060 2640 1065 2660
rect 1035 2610 1065 2640
rect 1035 2590 1040 2610
rect 1060 2590 1065 2610
rect 1035 2560 1065 2590
rect 1035 2540 1040 2560
rect 1060 2540 1065 2560
rect 1035 2510 1065 2540
rect 1035 2490 1040 2510
rect 1060 2490 1065 2510
rect 1035 2460 1065 2490
rect 1035 2440 1040 2460
rect 1060 2440 1065 2460
rect 1035 2410 1065 2440
rect 1035 2390 1040 2410
rect 1060 2390 1065 2410
rect 1035 2360 1065 2390
rect 1035 2340 1040 2360
rect 1060 2340 1065 2360
rect 1035 2330 1065 2340
rect 1095 2660 1125 2670
rect 1095 2640 1100 2660
rect 1120 2640 1125 2660
rect 1095 2610 1125 2640
rect 1095 2590 1100 2610
rect 1120 2590 1125 2610
rect 1095 2560 1125 2590
rect 1095 2540 1100 2560
rect 1120 2540 1125 2560
rect 1095 2510 1125 2540
rect 1095 2490 1100 2510
rect 1120 2490 1125 2510
rect 1095 2460 1125 2490
rect 1095 2440 1100 2460
rect 1120 2440 1125 2460
rect 1095 2410 1125 2440
rect 1095 2390 1100 2410
rect 1120 2390 1125 2410
rect 1095 2360 1125 2390
rect 1095 2340 1100 2360
rect 1120 2340 1125 2360
rect 1095 2330 1125 2340
rect 1155 2660 1225 2670
rect 1155 2640 1160 2660
rect 1180 2640 1200 2660
rect 1220 2640 1225 2660
rect 1155 2610 1225 2640
rect 1155 2590 1160 2610
rect 1180 2590 1200 2610
rect 1220 2590 1225 2610
rect 1155 2560 1225 2590
rect 1155 2540 1160 2560
rect 1180 2540 1200 2560
rect 1220 2540 1225 2560
rect 1155 2510 1225 2540
rect 1155 2490 1160 2510
rect 1180 2490 1200 2510
rect 1220 2490 1225 2510
rect 1155 2460 1225 2490
rect 1155 2440 1160 2460
rect 1180 2440 1200 2460
rect 1220 2440 1225 2460
rect 1155 2410 1225 2440
rect 1155 2390 1160 2410
rect 1180 2390 1200 2410
rect 1220 2390 1225 2410
rect 1155 2360 1225 2390
rect 1155 2340 1160 2360
rect 1180 2340 1200 2360
rect 1220 2340 1225 2360
rect 1155 2330 1225 2340
rect 1403 2660 1473 2670
rect 1403 2640 1408 2660
rect 1428 2640 1448 2660
rect 1468 2640 1473 2660
rect 1403 2610 1473 2640
rect 1403 2590 1408 2610
rect 1428 2590 1448 2610
rect 1468 2590 1473 2610
rect 1403 2560 1473 2590
rect 1403 2540 1408 2560
rect 1428 2540 1448 2560
rect 1468 2540 1473 2560
rect 1403 2510 1473 2540
rect 1403 2490 1408 2510
rect 1428 2490 1448 2510
rect 1468 2490 1473 2510
rect 1403 2460 1473 2490
rect 1403 2440 1408 2460
rect 1428 2440 1448 2460
rect 1468 2440 1473 2460
rect 1403 2410 1473 2440
rect 1403 2390 1408 2410
rect 1428 2390 1448 2410
rect 1468 2390 1473 2410
rect 1403 2360 1473 2390
rect 1403 2340 1408 2360
rect 1428 2340 1448 2360
rect 1468 2340 1473 2360
rect 1403 2330 1473 2340
rect 1503 2660 1533 2670
rect 1503 2640 1508 2660
rect 1528 2640 1533 2660
rect 1503 2610 1533 2640
rect 1503 2590 1508 2610
rect 1528 2590 1533 2610
rect 1503 2560 1533 2590
rect 1503 2540 1508 2560
rect 1528 2540 1533 2560
rect 1503 2510 1533 2540
rect 1503 2490 1508 2510
rect 1528 2490 1533 2510
rect 1503 2460 1533 2490
rect 1503 2440 1508 2460
rect 1528 2440 1533 2460
rect 1503 2410 1533 2440
rect 1503 2390 1508 2410
rect 1528 2390 1533 2410
rect 1503 2360 1533 2390
rect 1503 2340 1508 2360
rect 1528 2340 1533 2360
rect 1503 2330 1533 2340
rect 1563 2660 1593 2670
rect 1563 2640 1568 2660
rect 1588 2640 1593 2660
rect 1563 2610 1593 2640
rect 1563 2590 1568 2610
rect 1588 2590 1593 2610
rect 1563 2560 1593 2590
rect 1563 2540 1568 2560
rect 1588 2540 1593 2560
rect 1563 2510 1593 2540
rect 1563 2490 1568 2510
rect 1588 2490 1593 2510
rect 1563 2460 1593 2490
rect 1563 2440 1568 2460
rect 1588 2440 1593 2460
rect 1563 2410 1593 2440
rect 1563 2390 1568 2410
rect 1588 2390 1593 2410
rect 1563 2360 1593 2390
rect 1563 2340 1568 2360
rect 1588 2340 1593 2360
rect 1563 2330 1593 2340
rect 1623 2660 1693 2670
rect 1623 2640 1628 2660
rect 1648 2640 1668 2660
rect 1688 2640 1693 2660
rect 1623 2610 1693 2640
rect 1623 2590 1628 2610
rect 1648 2590 1668 2610
rect 1688 2590 1693 2610
rect 1623 2560 1693 2590
rect 1623 2540 1628 2560
rect 1648 2540 1668 2560
rect 1688 2540 1693 2560
rect 1623 2510 1693 2540
rect 1623 2490 1628 2510
rect 1648 2490 1668 2510
rect 1688 2490 1693 2510
rect 1623 2460 1693 2490
rect 1623 2440 1628 2460
rect 1648 2440 1668 2460
rect 1688 2440 1693 2460
rect 1623 2410 1693 2440
rect 1623 2390 1628 2410
rect 1648 2390 1668 2410
rect 1688 2390 1693 2410
rect 1623 2360 1693 2390
rect 1623 2340 1628 2360
rect 1648 2340 1668 2360
rect 1688 2340 1693 2360
rect 1623 2330 1693 2340
rect 95 2310 115 2330
rect 1573 2310 1593 2330
rect 75 2300 115 2310
rect 75 2280 85 2300
rect 105 2280 115 2300
rect 75 2270 115 2280
rect 139 2300 169 2310
rect 139 2280 144 2300
rect 164 2280 169 2300
rect 139 2270 169 2280
rect 609 2300 639 2310
rect 609 2280 614 2300
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1519 2300 1549 2310
rect 1519 2280 1524 2300
rect 1544 2280 1549 2300
rect 1519 2270 1549 2280
rect 1573 2300 1613 2310
rect 1573 2280 1583 2300
rect 1603 2280 1613 2300
rect 1573 2270 1613 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2125 -1125 2145
rect -1165 2115 -1125 2125
rect -1045 2145 -1005 2155
rect -1045 2125 -1035 2145
rect -1015 2125 -1005 2145
rect -1045 2115 -1005 2125
rect -925 2145 -885 2155
rect -925 2125 -915 2145
rect -895 2125 -885 2145
rect -925 2115 -885 2125
rect -805 2145 -765 2155
rect -805 2125 -795 2145
rect -775 2125 -765 2145
rect -805 2115 -765 2125
rect -685 2145 -645 2155
rect -685 2125 -675 2145
rect -655 2125 -645 2145
rect -685 2115 -645 2125
rect -565 2145 -525 2155
rect -565 2125 -555 2145
rect -535 2125 -525 2145
rect -565 2115 -525 2125
rect -445 2145 -405 2155
rect -445 2125 -435 2145
rect -415 2125 -405 2145
rect -445 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2125 0 2145
rect -40 2115 0 2125
rect 80 2145 120 2155
rect 80 2125 90 2145
rect 110 2125 120 2145
rect 80 2115 120 2125
rect 200 2145 240 2155
rect 200 2125 210 2145
rect 230 2125 240 2145
rect 200 2115 240 2125
rect 320 2145 360 2155
rect 320 2125 330 2145
rect 350 2125 360 2145
rect 320 2115 360 2125
rect 440 2145 480 2155
rect 440 2125 450 2145
rect 470 2125 480 2145
rect 440 2115 480 2125
rect 560 2145 600 2155
rect 560 2125 570 2145
rect 590 2125 600 2145
rect 560 2115 600 2125
rect 680 2145 720 2155
rect 680 2125 690 2145
rect 710 2125 720 2145
rect 680 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2125 1010 2145
rect 970 2115 1010 2125
rect 1090 2145 1130 2155
rect 1090 2125 1100 2145
rect 1120 2125 1130 2145
rect 1090 2115 1130 2125
rect 1210 2145 1250 2155
rect 1210 2125 1220 2145
rect 1240 2125 1250 2145
rect 1210 2115 1250 2125
rect 1330 2145 1370 2155
rect 1330 2125 1340 2145
rect 1360 2125 1370 2145
rect 1330 2115 1370 2125
rect 1450 2145 1490 2155
rect 1450 2125 1460 2145
rect 1480 2125 1490 2145
rect 1450 2115 1490 2125
rect 1570 2145 1610 2155
rect 1570 2125 1580 2145
rect 1600 2125 1610 2145
rect 1570 2115 1610 2125
rect 1690 2145 1730 2155
rect 1690 2125 1700 2145
rect 1720 2125 1730 2145
rect 1690 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2125 2135 2145
rect 2095 2115 2135 2125
rect 2215 2145 2255 2155
rect 2215 2125 2225 2145
rect 2245 2125 2255 2145
rect 2215 2115 2255 2125
rect 2335 2145 2375 2155
rect 2335 2125 2345 2145
rect 2365 2125 2375 2145
rect 2335 2115 2375 2125
rect 2455 2145 2495 2155
rect 2455 2125 2465 2145
rect 2485 2125 2495 2145
rect 2455 2115 2495 2125
rect 2575 2145 2615 2155
rect 2575 2125 2585 2145
rect 2605 2125 2615 2145
rect 2575 2115 2615 2125
rect 2695 2145 2735 2155
rect 2695 2125 2705 2145
rect 2725 2125 2735 2145
rect 2695 2115 2735 2125
rect 2815 2145 2855 2155
rect 2815 2125 2825 2145
rect 2845 2125 2855 2145
rect 2815 2115 2855 2125
rect -1155 2095 -1135 2115
rect -1035 2095 -1015 2115
rect -915 2095 -895 2115
rect -795 2095 -775 2115
rect -675 2095 -655 2115
rect -555 2095 -535 2115
rect -435 2095 -415 2115
rect -30 2095 -10 2115
rect 90 2095 110 2115
rect 210 2095 230 2115
rect 330 2095 350 2115
rect 450 2095 470 2115
rect 570 2095 590 2115
rect 690 2095 710 2115
rect 980 2095 1000 2115
rect 1100 2095 1120 2115
rect 1220 2095 1240 2115
rect 1340 2095 1360 2115
rect 1460 2095 1480 2115
rect 1580 2095 1600 2115
rect 1700 2095 1720 2115
rect 2105 2095 2125 2115
rect 2225 2095 2245 2115
rect 2345 2095 2365 2115
rect 2465 2095 2485 2115
rect 2585 2095 2605 2115
rect 2705 2095 2725 2115
rect 2825 2095 2845 2115
rect -1200 2085 -1130 2095
rect -1200 2065 -1195 2085
rect -1175 2065 -1155 2085
rect -1135 2065 -1130 2085
rect -1200 2035 -1130 2065
rect -1200 2015 -1195 2035
rect -1175 2015 -1155 2035
rect -1135 2015 -1130 2035
rect -1200 1985 -1130 2015
rect -1200 1965 -1195 1985
rect -1175 1965 -1155 1985
rect -1135 1965 -1130 1985
rect -1200 1935 -1130 1965
rect -1200 1915 -1195 1935
rect -1175 1915 -1155 1935
rect -1135 1915 -1130 1935
rect -1200 1885 -1130 1915
rect -1200 1865 -1195 1885
rect -1175 1865 -1155 1885
rect -1135 1865 -1130 1885
rect -1200 1835 -1130 1865
rect -1200 1815 -1195 1835
rect -1175 1815 -1155 1835
rect -1135 1815 -1130 1835
rect -1200 1785 -1130 1815
rect -1200 1765 -1195 1785
rect -1175 1765 -1155 1785
rect -1135 1765 -1130 1785
rect -1200 1755 -1130 1765
rect -1100 2085 -1070 2095
rect -1100 2065 -1095 2085
rect -1075 2065 -1070 2085
rect -1100 2035 -1070 2065
rect -1100 2015 -1095 2035
rect -1075 2015 -1070 2035
rect -1100 1985 -1070 2015
rect -1100 1965 -1095 1985
rect -1075 1965 -1070 1985
rect -1100 1935 -1070 1965
rect -1100 1915 -1095 1935
rect -1075 1915 -1070 1935
rect -1100 1885 -1070 1915
rect -1100 1865 -1095 1885
rect -1075 1865 -1070 1885
rect -1100 1835 -1070 1865
rect -1100 1815 -1095 1835
rect -1075 1815 -1070 1835
rect -1100 1785 -1070 1815
rect -1100 1765 -1095 1785
rect -1075 1765 -1070 1785
rect -1100 1755 -1070 1765
rect -1040 2085 -1010 2095
rect -1040 2065 -1035 2085
rect -1015 2065 -1010 2085
rect -1040 2035 -1010 2065
rect -1040 2015 -1035 2035
rect -1015 2015 -1010 2035
rect -1040 1985 -1010 2015
rect -1040 1965 -1035 1985
rect -1015 1965 -1010 1985
rect -1040 1935 -1010 1965
rect -1040 1915 -1035 1935
rect -1015 1915 -1010 1935
rect -1040 1885 -1010 1915
rect -1040 1865 -1035 1885
rect -1015 1865 -1010 1885
rect -1040 1835 -1010 1865
rect -1040 1815 -1035 1835
rect -1015 1815 -1010 1835
rect -1040 1785 -1010 1815
rect -1040 1765 -1035 1785
rect -1015 1765 -1010 1785
rect -1040 1755 -1010 1765
rect -980 2085 -950 2095
rect -980 2065 -975 2085
rect -955 2065 -950 2085
rect -980 2035 -950 2065
rect -980 2015 -975 2035
rect -955 2015 -950 2035
rect -980 1985 -950 2015
rect -980 1965 -975 1985
rect -955 1965 -950 1985
rect -980 1935 -950 1965
rect -980 1915 -975 1935
rect -955 1915 -950 1935
rect -980 1885 -950 1915
rect -980 1865 -975 1885
rect -955 1865 -950 1885
rect -980 1835 -950 1865
rect -980 1815 -975 1835
rect -955 1815 -950 1835
rect -980 1785 -950 1815
rect -980 1765 -975 1785
rect -955 1765 -950 1785
rect -980 1755 -950 1765
rect -920 2085 -890 2095
rect -920 2065 -915 2085
rect -895 2065 -890 2085
rect -920 2035 -890 2065
rect -920 2015 -915 2035
rect -895 2015 -890 2035
rect -920 1985 -890 2015
rect -920 1965 -915 1985
rect -895 1965 -890 1985
rect -920 1935 -890 1965
rect -920 1915 -915 1935
rect -895 1915 -890 1935
rect -920 1885 -890 1915
rect -920 1865 -915 1885
rect -895 1865 -890 1885
rect -920 1835 -890 1865
rect -920 1815 -915 1835
rect -895 1815 -890 1835
rect -920 1785 -890 1815
rect -920 1765 -915 1785
rect -895 1765 -890 1785
rect -920 1755 -890 1765
rect -860 2085 -830 2095
rect -860 2065 -855 2085
rect -835 2065 -830 2085
rect -860 2035 -830 2065
rect -860 2015 -855 2035
rect -835 2015 -830 2035
rect -860 1985 -830 2015
rect -860 1965 -855 1985
rect -835 1965 -830 1985
rect -860 1935 -830 1965
rect -860 1915 -855 1935
rect -835 1915 -830 1935
rect -860 1885 -830 1915
rect -860 1865 -855 1885
rect -835 1865 -830 1885
rect -860 1835 -830 1865
rect -860 1815 -855 1835
rect -835 1815 -830 1835
rect -860 1785 -830 1815
rect -860 1765 -855 1785
rect -835 1765 -830 1785
rect -860 1755 -830 1765
rect -800 2085 -770 2095
rect -800 2065 -795 2085
rect -775 2065 -770 2085
rect -800 2035 -770 2065
rect -800 2015 -795 2035
rect -775 2015 -770 2035
rect -800 1985 -770 2015
rect -800 1965 -795 1985
rect -775 1965 -770 1985
rect -800 1935 -770 1965
rect -800 1915 -795 1935
rect -775 1915 -770 1935
rect -800 1885 -770 1915
rect -800 1865 -795 1885
rect -775 1865 -770 1885
rect -800 1835 -770 1865
rect -800 1815 -795 1835
rect -775 1815 -770 1835
rect -800 1785 -770 1815
rect -800 1765 -795 1785
rect -775 1765 -770 1785
rect -800 1755 -770 1765
rect -740 2085 -710 2095
rect -740 2065 -735 2085
rect -715 2065 -710 2085
rect -740 2035 -710 2065
rect -740 2015 -735 2035
rect -715 2015 -710 2035
rect -740 1985 -710 2015
rect -740 1965 -735 1985
rect -715 1965 -710 1985
rect -740 1935 -710 1965
rect -740 1915 -735 1935
rect -715 1915 -710 1935
rect -740 1885 -710 1915
rect -740 1865 -735 1885
rect -715 1865 -710 1885
rect -740 1835 -710 1865
rect -740 1815 -735 1835
rect -715 1815 -710 1835
rect -740 1785 -710 1815
rect -740 1765 -735 1785
rect -715 1765 -710 1785
rect -740 1755 -710 1765
rect -680 2085 -650 2095
rect -680 2065 -675 2085
rect -655 2065 -650 2085
rect -680 2035 -650 2065
rect -680 2015 -675 2035
rect -655 2015 -650 2035
rect -680 1985 -650 2015
rect -680 1965 -675 1985
rect -655 1965 -650 1985
rect -680 1935 -650 1965
rect -680 1915 -675 1935
rect -655 1915 -650 1935
rect -680 1885 -650 1915
rect -680 1865 -675 1885
rect -655 1865 -650 1885
rect -680 1835 -650 1865
rect -680 1815 -675 1835
rect -655 1815 -650 1835
rect -680 1785 -650 1815
rect -680 1765 -675 1785
rect -655 1765 -650 1785
rect -680 1755 -650 1765
rect -620 2085 -590 2095
rect -620 2065 -615 2085
rect -595 2065 -590 2085
rect -620 2035 -590 2065
rect -620 2015 -615 2035
rect -595 2015 -590 2035
rect -620 1985 -590 2015
rect -620 1965 -615 1985
rect -595 1965 -590 1985
rect -620 1935 -590 1965
rect -620 1915 -615 1935
rect -595 1915 -590 1935
rect -620 1885 -590 1915
rect -620 1865 -615 1885
rect -595 1865 -590 1885
rect -620 1835 -590 1865
rect -620 1815 -615 1835
rect -595 1815 -590 1835
rect -620 1785 -590 1815
rect -620 1765 -615 1785
rect -595 1765 -590 1785
rect -620 1755 -590 1765
rect -560 2085 -530 2095
rect -560 2065 -555 2085
rect -535 2065 -530 2085
rect -560 2035 -530 2065
rect -560 2015 -555 2035
rect -535 2015 -530 2035
rect -560 1985 -530 2015
rect -560 1965 -555 1985
rect -535 1965 -530 1985
rect -560 1935 -530 1965
rect -560 1915 -555 1935
rect -535 1915 -530 1935
rect -560 1885 -530 1915
rect -560 1865 -555 1885
rect -535 1865 -530 1885
rect -560 1835 -530 1865
rect -560 1815 -555 1835
rect -535 1815 -530 1835
rect -560 1785 -530 1815
rect -560 1765 -555 1785
rect -535 1765 -530 1785
rect -560 1755 -530 1765
rect -500 2085 -470 2095
rect -500 2065 -495 2085
rect -475 2065 -470 2085
rect -500 2035 -470 2065
rect -500 2015 -495 2035
rect -475 2015 -470 2035
rect -500 1985 -470 2015
rect -500 1965 -495 1985
rect -475 1965 -470 1985
rect -500 1935 -470 1965
rect -500 1915 -495 1935
rect -475 1915 -470 1935
rect -500 1885 -470 1915
rect -500 1865 -495 1885
rect -475 1865 -470 1885
rect -500 1835 -470 1865
rect -500 1815 -495 1835
rect -475 1815 -470 1835
rect -500 1785 -470 1815
rect -500 1765 -495 1785
rect -475 1765 -470 1785
rect -500 1755 -470 1765
rect -440 2085 -370 2095
rect -440 2065 -435 2085
rect -415 2065 -395 2085
rect -375 2065 -370 2085
rect -440 2035 -370 2065
rect -440 2015 -435 2035
rect -415 2015 -395 2035
rect -375 2015 -370 2035
rect -440 1985 -370 2015
rect -440 1965 -435 1985
rect -415 1965 -395 1985
rect -375 1965 -370 1985
rect -440 1935 -370 1965
rect -440 1915 -435 1935
rect -415 1915 -395 1935
rect -375 1915 -370 1935
rect -440 1885 -370 1915
rect -440 1865 -435 1885
rect -415 1865 -395 1885
rect -375 1865 -370 1885
rect -440 1835 -370 1865
rect -440 1815 -435 1835
rect -415 1815 -395 1835
rect -375 1815 -370 1835
rect -440 1785 -370 1815
rect -440 1765 -435 1785
rect -415 1765 -395 1785
rect -375 1765 -370 1785
rect -440 1755 -370 1765
rect -75 2085 -5 2095
rect -75 2065 -70 2085
rect -50 2065 -30 2085
rect -10 2065 -5 2085
rect -75 2035 -5 2065
rect -75 2015 -70 2035
rect -50 2015 -30 2035
rect -10 2015 -5 2035
rect -75 1985 -5 2015
rect -75 1965 -70 1985
rect -50 1965 -30 1985
rect -10 1965 -5 1985
rect -75 1935 -5 1965
rect -75 1915 -70 1935
rect -50 1915 -30 1935
rect -10 1915 -5 1935
rect -75 1885 -5 1915
rect -75 1865 -70 1885
rect -50 1865 -30 1885
rect -10 1865 -5 1885
rect -75 1835 -5 1865
rect -75 1815 -70 1835
rect -50 1815 -30 1835
rect -10 1815 -5 1835
rect -75 1785 -5 1815
rect -75 1765 -70 1785
rect -50 1765 -30 1785
rect -10 1765 -5 1785
rect -75 1755 -5 1765
rect 25 2085 55 2095
rect 25 2065 30 2085
rect 50 2065 55 2085
rect 25 2035 55 2065
rect 25 2015 30 2035
rect 50 2015 55 2035
rect 25 1985 55 2015
rect 25 1965 30 1985
rect 50 1965 55 1985
rect 25 1935 55 1965
rect 25 1915 30 1935
rect 50 1915 55 1935
rect 25 1885 55 1915
rect 25 1865 30 1885
rect 50 1865 55 1885
rect 25 1835 55 1865
rect 25 1815 30 1835
rect 50 1815 55 1835
rect 25 1785 55 1815
rect 25 1765 30 1785
rect 50 1765 55 1785
rect 25 1755 55 1765
rect 85 2085 115 2095
rect 85 2065 90 2085
rect 110 2065 115 2085
rect 85 2035 115 2065
rect 85 2015 90 2035
rect 110 2015 115 2035
rect 85 1985 115 2015
rect 85 1965 90 1985
rect 110 1965 115 1985
rect 85 1935 115 1965
rect 85 1915 90 1935
rect 110 1915 115 1935
rect 85 1885 115 1915
rect 85 1865 90 1885
rect 110 1865 115 1885
rect 85 1835 115 1865
rect 85 1815 90 1835
rect 110 1815 115 1835
rect 85 1785 115 1815
rect 85 1765 90 1785
rect 110 1765 115 1785
rect 85 1755 115 1765
rect 145 2085 175 2095
rect 145 2065 150 2085
rect 170 2065 175 2085
rect 145 2035 175 2065
rect 145 2015 150 2035
rect 170 2015 175 2035
rect 145 1985 175 2015
rect 145 1965 150 1985
rect 170 1965 175 1985
rect 145 1935 175 1965
rect 145 1915 150 1935
rect 170 1915 175 1935
rect 145 1885 175 1915
rect 145 1865 150 1885
rect 170 1865 175 1885
rect 145 1835 175 1865
rect 145 1815 150 1835
rect 170 1815 175 1835
rect 145 1785 175 1815
rect 145 1765 150 1785
rect 170 1765 175 1785
rect 145 1755 175 1765
rect 205 2085 235 2095
rect 205 2065 210 2085
rect 230 2065 235 2085
rect 205 2035 235 2065
rect 205 2015 210 2035
rect 230 2015 235 2035
rect 205 1985 235 2015
rect 205 1965 210 1985
rect 230 1965 235 1985
rect 205 1935 235 1965
rect 205 1915 210 1935
rect 230 1915 235 1935
rect 205 1885 235 1915
rect 205 1865 210 1885
rect 230 1865 235 1885
rect 205 1835 235 1865
rect 205 1815 210 1835
rect 230 1815 235 1835
rect 205 1785 235 1815
rect 205 1765 210 1785
rect 230 1765 235 1785
rect 205 1755 235 1765
rect 265 2085 295 2095
rect 265 2065 270 2085
rect 290 2065 295 2085
rect 265 2035 295 2065
rect 265 2015 270 2035
rect 290 2015 295 2035
rect 265 1985 295 2015
rect 265 1965 270 1985
rect 290 1965 295 1985
rect 265 1935 295 1965
rect 265 1915 270 1935
rect 290 1915 295 1935
rect 265 1885 295 1915
rect 265 1865 270 1885
rect 290 1865 295 1885
rect 265 1835 295 1865
rect 265 1815 270 1835
rect 290 1815 295 1835
rect 265 1785 295 1815
rect 265 1765 270 1785
rect 290 1765 295 1785
rect 265 1755 295 1765
rect 325 2085 355 2095
rect 325 2065 330 2085
rect 350 2065 355 2085
rect 325 2035 355 2065
rect 325 2015 330 2035
rect 350 2015 355 2035
rect 325 1985 355 2015
rect 325 1965 330 1985
rect 350 1965 355 1985
rect 325 1935 355 1965
rect 325 1915 330 1935
rect 350 1915 355 1935
rect 325 1885 355 1915
rect 325 1865 330 1885
rect 350 1865 355 1885
rect 325 1835 355 1865
rect 325 1815 330 1835
rect 350 1815 355 1835
rect 325 1785 355 1815
rect 325 1765 330 1785
rect 350 1765 355 1785
rect 325 1755 355 1765
rect 385 2085 415 2095
rect 385 2065 390 2085
rect 410 2065 415 2085
rect 385 2035 415 2065
rect 385 2015 390 2035
rect 410 2015 415 2035
rect 385 1985 415 2015
rect 385 1965 390 1985
rect 410 1965 415 1985
rect 385 1935 415 1965
rect 385 1915 390 1935
rect 410 1915 415 1935
rect 385 1885 415 1915
rect 385 1865 390 1885
rect 410 1865 415 1885
rect 385 1835 415 1865
rect 385 1815 390 1835
rect 410 1815 415 1835
rect 385 1785 415 1815
rect 385 1765 390 1785
rect 410 1765 415 1785
rect 385 1755 415 1765
rect 445 2085 475 2095
rect 445 2065 450 2085
rect 470 2065 475 2085
rect 445 2035 475 2065
rect 445 2015 450 2035
rect 470 2015 475 2035
rect 445 1985 475 2015
rect 445 1965 450 1985
rect 470 1965 475 1985
rect 445 1935 475 1965
rect 445 1915 450 1935
rect 470 1915 475 1935
rect 445 1885 475 1915
rect 445 1865 450 1885
rect 470 1865 475 1885
rect 445 1835 475 1865
rect 445 1815 450 1835
rect 470 1815 475 1835
rect 445 1785 475 1815
rect 445 1765 450 1785
rect 470 1765 475 1785
rect 445 1755 475 1765
rect 505 2085 535 2095
rect 505 2065 510 2085
rect 530 2065 535 2085
rect 505 2035 535 2065
rect 505 2015 510 2035
rect 530 2015 535 2035
rect 505 1985 535 2015
rect 505 1965 510 1985
rect 530 1965 535 1985
rect 505 1935 535 1965
rect 505 1915 510 1935
rect 530 1915 535 1935
rect 505 1885 535 1915
rect 505 1865 510 1885
rect 530 1865 535 1885
rect 505 1835 535 1865
rect 505 1815 510 1835
rect 530 1815 535 1835
rect 505 1785 535 1815
rect 505 1765 510 1785
rect 530 1765 535 1785
rect 505 1755 535 1765
rect 565 2085 595 2095
rect 565 2065 570 2085
rect 590 2065 595 2085
rect 565 2035 595 2065
rect 565 2015 570 2035
rect 590 2015 595 2035
rect 565 1985 595 2015
rect 565 1965 570 1985
rect 590 1965 595 1985
rect 565 1935 595 1965
rect 565 1915 570 1935
rect 590 1915 595 1935
rect 565 1885 595 1915
rect 565 1865 570 1885
rect 590 1865 595 1885
rect 565 1835 595 1865
rect 565 1815 570 1835
rect 590 1815 595 1835
rect 565 1785 595 1815
rect 565 1765 570 1785
rect 590 1765 595 1785
rect 565 1755 595 1765
rect 625 2085 655 2095
rect 625 2065 630 2085
rect 650 2065 655 2085
rect 625 2035 655 2065
rect 625 2015 630 2035
rect 650 2015 655 2035
rect 625 1985 655 2015
rect 625 1965 630 1985
rect 650 1965 655 1985
rect 625 1935 655 1965
rect 625 1915 630 1935
rect 650 1915 655 1935
rect 625 1885 655 1915
rect 625 1865 630 1885
rect 650 1865 655 1885
rect 625 1835 655 1865
rect 625 1815 630 1835
rect 650 1815 655 1835
rect 625 1785 655 1815
rect 625 1765 630 1785
rect 650 1765 655 1785
rect 625 1755 655 1765
rect 685 2085 755 2095
rect 685 2065 690 2085
rect 710 2065 730 2085
rect 750 2065 755 2085
rect 685 2035 755 2065
rect 685 2015 690 2035
rect 710 2015 730 2035
rect 750 2015 755 2035
rect 685 1985 755 2015
rect 685 1965 690 1985
rect 710 1965 730 1985
rect 750 1965 755 1985
rect 685 1935 755 1965
rect 685 1915 690 1935
rect 710 1915 730 1935
rect 750 1915 755 1935
rect 685 1885 755 1915
rect 685 1865 690 1885
rect 710 1865 730 1885
rect 750 1865 755 1885
rect 685 1835 755 1865
rect 685 1815 690 1835
rect 710 1815 730 1835
rect 750 1815 755 1835
rect 685 1785 755 1815
rect 685 1765 690 1785
rect 710 1765 730 1785
rect 750 1765 755 1785
rect 685 1755 755 1765
rect 935 2085 1005 2095
rect 935 2065 940 2085
rect 960 2065 980 2085
rect 1000 2065 1005 2085
rect 935 2035 1005 2065
rect 935 2015 940 2035
rect 960 2015 980 2035
rect 1000 2015 1005 2035
rect 935 1985 1005 2015
rect 935 1965 940 1985
rect 960 1965 980 1985
rect 1000 1965 1005 1985
rect 935 1935 1005 1965
rect 935 1915 940 1935
rect 960 1915 980 1935
rect 1000 1915 1005 1935
rect 935 1885 1005 1915
rect 935 1865 940 1885
rect 960 1865 980 1885
rect 1000 1865 1005 1885
rect 935 1835 1005 1865
rect 935 1815 940 1835
rect 960 1815 980 1835
rect 1000 1815 1005 1835
rect 935 1785 1005 1815
rect 935 1765 940 1785
rect 960 1765 980 1785
rect 1000 1765 1005 1785
rect 935 1755 1005 1765
rect 1035 2085 1065 2095
rect 1035 2065 1040 2085
rect 1060 2065 1065 2085
rect 1035 2035 1065 2065
rect 1035 2015 1040 2035
rect 1060 2015 1065 2035
rect 1035 1985 1065 2015
rect 1035 1965 1040 1985
rect 1060 1965 1065 1985
rect 1035 1935 1065 1965
rect 1035 1915 1040 1935
rect 1060 1915 1065 1935
rect 1035 1885 1065 1915
rect 1035 1865 1040 1885
rect 1060 1865 1065 1885
rect 1035 1835 1065 1865
rect 1035 1815 1040 1835
rect 1060 1815 1065 1835
rect 1035 1785 1065 1815
rect 1035 1765 1040 1785
rect 1060 1765 1065 1785
rect 1035 1755 1065 1765
rect 1095 2085 1125 2095
rect 1095 2065 1100 2085
rect 1120 2065 1125 2085
rect 1095 2035 1125 2065
rect 1095 2015 1100 2035
rect 1120 2015 1125 2035
rect 1095 1985 1125 2015
rect 1095 1965 1100 1985
rect 1120 1965 1125 1985
rect 1095 1935 1125 1965
rect 1095 1915 1100 1935
rect 1120 1915 1125 1935
rect 1095 1885 1125 1915
rect 1095 1865 1100 1885
rect 1120 1865 1125 1885
rect 1095 1835 1125 1865
rect 1095 1815 1100 1835
rect 1120 1815 1125 1835
rect 1095 1785 1125 1815
rect 1095 1765 1100 1785
rect 1120 1765 1125 1785
rect 1095 1755 1125 1765
rect 1155 2085 1185 2095
rect 1155 2065 1160 2085
rect 1180 2065 1185 2085
rect 1155 2035 1185 2065
rect 1155 2015 1160 2035
rect 1180 2015 1185 2035
rect 1155 1985 1185 2015
rect 1155 1965 1160 1985
rect 1180 1965 1185 1985
rect 1155 1935 1185 1965
rect 1155 1915 1160 1935
rect 1180 1915 1185 1935
rect 1155 1885 1185 1915
rect 1155 1865 1160 1885
rect 1180 1865 1185 1885
rect 1155 1835 1185 1865
rect 1155 1815 1160 1835
rect 1180 1815 1185 1835
rect 1155 1785 1185 1815
rect 1155 1765 1160 1785
rect 1180 1765 1185 1785
rect 1155 1755 1185 1765
rect 1215 2085 1245 2095
rect 1215 2065 1220 2085
rect 1240 2065 1245 2085
rect 1215 2035 1245 2065
rect 1215 2015 1220 2035
rect 1240 2015 1245 2035
rect 1215 1985 1245 2015
rect 1215 1965 1220 1985
rect 1240 1965 1245 1985
rect 1215 1935 1245 1965
rect 1215 1915 1220 1935
rect 1240 1915 1245 1935
rect 1215 1885 1245 1915
rect 1215 1865 1220 1885
rect 1240 1865 1245 1885
rect 1215 1835 1245 1865
rect 1215 1815 1220 1835
rect 1240 1815 1245 1835
rect 1215 1785 1245 1815
rect 1215 1765 1220 1785
rect 1240 1765 1245 1785
rect 1215 1755 1245 1765
rect 1275 2085 1305 2095
rect 1275 2065 1280 2085
rect 1300 2065 1305 2085
rect 1275 2035 1305 2065
rect 1275 2015 1280 2035
rect 1300 2015 1305 2035
rect 1275 1985 1305 2015
rect 1275 1965 1280 1985
rect 1300 1965 1305 1985
rect 1275 1935 1305 1965
rect 1275 1915 1280 1935
rect 1300 1915 1305 1935
rect 1275 1885 1305 1915
rect 1275 1865 1280 1885
rect 1300 1865 1305 1885
rect 1275 1835 1305 1865
rect 1275 1815 1280 1835
rect 1300 1815 1305 1835
rect 1275 1785 1305 1815
rect 1275 1765 1280 1785
rect 1300 1765 1305 1785
rect 1275 1755 1305 1765
rect 1335 2085 1365 2095
rect 1335 2065 1340 2085
rect 1360 2065 1365 2085
rect 1335 2035 1365 2065
rect 1335 2015 1340 2035
rect 1360 2015 1365 2035
rect 1335 1985 1365 2015
rect 1335 1965 1340 1985
rect 1360 1965 1365 1985
rect 1335 1935 1365 1965
rect 1335 1915 1340 1935
rect 1360 1915 1365 1935
rect 1335 1885 1365 1915
rect 1335 1865 1340 1885
rect 1360 1865 1365 1885
rect 1335 1835 1365 1865
rect 1335 1815 1340 1835
rect 1360 1815 1365 1835
rect 1335 1785 1365 1815
rect 1335 1765 1340 1785
rect 1360 1765 1365 1785
rect 1335 1755 1365 1765
rect 1395 2085 1425 2095
rect 1395 2065 1400 2085
rect 1420 2065 1425 2085
rect 1395 2035 1425 2065
rect 1395 2015 1400 2035
rect 1420 2015 1425 2035
rect 1395 1985 1425 2015
rect 1395 1965 1400 1985
rect 1420 1965 1425 1985
rect 1395 1935 1425 1965
rect 1395 1915 1400 1935
rect 1420 1915 1425 1935
rect 1395 1885 1425 1915
rect 1395 1865 1400 1885
rect 1420 1865 1425 1885
rect 1395 1835 1425 1865
rect 1395 1815 1400 1835
rect 1420 1815 1425 1835
rect 1395 1785 1425 1815
rect 1395 1765 1400 1785
rect 1420 1765 1425 1785
rect 1395 1755 1425 1765
rect 1455 2085 1485 2095
rect 1455 2065 1460 2085
rect 1480 2065 1485 2085
rect 1455 2035 1485 2065
rect 1455 2015 1460 2035
rect 1480 2015 1485 2035
rect 1455 1985 1485 2015
rect 1455 1965 1460 1985
rect 1480 1965 1485 1985
rect 1455 1935 1485 1965
rect 1455 1915 1460 1935
rect 1480 1915 1485 1935
rect 1455 1885 1485 1915
rect 1455 1865 1460 1885
rect 1480 1865 1485 1885
rect 1455 1835 1485 1865
rect 1455 1815 1460 1835
rect 1480 1815 1485 1835
rect 1455 1785 1485 1815
rect 1455 1765 1460 1785
rect 1480 1765 1485 1785
rect 1455 1755 1485 1765
rect 1515 2085 1545 2095
rect 1515 2065 1520 2085
rect 1540 2065 1545 2085
rect 1515 2035 1545 2065
rect 1515 2015 1520 2035
rect 1540 2015 1545 2035
rect 1515 1985 1545 2015
rect 1515 1965 1520 1985
rect 1540 1965 1545 1985
rect 1515 1935 1545 1965
rect 1515 1915 1520 1935
rect 1540 1915 1545 1935
rect 1515 1885 1545 1915
rect 1515 1865 1520 1885
rect 1540 1865 1545 1885
rect 1515 1835 1545 1865
rect 1515 1815 1520 1835
rect 1540 1815 1545 1835
rect 1515 1785 1545 1815
rect 1515 1765 1520 1785
rect 1540 1765 1545 1785
rect 1515 1755 1545 1765
rect 1575 2085 1605 2095
rect 1575 2065 1580 2085
rect 1600 2065 1605 2085
rect 1575 2035 1605 2065
rect 1575 2015 1580 2035
rect 1600 2015 1605 2035
rect 1575 1985 1605 2015
rect 1575 1965 1580 1985
rect 1600 1965 1605 1985
rect 1575 1935 1605 1965
rect 1575 1915 1580 1935
rect 1600 1915 1605 1935
rect 1575 1885 1605 1915
rect 1575 1865 1580 1885
rect 1600 1865 1605 1885
rect 1575 1835 1605 1865
rect 1575 1815 1580 1835
rect 1600 1815 1605 1835
rect 1575 1785 1605 1815
rect 1575 1765 1580 1785
rect 1600 1765 1605 1785
rect 1575 1755 1605 1765
rect 1635 2085 1665 2095
rect 1635 2065 1640 2085
rect 1660 2065 1665 2085
rect 1635 2035 1665 2065
rect 1635 2015 1640 2035
rect 1660 2015 1665 2035
rect 1635 1985 1665 2015
rect 1635 1965 1640 1985
rect 1660 1965 1665 1985
rect 1635 1935 1665 1965
rect 1635 1915 1640 1935
rect 1660 1915 1665 1935
rect 1635 1885 1665 1915
rect 1635 1865 1640 1885
rect 1660 1865 1665 1885
rect 1635 1835 1665 1865
rect 1635 1815 1640 1835
rect 1660 1815 1665 1835
rect 1635 1785 1665 1815
rect 1635 1765 1640 1785
rect 1660 1765 1665 1785
rect 1635 1755 1665 1765
rect 1695 2085 1765 2095
rect 1695 2065 1700 2085
rect 1720 2065 1740 2085
rect 1760 2065 1765 2085
rect 1695 2035 1765 2065
rect 1695 2015 1700 2035
rect 1720 2015 1740 2035
rect 1760 2015 1765 2035
rect 1695 1985 1765 2015
rect 1695 1965 1700 1985
rect 1720 1965 1740 1985
rect 1760 1965 1765 1985
rect 1695 1935 1765 1965
rect 1695 1915 1700 1935
rect 1720 1915 1740 1935
rect 1760 1915 1765 1935
rect 1695 1885 1765 1915
rect 1695 1865 1700 1885
rect 1720 1865 1740 1885
rect 1760 1865 1765 1885
rect 1695 1835 1765 1865
rect 1695 1815 1700 1835
rect 1720 1815 1740 1835
rect 1760 1815 1765 1835
rect 1695 1785 1765 1815
rect 1695 1765 1700 1785
rect 1720 1765 1740 1785
rect 1760 1765 1765 1785
rect 1695 1755 1765 1765
rect 2060 2085 2130 2095
rect 2060 2065 2065 2085
rect 2085 2065 2105 2085
rect 2125 2065 2130 2085
rect 2060 2035 2130 2065
rect 2060 2015 2065 2035
rect 2085 2015 2105 2035
rect 2125 2015 2130 2035
rect 2060 1985 2130 2015
rect 2060 1965 2065 1985
rect 2085 1965 2105 1985
rect 2125 1965 2130 1985
rect 2060 1935 2130 1965
rect 2060 1915 2065 1935
rect 2085 1915 2105 1935
rect 2125 1915 2130 1935
rect 2060 1885 2130 1915
rect 2060 1865 2065 1885
rect 2085 1865 2105 1885
rect 2125 1865 2130 1885
rect 2060 1835 2130 1865
rect 2060 1815 2065 1835
rect 2085 1815 2105 1835
rect 2125 1815 2130 1835
rect 2060 1785 2130 1815
rect 2060 1765 2065 1785
rect 2085 1765 2105 1785
rect 2125 1765 2130 1785
rect 2060 1755 2130 1765
rect 2160 2085 2190 2095
rect 2160 2065 2165 2085
rect 2185 2065 2190 2085
rect 2160 2035 2190 2065
rect 2160 2015 2165 2035
rect 2185 2015 2190 2035
rect 2160 1985 2190 2015
rect 2160 1965 2165 1985
rect 2185 1965 2190 1985
rect 2160 1935 2190 1965
rect 2160 1915 2165 1935
rect 2185 1915 2190 1935
rect 2160 1885 2190 1915
rect 2160 1865 2165 1885
rect 2185 1865 2190 1885
rect 2160 1835 2190 1865
rect 2160 1815 2165 1835
rect 2185 1815 2190 1835
rect 2160 1785 2190 1815
rect 2160 1765 2165 1785
rect 2185 1765 2190 1785
rect 2160 1755 2190 1765
rect 2220 2085 2250 2095
rect 2220 2065 2225 2085
rect 2245 2065 2250 2085
rect 2220 2035 2250 2065
rect 2220 2015 2225 2035
rect 2245 2015 2250 2035
rect 2220 1985 2250 2015
rect 2220 1965 2225 1985
rect 2245 1965 2250 1985
rect 2220 1935 2250 1965
rect 2220 1915 2225 1935
rect 2245 1915 2250 1935
rect 2220 1885 2250 1915
rect 2220 1865 2225 1885
rect 2245 1865 2250 1885
rect 2220 1835 2250 1865
rect 2220 1815 2225 1835
rect 2245 1815 2250 1835
rect 2220 1785 2250 1815
rect 2220 1765 2225 1785
rect 2245 1765 2250 1785
rect 2220 1755 2250 1765
rect 2280 2085 2310 2095
rect 2280 2065 2285 2085
rect 2305 2065 2310 2085
rect 2280 2035 2310 2065
rect 2280 2015 2285 2035
rect 2305 2015 2310 2035
rect 2280 1985 2310 2015
rect 2280 1965 2285 1985
rect 2305 1965 2310 1985
rect 2280 1935 2310 1965
rect 2280 1915 2285 1935
rect 2305 1915 2310 1935
rect 2280 1885 2310 1915
rect 2280 1865 2285 1885
rect 2305 1865 2310 1885
rect 2280 1835 2310 1865
rect 2280 1815 2285 1835
rect 2305 1815 2310 1835
rect 2280 1785 2310 1815
rect 2280 1765 2285 1785
rect 2305 1765 2310 1785
rect 2280 1755 2310 1765
rect 2340 2085 2370 2095
rect 2340 2065 2345 2085
rect 2365 2065 2370 2085
rect 2340 2035 2370 2065
rect 2340 2015 2345 2035
rect 2365 2015 2370 2035
rect 2340 1985 2370 2015
rect 2340 1965 2345 1985
rect 2365 1965 2370 1985
rect 2340 1935 2370 1965
rect 2340 1915 2345 1935
rect 2365 1915 2370 1935
rect 2340 1885 2370 1915
rect 2340 1865 2345 1885
rect 2365 1865 2370 1885
rect 2340 1835 2370 1865
rect 2340 1815 2345 1835
rect 2365 1815 2370 1835
rect 2340 1785 2370 1815
rect 2340 1765 2345 1785
rect 2365 1765 2370 1785
rect 2340 1755 2370 1765
rect 2400 2085 2430 2095
rect 2400 2065 2405 2085
rect 2425 2065 2430 2085
rect 2400 2035 2430 2065
rect 2400 2015 2405 2035
rect 2425 2015 2430 2035
rect 2400 1985 2430 2015
rect 2400 1965 2405 1985
rect 2425 1965 2430 1985
rect 2400 1935 2430 1965
rect 2400 1915 2405 1935
rect 2425 1915 2430 1935
rect 2400 1885 2430 1915
rect 2400 1865 2405 1885
rect 2425 1865 2430 1885
rect 2400 1835 2430 1865
rect 2400 1815 2405 1835
rect 2425 1815 2430 1835
rect 2400 1785 2430 1815
rect 2400 1765 2405 1785
rect 2425 1765 2430 1785
rect 2400 1755 2430 1765
rect 2460 2085 2490 2095
rect 2460 2065 2465 2085
rect 2485 2065 2490 2085
rect 2460 2035 2490 2065
rect 2460 2015 2465 2035
rect 2485 2015 2490 2035
rect 2460 1985 2490 2015
rect 2460 1965 2465 1985
rect 2485 1965 2490 1985
rect 2460 1935 2490 1965
rect 2460 1915 2465 1935
rect 2485 1915 2490 1935
rect 2460 1885 2490 1915
rect 2460 1865 2465 1885
rect 2485 1865 2490 1885
rect 2460 1835 2490 1865
rect 2460 1815 2465 1835
rect 2485 1815 2490 1835
rect 2460 1785 2490 1815
rect 2460 1765 2465 1785
rect 2485 1765 2490 1785
rect 2460 1755 2490 1765
rect 2520 2085 2550 2095
rect 2520 2065 2525 2085
rect 2545 2065 2550 2085
rect 2520 2035 2550 2065
rect 2520 2015 2525 2035
rect 2545 2015 2550 2035
rect 2520 1985 2550 2015
rect 2520 1965 2525 1985
rect 2545 1965 2550 1985
rect 2520 1935 2550 1965
rect 2520 1915 2525 1935
rect 2545 1915 2550 1935
rect 2520 1885 2550 1915
rect 2520 1865 2525 1885
rect 2545 1865 2550 1885
rect 2520 1835 2550 1865
rect 2520 1815 2525 1835
rect 2545 1815 2550 1835
rect 2520 1785 2550 1815
rect 2520 1765 2525 1785
rect 2545 1765 2550 1785
rect 2520 1755 2550 1765
rect 2580 2085 2610 2095
rect 2580 2065 2585 2085
rect 2605 2065 2610 2085
rect 2580 2035 2610 2065
rect 2580 2015 2585 2035
rect 2605 2015 2610 2035
rect 2580 1985 2610 2015
rect 2580 1965 2585 1985
rect 2605 1965 2610 1985
rect 2580 1935 2610 1965
rect 2580 1915 2585 1935
rect 2605 1915 2610 1935
rect 2580 1885 2610 1915
rect 2580 1865 2585 1885
rect 2605 1865 2610 1885
rect 2580 1835 2610 1865
rect 2580 1815 2585 1835
rect 2605 1815 2610 1835
rect 2580 1785 2610 1815
rect 2580 1765 2585 1785
rect 2605 1765 2610 1785
rect 2580 1755 2610 1765
rect 2640 2085 2670 2095
rect 2640 2065 2645 2085
rect 2665 2065 2670 2085
rect 2640 2035 2670 2065
rect 2640 2015 2645 2035
rect 2665 2015 2670 2035
rect 2640 1985 2670 2015
rect 2640 1965 2645 1985
rect 2665 1965 2670 1985
rect 2640 1935 2670 1965
rect 2640 1915 2645 1935
rect 2665 1915 2670 1935
rect 2640 1885 2670 1915
rect 2640 1865 2645 1885
rect 2665 1865 2670 1885
rect 2640 1835 2670 1865
rect 2640 1815 2645 1835
rect 2665 1815 2670 1835
rect 2640 1785 2670 1815
rect 2640 1765 2645 1785
rect 2665 1765 2670 1785
rect 2640 1755 2670 1765
rect 2700 2085 2730 2095
rect 2700 2065 2705 2085
rect 2725 2065 2730 2085
rect 2700 2035 2730 2065
rect 2700 2015 2705 2035
rect 2725 2015 2730 2035
rect 2700 1985 2730 2015
rect 2700 1965 2705 1985
rect 2725 1965 2730 1985
rect 2700 1935 2730 1965
rect 2700 1915 2705 1935
rect 2725 1915 2730 1935
rect 2700 1885 2730 1915
rect 2700 1865 2705 1885
rect 2725 1865 2730 1885
rect 2700 1835 2730 1865
rect 2700 1815 2705 1835
rect 2725 1815 2730 1835
rect 2700 1785 2730 1815
rect 2700 1765 2705 1785
rect 2725 1765 2730 1785
rect 2700 1755 2730 1765
rect 2760 2085 2790 2095
rect 2760 2065 2765 2085
rect 2785 2065 2790 2085
rect 2760 2035 2790 2065
rect 2760 2015 2765 2035
rect 2785 2015 2790 2035
rect 2760 1985 2790 2015
rect 2760 1965 2765 1985
rect 2785 1965 2790 1985
rect 2760 1935 2790 1965
rect 2760 1915 2765 1935
rect 2785 1915 2790 1935
rect 2760 1885 2790 1915
rect 2760 1865 2765 1885
rect 2785 1865 2790 1885
rect 2760 1835 2790 1865
rect 2760 1815 2765 1835
rect 2785 1815 2790 1835
rect 2760 1785 2790 1815
rect 2760 1765 2765 1785
rect 2785 1765 2790 1785
rect 2760 1755 2790 1765
rect 2820 2085 2890 2095
rect 2820 2065 2825 2085
rect 2845 2065 2865 2085
rect 2885 2065 2890 2085
rect 2820 2035 2890 2065
rect 2820 2015 2825 2035
rect 2845 2015 2865 2035
rect 2885 2015 2890 2035
rect 2820 1985 2890 2015
rect 2820 1965 2825 1985
rect 2845 1965 2865 1985
rect 2885 1965 2890 1985
rect 2820 1935 2890 1965
rect 2820 1915 2825 1935
rect 2845 1915 2865 1935
rect 2885 1915 2890 1935
rect 2820 1885 2890 1915
rect 2820 1865 2825 1885
rect 2845 1865 2865 1885
rect 2885 1865 2890 1885
rect 2820 1835 2890 1865
rect 2820 1815 2825 1835
rect 2845 1815 2865 1835
rect 2885 1815 2890 1835
rect 2820 1785 2890 1815
rect 2820 1765 2825 1785
rect 2845 1765 2865 1785
rect 2885 1765 2890 1785
rect 2820 1755 2890 1765
rect -1095 1730 -1075 1755
rect -975 1730 -955 1755
rect -855 1730 -835 1755
rect -735 1730 -715 1755
rect -615 1730 -595 1755
rect -495 1730 -475 1755
rect 30 1730 50 1755
rect 150 1730 170 1755
rect 270 1730 290 1755
rect 390 1730 410 1755
rect 510 1730 530 1755
rect 630 1730 650 1755
rect 1040 1730 1060 1755
rect 1160 1730 1180 1755
rect 1280 1730 1300 1755
rect 1400 1730 1420 1755
rect 1520 1730 1540 1755
rect 1640 1730 1660 1755
rect 2165 1730 2185 1755
rect 2285 1730 2305 1755
rect 2405 1730 2425 1755
rect 2525 1730 2545 1755
rect 2645 1730 2665 1755
rect 2765 1730 2785 1755
rect -1105 1720 -1065 1730
rect -1105 1700 -1095 1720
rect -1075 1700 -1065 1720
rect -1105 1690 -1065 1700
rect -985 1720 -945 1730
rect -985 1700 -975 1720
rect -955 1700 -945 1720
rect -985 1690 -945 1700
rect -865 1720 -825 1730
rect -865 1700 -855 1720
rect -835 1700 -825 1720
rect -865 1690 -825 1700
rect -800 1720 -770 1730
rect -800 1700 -795 1720
rect -775 1700 -770 1720
rect -800 1690 -770 1700
rect -745 1720 -705 1730
rect -745 1700 -735 1720
rect -715 1700 -705 1720
rect -745 1690 -705 1700
rect -625 1720 -585 1730
rect -625 1700 -615 1720
rect -595 1700 -585 1720
rect -625 1690 -585 1700
rect -505 1720 -465 1730
rect -505 1700 -495 1720
rect -475 1700 -465 1720
rect -505 1690 -465 1700
rect 20 1720 60 1730
rect 20 1700 30 1720
rect 50 1700 60 1720
rect 20 1690 60 1700
rect 140 1720 180 1730
rect 140 1700 150 1720
rect 170 1700 180 1720
rect 140 1690 180 1700
rect 260 1720 300 1730
rect 260 1700 270 1720
rect 290 1700 300 1720
rect 260 1690 300 1700
rect 325 1720 355 1730
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 380 1720 420 1730
rect 380 1700 390 1720
rect 410 1700 420 1720
rect 380 1690 420 1700
rect 500 1720 540 1730
rect 500 1700 510 1720
rect 530 1700 540 1720
rect 500 1690 540 1700
rect 620 1720 660 1730
rect 620 1700 630 1720
rect 650 1700 660 1720
rect 620 1690 660 1700
rect 1030 1720 1070 1730
rect 1030 1700 1040 1720
rect 1060 1700 1070 1720
rect 1030 1690 1070 1700
rect 1150 1720 1190 1730
rect 1150 1700 1160 1720
rect 1180 1700 1190 1720
rect 1150 1690 1190 1700
rect 1270 1720 1310 1730
rect 1270 1700 1280 1720
rect 1300 1700 1310 1720
rect 1270 1690 1310 1700
rect 1335 1720 1365 1730
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 1390 1720 1430 1730
rect 1390 1700 1400 1720
rect 1420 1700 1430 1720
rect 1390 1690 1430 1700
rect 1510 1720 1550 1730
rect 1510 1700 1520 1720
rect 1540 1700 1550 1720
rect 1510 1690 1550 1700
rect 1630 1720 1670 1730
rect 1630 1700 1640 1720
rect 1660 1700 1670 1720
rect 1630 1690 1670 1700
rect 2155 1720 2195 1730
rect 2155 1700 2165 1720
rect 2185 1700 2195 1720
rect 2155 1690 2195 1700
rect 2275 1720 2315 1730
rect 2275 1700 2285 1720
rect 2305 1700 2315 1720
rect 2275 1690 2315 1700
rect 2395 1720 2435 1730
rect 2395 1700 2405 1720
rect 2425 1700 2435 1720
rect 2395 1690 2435 1700
rect 2460 1720 2490 1730
rect 2460 1700 2465 1720
rect 2485 1700 2490 1720
rect 2460 1690 2490 1700
rect 2515 1720 2555 1730
rect 2515 1700 2525 1720
rect 2545 1700 2555 1720
rect 2515 1690 2555 1700
rect 2635 1720 2675 1730
rect 2635 1700 2645 1720
rect 2665 1700 2675 1720
rect 2635 1690 2675 1700
rect 2755 1720 2795 1730
rect 2755 1700 2765 1720
rect 2785 1700 2795 1720
rect 2755 1690 2795 1700
rect 455 1575 495 1585
rect 455 1555 465 1575
rect 485 1555 495 1575
rect 455 1545 495 1555
rect 625 1575 655 1585
rect 625 1555 630 1575
rect 650 1555 655 1575
rect 625 1545 655 1555
rect 785 1575 825 1585
rect 785 1555 795 1575
rect 815 1555 825 1575
rect 785 1545 825 1555
rect 865 1575 905 1585
rect 865 1555 875 1575
rect 895 1555 905 1575
rect 865 1545 905 1555
rect 1035 1575 1065 1585
rect 1035 1555 1040 1575
rect 1060 1555 1065 1575
rect 1035 1545 1065 1555
rect 1195 1575 1235 1585
rect 1195 1555 1205 1575
rect 1225 1555 1235 1575
rect 1195 1545 1235 1555
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1460 -1095 1480
rect -1135 1450 -1095 1460
rect -1025 1480 -985 1490
rect -1025 1460 -1015 1480
rect -995 1460 -985 1480
rect -1025 1450 -985 1460
rect -915 1480 -875 1490
rect -915 1460 -905 1480
rect -885 1460 -875 1480
rect -915 1450 -875 1460
rect -805 1480 -765 1490
rect -805 1460 -795 1480
rect -775 1460 -765 1480
rect -805 1450 -765 1460
rect -695 1480 -655 1490
rect -695 1460 -685 1480
rect -665 1460 -655 1480
rect -695 1450 -655 1460
rect -585 1480 -545 1490
rect -585 1460 -575 1480
rect -555 1460 -545 1480
rect -585 1450 -545 1460
rect -475 1480 -435 1490
rect 465 1480 485 1545
rect 565 1530 605 1540
rect 565 1510 575 1530
rect 595 1510 605 1530
rect 565 1500 605 1510
rect 575 1480 595 1500
rect 630 1480 650 1545
rect 675 1530 715 1540
rect 675 1510 685 1530
rect 705 1510 715 1530
rect 675 1500 715 1510
rect 685 1480 705 1500
rect 795 1480 815 1545
rect 875 1480 895 1545
rect 975 1530 1015 1540
rect 975 1510 985 1530
rect 1005 1510 1015 1530
rect 975 1500 1015 1510
rect 985 1480 1005 1500
rect 1040 1480 1060 1545
rect 1085 1530 1125 1540
rect 1085 1510 1095 1530
rect 1115 1510 1125 1530
rect 1085 1500 1125 1510
rect 1095 1480 1115 1500
rect 1205 1480 1225 1545
rect 2125 1480 2165 1490
rect -475 1460 -465 1480
rect -445 1460 -435 1480
rect -475 1450 -435 1460
rect 420 1470 490 1480
rect 420 1450 425 1470
rect 445 1450 465 1470
rect 485 1450 490 1470
rect -1125 1430 -1105 1450
rect -1015 1430 -995 1450
rect -905 1430 -885 1450
rect -795 1430 -775 1450
rect -685 1430 -665 1450
rect -575 1430 -555 1450
rect -465 1430 -445 1450
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1170 1420 -1100 1430
rect -1170 1400 -1165 1420
rect -1145 1400 -1125 1420
rect -1105 1400 -1100 1420
rect -1170 1370 -1100 1400
rect -1170 1350 -1165 1370
rect -1145 1350 -1125 1370
rect -1105 1350 -1100 1370
rect -1170 1320 -1100 1350
rect -1170 1300 -1165 1320
rect -1145 1300 -1125 1320
rect -1105 1300 -1100 1320
rect -1170 1270 -1100 1300
rect -1170 1250 -1165 1270
rect -1145 1250 -1125 1270
rect -1105 1250 -1100 1270
rect -1170 1220 -1100 1250
rect -1170 1200 -1165 1220
rect -1145 1200 -1125 1220
rect -1105 1200 -1100 1220
rect -1170 1170 -1100 1200
rect -1170 1150 -1165 1170
rect -1145 1150 -1125 1170
rect -1105 1150 -1100 1170
rect -1170 1120 -1100 1150
rect -1170 1100 -1165 1120
rect -1145 1100 -1125 1120
rect -1105 1100 -1100 1120
rect -1170 1070 -1100 1100
rect -1170 1050 -1165 1070
rect -1145 1050 -1125 1070
rect -1105 1050 -1100 1070
rect -1170 1020 -1100 1050
rect -1170 1000 -1165 1020
rect -1145 1000 -1125 1020
rect -1105 1000 -1100 1020
rect -1170 970 -1100 1000
rect -1170 950 -1165 970
rect -1145 950 -1125 970
rect -1105 950 -1100 970
rect -1170 920 -1100 950
rect -1170 900 -1165 920
rect -1145 900 -1125 920
rect -1105 900 -1100 920
rect -1170 870 -1100 900
rect -1170 850 -1165 870
rect -1145 850 -1125 870
rect -1105 850 -1100 870
rect -1170 840 -1100 850
rect -1075 1420 -1045 1430
rect -1075 1400 -1070 1420
rect -1050 1400 -1045 1420
rect -1075 1370 -1045 1400
rect -1075 1350 -1070 1370
rect -1050 1350 -1045 1370
rect -1075 1320 -1045 1350
rect -1075 1300 -1070 1320
rect -1050 1300 -1045 1320
rect -1075 1270 -1045 1300
rect -1075 1250 -1070 1270
rect -1050 1250 -1045 1270
rect -1075 1220 -1045 1250
rect -1075 1200 -1070 1220
rect -1050 1200 -1045 1220
rect -1075 1170 -1045 1200
rect -1075 1150 -1070 1170
rect -1050 1150 -1045 1170
rect -1075 1120 -1045 1150
rect -1075 1100 -1070 1120
rect -1050 1100 -1045 1120
rect -1075 1070 -1045 1100
rect -1075 1050 -1070 1070
rect -1050 1050 -1045 1070
rect -1075 1020 -1045 1050
rect -1075 1000 -1070 1020
rect -1050 1000 -1045 1020
rect -1075 970 -1045 1000
rect -1075 950 -1070 970
rect -1050 950 -1045 970
rect -1075 920 -1045 950
rect -1075 900 -1070 920
rect -1050 900 -1045 920
rect -1075 870 -1045 900
rect -1075 850 -1070 870
rect -1050 850 -1045 870
rect -1075 840 -1045 850
rect -1020 1420 -990 1430
rect -1020 1400 -1015 1420
rect -995 1400 -990 1420
rect -1020 1370 -990 1400
rect -1020 1350 -1015 1370
rect -995 1350 -990 1370
rect -1020 1320 -990 1350
rect -1020 1300 -1015 1320
rect -995 1300 -990 1320
rect -1020 1270 -990 1300
rect -1020 1250 -1015 1270
rect -995 1250 -990 1270
rect -1020 1220 -990 1250
rect -1020 1200 -1015 1220
rect -995 1200 -990 1220
rect -1020 1170 -990 1200
rect -1020 1150 -1015 1170
rect -995 1150 -990 1170
rect -1020 1120 -990 1150
rect -1020 1100 -1015 1120
rect -995 1100 -990 1120
rect -1020 1070 -990 1100
rect -1020 1050 -1015 1070
rect -995 1050 -990 1070
rect -1020 1020 -990 1050
rect -1020 1000 -1015 1020
rect -995 1000 -990 1020
rect -1020 970 -990 1000
rect -1020 950 -1015 970
rect -995 950 -990 970
rect -1020 920 -990 950
rect -1020 900 -1015 920
rect -995 900 -990 920
rect -1020 870 -990 900
rect -1020 850 -1015 870
rect -995 850 -990 870
rect -1020 840 -990 850
rect -965 1420 -935 1430
rect -965 1400 -960 1420
rect -940 1400 -935 1420
rect -965 1370 -935 1400
rect -965 1350 -960 1370
rect -940 1350 -935 1370
rect -965 1320 -935 1350
rect -965 1300 -960 1320
rect -940 1300 -935 1320
rect -965 1270 -935 1300
rect -965 1250 -960 1270
rect -940 1250 -935 1270
rect -965 1220 -935 1250
rect -965 1200 -960 1220
rect -940 1200 -935 1220
rect -965 1170 -935 1200
rect -965 1150 -960 1170
rect -940 1150 -935 1170
rect -965 1120 -935 1150
rect -965 1100 -960 1120
rect -940 1100 -935 1120
rect -965 1070 -935 1100
rect -965 1050 -960 1070
rect -940 1050 -935 1070
rect -965 1020 -935 1050
rect -965 1000 -960 1020
rect -940 1000 -935 1020
rect -965 970 -935 1000
rect -965 950 -960 970
rect -940 950 -935 970
rect -965 920 -935 950
rect -965 900 -960 920
rect -940 900 -935 920
rect -965 870 -935 900
rect -965 850 -960 870
rect -940 850 -935 870
rect -965 840 -935 850
rect -910 1420 -880 1430
rect -910 1400 -905 1420
rect -885 1400 -880 1420
rect -910 1370 -880 1400
rect -910 1350 -905 1370
rect -885 1350 -880 1370
rect -910 1320 -880 1350
rect -910 1300 -905 1320
rect -885 1300 -880 1320
rect -910 1270 -880 1300
rect -910 1250 -905 1270
rect -885 1250 -880 1270
rect -910 1220 -880 1250
rect -910 1200 -905 1220
rect -885 1200 -880 1220
rect -910 1170 -880 1200
rect -910 1150 -905 1170
rect -885 1150 -880 1170
rect -910 1120 -880 1150
rect -910 1100 -905 1120
rect -885 1100 -880 1120
rect -910 1070 -880 1100
rect -910 1050 -905 1070
rect -885 1050 -880 1070
rect -910 1020 -880 1050
rect -910 1000 -905 1020
rect -885 1000 -880 1020
rect -910 970 -880 1000
rect -910 950 -905 970
rect -885 950 -880 970
rect -910 920 -880 950
rect -910 900 -905 920
rect -885 900 -880 920
rect -910 870 -880 900
rect -910 850 -905 870
rect -885 850 -880 870
rect -910 840 -880 850
rect -855 1420 -825 1430
rect -855 1400 -850 1420
rect -830 1400 -825 1420
rect -855 1370 -825 1400
rect -855 1350 -850 1370
rect -830 1350 -825 1370
rect -855 1320 -825 1350
rect -855 1300 -850 1320
rect -830 1300 -825 1320
rect -855 1270 -825 1300
rect -855 1250 -850 1270
rect -830 1250 -825 1270
rect -855 1220 -825 1250
rect -855 1200 -850 1220
rect -830 1200 -825 1220
rect -855 1170 -825 1200
rect -855 1150 -850 1170
rect -830 1150 -825 1170
rect -855 1120 -825 1150
rect -855 1100 -850 1120
rect -830 1100 -825 1120
rect -855 1070 -825 1100
rect -855 1050 -850 1070
rect -830 1050 -825 1070
rect -855 1020 -825 1050
rect -855 1000 -850 1020
rect -830 1000 -825 1020
rect -855 970 -825 1000
rect -855 950 -850 970
rect -830 950 -825 970
rect -855 920 -825 950
rect -855 900 -850 920
rect -830 900 -825 920
rect -855 870 -825 900
rect -855 850 -850 870
rect -830 850 -825 870
rect -855 840 -825 850
rect -800 1420 -770 1430
rect -800 1400 -795 1420
rect -775 1400 -770 1420
rect -800 1370 -770 1400
rect -800 1350 -795 1370
rect -775 1350 -770 1370
rect -800 1320 -770 1350
rect -800 1300 -795 1320
rect -775 1300 -770 1320
rect -800 1270 -770 1300
rect -800 1250 -795 1270
rect -775 1250 -770 1270
rect -800 1220 -770 1250
rect -800 1200 -795 1220
rect -775 1200 -770 1220
rect -800 1170 -770 1200
rect -800 1150 -795 1170
rect -775 1150 -770 1170
rect -800 1120 -770 1150
rect -800 1100 -795 1120
rect -775 1100 -770 1120
rect -800 1070 -770 1100
rect -800 1050 -795 1070
rect -775 1050 -770 1070
rect -800 1020 -770 1050
rect -800 1000 -795 1020
rect -775 1000 -770 1020
rect -800 970 -770 1000
rect -800 950 -795 970
rect -775 950 -770 970
rect -800 920 -770 950
rect -800 900 -795 920
rect -775 900 -770 920
rect -800 870 -770 900
rect -800 850 -795 870
rect -775 850 -770 870
rect -800 840 -770 850
rect -745 1420 -715 1430
rect -745 1400 -740 1420
rect -720 1400 -715 1420
rect -745 1370 -715 1400
rect -745 1350 -740 1370
rect -720 1350 -715 1370
rect -745 1320 -715 1350
rect -745 1300 -740 1320
rect -720 1300 -715 1320
rect -745 1270 -715 1300
rect -745 1250 -740 1270
rect -720 1250 -715 1270
rect -745 1220 -715 1250
rect -745 1200 -740 1220
rect -720 1200 -715 1220
rect -745 1170 -715 1200
rect -745 1150 -740 1170
rect -720 1150 -715 1170
rect -745 1120 -715 1150
rect -745 1100 -740 1120
rect -720 1100 -715 1120
rect -745 1070 -715 1100
rect -745 1050 -740 1070
rect -720 1050 -715 1070
rect -745 1020 -715 1050
rect -745 1000 -740 1020
rect -720 1000 -715 1020
rect -745 970 -715 1000
rect -745 950 -740 970
rect -720 950 -715 970
rect -745 920 -715 950
rect -745 900 -740 920
rect -720 900 -715 920
rect -745 870 -715 900
rect -745 850 -740 870
rect -720 850 -715 870
rect -745 840 -715 850
rect -690 1420 -660 1430
rect -690 1400 -685 1420
rect -665 1400 -660 1420
rect -690 1370 -660 1400
rect -690 1350 -685 1370
rect -665 1350 -660 1370
rect -690 1320 -660 1350
rect -690 1300 -685 1320
rect -665 1300 -660 1320
rect -690 1270 -660 1300
rect -690 1250 -685 1270
rect -665 1250 -660 1270
rect -690 1220 -660 1250
rect -690 1200 -685 1220
rect -665 1200 -660 1220
rect -690 1170 -660 1200
rect -690 1150 -685 1170
rect -665 1150 -660 1170
rect -690 1120 -660 1150
rect -690 1100 -685 1120
rect -665 1100 -660 1120
rect -690 1070 -660 1100
rect -690 1050 -685 1070
rect -665 1050 -660 1070
rect -690 1020 -660 1050
rect -690 1000 -685 1020
rect -665 1000 -660 1020
rect -690 970 -660 1000
rect -690 950 -685 970
rect -665 950 -660 970
rect -690 920 -660 950
rect -690 900 -685 920
rect -665 900 -660 920
rect -690 870 -660 900
rect -690 850 -685 870
rect -665 850 -660 870
rect -690 840 -660 850
rect -635 1420 -605 1430
rect -635 1400 -630 1420
rect -610 1400 -605 1420
rect -635 1370 -605 1400
rect -635 1350 -630 1370
rect -610 1350 -605 1370
rect -635 1320 -605 1350
rect -635 1300 -630 1320
rect -610 1300 -605 1320
rect -635 1270 -605 1300
rect -635 1250 -630 1270
rect -610 1250 -605 1270
rect -635 1220 -605 1250
rect -635 1200 -630 1220
rect -610 1200 -605 1220
rect -635 1170 -605 1200
rect -635 1150 -630 1170
rect -610 1150 -605 1170
rect -635 1120 -605 1150
rect -635 1100 -630 1120
rect -610 1100 -605 1120
rect -635 1070 -605 1100
rect -635 1050 -630 1070
rect -610 1050 -605 1070
rect -635 1020 -605 1050
rect -635 1000 -630 1020
rect -610 1000 -605 1020
rect -635 970 -605 1000
rect -635 950 -630 970
rect -610 950 -605 970
rect -635 920 -605 950
rect -635 900 -630 920
rect -610 900 -605 920
rect -635 870 -605 900
rect -635 850 -630 870
rect -610 850 -605 870
rect -635 840 -605 850
rect -580 1420 -550 1430
rect -580 1400 -575 1420
rect -555 1400 -550 1420
rect -580 1370 -550 1400
rect -580 1350 -575 1370
rect -555 1350 -550 1370
rect -580 1320 -550 1350
rect -580 1300 -575 1320
rect -555 1300 -550 1320
rect -580 1270 -550 1300
rect -580 1250 -575 1270
rect -555 1250 -550 1270
rect -580 1220 -550 1250
rect -580 1200 -575 1220
rect -555 1200 -550 1220
rect -580 1170 -550 1200
rect -580 1150 -575 1170
rect -555 1150 -550 1170
rect -580 1120 -550 1150
rect -580 1100 -575 1120
rect -555 1100 -550 1120
rect -580 1070 -550 1100
rect -580 1050 -575 1070
rect -555 1050 -550 1070
rect -580 1020 -550 1050
rect -580 1000 -575 1020
rect -555 1000 -550 1020
rect -580 970 -550 1000
rect -580 950 -575 970
rect -555 950 -550 970
rect -580 920 -550 950
rect -580 900 -575 920
rect -555 900 -550 920
rect -580 870 -550 900
rect -580 850 -575 870
rect -555 850 -550 870
rect -580 840 -550 850
rect -525 1420 -495 1430
rect -525 1400 -520 1420
rect -500 1400 -495 1420
rect -525 1370 -495 1400
rect -525 1350 -520 1370
rect -500 1350 -495 1370
rect -525 1320 -495 1350
rect -525 1300 -520 1320
rect -500 1300 -495 1320
rect -525 1270 -495 1300
rect -525 1250 -520 1270
rect -500 1250 -495 1270
rect -525 1220 -495 1250
rect -525 1200 -520 1220
rect -500 1200 -495 1220
rect -525 1170 -495 1200
rect -525 1150 -520 1170
rect -500 1150 -495 1170
rect -525 1120 -495 1150
rect -525 1100 -520 1120
rect -500 1100 -495 1120
rect -525 1070 -495 1100
rect -525 1050 -520 1070
rect -500 1050 -495 1070
rect -525 1020 -495 1050
rect -525 1000 -520 1020
rect -500 1000 -495 1020
rect -525 970 -495 1000
rect -525 950 -520 970
rect -500 950 -495 970
rect -525 920 -495 950
rect -525 900 -520 920
rect -500 900 -495 920
rect -525 870 -495 900
rect -525 850 -520 870
rect -500 850 -495 870
rect -525 840 -495 850
rect -470 1420 -400 1430
rect -470 1400 -465 1420
rect -445 1400 -425 1420
rect -405 1400 -400 1420
rect -470 1370 -400 1400
rect -470 1350 -465 1370
rect -445 1350 -425 1370
rect -405 1350 -400 1370
rect -470 1320 -400 1350
rect -470 1300 -465 1320
rect -445 1300 -425 1320
rect -405 1300 -400 1320
rect -470 1270 -400 1300
rect -470 1250 -465 1270
rect -445 1250 -425 1270
rect -405 1250 -400 1270
rect -470 1220 -400 1250
rect 420 1420 490 1450
rect 420 1400 425 1420
rect 445 1400 465 1420
rect 485 1400 490 1420
rect 420 1370 490 1400
rect 420 1350 425 1370
rect 445 1350 465 1370
rect 485 1350 490 1370
rect 420 1320 490 1350
rect 420 1300 425 1320
rect 445 1300 465 1320
rect 485 1300 490 1320
rect 420 1270 490 1300
rect 420 1250 425 1270
rect 445 1250 465 1270
rect 485 1250 490 1270
rect 420 1240 490 1250
rect 515 1470 545 1480
rect 515 1450 520 1470
rect 540 1450 545 1470
rect 515 1420 545 1450
rect 515 1400 520 1420
rect 540 1400 545 1420
rect 515 1370 545 1400
rect 515 1350 520 1370
rect 540 1350 545 1370
rect 515 1320 545 1350
rect 515 1300 520 1320
rect 540 1300 545 1320
rect 515 1270 545 1300
rect 515 1250 520 1270
rect 540 1250 545 1270
rect 515 1240 545 1250
rect 570 1470 600 1480
rect 570 1450 575 1470
rect 595 1450 600 1470
rect 570 1420 600 1450
rect 570 1400 575 1420
rect 595 1400 600 1420
rect 570 1370 600 1400
rect 570 1350 575 1370
rect 595 1350 600 1370
rect 570 1320 600 1350
rect 570 1300 575 1320
rect 595 1300 600 1320
rect 570 1270 600 1300
rect 570 1250 575 1270
rect 595 1250 600 1270
rect 570 1240 600 1250
rect 625 1470 655 1480
rect 625 1450 630 1470
rect 650 1450 655 1470
rect 625 1420 655 1450
rect 625 1400 630 1420
rect 650 1400 655 1420
rect 625 1370 655 1400
rect 625 1350 630 1370
rect 650 1350 655 1370
rect 625 1320 655 1350
rect 625 1300 630 1320
rect 650 1300 655 1320
rect 625 1270 655 1300
rect 625 1250 630 1270
rect 650 1250 655 1270
rect 625 1240 655 1250
rect 680 1470 710 1480
rect 680 1450 685 1470
rect 705 1450 710 1470
rect 680 1420 710 1450
rect 680 1400 685 1420
rect 705 1400 710 1420
rect 680 1370 710 1400
rect 680 1350 685 1370
rect 705 1350 710 1370
rect 680 1320 710 1350
rect 680 1300 685 1320
rect 705 1300 710 1320
rect 680 1270 710 1300
rect 680 1250 685 1270
rect 705 1250 710 1270
rect 680 1240 710 1250
rect 735 1470 765 1480
rect 735 1450 740 1470
rect 760 1450 765 1470
rect 735 1420 765 1450
rect 735 1400 740 1420
rect 760 1400 765 1420
rect 735 1370 765 1400
rect 735 1350 740 1370
rect 760 1350 765 1370
rect 735 1320 765 1350
rect 735 1300 740 1320
rect 760 1300 765 1320
rect 735 1270 765 1300
rect 735 1250 740 1270
rect 760 1250 765 1270
rect 735 1240 765 1250
rect 790 1470 900 1480
rect 790 1450 795 1470
rect 815 1450 835 1470
rect 855 1450 875 1470
rect 895 1450 900 1470
rect 790 1420 900 1450
rect 790 1400 795 1420
rect 815 1400 835 1420
rect 855 1400 875 1420
rect 895 1400 900 1420
rect 790 1370 900 1400
rect 790 1350 795 1370
rect 815 1350 835 1370
rect 855 1350 875 1370
rect 895 1350 900 1370
rect 790 1320 900 1350
rect 790 1300 795 1320
rect 815 1300 835 1320
rect 855 1300 875 1320
rect 895 1300 900 1320
rect 790 1270 900 1300
rect 790 1250 795 1270
rect 815 1250 835 1270
rect 855 1250 875 1270
rect 895 1250 900 1270
rect 790 1240 900 1250
rect 925 1470 955 1480
rect 925 1450 930 1470
rect 950 1450 955 1470
rect 925 1420 955 1450
rect 925 1400 930 1420
rect 950 1400 955 1420
rect 925 1370 955 1400
rect 925 1350 930 1370
rect 950 1350 955 1370
rect 925 1320 955 1350
rect 925 1300 930 1320
rect 950 1300 955 1320
rect 925 1270 955 1300
rect 925 1250 930 1270
rect 950 1250 955 1270
rect 925 1240 955 1250
rect 980 1470 1010 1480
rect 980 1450 985 1470
rect 1005 1450 1010 1470
rect 980 1420 1010 1450
rect 980 1400 985 1420
rect 1005 1400 1010 1420
rect 980 1370 1010 1400
rect 980 1350 985 1370
rect 1005 1350 1010 1370
rect 980 1320 1010 1350
rect 980 1300 985 1320
rect 1005 1300 1010 1320
rect 980 1270 1010 1300
rect 980 1250 985 1270
rect 1005 1250 1010 1270
rect 980 1240 1010 1250
rect 1035 1470 1065 1480
rect 1035 1450 1040 1470
rect 1060 1450 1065 1470
rect 1035 1420 1065 1450
rect 1035 1400 1040 1420
rect 1060 1400 1065 1420
rect 1035 1370 1065 1400
rect 1035 1350 1040 1370
rect 1060 1350 1065 1370
rect 1035 1320 1065 1350
rect 1035 1300 1040 1320
rect 1060 1300 1065 1320
rect 1035 1270 1065 1300
rect 1035 1250 1040 1270
rect 1060 1250 1065 1270
rect 1035 1240 1065 1250
rect 1090 1470 1120 1480
rect 1090 1450 1095 1470
rect 1115 1450 1120 1470
rect 1090 1420 1120 1450
rect 1090 1400 1095 1420
rect 1115 1400 1120 1420
rect 1090 1370 1120 1400
rect 1090 1350 1095 1370
rect 1115 1350 1120 1370
rect 1090 1320 1120 1350
rect 1090 1300 1095 1320
rect 1115 1300 1120 1320
rect 1090 1270 1120 1300
rect 1090 1250 1095 1270
rect 1115 1250 1120 1270
rect 1090 1240 1120 1250
rect 1145 1470 1175 1480
rect 1145 1450 1150 1470
rect 1170 1450 1175 1470
rect 1145 1420 1175 1450
rect 1145 1400 1150 1420
rect 1170 1400 1175 1420
rect 1145 1370 1175 1400
rect 1145 1350 1150 1370
rect 1170 1350 1175 1370
rect 1145 1320 1175 1350
rect 1145 1300 1150 1320
rect 1170 1300 1175 1320
rect 1145 1270 1175 1300
rect 1145 1250 1150 1270
rect 1170 1250 1175 1270
rect 1145 1240 1175 1250
rect 1200 1470 1270 1480
rect 1200 1450 1205 1470
rect 1225 1450 1245 1470
rect 1265 1450 1270 1470
rect 2125 1460 2135 1480
rect 2155 1460 2165 1480
rect 2125 1450 2165 1460
rect 2235 1480 2275 1490
rect 2235 1460 2245 1480
rect 2265 1460 2275 1480
rect 2235 1450 2275 1460
rect 2345 1480 2385 1490
rect 2345 1460 2355 1480
rect 2375 1460 2385 1480
rect 2345 1450 2385 1460
rect 2455 1480 2495 1490
rect 2455 1460 2465 1480
rect 2485 1460 2495 1480
rect 2455 1450 2495 1460
rect 2565 1480 2605 1490
rect 2565 1460 2575 1480
rect 2595 1460 2605 1480
rect 2565 1450 2605 1460
rect 2675 1480 2715 1490
rect 2675 1460 2685 1480
rect 2705 1460 2715 1480
rect 2675 1450 2715 1460
rect 2785 1480 2825 1490
rect 2785 1460 2795 1480
rect 2815 1460 2825 1480
rect 2785 1450 2825 1460
rect 1200 1420 1270 1450
rect 2135 1430 2155 1450
rect 2245 1430 2265 1450
rect 2355 1430 2375 1450
rect 2465 1430 2485 1450
rect 2575 1430 2595 1450
rect 2685 1430 2705 1450
rect 2795 1430 2815 1450
rect 1200 1400 1205 1420
rect 1225 1400 1245 1420
rect 1265 1400 1270 1420
rect 1200 1370 1270 1400
rect 1200 1350 1205 1370
rect 1225 1350 1245 1370
rect 1265 1350 1270 1370
rect 1200 1320 1270 1350
rect 1200 1300 1205 1320
rect 1225 1300 1245 1320
rect 1265 1300 1270 1320
rect 1200 1270 1270 1300
rect 1200 1250 1205 1270
rect 1225 1250 1245 1270
rect 1265 1250 1270 1270
rect 1200 1240 1270 1250
rect 2090 1420 2160 1430
rect 2090 1400 2095 1420
rect 2115 1400 2135 1420
rect 2155 1400 2160 1420
rect 2090 1370 2160 1400
rect 2090 1350 2095 1370
rect 2115 1350 2135 1370
rect 2155 1350 2160 1370
rect 2090 1320 2160 1350
rect 2090 1300 2095 1320
rect 2115 1300 2135 1320
rect 2155 1300 2160 1320
rect 2090 1270 2160 1300
rect 2090 1250 2095 1270
rect 2115 1250 2135 1270
rect 2155 1250 2160 1270
rect 515 1230 535 1240
rect -470 1200 -465 1220
rect -445 1200 -425 1220
rect -405 1200 -400 1220
rect -470 1170 -400 1200
rect 505 1220 535 1230
rect 745 1230 765 1240
rect 925 1230 945 1240
rect 745 1220 775 1230
rect 505 1200 510 1220
rect 530 1200 535 1220
rect 505 1190 535 1200
rect 552 1210 582 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1210 660 1220
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 698 1210 728 1220
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 745 1200 750 1220
rect 770 1200 775 1220
rect 745 1190 775 1200
rect 915 1220 945 1230
rect 1155 1230 1175 1240
rect 1155 1220 1185 1230
rect 915 1200 920 1220
rect 940 1200 945 1220
rect 915 1190 945 1200
rect 962 1210 992 1220
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 698 1180 728 1190
rect 962 1180 992 1190
rect 1030 1210 1070 1220
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1108 1210 1138 1220
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1155 1200 1160 1220
rect 1180 1200 1185 1220
rect 1155 1190 1185 1200
rect 2090 1220 2160 1250
rect 2090 1200 2095 1220
rect 2115 1200 2135 1220
rect 2155 1200 2160 1220
rect 1108 1180 1138 1190
rect -470 1150 -465 1170
rect -445 1150 -425 1170
rect -405 1150 -400 1170
rect 2090 1170 2160 1200
rect -470 1120 -400 1150
rect 545 1150 585 1160
rect 545 1130 555 1150
rect 575 1130 585 1150
rect 545 1120 585 1130
rect 1105 1150 1145 1160
rect 1105 1130 1115 1150
rect 1135 1130 1145 1150
rect 1105 1120 1145 1130
rect 2090 1150 2095 1170
rect 2115 1150 2135 1170
rect 2155 1150 2160 1170
rect 2090 1120 2160 1150
rect -470 1100 -465 1120
rect -445 1100 -425 1120
rect -405 1100 -400 1120
rect -470 1070 -400 1100
rect -470 1050 -465 1070
rect -445 1050 -425 1070
rect -405 1050 -400 1070
rect -470 1020 -400 1050
rect -470 1000 -465 1020
rect -445 1000 -425 1020
rect -405 1000 -400 1020
rect -470 970 -400 1000
rect -470 950 -465 970
rect -445 950 -425 970
rect -405 950 -400 970
rect -470 920 -400 950
rect 2090 1100 2095 1120
rect 2115 1100 2135 1120
rect 2155 1100 2160 1120
rect 2090 1070 2160 1100
rect 2090 1050 2095 1070
rect 2115 1050 2135 1070
rect 2155 1050 2160 1070
rect 2090 1020 2160 1050
rect 2090 1000 2095 1020
rect 2115 1000 2135 1020
rect 2155 1000 2160 1020
rect 2090 970 2160 1000
rect 2090 950 2095 970
rect 2115 950 2135 970
rect 2155 950 2160 970
rect -470 900 -465 920
rect -445 900 -425 920
rect -405 900 -400 920
rect 780 920 835 930
rect -470 870 -400 900
rect -50 900 -10 910
rect -50 880 -40 900
rect -20 880 -10 900
rect -50 870 -10 880
rect 60 900 100 910
rect 60 880 70 900
rect 90 880 100 900
rect 60 870 100 880
rect 170 900 210 910
rect 170 880 180 900
rect 200 880 210 900
rect 170 870 210 880
rect 230 900 260 910
rect 230 880 235 900
rect 255 880 260 900
rect 230 870 260 880
rect 280 900 320 910
rect 280 880 290 900
rect 310 880 320 900
rect 280 870 320 880
rect 390 900 430 910
rect 390 880 400 900
rect 420 880 430 900
rect 390 870 430 880
rect 500 900 540 910
rect 500 880 510 900
rect 530 880 540 900
rect 500 870 540 880
rect 780 900 805 920
rect 825 900 835 920
rect 780 890 835 900
rect 880 920 920 930
rect 880 900 890 920
rect 910 900 920 920
rect 2090 920 2160 950
rect 880 890 920 900
rect 1150 900 1190 910
rect 780 870 800 890
rect 890 870 910 890
rect 1150 880 1160 900
rect 1180 880 1190 900
rect 1150 870 1190 880
rect 1260 900 1300 910
rect 1260 880 1270 900
rect 1290 880 1300 900
rect 1260 870 1300 880
rect 1370 900 1410 910
rect 1370 880 1380 900
rect 1400 880 1410 900
rect 1370 870 1410 880
rect 1430 900 1460 910
rect 1430 880 1435 900
rect 1455 880 1460 900
rect 1430 870 1460 880
rect 1480 900 1520 910
rect 1480 880 1490 900
rect 1510 880 1520 900
rect 1480 870 1520 880
rect 1590 900 1630 910
rect 1590 880 1600 900
rect 1620 880 1630 900
rect 1590 870 1630 880
rect 1700 900 1740 910
rect 1700 880 1710 900
rect 1730 880 1740 900
rect 1700 870 1740 880
rect 2090 900 2095 920
rect 2115 900 2135 920
rect 2155 900 2160 920
rect 2090 870 2160 900
rect -470 850 -465 870
rect -445 850 -425 870
rect -405 850 -400 870
rect -470 840 -400 850
rect -40 845 -20 870
rect 70 845 90 870
rect 180 845 200 870
rect 290 845 310 870
rect 400 845 420 870
rect 510 845 530 870
rect 680 860 750 870
rect -1501 815 -1360 825
rect -1070 815 -1050 840
rect -960 815 -940 840
rect -850 815 -830 840
rect -740 815 -720 840
rect -630 815 -610 840
rect -520 815 -500 840
rect -140 835 -70 845
rect -140 815 -135 835
rect -115 815 -95 835
rect -75 815 -70 835
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -1080 805 -1040 815
rect -1080 785 -1070 805
rect -1050 785 -1040 805
rect -1080 775 -1040 785
rect -970 805 -930 815
rect -970 785 -960 805
rect -940 785 -930 805
rect -970 775 -930 785
rect -860 805 -820 815
rect -860 785 -850 805
rect -830 785 -820 805
rect -860 775 -820 785
rect -800 800 -770 810
rect -800 780 -795 800
rect -775 780 -770 800
rect -800 770 -770 780
rect -750 805 -710 815
rect -750 785 -740 805
rect -720 785 -710 805
rect -750 775 -710 785
rect -640 805 -600 815
rect -640 785 -630 805
rect -610 785 -600 805
rect -640 775 -600 785
rect -530 805 -490 815
rect -530 785 -520 805
rect -500 785 -490 805
rect -530 775 -490 785
rect -140 785 -70 815
rect -140 765 -135 785
rect -115 765 -95 785
rect -75 765 -70 785
rect -140 735 -70 765
rect -140 715 -135 735
rect -115 715 -95 735
rect -75 715 -70 735
rect -140 705 -70 715
rect -45 835 -15 845
rect -45 815 -40 835
rect -20 815 -15 835
rect -45 785 -15 815
rect -45 765 -40 785
rect -20 765 -15 785
rect -45 735 -15 765
rect -45 715 -40 735
rect -20 715 -15 735
rect -45 705 -15 715
rect 10 835 40 845
rect 10 815 15 835
rect 35 815 40 835
rect 10 785 40 815
rect 10 765 15 785
rect 35 765 40 785
rect 10 735 40 765
rect 10 715 15 735
rect 35 715 40 735
rect 10 705 40 715
rect 65 835 95 845
rect 65 815 70 835
rect 90 815 95 835
rect 65 785 95 815
rect 65 765 70 785
rect 90 765 95 785
rect 65 735 95 765
rect 65 715 70 735
rect 90 715 95 735
rect 65 705 95 715
rect 120 835 150 845
rect 120 815 125 835
rect 145 815 150 835
rect 120 785 150 815
rect 120 765 125 785
rect 145 765 150 785
rect 120 735 150 765
rect 120 715 125 735
rect 145 715 150 735
rect 120 705 150 715
rect 175 835 205 845
rect 175 815 180 835
rect 200 815 205 835
rect 175 785 205 815
rect 175 765 180 785
rect 200 765 205 785
rect 175 735 205 765
rect 175 715 180 735
rect 200 715 205 735
rect 175 705 205 715
rect 230 835 260 845
rect 230 815 235 835
rect 255 815 260 835
rect 230 785 260 815
rect 230 765 235 785
rect 255 765 260 785
rect 230 735 260 765
rect 230 715 235 735
rect 255 715 260 735
rect 230 705 260 715
rect 285 835 315 845
rect 285 815 290 835
rect 310 815 315 835
rect 285 785 315 815
rect 285 765 290 785
rect 310 765 315 785
rect 285 735 315 765
rect 285 715 290 735
rect 310 715 315 735
rect 285 705 315 715
rect 340 835 370 845
rect 340 815 345 835
rect 365 815 370 835
rect 340 785 370 815
rect 340 765 345 785
rect 365 765 370 785
rect 340 735 370 765
rect 340 715 345 735
rect 365 715 370 735
rect 340 705 370 715
rect 395 835 425 845
rect 395 815 400 835
rect 420 815 425 835
rect 395 785 425 815
rect 395 765 400 785
rect 420 765 425 785
rect 395 735 425 765
rect 395 715 400 735
rect 420 715 425 735
rect 395 705 425 715
rect 450 835 480 845
rect 450 815 455 835
rect 475 815 480 835
rect 450 785 480 815
rect 450 765 455 785
rect 475 765 480 785
rect 450 735 480 765
rect 450 715 455 735
rect 475 715 480 735
rect 450 705 480 715
rect 505 835 535 845
rect 505 815 510 835
rect 530 815 535 835
rect 505 785 535 815
rect 505 765 510 785
rect 530 765 535 785
rect 505 735 535 765
rect 505 715 510 735
rect 530 715 535 735
rect 505 705 535 715
rect 560 835 630 845
rect 560 815 565 835
rect 585 815 605 835
rect 625 815 630 835
rect 560 785 630 815
rect 560 765 565 785
rect 585 765 605 785
rect 625 765 630 785
rect 560 735 630 765
rect 560 715 565 735
rect 585 715 605 735
rect 625 715 630 735
rect 560 705 630 715
rect 680 840 685 860
rect 705 840 725 860
rect 745 840 750 860
rect 680 810 750 840
rect 680 790 685 810
rect 705 790 725 810
rect 745 790 750 810
rect 680 760 750 790
rect 680 740 685 760
rect 705 740 725 760
rect 745 740 750 760
rect 680 710 750 740
rect -95 685 -75 705
rect 15 685 35 705
rect 125 685 145 705
rect 235 685 255 705
rect 345 685 365 705
rect 455 685 475 705
rect 565 685 585 705
rect 680 690 685 710
rect 705 690 725 710
rect 745 690 750 710
rect -100 675 -70 685
rect -1145 665 -1105 675
rect -1145 645 -1135 665
rect -1115 645 -1105 665
rect -1145 635 -1105 645
rect -1080 665 -1040 675
rect -1080 645 -1070 665
rect -1050 645 -1040 665
rect -1080 635 -1040 645
rect -970 665 -930 675
rect -970 645 -960 665
rect -940 645 -930 665
rect -970 635 -930 645
rect -860 665 -820 675
rect -860 645 -850 665
rect -830 645 -820 665
rect -860 635 -820 645
rect -750 665 -710 675
rect -750 645 -740 665
rect -720 645 -710 665
rect -750 635 -710 645
rect -640 665 -600 675
rect -640 645 -630 665
rect -610 645 -600 665
rect -640 635 -600 645
rect -530 665 -490 675
rect -530 645 -520 665
rect -500 645 -490 665
rect -530 635 -490 645
rect -465 665 -425 675
rect -465 645 -455 665
rect -435 645 -425 665
rect -100 655 -95 675
rect -75 655 -70 675
rect -100 645 -70 655
rect 5 675 45 685
rect 5 655 15 675
rect 35 655 45 675
rect 5 645 45 655
rect 115 675 155 685
rect 115 655 125 675
rect 145 655 155 675
rect 115 645 155 655
rect 225 675 265 685
rect 225 655 235 675
rect 255 655 265 675
rect 225 645 265 655
rect 335 675 375 685
rect 335 655 345 675
rect 365 655 375 675
rect 335 645 375 655
rect 445 675 485 685
rect 445 655 455 675
rect 475 655 485 675
rect 445 645 485 655
rect 560 675 590 685
rect 560 655 565 675
rect 585 655 590 675
rect 560 645 590 655
rect 680 660 750 690
rect -465 635 -425 645
rect 680 640 685 660
rect 705 640 725 660
rect 745 640 750 660
rect -1125 615 -1105 635
rect -1070 615 -1050 635
rect -960 615 -940 635
rect -850 615 -830 635
rect -740 615 -720 635
rect -630 615 -610 635
rect -520 615 -500 635
rect -465 615 -445 635
rect 680 630 750 640
rect 775 860 805 870
rect 775 840 780 860
rect 800 840 805 860
rect 775 810 805 840
rect 775 790 780 810
rect 800 790 805 810
rect 775 760 805 790
rect 775 740 780 760
rect 800 740 805 760
rect 775 710 805 740
rect 775 690 780 710
rect 800 690 805 710
rect 775 660 805 690
rect 775 640 780 660
rect 800 640 805 660
rect 775 630 805 640
rect 830 860 860 870
rect 830 840 835 860
rect 855 840 860 860
rect 830 810 860 840
rect 830 790 835 810
rect 855 790 860 810
rect 830 760 860 790
rect 830 740 835 760
rect 855 740 860 760
rect 830 710 860 740
rect 830 690 835 710
rect 855 690 860 710
rect 830 660 860 690
rect 830 640 835 660
rect 855 640 860 660
rect 830 630 860 640
rect 885 860 915 870
rect 885 840 890 860
rect 910 840 915 860
rect 885 810 915 840
rect 885 790 890 810
rect 910 790 915 810
rect 885 760 915 790
rect 885 740 890 760
rect 910 740 915 760
rect 885 710 915 740
rect 885 690 890 710
rect 910 690 915 710
rect 885 660 915 690
rect 885 640 890 660
rect 910 640 915 660
rect 885 630 915 640
rect 940 860 1010 870
rect 940 840 945 860
rect 965 840 985 860
rect 1005 840 1010 860
rect 1160 845 1180 870
rect 1270 845 1290 870
rect 1380 845 1400 870
rect 1490 845 1510 870
rect 1600 845 1620 870
rect 1710 845 1730 870
rect 2090 850 2095 870
rect 2115 850 2135 870
rect 2155 850 2160 870
rect 940 810 1010 840
rect 940 790 945 810
rect 965 790 985 810
rect 1005 790 1010 810
rect 940 760 1010 790
rect 940 740 945 760
rect 965 740 985 760
rect 1005 740 1010 760
rect 940 710 1010 740
rect 940 690 945 710
rect 965 690 985 710
rect 1005 690 1010 710
rect 1060 835 1130 845
rect 1060 815 1065 835
rect 1085 815 1105 835
rect 1125 815 1130 835
rect 1060 785 1130 815
rect 1060 765 1065 785
rect 1085 765 1105 785
rect 1125 765 1130 785
rect 1060 735 1130 765
rect 1060 715 1065 735
rect 1085 715 1105 735
rect 1125 715 1130 735
rect 1060 705 1130 715
rect 1155 835 1185 845
rect 1155 815 1160 835
rect 1180 815 1185 835
rect 1155 785 1185 815
rect 1155 765 1160 785
rect 1180 765 1185 785
rect 1155 735 1185 765
rect 1155 715 1160 735
rect 1180 715 1185 735
rect 1155 705 1185 715
rect 1210 835 1240 845
rect 1210 815 1215 835
rect 1235 815 1240 835
rect 1210 785 1240 815
rect 1210 765 1215 785
rect 1235 765 1240 785
rect 1210 735 1240 765
rect 1210 715 1215 735
rect 1235 715 1240 735
rect 1210 705 1240 715
rect 1265 835 1295 845
rect 1265 815 1270 835
rect 1290 815 1295 835
rect 1265 785 1295 815
rect 1265 765 1270 785
rect 1290 765 1295 785
rect 1265 735 1295 765
rect 1265 715 1270 735
rect 1290 715 1295 735
rect 1265 705 1295 715
rect 1320 835 1350 845
rect 1320 815 1325 835
rect 1345 815 1350 835
rect 1320 785 1350 815
rect 1320 765 1325 785
rect 1345 765 1350 785
rect 1320 735 1350 765
rect 1320 715 1325 735
rect 1345 715 1350 735
rect 1320 705 1350 715
rect 1375 835 1405 845
rect 1375 815 1380 835
rect 1400 815 1405 835
rect 1375 785 1405 815
rect 1375 765 1380 785
rect 1400 765 1405 785
rect 1375 735 1405 765
rect 1375 715 1380 735
rect 1400 715 1405 735
rect 1375 705 1405 715
rect 1430 835 1460 845
rect 1430 815 1435 835
rect 1455 815 1460 835
rect 1430 785 1460 815
rect 1430 765 1435 785
rect 1455 765 1460 785
rect 1430 735 1460 765
rect 1430 715 1435 735
rect 1455 715 1460 735
rect 1430 705 1460 715
rect 1485 835 1515 845
rect 1485 815 1490 835
rect 1510 815 1515 835
rect 1485 785 1515 815
rect 1485 765 1490 785
rect 1510 765 1515 785
rect 1485 735 1515 765
rect 1485 715 1490 735
rect 1510 715 1515 735
rect 1485 705 1515 715
rect 1540 835 1570 845
rect 1540 815 1545 835
rect 1565 815 1570 835
rect 1540 785 1570 815
rect 1540 765 1545 785
rect 1565 765 1570 785
rect 1540 735 1570 765
rect 1540 715 1545 735
rect 1565 715 1570 735
rect 1540 705 1570 715
rect 1595 835 1625 845
rect 1595 815 1600 835
rect 1620 815 1625 835
rect 1595 785 1625 815
rect 1595 765 1600 785
rect 1620 765 1625 785
rect 1595 735 1625 765
rect 1595 715 1600 735
rect 1620 715 1625 735
rect 1595 705 1625 715
rect 1650 835 1680 845
rect 1650 815 1655 835
rect 1675 815 1680 835
rect 1650 785 1680 815
rect 1650 765 1655 785
rect 1675 765 1680 785
rect 1650 735 1680 765
rect 1650 715 1655 735
rect 1675 715 1680 735
rect 1650 705 1680 715
rect 1705 835 1735 845
rect 1705 815 1710 835
rect 1730 815 1735 835
rect 1705 785 1735 815
rect 1705 765 1710 785
rect 1730 765 1735 785
rect 1705 735 1735 765
rect 1705 715 1710 735
rect 1730 715 1735 735
rect 1705 705 1735 715
rect 1760 835 1830 845
rect 2090 840 2160 850
rect 2185 1420 2215 1430
rect 2185 1400 2190 1420
rect 2210 1400 2215 1420
rect 2185 1370 2215 1400
rect 2185 1350 2190 1370
rect 2210 1350 2215 1370
rect 2185 1320 2215 1350
rect 2185 1300 2190 1320
rect 2210 1300 2215 1320
rect 2185 1270 2215 1300
rect 2185 1250 2190 1270
rect 2210 1250 2215 1270
rect 2185 1220 2215 1250
rect 2185 1200 2190 1220
rect 2210 1200 2215 1220
rect 2185 1170 2215 1200
rect 2185 1150 2190 1170
rect 2210 1150 2215 1170
rect 2185 1120 2215 1150
rect 2185 1100 2190 1120
rect 2210 1100 2215 1120
rect 2185 1070 2215 1100
rect 2185 1050 2190 1070
rect 2210 1050 2215 1070
rect 2185 1020 2215 1050
rect 2185 1000 2190 1020
rect 2210 1000 2215 1020
rect 2185 970 2215 1000
rect 2185 950 2190 970
rect 2210 950 2215 970
rect 2185 920 2215 950
rect 2185 900 2190 920
rect 2210 900 2215 920
rect 2185 870 2215 900
rect 2185 850 2190 870
rect 2210 850 2215 870
rect 2185 840 2215 850
rect 2240 1420 2270 1430
rect 2240 1400 2245 1420
rect 2265 1400 2270 1420
rect 2240 1370 2270 1400
rect 2240 1350 2245 1370
rect 2265 1350 2270 1370
rect 2240 1320 2270 1350
rect 2240 1300 2245 1320
rect 2265 1300 2270 1320
rect 2240 1270 2270 1300
rect 2240 1250 2245 1270
rect 2265 1250 2270 1270
rect 2240 1220 2270 1250
rect 2240 1200 2245 1220
rect 2265 1200 2270 1220
rect 2240 1170 2270 1200
rect 2240 1150 2245 1170
rect 2265 1150 2270 1170
rect 2240 1120 2270 1150
rect 2240 1100 2245 1120
rect 2265 1100 2270 1120
rect 2240 1070 2270 1100
rect 2240 1050 2245 1070
rect 2265 1050 2270 1070
rect 2240 1020 2270 1050
rect 2240 1000 2245 1020
rect 2265 1000 2270 1020
rect 2240 970 2270 1000
rect 2240 950 2245 970
rect 2265 950 2270 970
rect 2240 920 2270 950
rect 2240 900 2245 920
rect 2265 900 2270 920
rect 2240 870 2270 900
rect 2240 850 2245 870
rect 2265 850 2270 870
rect 2240 840 2270 850
rect 2295 1420 2325 1430
rect 2295 1400 2300 1420
rect 2320 1400 2325 1420
rect 2295 1370 2325 1400
rect 2295 1350 2300 1370
rect 2320 1350 2325 1370
rect 2295 1320 2325 1350
rect 2295 1300 2300 1320
rect 2320 1300 2325 1320
rect 2295 1270 2325 1300
rect 2295 1250 2300 1270
rect 2320 1250 2325 1270
rect 2295 1220 2325 1250
rect 2295 1200 2300 1220
rect 2320 1200 2325 1220
rect 2295 1170 2325 1200
rect 2295 1150 2300 1170
rect 2320 1150 2325 1170
rect 2295 1120 2325 1150
rect 2295 1100 2300 1120
rect 2320 1100 2325 1120
rect 2295 1070 2325 1100
rect 2295 1050 2300 1070
rect 2320 1050 2325 1070
rect 2295 1020 2325 1050
rect 2295 1000 2300 1020
rect 2320 1000 2325 1020
rect 2295 970 2325 1000
rect 2295 950 2300 970
rect 2320 950 2325 970
rect 2295 920 2325 950
rect 2295 900 2300 920
rect 2320 900 2325 920
rect 2295 870 2325 900
rect 2295 850 2300 870
rect 2320 850 2325 870
rect 2295 840 2325 850
rect 2350 1420 2380 1430
rect 2350 1400 2355 1420
rect 2375 1400 2380 1420
rect 2350 1370 2380 1400
rect 2350 1350 2355 1370
rect 2375 1350 2380 1370
rect 2350 1320 2380 1350
rect 2350 1300 2355 1320
rect 2375 1300 2380 1320
rect 2350 1270 2380 1300
rect 2350 1250 2355 1270
rect 2375 1250 2380 1270
rect 2350 1220 2380 1250
rect 2350 1200 2355 1220
rect 2375 1200 2380 1220
rect 2350 1170 2380 1200
rect 2350 1150 2355 1170
rect 2375 1150 2380 1170
rect 2350 1120 2380 1150
rect 2350 1100 2355 1120
rect 2375 1100 2380 1120
rect 2350 1070 2380 1100
rect 2350 1050 2355 1070
rect 2375 1050 2380 1070
rect 2350 1020 2380 1050
rect 2350 1000 2355 1020
rect 2375 1000 2380 1020
rect 2350 970 2380 1000
rect 2350 950 2355 970
rect 2375 950 2380 970
rect 2350 920 2380 950
rect 2350 900 2355 920
rect 2375 900 2380 920
rect 2350 870 2380 900
rect 2350 850 2355 870
rect 2375 850 2380 870
rect 2350 840 2380 850
rect 2405 1420 2435 1430
rect 2405 1400 2410 1420
rect 2430 1400 2435 1420
rect 2405 1370 2435 1400
rect 2405 1350 2410 1370
rect 2430 1350 2435 1370
rect 2405 1320 2435 1350
rect 2405 1300 2410 1320
rect 2430 1300 2435 1320
rect 2405 1270 2435 1300
rect 2405 1250 2410 1270
rect 2430 1250 2435 1270
rect 2405 1220 2435 1250
rect 2405 1200 2410 1220
rect 2430 1200 2435 1220
rect 2405 1170 2435 1200
rect 2405 1150 2410 1170
rect 2430 1150 2435 1170
rect 2405 1120 2435 1150
rect 2405 1100 2410 1120
rect 2430 1100 2435 1120
rect 2405 1070 2435 1100
rect 2405 1050 2410 1070
rect 2430 1050 2435 1070
rect 2405 1020 2435 1050
rect 2405 1000 2410 1020
rect 2430 1000 2435 1020
rect 2405 970 2435 1000
rect 2405 950 2410 970
rect 2430 950 2435 970
rect 2405 920 2435 950
rect 2405 900 2410 920
rect 2430 900 2435 920
rect 2405 870 2435 900
rect 2405 850 2410 870
rect 2430 850 2435 870
rect 2405 840 2435 850
rect 2460 1420 2490 1430
rect 2460 1400 2465 1420
rect 2485 1400 2490 1420
rect 2460 1370 2490 1400
rect 2460 1350 2465 1370
rect 2485 1350 2490 1370
rect 2460 1320 2490 1350
rect 2460 1300 2465 1320
rect 2485 1300 2490 1320
rect 2460 1270 2490 1300
rect 2460 1250 2465 1270
rect 2485 1250 2490 1270
rect 2460 1220 2490 1250
rect 2460 1200 2465 1220
rect 2485 1200 2490 1220
rect 2460 1170 2490 1200
rect 2460 1150 2465 1170
rect 2485 1150 2490 1170
rect 2460 1120 2490 1150
rect 2460 1100 2465 1120
rect 2485 1100 2490 1120
rect 2460 1070 2490 1100
rect 2460 1050 2465 1070
rect 2485 1050 2490 1070
rect 2460 1020 2490 1050
rect 2460 1000 2465 1020
rect 2485 1000 2490 1020
rect 2460 970 2490 1000
rect 2460 950 2465 970
rect 2485 950 2490 970
rect 2460 920 2490 950
rect 2460 900 2465 920
rect 2485 900 2490 920
rect 2460 870 2490 900
rect 2460 850 2465 870
rect 2485 850 2490 870
rect 2460 840 2490 850
rect 2515 1420 2545 1430
rect 2515 1400 2520 1420
rect 2540 1400 2545 1420
rect 2515 1370 2545 1400
rect 2515 1350 2520 1370
rect 2540 1350 2545 1370
rect 2515 1320 2545 1350
rect 2515 1300 2520 1320
rect 2540 1300 2545 1320
rect 2515 1270 2545 1300
rect 2515 1250 2520 1270
rect 2540 1250 2545 1270
rect 2515 1220 2545 1250
rect 2515 1200 2520 1220
rect 2540 1200 2545 1220
rect 2515 1170 2545 1200
rect 2515 1150 2520 1170
rect 2540 1150 2545 1170
rect 2515 1120 2545 1150
rect 2515 1100 2520 1120
rect 2540 1100 2545 1120
rect 2515 1070 2545 1100
rect 2515 1050 2520 1070
rect 2540 1050 2545 1070
rect 2515 1020 2545 1050
rect 2515 1000 2520 1020
rect 2540 1000 2545 1020
rect 2515 970 2545 1000
rect 2515 950 2520 970
rect 2540 950 2545 970
rect 2515 920 2545 950
rect 2515 900 2520 920
rect 2540 900 2545 920
rect 2515 870 2545 900
rect 2515 850 2520 870
rect 2540 850 2545 870
rect 2515 840 2545 850
rect 2570 1420 2600 1430
rect 2570 1400 2575 1420
rect 2595 1400 2600 1420
rect 2570 1370 2600 1400
rect 2570 1350 2575 1370
rect 2595 1350 2600 1370
rect 2570 1320 2600 1350
rect 2570 1300 2575 1320
rect 2595 1300 2600 1320
rect 2570 1270 2600 1300
rect 2570 1250 2575 1270
rect 2595 1250 2600 1270
rect 2570 1220 2600 1250
rect 2570 1200 2575 1220
rect 2595 1200 2600 1220
rect 2570 1170 2600 1200
rect 2570 1150 2575 1170
rect 2595 1150 2600 1170
rect 2570 1120 2600 1150
rect 2570 1100 2575 1120
rect 2595 1100 2600 1120
rect 2570 1070 2600 1100
rect 2570 1050 2575 1070
rect 2595 1050 2600 1070
rect 2570 1020 2600 1050
rect 2570 1000 2575 1020
rect 2595 1000 2600 1020
rect 2570 970 2600 1000
rect 2570 950 2575 970
rect 2595 950 2600 970
rect 2570 920 2600 950
rect 2570 900 2575 920
rect 2595 900 2600 920
rect 2570 870 2600 900
rect 2570 850 2575 870
rect 2595 850 2600 870
rect 2570 840 2600 850
rect 2625 1420 2655 1430
rect 2625 1400 2630 1420
rect 2650 1400 2655 1420
rect 2625 1370 2655 1400
rect 2625 1350 2630 1370
rect 2650 1350 2655 1370
rect 2625 1320 2655 1350
rect 2625 1300 2630 1320
rect 2650 1300 2655 1320
rect 2625 1270 2655 1300
rect 2625 1250 2630 1270
rect 2650 1250 2655 1270
rect 2625 1220 2655 1250
rect 2625 1200 2630 1220
rect 2650 1200 2655 1220
rect 2625 1170 2655 1200
rect 2625 1150 2630 1170
rect 2650 1150 2655 1170
rect 2625 1120 2655 1150
rect 2625 1100 2630 1120
rect 2650 1100 2655 1120
rect 2625 1070 2655 1100
rect 2625 1050 2630 1070
rect 2650 1050 2655 1070
rect 2625 1020 2655 1050
rect 2625 1000 2630 1020
rect 2650 1000 2655 1020
rect 2625 970 2655 1000
rect 2625 950 2630 970
rect 2650 950 2655 970
rect 2625 920 2655 950
rect 2625 900 2630 920
rect 2650 900 2655 920
rect 2625 870 2655 900
rect 2625 850 2630 870
rect 2650 850 2655 870
rect 2625 840 2655 850
rect 2680 1420 2710 1430
rect 2680 1400 2685 1420
rect 2705 1400 2710 1420
rect 2680 1370 2710 1400
rect 2680 1350 2685 1370
rect 2705 1350 2710 1370
rect 2680 1320 2710 1350
rect 2680 1300 2685 1320
rect 2705 1300 2710 1320
rect 2680 1270 2710 1300
rect 2680 1250 2685 1270
rect 2705 1250 2710 1270
rect 2680 1220 2710 1250
rect 2680 1200 2685 1220
rect 2705 1200 2710 1220
rect 2680 1170 2710 1200
rect 2680 1150 2685 1170
rect 2705 1150 2710 1170
rect 2680 1120 2710 1150
rect 2680 1100 2685 1120
rect 2705 1100 2710 1120
rect 2680 1070 2710 1100
rect 2680 1050 2685 1070
rect 2705 1050 2710 1070
rect 2680 1020 2710 1050
rect 2680 1000 2685 1020
rect 2705 1000 2710 1020
rect 2680 970 2710 1000
rect 2680 950 2685 970
rect 2705 950 2710 970
rect 2680 920 2710 950
rect 2680 900 2685 920
rect 2705 900 2710 920
rect 2680 870 2710 900
rect 2680 850 2685 870
rect 2705 850 2710 870
rect 2680 840 2710 850
rect 2735 1420 2765 1430
rect 2735 1400 2740 1420
rect 2760 1400 2765 1420
rect 2735 1370 2765 1400
rect 2735 1350 2740 1370
rect 2760 1350 2765 1370
rect 2735 1320 2765 1350
rect 2735 1300 2740 1320
rect 2760 1300 2765 1320
rect 2735 1270 2765 1300
rect 2735 1250 2740 1270
rect 2760 1250 2765 1270
rect 2735 1220 2765 1250
rect 2735 1200 2740 1220
rect 2760 1200 2765 1220
rect 2735 1170 2765 1200
rect 2735 1150 2740 1170
rect 2760 1150 2765 1170
rect 2735 1120 2765 1150
rect 2735 1100 2740 1120
rect 2760 1100 2765 1120
rect 2735 1070 2765 1100
rect 2735 1050 2740 1070
rect 2760 1050 2765 1070
rect 2735 1020 2765 1050
rect 2735 1000 2740 1020
rect 2760 1000 2765 1020
rect 2735 970 2765 1000
rect 2735 950 2740 970
rect 2760 950 2765 970
rect 2735 920 2765 950
rect 2735 900 2740 920
rect 2760 900 2765 920
rect 2735 870 2765 900
rect 2735 850 2740 870
rect 2760 850 2765 870
rect 2735 840 2765 850
rect 2790 1420 2860 1430
rect 2790 1400 2795 1420
rect 2815 1400 2835 1420
rect 2855 1400 2860 1420
rect 2790 1370 2860 1400
rect 2790 1350 2795 1370
rect 2815 1350 2835 1370
rect 2855 1350 2860 1370
rect 2790 1320 2860 1350
rect 2790 1300 2795 1320
rect 2815 1300 2835 1320
rect 2855 1300 2860 1320
rect 2790 1270 2860 1300
rect 2790 1250 2795 1270
rect 2815 1250 2835 1270
rect 2855 1250 2860 1270
rect 2790 1220 2860 1250
rect 2790 1200 2795 1220
rect 2815 1200 2835 1220
rect 2855 1200 2860 1220
rect 2790 1170 2860 1200
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2790 1150 2795 1170
rect 2815 1150 2835 1170
rect 2855 1150 2860 1170
rect 2790 1120 2860 1150
rect 2790 1100 2795 1120
rect 2815 1100 2835 1120
rect 2855 1100 2860 1120
rect 2790 1070 2860 1100
rect 2790 1050 2795 1070
rect 2815 1050 2835 1070
rect 2855 1050 2860 1070
rect 2790 1020 2860 1050
rect 2790 1000 2795 1020
rect 2815 1000 2835 1020
rect 2855 1000 2860 1020
rect 2790 970 2860 1000
rect 2790 950 2795 970
rect 2815 950 2835 970
rect 2855 950 2860 970
rect 2790 920 2860 950
rect 2790 900 2795 920
rect 2815 900 2835 920
rect 2855 900 2860 920
rect 2790 870 2860 900
rect 2790 850 2795 870
rect 2815 850 2835 870
rect 2855 850 2860 870
rect 2790 840 2860 850
rect 1760 815 1765 835
rect 1785 815 1805 835
rect 1825 815 1830 835
rect 2190 815 2210 840
rect 2300 815 2320 840
rect 2410 815 2430 840
rect 2520 815 2540 840
rect 2630 815 2650 840
rect 2740 815 2760 840
rect 3050 815 3191 825
rect 1760 785 1830 815
rect 1760 765 1765 785
rect 1785 765 1805 785
rect 1825 765 1830 785
rect 2180 805 2220 815
rect 2180 785 2190 805
rect 2210 785 2220 805
rect 2180 775 2220 785
rect 2290 805 2330 815
rect 2290 785 2300 805
rect 2320 785 2330 805
rect 2290 775 2330 785
rect 2400 805 2440 815
rect 2400 785 2410 805
rect 2430 785 2440 805
rect 2400 775 2440 785
rect 2460 800 2490 810
rect 2460 780 2465 800
rect 2485 780 2490 800
rect 2460 770 2490 780
rect 2510 805 2550 815
rect 2510 785 2520 805
rect 2540 785 2550 805
rect 2510 775 2550 785
rect 2620 805 2660 815
rect 2620 785 2630 805
rect 2650 785 2660 805
rect 2620 775 2660 785
rect 2730 805 2770 815
rect 2730 785 2740 805
rect 2760 785 2770 805
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2730 775 2770 785
rect 1760 735 1830 765
rect 1760 715 1765 735
rect 1785 715 1805 735
rect 1825 715 1830 735
rect 1760 705 1830 715
rect 940 660 1010 690
rect 1105 685 1125 705
rect 1215 685 1235 705
rect 1325 685 1345 705
rect 1435 685 1455 705
rect 1545 685 1565 705
rect 1655 685 1675 705
rect 1765 685 1785 705
rect 940 640 945 660
rect 965 640 985 660
rect 1005 640 1010 660
rect 1100 675 1130 685
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1100 645 1130 655
rect 1205 675 1245 685
rect 1205 655 1215 675
rect 1235 655 1245 675
rect 1205 645 1245 655
rect 1315 675 1355 685
rect 1315 655 1325 675
rect 1345 655 1355 675
rect 1315 645 1355 655
rect 1425 675 1465 685
rect 1425 655 1435 675
rect 1455 655 1465 675
rect 1425 645 1465 655
rect 1535 675 1575 685
rect 1535 655 1545 675
rect 1565 655 1575 675
rect 1535 645 1575 655
rect 1645 675 1685 685
rect 1645 655 1655 675
rect 1675 655 1685 675
rect 1645 645 1685 655
rect 1760 675 1790 685
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2115 665 2155 675
rect 2115 645 2125 665
rect 2145 645 2155 665
rect 940 630 1010 640
rect 2115 635 2155 645
rect 2180 665 2220 675
rect 2180 645 2190 665
rect 2210 645 2220 665
rect 2180 635 2220 645
rect 2290 665 2330 675
rect 2290 645 2300 665
rect 2320 645 2330 665
rect 2290 635 2330 645
rect 2400 665 2440 675
rect 2400 645 2410 665
rect 2430 645 2440 665
rect 2400 635 2440 645
rect 2510 665 2550 675
rect 2510 645 2520 665
rect 2540 645 2550 665
rect 2510 635 2550 645
rect 2620 665 2660 675
rect 2620 645 2630 665
rect 2650 645 2660 665
rect 2620 635 2660 645
rect 2730 665 2770 675
rect 2730 645 2740 665
rect 2760 645 2770 665
rect 2730 635 2770 645
rect 2795 665 2835 675
rect 2795 645 2805 665
rect 2825 645 2835 665
rect 2795 635 2835 645
rect -1170 605 -1100 615
rect -1170 585 -1165 605
rect -1145 585 -1125 605
rect -1105 585 -1100 605
rect -1490 537 -1275 572
rect -1490 517 -1455 537
rect -1310 517 -1275 537
rect -1395 467 -1370 517
rect -1170 555 -1100 585
rect -1170 535 -1165 555
rect -1145 535 -1125 555
rect -1105 535 -1100 555
rect -1170 505 -1100 535
rect -1170 485 -1165 505
rect -1145 485 -1125 505
rect -1105 485 -1100 505
rect -1170 455 -1100 485
rect -1170 435 -1165 455
rect -1145 435 -1125 455
rect -1105 435 -1100 455
rect -1170 425 -1100 435
rect -1075 605 -1045 615
rect -1075 585 -1070 605
rect -1050 585 -1045 605
rect -1075 555 -1045 585
rect -1075 535 -1070 555
rect -1050 535 -1045 555
rect -1075 505 -1045 535
rect -1075 485 -1070 505
rect -1050 485 -1045 505
rect -1075 455 -1045 485
rect -1075 435 -1070 455
rect -1050 435 -1045 455
rect -1075 425 -1045 435
rect -1020 605 -990 615
rect -1020 585 -1015 605
rect -995 585 -990 605
rect -1020 555 -990 585
rect -1020 535 -1015 555
rect -995 535 -990 555
rect -1020 505 -990 535
rect -1020 485 -1015 505
rect -995 485 -990 505
rect -1020 455 -990 485
rect -1020 435 -1015 455
rect -995 435 -990 455
rect -1020 425 -990 435
rect -965 605 -935 615
rect -965 585 -960 605
rect -940 585 -935 605
rect -965 555 -935 585
rect -965 535 -960 555
rect -940 535 -935 555
rect -965 505 -935 535
rect -965 485 -960 505
rect -940 485 -935 505
rect -965 455 -935 485
rect -965 435 -960 455
rect -940 435 -935 455
rect -965 425 -935 435
rect -910 605 -880 615
rect -910 585 -905 605
rect -885 585 -880 605
rect -910 555 -880 585
rect -910 535 -905 555
rect -885 535 -880 555
rect -910 505 -880 535
rect -910 485 -905 505
rect -885 485 -880 505
rect -910 455 -880 485
rect -910 435 -905 455
rect -885 435 -880 455
rect -910 425 -880 435
rect -855 605 -825 615
rect -855 585 -850 605
rect -830 585 -825 605
rect -855 555 -825 585
rect -855 535 -850 555
rect -830 535 -825 555
rect -855 505 -825 535
rect -855 485 -850 505
rect -830 485 -825 505
rect -855 455 -825 485
rect -855 435 -850 455
rect -830 435 -825 455
rect -855 425 -825 435
rect -800 605 -770 615
rect -800 585 -795 605
rect -775 585 -770 605
rect -800 555 -770 585
rect -800 535 -795 555
rect -775 535 -770 555
rect -800 505 -770 535
rect -800 485 -795 505
rect -775 485 -770 505
rect -800 455 -770 485
rect -800 435 -795 455
rect -775 435 -770 455
rect -800 425 -770 435
rect -745 605 -715 615
rect -745 585 -740 605
rect -720 585 -715 605
rect -745 555 -715 585
rect -745 535 -740 555
rect -720 535 -715 555
rect -745 505 -715 535
rect -745 485 -740 505
rect -720 485 -715 505
rect -745 455 -715 485
rect -745 435 -740 455
rect -720 435 -715 455
rect -745 425 -715 435
rect -690 605 -660 615
rect -690 585 -685 605
rect -665 585 -660 605
rect -690 555 -660 585
rect -690 535 -685 555
rect -665 535 -660 555
rect -690 505 -660 535
rect -690 485 -685 505
rect -665 485 -660 505
rect -690 455 -660 485
rect -690 435 -685 455
rect -665 435 -660 455
rect -690 425 -660 435
rect -635 605 -605 615
rect -635 585 -630 605
rect -610 585 -605 605
rect -635 555 -605 585
rect -635 535 -630 555
rect -610 535 -605 555
rect -635 505 -605 535
rect -635 485 -630 505
rect -610 485 -605 505
rect -635 455 -605 485
rect -635 435 -630 455
rect -610 435 -605 455
rect -635 425 -605 435
rect -580 605 -550 615
rect -580 585 -575 605
rect -555 585 -550 605
rect -580 555 -550 585
rect -580 535 -575 555
rect -555 535 -550 555
rect -580 505 -550 535
rect -580 485 -575 505
rect -555 485 -550 505
rect -580 455 -550 485
rect -580 435 -575 455
rect -555 435 -550 455
rect -580 425 -550 435
rect -525 605 -495 615
rect -525 585 -520 605
rect -500 585 -495 605
rect -525 555 -495 585
rect -525 535 -520 555
rect -500 535 -495 555
rect -525 505 -495 535
rect -525 485 -520 505
rect -500 485 -495 505
rect -525 455 -495 485
rect -525 435 -520 455
rect -500 435 -495 455
rect -525 425 -495 435
rect -470 605 -400 615
rect 725 610 745 630
rect 835 610 855 630
rect 945 610 965 630
rect 2135 615 2155 635
rect 2190 615 2210 635
rect 2300 615 2320 635
rect 2410 615 2430 635
rect 2520 615 2540 635
rect 2630 615 2650 635
rect 2740 615 2760 635
rect 2795 615 2815 635
rect -470 585 -465 605
rect -445 585 -425 605
rect -405 585 -400 605
rect -470 555 -400 585
rect 715 600 755 610
rect 715 580 725 600
rect 745 580 755 600
rect 715 570 755 580
rect 825 600 865 610
rect 825 580 835 600
rect 855 580 865 600
rect 825 570 865 580
rect 935 600 975 610
rect 935 580 945 600
rect 965 580 975 600
rect 935 570 975 580
rect 2090 605 2160 615
rect 2090 585 2095 605
rect 2115 585 2135 605
rect 2155 585 2160 605
rect -470 535 -465 555
rect -445 535 -425 555
rect -405 535 -400 555
rect -470 505 -400 535
rect -50 550 -10 560
rect -50 530 -40 550
rect -20 530 -10 550
rect -50 520 -10 530
rect 60 550 100 560
rect 60 530 70 550
rect 90 530 100 550
rect 60 520 100 530
rect 170 550 210 560
rect 170 530 180 550
rect 200 530 210 550
rect 230 530 260 570
rect 280 550 320 560
rect 280 530 290 550
rect 310 530 320 550
rect 170 520 210 530
rect 280 520 320 530
rect 390 550 430 560
rect 390 530 400 550
rect 420 530 430 550
rect 390 520 430 530
rect 500 550 540 560
rect 500 530 510 550
rect 530 530 540 550
rect 500 520 540 530
rect 1150 550 1190 560
rect 1150 530 1160 550
rect 1180 530 1190 550
rect 1150 520 1190 530
rect 1260 550 1300 560
rect 1260 530 1270 550
rect 1290 530 1300 550
rect 1260 520 1300 530
rect 1370 550 1410 560
rect 1370 530 1380 550
rect 1400 530 1410 550
rect 1430 530 1460 570
rect 1480 550 1520 560
rect 1480 530 1490 550
rect 1510 530 1520 550
rect 1370 520 1410 530
rect 1480 520 1520 530
rect 1590 550 1630 560
rect 1590 530 1600 550
rect 1620 530 1630 550
rect 1590 520 1630 530
rect 1700 550 1740 560
rect 1700 530 1710 550
rect 1730 530 1740 550
rect 1700 520 1740 530
rect 2090 555 2160 585
rect 2090 535 2095 555
rect 2115 535 2135 555
rect 2155 535 2160 555
rect -470 485 -465 505
rect -445 485 -425 505
rect -405 485 -400 505
rect -470 455 -400 485
rect -470 435 -465 455
rect -445 435 -425 455
rect -405 435 -400 455
rect -40 450 -20 520
rect 70 450 90 520
rect 180 450 200 520
rect 230 500 260 510
rect 230 480 235 500
rect 255 480 260 500
rect 230 470 260 480
rect 290 450 310 520
rect 400 450 420 520
rect 510 450 530 520
rect 715 500 755 510
rect 715 480 725 500
rect 745 480 755 500
rect 715 470 755 480
rect 795 500 825 510
rect 795 480 800 500
rect 820 480 825 500
rect 795 470 825 480
rect 865 500 895 510
rect 865 480 870 500
rect 890 480 895 500
rect 865 470 895 480
rect 935 500 975 510
rect 935 480 945 500
rect 965 480 975 500
rect 935 470 975 480
rect 725 450 745 470
rect 945 450 965 470
rect 1160 450 1180 520
rect 1270 450 1290 520
rect 1380 450 1400 520
rect 1430 500 1460 510
rect 1430 480 1435 500
rect 1455 480 1460 500
rect 1430 470 1460 480
rect 1490 450 1510 520
rect 1600 450 1620 520
rect 1710 450 1730 520
rect 2090 505 2160 535
rect 2090 485 2095 505
rect 2115 485 2135 505
rect 2155 485 2160 505
rect 2090 455 2160 485
rect -470 425 -400 435
rect -140 440 -70 450
rect -1015 400 -995 425
rect -905 400 -885 425
rect -795 400 -775 425
rect -685 400 -665 425
rect -575 400 -555 425
rect -140 420 -135 440
rect -115 420 -95 440
rect -75 420 -70 440
rect -1025 390 -985 400
rect -1025 370 -1015 390
rect -995 370 -985 390
rect -1025 360 -985 370
rect -915 390 -875 400
rect -915 370 -905 390
rect -885 370 -875 390
rect -915 360 -875 370
rect -805 390 -765 400
rect -805 370 -795 390
rect -775 370 -765 390
rect -805 360 -765 370
rect -745 390 -715 400
rect -745 370 -740 390
rect -720 370 -715 390
rect -745 360 -715 370
rect -695 390 -655 400
rect -695 370 -685 390
rect -665 370 -655 390
rect -695 360 -655 370
rect -585 390 -545 400
rect -585 370 -575 390
rect -555 370 -545 390
rect -585 360 -545 370
rect -140 390 -70 420
rect -140 370 -135 390
rect -115 370 -95 390
rect -75 370 -70 390
rect -140 340 -70 370
rect -140 320 -135 340
rect -115 320 -95 340
rect -75 320 -70 340
rect -140 310 -70 320
rect -45 440 -15 450
rect -45 420 -40 440
rect -20 420 -15 440
rect -45 390 -15 420
rect -45 370 -40 390
rect -20 370 -15 390
rect -45 340 -15 370
rect -45 320 -40 340
rect -20 320 -15 340
rect -45 310 -15 320
rect 10 440 40 450
rect 10 420 15 440
rect 35 420 40 440
rect 10 390 40 420
rect 10 370 15 390
rect 35 370 40 390
rect 10 340 40 370
rect 10 320 15 340
rect 35 320 40 340
rect 10 310 40 320
rect 65 440 95 450
rect 65 420 70 440
rect 90 420 95 440
rect 65 390 95 420
rect 65 370 70 390
rect 90 370 95 390
rect 65 340 95 370
rect 65 320 70 340
rect 90 320 95 340
rect 65 310 95 320
rect 120 440 150 450
rect 120 420 125 440
rect 145 420 150 440
rect 120 390 150 420
rect 120 370 125 390
rect 145 370 150 390
rect 120 340 150 370
rect 120 320 125 340
rect 145 320 150 340
rect 120 310 150 320
rect 175 440 205 450
rect 175 420 180 440
rect 200 420 205 440
rect 175 390 205 420
rect 175 370 180 390
rect 200 370 205 390
rect 175 340 205 370
rect 175 320 180 340
rect 200 320 205 340
rect 175 310 205 320
rect 230 440 260 450
rect 230 420 235 440
rect 255 420 260 440
rect 230 390 260 420
rect 230 370 235 390
rect 255 370 260 390
rect 230 340 260 370
rect 230 320 235 340
rect 255 320 260 340
rect 230 310 260 320
rect 285 440 315 450
rect 285 420 290 440
rect 310 420 315 440
rect 285 390 315 420
rect 285 370 290 390
rect 310 370 315 390
rect 285 340 315 370
rect 285 320 290 340
rect 310 320 315 340
rect 285 310 315 320
rect 340 440 370 450
rect 340 420 345 440
rect 365 420 370 440
rect 340 390 370 420
rect 340 370 345 390
rect 365 370 370 390
rect 340 340 370 370
rect 340 320 345 340
rect 365 320 370 340
rect 340 310 370 320
rect 395 440 425 450
rect 395 420 400 440
rect 420 420 425 440
rect 395 390 425 420
rect 395 370 400 390
rect 420 370 425 390
rect 395 340 425 370
rect 395 320 400 340
rect 420 320 425 340
rect 395 310 425 320
rect 450 440 480 450
rect 450 420 455 440
rect 475 420 480 440
rect 450 390 480 420
rect 450 370 455 390
rect 475 370 480 390
rect 450 340 480 370
rect 450 320 455 340
rect 475 320 480 340
rect 450 310 480 320
rect 505 440 535 450
rect 505 420 510 440
rect 530 420 535 440
rect 505 390 535 420
rect 505 370 510 390
rect 530 370 535 390
rect 505 340 535 370
rect 505 320 510 340
rect 530 320 535 340
rect 505 310 535 320
rect 560 440 630 450
rect 560 420 565 440
rect 585 420 605 440
rect 625 420 630 440
rect 560 390 630 420
rect 560 370 565 390
rect 585 370 605 390
rect 625 370 630 390
rect 560 340 630 370
rect 560 320 565 340
rect 585 320 605 340
rect 625 320 630 340
rect 560 310 630 320
rect 680 440 750 450
rect 680 420 685 440
rect 705 420 725 440
rect 745 420 750 440
rect 680 390 750 420
rect 680 370 685 390
rect 705 370 725 390
rect 745 370 750 390
rect 680 340 750 370
rect 680 320 685 340
rect 705 320 725 340
rect 745 320 750 340
rect 680 310 750 320
rect 775 440 805 450
rect 775 420 780 440
rect 800 420 805 440
rect 775 390 805 420
rect 775 370 780 390
rect 800 370 805 390
rect 775 340 805 370
rect 775 320 780 340
rect 800 320 805 340
rect 775 310 805 320
rect 830 440 860 450
rect 830 420 835 440
rect 855 420 860 440
rect 830 390 860 420
rect 830 370 835 390
rect 855 370 860 390
rect 830 340 860 370
rect 830 320 835 340
rect 855 320 860 340
rect 830 310 860 320
rect 885 440 915 450
rect 885 420 890 440
rect 910 420 915 440
rect 885 390 915 420
rect 885 370 890 390
rect 910 370 915 390
rect 885 340 915 370
rect 885 320 890 340
rect 910 320 915 340
rect 885 310 915 320
rect 940 440 1010 450
rect 940 420 945 440
rect 965 420 985 440
rect 1005 420 1010 440
rect 940 390 1010 420
rect 940 370 945 390
rect 965 370 985 390
rect 1005 370 1010 390
rect 940 340 1010 370
rect 940 320 945 340
rect 965 320 985 340
rect 1005 320 1010 340
rect 940 310 1010 320
rect 1060 440 1130 450
rect 1060 420 1065 440
rect 1085 420 1105 440
rect 1125 420 1130 440
rect 1060 390 1130 420
rect 1060 370 1065 390
rect 1085 370 1105 390
rect 1125 370 1130 390
rect 1060 340 1130 370
rect 1060 320 1065 340
rect 1085 320 1105 340
rect 1125 320 1130 340
rect 1060 310 1130 320
rect 1155 440 1185 450
rect 1155 420 1160 440
rect 1180 420 1185 440
rect 1155 390 1185 420
rect 1155 370 1160 390
rect 1180 370 1185 390
rect 1155 340 1185 370
rect 1155 320 1160 340
rect 1180 320 1185 340
rect 1155 310 1185 320
rect 1210 440 1240 450
rect 1210 420 1215 440
rect 1235 420 1240 440
rect 1210 390 1240 420
rect 1210 370 1215 390
rect 1235 370 1240 390
rect 1210 340 1240 370
rect 1210 320 1215 340
rect 1235 320 1240 340
rect 1210 310 1240 320
rect 1265 440 1295 450
rect 1265 420 1270 440
rect 1290 420 1295 440
rect 1265 390 1295 420
rect 1265 370 1270 390
rect 1290 370 1295 390
rect 1265 340 1295 370
rect 1265 320 1270 340
rect 1290 320 1295 340
rect 1265 310 1295 320
rect 1320 440 1350 450
rect 1320 420 1325 440
rect 1345 420 1350 440
rect 1320 390 1350 420
rect 1320 370 1325 390
rect 1345 370 1350 390
rect 1320 340 1350 370
rect 1320 320 1325 340
rect 1345 320 1350 340
rect 1320 310 1350 320
rect 1375 440 1405 450
rect 1375 420 1380 440
rect 1400 420 1405 440
rect 1375 390 1405 420
rect 1375 370 1380 390
rect 1400 370 1405 390
rect 1375 340 1405 370
rect 1375 320 1380 340
rect 1400 320 1405 340
rect 1375 310 1405 320
rect 1430 440 1460 450
rect 1430 420 1435 440
rect 1455 420 1460 440
rect 1430 390 1460 420
rect 1430 370 1435 390
rect 1455 370 1460 390
rect 1430 340 1460 370
rect 1430 320 1435 340
rect 1455 320 1460 340
rect 1430 310 1460 320
rect 1485 440 1515 450
rect 1485 420 1490 440
rect 1510 420 1515 440
rect 1485 390 1515 420
rect 1485 370 1490 390
rect 1510 370 1515 390
rect 1485 340 1515 370
rect 1485 320 1490 340
rect 1510 320 1515 340
rect 1485 310 1515 320
rect 1540 440 1570 450
rect 1540 420 1545 440
rect 1565 420 1570 440
rect 1540 390 1570 420
rect 1540 370 1545 390
rect 1565 370 1570 390
rect 1540 340 1570 370
rect 1540 320 1545 340
rect 1565 320 1570 340
rect 1540 310 1570 320
rect 1595 440 1625 450
rect 1595 420 1600 440
rect 1620 420 1625 440
rect 1595 390 1625 420
rect 1595 370 1600 390
rect 1620 370 1625 390
rect 1595 340 1625 370
rect 1595 320 1600 340
rect 1620 320 1625 340
rect 1595 310 1625 320
rect 1650 440 1680 450
rect 1650 420 1655 440
rect 1675 420 1680 440
rect 1650 390 1680 420
rect 1650 370 1655 390
rect 1675 370 1680 390
rect 1650 340 1680 370
rect 1650 320 1655 340
rect 1675 320 1680 340
rect 1650 310 1680 320
rect 1705 440 1735 450
rect 1705 420 1710 440
rect 1730 420 1735 440
rect 1705 390 1735 420
rect 1705 370 1710 390
rect 1730 370 1735 390
rect 1705 340 1735 370
rect 1705 320 1710 340
rect 1730 320 1735 340
rect 1705 310 1735 320
rect 1760 440 1835 450
rect 1760 420 1765 440
rect 1785 420 1805 440
rect 1825 420 1835 440
rect 2090 435 2095 455
rect 2115 435 2135 455
rect 2155 435 2160 455
rect 2090 425 2160 435
rect 2185 605 2215 615
rect 2185 585 2190 605
rect 2210 585 2215 605
rect 2185 555 2215 585
rect 2185 535 2190 555
rect 2210 535 2215 555
rect 2185 505 2215 535
rect 2185 485 2190 505
rect 2210 485 2215 505
rect 2185 455 2215 485
rect 2185 435 2190 455
rect 2210 435 2215 455
rect 2185 425 2215 435
rect 2240 605 2270 615
rect 2240 585 2245 605
rect 2265 585 2270 605
rect 2240 555 2270 585
rect 2240 535 2245 555
rect 2265 535 2270 555
rect 2240 505 2270 535
rect 2240 485 2245 505
rect 2265 485 2270 505
rect 2240 455 2270 485
rect 2240 435 2245 455
rect 2265 435 2270 455
rect 2240 425 2270 435
rect 2295 605 2325 615
rect 2295 585 2300 605
rect 2320 585 2325 605
rect 2295 555 2325 585
rect 2295 535 2300 555
rect 2320 535 2325 555
rect 2295 505 2325 535
rect 2295 485 2300 505
rect 2320 485 2325 505
rect 2295 455 2325 485
rect 2295 435 2300 455
rect 2320 435 2325 455
rect 2295 425 2325 435
rect 2350 605 2380 615
rect 2350 585 2355 605
rect 2375 585 2380 605
rect 2350 555 2380 585
rect 2350 535 2355 555
rect 2375 535 2380 555
rect 2350 505 2380 535
rect 2350 485 2355 505
rect 2375 485 2380 505
rect 2350 455 2380 485
rect 2350 435 2355 455
rect 2375 435 2380 455
rect 2350 425 2380 435
rect 2405 605 2435 615
rect 2405 585 2410 605
rect 2430 585 2435 605
rect 2405 555 2435 585
rect 2405 535 2410 555
rect 2430 535 2435 555
rect 2405 505 2435 535
rect 2405 485 2410 505
rect 2430 485 2435 505
rect 2405 455 2435 485
rect 2405 435 2410 455
rect 2430 435 2435 455
rect 2405 425 2435 435
rect 2460 605 2490 615
rect 2460 585 2465 605
rect 2485 585 2490 605
rect 2460 555 2490 585
rect 2460 535 2465 555
rect 2485 535 2490 555
rect 2460 505 2490 535
rect 2460 485 2465 505
rect 2485 485 2490 505
rect 2460 455 2490 485
rect 2460 435 2465 455
rect 2485 435 2490 455
rect 2460 425 2490 435
rect 2515 605 2545 615
rect 2515 585 2520 605
rect 2540 585 2545 605
rect 2515 555 2545 585
rect 2515 535 2520 555
rect 2540 535 2545 555
rect 2515 505 2545 535
rect 2515 485 2520 505
rect 2540 485 2545 505
rect 2515 455 2545 485
rect 2515 435 2520 455
rect 2540 435 2545 455
rect 2515 425 2545 435
rect 2570 605 2600 615
rect 2570 585 2575 605
rect 2595 585 2600 605
rect 2570 555 2600 585
rect 2570 535 2575 555
rect 2595 535 2600 555
rect 2570 505 2600 535
rect 2570 485 2575 505
rect 2595 485 2600 505
rect 2570 455 2600 485
rect 2570 435 2575 455
rect 2595 435 2600 455
rect 2570 425 2600 435
rect 2625 605 2655 615
rect 2625 585 2630 605
rect 2650 585 2655 605
rect 2625 555 2655 585
rect 2625 535 2630 555
rect 2650 535 2655 555
rect 2625 505 2655 535
rect 2625 485 2630 505
rect 2650 485 2655 505
rect 2625 455 2655 485
rect 2625 435 2630 455
rect 2650 435 2655 455
rect 2625 425 2655 435
rect 2680 605 2710 615
rect 2680 585 2685 605
rect 2705 585 2710 605
rect 2680 555 2710 585
rect 2680 535 2685 555
rect 2705 535 2710 555
rect 2680 505 2710 535
rect 2680 485 2685 505
rect 2705 485 2710 505
rect 2680 455 2710 485
rect 2680 435 2685 455
rect 2705 435 2710 455
rect 2680 425 2710 435
rect 2735 605 2765 615
rect 2735 585 2740 605
rect 2760 585 2765 605
rect 2735 555 2765 585
rect 2735 535 2740 555
rect 2760 535 2765 555
rect 2735 505 2765 535
rect 2735 485 2740 505
rect 2760 485 2765 505
rect 2735 455 2765 485
rect 2735 435 2740 455
rect 2760 435 2765 455
rect 2735 425 2765 435
rect 2790 605 2860 615
rect 2790 585 2795 605
rect 2815 585 2835 605
rect 2855 585 2860 605
rect 2790 555 2860 585
rect 2790 535 2795 555
rect 2815 535 2835 555
rect 2855 535 2860 555
rect 2790 505 2860 535
rect 2790 485 2795 505
rect 2815 485 2835 505
rect 2855 485 2860 505
rect 2790 455 2860 485
rect 2790 435 2795 455
rect 2815 435 2835 455
rect 2855 435 2860 455
rect 2790 425 2860 435
rect 2965 537 3180 572
rect 2965 517 3000 537
rect 3145 517 3180 537
rect 1760 390 1835 420
rect 2245 400 2265 425
rect 2355 400 2375 425
rect 2465 400 2485 425
rect 2575 400 2595 425
rect 2685 400 2705 425
rect 1760 370 1765 390
rect 1785 370 1805 390
rect 1825 370 1835 390
rect 1760 340 1835 370
rect 2235 390 2275 400
rect 2235 370 2245 390
rect 2265 370 2275 390
rect 2235 360 2275 370
rect 2345 390 2385 400
rect 2345 370 2355 390
rect 2375 370 2385 390
rect 2345 360 2385 370
rect 2405 390 2435 400
rect 2405 370 2410 390
rect 2430 370 2435 390
rect 2405 360 2435 370
rect 2455 390 2495 400
rect 2455 370 2465 390
rect 2485 370 2495 390
rect 2455 360 2495 370
rect 2565 390 2605 400
rect 2565 370 2575 390
rect 2595 370 2605 390
rect 2565 360 2605 370
rect 2675 390 2715 400
rect 2675 370 2685 390
rect 2705 370 2715 390
rect 2675 360 2715 370
rect 1760 320 1765 340
rect 1785 320 1805 340
rect 1825 320 1835 340
rect 1760 310 1835 320
rect -95 290 -75 310
rect 15 290 35 310
rect 125 290 145 310
rect 235 290 255 310
rect 345 290 365 310
rect 455 290 475 310
rect 605 290 625 310
rect 780 290 800 310
rect 835 290 855 310
rect 890 290 910 310
rect 1065 290 1085 310
rect 1215 290 1235 310
rect 1325 290 1345 310
rect 1435 290 1455 310
rect 1545 290 1565 310
rect 1655 290 1675 310
rect 1765 290 1785 310
rect 3060 467 3085 517
rect -1025 280 -985 290
rect -1025 260 -1015 280
rect -995 260 -985 280
rect -1025 250 -985 260
rect -915 280 -875 290
rect -915 260 -905 280
rect -885 260 -875 280
rect -915 250 -875 260
rect -805 280 -765 290
rect -805 260 -795 280
rect -775 260 -765 280
rect -805 250 -765 260
rect -745 280 -715 290
rect -745 260 -740 280
rect -720 260 -715 280
rect -745 250 -715 260
rect -695 280 -655 290
rect -695 260 -685 280
rect -665 260 -655 280
rect -695 250 -655 260
rect -585 280 -545 290
rect -585 260 -575 280
rect -555 260 -545 280
rect -585 250 -545 260
rect -100 280 -70 290
rect -100 260 -95 280
rect -75 260 -70 280
rect -100 250 -70 260
rect 5 280 45 290
rect 5 260 15 280
rect 35 260 45 280
rect 5 250 45 260
rect 115 280 155 290
rect 115 260 125 280
rect 145 260 155 280
rect 115 250 155 260
rect 225 280 265 290
rect 225 260 235 280
rect 255 260 265 280
rect 225 250 265 260
rect 335 280 375 290
rect 335 260 345 280
rect 365 260 375 280
rect 335 250 375 260
rect 445 280 485 290
rect 445 260 455 280
rect 475 260 485 280
rect 445 250 485 260
rect 600 280 630 290
rect 600 260 605 280
rect 625 260 630 280
rect 600 250 630 260
rect 775 280 805 290
rect 775 260 780 280
rect 800 260 805 280
rect 775 250 805 260
rect 830 280 860 290
rect 830 260 835 280
rect 855 260 860 280
rect 830 250 860 260
rect 885 280 915 290
rect 885 260 890 280
rect 910 260 915 280
rect 885 250 915 260
rect 1060 280 1090 290
rect 1060 260 1065 280
rect 1085 260 1090 280
rect 1060 250 1090 260
rect 1205 280 1245 290
rect 1205 260 1215 280
rect 1235 260 1245 280
rect 1205 250 1245 260
rect 1315 280 1355 290
rect 1315 260 1325 280
rect 1345 260 1355 280
rect 1315 250 1355 260
rect 1425 280 1465 290
rect 1425 260 1435 280
rect 1455 260 1465 280
rect 1425 250 1465 260
rect 1535 280 1575 290
rect 1535 260 1545 280
rect 1565 260 1575 280
rect 1535 250 1575 260
rect 1645 280 1685 290
rect 1645 260 1655 280
rect 1675 260 1685 280
rect 1645 250 1685 260
rect 1760 280 1790 290
rect 1760 260 1765 280
rect 1785 260 1790 280
rect 1760 250 1790 260
rect 2235 280 2275 290
rect 2235 260 2245 280
rect 2265 260 2275 280
rect 2235 250 2275 260
rect 2345 280 2385 290
rect 2345 260 2355 280
rect 2375 260 2385 280
rect 2345 250 2385 260
rect 2405 280 2435 290
rect 2405 260 2410 280
rect 2430 260 2435 280
rect 2405 250 2435 260
rect 2455 280 2495 290
rect 2455 260 2465 280
rect 2485 260 2495 280
rect 2455 250 2495 260
rect 2565 280 2605 290
rect 2565 260 2575 280
rect 2595 260 2605 280
rect 2565 250 2605 260
rect 2675 280 2715 290
rect 2675 260 2685 280
rect 2705 260 2715 280
rect 2675 250 2715 260
rect -1015 225 -995 250
rect -905 225 -885 250
rect -795 225 -775 250
rect -685 225 -665 250
rect -575 225 -555 250
rect 2245 225 2265 250
rect 2355 225 2375 250
rect 2465 225 2485 250
rect 2575 225 2595 250
rect 2685 225 2705 250
rect -1170 215 -1100 225
rect -1170 195 -1165 215
rect -1145 195 -1125 215
rect -1105 195 -1100 215
rect -1170 165 -1100 195
rect -1170 145 -1165 165
rect -1145 145 -1125 165
rect -1105 145 -1100 165
rect -1490 -93 -1455 -85
rect -1490 -113 -1485 -93
rect -1460 -113 -1455 -93
rect -1490 -120 -1455 -113
rect -1430 -93 -1395 -85
rect -1430 -113 -1425 -93
rect -1400 -113 -1395 -93
rect -1430 -120 -1395 -113
rect -1370 -93 -1335 -85
rect -1370 -113 -1365 -93
rect -1340 -113 -1335 -93
rect -1370 -120 -1335 -113
rect -1170 115 -1100 145
rect -1170 95 -1165 115
rect -1145 95 -1125 115
rect -1105 95 -1100 115
rect -1170 65 -1100 95
rect -1170 45 -1165 65
rect -1145 45 -1125 65
rect -1105 45 -1100 65
rect -1170 15 -1100 45
rect -1170 -5 -1165 15
rect -1145 -5 -1125 15
rect -1105 -5 -1100 15
rect -1170 -35 -1100 -5
rect -1170 -55 -1165 -35
rect -1145 -55 -1125 -35
rect -1105 -55 -1100 -35
rect -1170 -65 -1100 -55
rect -1075 215 -1045 225
rect -1075 195 -1070 215
rect -1050 195 -1045 215
rect -1075 165 -1045 195
rect -1075 145 -1070 165
rect -1050 145 -1045 165
rect -1075 115 -1045 145
rect -1075 95 -1070 115
rect -1050 95 -1045 115
rect -1075 65 -1045 95
rect -1075 45 -1070 65
rect -1050 45 -1045 65
rect -1075 15 -1045 45
rect -1075 -5 -1070 15
rect -1050 -5 -1045 15
rect -1075 -35 -1045 -5
rect -1075 -55 -1070 -35
rect -1050 -55 -1045 -35
rect -1075 -65 -1045 -55
rect -1020 215 -990 225
rect -1020 195 -1015 215
rect -995 195 -990 215
rect -1020 165 -990 195
rect -1020 145 -1015 165
rect -995 145 -990 165
rect -1020 115 -990 145
rect -1020 95 -1015 115
rect -995 95 -990 115
rect -1020 65 -990 95
rect -1020 45 -1015 65
rect -995 45 -990 65
rect -1020 15 -990 45
rect -1020 -5 -1015 15
rect -995 -5 -990 15
rect -1020 -35 -990 -5
rect -1020 -55 -1015 -35
rect -995 -55 -990 -35
rect -1020 -65 -990 -55
rect -965 215 -935 225
rect -965 195 -960 215
rect -940 195 -935 215
rect -965 165 -935 195
rect -965 145 -960 165
rect -940 145 -935 165
rect -965 115 -935 145
rect -965 95 -960 115
rect -940 95 -935 115
rect -965 65 -935 95
rect -965 45 -960 65
rect -940 45 -935 65
rect -965 15 -935 45
rect -965 -5 -960 15
rect -940 -5 -935 15
rect -965 -35 -935 -5
rect -965 -55 -960 -35
rect -940 -55 -935 -35
rect -965 -65 -935 -55
rect -910 215 -880 225
rect -910 195 -905 215
rect -885 195 -880 215
rect -910 165 -880 195
rect -910 145 -905 165
rect -885 145 -880 165
rect -910 115 -880 145
rect -910 95 -905 115
rect -885 95 -880 115
rect -910 65 -880 95
rect -910 45 -905 65
rect -885 45 -880 65
rect -910 15 -880 45
rect -910 -5 -905 15
rect -885 -5 -880 15
rect -910 -35 -880 -5
rect -910 -55 -905 -35
rect -885 -55 -880 -35
rect -910 -65 -880 -55
rect -855 215 -825 225
rect -855 195 -850 215
rect -830 195 -825 215
rect -855 165 -825 195
rect -855 145 -850 165
rect -830 145 -825 165
rect -855 115 -825 145
rect -855 95 -850 115
rect -830 95 -825 115
rect -855 65 -825 95
rect -855 45 -850 65
rect -830 45 -825 65
rect -855 15 -825 45
rect -855 -5 -850 15
rect -830 -5 -825 15
rect -855 -35 -825 -5
rect -855 -55 -850 -35
rect -830 -55 -825 -35
rect -855 -65 -825 -55
rect -800 215 -770 225
rect -800 195 -795 215
rect -775 195 -770 215
rect -800 165 -770 195
rect -800 145 -795 165
rect -775 145 -770 165
rect -800 115 -770 145
rect -800 95 -795 115
rect -775 95 -770 115
rect -800 65 -770 95
rect -800 45 -795 65
rect -775 45 -770 65
rect -800 15 -770 45
rect -800 -5 -795 15
rect -775 -5 -770 15
rect -800 -35 -770 -5
rect -800 -55 -795 -35
rect -775 -55 -770 -35
rect -800 -65 -770 -55
rect -745 215 -715 225
rect -745 195 -740 215
rect -720 195 -715 215
rect -745 165 -715 195
rect -745 145 -740 165
rect -720 145 -715 165
rect -745 115 -715 145
rect -745 95 -740 115
rect -720 95 -715 115
rect -745 65 -715 95
rect -745 45 -740 65
rect -720 45 -715 65
rect -745 15 -715 45
rect -745 -5 -740 15
rect -720 -5 -715 15
rect -745 -35 -715 -5
rect -745 -55 -740 -35
rect -720 -55 -715 -35
rect -745 -65 -715 -55
rect -690 215 -660 225
rect -690 195 -685 215
rect -665 195 -660 215
rect -690 165 -660 195
rect -690 145 -685 165
rect -665 145 -660 165
rect -690 115 -660 145
rect -690 95 -685 115
rect -665 95 -660 115
rect -690 65 -660 95
rect -690 45 -685 65
rect -665 45 -660 65
rect -690 15 -660 45
rect -690 -5 -685 15
rect -665 -5 -660 15
rect -690 -35 -660 -5
rect -690 -55 -685 -35
rect -665 -55 -660 -35
rect -690 -65 -660 -55
rect -635 215 -605 225
rect -635 195 -630 215
rect -610 195 -605 215
rect -635 165 -605 195
rect -635 145 -630 165
rect -610 145 -605 165
rect -635 115 -605 145
rect -635 95 -630 115
rect -610 95 -605 115
rect -635 65 -605 95
rect -635 45 -630 65
rect -610 45 -605 65
rect -635 15 -605 45
rect -635 -5 -630 15
rect -610 -5 -605 15
rect -635 -35 -605 -5
rect -635 -55 -630 -35
rect -610 -55 -605 -35
rect -635 -65 -605 -55
rect -580 215 -550 225
rect -580 195 -575 215
rect -555 195 -550 215
rect -580 165 -550 195
rect -580 145 -575 165
rect -555 145 -550 165
rect -580 115 -550 145
rect -580 95 -575 115
rect -555 95 -550 115
rect -580 65 -550 95
rect -580 45 -575 65
rect -555 45 -550 65
rect -580 15 -550 45
rect -580 -5 -575 15
rect -555 -5 -550 15
rect -580 -35 -550 -5
rect -580 -55 -575 -35
rect -555 -55 -550 -35
rect -580 -65 -550 -55
rect -525 215 -495 225
rect -525 195 -520 215
rect -500 195 -495 215
rect -525 165 -495 195
rect -525 145 -520 165
rect -500 145 -495 165
rect -525 115 -495 145
rect -525 95 -520 115
rect -500 95 -495 115
rect -525 65 -495 95
rect -525 45 -520 65
rect -500 45 -495 65
rect -525 15 -495 45
rect -525 -5 -520 15
rect -500 -5 -495 15
rect -525 -35 -495 -5
rect -525 -55 -520 -35
rect -500 -55 -495 -35
rect -525 -65 -495 -55
rect -470 215 -400 225
rect -470 195 -465 215
rect -445 195 -425 215
rect -405 195 -400 215
rect -470 165 -400 195
rect -470 145 -465 165
rect -445 145 -425 165
rect -405 145 -400 165
rect -470 115 -400 145
rect -470 95 -465 115
rect -445 95 -425 115
rect -405 95 -400 115
rect -470 65 -400 95
rect -470 45 -465 65
rect -445 45 -425 65
rect -405 45 -400 65
rect -470 15 -400 45
rect 2090 215 2160 225
rect 2090 195 2095 215
rect 2115 195 2135 215
rect 2155 195 2160 215
rect 2090 165 2160 195
rect 2090 145 2095 165
rect 2115 145 2135 165
rect 2155 145 2160 165
rect 2090 115 2160 145
rect 2090 95 2095 115
rect 2115 95 2135 115
rect 2155 95 2160 115
rect 2090 65 2160 95
rect 2090 45 2095 65
rect 2115 45 2135 65
rect 2155 45 2160 65
rect -470 -5 -465 15
rect -445 -5 -425 15
rect -405 -5 -400 15
rect -470 -35 -400 -5
rect 775 5 805 15
rect 775 -15 780 5
rect 800 -15 805 5
rect 775 -25 805 -15
rect 830 10 860 20
rect 2090 15 2160 45
rect 830 -10 835 10
rect 855 -10 860 10
rect 830 -20 860 -10
rect 885 5 915 15
rect 885 -15 890 5
rect 910 -15 915 5
rect 885 -25 915 -15
rect 2090 -5 2095 15
rect 2115 -5 2135 15
rect 2155 -5 2160 15
rect -470 -55 -465 -35
rect -445 -55 -425 -35
rect -405 -55 -400 -35
rect 780 -45 800 -25
rect 890 -45 910 -25
rect 2090 -35 2160 -5
rect -470 -65 -400 -55
rect 680 -55 750 -45
rect -1125 -85 -1105 -65
rect -1070 -85 -1050 -65
rect -960 -85 -940 -65
rect -850 -85 -830 -65
rect -740 -85 -720 -65
rect -630 -85 -610 -65
rect -520 -85 -500 -65
rect -465 -85 -445 -65
rect 680 -75 685 -55
rect 705 -75 725 -55
rect 745 -75 750 -55
rect -1310 -93 -1275 -85
rect -1310 -113 -1305 -93
rect -1280 -113 -1275 -93
rect -1310 -120 -1275 -113
rect -1145 -95 -1105 -85
rect -1145 -115 -1135 -95
rect -1115 -115 -1105 -95
rect -1145 -125 -1105 -115
rect -1080 -95 -1040 -85
rect -1080 -115 -1070 -95
rect -1050 -115 -1040 -95
rect -1080 -125 -1040 -115
rect -970 -95 -930 -85
rect -970 -115 -960 -95
rect -940 -115 -930 -95
rect -970 -125 -930 -115
rect -860 -95 -820 -85
rect -860 -115 -850 -95
rect -830 -115 -820 -95
rect -860 -125 -820 -115
rect -750 -95 -710 -85
rect -750 -115 -740 -95
rect -720 -115 -710 -95
rect -750 -125 -710 -115
rect -640 -95 -600 -85
rect -640 -115 -630 -95
rect -610 -115 -600 -95
rect -640 -125 -600 -115
rect -530 -95 -490 -85
rect -530 -115 -520 -95
rect -500 -115 -490 -95
rect -530 -125 -490 -115
rect -465 -95 -425 -85
rect -465 -115 -455 -95
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect 680 -105 750 -75
rect 680 -125 685 -105
rect 705 -125 725 -105
rect 745 -125 750 -105
rect 680 -155 750 -125
rect 680 -175 685 -155
rect 705 -175 725 -155
rect 745 -175 750 -155
rect 680 -205 750 -175
rect 680 -225 685 -205
rect 705 -225 725 -205
rect 745 -225 750 -205
rect 680 -255 750 -225
rect 680 -275 685 -255
rect 705 -275 725 -255
rect 745 -275 750 -255
rect 680 -285 750 -275
rect 775 -55 805 -45
rect 775 -75 780 -55
rect 800 -75 805 -55
rect 775 -105 805 -75
rect 775 -125 780 -105
rect 800 -125 805 -105
rect 775 -155 805 -125
rect 775 -175 780 -155
rect 800 -175 805 -155
rect 775 -205 805 -175
rect 775 -225 780 -205
rect 800 -225 805 -205
rect 775 -255 805 -225
rect 775 -275 780 -255
rect 800 -275 805 -255
rect 775 -285 805 -275
rect 830 -55 860 -45
rect 830 -75 835 -55
rect 855 -75 860 -55
rect 830 -105 860 -75
rect 830 -125 835 -105
rect 855 -125 860 -105
rect 830 -155 860 -125
rect 830 -175 835 -155
rect 855 -175 860 -155
rect 830 -205 860 -175
rect 830 -225 835 -205
rect 855 -225 860 -205
rect 830 -255 860 -225
rect 830 -275 835 -255
rect 855 -275 860 -255
rect 830 -285 860 -275
rect 885 -55 915 -45
rect 885 -75 890 -55
rect 910 -75 915 -55
rect 885 -105 915 -75
rect 885 -125 890 -105
rect 910 -125 915 -105
rect 885 -155 915 -125
rect 885 -175 890 -155
rect 910 -175 915 -155
rect 885 -205 915 -175
rect 885 -225 890 -205
rect 910 -225 915 -205
rect 885 -255 915 -225
rect 885 -275 890 -255
rect 910 -275 915 -255
rect 885 -285 915 -275
rect 940 -55 1010 -45
rect 940 -75 945 -55
rect 965 -75 985 -55
rect 1005 -75 1010 -55
rect 2090 -55 2095 -35
rect 2115 -55 2135 -35
rect 2155 -55 2160 -35
rect 2090 -65 2160 -55
rect 2185 215 2215 225
rect 2185 195 2190 215
rect 2210 195 2215 215
rect 2185 165 2215 195
rect 2185 145 2190 165
rect 2210 145 2215 165
rect 2185 115 2215 145
rect 2185 95 2190 115
rect 2210 95 2215 115
rect 2185 65 2215 95
rect 2185 45 2190 65
rect 2210 45 2215 65
rect 2185 15 2215 45
rect 2185 -5 2190 15
rect 2210 -5 2215 15
rect 2185 -35 2215 -5
rect 2185 -55 2190 -35
rect 2210 -55 2215 -35
rect 2185 -65 2215 -55
rect 2240 215 2270 225
rect 2240 195 2245 215
rect 2265 195 2270 215
rect 2240 165 2270 195
rect 2240 145 2245 165
rect 2265 145 2270 165
rect 2240 115 2270 145
rect 2240 95 2245 115
rect 2265 95 2270 115
rect 2240 65 2270 95
rect 2240 45 2245 65
rect 2265 45 2270 65
rect 2240 15 2270 45
rect 2240 -5 2245 15
rect 2265 -5 2270 15
rect 2240 -35 2270 -5
rect 2240 -55 2245 -35
rect 2265 -55 2270 -35
rect 2240 -65 2270 -55
rect 2295 215 2325 225
rect 2295 195 2300 215
rect 2320 195 2325 215
rect 2295 165 2325 195
rect 2295 145 2300 165
rect 2320 145 2325 165
rect 2295 115 2325 145
rect 2295 95 2300 115
rect 2320 95 2325 115
rect 2295 65 2325 95
rect 2295 45 2300 65
rect 2320 45 2325 65
rect 2295 15 2325 45
rect 2295 -5 2300 15
rect 2320 -5 2325 15
rect 2295 -35 2325 -5
rect 2295 -55 2300 -35
rect 2320 -55 2325 -35
rect 2295 -65 2325 -55
rect 2350 215 2380 225
rect 2350 195 2355 215
rect 2375 195 2380 215
rect 2350 165 2380 195
rect 2350 145 2355 165
rect 2375 145 2380 165
rect 2350 115 2380 145
rect 2350 95 2355 115
rect 2375 95 2380 115
rect 2350 65 2380 95
rect 2350 45 2355 65
rect 2375 45 2380 65
rect 2350 15 2380 45
rect 2350 -5 2355 15
rect 2375 -5 2380 15
rect 2350 -35 2380 -5
rect 2350 -55 2355 -35
rect 2375 -55 2380 -35
rect 2350 -65 2380 -55
rect 2405 215 2435 225
rect 2405 195 2410 215
rect 2430 195 2435 215
rect 2405 165 2435 195
rect 2405 145 2410 165
rect 2430 145 2435 165
rect 2405 115 2435 145
rect 2405 95 2410 115
rect 2430 95 2435 115
rect 2405 65 2435 95
rect 2405 45 2410 65
rect 2430 45 2435 65
rect 2405 15 2435 45
rect 2405 -5 2410 15
rect 2430 -5 2435 15
rect 2405 -35 2435 -5
rect 2405 -55 2410 -35
rect 2430 -55 2435 -35
rect 2405 -65 2435 -55
rect 2460 215 2490 225
rect 2460 195 2465 215
rect 2485 195 2490 215
rect 2460 165 2490 195
rect 2460 145 2465 165
rect 2485 145 2490 165
rect 2460 115 2490 145
rect 2460 95 2465 115
rect 2485 95 2490 115
rect 2460 65 2490 95
rect 2460 45 2465 65
rect 2485 45 2490 65
rect 2460 15 2490 45
rect 2460 -5 2465 15
rect 2485 -5 2490 15
rect 2460 -35 2490 -5
rect 2460 -55 2465 -35
rect 2485 -55 2490 -35
rect 2460 -65 2490 -55
rect 2515 215 2545 225
rect 2515 195 2520 215
rect 2540 195 2545 215
rect 2515 165 2545 195
rect 2515 145 2520 165
rect 2540 145 2545 165
rect 2515 115 2545 145
rect 2515 95 2520 115
rect 2540 95 2545 115
rect 2515 65 2545 95
rect 2515 45 2520 65
rect 2540 45 2545 65
rect 2515 15 2545 45
rect 2515 -5 2520 15
rect 2540 -5 2545 15
rect 2515 -35 2545 -5
rect 2515 -55 2520 -35
rect 2540 -55 2545 -35
rect 2515 -65 2545 -55
rect 2570 215 2600 225
rect 2570 195 2575 215
rect 2595 195 2600 215
rect 2570 165 2600 195
rect 2570 145 2575 165
rect 2595 145 2600 165
rect 2570 115 2600 145
rect 2570 95 2575 115
rect 2595 95 2600 115
rect 2570 65 2600 95
rect 2570 45 2575 65
rect 2595 45 2600 65
rect 2570 15 2600 45
rect 2570 -5 2575 15
rect 2595 -5 2600 15
rect 2570 -35 2600 -5
rect 2570 -55 2575 -35
rect 2595 -55 2600 -35
rect 2570 -65 2600 -55
rect 2625 215 2655 225
rect 2625 195 2630 215
rect 2650 195 2655 215
rect 2625 165 2655 195
rect 2625 145 2630 165
rect 2650 145 2655 165
rect 2625 115 2655 145
rect 2625 95 2630 115
rect 2650 95 2655 115
rect 2625 65 2655 95
rect 2625 45 2630 65
rect 2650 45 2655 65
rect 2625 15 2655 45
rect 2625 -5 2630 15
rect 2650 -5 2655 15
rect 2625 -35 2655 -5
rect 2625 -55 2630 -35
rect 2650 -55 2655 -35
rect 2625 -65 2655 -55
rect 2680 215 2710 225
rect 2680 195 2685 215
rect 2705 195 2710 215
rect 2680 165 2710 195
rect 2680 145 2685 165
rect 2705 145 2710 165
rect 2680 115 2710 145
rect 2680 95 2685 115
rect 2705 95 2710 115
rect 2680 65 2710 95
rect 2680 45 2685 65
rect 2705 45 2710 65
rect 2680 15 2710 45
rect 2680 -5 2685 15
rect 2705 -5 2710 15
rect 2680 -35 2710 -5
rect 2680 -55 2685 -35
rect 2705 -55 2710 -35
rect 2680 -65 2710 -55
rect 2735 215 2765 225
rect 2735 195 2740 215
rect 2760 195 2765 215
rect 2735 165 2765 195
rect 2735 145 2740 165
rect 2760 145 2765 165
rect 2735 115 2765 145
rect 2735 95 2740 115
rect 2760 95 2765 115
rect 2735 65 2765 95
rect 2735 45 2740 65
rect 2760 45 2765 65
rect 2735 15 2765 45
rect 2735 -5 2740 15
rect 2760 -5 2765 15
rect 2735 -35 2765 -5
rect 2735 -55 2740 -35
rect 2760 -55 2765 -35
rect 2735 -65 2765 -55
rect 2790 215 2860 225
rect 2790 195 2795 215
rect 2815 195 2835 215
rect 2855 195 2860 215
rect 2790 165 2860 195
rect 2790 145 2795 165
rect 2815 145 2835 165
rect 2855 145 2860 165
rect 2790 115 2860 145
rect 2790 95 2795 115
rect 2815 95 2835 115
rect 2855 95 2860 115
rect 2790 65 2860 95
rect 2790 45 2795 65
rect 2815 45 2835 65
rect 2855 45 2860 65
rect 2790 15 2860 45
rect 2790 -5 2795 15
rect 2815 -5 2835 15
rect 2855 -5 2860 15
rect 2790 -35 2860 -5
rect 2790 -55 2795 -35
rect 2815 -55 2835 -35
rect 2855 -55 2860 -35
rect 2790 -65 2860 -55
rect 940 -105 1010 -75
rect 2135 -85 2155 -65
rect 2190 -85 2210 -65
rect 2300 -85 2320 -65
rect 2410 -85 2430 -65
rect 2520 -85 2540 -65
rect 2630 -85 2650 -65
rect 2740 -85 2760 -65
rect 2795 -85 2815 -65
rect 940 -125 945 -105
rect 965 -125 985 -105
rect 1005 -125 1010 -105
rect 2115 -95 2155 -85
rect 2115 -115 2125 -95
rect 2145 -115 2155 -95
rect 2115 -125 2155 -115
rect 2180 -95 2220 -85
rect 2180 -115 2190 -95
rect 2210 -115 2220 -95
rect 2180 -125 2220 -115
rect 2290 -95 2330 -85
rect 2290 -115 2300 -95
rect 2320 -115 2330 -95
rect 2290 -125 2330 -115
rect 2400 -95 2440 -85
rect 2400 -115 2410 -95
rect 2430 -115 2440 -95
rect 2400 -125 2440 -115
rect 2510 -95 2550 -85
rect 2510 -115 2520 -95
rect 2540 -115 2550 -95
rect 2510 -125 2550 -115
rect 2620 -95 2660 -85
rect 2620 -115 2630 -95
rect 2650 -115 2660 -95
rect 2620 -125 2660 -115
rect 2730 -95 2770 -85
rect 2730 -115 2740 -95
rect 2760 -115 2770 -95
rect 2730 -125 2770 -115
rect 2795 -95 2835 -85
rect 2795 -115 2805 -95
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect 2965 -93 3000 -85
rect 2965 -113 2970 -93
rect 2995 -113 3000 -93
rect 2965 -120 3000 -113
rect 3025 -93 3060 -85
rect 3025 -113 3030 -93
rect 3055 -113 3060 -93
rect 3025 -120 3060 -113
rect 3085 -93 3120 -85
rect 3085 -113 3090 -93
rect 3115 -113 3120 -93
rect 3085 -120 3120 -113
rect 3145 -93 3180 -85
rect 3145 -113 3150 -93
rect 3175 -113 3180 -93
rect 3145 -120 3180 -113
rect 940 -155 1010 -125
rect 940 -175 945 -155
rect 965 -175 985 -155
rect 1005 -175 1010 -155
rect 940 -205 1010 -175
rect 940 -225 945 -205
rect 965 -225 985 -205
rect 1005 -225 1010 -205
rect 940 -255 1010 -225
rect 940 -275 945 -255
rect 965 -275 985 -255
rect 1005 -275 1010 -255
rect 940 -285 1010 -275
rect -925 -305 -885 -295
rect -925 -325 -915 -305
rect -895 -325 -885 -305
rect -925 -335 -885 -325
rect -725 -305 -685 -295
rect -725 -325 -715 -305
rect -695 -325 -685 -305
rect -725 -335 -685 -325
rect -625 -305 -585 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -335 -585 -325
rect -525 -305 -485 -295
rect 725 -305 745 -285
rect 835 -305 855 -285
rect 945 -305 965 -285
rect 2175 -305 2215 -295
rect -525 -325 -515 -305
rect -495 -325 -485 -305
rect -525 -335 -485 -325
rect 715 -315 755 -305
rect 715 -335 725 -315
rect 745 -335 755 -315
rect -915 -360 -895 -335
rect -715 -360 -695 -335
rect -515 -360 -495 -335
rect 715 -345 755 -335
rect 825 -315 865 -305
rect 825 -335 835 -315
rect 855 -335 865 -315
rect 825 -345 865 -335
rect 935 -315 975 -305
rect 935 -335 945 -315
rect 965 -335 975 -315
rect 2175 -325 2185 -305
rect 2205 -325 2215 -305
rect 2175 -335 2215 -325
rect 2275 -305 2315 -295
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -335 2315 -325
rect 2375 -305 2415 -295
rect 2375 -325 2385 -305
rect 2405 -325 2415 -305
rect 2375 -335 2415 -325
rect 2575 -305 2615 -295
rect 2575 -325 2585 -305
rect 2605 -325 2615 -305
rect 2575 -335 2615 -325
rect 935 -345 975 -335
rect 2185 -360 2205 -335
rect 2385 -360 2405 -335
rect 2585 -360 2605 -335
rect -1060 -370 -990 -360
rect -1210 -387 -1175 -380
rect -1210 -407 -1205 -387
rect -1180 -407 -1175 -387
rect -1210 -415 -1175 -407
rect -1150 -387 -1115 -380
rect -1150 -407 -1145 -387
rect -1120 -407 -1115 -387
rect -1150 -415 -1115 -407
rect -1060 -390 -1055 -370
rect -1035 -390 -1015 -370
rect -995 -390 -990 -370
rect -1060 -420 -990 -390
rect -1060 -440 -1055 -420
rect -1035 -440 -1015 -420
rect -995 -440 -990 -420
rect -1060 -470 -990 -440
rect -1060 -490 -1055 -470
rect -1035 -490 -1015 -470
rect -995 -490 -990 -470
rect -1060 -520 -990 -490
rect -1060 -540 -1055 -520
rect -1035 -540 -1015 -520
rect -995 -540 -990 -520
rect -1060 -570 -990 -540
rect -1060 -590 -1055 -570
rect -1035 -590 -1015 -570
rect -995 -590 -990 -570
rect -1060 -620 -990 -590
rect -1060 -640 -1055 -620
rect -1035 -640 -1015 -620
rect -995 -640 -990 -620
rect -1060 -670 -990 -640
rect -1060 -690 -1055 -670
rect -1035 -690 -1015 -670
rect -995 -690 -990 -670
rect -1060 -720 -990 -690
rect -1060 -740 -1055 -720
rect -1035 -740 -1015 -720
rect -995 -740 -990 -720
rect -1060 -770 -990 -740
rect -1060 -790 -1055 -770
rect -1035 -790 -1015 -770
rect -995 -790 -990 -770
rect -1060 -820 -990 -790
rect -1060 -840 -1055 -820
rect -1035 -840 -1015 -820
rect -995 -840 -990 -820
rect -1060 -870 -990 -840
rect -1175 -1105 -1150 -1055
rect -1060 -890 -1055 -870
rect -1035 -890 -1015 -870
rect -995 -890 -990 -870
rect -1060 -920 -990 -890
rect -1060 -940 -1055 -920
rect -1035 -940 -1015 -920
rect -995 -940 -990 -920
rect -1060 -970 -990 -940
rect -1060 -990 -1055 -970
rect -1035 -990 -1015 -970
rect -995 -990 -990 -970
rect -1060 -1020 -990 -990
rect -1060 -1040 -1055 -1020
rect -1035 -1040 -1015 -1020
rect -995 -1040 -990 -1020
rect -1060 -1050 -990 -1040
rect -920 -370 -890 -360
rect -920 -390 -915 -370
rect -895 -390 -890 -370
rect -920 -420 -890 -390
rect -920 -440 -915 -420
rect -895 -440 -890 -420
rect -920 -470 -890 -440
rect -920 -490 -915 -470
rect -895 -490 -890 -470
rect -920 -520 -890 -490
rect -920 -540 -915 -520
rect -895 -540 -890 -520
rect -920 -570 -890 -540
rect -920 -590 -915 -570
rect -895 -590 -890 -570
rect -920 -620 -890 -590
rect -920 -640 -915 -620
rect -895 -640 -890 -620
rect -920 -670 -890 -640
rect -920 -690 -915 -670
rect -895 -690 -890 -670
rect -920 -720 -890 -690
rect -920 -740 -915 -720
rect -895 -740 -890 -720
rect -920 -770 -890 -740
rect -920 -790 -915 -770
rect -895 -790 -890 -770
rect -920 -820 -890 -790
rect -920 -840 -915 -820
rect -895 -840 -890 -820
rect -920 -870 -890 -840
rect -920 -890 -915 -870
rect -895 -890 -890 -870
rect -920 -920 -890 -890
rect -920 -940 -915 -920
rect -895 -940 -890 -920
rect -920 -970 -890 -940
rect -920 -990 -915 -970
rect -895 -990 -890 -970
rect -920 -1020 -890 -990
rect -920 -1040 -915 -1020
rect -895 -1040 -890 -1020
rect -920 -1050 -890 -1040
rect -820 -370 -790 -360
rect -820 -390 -815 -370
rect -795 -390 -790 -370
rect -820 -420 -790 -390
rect -820 -440 -815 -420
rect -795 -440 -790 -420
rect -820 -470 -790 -440
rect -820 -490 -815 -470
rect -795 -490 -790 -470
rect -820 -520 -790 -490
rect -820 -540 -815 -520
rect -795 -540 -790 -520
rect -820 -570 -790 -540
rect -820 -590 -815 -570
rect -795 -590 -790 -570
rect -820 -620 -790 -590
rect -820 -640 -815 -620
rect -795 -640 -790 -620
rect -820 -670 -790 -640
rect -820 -690 -815 -670
rect -795 -690 -790 -670
rect -820 -720 -790 -690
rect -820 -740 -815 -720
rect -795 -740 -790 -720
rect -820 -770 -790 -740
rect -820 -790 -815 -770
rect -795 -790 -790 -770
rect -820 -820 -790 -790
rect -820 -840 -815 -820
rect -795 -840 -790 -820
rect -820 -870 -790 -840
rect -820 -890 -815 -870
rect -795 -890 -790 -870
rect -820 -920 -790 -890
rect -820 -940 -815 -920
rect -795 -940 -790 -920
rect -820 -970 -790 -940
rect -820 -990 -815 -970
rect -795 -990 -790 -970
rect -820 -1020 -790 -990
rect -820 -1040 -815 -1020
rect -795 -1040 -790 -1020
rect -820 -1050 -790 -1040
rect -720 -370 -690 -360
rect -720 -390 -715 -370
rect -695 -390 -690 -370
rect -720 -420 -690 -390
rect -720 -440 -715 -420
rect -695 -440 -690 -420
rect -720 -470 -690 -440
rect -720 -490 -715 -470
rect -695 -490 -690 -470
rect -720 -520 -690 -490
rect -720 -540 -715 -520
rect -695 -540 -690 -520
rect -720 -570 -690 -540
rect -720 -590 -715 -570
rect -695 -590 -690 -570
rect -720 -620 -690 -590
rect -720 -640 -715 -620
rect -695 -640 -690 -620
rect -720 -670 -690 -640
rect -720 -690 -715 -670
rect -695 -690 -690 -670
rect -720 -720 -690 -690
rect -720 -740 -715 -720
rect -695 -740 -690 -720
rect -720 -770 -690 -740
rect -720 -790 -715 -770
rect -695 -790 -690 -770
rect -720 -820 -690 -790
rect -720 -840 -715 -820
rect -695 -840 -690 -820
rect -720 -870 -690 -840
rect -720 -890 -715 -870
rect -695 -890 -690 -870
rect -720 -920 -690 -890
rect -720 -940 -715 -920
rect -695 -940 -690 -920
rect -720 -970 -690 -940
rect -720 -990 -715 -970
rect -695 -990 -690 -970
rect -720 -1020 -690 -990
rect -720 -1040 -715 -1020
rect -695 -1040 -690 -1020
rect -720 -1050 -690 -1040
rect -620 -370 -590 -360
rect -620 -390 -615 -370
rect -595 -390 -590 -370
rect -620 -420 -590 -390
rect -620 -440 -615 -420
rect -595 -440 -590 -420
rect -620 -470 -590 -440
rect -620 -490 -615 -470
rect -595 -490 -590 -470
rect -620 -520 -590 -490
rect -620 -540 -615 -520
rect -595 -540 -590 -520
rect -620 -570 -590 -540
rect -620 -590 -615 -570
rect -595 -590 -590 -570
rect -620 -620 -590 -590
rect -620 -640 -615 -620
rect -595 -640 -590 -620
rect -620 -670 -590 -640
rect -620 -690 -615 -670
rect -595 -690 -590 -670
rect -620 -720 -590 -690
rect -620 -740 -615 -720
rect -595 -740 -590 -720
rect -620 -770 -590 -740
rect -620 -790 -615 -770
rect -595 -790 -590 -770
rect -620 -820 -590 -790
rect -620 -840 -615 -820
rect -595 -840 -590 -820
rect -620 -870 -590 -840
rect -620 -890 -615 -870
rect -595 -890 -590 -870
rect -620 -920 -590 -890
rect -620 -940 -615 -920
rect -595 -940 -590 -920
rect -620 -970 -590 -940
rect -620 -990 -615 -970
rect -595 -990 -590 -970
rect -620 -1020 -590 -990
rect -620 -1040 -615 -1020
rect -595 -1040 -590 -1020
rect -620 -1050 -590 -1040
rect -520 -370 -490 -360
rect -520 -390 -515 -370
rect -495 -390 -490 -370
rect -520 -420 -490 -390
rect -520 -440 -515 -420
rect -495 -440 -490 -420
rect -520 -470 -490 -440
rect -520 -490 -515 -470
rect -495 -490 -490 -470
rect -520 -520 -490 -490
rect -520 -540 -515 -520
rect -495 -540 -490 -520
rect -520 -570 -490 -540
rect -520 -590 -515 -570
rect -495 -590 -490 -570
rect -520 -620 -490 -590
rect -520 -640 -515 -620
rect -495 -640 -490 -620
rect -520 -670 -490 -640
rect -520 -690 -515 -670
rect -495 -690 -490 -670
rect -520 -720 -490 -690
rect -520 -740 -515 -720
rect -495 -740 -490 -720
rect -520 -770 -490 -740
rect -520 -790 -515 -770
rect -495 -790 -490 -770
rect -520 -820 -490 -790
rect -520 -840 -515 -820
rect -495 -840 -490 -820
rect -520 -870 -490 -840
rect -520 -890 -515 -870
rect -495 -890 -490 -870
rect -520 -920 -490 -890
rect -520 -940 -515 -920
rect -495 -940 -490 -920
rect -520 -970 -490 -940
rect -520 -990 -515 -970
rect -495 -990 -490 -970
rect -520 -1020 -490 -990
rect -520 -1040 -515 -1020
rect -495 -1040 -490 -1020
rect -520 -1050 -490 -1040
rect -420 -370 -350 -360
rect -420 -390 -415 -370
rect -395 -390 -375 -370
rect -355 -390 -350 -370
rect -420 -420 -350 -390
rect -420 -440 -415 -420
rect -395 -440 -375 -420
rect -355 -440 -350 -420
rect -420 -470 -350 -440
rect -420 -490 -415 -470
rect -395 -490 -375 -470
rect -355 -490 -350 -470
rect 2040 -370 2110 -360
rect 2040 -390 2045 -370
rect 2065 -390 2085 -370
rect 2105 -390 2110 -370
rect 2040 -420 2110 -390
rect 2040 -440 2045 -420
rect 2065 -440 2085 -420
rect 2105 -440 2110 -420
rect 2040 -470 2110 -440
rect -420 -520 -350 -490
rect 385 -485 425 -475
rect 385 -505 395 -485
rect 415 -505 425 -485
rect 385 -515 425 -505
rect 445 -485 475 -475
rect 445 -505 450 -485
rect 470 -505 475 -485
rect 445 -515 475 -505
rect 495 -485 535 -475
rect 495 -505 505 -485
rect 525 -505 535 -485
rect 495 -515 535 -505
rect 605 -485 645 -475
rect 605 -505 615 -485
rect 635 -505 645 -485
rect 605 -515 645 -505
rect 715 -485 755 -475
rect 715 -505 725 -485
rect 745 -505 755 -485
rect 715 -515 755 -505
rect 825 -485 865 -475
rect 825 -505 835 -485
rect 855 -505 865 -485
rect 825 -515 865 -505
rect 935 -485 975 -475
rect 935 -505 945 -485
rect 965 -505 975 -485
rect 935 -515 975 -505
rect 1045 -485 1085 -475
rect 1045 -505 1055 -485
rect 1075 -505 1085 -485
rect 1045 -515 1085 -505
rect 1155 -485 1195 -475
rect 1155 -505 1165 -485
rect 1185 -505 1195 -485
rect 1155 -515 1195 -505
rect 1265 -485 1305 -475
rect 1265 -505 1275 -485
rect 1295 -505 1305 -485
rect 1265 -515 1305 -505
rect 1341 -485 1371 -475
rect 1341 -505 1346 -485
rect 1366 -505 1371 -485
rect 1341 -515 1371 -505
rect 1390 -485 1430 -475
rect 1390 -505 1400 -485
rect 1420 -505 1430 -485
rect 1390 -515 1430 -505
rect 2040 -490 2045 -470
rect 2065 -490 2085 -470
rect 2105 -490 2110 -470
rect -420 -540 -415 -520
rect -395 -540 -375 -520
rect -355 -540 -350 -520
rect 395 -540 415 -515
rect 505 -540 525 -515
rect 615 -540 635 -515
rect 725 -540 745 -515
rect 835 -540 855 -515
rect 945 -540 965 -515
rect 1055 -540 1075 -515
rect 1165 -540 1185 -515
rect 1275 -540 1295 -515
rect 1390 -540 1410 -515
rect 2040 -520 2110 -490
rect 2040 -540 2045 -520
rect 2065 -540 2085 -520
rect 2105 -540 2110 -520
rect -420 -570 -350 -540
rect -420 -590 -415 -570
rect -395 -590 -375 -570
rect -355 -590 -350 -570
rect -420 -620 -350 -590
rect -420 -640 -415 -620
rect -395 -640 -375 -620
rect -355 -640 -350 -620
rect -420 -670 -350 -640
rect -420 -690 -415 -670
rect -395 -690 -375 -670
rect -355 -690 -350 -670
rect -420 -720 -350 -690
rect -420 -740 -415 -720
rect -395 -740 -375 -720
rect -355 -740 -350 -720
rect -420 -770 -350 -740
rect -420 -790 -415 -770
rect -395 -790 -375 -770
rect -355 -790 -350 -770
rect 240 -550 310 -540
rect 240 -570 245 -550
rect 265 -570 285 -550
rect 305 -570 310 -550
rect 240 -600 310 -570
rect 240 -620 245 -600
rect 265 -620 285 -600
rect 305 -620 310 -600
rect 240 -650 310 -620
rect 240 -670 245 -650
rect 265 -670 285 -650
rect 305 -670 310 -650
rect 240 -700 310 -670
rect 240 -720 245 -700
rect 265 -720 285 -700
rect 305 -720 310 -700
rect 240 -750 310 -720
rect 240 -770 245 -750
rect 265 -770 285 -750
rect 305 -770 310 -750
rect 240 -780 310 -770
rect 335 -550 365 -540
rect 335 -570 340 -550
rect 360 -570 365 -550
rect 335 -600 365 -570
rect 335 -620 340 -600
rect 360 -620 365 -600
rect 335 -650 365 -620
rect 335 -670 340 -650
rect 360 -670 365 -650
rect 335 -700 365 -670
rect 335 -720 340 -700
rect 360 -720 365 -700
rect 335 -750 365 -720
rect 335 -770 340 -750
rect 360 -770 365 -750
rect 335 -780 365 -770
rect 390 -550 420 -540
rect 390 -570 395 -550
rect 415 -570 420 -550
rect 390 -600 420 -570
rect 390 -620 395 -600
rect 415 -620 420 -600
rect 390 -650 420 -620
rect 390 -670 395 -650
rect 415 -670 420 -650
rect 390 -700 420 -670
rect 390 -720 395 -700
rect 415 -720 420 -700
rect 390 -750 420 -720
rect 390 -770 395 -750
rect 415 -770 420 -750
rect 390 -780 420 -770
rect 445 -550 475 -540
rect 445 -570 450 -550
rect 470 -570 475 -550
rect 445 -600 475 -570
rect 445 -620 450 -600
rect 470 -620 475 -600
rect 445 -650 475 -620
rect 445 -670 450 -650
rect 470 -670 475 -650
rect 445 -700 475 -670
rect 445 -720 450 -700
rect 470 -720 475 -700
rect 445 -750 475 -720
rect 445 -770 450 -750
rect 470 -770 475 -750
rect 445 -780 475 -770
rect 500 -550 530 -540
rect 500 -570 505 -550
rect 525 -570 530 -550
rect 500 -600 530 -570
rect 500 -620 505 -600
rect 525 -620 530 -600
rect 500 -650 530 -620
rect 500 -670 505 -650
rect 525 -670 530 -650
rect 500 -700 530 -670
rect 500 -720 505 -700
rect 525 -720 530 -700
rect 500 -750 530 -720
rect 500 -770 505 -750
rect 525 -770 530 -750
rect 500 -780 530 -770
rect 555 -550 585 -540
rect 555 -570 560 -550
rect 580 -570 585 -550
rect 555 -600 585 -570
rect 555 -620 560 -600
rect 580 -620 585 -600
rect 555 -650 585 -620
rect 555 -670 560 -650
rect 580 -670 585 -650
rect 555 -700 585 -670
rect 555 -720 560 -700
rect 580 -720 585 -700
rect 555 -750 585 -720
rect 555 -770 560 -750
rect 580 -770 585 -750
rect 555 -780 585 -770
rect 610 -550 640 -540
rect 610 -570 615 -550
rect 635 -570 640 -550
rect 610 -600 640 -570
rect 610 -620 615 -600
rect 635 -620 640 -600
rect 610 -650 640 -620
rect 610 -670 615 -650
rect 635 -670 640 -650
rect 610 -700 640 -670
rect 610 -720 615 -700
rect 635 -720 640 -700
rect 610 -750 640 -720
rect 610 -770 615 -750
rect 635 -770 640 -750
rect 610 -780 640 -770
rect 665 -550 695 -540
rect 665 -570 670 -550
rect 690 -570 695 -550
rect 665 -600 695 -570
rect 665 -620 670 -600
rect 690 -620 695 -600
rect 665 -650 695 -620
rect 665 -670 670 -650
rect 690 -670 695 -650
rect 665 -700 695 -670
rect 665 -720 670 -700
rect 690 -720 695 -700
rect 665 -750 695 -720
rect 665 -770 670 -750
rect 690 -770 695 -750
rect 665 -780 695 -770
rect 720 -550 750 -540
rect 720 -570 725 -550
rect 745 -570 750 -550
rect 720 -600 750 -570
rect 720 -620 725 -600
rect 745 -620 750 -600
rect 720 -650 750 -620
rect 720 -670 725 -650
rect 745 -670 750 -650
rect 720 -700 750 -670
rect 720 -720 725 -700
rect 745 -720 750 -700
rect 720 -750 750 -720
rect 720 -770 725 -750
rect 745 -770 750 -750
rect 720 -780 750 -770
rect 775 -550 805 -540
rect 775 -570 780 -550
rect 800 -570 805 -550
rect 775 -600 805 -570
rect 775 -620 780 -600
rect 800 -620 805 -600
rect 775 -650 805 -620
rect 775 -670 780 -650
rect 800 -670 805 -650
rect 775 -700 805 -670
rect 775 -720 780 -700
rect 800 -720 805 -700
rect 775 -750 805 -720
rect 775 -770 780 -750
rect 800 -770 805 -750
rect 775 -780 805 -770
rect 830 -550 860 -540
rect 830 -570 835 -550
rect 855 -570 860 -550
rect 830 -600 860 -570
rect 830 -620 835 -600
rect 855 -620 860 -600
rect 830 -650 860 -620
rect 830 -670 835 -650
rect 855 -670 860 -650
rect 830 -700 860 -670
rect 830 -720 835 -700
rect 855 -720 860 -700
rect 830 -750 860 -720
rect 830 -770 835 -750
rect 855 -770 860 -750
rect 830 -780 860 -770
rect 885 -550 915 -540
rect 885 -570 890 -550
rect 910 -570 915 -550
rect 885 -600 915 -570
rect 885 -620 890 -600
rect 910 -620 915 -600
rect 885 -650 915 -620
rect 885 -670 890 -650
rect 910 -670 915 -650
rect 885 -700 915 -670
rect 885 -720 890 -700
rect 910 -720 915 -700
rect 885 -750 915 -720
rect 885 -770 890 -750
rect 910 -770 915 -750
rect 885 -780 915 -770
rect 940 -550 970 -540
rect 940 -570 945 -550
rect 965 -570 970 -550
rect 940 -600 970 -570
rect 940 -620 945 -600
rect 965 -620 970 -600
rect 940 -650 970 -620
rect 940 -670 945 -650
rect 965 -670 970 -650
rect 940 -700 970 -670
rect 940 -720 945 -700
rect 965 -720 970 -700
rect 940 -750 970 -720
rect 940 -770 945 -750
rect 965 -770 970 -750
rect 940 -780 970 -770
rect 995 -550 1025 -540
rect 995 -570 1000 -550
rect 1020 -570 1025 -550
rect 995 -600 1025 -570
rect 995 -620 1000 -600
rect 1020 -620 1025 -600
rect 995 -650 1025 -620
rect 995 -670 1000 -650
rect 1020 -670 1025 -650
rect 995 -700 1025 -670
rect 995 -720 1000 -700
rect 1020 -720 1025 -700
rect 995 -750 1025 -720
rect 995 -770 1000 -750
rect 1020 -770 1025 -750
rect 995 -780 1025 -770
rect 1050 -550 1080 -540
rect 1050 -570 1055 -550
rect 1075 -570 1080 -550
rect 1050 -600 1080 -570
rect 1050 -620 1055 -600
rect 1075 -620 1080 -600
rect 1050 -650 1080 -620
rect 1050 -670 1055 -650
rect 1075 -670 1080 -650
rect 1050 -700 1080 -670
rect 1050 -720 1055 -700
rect 1075 -720 1080 -700
rect 1050 -750 1080 -720
rect 1050 -770 1055 -750
rect 1075 -770 1080 -750
rect 1050 -780 1080 -770
rect 1105 -550 1135 -540
rect 1105 -570 1110 -550
rect 1130 -570 1135 -550
rect 1105 -600 1135 -570
rect 1105 -620 1110 -600
rect 1130 -620 1135 -600
rect 1105 -650 1135 -620
rect 1105 -670 1110 -650
rect 1130 -670 1135 -650
rect 1105 -700 1135 -670
rect 1105 -720 1110 -700
rect 1130 -720 1135 -700
rect 1105 -750 1135 -720
rect 1105 -770 1110 -750
rect 1130 -770 1135 -750
rect 1105 -780 1135 -770
rect 1160 -550 1190 -540
rect 1160 -570 1165 -550
rect 1185 -570 1190 -550
rect 1160 -600 1190 -570
rect 1160 -620 1165 -600
rect 1185 -620 1190 -600
rect 1160 -650 1190 -620
rect 1160 -670 1165 -650
rect 1185 -670 1190 -650
rect 1160 -700 1190 -670
rect 1160 -720 1165 -700
rect 1185 -720 1190 -700
rect 1160 -750 1190 -720
rect 1160 -770 1165 -750
rect 1185 -770 1190 -750
rect 1160 -780 1190 -770
rect 1215 -550 1245 -540
rect 1215 -570 1220 -550
rect 1240 -570 1245 -550
rect 1215 -600 1245 -570
rect 1215 -620 1220 -600
rect 1240 -620 1245 -600
rect 1215 -650 1245 -620
rect 1215 -670 1220 -650
rect 1240 -670 1245 -650
rect 1215 -700 1245 -670
rect 1215 -720 1220 -700
rect 1240 -720 1245 -700
rect 1215 -750 1245 -720
rect 1215 -770 1220 -750
rect 1240 -770 1245 -750
rect 1215 -780 1245 -770
rect 1270 -550 1300 -540
rect 1270 -570 1275 -550
rect 1295 -570 1300 -550
rect 1270 -600 1300 -570
rect 1270 -620 1275 -600
rect 1295 -620 1300 -600
rect 1270 -650 1300 -620
rect 1270 -670 1275 -650
rect 1295 -670 1300 -650
rect 1270 -700 1300 -670
rect 1270 -720 1275 -700
rect 1295 -720 1300 -700
rect 1270 -750 1300 -720
rect 1270 -770 1275 -750
rect 1295 -770 1300 -750
rect 1270 -780 1300 -770
rect 1325 -550 1355 -540
rect 1325 -570 1330 -550
rect 1350 -570 1355 -550
rect 1325 -600 1355 -570
rect 1325 -620 1330 -600
rect 1350 -620 1355 -600
rect 1325 -650 1355 -620
rect 1325 -670 1330 -650
rect 1350 -670 1355 -650
rect 1325 -700 1355 -670
rect 1325 -720 1330 -700
rect 1350 -720 1355 -700
rect 1325 -750 1355 -720
rect 1325 -770 1330 -750
rect 1350 -770 1355 -750
rect 1325 -780 1355 -770
rect 1380 -550 1410 -540
rect 1380 -570 1385 -550
rect 1405 -570 1410 -550
rect 1380 -600 1410 -570
rect 1380 -620 1385 -600
rect 1405 -620 1410 -600
rect 1380 -650 1410 -620
rect 1380 -670 1385 -650
rect 1405 -670 1410 -650
rect 1380 -700 1410 -670
rect 1380 -720 1385 -700
rect 1405 -720 1410 -700
rect 1380 -750 1410 -720
rect 1380 -770 1385 -750
rect 1405 -770 1410 -750
rect 1380 -780 1410 -770
rect 1435 -550 1505 -540
rect 1435 -570 1440 -550
rect 1460 -570 1480 -550
rect 1500 -570 1505 -550
rect 1435 -600 1505 -570
rect 1435 -620 1440 -600
rect 1460 -620 1480 -600
rect 1500 -620 1505 -600
rect 1435 -650 1505 -620
rect 1435 -670 1440 -650
rect 1460 -670 1480 -650
rect 1500 -670 1505 -650
rect 1435 -700 1505 -670
rect 1435 -720 1440 -700
rect 1460 -720 1480 -700
rect 1500 -720 1505 -700
rect 1435 -750 1505 -720
rect 1435 -770 1440 -750
rect 1460 -770 1480 -750
rect 1500 -770 1505 -750
rect 1435 -780 1505 -770
rect 2040 -570 2110 -540
rect 2040 -590 2045 -570
rect 2065 -590 2085 -570
rect 2105 -590 2110 -570
rect 2040 -620 2110 -590
rect 2040 -640 2045 -620
rect 2065 -640 2085 -620
rect 2105 -640 2110 -620
rect 2040 -670 2110 -640
rect 2040 -690 2045 -670
rect 2065 -690 2085 -670
rect 2105 -690 2110 -670
rect 2040 -720 2110 -690
rect 2040 -740 2045 -720
rect 2065 -740 2085 -720
rect 2105 -740 2110 -720
rect 2040 -770 2110 -740
rect -420 -820 -350 -790
rect 285 -800 305 -780
rect 340 -800 360 -780
rect 450 -800 470 -780
rect 560 -800 580 -780
rect 670 -800 690 -780
rect 780 -800 800 -780
rect 890 -800 910 -780
rect 1000 -800 1020 -780
rect 1110 -800 1130 -780
rect 1220 -800 1240 -780
rect 1330 -800 1350 -780
rect 1440 -800 1460 -780
rect 2040 -790 2045 -770
rect 2065 -790 2085 -770
rect 2105 -790 2110 -770
rect -420 -840 -415 -820
rect -395 -840 -375 -820
rect -355 -840 -350 -820
rect 265 -810 305 -800
rect 265 -830 275 -810
rect 295 -830 305 -810
rect 265 -840 305 -830
rect 330 -810 370 -800
rect 330 -830 340 -810
rect 360 -830 370 -810
rect 330 -840 370 -830
rect 440 -810 480 -800
rect 440 -830 450 -810
rect 470 -830 480 -810
rect 440 -840 480 -830
rect 550 -810 590 -800
rect 550 -830 560 -810
rect 580 -830 590 -810
rect 550 -840 590 -830
rect 660 -810 700 -800
rect 660 -830 670 -810
rect 690 -830 700 -810
rect 660 -840 700 -830
rect 770 -810 810 -800
rect 770 -830 780 -810
rect 800 -830 810 -810
rect 770 -840 810 -830
rect 880 -810 920 -800
rect 880 -830 890 -810
rect 910 -830 920 -810
rect 880 -840 920 -830
rect 990 -810 1030 -800
rect 990 -830 1000 -810
rect 1020 -830 1030 -810
rect 990 -840 1030 -830
rect 1100 -810 1140 -800
rect 1100 -830 1110 -810
rect 1130 -830 1140 -810
rect 1100 -840 1140 -830
rect 1210 -810 1250 -800
rect 1210 -830 1220 -810
rect 1240 -830 1250 -810
rect 1210 -840 1250 -830
rect 1320 -810 1360 -800
rect 1320 -830 1330 -810
rect 1350 -830 1360 -810
rect 1320 -840 1360 -830
rect 1430 -810 1470 -800
rect 1430 -830 1440 -810
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 2040 -820 2110 -790
rect 2040 -840 2045 -820
rect 2065 -840 2085 -820
rect 2105 -840 2110 -820
rect -420 -870 -350 -840
rect -420 -890 -415 -870
rect -395 -890 -375 -870
rect -355 -890 -350 -870
rect -420 -920 -350 -890
rect 1315 -870 1355 -860
rect 1315 -890 1325 -870
rect 1345 -890 1355 -870
rect -420 -940 -415 -920
rect -395 -940 -375 -920
rect -355 -940 -350 -920
rect 550 -905 590 -895
rect 550 -925 560 -905
rect 580 -925 590 -905
rect 550 -935 590 -925
rect 660 -905 700 -895
rect 660 -925 670 -905
rect 690 -925 700 -905
rect 660 -935 700 -925
rect 770 -905 810 -895
rect 770 -925 780 -905
rect 800 -925 810 -905
rect 770 -935 810 -925
rect 1005 -905 1045 -895
rect 1005 -925 1015 -905
rect 1035 -925 1045 -905
rect 1005 -935 1045 -925
rect 1125 -905 1165 -895
rect 1125 -925 1135 -905
rect 1155 -925 1165 -905
rect 1125 -935 1165 -925
rect 1255 -905 1295 -895
rect 1255 -925 1265 -905
rect 1285 -925 1295 -905
rect 1255 -935 1295 -925
rect 1315 -900 1355 -890
rect 2040 -870 2110 -840
rect 2040 -890 2045 -870
rect 2065 -890 2085 -870
rect 2105 -890 2110 -870
rect -420 -970 -350 -940
rect 560 -955 580 -935
rect 670 -955 690 -935
rect 780 -955 800 -935
rect 1315 -955 1335 -900
rect -420 -990 -415 -970
rect -395 -990 -375 -970
rect -355 -990 -350 -970
rect -420 -1020 -350 -990
rect -420 -1040 -415 -1020
rect -395 -1040 -375 -1020
rect -355 -1040 -350 -1020
rect -420 -1050 -350 -1040
rect 460 -965 530 -955
rect 460 -985 465 -965
rect 485 -985 505 -965
rect 525 -985 530 -965
rect 460 -1015 530 -985
rect 460 -1035 465 -1015
rect 485 -1035 505 -1015
rect 525 -1035 530 -1015
rect -1015 -1070 -995 -1050
rect -815 -1070 -795 -1050
rect -615 -1070 -595 -1050
rect -415 -1070 -395 -1050
rect 460 -1065 530 -1035
rect -1025 -1080 -985 -1070
rect -1025 -1100 -1015 -1080
rect -995 -1100 -985 -1080
rect -1025 -1110 -985 -1100
rect -825 -1080 -785 -1070
rect -825 -1100 -815 -1080
rect -795 -1100 -785 -1080
rect -825 -1110 -785 -1100
rect -625 -1080 -585 -1070
rect -625 -1100 -615 -1080
rect -595 -1100 -585 -1080
rect -625 -1110 -585 -1100
rect -425 -1080 -385 -1070
rect -425 -1100 -415 -1080
rect -395 -1100 -385 -1080
rect 460 -1085 465 -1065
rect 485 -1085 505 -1065
rect 525 -1085 530 -1065
rect 460 -1095 530 -1085
rect 555 -965 585 -955
rect 555 -985 560 -965
rect 580 -985 585 -965
rect 555 -1015 585 -985
rect 555 -1035 560 -1015
rect 580 -1035 585 -1015
rect 555 -1065 585 -1035
rect 555 -1085 560 -1065
rect 580 -1085 585 -1065
rect 555 -1095 585 -1085
rect 610 -965 640 -955
rect 610 -985 615 -965
rect 635 -985 640 -965
rect 610 -1015 640 -985
rect 610 -1035 615 -1015
rect 635 -1035 640 -1015
rect 610 -1065 640 -1035
rect 610 -1085 615 -1065
rect 635 -1085 640 -1065
rect 610 -1095 640 -1085
rect 665 -965 695 -955
rect 665 -985 670 -965
rect 690 -985 695 -965
rect 665 -1015 695 -985
rect 665 -1035 670 -1015
rect 690 -1035 695 -1015
rect 665 -1065 695 -1035
rect 665 -1085 670 -1065
rect 690 -1085 695 -1065
rect 665 -1095 695 -1085
rect 720 -965 750 -955
rect 720 -985 725 -965
rect 745 -985 750 -965
rect 720 -1015 750 -985
rect 720 -1035 725 -1015
rect 745 -1035 750 -1015
rect 720 -1065 750 -1035
rect 720 -1085 725 -1065
rect 745 -1085 750 -1065
rect 720 -1095 750 -1085
rect 775 -965 805 -955
rect 775 -985 780 -965
rect 800 -985 805 -965
rect 775 -1015 805 -985
rect 775 -1035 780 -1015
rect 800 -1035 805 -1015
rect 775 -1065 805 -1035
rect 775 -1085 780 -1065
rect 800 -1085 805 -1065
rect 775 -1095 805 -1085
rect 830 -965 900 -955
rect 830 -985 835 -965
rect 855 -985 875 -965
rect 895 -985 900 -965
rect 830 -1015 900 -985
rect 965 -965 995 -955
rect 965 -985 970 -965
rect 990 -985 995 -965
rect 965 -1005 995 -985
rect 830 -1035 835 -1015
rect 855 -1035 875 -1015
rect 895 -1035 900 -1015
rect 830 -1065 900 -1035
rect 925 -1015 995 -1005
rect 925 -1035 935 -1015
rect 955 -1035 970 -1015
rect 990 -1035 995 -1015
rect 925 -1045 995 -1035
rect 830 -1085 835 -1065
rect 855 -1085 875 -1065
rect 895 -1085 900 -1065
rect 830 -1095 900 -1085
rect 965 -1065 995 -1045
rect 965 -1085 970 -1065
rect 990 -1085 995 -1065
rect 965 -1095 995 -1085
rect 1305 -965 1335 -955
rect 1305 -985 1310 -965
rect 1330 -985 1335 -965
rect 1305 -1015 1335 -985
rect 1305 -1035 1310 -1015
rect 1330 -1035 1335 -1015
rect 1305 -1065 1335 -1035
rect 2040 -920 2110 -890
rect 2040 -940 2045 -920
rect 2065 -940 2085 -920
rect 2105 -940 2110 -920
rect 2040 -970 2110 -940
rect 2040 -990 2045 -970
rect 2065 -990 2085 -970
rect 2105 -990 2110 -970
rect 2040 -1020 2110 -990
rect 2040 -1040 2045 -1020
rect 2065 -1040 2085 -1020
rect 2105 -1040 2110 -1020
rect 2040 -1050 2110 -1040
rect 2180 -370 2210 -360
rect 2180 -390 2185 -370
rect 2205 -390 2210 -370
rect 2180 -420 2210 -390
rect 2180 -440 2185 -420
rect 2205 -440 2210 -420
rect 2180 -470 2210 -440
rect 2180 -490 2185 -470
rect 2205 -490 2210 -470
rect 2180 -520 2210 -490
rect 2180 -540 2185 -520
rect 2205 -540 2210 -520
rect 2180 -570 2210 -540
rect 2180 -590 2185 -570
rect 2205 -590 2210 -570
rect 2180 -620 2210 -590
rect 2180 -640 2185 -620
rect 2205 -640 2210 -620
rect 2180 -670 2210 -640
rect 2180 -690 2185 -670
rect 2205 -690 2210 -670
rect 2180 -720 2210 -690
rect 2180 -740 2185 -720
rect 2205 -740 2210 -720
rect 2180 -770 2210 -740
rect 2180 -790 2185 -770
rect 2205 -790 2210 -770
rect 2180 -820 2210 -790
rect 2180 -840 2185 -820
rect 2205 -840 2210 -820
rect 2180 -870 2210 -840
rect 2180 -890 2185 -870
rect 2205 -890 2210 -870
rect 2180 -920 2210 -890
rect 2180 -940 2185 -920
rect 2205 -940 2210 -920
rect 2180 -970 2210 -940
rect 2180 -990 2185 -970
rect 2205 -990 2210 -970
rect 2180 -1020 2210 -990
rect 2180 -1040 2185 -1020
rect 2205 -1040 2210 -1020
rect 2180 -1050 2210 -1040
rect 2280 -370 2310 -360
rect 2280 -390 2285 -370
rect 2305 -390 2310 -370
rect 2280 -420 2310 -390
rect 2280 -440 2285 -420
rect 2305 -440 2310 -420
rect 2280 -470 2310 -440
rect 2280 -490 2285 -470
rect 2305 -490 2310 -470
rect 2280 -520 2310 -490
rect 2280 -540 2285 -520
rect 2305 -540 2310 -520
rect 2280 -570 2310 -540
rect 2280 -590 2285 -570
rect 2305 -590 2310 -570
rect 2280 -620 2310 -590
rect 2280 -640 2285 -620
rect 2305 -640 2310 -620
rect 2280 -670 2310 -640
rect 2280 -690 2285 -670
rect 2305 -690 2310 -670
rect 2280 -720 2310 -690
rect 2280 -740 2285 -720
rect 2305 -740 2310 -720
rect 2280 -770 2310 -740
rect 2280 -790 2285 -770
rect 2305 -790 2310 -770
rect 2280 -820 2310 -790
rect 2280 -840 2285 -820
rect 2305 -840 2310 -820
rect 2280 -870 2310 -840
rect 2280 -890 2285 -870
rect 2305 -890 2310 -870
rect 2280 -920 2310 -890
rect 2280 -940 2285 -920
rect 2305 -940 2310 -920
rect 2280 -970 2310 -940
rect 2280 -990 2285 -970
rect 2305 -990 2310 -970
rect 2280 -1020 2310 -990
rect 2280 -1040 2285 -1020
rect 2305 -1040 2310 -1020
rect 2280 -1050 2310 -1040
rect 2380 -370 2410 -360
rect 2380 -390 2385 -370
rect 2405 -390 2410 -370
rect 2380 -420 2410 -390
rect 2380 -440 2385 -420
rect 2405 -440 2410 -420
rect 2380 -470 2410 -440
rect 2380 -490 2385 -470
rect 2405 -490 2410 -470
rect 2380 -520 2410 -490
rect 2380 -540 2385 -520
rect 2405 -540 2410 -520
rect 2380 -570 2410 -540
rect 2380 -590 2385 -570
rect 2405 -590 2410 -570
rect 2380 -620 2410 -590
rect 2380 -640 2385 -620
rect 2405 -640 2410 -620
rect 2380 -670 2410 -640
rect 2380 -690 2385 -670
rect 2405 -690 2410 -670
rect 2380 -720 2410 -690
rect 2380 -740 2385 -720
rect 2405 -740 2410 -720
rect 2380 -770 2410 -740
rect 2380 -790 2385 -770
rect 2405 -790 2410 -770
rect 2380 -820 2410 -790
rect 2380 -840 2385 -820
rect 2405 -840 2410 -820
rect 2380 -870 2410 -840
rect 2380 -890 2385 -870
rect 2405 -890 2410 -870
rect 2380 -920 2410 -890
rect 2380 -940 2385 -920
rect 2405 -940 2410 -920
rect 2380 -970 2410 -940
rect 2380 -990 2385 -970
rect 2405 -990 2410 -970
rect 2380 -1020 2410 -990
rect 2380 -1040 2385 -1020
rect 2405 -1040 2410 -1020
rect 2380 -1050 2410 -1040
rect 2480 -370 2510 -360
rect 2480 -390 2485 -370
rect 2505 -390 2510 -370
rect 2480 -420 2510 -390
rect 2480 -440 2485 -420
rect 2505 -440 2510 -420
rect 2480 -470 2510 -440
rect 2480 -490 2485 -470
rect 2505 -490 2510 -470
rect 2480 -520 2510 -490
rect 2480 -540 2485 -520
rect 2505 -540 2510 -520
rect 2480 -570 2510 -540
rect 2480 -590 2485 -570
rect 2505 -590 2510 -570
rect 2480 -620 2510 -590
rect 2480 -640 2485 -620
rect 2505 -640 2510 -620
rect 2480 -670 2510 -640
rect 2480 -690 2485 -670
rect 2505 -690 2510 -670
rect 2480 -720 2510 -690
rect 2480 -740 2485 -720
rect 2505 -740 2510 -720
rect 2480 -770 2510 -740
rect 2480 -790 2485 -770
rect 2505 -790 2510 -770
rect 2480 -820 2510 -790
rect 2480 -840 2485 -820
rect 2505 -840 2510 -820
rect 2480 -870 2510 -840
rect 2480 -890 2485 -870
rect 2505 -890 2510 -870
rect 2480 -920 2510 -890
rect 2480 -940 2485 -920
rect 2505 -940 2510 -920
rect 2480 -970 2510 -940
rect 2480 -990 2485 -970
rect 2505 -990 2510 -970
rect 2480 -1020 2510 -990
rect 2480 -1040 2485 -1020
rect 2505 -1040 2510 -1020
rect 2480 -1050 2510 -1040
rect 2580 -370 2610 -360
rect 2580 -390 2585 -370
rect 2605 -390 2610 -370
rect 2580 -420 2610 -390
rect 2580 -440 2585 -420
rect 2605 -440 2610 -420
rect 2580 -470 2610 -440
rect 2580 -490 2585 -470
rect 2605 -490 2610 -470
rect 2580 -520 2610 -490
rect 2580 -540 2585 -520
rect 2605 -540 2610 -520
rect 2580 -570 2610 -540
rect 2580 -590 2585 -570
rect 2605 -590 2610 -570
rect 2580 -620 2610 -590
rect 2580 -640 2585 -620
rect 2605 -640 2610 -620
rect 2580 -670 2610 -640
rect 2580 -690 2585 -670
rect 2605 -690 2610 -670
rect 2580 -720 2610 -690
rect 2580 -740 2585 -720
rect 2605 -740 2610 -720
rect 2580 -770 2610 -740
rect 2580 -790 2585 -770
rect 2605 -790 2610 -770
rect 2580 -820 2610 -790
rect 2580 -840 2585 -820
rect 2605 -840 2610 -820
rect 2580 -870 2610 -840
rect 2580 -890 2585 -870
rect 2605 -890 2610 -870
rect 2580 -920 2610 -890
rect 2580 -940 2585 -920
rect 2605 -940 2610 -920
rect 2580 -970 2610 -940
rect 2580 -990 2585 -970
rect 2605 -990 2610 -970
rect 2580 -1020 2610 -990
rect 2580 -1040 2585 -1020
rect 2605 -1040 2610 -1020
rect 2580 -1050 2610 -1040
rect 2680 -370 2750 -360
rect 2680 -390 2685 -370
rect 2705 -390 2725 -370
rect 2745 -390 2750 -370
rect 2680 -420 2750 -390
rect 2680 -440 2685 -420
rect 2705 -440 2725 -420
rect 2745 -440 2750 -420
rect 2680 -470 2750 -440
rect 2680 -490 2685 -470
rect 2705 -490 2725 -470
rect 2745 -490 2750 -470
rect 2680 -520 2750 -490
rect 2680 -540 2685 -520
rect 2705 -540 2725 -520
rect 2745 -540 2750 -520
rect 2680 -570 2750 -540
rect 2680 -590 2685 -570
rect 2705 -590 2725 -570
rect 2745 -590 2750 -570
rect 2680 -620 2750 -590
rect 2680 -640 2685 -620
rect 2705 -640 2725 -620
rect 2745 -640 2750 -620
rect 2805 -387 2840 -380
rect 2805 -407 2810 -387
rect 2835 -407 2840 -387
rect 2805 -415 2840 -407
rect 2865 -387 2900 -380
rect 2865 -407 2870 -387
rect 2895 -407 2900 -387
rect 2865 -415 2900 -407
rect 2680 -670 2750 -640
rect 2680 -690 2685 -670
rect 2705 -690 2725 -670
rect 2745 -690 2750 -670
rect 2680 -720 2750 -690
rect 2680 -740 2685 -720
rect 2705 -740 2725 -720
rect 2745 -740 2750 -720
rect 2680 -770 2750 -740
rect 2680 -790 2685 -770
rect 2705 -790 2725 -770
rect 2745 -790 2750 -770
rect 2680 -820 2750 -790
rect 2680 -840 2685 -820
rect 2705 -840 2725 -820
rect 2745 -840 2750 -820
rect 2680 -870 2750 -840
rect 2680 -890 2685 -870
rect 2705 -890 2725 -870
rect 2745 -890 2750 -870
rect 2680 -920 2750 -890
rect 2680 -940 2685 -920
rect 2705 -940 2725 -920
rect 2745 -940 2750 -920
rect 2680 -970 2750 -940
rect 2680 -990 2685 -970
rect 2705 -990 2725 -970
rect 2745 -990 2750 -970
rect 2680 -1020 2750 -990
rect 2680 -1040 2685 -1020
rect 2705 -1040 2725 -1020
rect 2745 -1040 2750 -1020
rect 2680 -1050 2750 -1040
rect 1305 -1085 1310 -1065
rect 1330 -1085 1335 -1065
rect 2085 -1070 2105 -1050
rect 2285 -1070 2305 -1050
rect 2485 -1070 2505 -1050
rect 2685 -1070 2705 -1050
rect 1305 -1095 1335 -1085
rect 2075 -1080 2115 -1070
rect -425 -1110 -385 -1100
rect 500 -1125 530 -1095
rect 615 -1115 635 -1095
rect 725 -1115 745 -1095
rect 500 -1145 505 -1125
rect 525 -1145 530 -1125
rect 500 -1155 530 -1145
rect 605 -1125 645 -1115
rect 605 -1145 615 -1125
rect 635 -1145 645 -1125
rect 605 -1155 645 -1145
rect 715 -1125 755 -1115
rect 715 -1145 725 -1125
rect 745 -1145 755 -1125
rect 715 -1155 755 -1145
rect 830 -1125 860 -1095
rect 2075 -1100 2085 -1080
rect 2105 -1100 2115 -1080
rect 2075 -1110 2115 -1100
rect 2275 -1080 2315 -1070
rect 2275 -1100 2285 -1080
rect 2305 -1100 2315 -1080
rect 2275 -1110 2315 -1100
rect 2475 -1080 2515 -1070
rect 2475 -1100 2485 -1080
rect 2505 -1100 2515 -1080
rect 2475 -1110 2515 -1100
rect 2675 -1080 2715 -1070
rect 2675 -1100 2685 -1080
rect 2705 -1100 2715 -1080
rect 2675 -1110 2715 -1100
rect 2840 -1105 2865 -1055
rect 830 -1145 835 -1125
rect 855 -1145 860 -1125
rect 830 -1155 860 -1145
<< viali >>
rect 40 2700 60 2720
rect 160 2700 180 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1040 2700 1060 2720
rect 1100 2700 1120 2720
rect 1160 2700 1180 2720
rect 1448 2700 1468 2720
rect 1508 2700 1528 2720
rect 1628 2700 1648 2720
rect 510 2530 530 2550
rect 570 2530 590 2550
rect 630 2530 650 2550
rect 690 2530 710 2550
rect 85 2280 105 2300
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1524 2280 1544 2300
rect 1583 2280 1603 2300
rect -1155 2125 -1135 2145
rect -1035 2125 -1015 2145
rect -915 2125 -895 2145
rect -795 2125 -775 2145
rect -675 2125 -655 2145
rect -555 2125 -535 2145
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 90 2125 110 2145
rect 210 2125 230 2145
rect 330 2125 350 2145
rect 450 2125 470 2145
rect 570 2125 590 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1100 2125 1120 2145
rect 1220 2125 1240 2145
rect 1340 2125 1360 2145
rect 1460 2125 1480 2145
rect 1580 2125 1600 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect 2225 2125 2245 2145
rect 2345 2125 2365 2145
rect 2465 2125 2485 2145
rect 2585 2125 2605 2145
rect 2705 2125 2725 2145
rect 2825 2125 2845 2145
rect -1095 1700 -1075 1720
rect -975 1700 -955 1720
rect -855 1700 -835 1720
rect -795 1700 -775 1720
rect -735 1700 -715 1720
rect -615 1700 -595 1720
rect -495 1700 -475 1720
rect 30 1700 50 1720
rect 150 1700 170 1720
rect 270 1700 290 1720
rect 330 1700 350 1720
rect 390 1700 410 1720
rect 510 1700 530 1720
rect 630 1700 650 1720
rect 1040 1700 1060 1720
rect 1160 1700 1180 1720
rect 1280 1700 1300 1720
rect 1340 1700 1360 1720
rect 1400 1700 1420 1720
rect 1520 1700 1540 1720
rect 1640 1700 1660 1720
rect 2165 1700 2185 1720
rect 2285 1700 2305 1720
rect 2405 1700 2425 1720
rect 2465 1700 2485 1720
rect 2525 1700 2545 1720
rect 2645 1700 2665 1720
rect 2765 1700 2785 1720
rect 465 1555 485 1575
rect 630 1555 650 1575
rect 795 1555 815 1575
rect 875 1555 895 1575
rect 1040 1555 1060 1575
rect 1205 1555 1225 1575
rect -1125 1460 -1105 1480
rect -1015 1460 -995 1480
rect -905 1460 -885 1480
rect -795 1460 -775 1480
rect -685 1460 -665 1480
rect -575 1460 -555 1480
rect 575 1510 595 1530
rect 685 1510 705 1530
rect 985 1510 1005 1530
rect 1095 1510 1115 1530
rect -465 1460 -445 1480
rect -1495 1400 -1475 1420
rect -1440 1400 -1420 1420
rect -1385 1400 -1365 1420
rect 2135 1460 2155 1480
rect 2245 1460 2265 1480
rect 2355 1460 2375 1480
rect 2465 1460 2485 1480
rect 2575 1460 2595 1480
rect 2685 1460 2705 1480
rect 2795 1460 2815 1480
rect 510 1200 530 1220
rect 557 1190 577 1210
rect 630 1190 650 1210
rect 703 1190 723 1210
rect 750 1200 770 1220
rect 920 1200 940 1220
rect 967 1190 987 1210
rect 1040 1190 1060 1210
rect 1113 1190 1133 1210
rect 1160 1200 1180 1220
rect 555 1130 575 1150
rect 1115 1130 1135 1150
rect -40 880 -20 900
rect 70 880 90 900
rect 180 880 200 900
rect 235 880 255 900
rect 290 880 310 900
rect 400 880 420 900
rect 510 880 530 900
rect 805 900 825 920
rect 890 900 910 920
rect 1160 880 1180 900
rect 1270 880 1290 900
rect 1380 880 1400 900
rect 1435 880 1455 900
rect 1490 880 1510 900
rect 1600 880 1620 900
rect 1710 880 1730 900
rect -1495 795 -1475 815
rect -1440 795 -1420 815
rect -1385 795 -1365 815
rect -1070 785 -1050 805
rect -960 785 -940 805
rect -850 785 -830 805
rect -795 780 -775 800
rect -740 785 -720 805
rect -630 785 -610 805
rect -520 785 -500 805
rect -1135 645 -1115 665
rect -1070 645 -1050 665
rect -960 645 -940 665
rect -850 645 -830 665
rect -740 645 -720 665
rect -630 645 -610 665
rect -520 645 -500 665
rect -455 645 -435 665
rect -95 655 -75 675
rect 15 655 35 675
rect 125 655 145 675
rect 235 655 255 675
rect 345 655 365 675
rect 455 655 475 675
rect 565 655 585 675
rect 3055 1400 3075 1420
rect 3110 1400 3130 1420
rect 3165 1400 3185 1420
rect 2190 785 2210 805
rect 2300 785 2320 805
rect 2410 785 2430 805
rect 2465 780 2485 800
rect 2520 785 2540 805
rect 2630 785 2650 805
rect 2740 785 2760 805
rect 3055 795 3075 815
rect 3110 795 3130 815
rect 3165 795 3185 815
rect 1105 655 1125 675
rect 1215 655 1235 675
rect 1325 655 1345 675
rect 1435 655 1455 675
rect 1545 655 1565 675
rect 1655 655 1675 675
rect 1765 655 1785 675
rect 2125 645 2145 665
rect 2190 645 2210 665
rect 2300 645 2320 665
rect 2410 645 2430 665
rect 2520 645 2540 665
rect 2630 645 2650 665
rect 2740 645 2760 665
rect 2805 645 2825 665
rect 725 580 745 600
rect 835 580 855 600
rect 945 580 965 600
rect -40 530 -20 550
rect 70 530 90 550
rect 180 530 200 550
rect 290 530 310 550
rect 400 530 420 550
rect 510 530 530 550
rect 1160 530 1180 550
rect 1270 530 1290 550
rect 1380 530 1400 550
rect 1490 530 1510 550
rect 1600 530 1620 550
rect 1710 530 1730 550
rect 235 480 255 500
rect 725 480 745 500
rect 800 480 820 500
rect 870 480 890 500
rect 945 480 965 500
rect 1435 480 1455 500
rect -1015 370 -995 390
rect -905 370 -885 390
rect -795 370 -775 390
rect -740 370 -720 390
rect -685 370 -665 390
rect -575 370 -555 390
rect 2245 370 2265 390
rect 2355 370 2375 390
rect 2410 370 2430 390
rect 2465 370 2485 390
rect 2575 370 2595 390
rect 2685 370 2705 390
rect -1015 260 -995 280
rect -905 260 -885 280
rect -795 260 -775 280
rect -740 260 -720 280
rect -685 260 -665 280
rect -575 260 -555 280
rect -95 260 -75 280
rect 15 260 35 280
rect 125 260 145 280
rect 235 260 255 280
rect 345 260 365 280
rect 455 260 475 280
rect 605 260 625 280
rect 780 260 800 280
rect 835 260 855 280
rect 890 260 910 280
rect 1065 260 1085 280
rect 1215 260 1235 280
rect 1325 260 1345 280
rect 1435 260 1455 280
rect 1545 260 1565 280
rect 1655 260 1675 280
rect 1765 260 1785 280
rect 2245 260 2265 280
rect 2355 260 2375 280
rect 2410 260 2430 280
rect 2465 260 2485 280
rect 2575 260 2595 280
rect 2685 260 2705 280
rect -1485 -113 -1460 -93
rect -1425 -113 -1400 -93
rect -1365 -113 -1340 -93
rect 780 -15 800 5
rect 835 -10 855 10
rect 890 -15 910 5
rect -1305 -113 -1280 -93
rect -1135 -115 -1115 -95
rect -1070 -115 -1050 -95
rect -960 -115 -940 -95
rect -850 -115 -830 -95
rect -740 -115 -720 -95
rect -630 -115 -610 -95
rect -520 -115 -500 -95
rect -455 -115 -435 -95
rect 2125 -115 2145 -95
rect 2190 -115 2210 -95
rect 2300 -115 2320 -95
rect 2410 -115 2430 -95
rect 2520 -115 2540 -95
rect 2630 -115 2650 -95
rect 2740 -115 2760 -95
rect 2805 -115 2825 -95
rect 2970 -113 2995 -93
rect 3030 -113 3055 -93
rect 3090 -113 3115 -93
rect 3150 -113 3175 -93
rect -915 -325 -895 -305
rect -715 -325 -695 -305
rect -615 -325 -595 -305
rect -515 -325 -495 -305
rect 725 -335 745 -315
rect 835 -335 855 -315
rect 945 -335 965 -315
rect 2185 -325 2205 -305
rect 2285 -325 2305 -305
rect 2385 -325 2405 -305
rect 2585 -325 2605 -305
rect -1205 -407 -1180 -387
rect -1145 -407 -1120 -387
rect 395 -505 415 -485
rect 450 -505 470 -485
rect 505 -505 525 -485
rect 615 -505 635 -485
rect 725 -505 745 -485
rect 835 -505 855 -485
rect 945 -505 965 -485
rect 1055 -505 1075 -485
rect 1165 -505 1185 -485
rect 1275 -505 1295 -485
rect 1346 -505 1366 -485
rect 1400 -505 1420 -485
rect 275 -830 295 -810
rect 340 -830 360 -810
rect 450 -830 470 -810
rect 560 -830 580 -810
rect 670 -830 690 -810
rect 780 -830 800 -810
rect 890 -830 910 -810
rect 1000 -830 1020 -810
rect 1110 -830 1130 -810
rect 1220 -830 1240 -810
rect 1330 -830 1350 -810
rect 1440 -830 1460 -810
rect 1325 -890 1345 -870
rect 560 -925 580 -905
rect 670 -925 690 -905
rect 780 -925 800 -905
rect 1015 -925 1035 -905
rect 1135 -925 1155 -905
rect 1265 -925 1285 -905
rect -1015 -1100 -995 -1080
rect -815 -1100 -795 -1080
rect -615 -1100 -595 -1080
rect -415 -1100 -395 -1080
rect 935 -1035 955 -1015
rect 2810 -407 2835 -387
rect 2870 -407 2895 -387
rect 505 -1145 525 -1125
rect 615 -1145 635 -1125
rect 725 -1145 745 -1125
rect 2085 -1100 2105 -1080
rect 2285 -1100 2305 -1080
rect 2485 -1100 2505 -1080
rect 2685 -1100 2705 -1080
rect 835 -1145 855 -1125
<< metal1 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 150 2780 190 2785
rect 150 2750 155 2780
rect 185 2750 190 2780
rect 150 2745 190 2750
rect 620 2780 660 2785
rect 620 2750 625 2780
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 160 2730 180 2745
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2695 70 2725
rect 30 2690 70 2695
rect 150 2725 190 2730
rect 150 2695 155 2725
rect 185 2695 190 2725
rect 150 2690 190 2695
rect 210 2725 250 2730
rect 210 2695 215 2725
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 630 2560 650 2745
rect 835 2730 855 4240
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2750 1070 2780
rect 1030 2745 1070 2750
rect 1498 2780 1538 2785
rect 1498 2750 1503 2780
rect 1533 2750 1538 2780
rect 1498 2745 1538 2750
rect 1040 2730 1060 2745
rect 1508 2730 1528 2745
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2695 865 2725
rect 825 2690 865 2695
rect 970 2725 1010 2730
rect 970 2695 975 2725
rect 1005 2695 1010 2725
rect 970 2690 1010 2695
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 1035 2690 1065 2700
rect 1090 2725 1130 2730
rect 1090 2695 1095 2725
rect 1125 2695 1130 2725
rect 1090 2690 1130 2695
rect 1150 2725 1190 2730
rect 1150 2695 1155 2725
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1438 2725 1478 2730
rect 1438 2695 1443 2725
rect 1473 2695 1478 2725
rect 1438 2690 1478 2695
rect 1498 2725 1538 2730
rect 1498 2695 1503 2725
rect 1533 2695 1538 2725
rect 1498 2690 1538 2695
rect 1618 2725 1658 2730
rect 1618 2695 1623 2725
rect 1653 2695 1658 2725
rect 1618 2690 1658 2695
rect 835 2560 855 2690
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2525 540 2555
rect 500 2520 540 2525
rect 560 2555 600 2560
rect 560 2525 565 2555
rect 595 2525 600 2555
rect 560 2520 600 2525
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 625 2520 655 2530
rect 680 2555 720 2560
rect 680 2525 685 2555
rect 715 2525 720 2555
rect 680 2520 720 2525
rect 825 2555 865 2560
rect 825 2525 830 2555
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2275 115 2305
rect 75 2270 115 2275
rect 139 2305 169 2310
rect 139 2270 169 2275
rect 609 2305 639 2310
rect 609 2270 639 2275
rect 770 2305 810 2310
rect 770 2275 775 2305
rect 805 2275 810 2305
rect 770 2270 810 2275
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2175 -765 2205
rect -805 2170 -765 2175
rect -235 2205 -195 2210
rect -235 2175 -230 2205
rect -200 2175 -195 2205
rect -235 2170 -195 2175
rect -795 2155 -775 2170
rect -1165 2150 -1125 2155
rect -1165 2120 -1160 2150
rect -1130 2120 -1125 2150
rect -1165 2115 -1125 2120
rect -1045 2150 -1005 2155
rect -1045 2120 -1040 2150
rect -1010 2120 -1005 2150
rect -1045 2115 -1005 2120
rect -925 2150 -885 2155
rect -925 2120 -920 2150
rect -890 2120 -885 2150
rect -925 2115 -885 2120
rect -805 2150 -765 2155
rect -805 2120 -800 2150
rect -770 2120 -765 2150
rect -805 2115 -765 2120
rect -685 2150 -645 2155
rect -685 2120 -680 2150
rect -650 2120 -645 2150
rect -685 2115 -645 2120
rect -565 2150 -525 2155
rect -565 2120 -560 2150
rect -530 2120 -525 2150
rect -565 2115 -525 2120
rect -445 2150 -405 2155
rect -445 2120 -440 2150
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2120 -240 2150
rect -280 2115 -240 2120
rect -270 1730 -250 2115
rect -1105 1725 -1065 1730
rect -1105 1695 -1100 1725
rect -1070 1695 -1065 1725
rect -1105 1690 -1065 1695
rect -985 1725 -945 1730
rect -985 1695 -980 1725
rect -950 1695 -945 1725
rect -985 1690 -945 1695
rect -865 1725 -825 1730
rect -865 1695 -860 1725
rect -830 1695 -825 1725
rect -865 1690 -825 1695
rect -800 1720 -770 1730
rect -800 1700 -795 1720
rect -775 1700 -770 1720
rect -800 1690 -770 1700
rect -745 1725 -705 1730
rect -745 1695 -740 1725
rect -710 1695 -705 1725
rect -745 1690 -705 1695
rect -625 1725 -585 1730
rect -625 1695 -620 1725
rect -590 1695 -585 1725
rect -625 1690 -585 1695
rect -505 1725 -465 1730
rect -505 1695 -500 1725
rect -470 1695 -465 1725
rect -505 1690 -465 1695
rect -280 1725 -240 1730
rect -280 1695 -275 1725
rect -245 1695 -240 1725
rect -280 1690 -240 1695
rect -795 1630 -775 1690
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1640 -330 1670
rect -370 1635 -330 1640
rect -805 1625 -765 1630
rect -805 1595 -800 1625
rect -770 1595 -765 1625
rect -805 1590 -765 1595
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -1440 1430 -1420 1505
rect -1135 1485 -1095 1490
rect -1135 1455 -1130 1485
rect -1100 1455 -1095 1485
rect -1135 1450 -1095 1455
rect -1025 1485 -985 1490
rect -1025 1455 -1020 1485
rect -990 1455 -985 1485
rect -1025 1450 -985 1455
rect -915 1485 -875 1490
rect -915 1455 -910 1485
rect -880 1455 -875 1485
rect -915 1450 -875 1455
rect -805 1485 -765 1490
rect -805 1455 -800 1485
rect -770 1455 -765 1485
rect -805 1450 -765 1455
rect -695 1485 -655 1490
rect -695 1455 -690 1485
rect -660 1455 -655 1485
rect -695 1450 -655 1455
rect -585 1485 -545 1490
rect -585 1455 -580 1485
rect -550 1455 -545 1485
rect -585 1450 -545 1455
rect -475 1485 -435 1490
rect -475 1455 -470 1485
rect -440 1455 -435 1485
rect -475 1450 -435 1455
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -360 965 -340 1635
rect -225 1490 -205 2170
rect -40 2150 0 2155
rect -40 2120 -35 2150
rect -5 2120 0 2150
rect -40 2115 0 2120
rect 80 2150 120 2155
rect 80 2120 85 2150
rect 115 2120 120 2150
rect 80 2115 120 2120
rect 200 2150 240 2155
rect 200 2120 205 2150
rect 235 2120 240 2150
rect 200 2115 240 2120
rect 320 2150 360 2155
rect 320 2120 325 2150
rect 355 2120 360 2150
rect 320 2115 360 2120
rect 440 2150 480 2155
rect 440 2120 445 2150
rect 475 2120 480 2150
rect 440 2115 480 2120
rect 560 2150 600 2155
rect 560 2120 565 2150
rect 595 2120 600 2150
rect 560 2115 600 2120
rect 680 2150 720 2155
rect 680 2120 685 2150
rect 715 2120 720 2150
rect 680 2115 720 2120
rect 20 1725 60 1730
rect 20 1695 25 1725
rect 55 1695 60 1725
rect 20 1690 60 1695
rect 140 1725 180 1730
rect 140 1695 145 1725
rect 175 1695 180 1725
rect 140 1690 180 1695
rect 260 1725 300 1730
rect 260 1695 265 1725
rect 295 1695 300 1725
rect 260 1690 300 1695
rect 325 1720 355 1730
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 380 1725 420 1730
rect 380 1695 385 1725
rect 415 1695 420 1725
rect 380 1690 420 1695
rect 500 1725 540 1730
rect 500 1695 505 1725
rect 535 1695 540 1725
rect 500 1690 540 1695
rect 620 1725 660 1730
rect 620 1695 625 1725
rect 655 1695 660 1725
rect 620 1690 660 1695
rect 30 1675 50 1690
rect 330 1675 350 1690
rect 790 1675 810 2270
rect 835 2210 855 2520
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1519 2305 1549 2310
rect 1519 2270 1549 2275
rect 1573 2300 1613 2310
rect 1573 2280 1583 2300
rect 1603 2280 1613 2300
rect 1573 2270 1613 2280
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2230 920 2260
rect 1055 2255 1075 2270
rect 1583 2255 1603 2270
rect 880 2225 920 2230
rect 1045 2250 1085 2255
rect 825 2205 865 2210
rect 825 2175 830 2205
rect 860 2175 865 2205
rect 825 2170 865 2175
rect 20 1670 60 1675
rect 20 1640 25 1670
rect 55 1640 60 1670
rect 20 1635 60 1640
rect 320 1670 360 1675
rect 320 1640 325 1670
rect 355 1640 360 1670
rect 320 1635 360 1640
rect 780 1670 820 1675
rect 780 1640 785 1670
rect 815 1640 820 1670
rect 780 1635 820 1640
rect 880 1630 900 2225
rect 1045 2220 1050 2250
rect 1080 2220 1085 2250
rect 1045 2215 1085 2220
rect 1573 2250 1613 2255
rect 1573 2220 1578 2250
rect 1608 2220 1613 2250
rect 1573 2215 1613 2220
rect 1885 2205 1925 2210
rect 1885 2175 1890 2205
rect 1920 2175 1925 2205
rect 1885 2170 1925 2175
rect 2455 2205 2495 2210
rect 2455 2175 2460 2205
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2120 1010 2150
rect 970 2115 1010 2120
rect 1090 2150 1130 2155
rect 1090 2120 1095 2150
rect 1125 2120 1130 2150
rect 1090 2115 1130 2120
rect 1210 2150 1250 2155
rect 1210 2120 1215 2150
rect 1245 2120 1250 2150
rect 1210 2115 1250 2120
rect 1330 2150 1370 2155
rect 1330 2120 1335 2150
rect 1365 2120 1370 2150
rect 1330 2115 1370 2120
rect 1450 2150 1490 2155
rect 1450 2120 1455 2150
rect 1485 2120 1490 2150
rect 1450 2115 1490 2120
rect 1570 2150 1610 2155
rect 1570 2120 1575 2150
rect 1605 2120 1610 2150
rect 1570 2115 1610 2120
rect 1690 2150 1730 2155
rect 1690 2120 1695 2150
rect 1725 2120 1730 2150
rect 1690 2115 1730 2120
rect 1030 1725 1070 1730
rect 1030 1695 1035 1725
rect 1065 1695 1070 1725
rect 1030 1690 1070 1695
rect 1150 1725 1190 1730
rect 1150 1695 1155 1725
rect 1185 1695 1190 1725
rect 1150 1690 1190 1695
rect 1270 1725 1310 1730
rect 1270 1695 1275 1725
rect 1305 1695 1310 1725
rect 1270 1690 1310 1695
rect 1335 1720 1365 1730
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 1390 1725 1430 1730
rect 1390 1695 1395 1725
rect 1425 1695 1430 1725
rect 1390 1690 1430 1695
rect 1510 1725 1550 1730
rect 1510 1695 1515 1725
rect 1545 1695 1550 1725
rect 1510 1690 1550 1695
rect 1630 1725 1670 1730
rect 1630 1695 1635 1725
rect 1665 1695 1670 1725
rect 1630 1690 1670 1695
rect 1340 1675 1360 1690
rect 1640 1675 1660 1690
rect 1330 1670 1370 1675
rect 1330 1640 1335 1670
rect 1365 1640 1370 1670
rect 1330 1635 1370 1640
rect 1630 1670 1670 1675
rect 1630 1640 1635 1670
rect 1665 1640 1670 1670
rect 1630 1635 1670 1640
rect 870 1600 875 1630
rect 905 1600 910 1630
rect 1895 1585 1915 2170
rect 2465 2155 2485 2170
rect 1930 2150 1970 2155
rect 1930 2120 1935 2150
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2120 2135 2150
rect 2095 2115 2135 2120
rect 2215 2150 2255 2155
rect 2215 2120 2220 2150
rect 2250 2120 2255 2150
rect 2215 2115 2255 2120
rect 2335 2150 2375 2155
rect 2335 2120 2340 2150
rect 2370 2120 2375 2150
rect 2335 2115 2375 2120
rect 2455 2150 2495 2155
rect 2455 2120 2460 2150
rect 2490 2120 2495 2150
rect 2455 2115 2495 2120
rect 2575 2150 2615 2155
rect 2575 2120 2580 2150
rect 2610 2120 2615 2150
rect 2575 2115 2615 2120
rect 2695 2150 2735 2155
rect 2695 2120 2700 2150
rect 2730 2120 2735 2150
rect 2695 2115 2735 2120
rect 2815 2150 2855 2155
rect 2815 2120 2820 2150
rect 2850 2120 2855 2150
rect 2815 2115 2855 2120
rect 1940 1730 1960 2115
rect 1930 1725 1970 1730
rect 1930 1695 1935 1725
rect 1965 1695 1970 1725
rect 1930 1690 1970 1695
rect 2155 1725 2195 1730
rect 2155 1695 2160 1725
rect 2190 1695 2195 1725
rect 2155 1690 2195 1695
rect 2275 1725 2315 1730
rect 2275 1695 2280 1725
rect 2310 1695 2315 1725
rect 2275 1690 2315 1695
rect 2395 1725 2435 1730
rect 2395 1695 2400 1725
rect 2430 1695 2435 1725
rect 2395 1690 2435 1695
rect 2460 1720 2490 1730
rect 2460 1700 2465 1720
rect 2485 1700 2490 1720
rect 2460 1690 2490 1700
rect 2515 1725 2555 1730
rect 2515 1695 2520 1725
rect 2550 1695 2555 1725
rect 2515 1690 2555 1695
rect 2635 1725 2675 1730
rect 2635 1695 2640 1725
rect 2670 1695 2675 1725
rect 2635 1690 2675 1695
rect 2755 1725 2795 1730
rect 2755 1695 2760 1725
rect 2790 1695 2795 1725
rect 2755 1690 2795 1695
rect 2020 1670 2060 1675
rect 2020 1640 2025 1670
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect 455 1580 495 1585
rect 455 1550 460 1580
rect 490 1550 495 1580
rect 455 1545 495 1550
rect 625 1580 655 1585
rect 625 1545 655 1550
rect 785 1580 825 1585
rect 785 1550 790 1580
rect 820 1550 825 1580
rect 785 1545 825 1550
rect 865 1580 905 1585
rect 865 1550 870 1580
rect 900 1550 905 1580
rect 865 1545 905 1550
rect 1035 1580 1065 1585
rect 1035 1545 1065 1550
rect 1195 1580 1235 1585
rect 1195 1550 1200 1580
rect 1230 1550 1235 1580
rect 1195 1545 1235 1550
rect 1885 1580 1925 1585
rect 1885 1550 1890 1580
rect 1920 1550 1925 1580
rect 1885 1545 1925 1550
rect 565 1535 605 1540
rect 565 1505 570 1535
rect 600 1505 605 1535
rect 565 1500 605 1505
rect 675 1535 715 1540
rect 675 1505 680 1535
rect 710 1505 715 1535
rect 675 1500 715 1505
rect 975 1535 1015 1540
rect 975 1505 980 1535
rect 1010 1505 1015 1535
rect 975 1500 1015 1505
rect 1085 1535 1125 1540
rect 1085 1505 1090 1535
rect 1120 1505 1125 1535
rect 1085 1500 1125 1505
rect 1895 1490 1915 1545
rect -235 1485 -195 1490
rect -235 1455 -230 1485
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 1885 1485 1925 1490
rect 1885 1455 1890 1485
rect 1920 1455 1925 1485
rect 1885 1450 1925 1455
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1075 -285 1105
rect -325 1070 -285 1075
rect -370 960 -330 965
rect -370 930 -365 960
rect -335 930 -330 960
rect -370 925 -330 930
rect -1501 815 -1360 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -1080 810 -1040 815
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 730 -1500 760
rect -1540 725 -1500 730
rect -1530 360 -1510 725
rect -1440 720 -1420 785
rect -1080 780 -1075 810
rect -1045 780 -1040 810
rect -1080 775 -1040 780
rect -970 810 -930 815
rect -970 780 -965 810
rect -935 780 -930 810
rect -970 775 -930 780
rect -860 810 -820 815
rect -750 810 -710 815
rect -860 780 -855 810
rect -825 780 -820 810
rect -860 775 -820 780
rect -800 800 -770 810
rect -800 780 -795 800
rect -775 780 -770 800
rect -960 760 -940 775
rect -800 770 -770 780
rect -750 780 -745 810
rect -715 780 -710 810
rect -750 775 -710 780
rect -640 810 -600 815
rect -640 780 -635 810
rect -605 780 -600 810
rect -640 775 -600 780
rect -530 810 -490 815
rect -530 780 -525 810
rect -495 780 -490 810
rect -530 775 -490 780
rect -970 730 -965 760
rect -935 730 -930 760
rect -795 720 -775 770
rect -530 730 -525 760
rect -495 730 -490 760
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 685 -1410 715
rect -1450 680 -1410 685
rect -805 715 -765 720
rect -805 685 -800 715
rect -770 685 -765 715
rect -805 680 -765 685
rect -520 675 -500 730
rect -360 720 -340 925
rect -370 715 -330 720
rect -370 685 -365 715
rect -335 685 -330 715
rect -370 680 -330 685
rect -1145 670 -1105 675
rect -1145 640 -1140 670
rect -1110 640 -1105 670
rect -1145 635 -1105 640
rect -1080 670 -1040 675
rect -1080 640 -1075 670
rect -1045 640 -1040 670
rect -1080 635 -1040 640
rect -970 670 -930 675
rect -970 640 -965 670
rect -935 640 -930 670
rect -970 635 -930 640
rect -860 670 -820 675
rect -860 640 -855 670
rect -825 640 -820 670
rect -860 635 -820 640
rect -750 670 -710 675
rect -750 640 -745 670
rect -715 640 -710 670
rect -750 635 -710 640
rect -640 670 -600 675
rect -640 640 -635 670
rect -605 640 -600 670
rect -640 635 -600 640
rect -530 670 -490 675
rect -530 640 -525 670
rect -495 640 -490 670
rect -530 635 -490 640
rect -465 670 -425 675
rect -465 640 -460 670
rect -430 640 -425 670
rect -465 635 -425 640
rect -1270 395 -1230 400
rect -1270 365 -1265 395
rect -1235 365 -1230 395
rect -1270 360 -1230 365
rect -1025 395 -985 400
rect -1025 365 -1020 395
rect -990 365 -985 395
rect -1025 360 -985 365
rect -915 395 -875 400
rect -915 365 -910 395
rect -880 365 -875 395
rect -915 360 -875 365
rect -805 395 -765 400
rect -805 365 -800 395
rect -770 365 -765 395
rect -805 360 -765 365
rect -745 390 -715 400
rect -745 370 -740 390
rect -720 370 -715 390
rect -745 360 -715 370
rect -695 395 -655 400
rect -695 365 -690 395
rect -660 365 -655 395
rect -695 360 -655 365
rect -585 395 -545 400
rect -585 365 -580 395
rect -550 365 -545 395
rect -585 360 -545 365
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect -1545 310 -1495 320
rect -1530 -295 -1510 310
rect -1490 -120 -1486 -85
rect -1459 -120 -1455 -85
rect -1430 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -120 -1275 -85
rect -1485 -185 -1460 -120
rect -1370 -145 -1335 -120
rect -1260 -140 -1240 360
rect -740 345 -720 360
rect -360 345 -340 680
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 310 -710 340
rect -750 305 -710 310
rect -370 340 -330 345
rect -370 310 -365 340
rect -335 310 -330 340
rect -370 305 -330 310
rect -740 290 -720 305
rect -1225 285 -1185 290
rect -1225 255 -1220 285
rect -1190 255 -1185 285
rect -1225 250 -1185 255
rect -1025 285 -985 290
rect -1025 255 -1020 285
rect -990 255 -985 285
rect -1025 250 -985 255
rect -915 285 -875 290
rect -915 255 -910 285
rect -880 255 -875 285
rect -915 250 -875 255
rect -805 285 -765 290
rect -805 255 -800 285
rect -770 255 -765 285
rect -805 250 -765 255
rect -745 280 -715 290
rect -745 260 -740 280
rect -720 260 -715 280
rect -745 250 -715 260
rect -695 285 -655 290
rect -695 255 -690 285
rect -660 255 -655 285
rect -695 250 -655 255
rect -585 285 -545 290
rect -585 255 -580 285
rect -550 255 -545 285
rect -585 250 -545 255
rect -1215 -85 -1195 250
rect -1225 -90 -1185 -85
rect -1225 -120 -1220 -90
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -1145 -95 -1105 -85
rect -1145 -115 -1135 -95
rect -1115 -115 -1105 -95
rect -1145 -125 -1105 -115
rect -1080 -90 -1040 -85
rect -1080 -120 -1075 -90
rect -1045 -120 -1040 -90
rect -1080 -125 -1040 -120
rect -970 -90 -930 -85
rect -970 -120 -965 -90
rect -935 -120 -930 -90
rect -970 -125 -930 -120
rect -860 -90 -820 -85
rect -860 -120 -855 -90
rect -825 -120 -820 -90
rect -860 -125 -820 -120
rect -750 -90 -710 -85
rect -750 -120 -745 -90
rect -715 -120 -710 -90
rect -750 -125 -710 -120
rect -640 -90 -600 -85
rect -640 -120 -635 -90
rect -605 -120 -600 -90
rect -640 -125 -600 -120
rect -530 -90 -490 -85
rect -530 -120 -525 -90
rect -495 -120 -490 -90
rect -530 -125 -490 -120
rect -465 -95 -425 -85
rect -465 -115 -455 -95
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect -1135 -140 -1115 -125
rect -455 -140 -435 -125
rect -1370 -180 -1335 -175
rect -1270 -145 -1230 -140
rect -1270 -175 -1265 -145
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1145 -145 -1105 -140
rect -1145 -175 -1140 -145
rect -1110 -175 -1105 -145
rect -1145 -180 -1105 -175
rect -465 -145 -425 -140
rect -465 -175 -460 -145
rect -430 -175 -425 -145
rect -465 -180 -425 -175
rect -1490 -190 -1455 -185
rect -315 -190 -295 1070
rect -280 770 -240 775
rect -280 740 -275 770
rect -245 740 -240 770
rect -280 735 -240 740
rect -270 -140 -250 735
rect -225 675 -205 1450
rect 505 1225 535 1230
rect 745 1225 775 1230
rect 505 1190 535 1195
rect 552 1210 582 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1215 660 1220
rect 620 1185 625 1215
rect 655 1185 660 1215
rect 620 1180 660 1185
rect 698 1210 728 1220
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 745 1190 775 1195
rect 915 1220 945 1230
rect 1155 1220 1185 1230
rect 915 1200 920 1220
rect 940 1200 945 1220
rect 915 1190 945 1200
rect 962 1210 992 1220
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 698 1180 728 1190
rect 555 1160 575 1180
rect 545 1155 585 1160
rect 545 1125 550 1155
rect 580 1125 585 1155
rect 545 1120 585 1125
rect 705 1110 725 1180
rect 690 1105 730 1110
rect 690 1075 695 1105
rect 725 1075 730 1105
rect 690 1070 730 1075
rect 915 1065 935 1190
rect 962 1180 992 1190
rect 1030 1215 1070 1220
rect 1030 1185 1035 1215
rect 1065 1185 1070 1215
rect 1030 1180 1070 1185
rect 1108 1210 1138 1220
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1155 1200 1160 1220
rect 1180 1200 1185 1220
rect 1155 1190 1185 1200
rect 1108 1180 1138 1190
rect 965 1110 985 1180
rect 1115 1160 1135 1180
rect 1105 1155 1145 1160
rect 1105 1125 1110 1155
rect 1140 1125 1145 1155
rect 1105 1120 1145 1125
rect 960 1105 1000 1110
rect 960 1075 965 1105
rect 995 1075 1000 1105
rect 960 1070 1000 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1030 835 1060
rect 795 1025 835 1030
rect 905 1060 945 1065
rect 905 1030 910 1060
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 805 1010 825 1025
rect 1165 1020 1185 1190
rect 1155 1015 1195 1020
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 975 920 1005
rect 1155 985 1160 1015
rect 1190 985 1195 1015
rect 1155 980 1195 985
rect 1840 1005 1880 1010
rect 880 970 920 975
rect 1840 975 1845 1005
rect 1875 975 1880 1005
rect 1840 970 1880 975
rect -50 960 -10 965
rect -50 930 -45 960
rect -15 930 -10 960
rect -50 925 -10 930
rect 60 960 100 965
rect 60 930 65 960
rect 95 930 100 960
rect 60 925 100 930
rect 170 960 210 965
rect 170 930 175 960
rect 205 930 210 960
rect 170 925 210 930
rect 280 960 320 965
rect 280 930 285 960
rect 315 930 320 960
rect 280 925 320 930
rect 390 960 430 965
rect 390 930 395 960
rect 425 930 430 960
rect 390 925 430 930
rect 500 960 540 965
rect 500 930 505 960
rect 535 930 540 960
rect 805 930 825 970
rect 890 930 910 970
rect 1150 960 1190 965
rect 1150 930 1155 960
rect 1185 930 1190 960
rect 500 925 540 930
rect -40 910 -20 925
rect 70 910 90 925
rect 180 910 200 925
rect 290 910 310 925
rect 400 910 420 925
rect 510 910 530 925
rect 795 920 835 930
rect -180 905 -140 910
rect -180 875 -175 905
rect -145 875 -140 905
rect -180 870 -140 875
rect -50 900 -10 910
rect -50 880 -40 900
rect -20 880 -10 900
rect -50 870 -10 880
rect 60 900 100 910
rect 60 880 70 900
rect 90 880 100 900
rect 60 870 100 880
rect 170 900 210 910
rect 170 880 180 900
rect 200 880 210 900
rect 170 870 210 880
rect 230 905 260 910
rect 230 870 260 875
rect 280 900 320 910
rect 280 880 290 900
rect 310 880 320 900
rect 280 870 320 880
rect 390 900 430 910
rect 390 880 400 900
rect 420 880 430 900
rect 390 870 430 880
rect 500 900 540 910
rect 500 880 510 900
rect 530 880 540 900
rect 795 900 805 920
rect 825 900 835 920
rect 795 890 835 900
rect 880 920 920 930
rect 1150 925 1190 930
rect 1260 960 1300 965
rect 1260 930 1265 960
rect 1295 930 1300 960
rect 1260 925 1300 930
rect 1370 960 1410 965
rect 1370 930 1375 960
rect 1405 930 1410 960
rect 1370 925 1410 930
rect 1480 960 1520 965
rect 1480 930 1485 960
rect 1515 930 1520 960
rect 1480 925 1520 930
rect 1590 960 1630 965
rect 1590 930 1595 960
rect 1625 930 1630 960
rect 1590 925 1630 930
rect 1700 960 1740 965
rect 1700 930 1705 960
rect 1735 930 1740 960
rect 1700 925 1740 930
rect 880 900 890 920
rect 910 900 920 920
rect 1160 910 1180 925
rect 1270 910 1290 925
rect 1380 910 1400 925
rect 1490 910 1510 925
rect 1600 910 1620 925
rect 1710 910 1730 925
rect 880 890 920 900
rect 1150 900 1190 910
rect 500 870 540 880
rect 1150 880 1160 900
rect 1180 880 1190 900
rect 1150 870 1190 880
rect 1260 900 1300 910
rect 1260 880 1270 900
rect 1290 880 1300 900
rect 1260 870 1300 880
rect 1370 900 1410 910
rect 1370 880 1380 900
rect 1400 880 1410 900
rect 1370 870 1410 880
rect 1430 905 1460 910
rect 1430 870 1460 875
rect 1480 900 1520 910
rect 1480 880 1490 900
rect 1510 880 1520 900
rect 1480 870 1520 880
rect 1590 900 1630 910
rect 1590 880 1600 900
rect 1620 880 1630 900
rect 1590 870 1630 880
rect 1700 900 1740 910
rect 1700 880 1710 900
rect 1730 880 1740 900
rect 1700 870 1740 880
rect -235 670 -195 675
rect -235 640 -230 670
rect -200 640 -195 670
rect -235 635 -195 640
rect -225 -85 -205 635
rect -235 -90 -195 -85
rect -235 -120 -230 -90
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect -280 -145 -240 -140
rect -280 -175 -275 -145
rect -245 -175 -240 -145
rect -1490 -225 -1455 -220
rect -325 -220 -320 -190
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect -1210 -245 -1175 -240
rect -1210 -280 -1175 -275
rect -625 -245 -585 -240
rect -625 -275 -620 -245
rect -590 -275 -585 -245
rect -625 -280 -585 -275
rect -1540 -300 -1500 -295
rect -1540 -330 -1535 -300
rect -1505 -330 -1500 -300
rect -1540 -335 -1500 -330
rect -1205 -380 -1180 -280
rect -615 -295 -595 -280
rect -1150 -300 -1115 -295
rect -1150 -335 -1115 -330
rect -925 -300 -885 -295
rect -925 -330 -920 -300
rect -890 -330 -885 -300
rect -925 -335 -885 -330
rect -725 -300 -685 -295
rect -725 -330 -720 -300
rect -690 -330 -685 -300
rect -725 -335 -685 -330
rect -625 -305 -585 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -335 -585 -325
rect -525 -300 -485 -295
rect -525 -330 -520 -300
rect -490 -330 -485 -300
rect -525 -335 -485 -330
rect -1145 -380 -1120 -335
rect -1210 -415 -1206 -380
rect -1179 -415 -1175 -380
rect -1150 -415 -1146 -380
rect -1119 -415 -1115 -380
rect -1025 -1075 -985 -1070
rect -1025 -1105 -1020 -1075
rect -990 -1105 -985 -1075
rect -1025 -1110 -985 -1105
rect -825 -1075 -785 -1070
rect -825 -1105 -820 -1075
rect -790 -1105 -785 -1075
rect -825 -1110 -785 -1105
rect -725 -1075 -685 -1070
rect -725 -1105 -720 -1075
rect -690 -1105 -685 -1075
rect -725 -1110 -685 -1105
rect -625 -1075 -585 -1070
rect -625 -1105 -620 -1075
rect -590 -1105 -585 -1075
rect -625 -1110 -585 -1105
rect -425 -1075 -385 -1070
rect -425 -1105 -420 -1075
rect -390 -1105 -385 -1075
rect -425 -1110 -385 -1105
rect -715 -1170 -695 -1110
rect -270 -1170 -250 -175
rect -235 -245 -195 -240
rect -235 -275 -230 -245
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect -225 -350 -205 -280
rect -235 -355 -195 -350
rect -235 -385 -230 -355
rect -200 -385 -195 -355
rect -235 -390 -195 -385
rect -180 -895 -160 870
rect -100 675 -70 685
rect -100 655 -95 675
rect -75 655 -70 675
rect -100 645 -70 655
rect 5 680 45 685
rect 5 650 10 680
rect 40 650 45 680
rect 5 645 45 650
rect 115 680 155 685
rect 115 650 120 680
rect 150 650 155 680
rect 115 645 155 650
rect 225 680 265 685
rect 225 650 230 680
rect 260 650 265 680
rect 225 645 265 650
rect 335 680 375 685
rect 335 650 340 680
rect 370 650 375 680
rect 335 645 375 650
rect 445 680 485 685
rect 445 650 450 680
rect 480 650 485 680
rect 445 645 485 650
rect 560 675 590 685
rect 560 655 565 675
rect 585 655 590 675
rect 560 645 590 655
rect 1100 675 1130 685
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1100 645 1130 655
rect 1205 680 1245 685
rect 1205 650 1210 680
rect 1240 650 1245 680
rect 1205 645 1245 650
rect 1315 680 1355 685
rect 1315 650 1320 680
rect 1350 650 1355 680
rect 1315 645 1355 650
rect 1425 680 1465 685
rect 1425 650 1430 680
rect 1460 650 1465 680
rect 1425 645 1465 650
rect 1535 680 1575 685
rect 1535 650 1540 680
rect 1570 650 1575 680
rect 1535 645 1575 650
rect 1645 680 1685 685
rect 1645 650 1650 680
rect 1680 650 1685 680
rect 1645 645 1685 650
rect 1760 675 1790 685
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1760 645 1790 655
rect -95 630 -75 645
rect -105 625 -65 630
rect -105 595 -100 625
rect -70 595 -65 625
rect -105 590 -65 595
rect 235 570 255 645
rect 565 630 585 645
rect 1105 630 1125 645
rect 555 625 595 630
rect 555 595 560 625
rect 590 595 595 625
rect 1095 625 1135 630
rect 555 590 595 595
rect 715 605 755 610
rect 715 575 720 605
rect 750 575 755 605
rect 715 570 755 575
rect 825 605 865 610
rect 825 575 830 605
rect 860 575 865 605
rect 825 570 865 575
rect 935 605 975 610
rect 935 575 940 605
rect 970 575 975 605
rect 1095 595 1100 625
rect 1130 595 1135 625
rect 1095 590 1135 595
rect 935 570 975 575
rect 1435 570 1455 645
rect 1765 630 1785 645
rect 1755 625 1795 630
rect 1755 595 1760 625
rect 1790 595 1795 625
rect 1755 590 1795 595
rect 230 565 260 570
rect -50 555 -10 560
rect -50 525 -45 555
rect -15 525 -10 555
rect -50 520 -10 525
rect 60 555 100 560
rect 60 525 65 555
rect 95 525 100 555
rect 60 520 100 525
rect 170 555 210 560
rect 170 525 175 555
rect 205 525 210 555
rect 230 530 260 535
rect 280 555 320 560
rect 170 520 210 525
rect 280 525 285 555
rect 315 525 320 555
rect 280 520 320 525
rect 390 555 430 560
rect 390 525 395 555
rect 425 525 430 555
rect 390 520 430 525
rect 500 555 540 560
rect 500 525 505 555
rect 535 525 540 555
rect 500 520 540 525
rect 725 510 745 570
rect 945 510 965 570
rect 1430 565 1460 570
rect 1150 555 1190 560
rect 1150 525 1155 555
rect 1185 525 1190 555
rect 1150 520 1190 525
rect 1260 555 1300 560
rect 1260 525 1265 555
rect 1295 525 1300 555
rect 1260 520 1300 525
rect 1370 555 1410 560
rect 1370 525 1375 555
rect 1405 525 1410 555
rect 1430 530 1460 535
rect 1480 555 1520 560
rect 1370 520 1410 525
rect 1480 525 1485 555
rect 1515 525 1520 555
rect 1480 520 1520 525
rect 1590 555 1630 560
rect 1590 525 1595 555
rect 1625 525 1630 555
rect 1590 520 1630 525
rect 1700 555 1740 560
rect 1700 525 1705 555
rect 1735 525 1740 555
rect 1700 520 1740 525
rect 230 505 260 510
rect 230 470 260 475
rect 715 500 755 510
rect 715 480 725 500
rect 745 480 755 500
rect 715 470 755 480
rect 795 505 825 510
rect 795 470 825 475
rect 865 505 895 510
rect 865 470 895 475
rect 935 500 975 510
rect 935 480 945 500
rect 965 480 975 500
rect 935 470 975 480
rect 1430 505 1460 510
rect 1430 470 1460 475
rect -100 280 -70 290
rect -100 260 -95 280
rect -75 260 -70 280
rect -100 250 -70 260
rect 5 285 45 290
rect 5 255 10 285
rect 40 255 45 285
rect 5 250 45 255
rect 115 285 155 290
rect 115 255 120 285
rect 150 255 155 285
rect 115 250 155 255
rect 225 285 265 290
rect 225 255 230 285
rect 260 255 265 285
rect 225 250 265 255
rect 335 285 375 290
rect 335 255 340 285
rect 370 255 375 285
rect 335 250 375 255
rect 445 285 485 290
rect 445 255 450 285
rect 480 255 485 285
rect 445 250 485 255
rect 600 280 630 290
rect 600 260 605 280
rect 625 260 630 280
rect 600 250 630 260
rect 775 280 805 290
rect 775 260 780 280
rect 800 260 805 280
rect 775 250 805 260
rect 830 280 860 290
rect 830 260 835 280
rect 855 260 860 280
rect 830 250 860 260
rect 885 280 915 290
rect 885 260 890 280
rect 910 260 915 280
rect 885 250 915 260
rect 1060 280 1090 290
rect 1060 260 1065 280
rect 1085 260 1090 280
rect 1060 250 1090 260
rect 1205 285 1245 290
rect 1205 255 1210 285
rect 1240 255 1245 285
rect 1205 250 1245 255
rect 1265 285 1295 290
rect 1265 250 1295 255
rect 1315 285 1355 290
rect 1315 255 1320 285
rect 1350 255 1355 285
rect 1315 250 1355 255
rect 1425 285 1465 290
rect 1425 255 1430 285
rect 1460 255 1465 285
rect 1425 250 1465 255
rect 1535 285 1575 290
rect 1535 255 1540 285
rect 1570 255 1575 285
rect 1535 250 1575 255
rect 1645 285 1685 290
rect 1645 255 1650 285
rect 1680 255 1685 285
rect 1645 250 1685 255
rect 1760 280 1790 290
rect 1760 260 1765 280
rect 1785 260 1790 280
rect 1760 250 1790 260
rect -95 -305 -75 250
rect 440 15 480 20
rect 440 -15 445 15
rect 475 -15 480 15
rect 440 -20 480 -15
rect -105 -310 -65 -305
rect -105 -340 -100 -310
rect -70 -340 -65 -310
rect -105 -345 -65 -340
rect 450 -475 470 -20
rect 605 -305 625 250
rect 780 235 800 250
rect 780 230 820 235
rect 780 200 785 230
rect 815 200 820 230
rect 780 195 820 200
rect 795 125 815 195
rect 835 180 855 250
rect 890 235 910 250
rect 870 230 910 235
rect 870 200 875 230
rect 905 200 910 230
rect 870 195 910 200
rect 835 175 895 180
rect 835 145 860 175
rect 890 145 895 175
rect 835 140 895 145
rect 795 120 855 125
rect 795 90 800 120
rect 830 90 855 120
rect 795 85 855 90
rect 780 65 820 70
rect 780 35 785 65
rect 815 35 820 65
rect 780 30 820 35
rect 780 15 800 30
rect 835 20 855 85
rect 875 70 895 140
rect 870 65 910 70
rect 870 35 875 65
rect 905 35 910 65
rect 870 30 910 35
rect 830 15 860 20
rect 890 15 910 30
rect 775 5 805 15
rect 775 -15 780 5
rect 800 -15 805 5
rect 775 -25 805 -15
rect 830 -20 860 -15
rect 885 5 915 15
rect 885 -15 890 5
rect 910 -15 915 5
rect 885 -25 915 -15
rect 1065 -305 1085 250
rect 595 -310 635 -305
rect 595 -340 600 -310
rect 630 -340 635 -310
rect 595 -345 635 -340
rect 715 -310 755 -305
rect 715 -340 720 -310
rect 750 -340 755 -310
rect 715 -345 755 -340
rect 825 -310 865 -305
rect 825 -340 830 -310
rect 860 -340 865 -310
rect 825 -345 865 -340
rect 935 -310 975 -305
rect 935 -340 940 -310
rect 970 -340 975 -310
rect 935 -345 975 -340
rect 1065 -310 1105 -305
rect 1065 -340 1070 -310
rect 1100 -340 1105 -310
rect 1065 -345 1105 -340
rect 1270 -475 1290 250
rect 1760 -305 1780 250
rect 1750 -310 1790 -305
rect 1750 -340 1755 -310
rect 1785 -340 1790 -310
rect 1750 -345 1790 -340
rect 1850 -420 1870 970
rect 1895 675 1915 1450
rect 1975 1105 2015 1110
rect 1975 1075 1980 1105
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 1930 770 1970 775
rect 1930 740 1935 770
rect 1965 740 1970 770
rect 1930 735 1970 740
rect 1885 670 1925 675
rect 1885 640 1890 670
rect 1920 640 1925 670
rect 1885 635 1925 640
rect 1895 -85 1915 635
rect 1940 620 1960 735
rect 1930 615 1970 620
rect 1930 585 1935 615
rect 1965 585 1970 615
rect 1930 580 1970 585
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -120 1925 -90
rect 1885 -125 1925 -120
rect 1940 -140 1960 580
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -175 1970 -145
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -275 1925 -245
rect 1885 -280 1925 -275
rect 1895 -350 1915 -280
rect 1940 -305 1960 -175
rect 1985 -190 2005 1070
rect 2030 965 2050 1635
rect 2465 1630 2485 1690
rect 2455 1625 2495 1630
rect 2455 1595 2460 1625
rect 2490 1595 2495 1625
rect 2455 1590 2495 1595
rect 3100 1490 3140 1495
rect 2125 1485 2165 1490
rect 2125 1455 2130 1485
rect 2160 1455 2165 1485
rect 2125 1450 2165 1455
rect 2235 1485 2275 1490
rect 2235 1455 2240 1485
rect 2270 1455 2275 1485
rect 2235 1450 2275 1455
rect 2345 1485 2385 1490
rect 2345 1455 2350 1485
rect 2380 1455 2385 1485
rect 2345 1450 2385 1455
rect 2455 1485 2495 1490
rect 2455 1455 2460 1485
rect 2490 1455 2495 1485
rect 2455 1450 2495 1455
rect 2565 1485 2605 1490
rect 2565 1455 2570 1485
rect 2600 1455 2605 1485
rect 2565 1450 2605 1455
rect 2675 1485 2715 1490
rect 2675 1455 2680 1485
rect 2710 1455 2715 1485
rect 2675 1450 2715 1455
rect 2785 1485 2825 1490
rect 2785 1455 2790 1485
rect 2820 1455 2825 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2785 1450 2825 1455
rect 3110 1430 3130 1455
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2020 960 2060 965
rect 2020 930 2025 960
rect 2055 930 2060 960
rect 2020 925 2060 930
rect 2030 720 2050 925
rect 3050 815 3191 825
rect 2180 810 2220 815
rect 2180 780 2185 810
rect 2215 780 2220 810
rect 2180 775 2220 780
rect 2290 810 2330 815
rect 2290 780 2295 810
rect 2325 780 2330 810
rect 2290 775 2330 780
rect 2400 810 2440 815
rect 2510 810 2550 815
rect 2400 780 2405 810
rect 2435 780 2440 810
rect 2400 775 2440 780
rect 2460 800 2490 810
rect 2460 780 2465 800
rect 2485 780 2490 800
rect 2460 770 2490 780
rect 2510 780 2515 810
rect 2545 780 2550 810
rect 2510 775 2550 780
rect 2620 810 2660 815
rect 2620 780 2625 810
rect 2655 780 2660 810
rect 2620 775 2660 780
rect 2730 810 2770 815
rect 2730 780 2735 810
rect 2765 780 2770 810
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2730 775 2770 780
rect 2180 730 2185 760
rect 2215 730 2220 760
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 685 2060 715
rect 2020 680 2060 685
rect 2030 345 2050 680
rect 2190 675 2210 730
rect 2465 720 2485 770
rect 2630 760 2650 775
rect 2620 730 2625 760
rect 2655 730 2660 760
rect 3110 720 3130 785
rect 3190 760 3230 765
rect 3190 730 3195 760
rect 3225 730 3230 760
rect 3190 725 3230 730
rect 2455 715 2495 720
rect 2455 685 2460 715
rect 2490 685 2495 715
rect 2455 680 2495 685
rect 3100 715 3140 720
rect 3100 685 3105 715
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 2115 670 2155 675
rect 2115 640 2120 670
rect 2150 640 2155 670
rect 2115 635 2155 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 640 2220 670
rect 2180 635 2220 640
rect 2290 670 2330 675
rect 2290 640 2295 670
rect 2325 640 2330 670
rect 2290 635 2330 640
rect 2400 670 2440 675
rect 2400 640 2405 670
rect 2435 640 2440 670
rect 2400 635 2440 640
rect 2510 670 2550 675
rect 2510 640 2515 670
rect 2545 640 2550 670
rect 2510 635 2550 640
rect 2620 670 2660 675
rect 2620 640 2625 670
rect 2655 640 2660 670
rect 2620 635 2660 640
rect 2730 670 2770 675
rect 2730 640 2735 670
rect 2765 640 2770 670
rect 2730 635 2770 640
rect 2795 670 2835 675
rect 2795 640 2800 670
rect 2830 640 2835 670
rect 2795 635 2835 640
rect 2235 395 2275 400
rect 2235 365 2240 395
rect 2270 365 2275 395
rect 2235 360 2275 365
rect 2345 395 2385 400
rect 2345 365 2350 395
rect 2380 365 2385 395
rect 2345 360 2385 365
rect 2405 390 2435 400
rect 2405 370 2410 390
rect 2430 370 2435 390
rect 2405 360 2435 370
rect 2455 395 2495 400
rect 2455 365 2460 395
rect 2490 365 2495 395
rect 2455 360 2495 365
rect 2565 395 2605 400
rect 2565 365 2570 395
rect 2600 365 2605 395
rect 2565 360 2605 365
rect 2675 395 2715 400
rect 2675 365 2680 395
rect 2710 365 2715 395
rect 2675 360 2715 365
rect 2920 395 2960 400
rect 2920 365 2925 395
rect 2955 365 2960 395
rect 2920 360 2960 365
rect 3200 360 3220 725
rect 2410 345 2430 360
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 310 2060 340
rect 2020 305 2060 310
rect 2400 340 2440 345
rect 2400 310 2405 340
rect 2435 310 2440 340
rect 2400 305 2440 310
rect 2410 290 2430 305
rect 2235 285 2275 290
rect 2235 255 2240 285
rect 2270 255 2275 285
rect 2235 250 2275 255
rect 2345 285 2385 290
rect 2345 255 2350 285
rect 2380 255 2385 285
rect 2345 250 2385 255
rect 2405 280 2435 290
rect 2405 260 2410 280
rect 2430 260 2435 280
rect 2405 250 2435 260
rect 2455 285 2495 290
rect 2455 255 2460 285
rect 2490 255 2495 285
rect 2455 250 2495 255
rect 2565 285 2605 290
rect 2565 255 2570 285
rect 2600 255 2605 285
rect 2565 250 2605 255
rect 2675 285 2715 290
rect 2675 255 2680 285
rect 2710 255 2715 285
rect 2675 250 2715 255
rect 2875 285 2915 290
rect 2875 255 2880 285
rect 2910 255 2915 285
rect 2875 250 2915 255
rect 2885 -85 2905 250
rect 2115 -95 2155 -85
rect 2115 -115 2125 -95
rect 2145 -115 2155 -95
rect 2115 -125 2155 -115
rect 2180 -90 2220 -85
rect 2180 -120 2185 -90
rect 2215 -120 2220 -90
rect 2180 -125 2220 -120
rect 2290 -90 2330 -85
rect 2290 -120 2295 -90
rect 2325 -120 2330 -90
rect 2290 -125 2330 -120
rect 2400 -90 2440 -85
rect 2400 -120 2405 -90
rect 2435 -120 2440 -90
rect 2400 -125 2440 -120
rect 2510 -90 2550 -85
rect 2510 -120 2515 -90
rect 2545 -120 2550 -90
rect 2510 -125 2550 -120
rect 2620 -90 2660 -85
rect 2620 -120 2625 -90
rect 2655 -120 2660 -90
rect 2620 -125 2660 -120
rect 2730 -90 2770 -85
rect 2730 -120 2735 -90
rect 2765 -120 2770 -90
rect 2730 -125 2770 -120
rect 2795 -95 2835 -85
rect 2795 -115 2805 -95
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -120 2915 -90
rect 2875 -125 2915 -120
rect 2125 -140 2145 -125
rect 2805 -140 2825 -125
rect 2930 -140 2950 360
rect 3185 350 3235 360
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2965 -120 2969 -85
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3120 -85
rect 3145 -120 3149 -85
rect 3176 -120 3180 -85
rect 2115 -145 2155 -140
rect 2115 -175 2120 -145
rect 2150 -175 2155 -145
rect 2115 -180 2155 -175
rect 2795 -145 2835 -140
rect 2795 -175 2800 -145
rect 2830 -175 2835 -145
rect 2795 -180 2835 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -175 2960 -145
rect 2920 -180 2960 -175
rect 3025 -145 3060 -120
rect 3025 -180 3060 -175
rect 3150 -185 3175 -120
rect 3145 -190 3180 -185
rect 1975 -220 1980 -190
rect 2010 -220 2015 -190
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect 2275 -245 2315 -240
rect 2275 -275 2280 -245
rect 2310 -275 2315 -245
rect 2275 -280 2315 -275
rect 2865 -245 2900 -240
rect 2865 -280 2900 -275
rect 2285 -295 2305 -280
rect 2175 -300 2215 -295
rect 1940 -310 1980 -305
rect 1940 -340 1945 -310
rect 1975 -340 1980 -310
rect 2175 -330 2180 -300
rect 2210 -330 2215 -300
rect 2175 -335 2215 -330
rect 2275 -305 2315 -295
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -335 2315 -325
rect 2375 -300 2415 -295
rect 2375 -330 2380 -300
rect 2410 -330 2415 -300
rect 2375 -335 2415 -330
rect 2575 -300 2615 -295
rect 2575 -330 2580 -300
rect 2610 -330 2615 -300
rect 2575 -335 2615 -330
rect 2805 -300 2840 -295
rect 2805 -335 2840 -330
rect 1940 -345 1980 -340
rect 1885 -355 1925 -350
rect 1885 -385 1890 -355
rect 1920 -385 1925 -355
rect 1885 -390 1925 -385
rect 1335 -425 1375 -420
rect 1335 -455 1340 -425
rect 1370 -455 1375 -425
rect 1335 -460 1375 -455
rect 1840 -425 1880 -420
rect 1840 -455 1845 -425
rect 1875 -455 1880 -425
rect 1840 -460 1880 -455
rect 1345 -475 1365 -460
rect 190 -480 230 -475
rect 190 -510 195 -480
rect 225 -510 230 -480
rect 190 -515 230 -510
rect 385 -480 425 -475
rect 385 -510 390 -480
rect 420 -510 425 -480
rect 385 -515 425 -510
rect 445 -485 475 -475
rect 445 -505 450 -485
rect 470 -505 475 -485
rect 445 -515 475 -505
rect 495 -480 535 -475
rect 495 -510 500 -480
rect 530 -510 535 -480
rect 495 -515 535 -510
rect 605 -480 645 -475
rect 605 -510 610 -480
rect 640 -510 645 -480
rect 605 -515 645 -510
rect 715 -480 755 -475
rect 715 -510 720 -480
rect 750 -510 755 -480
rect 715 -515 755 -510
rect 825 -480 865 -475
rect 825 -510 830 -480
rect 860 -510 865 -480
rect 825 -515 865 -510
rect 935 -480 975 -475
rect 935 -510 940 -480
rect 970 -510 975 -480
rect 935 -515 975 -510
rect 1045 -480 1085 -475
rect 1045 -510 1050 -480
rect 1080 -510 1085 -480
rect 1045 -515 1085 -510
rect 1155 -480 1195 -475
rect 1155 -510 1160 -480
rect 1190 -510 1195 -480
rect 1155 -515 1195 -510
rect 1265 -480 1305 -475
rect 1265 -510 1270 -480
rect 1300 -510 1305 -480
rect 1265 -515 1305 -510
rect 1341 -485 1371 -475
rect 1341 -505 1346 -485
rect 1366 -505 1371 -485
rect 1341 -515 1371 -505
rect 1390 -480 1430 -475
rect 1390 -510 1395 -480
rect 1425 -510 1430 -480
rect 1390 -515 1430 -510
rect 200 -850 220 -515
rect 1940 -800 1960 -345
rect 2810 -380 2835 -335
rect 2870 -380 2895 -280
rect 3200 -295 3220 310
rect 3190 -300 3230 -295
rect 3190 -330 3195 -300
rect 3225 -330 3230 -300
rect 3190 -335 3230 -330
rect 2805 -415 2809 -380
rect 2836 -415 2840 -380
rect 2865 -415 2869 -380
rect 2896 -415 2900 -380
rect 265 -805 305 -800
rect 265 -835 270 -805
rect 300 -835 305 -805
rect 265 -840 305 -835
rect 330 -805 370 -800
rect 330 -835 335 -805
rect 365 -835 370 -805
rect 330 -840 370 -835
rect 440 -805 480 -800
rect 440 -835 445 -805
rect 475 -835 480 -805
rect 440 -840 480 -835
rect 550 -805 590 -800
rect 550 -835 555 -805
rect 585 -835 590 -805
rect 550 -840 590 -835
rect 660 -805 700 -800
rect 660 -835 665 -805
rect 695 -835 700 -805
rect 660 -840 700 -835
rect 770 -805 810 -800
rect 770 -835 775 -805
rect 805 -835 810 -805
rect 770 -840 810 -835
rect 880 -805 920 -800
rect 880 -835 885 -805
rect 915 -835 920 -805
rect 880 -840 920 -835
rect 990 -805 1030 -800
rect 990 -835 995 -805
rect 1025 -835 1030 -805
rect 990 -840 1030 -835
rect 1100 -805 1140 -800
rect 1100 -835 1105 -805
rect 1135 -835 1140 -805
rect 1100 -840 1140 -835
rect 1210 -805 1250 -800
rect 1210 -835 1215 -805
rect 1245 -835 1250 -805
rect 1210 -840 1250 -835
rect 1320 -805 1360 -800
rect 1320 -835 1325 -805
rect 1355 -835 1360 -805
rect 1320 -840 1360 -835
rect 1430 -805 1470 -800
rect 1430 -835 1435 -805
rect 1465 -835 1470 -805
rect 1430 -840 1470 -835
rect 1930 -805 1970 -800
rect 1930 -835 1935 -805
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect 190 -855 230 -850
rect 190 -885 195 -855
rect 225 -885 230 -855
rect 190 -890 230 -885
rect 1315 -865 1355 -860
rect 1315 -895 1320 -865
rect 1350 -895 1355 -865
rect -190 -900 -150 -895
rect -190 -930 -185 -900
rect -155 -930 -150 -900
rect -190 -935 -150 -930
rect 550 -900 590 -895
rect 550 -930 555 -900
rect 585 -930 590 -900
rect 550 -935 590 -930
rect 660 -900 700 -895
rect 660 -930 665 -900
rect 695 -930 700 -900
rect 660 -935 700 -930
rect 770 -900 810 -895
rect 770 -930 775 -900
rect 805 -930 810 -900
rect 770 -935 810 -930
rect 1005 -900 1045 -895
rect 1005 -930 1010 -900
rect 1040 -930 1045 -900
rect 1005 -935 1045 -930
rect 1125 -900 1165 -895
rect 1125 -930 1130 -900
rect 1160 -930 1165 -900
rect 1125 -935 1165 -930
rect 1255 -900 1295 -895
rect 1315 -900 1355 -895
rect 1255 -930 1260 -900
rect 1290 -930 1295 -900
rect 1255 -935 1295 -930
rect 925 -1010 965 -1005
rect 925 -1040 930 -1010
rect 960 -1040 965 -1010
rect 925 -1045 965 -1040
rect 935 -1115 955 -1045
rect 500 -1125 530 -1115
rect 500 -1145 505 -1125
rect 525 -1145 530 -1125
rect 500 -1155 530 -1145
rect 605 -1120 645 -1115
rect 605 -1150 610 -1120
rect 640 -1150 645 -1120
rect 605 -1155 645 -1150
rect 715 -1120 755 -1115
rect 715 -1150 720 -1120
rect 750 -1150 755 -1120
rect 715 -1155 755 -1150
rect 830 -1125 860 -1115
rect 830 -1145 835 -1125
rect 855 -1145 860 -1125
rect 830 -1155 860 -1145
rect 925 -1120 965 -1115
rect 925 -1150 930 -1120
rect 960 -1150 965 -1120
rect 925 -1155 965 -1150
rect 505 -1170 525 -1155
rect 835 -1170 855 -1155
rect 1940 -1170 1960 -840
rect 2075 -1075 2115 -1070
rect 2075 -1105 2080 -1075
rect 2110 -1105 2115 -1075
rect 2075 -1110 2115 -1105
rect 2275 -1075 2315 -1070
rect 2275 -1105 2280 -1075
rect 2310 -1105 2315 -1075
rect 2275 -1110 2315 -1105
rect 2375 -1075 2415 -1070
rect 2375 -1105 2380 -1075
rect 2410 -1105 2415 -1075
rect 2375 -1110 2415 -1105
rect 2475 -1075 2515 -1070
rect 2475 -1105 2480 -1075
rect 2510 -1105 2515 -1075
rect 2475 -1110 2515 -1105
rect 2675 -1075 2715 -1070
rect 2675 -1105 2680 -1075
rect 2710 -1105 2715 -1075
rect 2675 -1110 2715 -1105
rect 2385 -1170 2405 -1110
rect -725 -1175 -685 -1170
rect -725 -1205 -720 -1175
rect -690 -1205 -685 -1175
rect -725 -1210 -685 -1205
rect -280 -1175 -240 -1170
rect -280 -1205 -275 -1175
rect -245 -1205 -240 -1175
rect -280 -1210 -240 -1205
rect 495 -1175 535 -1170
rect 495 -1205 500 -1175
rect 530 -1205 535 -1175
rect 495 -1210 535 -1205
rect 825 -1175 865 -1170
rect 825 -1205 830 -1175
rect 860 -1205 865 -1175
rect 825 -1210 865 -1205
rect 1930 -1175 1970 -1170
rect 1930 -1205 1935 -1175
rect 1965 -1205 1970 -1175
rect 1930 -1210 1970 -1205
rect 2375 -1175 2415 -1170
rect 2375 -1205 2380 -1175
rect 2410 -1205 2415 -1175
rect 2375 -1210 2415 -1205
rect 835 -2420 855 -1210
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via1 >>
rect 830 4245 860 4275
rect 155 2750 185 2780
rect 625 2750 655 2780
rect 35 2720 65 2725
rect 35 2700 40 2720
rect 40 2700 60 2720
rect 60 2700 65 2720
rect 35 2695 65 2700
rect 155 2720 185 2725
rect 155 2700 160 2720
rect 160 2700 180 2720
rect 180 2700 185 2720
rect 155 2695 185 2700
rect 215 2720 245 2725
rect 215 2700 220 2720
rect 220 2700 240 2720
rect 240 2700 245 2720
rect 215 2695 245 2700
rect 1035 2750 1065 2780
rect 1503 2750 1533 2780
rect 830 2695 860 2725
rect 975 2720 1005 2725
rect 975 2700 980 2720
rect 980 2700 1000 2720
rect 1000 2700 1005 2720
rect 975 2695 1005 2700
rect 1095 2720 1125 2725
rect 1095 2700 1100 2720
rect 1100 2700 1120 2720
rect 1120 2700 1125 2720
rect 1095 2695 1125 2700
rect 1155 2720 1185 2725
rect 1155 2700 1160 2720
rect 1160 2700 1180 2720
rect 1180 2700 1185 2720
rect 1155 2695 1185 2700
rect 1443 2720 1473 2725
rect 1443 2700 1448 2720
rect 1448 2700 1468 2720
rect 1468 2700 1473 2720
rect 1443 2695 1473 2700
rect 1503 2720 1533 2725
rect 1503 2700 1508 2720
rect 1508 2700 1528 2720
rect 1528 2700 1533 2720
rect 1503 2695 1533 2700
rect 1623 2720 1653 2725
rect 1623 2700 1628 2720
rect 1628 2700 1648 2720
rect 1648 2700 1653 2720
rect 1623 2695 1653 2700
rect 505 2550 535 2555
rect 505 2530 510 2550
rect 510 2530 530 2550
rect 530 2530 535 2550
rect 505 2525 535 2530
rect 565 2550 595 2555
rect 565 2530 570 2550
rect 570 2530 590 2550
rect 590 2530 595 2550
rect 565 2525 595 2530
rect 685 2550 715 2555
rect 685 2530 690 2550
rect 690 2530 710 2550
rect 710 2530 715 2550
rect 685 2525 715 2530
rect 830 2525 860 2555
rect 80 2300 110 2305
rect 80 2280 85 2300
rect 85 2280 105 2300
rect 105 2280 110 2300
rect 80 2275 110 2280
rect 139 2300 169 2305
rect 139 2280 144 2300
rect 144 2280 164 2300
rect 164 2280 169 2300
rect 139 2275 169 2280
rect 609 2300 639 2305
rect 609 2280 614 2300
rect 614 2280 634 2300
rect 634 2280 639 2300
rect 609 2275 639 2280
rect 775 2275 805 2305
rect -800 2175 -770 2205
rect -230 2175 -200 2205
rect -1160 2145 -1130 2150
rect -1160 2125 -1155 2145
rect -1155 2125 -1135 2145
rect -1135 2125 -1130 2145
rect -1160 2120 -1130 2125
rect -1040 2145 -1010 2150
rect -1040 2125 -1035 2145
rect -1035 2125 -1015 2145
rect -1015 2125 -1010 2145
rect -1040 2120 -1010 2125
rect -920 2145 -890 2150
rect -920 2125 -915 2145
rect -915 2125 -895 2145
rect -895 2125 -890 2145
rect -920 2120 -890 2125
rect -800 2145 -770 2150
rect -800 2125 -795 2145
rect -795 2125 -775 2145
rect -775 2125 -770 2145
rect -800 2120 -770 2125
rect -680 2145 -650 2150
rect -680 2125 -675 2145
rect -675 2125 -655 2145
rect -655 2125 -650 2145
rect -680 2120 -650 2125
rect -560 2145 -530 2150
rect -560 2125 -555 2145
rect -555 2125 -535 2145
rect -535 2125 -530 2145
rect -560 2120 -530 2125
rect -440 2145 -410 2150
rect -440 2125 -435 2145
rect -435 2125 -415 2145
rect -415 2125 -410 2145
rect -440 2120 -410 2125
rect -275 2120 -245 2150
rect -1100 1720 -1070 1725
rect -1100 1700 -1095 1720
rect -1095 1700 -1075 1720
rect -1075 1700 -1070 1720
rect -1100 1695 -1070 1700
rect -980 1720 -950 1725
rect -980 1700 -975 1720
rect -975 1700 -955 1720
rect -955 1700 -950 1720
rect -980 1695 -950 1700
rect -860 1720 -830 1725
rect -860 1700 -855 1720
rect -855 1700 -835 1720
rect -835 1700 -830 1720
rect -860 1695 -830 1700
rect -740 1720 -710 1725
rect -740 1700 -735 1720
rect -735 1700 -715 1720
rect -715 1700 -710 1720
rect -740 1695 -710 1700
rect -620 1720 -590 1725
rect -620 1700 -615 1720
rect -615 1700 -595 1720
rect -595 1700 -590 1720
rect -620 1695 -590 1700
rect -500 1720 -470 1725
rect -500 1700 -495 1720
rect -495 1700 -475 1720
rect -475 1700 -470 1720
rect -500 1695 -470 1700
rect -275 1695 -245 1725
rect -365 1640 -335 1670
rect -800 1595 -770 1625
rect -1445 1510 -1415 1540
rect -1130 1480 -1100 1485
rect -1130 1460 -1125 1480
rect -1125 1460 -1105 1480
rect -1105 1460 -1100 1480
rect -1130 1455 -1100 1460
rect -1020 1480 -990 1485
rect -1020 1460 -1015 1480
rect -1015 1460 -995 1480
rect -995 1460 -990 1480
rect -1020 1455 -990 1460
rect -910 1480 -880 1485
rect -910 1460 -905 1480
rect -905 1460 -885 1480
rect -885 1460 -880 1480
rect -910 1455 -880 1460
rect -800 1480 -770 1485
rect -800 1460 -795 1480
rect -795 1460 -775 1480
rect -775 1460 -770 1480
rect -800 1455 -770 1460
rect -690 1480 -660 1485
rect -690 1460 -685 1480
rect -685 1460 -665 1480
rect -665 1460 -660 1480
rect -690 1455 -660 1460
rect -580 1480 -550 1485
rect -580 1460 -575 1480
rect -575 1460 -555 1480
rect -555 1460 -550 1480
rect -580 1455 -550 1460
rect -470 1480 -440 1485
rect -470 1460 -465 1480
rect -465 1460 -445 1480
rect -445 1460 -440 1480
rect -470 1455 -440 1460
rect -35 2145 -5 2150
rect -35 2125 -30 2145
rect -30 2125 -10 2145
rect -10 2125 -5 2145
rect -35 2120 -5 2125
rect 85 2145 115 2150
rect 85 2125 90 2145
rect 90 2125 110 2145
rect 110 2125 115 2145
rect 85 2120 115 2125
rect 205 2145 235 2150
rect 205 2125 210 2145
rect 210 2125 230 2145
rect 230 2125 235 2145
rect 205 2120 235 2125
rect 325 2145 355 2150
rect 325 2125 330 2145
rect 330 2125 350 2145
rect 350 2125 355 2145
rect 325 2120 355 2125
rect 445 2145 475 2150
rect 445 2125 450 2145
rect 450 2125 470 2145
rect 470 2125 475 2145
rect 445 2120 475 2125
rect 565 2145 595 2150
rect 565 2125 570 2145
rect 570 2125 590 2145
rect 590 2125 595 2145
rect 565 2120 595 2125
rect 685 2145 715 2150
rect 685 2125 690 2145
rect 690 2125 710 2145
rect 710 2125 715 2145
rect 685 2120 715 2125
rect 25 1720 55 1725
rect 25 1700 30 1720
rect 30 1700 50 1720
rect 50 1700 55 1720
rect 25 1695 55 1700
rect 145 1720 175 1725
rect 145 1700 150 1720
rect 150 1700 170 1720
rect 170 1700 175 1720
rect 145 1695 175 1700
rect 265 1720 295 1725
rect 265 1700 270 1720
rect 270 1700 290 1720
rect 290 1700 295 1720
rect 265 1695 295 1700
rect 385 1720 415 1725
rect 385 1700 390 1720
rect 390 1700 410 1720
rect 410 1700 415 1720
rect 385 1695 415 1700
rect 505 1720 535 1725
rect 505 1700 510 1720
rect 510 1700 530 1720
rect 530 1700 535 1720
rect 505 1695 535 1700
rect 625 1720 655 1725
rect 625 1700 630 1720
rect 630 1700 650 1720
rect 650 1700 655 1720
rect 625 1695 655 1700
rect 1519 2300 1549 2305
rect 1519 2280 1524 2300
rect 1524 2280 1544 2300
rect 1544 2280 1549 2300
rect 1519 2275 1549 2280
rect 885 2230 915 2260
rect 830 2175 860 2205
rect 25 1640 55 1670
rect 325 1640 355 1670
rect 785 1640 815 1670
rect 1050 2220 1080 2250
rect 1578 2220 1608 2250
rect 1890 2175 1920 2205
rect 2460 2175 2490 2205
rect 975 2145 1005 2150
rect 975 2125 980 2145
rect 980 2125 1000 2145
rect 1000 2125 1005 2145
rect 975 2120 1005 2125
rect 1095 2145 1125 2150
rect 1095 2125 1100 2145
rect 1100 2125 1120 2145
rect 1120 2125 1125 2145
rect 1095 2120 1125 2125
rect 1215 2145 1245 2150
rect 1215 2125 1220 2145
rect 1220 2125 1240 2145
rect 1240 2125 1245 2145
rect 1215 2120 1245 2125
rect 1335 2145 1365 2150
rect 1335 2125 1340 2145
rect 1340 2125 1360 2145
rect 1360 2125 1365 2145
rect 1335 2120 1365 2125
rect 1455 2145 1485 2150
rect 1455 2125 1460 2145
rect 1460 2125 1480 2145
rect 1480 2125 1485 2145
rect 1455 2120 1485 2125
rect 1575 2145 1605 2150
rect 1575 2125 1580 2145
rect 1580 2125 1600 2145
rect 1600 2125 1605 2145
rect 1575 2120 1605 2125
rect 1695 2145 1725 2150
rect 1695 2125 1700 2145
rect 1700 2125 1720 2145
rect 1720 2125 1725 2145
rect 1695 2120 1725 2125
rect 1035 1720 1065 1725
rect 1035 1700 1040 1720
rect 1040 1700 1060 1720
rect 1060 1700 1065 1720
rect 1035 1695 1065 1700
rect 1155 1720 1185 1725
rect 1155 1700 1160 1720
rect 1160 1700 1180 1720
rect 1180 1700 1185 1720
rect 1155 1695 1185 1700
rect 1275 1720 1305 1725
rect 1275 1700 1280 1720
rect 1280 1700 1300 1720
rect 1300 1700 1305 1720
rect 1275 1695 1305 1700
rect 1395 1720 1425 1725
rect 1395 1700 1400 1720
rect 1400 1700 1420 1720
rect 1420 1700 1425 1720
rect 1395 1695 1425 1700
rect 1515 1720 1545 1725
rect 1515 1700 1520 1720
rect 1520 1700 1540 1720
rect 1540 1700 1545 1720
rect 1515 1695 1545 1700
rect 1635 1720 1665 1725
rect 1635 1700 1640 1720
rect 1640 1700 1660 1720
rect 1660 1700 1665 1720
rect 1635 1695 1665 1700
rect 1335 1640 1365 1670
rect 1635 1640 1665 1670
rect 875 1600 905 1630
rect 1935 2120 1965 2150
rect 2100 2145 2130 2150
rect 2100 2125 2105 2145
rect 2105 2125 2125 2145
rect 2125 2125 2130 2145
rect 2100 2120 2130 2125
rect 2220 2145 2250 2150
rect 2220 2125 2225 2145
rect 2225 2125 2245 2145
rect 2245 2125 2250 2145
rect 2220 2120 2250 2125
rect 2340 2145 2370 2150
rect 2340 2125 2345 2145
rect 2345 2125 2365 2145
rect 2365 2125 2370 2145
rect 2340 2120 2370 2125
rect 2460 2145 2490 2150
rect 2460 2125 2465 2145
rect 2465 2125 2485 2145
rect 2485 2125 2490 2145
rect 2460 2120 2490 2125
rect 2580 2145 2610 2150
rect 2580 2125 2585 2145
rect 2585 2125 2605 2145
rect 2605 2125 2610 2145
rect 2580 2120 2610 2125
rect 2700 2145 2730 2150
rect 2700 2125 2705 2145
rect 2705 2125 2725 2145
rect 2725 2125 2730 2145
rect 2700 2120 2730 2125
rect 2820 2145 2850 2150
rect 2820 2125 2825 2145
rect 2825 2125 2845 2145
rect 2845 2125 2850 2145
rect 2820 2120 2850 2125
rect 1935 1695 1965 1725
rect 2160 1720 2190 1725
rect 2160 1700 2165 1720
rect 2165 1700 2185 1720
rect 2185 1700 2190 1720
rect 2160 1695 2190 1700
rect 2280 1720 2310 1725
rect 2280 1700 2285 1720
rect 2285 1700 2305 1720
rect 2305 1700 2310 1720
rect 2280 1695 2310 1700
rect 2400 1720 2430 1725
rect 2400 1700 2405 1720
rect 2405 1700 2425 1720
rect 2425 1700 2430 1720
rect 2400 1695 2430 1700
rect 2520 1720 2550 1725
rect 2520 1700 2525 1720
rect 2525 1700 2545 1720
rect 2545 1700 2550 1720
rect 2520 1695 2550 1700
rect 2640 1720 2670 1725
rect 2640 1700 2645 1720
rect 2645 1700 2665 1720
rect 2665 1700 2670 1720
rect 2640 1695 2670 1700
rect 2760 1720 2790 1725
rect 2760 1700 2765 1720
rect 2765 1700 2785 1720
rect 2785 1700 2790 1720
rect 2760 1695 2790 1700
rect 2025 1640 2055 1670
rect 460 1575 490 1580
rect 460 1555 465 1575
rect 465 1555 485 1575
rect 485 1555 490 1575
rect 460 1550 490 1555
rect 625 1575 655 1580
rect 625 1555 630 1575
rect 630 1555 650 1575
rect 650 1555 655 1575
rect 625 1550 655 1555
rect 790 1575 820 1580
rect 790 1555 795 1575
rect 795 1555 815 1575
rect 815 1555 820 1575
rect 790 1550 820 1555
rect 870 1575 900 1580
rect 870 1555 875 1575
rect 875 1555 895 1575
rect 895 1555 900 1575
rect 870 1550 900 1555
rect 1035 1575 1065 1580
rect 1035 1555 1040 1575
rect 1040 1555 1060 1575
rect 1060 1555 1065 1575
rect 1035 1550 1065 1555
rect 1200 1575 1230 1580
rect 1200 1555 1205 1575
rect 1205 1555 1225 1575
rect 1225 1555 1230 1575
rect 1200 1550 1230 1555
rect 1890 1550 1920 1580
rect 570 1530 600 1535
rect 570 1510 575 1530
rect 575 1510 595 1530
rect 595 1510 600 1530
rect 570 1505 600 1510
rect 680 1530 710 1535
rect 680 1510 685 1530
rect 685 1510 705 1530
rect 705 1510 710 1530
rect 680 1505 710 1510
rect 980 1530 1010 1535
rect 980 1510 985 1530
rect 985 1510 1005 1530
rect 1005 1510 1010 1530
rect 980 1505 1010 1510
rect 1090 1530 1120 1535
rect 1090 1510 1095 1530
rect 1095 1510 1115 1530
rect 1115 1510 1120 1530
rect 1090 1505 1120 1510
rect -230 1455 -200 1485
rect 1890 1455 1920 1485
rect -320 1075 -290 1105
rect -365 930 -335 960
rect -1535 730 -1505 760
rect -1075 805 -1045 810
rect -1075 785 -1070 805
rect -1070 785 -1050 805
rect -1050 785 -1045 805
rect -1075 780 -1045 785
rect -965 805 -935 810
rect -965 785 -960 805
rect -960 785 -940 805
rect -940 785 -935 805
rect -965 780 -935 785
rect -855 805 -825 810
rect -855 785 -850 805
rect -850 785 -830 805
rect -830 785 -825 805
rect -855 780 -825 785
rect -745 805 -715 810
rect -745 785 -740 805
rect -740 785 -720 805
rect -720 785 -715 805
rect -745 780 -715 785
rect -635 805 -605 810
rect -635 785 -630 805
rect -630 785 -610 805
rect -610 785 -605 805
rect -635 780 -605 785
rect -525 805 -495 810
rect -525 785 -520 805
rect -520 785 -500 805
rect -500 785 -495 805
rect -525 780 -495 785
rect -965 730 -935 760
rect -525 730 -495 760
rect -1445 685 -1415 715
rect -800 685 -770 715
rect -365 685 -335 715
rect -1140 665 -1110 670
rect -1140 645 -1135 665
rect -1135 645 -1115 665
rect -1115 645 -1110 665
rect -1140 640 -1110 645
rect -1075 665 -1045 670
rect -1075 645 -1070 665
rect -1070 645 -1050 665
rect -1050 645 -1045 665
rect -1075 640 -1045 645
rect -965 665 -935 670
rect -965 645 -960 665
rect -960 645 -940 665
rect -940 645 -935 665
rect -965 640 -935 645
rect -855 665 -825 670
rect -855 645 -850 665
rect -850 645 -830 665
rect -830 645 -825 665
rect -855 640 -825 645
rect -745 665 -715 670
rect -745 645 -740 665
rect -740 645 -720 665
rect -720 645 -715 665
rect -745 640 -715 645
rect -635 665 -605 670
rect -635 645 -630 665
rect -630 645 -610 665
rect -610 645 -605 665
rect -635 640 -605 645
rect -525 665 -495 670
rect -525 645 -520 665
rect -520 645 -500 665
rect -500 645 -495 665
rect -525 640 -495 645
rect -460 665 -430 670
rect -460 645 -455 665
rect -455 645 -435 665
rect -435 645 -430 665
rect -460 640 -430 645
rect -1265 365 -1235 395
rect -1020 390 -990 395
rect -1020 370 -1015 390
rect -1015 370 -995 390
rect -995 370 -990 390
rect -1020 365 -990 370
rect -910 390 -880 395
rect -910 370 -905 390
rect -905 370 -885 390
rect -885 370 -880 390
rect -910 365 -880 370
rect -800 390 -770 395
rect -800 370 -795 390
rect -795 370 -775 390
rect -775 370 -770 390
rect -800 365 -770 370
rect -690 390 -660 395
rect -690 370 -685 390
rect -685 370 -665 390
rect -665 370 -660 390
rect -690 365 -660 370
rect -580 390 -550 395
rect -580 370 -575 390
rect -575 370 -555 390
rect -555 370 -550 390
rect -580 365 -550 370
rect -1535 320 -1505 350
rect -1486 -93 -1459 -85
rect -1486 -113 -1485 -93
rect -1485 -113 -1460 -93
rect -1460 -113 -1459 -93
rect -1486 -120 -1459 -113
rect -1426 -93 -1399 -85
rect -1426 -113 -1425 -93
rect -1425 -113 -1400 -93
rect -1400 -113 -1399 -93
rect -1426 -120 -1399 -113
rect -1366 -93 -1339 -85
rect -1366 -113 -1365 -93
rect -1365 -113 -1340 -93
rect -1340 -113 -1339 -93
rect -1366 -120 -1339 -113
rect -1306 -93 -1279 -85
rect -1306 -113 -1305 -93
rect -1305 -113 -1280 -93
rect -1280 -113 -1279 -93
rect -1306 -120 -1279 -113
rect -745 310 -715 340
rect -365 310 -335 340
rect -1220 255 -1190 285
rect -1020 280 -990 285
rect -1020 260 -1015 280
rect -1015 260 -995 280
rect -995 260 -990 280
rect -1020 255 -990 260
rect -910 280 -880 285
rect -910 260 -905 280
rect -905 260 -885 280
rect -885 260 -880 280
rect -910 255 -880 260
rect -800 280 -770 285
rect -800 260 -795 280
rect -795 260 -775 280
rect -775 260 -770 280
rect -800 255 -770 260
rect -690 280 -660 285
rect -690 260 -685 280
rect -685 260 -665 280
rect -665 260 -660 280
rect -690 255 -660 260
rect -580 280 -550 285
rect -580 260 -575 280
rect -575 260 -555 280
rect -555 260 -550 280
rect -580 255 -550 260
rect -1220 -120 -1190 -90
rect -1075 -95 -1045 -90
rect -1075 -115 -1070 -95
rect -1070 -115 -1050 -95
rect -1050 -115 -1045 -95
rect -1075 -120 -1045 -115
rect -965 -95 -935 -90
rect -965 -115 -960 -95
rect -960 -115 -940 -95
rect -940 -115 -935 -95
rect -965 -120 -935 -115
rect -855 -95 -825 -90
rect -855 -115 -850 -95
rect -850 -115 -830 -95
rect -830 -115 -825 -95
rect -855 -120 -825 -115
rect -745 -95 -715 -90
rect -745 -115 -740 -95
rect -740 -115 -720 -95
rect -720 -115 -715 -95
rect -745 -120 -715 -115
rect -635 -95 -605 -90
rect -635 -115 -630 -95
rect -630 -115 -610 -95
rect -610 -115 -605 -95
rect -635 -120 -605 -115
rect -525 -95 -495 -90
rect -525 -115 -520 -95
rect -520 -115 -500 -95
rect -500 -115 -495 -95
rect -525 -120 -495 -115
rect -1370 -175 -1335 -145
rect -1265 -175 -1235 -145
rect -1140 -175 -1110 -145
rect -460 -175 -430 -145
rect -275 740 -245 770
rect 505 1220 535 1225
rect 745 1220 775 1225
rect 505 1200 510 1220
rect 510 1200 530 1220
rect 530 1200 535 1220
rect 505 1195 535 1200
rect 625 1210 655 1215
rect 625 1190 630 1210
rect 630 1190 650 1210
rect 650 1190 655 1210
rect 625 1185 655 1190
rect 745 1200 750 1220
rect 750 1200 770 1220
rect 770 1200 775 1220
rect 745 1195 775 1200
rect 550 1150 580 1155
rect 550 1130 555 1150
rect 555 1130 575 1150
rect 575 1130 580 1150
rect 550 1125 580 1130
rect 695 1075 725 1105
rect 1035 1210 1065 1215
rect 1035 1190 1040 1210
rect 1040 1190 1060 1210
rect 1060 1190 1065 1210
rect 1035 1185 1065 1190
rect 1110 1150 1140 1155
rect 1110 1130 1115 1150
rect 1115 1130 1135 1150
rect 1135 1130 1140 1150
rect 1110 1125 1140 1130
rect 965 1075 995 1105
rect 800 1030 830 1060
rect 910 1030 940 1060
rect 800 975 830 1005
rect 885 975 915 1005
rect 1160 985 1190 1015
rect 1845 975 1875 1005
rect -45 930 -15 960
rect 65 930 95 960
rect 175 930 205 960
rect 285 930 315 960
rect 395 930 425 960
rect 505 930 535 960
rect 1155 930 1185 960
rect -175 875 -145 905
rect 230 900 260 905
rect 230 880 235 900
rect 235 880 255 900
rect 255 880 260 900
rect 230 875 260 880
rect 1265 930 1295 960
rect 1375 930 1405 960
rect 1485 930 1515 960
rect 1595 930 1625 960
rect 1705 930 1735 960
rect 1430 900 1460 905
rect 1430 880 1435 900
rect 1435 880 1455 900
rect 1455 880 1460 900
rect 1430 875 1460 880
rect -230 640 -200 670
rect -230 -120 -200 -90
rect -275 -175 -245 -145
rect -1490 -220 -1455 -190
rect -320 -220 -290 -190
rect -1210 -275 -1175 -245
rect -620 -275 -590 -245
rect -1535 -330 -1505 -300
rect -1150 -330 -1115 -300
rect -920 -305 -890 -300
rect -920 -325 -915 -305
rect -915 -325 -895 -305
rect -895 -325 -890 -305
rect -920 -330 -890 -325
rect -720 -305 -690 -300
rect -720 -325 -715 -305
rect -715 -325 -695 -305
rect -695 -325 -690 -305
rect -720 -330 -690 -325
rect -520 -305 -490 -300
rect -520 -325 -515 -305
rect -515 -325 -495 -305
rect -495 -325 -490 -305
rect -520 -330 -490 -325
rect -1206 -387 -1179 -380
rect -1206 -407 -1205 -387
rect -1205 -407 -1180 -387
rect -1180 -407 -1179 -387
rect -1206 -415 -1179 -407
rect -1146 -387 -1119 -380
rect -1146 -407 -1145 -387
rect -1145 -407 -1120 -387
rect -1120 -407 -1119 -387
rect -1146 -415 -1119 -407
rect -1020 -1080 -990 -1075
rect -1020 -1100 -1015 -1080
rect -1015 -1100 -995 -1080
rect -995 -1100 -990 -1080
rect -1020 -1105 -990 -1100
rect -820 -1080 -790 -1075
rect -820 -1100 -815 -1080
rect -815 -1100 -795 -1080
rect -795 -1100 -790 -1080
rect -820 -1105 -790 -1100
rect -720 -1105 -690 -1075
rect -620 -1080 -590 -1075
rect -620 -1100 -615 -1080
rect -615 -1100 -595 -1080
rect -595 -1100 -590 -1080
rect -620 -1105 -590 -1100
rect -420 -1080 -390 -1075
rect -420 -1100 -415 -1080
rect -415 -1100 -395 -1080
rect -395 -1100 -390 -1080
rect -420 -1105 -390 -1100
rect -230 -275 -200 -245
rect -230 -385 -200 -355
rect 10 675 40 680
rect 10 655 15 675
rect 15 655 35 675
rect 35 655 40 675
rect 10 650 40 655
rect 120 675 150 680
rect 120 655 125 675
rect 125 655 145 675
rect 145 655 150 675
rect 120 650 150 655
rect 230 675 260 680
rect 230 655 235 675
rect 235 655 255 675
rect 255 655 260 675
rect 230 650 260 655
rect 340 675 370 680
rect 340 655 345 675
rect 345 655 365 675
rect 365 655 370 675
rect 340 650 370 655
rect 450 675 480 680
rect 450 655 455 675
rect 455 655 475 675
rect 475 655 480 675
rect 450 650 480 655
rect 1210 675 1240 680
rect 1210 655 1215 675
rect 1215 655 1235 675
rect 1235 655 1240 675
rect 1210 650 1240 655
rect 1320 675 1350 680
rect 1320 655 1325 675
rect 1325 655 1345 675
rect 1345 655 1350 675
rect 1320 650 1350 655
rect 1430 675 1460 680
rect 1430 655 1435 675
rect 1435 655 1455 675
rect 1455 655 1460 675
rect 1430 650 1460 655
rect 1540 675 1570 680
rect 1540 655 1545 675
rect 1545 655 1565 675
rect 1565 655 1570 675
rect 1540 650 1570 655
rect 1650 675 1680 680
rect 1650 655 1655 675
rect 1655 655 1675 675
rect 1675 655 1680 675
rect 1650 650 1680 655
rect -100 595 -70 625
rect 560 595 590 625
rect 720 600 750 605
rect 720 580 725 600
rect 725 580 745 600
rect 745 580 750 600
rect 720 575 750 580
rect 830 600 860 605
rect 830 580 835 600
rect 835 580 855 600
rect 855 580 860 600
rect 830 575 860 580
rect 940 600 970 605
rect 940 580 945 600
rect 945 580 965 600
rect 965 580 970 600
rect 940 575 970 580
rect 1100 595 1130 625
rect 1760 595 1790 625
rect -45 550 -15 555
rect -45 530 -40 550
rect -40 530 -20 550
rect -20 530 -15 550
rect -45 525 -15 530
rect 65 550 95 555
rect 65 530 70 550
rect 70 530 90 550
rect 90 530 95 550
rect 65 525 95 530
rect 175 550 205 555
rect 175 530 180 550
rect 180 530 200 550
rect 200 530 205 550
rect 175 525 205 530
rect 230 535 260 565
rect 285 550 315 555
rect 285 530 290 550
rect 290 530 310 550
rect 310 530 315 550
rect 285 525 315 530
rect 395 550 425 555
rect 395 530 400 550
rect 400 530 420 550
rect 420 530 425 550
rect 395 525 425 530
rect 505 550 535 555
rect 505 530 510 550
rect 510 530 530 550
rect 530 530 535 550
rect 505 525 535 530
rect 1155 550 1185 555
rect 1155 530 1160 550
rect 1160 530 1180 550
rect 1180 530 1185 550
rect 1155 525 1185 530
rect 1265 550 1295 555
rect 1265 530 1270 550
rect 1270 530 1290 550
rect 1290 530 1295 550
rect 1265 525 1295 530
rect 1375 550 1405 555
rect 1375 530 1380 550
rect 1380 530 1400 550
rect 1400 530 1405 550
rect 1375 525 1405 530
rect 1430 535 1460 565
rect 1485 550 1515 555
rect 1485 530 1490 550
rect 1490 530 1510 550
rect 1510 530 1515 550
rect 1485 525 1515 530
rect 1595 550 1625 555
rect 1595 530 1600 550
rect 1600 530 1620 550
rect 1620 530 1625 550
rect 1595 525 1625 530
rect 1705 550 1735 555
rect 1705 530 1710 550
rect 1710 530 1730 550
rect 1730 530 1735 550
rect 1705 525 1735 530
rect 230 500 260 505
rect 230 480 235 500
rect 235 480 255 500
rect 255 480 260 500
rect 230 475 260 480
rect 795 500 825 505
rect 795 480 800 500
rect 800 480 820 500
rect 820 480 825 500
rect 795 475 825 480
rect 865 500 895 505
rect 865 480 870 500
rect 870 480 890 500
rect 890 480 895 500
rect 865 475 895 480
rect 1430 500 1460 505
rect 1430 480 1435 500
rect 1435 480 1455 500
rect 1455 480 1460 500
rect 1430 475 1460 480
rect 10 280 40 285
rect 10 260 15 280
rect 15 260 35 280
rect 35 260 40 280
rect 10 255 40 260
rect 120 280 150 285
rect 120 260 125 280
rect 125 260 145 280
rect 145 260 150 280
rect 120 255 150 260
rect 230 280 260 285
rect 230 260 235 280
rect 235 260 255 280
rect 255 260 260 280
rect 230 255 260 260
rect 340 280 370 285
rect 340 260 345 280
rect 345 260 365 280
rect 365 260 370 280
rect 340 255 370 260
rect 450 280 480 285
rect 450 260 455 280
rect 455 260 475 280
rect 475 260 480 280
rect 450 255 480 260
rect 1210 280 1240 285
rect 1210 260 1215 280
rect 1215 260 1235 280
rect 1235 260 1240 280
rect 1210 255 1240 260
rect 1265 255 1295 285
rect 1320 280 1350 285
rect 1320 260 1325 280
rect 1325 260 1345 280
rect 1345 260 1350 280
rect 1320 255 1350 260
rect 1430 280 1460 285
rect 1430 260 1435 280
rect 1435 260 1455 280
rect 1455 260 1460 280
rect 1430 255 1460 260
rect 1540 280 1570 285
rect 1540 260 1545 280
rect 1545 260 1565 280
rect 1565 260 1570 280
rect 1540 255 1570 260
rect 1650 280 1680 285
rect 1650 260 1655 280
rect 1655 260 1675 280
rect 1675 260 1680 280
rect 1650 255 1680 260
rect 445 -15 475 15
rect -100 -340 -70 -310
rect 785 200 815 230
rect 875 200 905 230
rect 860 145 890 175
rect 800 90 830 120
rect 785 35 815 65
rect 875 35 905 65
rect 830 10 860 15
rect 830 -10 835 10
rect 835 -10 855 10
rect 855 -10 860 10
rect 830 -15 860 -10
rect 600 -340 630 -310
rect 720 -315 750 -310
rect 720 -335 725 -315
rect 725 -335 745 -315
rect 745 -335 750 -315
rect 720 -340 750 -335
rect 830 -315 860 -310
rect 830 -335 835 -315
rect 835 -335 855 -315
rect 855 -335 860 -315
rect 830 -340 860 -335
rect 940 -315 970 -310
rect 940 -335 945 -315
rect 945 -335 965 -315
rect 965 -335 970 -315
rect 940 -340 970 -335
rect 1070 -340 1100 -310
rect 1755 -340 1785 -310
rect 1980 1075 2010 1105
rect 1935 740 1965 770
rect 1890 640 1920 670
rect 1935 585 1965 615
rect 1890 -120 1920 -90
rect 1935 -175 1965 -145
rect 1890 -275 1920 -245
rect 2460 1595 2490 1625
rect 2130 1480 2160 1485
rect 2130 1460 2135 1480
rect 2135 1460 2155 1480
rect 2155 1460 2160 1480
rect 2130 1455 2160 1460
rect 2240 1480 2270 1485
rect 2240 1460 2245 1480
rect 2245 1460 2265 1480
rect 2265 1460 2270 1480
rect 2240 1455 2270 1460
rect 2350 1480 2380 1485
rect 2350 1460 2355 1480
rect 2355 1460 2375 1480
rect 2375 1460 2380 1480
rect 2350 1455 2380 1460
rect 2460 1480 2490 1485
rect 2460 1460 2465 1480
rect 2465 1460 2485 1480
rect 2485 1460 2490 1480
rect 2460 1455 2490 1460
rect 2570 1480 2600 1485
rect 2570 1460 2575 1480
rect 2575 1460 2595 1480
rect 2595 1460 2600 1480
rect 2570 1455 2600 1460
rect 2680 1480 2710 1485
rect 2680 1460 2685 1480
rect 2685 1460 2705 1480
rect 2705 1460 2710 1480
rect 2680 1455 2710 1460
rect 2790 1480 2820 1485
rect 2790 1460 2795 1480
rect 2795 1460 2815 1480
rect 2815 1460 2820 1480
rect 2790 1455 2820 1460
rect 3105 1460 3135 1490
rect 2025 930 2055 960
rect 2185 805 2215 810
rect 2185 785 2190 805
rect 2190 785 2210 805
rect 2210 785 2215 805
rect 2185 780 2215 785
rect 2295 805 2325 810
rect 2295 785 2300 805
rect 2300 785 2320 805
rect 2320 785 2325 805
rect 2295 780 2325 785
rect 2405 805 2435 810
rect 2405 785 2410 805
rect 2410 785 2430 805
rect 2430 785 2435 805
rect 2405 780 2435 785
rect 2515 805 2545 810
rect 2515 785 2520 805
rect 2520 785 2540 805
rect 2540 785 2545 805
rect 2515 780 2545 785
rect 2625 805 2655 810
rect 2625 785 2630 805
rect 2630 785 2650 805
rect 2650 785 2655 805
rect 2625 780 2655 785
rect 2735 805 2765 810
rect 2735 785 2740 805
rect 2740 785 2760 805
rect 2760 785 2765 805
rect 2735 780 2765 785
rect 2185 730 2215 760
rect 2025 685 2055 715
rect 2625 730 2655 760
rect 3195 730 3225 760
rect 2460 685 2490 715
rect 3105 685 3135 715
rect 2120 665 2150 670
rect 2120 645 2125 665
rect 2125 645 2145 665
rect 2145 645 2150 665
rect 2120 640 2150 645
rect 2185 665 2215 670
rect 2185 645 2190 665
rect 2190 645 2210 665
rect 2210 645 2215 665
rect 2185 640 2215 645
rect 2295 665 2325 670
rect 2295 645 2300 665
rect 2300 645 2320 665
rect 2320 645 2325 665
rect 2295 640 2325 645
rect 2405 665 2435 670
rect 2405 645 2410 665
rect 2410 645 2430 665
rect 2430 645 2435 665
rect 2405 640 2435 645
rect 2515 665 2545 670
rect 2515 645 2520 665
rect 2520 645 2540 665
rect 2540 645 2545 665
rect 2515 640 2545 645
rect 2625 665 2655 670
rect 2625 645 2630 665
rect 2630 645 2650 665
rect 2650 645 2655 665
rect 2625 640 2655 645
rect 2735 665 2765 670
rect 2735 645 2740 665
rect 2740 645 2760 665
rect 2760 645 2765 665
rect 2735 640 2765 645
rect 2800 665 2830 670
rect 2800 645 2805 665
rect 2805 645 2825 665
rect 2825 645 2830 665
rect 2800 640 2830 645
rect 2240 390 2270 395
rect 2240 370 2245 390
rect 2245 370 2265 390
rect 2265 370 2270 390
rect 2240 365 2270 370
rect 2350 390 2380 395
rect 2350 370 2355 390
rect 2355 370 2375 390
rect 2375 370 2380 390
rect 2350 365 2380 370
rect 2460 390 2490 395
rect 2460 370 2465 390
rect 2465 370 2485 390
rect 2485 370 2490 390
rect 2460 365 2490 370
rect 2570 390 2600 395
rect 2570 370 2575 390
rect 2575 370 2595 390
rect 2595 370 2600 390
rect 2570 365 2600 370
rect 2680 390 2710 395
rect 2680 370 2685 390
rect 2685 370 2705 390
rect 2705 370 2710 390
rect 2680 365 2710 370
rect 2925 365 2955 395
rect 2025 310 2055 340
rect 2405 310 2435 340
rect 2240 280 2270 285
rect 2240 260 2245 280
rect 2245 260 2265 280
rect 2265 260 2270 280
rect 2240 255 2270 260
rect 2350 280 2380 285
rect 2350 260 2355 280
rect 2355 260 2375 280
rect 2375 260 2380 280
rect 2350 255 2380 260
rect 2460 280 2490 285
rect 2460 260 2465 280
rect 2465 260 2485 280
rect 2485 260 2490 280
rect 2460 255 2490 260
rect 2570 280 2600 285
rect 2570 260 2575 280
rect 2575 260 2595 280
rect 2595 260 2600 280
rect 2570 255 2600 260
rect 2680 280 2710 285
rect 2680 260 2685 280
rect 2685 260 2705 280
rect 2705 260 2710 280
rect 2680 255 2710 260
rect 2880 255 2910 285
rect 2185 -95 2215 -90
rect 2185 -115 2190 -95
rect 2190 -115 2210 -95
rect 2210 -115 2215 -95
rect 2185 -120 2215 -115
rect 2295 -95 2325 -90
rect 2295 -115 2300 -95
rect 2300 -115 2320 -95
rect 2320 -115 2325 -95
rect 2295 -120 2325 -115
rect 2405 -95 2435 -90
rect 2405 -115 2410 -95
rect 2410 -115 2430 -95
rect 2430 -115 2435 -95
rect 2405 -120 2435 -115
rect 2515 -95 2545 -90
rect 2515 -115 2520 -95
rect 2520 -115 2540 -95
rect 2540 -115 2545 -95
rect 2515 -120 2545 -115
rect 2625 -95 2655 -90
rect 2625 -115 2630 -95
rect 2630 -115 2650 -95
rect 2650 -115 2655 -95
rect 2625 -120 2655 -115
rect 2735 -95 2765 -90
rect 2735 -115 2740 -95
rect 2740 -115 2760 -95
rect 2760 -115 2765 -95
rect 2735 -120 2765 -115
rect 2880 -120 2910 -90
rect 3195 320 3225 350
rect 2969 -93 2996 -85
rect 2969 -113 2970 -93
rect 2970 -113 2995 -93
rect 2995 -113 2996 -93
rect 2969 -120 2996 -113
rect 3029 -93 3056 -85
rect 3029 -113 3030 -93
rect 3030 -113 3055 -93
rect 3055 -113 3056 -93
rect 3029 -120 3056 -113
rect 3089 -93 3116 -85
rect 3089 -113 3090 -93
rect 3090 -113 3115 -93
rect 3115 -113 3116 -93
rect 3089 -120 3116 -113
rect 3149 -93 3176 -85
rect 3149 -113 3150 -93
rect 3150 -113 3175 -93
rect 3175 -113 3176 -93
rect 3149 -120 3176 -113
rect 2120 -175 2150 -145
rect 2800 -175 2830 -145
rect 2925 -175 2955 -145
rect 3025 -175 3060 -145
rect 1980 -220 2010 -190
rect 3145 -220 3180 -190
rect 2280 -275 2310 -245
rect 2865 -275 2900 -245
rect 1945 -340 1975 -310
rect 2180 -305 2210 -300
rect 2180 -325 2185 -305
rect 2185 -325 2205 -305
rect 2205 -325 2210 -305
rect 2180 -330 2210 -325
rect 2380 -305 2410 -300
rect 2380 -325 2385 -305
rect 2385 -325 2405 -305
rect 2405 -325 2410 -305
rect 2380 -330 2410 -325
rect 2580 -305 2610 -300
rect 2580 -325 2585 -305
rect 2585 -325 2605 -305
rect 2605 -325 2610 -305
rect 2580 -330 2610 -325
rect 2805 -330 2840 -300
rect 1890 -385 1920 -355
rect 1340 -455 1370 -425
rect 1845 -455 1875 -425
rect 195 -510 225 -480
rect 390 -485 420 -480
rect 390 -505 395 -485
rect 395 -505 415 -485
rect 415 -505 420 -485
rect 390 -510 420 -505
rect 500 -485 530 -480
rect 500 -505 505 -485
rect 505 -505 525 -485
rect 525 -505 530 -485
rect 500 -510 530 -505
rect 610 -485 640 -480
rect 610 -505 615 -485
rect 615 -505 635 -485
rect 635 -505 640 -485
rect 610 -510 640 -505
rect 720 -485 750 -480
rect 720 -505 725 -485
rect 725 -505 745 -485
rect 745 -505 750 -485
rect 720 -510 750 -505
rect 830 -485 860 -480
rect 830 -505 835 -485
rect 835 -505 855 -485
rect 855 -505 860 -485
rect 830 -510 860 -505
rect 940 -485 970 -480
rect 940 -505 945 -485
rect 945 -505 965 -485
rect 965 -505 970 -485
rect 940 -510 970 -505
rect 1050 -485 1080 -480
rect 1050 -505 1055 -485
rect 1055 -505 1075 -485
rect 1075 -505 1080 -485
rect 1050 -510 1080 -505
rect 1160 -485 1190 -480
rect 1160 -505 1165 -485
rect 1165 -505 1185 -485
rect 1185 -505 1190 -485
rect 1160 -510 1190 -505
rect 1270 -485 1300 -480
rect 1270 -505 1275 -485
rect 1275 -505 1295 -485
rect 1295 -505 1300 -485
rect 1270 -510 1300 -505
rect 1395 -485 1425 -480
rect 1395 -505 1400 -485
rect 1400 -505 1420 -485
rect 1420 -505 1425 -485
rect 1395 -510 1425 -505
rect 3195 -330 3225 -300
rect 2809 -387 2836 -380
rect 2809 -407 2810 -387
rect 2810 -407 2835 -387
rect 2835 -407 2836 -387
rect 2809 -415 2836 -407
rect 2869 -387 2896 -380
rect 2869 -407 2870 -387
rect 2870 -407 2895 -387
rect 2895 -407 2896 -387
rect 2869 -415 2896 -407
rect 270 -810 300 -805
rect 270 -830 275 -810
rect 275 -830 295 -810
rect 295 -830 300 -810
rect 270 -835 300 -830
rect 335 -810 365 -805
rect 335 -830 340 -810
rect 340 -830 360 -810
rect 360 -830 365 -810
rect 335 -835 365 -830
rect 445 -810 475 -805
rect 445 -830 450 -810
rect 450 -830 470 -810
rect 470 -830 475 -810
rect 445 -835 475 -830
rect 555 -810 585 -805
rect 555 -830 560 -810
rect 560 -830 580 -810
rect 580 -830 585 -810
rect 555 -835 585 -830
rect 665 -810 695 -805
rect 665 -830 670 -810
rect 670 -830 690 -810
rect 690 -830 695 -810
rect 665 -835 695 -830
rect 775 -810 805 -805
rect 775 -830 780 -810
rect 780 -830 800 -810
rect 800 -830 805 -810
rect 775 -835 805 -830
rect 885 -810 915 -805
rect 885 -830 890 -810
rect 890 -830 910 -810
rect 910 -830 915 -810
rect 885 -835 915 -830
rect 995 -810 1025 -805
rect 995 -830 1000 -810
rect 1000 -830 1020 -810
rect 1020 -830 1025 -810
rect 995 -835 1025 -830
rect 1105 -810 1135 -805
rect 1105 -830 1110 -810
rect 1110 -830 1130 -810
rect 1130 -830 1135 -810
rect 1105 -835 1135 -830
rect 1215 -810 1245 -805
rect 1215 -830 1220 -810
rect 1220 -830 1240 -810
rect 1240 -830 1245 -810
rect 1215 -835 1245 -830
rect 1325 -810 1355 -805
rect 1325 -830 1330 -810
rect 1330 -830 1350 -810
rect 1350 -830 1355 -810
rect 1325 -835 1355 -830
rect 1435 -810 1465 -805
rect 1435 -830 1440 -810
rect 1440 -830 1460 -810
rect 1460 -830 1465 -810
rect 1435 -835 1465 -830
rect 1935 -835 1965 -805
rect 195 -885 225 -855
rect 1320 -870 1350 -865
rect 1320 -890 1325 -870
rect 1325 -890 1345 -870
rect 1345 -890 1350 -870
rect 1320 -895 1350 -890
rect -185 -930 -155 -900
rect 555 -905 585 -900
rect 555 -925 560 -905
rect 560 -925 580 -905
rect 580 -925 585 -905
rect 555 -930 585 -925
rect 665 -905 695 -900
rect 665 -925 670 -905
rect 670 -925 690 -905
rect 690 -925 695 -905
rect 665 -930 695 -925
rect 775 -905 805 -900
rect 775 -925 780 -905
rect 780 -925 800 -905
rect 800 -925 805 -905
rect 775 -930 805 -925
rect 1010 -905 1040 -900
rect 1010 -925 1015 -905
rect 1015 -925 1035 -905
rect 1035 -925 1040 -905
rect 1010 -930 1040 -925
rect 1130 -905 1160 -900
rect 1130 -925 1135 -905
rect 1135 -925 1155 -905
rect 1155 -925 1160 -905
rect 1130 -930 1160 -925
rect 1260 -905 1290 -900
rect 1260 -925 1265 -905
rect 1265 -925 1285 -905
rect 1285 -925 1290 -905
rect 1260 -930 1290 -925
rect 930 -1015 960 -1010
rect 930 -1035 935 -1015
rect 935 -1035 955 -1015
rect 955 -1035 960 -1015
rect 930 -1040 960 -1035
rect 610 -1125 640 -1120
rect 610 -1145 615 -1125
rect 615 -1145 635 -1125
rect 635 -1145 640 -1125
rect 610 -1150 640 -1145
rect 720 -1125 750 -1120
rect 720 -1145 725 -1125
rect 725 -1145 745 -1125
rect 745 -1145 750 -1125
rect 720 -1150 750 -1145
rect 930 -1150 960 -1120
rect 2080 -1080 2110 -1075
rect 2080 -1100 2085 -1080
rect 2085 -1100 2105 -1080
rect 2105 -1100 2110 -1080
rect 2080 -1105 2110 -1100
rect 2280 -1080 2310 -1075
rect 2280 -1100 2285 -1080
rect 2285 -1100 2305 -1080
rect 2305 -1100 2310 -1080
rect 2280 -1105 2310 -1100
rect 2380 -1105 2410 -1075
rect 2480 -1080 2510 -1075
rect 2480 -1100 2485 -1080
rect 2485 -1100 2505 -1080
rect 2505 -1100 2510 -1080
rect 2480 -1105 2510 -1100
rect 2680 -1080 2710 -1075
rect 2680 -1100 2685 -1080
rect 2685 -1100 2705 -1080
rect 2705 -1100 2710 -1080
rect 2680 -1105 2710 -1100
rect -720 -1205 -690 -1175
rect -275 -1205 -245 -1175
rect 500 -1205 530 -1175
rect 830 -1205 860 -1175
rect 1935 -1205 1965 -1175
rect 2380 -1205 2410 -1175
rect 830 -2455 860 -2425
<< metal2 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 150 2780 190 2785
rect 150 2750 155 2780
rect 185 2775 190 2780
rect 620 2780 660 2785
rect 620 2775 625 2780
rect 185 2755 625 2775
rect 185 2750 190 2755
rect 150 2745 190 2750
rect 620 2750 625 2755
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2775 1070 2780
rect 1498 2780 1538 2785
rect 1498 2775 1503 2780
rect 1065 2755 1503 2775
rect 1065 2750 1070 2755
rect 1030 2745 1070 2750
rect 1498 2750 1503 2755
rect 1533 2750 1538 2780
rect 1498 2745 1538 2750
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2720 70 2725
rect 150 2725 190 2730
rect 150 2720 155 2725
rect 65 2700 155 2720
rect 65 2695 70 2700
rect 30 2690 70 2695
rect 150 2695 155 2700
rect 185 2720 190 2725
rect 210 2725 250 2730
rect 210 2720 215 2725
rect 185 2700 215 2720
rect 185 2695 190 2700
rect 150 2690 190 2695
rect 210 2695 215 2700
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2720 865 2725
rect 970 2725 1010 2730
rect 970 2720 975 2725
rect 860 2700 975 2720
rect 860 2695 865 2700
rect 825 2690 865 2695
rect 970 2695 975 2700
rect 1005 2720 1010 2725
rect 1090 2725 1130 2730
rect 1090 2720 1095 2725
rect 1005 2700 1095 2720
rect 1005 2695 1010 2700
rect 970 2690 1010 2695
rect 1090 2695 1095 2700
rect 1125 2720 1130 2725
rect 1150 2725 1190 2730
rect 1150 2720 1155 2725
rect 1125 2700 1155 2720
rect 1125 2695 1130 2700
rect 1090 2690 1130 2695
rect 1150 2695 1155 2700
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1438 2725 1478 2730
rect 1438 2695 1443 2725
rect 1473 2720 1478 2725
rect 1498 2725 1538 2730
rect 1498 2720 1503 2725
rect 1473 2700 1503 2720
rect 1473 2695 1478 2700
rect 1438 2690 1478 2695
rect 1498 2695 1503 2700
rect 1533 2720 1538 2725
rect 1618 2725 1658 2730
rect 1618 2720 1623 2725
rect 1533 2700 1623 2720
rect 1533 2695 1538 2700
rect 1498 2690 1538 2695
rect 1618 2695 1623 2700
rect 1653 2695 1658 2725
rect 1618 2690 1658 2695
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2550 540 2555
rect 560 2555 600 2560
rect 560 2550 565 2555
rect 535 2530 565 2550
rect 535 2525 540 2530
rect 500 2520 540 2525
rect 560 2525 565 2530
rect 595 2550 600 2555
rect 680 2555 720 2560
rect 680 2550 685 2555
rect 595 2530 685 2550
rect 595 2525 600 2530
rect 560 2520 600 2525
rect 680 2525 685 2530
rect 715 2550 720 2555
rect 825 2555 865 2560
rect 825 2550 830 2555
rect 715 2530 830 2550
rect 715 2525 720 2530
rect 680 2520 720 2525
rect 825 2525 830 2530
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2300 115 2305
rect 139 2305 169 2310
rect 110 2280 139 2300
rect 110 2275 115 2280
rect 75 2270 115 2275
rect 609 2305 639 2310
rect 169 2280 609 2300
rect 139 2270 169 2275
rect 770 2305 810 2310
rect 770 2300 775 2305
rect 639 2280 775 2300
rect 609 2270 639 2275
rect 770 2275 775 2280
rect 805 2300 810 2305
rect 1519 2305 1549 2310
rect 805 2280 1519 2300
rect 805 2275 810 2280
rect 770 2270 810 2275
rect 1519 2270 1549 2275
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2245 920 2260
rect 1045 2250 1085 2255
rect 1045 2245 1050 2250
rect 915 2230 1050 2245
rect 880 2225 1050 2230
rect 1045 2220 1050 2225
rect 1080 2245 1085 2250
rect 1573 2250 1613 2255
rect 1573 2245 1578 2250
rect 1080 2225 1578 2245
rect 1080 2220 1085 2225
rect 1045 2215 1085 2220
rect 1573 2220 1578 2225
rect 1608 2220 1613 2250
rect 1573 2215 1613 2220
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2200 -765 2205
rect -235 2205 -195 2210
rect -235 2200 -230 2205
rect -770 2180 -230 2200
rect -770 2175 -765 2180
rect -805 2170 -765 2175
rect -235 2175 -230 2180
rect -200 2200 -195 2205
rect 825 2205 865 2210
rect 825 2200 830 2205
rect -200 2180 830 2200
rect -200 2175 -195 2180
rect -235 2170 -195 2175
rect 825 2175 830 2180
rect 860 2200 865 2205
rect 1885 2205 1925 2210
rect 1885 2200 1890 2205
rect 860 2180 1890 2200
rect 860 2175 865 2180
rect 825 2170 865 2175
rect 1885 2175 1890 2180
rect 1920 2200 1925 2205
rect 2455 2205 2495 2210
rect 2455 2200 2460 2205
rect 1920 2180 2460 2200
rect 1920 2175 1925 2180
rect 1885 2170 1925 2175
rect 2455 2175 2460 2180
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect -1165 2150 -1125 2155
rect -1165 2120 -1160 2150
rect -1130 2145 -1125 2150
rect -1045 2150 -1005 2155
rect -1045 2145 -1040 2150
rect -1130 2125 -1040 2145
rect -1130 2120 -1125 2125
rect -1165 2115 -1125 2120
rect -1045 2120 -1040 2125
rect -1010 2145 -1005 2150
rect -925 2150 -885 2155
rect -925 2145 -920 2150
rect -1010 2125 -920 2145
rect -1010 2120 -1005 2125
rect -1045 2115 -1005 2120
rect -925 2120 -920 2125
rect -890 2145 -885 2150
rect -805 2150 -765 2155
rect -805 2145 -800 2150
rect -890 2125 -800 2145
rect -890 2120 -885 2125
rect -925 2115 -885 2120
rect -805 2120 -800 2125
rect -770 2145 -765 2150
rect -685 2150 -645 2155
rect -685 2145 -680 2150
rect -770 2125 -680 2145
rect -770 2120 -765 2125
rect -805 2115 -765 2120
rect -685 2120 -680 2125
rect -650 2145 -645 2150
rect -565 2150 -525 2155
rect -565 2145 -560 2150
rect -650 2125 -560 2145
rect -650 2120 -645 2125
rect -685 2115 -645 2120
rect -565 2120 -560 2125
rect -530 2145 -525 2150
rect -445 2150 -405 2155
rect -445 2145 -440 2150
rect -530 2125 -440 2145
rect -530 2120 -525 2125
rect -565 2115 -525 2120
rect -445 2120 -440 2125
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2145 -240 2150
rect -40 2150 0 2155
rect -40 2145 -35 2150
rect -245 2125 -35 2145
rect -245 2120 -240 2125
rect -280 2115 -240 2120
rect -40 2120 -35 2125
rect -5 2145 0 2150
rect 80 2150 120 2155
rect 80 2145 85 2150
rect -5 2125 85 2145
rect -5 2120 0 2125
rect -40 2115 0 2120
rect 80 2120 85 2125
rect 115 2145 120 2150
rect 200 2150 240 2155
rect 200 2145 205 2150
rect 115 2125 205 2145
rect 115 2120 120 2125
rect 80 2115 120 2120
rect 200 2120 205 2125
rect 235 2145 240 2150
rect 320 2150 360 2155
rect 320 2145 325 2150
rect 235 2125 325 2145
rect 235 2120 240 2125
rect 200 2115 240 2120
rect 320 2120 325 2125
rect 355 2145 360 2150
rect 440 2150 480 2155
rect 440 2145 445 2150
rect 355 2125 445 2145
rect 355 2120 360 2125
rect 320 2115 360 2120
rect 440 2120 445 2125
rect 475 2145 480 2150
rect 560 2150 600 2155
rect 560 2145 565 2150
rect 475 2125 565 2145
rect 475 2120 480 2125
rect 440 2115 480 2120
rect 560 2120 565 2125
rect 595 2145 600 2150
rect 680 2150 720 2155
rect 680 2145 685 2150
rect 595 2125 685 2145
rect 595 2120 600 2125
rect 560 2115 600 2120
rect 680 2120 685 2125
rect 715 2120 720 2150
rect 680 2115 720 2120
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2145 1010 2150
rect 1090 2150 1130 2155
rect 1090 2145 1095 2150
rect 1005 2125 1095 2145
rect 1005 2120 1010 2125
rect 970 2115 1010 2120
rect 1090 2120 1095 2125
rect 1125 2145 1130 2150
rect 1210 2150 1250 2155
rect 1210 2145 1215 2150
rect 1125 2125 1215 2145
rect 1125 2120 1130 2125
rect 1090 2115 1130 2120
rect 1210 2120 1215 2125
rect 1245 2145 1250 2150
rect 1330 2150 1370 2155
rect 1330 2145 1335 2150
rect 1245 2125 1335 2145
rect 1245 2120 1250 2125
rect 1210 2115 1250 2120
rect 1330 2120 1335 2125
rect 1365 2145 1370 2150
rect 1450 2150 1490 2155
rect 1450 2145 1455 2150
rect 1365 2125 1455 2145
rect 1365 2120 1370 2125
rect 1330 2115 1370 2120
rect 1450 2120 1455 2125
rect 1485 2145 1490 2150
rect 1570 2150 1610 2155
rect 1570 2145 1575 2150
rect 1485 2125 1575 2145
rect 1485 2120 1490 2125
rect 1450 2115 1490 2120
rect 1570 2120 1575 2125
rect 1605 2145 1610 2150
rect 1690 2150 1730 2155
rect 1690 2145 1695 2150
rect 1605 2125 1695 2145
rect 1605 2120 1610 2125
rect 1570 2115 1610 2120
rect 1690 2120 1695 2125
rect 1725 2145 1730 2150
rect 1930 2150 1970 2155
rect 1930 2145 1935 2150
rect 1725 2125 1935 2145
rect 1725 2120 1730 2125
rect 1690 2115 1730 2120
rect 1930 2120 1935 2125
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2145 2135 2150
rect 2215 2150 2255 2155
rect 2215 2145 2220 2150
rect 2130 2125 2220 2145
rect 2130 2120 2135 2125
rect 2095 2115 2135 2120
rect 2215 2120 2220 2125
rect 2250 2145 2255 2150
rect 2335 2150 2375 2155
rect 2335 2145 2340 2150
rect 2250 2125 2340 2145
rect 2250 2120 2255 2125
rect 2215 2115 2255 2120
rect 2335 2120 2340 2125
rect 2370 2145 2375 2150
rect 2455 2150 2495 2155
rect 2455 2145 2460 2150
rect 2370 2125 2460 2145
rect 2370 2120 2375 2125
rect 2335 2115 2375 2120
rect 2455 2120 2460 2125
rect 2490 2145 2495 2150
rect 2575 2150 2615 2155
rect 2575 2145 2580 2150
rect 2490 2125 2580 2145
rect 2490 2120 2495 2125
rect 2455 2115 2495 2120
rect 2575 2120 2580 2125
rect 2610 2145 2615 2150
rect 2695 2150 2735 2155
rect 2695 2145 2700 2150
rect 2610 2125 2700 2145
rect 2610 2120 2615 2125
rect 2575 2115 2615 2120
rect 2695 2120 2700 2125
rect 2730 2145 2735 2150
rect 2815 2150 2855 2155
rect 2815 2145 2820 2150
rect 2730 2125 2820 2145
rect 2730 2120 2735 2125
rect 2695 2115 2735 2120
rect 2815 2120 2820 2125
rect 2850 2120 2855 2150
rect 2815 2115 2855 2120
rect -1105 1725 -1065 1730
rect -1105 1695 -1100 1725
rect -1070 1720 -1065 1725
rect -985 1725 -945 1730
rect -985 1720 -980 1725
rect -1070 1700 -980 1720
rect -1070 1695 -1065 1700
rect -1105 1690 -1065 1695
rect -985 1695 -980 1700
rect -950 1720 -945 1725
rect -865 1725 -825 1730
rect -865 1720 -860 1725
rect -950 1700 -860 1720
rect -950 1695 -945 1700
rect -985 1690 -945 1695
rect -865 1695 -860 1700
rect -830 1720 -825 1725
rect -745 1725 -705 1730
rect -745 1720 -740 1725
rect -830 1700 -740 1720
rect -830 1695 -825 1700
rect -865 1690 -825 1695
rect -745 1695 -740 1700
rect -710 1720 -705 1725
rect -625 1725 -585 1730
rect -625 1720 -620 1725
rect -710 1700 -620 1720
rect -710 1695 -705 1700
rect -745 1690 -705 1695
rect -625 1695 -620 1700
rect -590 1720 -585 1725
rect -505 1725 -465 1730
rect -505 1720 -500 1725
rect -590 1700 -500 1720
rect -590 1695 -585 1700
rect -625 1690 -585 1695
rect -505 1695 -500 1700
rect -470 1720 -465 1725
rect -280 1725 -240 1730
rect -280 1720 -275 1725
rect -470 1700 -275 1720
rect -470 1695 -465 1700
rect -505 1690 -465 1695
rect -280 1695 -275 1700
rect -245 1695 -240 1725
rect -280 1690 -240 1695
rect 20 1725 60 1730
rect 20 1695 25 1725
rect 55 1720 60 1725
rect 140 1725 180 1730
rect 140 1720 145 1725
rect 55 1700 145 1720
rect 55 1695 60 1700
rect 20 1690 60 1695
rect 140 1695 145 1700
rect 175 1720 180 1725
rect 260 1725 300 1730
rect 260 1720 265 1725
rect 175 1700 265 1720
rect 175 1695 180 1700
rect 140 1690 180 1695
rect 260 1695 265 1700
rect 295 1720 300 1725
rect 380 1725 420 1730
rect 380 1720 385 1725
rect 295 1700 385 1720
rect 295 1695 300 1700
rect 260 1690 300 1695
rect 380 1695 385 1700
rect 415 1720 420 1725
rect 500 1725 540 1730
rect 500 1720 505 1725
rect 415 1700 505 1720
rect 415 1695 420 1700
rect 380 1690 420 1695
rect 500 1695 505 1700
rect 535 1720 540 1725
rect 620 1725 660 1730
rect 620 1720 625 1725
rect 535 1700 625 1720
rect 535 1695 540 1700
rect 500 1690 540 1695
rect 620 1695 625 1700
rect 655 1695 660 1725
rect 620 1690 660 1695
rect 1030 1725 1070 1730
rect 1030 1695 1035 1725
rect 1065 1720 1070 1725
rect 1150 1725 1190 1730
rect 1150 1720 1155 1725
rect 1065 1700 1155 1720
rect 1065 1695 1070 1700
rect 1030 1690 1070 1695
rect 1150 1695 1155 1700
rect 1185 1720 1190 1725
rect 1270 1725 1310 1730
rect 1270 1720 1275 1725
rect 1185 1700 1275 1720
rect 1185 1695 1190 1700
rect 1150 1690 1190 1695
rect 1270 1695 1275 1700
rect 1305 1720 1310 1725
rect 1390 1725 1430 1730
rect 1390 1720 1395 1725
rect 1305 1700 1395 1720
rect 1305 1695 1310 1700
rect 1270 1690 1310 1695
rect 1390 1695 1395 1700
rect 1425 1720 1430 1725
rect 1510 1725 1550 1730
rect 1510 1720 1515 1725
rect 1425 1700 1515 1720
rect 1425 1695 1430 1700
rect 1390 1690 1430 1695
rect 1510 1695 1515 1700
rect 1545 1720 1550 1725
rect 1630 1725 1670 1730
rect 1630 1720 1635 1725
rect 1545 1700 1635 1720
rect 1545 1695 1550 1700
rect 1510 1690 1550 1695
rect 1630 1695 1635 1700
rect 1665 1695 1670 1725
rect 1630 1690 1670 1695
rect 1930 1725 1970 1730
rect 1930 1695 1935 1725
rect 1965 1720 1970 1725
rect 2155 1725 2195 1730
rect 2155 1720 2160 1725
rect 1965 1700 2160 1720
rect 1965 1695 1970 1700
rect 1930 1690 1970 1695
rect 2155 1695 2160 1700
rect 2190 1720 2195 1725
rect 2275 1725 2315 1730
rect 2275 1720 2280 1725
rect 2190 1700 2280 1720
rect 2190 1695 2195 1700
rect 2155 1690 2195 1695
rect 2275 1695 2280 1700
rect 2310 1720 2315 1725
rect 2395 1725 2435 1730
rect 2395 1720 2400 1725
rect 2310 1700 2400 1720
rect 2310 1695 2315 1700
rect 2275 1690 2315 1695
rect 2395 1695 2400 1700
rect 2430 1720 2435 1725
rect 2515 1725 2555 1730
rect 2515 1720 2520 1725
rect 2430 1700 2520 1720
rect 2430 1695 2435 1700
rect 2395 1690 2435 1695
rect 2515 1695 2520 1700
rect 2550 1720 2555 1725
rect 2635 1725 2675 1730
rect 2635 1720 2640 1725
rect 2550 1700 2640 1720
rect 2550 1695 2555 1700
rect 2515 1690 2555 1695
rect 2635 1695 2640 1700
rect 2670 1720 2675 1725
rect 2755 1725 2795 1730
rect 2755 1720 2760 1725
rect 2670 1700 2760 1720
rect 2670 1695 2675 1700
rect 2635 1690 2675 1695
rect 2755 1695 2760 1700
rect 2790 1695 2795 1725
rect 2755 1690 2795 1695
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1665 -330 1670
rect 20 1670 60 1675
rect 20 1665 25 1670
rect -335 1645 25 1665
rect -335 1640 -330 1645
rect -370 1635 -330 1640
rect 20 1640 25 1645
rect 55 1640 60 1670
rect 20 1635 60 1640
rect 320 1670 360 1675
rect 320 1640 325 1670
rect 355 1665 360 1670
rect 780 1670 820 1675
rect 780 1665 785 1670
rect 355 1645 785 1665
rect 355 1640 360 1645
rect 320 1635 360 1640
rect 780 1640 785 1645
rect 815 1665 820 1670
rect 1330 1670 1370 1675
rect 1330 1665 1335 1670
rect 815 1645 1335 1665
rect 815 1640 820 1645
rect 780 1635 820 1640
rect 1330 1640 1335 1645
rect 1365 1640 1370 1670
rect 1330 1635 1370 1640
rect 1630 1670 1670 1675
rect 1630 1640 1635 1670
rect 1665 1665 1670 1670
rect 2020 1670 2060 1675
rect 2020 1665 2025 1670
rect 1665 1645 2025 1665
rect 1665 1640 1670 1645
rect 1630 1635 1670 1640
rect 2020 1640 2025 1645
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect -805 1625 -765 1630
rect -805 1595 -800 1625
rect -770 1620 -765 1625
rect 870 1620 875 1630
rect -770 1600 875 1620
rect 905 1620 910 1630
rect 2455 1625 2495 1630
rect 2455 1620 2460 1625
rect 905 1600 2460 1620
rect -770 1595 -765 1600
rect -805 1590 -765 1595
rect 2455 1595 2460 1600
rect 2490 1595 2495 1625
rect 2455 1590 2495 1595
rect 455 1580 495 1585
rect 455 1550 460 1580
rect 490 1575 495 1580
rect 625 1580 655 1585
rect 490 1555 625 1575
rect 490 1550 495 1555
rect 455 1545 495 1550
rect 785 1580 825 1585
rect 785 1575 790 1580
rect 655 1555 790 1575
rect 625 1545 655 1550
rect 785 1550 790 1555
rect 820 1575 825 1580
rect 865 1580 905 1585
rect 865 1575 870 1580
rect 820 1555 870 1575
rect 820 1550 825 1555
rect 785 1545 825 1550
rect 865 1550 870 1555
rect 900 1575 905 1580
rect 1035 1580 1065 1585
rect 900 1555 1035 1575
rect 900 1550 905 1555
rect 865 1545 905 1550
rect 1195 1580 1235 1585
rect 1195 1575 1200 1580
rect 1065 1555 1200 1575
rect 1035 1545 1065 1550
rect 1195 1550 1200 1555
rect 1230 1575 1235 1580
rect 1885 1580 1925 1585
rect 1885 1575 1890 1580
rect 1230 1555 1890 1575
rect 1230 1550 1235 1555
rect 1195 1545 1235 1550
rect 1885 1550 1890 1555
rect 1920 1550 1925 1580
rect 1885 1545 1925 1550
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect 565 1535 605 1540
rect 565 1505 570 1535
rect 600 1530 605 1535
rect 675 1535 715 1540
rect 675 1530 680 1535
rect 600 1510 680 1530
rect 600 1505 605 1510
rect 565 1500 605 1505
rect 675 1505 680 1510
rect 710 1505 715 1535
rect 675 1500 715 1505
rect 975 1535 1015 1540
rect 975 1505 980 1535
rect 1010 1530 1015 1535
rect 1085 1535 1125 1540
rect 1085 1530 1090 1535
rect 1010 1510 1090 1530
rect 1010 1505 1015 1510
rect 975 1500 1015 1505
rect 1085 1505 1090 1510
rect 1120 1505 1125 1535
rect 1085 1500 1125 1505
rect 3100 1490 3140 1495
rect -1135 1485 -1095 1490
rect -1135 1455 -1130 1485
rect -1100 1480 -1095 1485
rect -1025 1485 -985 1490
rect -1025 1480 -1020 1485
rect -1100 1460 -1020 1480
rect -1100 1455 -1095 1460
rect -1135 1450 -1095 1455
rect -1025 1455 -1020 1460
rect -990 1480 -985 1485
rect -915 1485 -875 1490
rect -915 1480 -910 1485
rect -990 1460 -910 1480
rect -990 1455 -985 1460
rect -1025 1450 -985 1455
rect -915 1455 -910 1460
rect -880 1480 -875 1485
rect -805 1485 -765 1490
rect -805 1480 -800 1485
rect -880 1460 -800 1480
rect -880 1455 -875 1460
rect -915 1450 -875 1455
rect -805 1455 -800 1460
rect -770 1480 -765 1485
rect -695 1485 -655 1490
rect -695 1480 -690 1485
rect -770 1460 -690 1480
rect -770 1455 -765 1460
rect -805 1450 -765 1455
rect -695 1455 -690 1460
rect -660 1480 -655 1485
rect -585 1485 -545 1490
rect -585 1480 -580 1485
rect -660 1460 -580 1480
rect -660 1455 -655 1460
rect -695 1450 -655 1455
rect -585 1455 -580 1460
rect -550 1480 -545 1485
rect -475 1485 -435 1490
rect -475 1480 -470 1485
rect -550 1460 -470 1480
rect -550 1455 -545 1460
rect -585 1450 -545 1455
rect -475 1455 -470 1460
rect -440 1480 -435 1485
rect -235 1485 -195 1490
rect -235 1480 -230 1485
rect -440 1460 -230 1480
rect -440 1455 -435 1460
rect -475 1450 -435 1455
rect -235 1455 -230 1460
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 1885 1485 1925 1490
rect 1885 1455 1890 1485
rect 1920 1480 1925 1485
rect 2125 1485 2165 1490
rect 2125 1480 2130 1485
rect 1920 1460 2130 1480
rect 1920 1455 1925 1460
rect 1885 1450 1925 1455
rect 2125 1455 2130 1460
rect 2160 1480 2165 1485
rect 2235 1485 2275 1490
rect 2235 1480 2240 1485
rect 2160 1460 2240 1480
rect 2160 1455 2165 1460
rect 2125 1450 2165 1455
rect 2235 1455 2240 1460
rect 2270 1480 2275 1485
rect 2345 1485 2385 1490
rect 2345 1480 2350 1485
rect 2270 1460 2350 1480
rect 2270 1455 2275 1460
rect 2235 1450 2275 1455
rect 2345 1455 2350 1460
rect 2380 1480 2385 1485
rect 2455 1485 2495 1490
rect 2455 1480 2460 1485
rect 2380 1460 2460 1480
rect 2380 1455 2385 1460
rect 2345 1450 2385 1455
rect 2455 1455 2460 1460
rect 2490 1480 2495 1485
rect 2565 1485 2605 1490
rect 2565 1480 2570 1485
rect 2490 1460 2570 1480
rect 2490 1455 2495 1460
rect 2455 1450 2495 1455
rect 2565 1455 2570 1460
rect 2600 1480 2605 1485
rect 2675 1485 2715 1490
rect 2675 1480 2680 1485
rect 2600 1460 2680 1480
rect 2600 1455 2605 1460
rect 2565 1450 2605 1455
rect 2675 1455 2680 1460
rect 2710 1480 2715 1485
rect 2785 1485 2825 1490
rect 2785 1480 2790 1485
rect 2710 1460 2790 1480
rect 2710 1455 2715 1460
rect 2675 1450 2715 1455
rect 2785 1455 2790 1460
rect 2820 1455 2825 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2785 1450 2825 1455
rect 505 1225 535 1230
rect 745 1225 775 1230
rect 620 1215 660 1220
rect 620 1210 625 1215
rect 535 1195 625 1210
rect 505 1190 625 1195
rect 620 1185 625 1190
rect 655 1210 660 1215
rect 655 1195 745 1210
rect 1030 1215 1070 1220
rect 1030 1210 1035 1215
rect 775 1195 1035 1210
rect 655 1190 1035 1195
rect 655 1185 660 1190
rect 620 1180 660 1185
rect 1030 1185 1035 1190
rect 1065 1210 1070 1215
rect 1065 1190 1075 1210
rect 1065 1185 1070 1190
rect 1030 1180 1070 1185
rect 545 1155 585 1160
rect 545 1150 550 1155
rect 310 1130 550 1150
rect 545 1125 550 1130
rect 580 1150 585 1155
rect 1105 1155 1145 1160
rect 1105 1150 1110 1155
rect 580 1130 1110 1150
rect 580 1125 585 1130
rect 545 1120 585 1125
rect 1105 1125 1110 1130
rect 1140 1125 1145 1155
rect 1105 1120 1145 1125
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1100 -285 1105
rect 690 1105 730 1110
rect 690 1100 695 1105
rect -290 1080 695 1100
rect -290 1075 -285 1080
rect -325 1070 -285 1075
rect 690 1075 695 1080
rect 725 1100 730 1105
rect 960 1105 1000 1110
rect 960 1100 965 1105
rect 725 1080 965 1100
rect 725 1075 730 1080
rect 690 1070 730 1075
rect 960 1075 965 1080
rect 995 1100 1000 1105
rect 1975 1105 2015 1110
rect 1975 1100 1980 1105
rect 995 1080 1980 1100
rect 995 1075 1000 1080
rect 960 1070 1000 1075
rect 1975 1075 1980 1080
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1055 835 1060
rect 905 1060 945 1065
rect 905 1055 910 1060
rect 830 1035 910 1055
rect 830 1030 835 1035
rect 795 1025 835 1030
rect 905 1030 910 1035
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 1155 1015 1195 1020
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 1000 920 1005
rect 1155 1000 1160 1015
rect 915 985 1160 1000
rect 1190 1000 1195 1015
rect 1840 1005 1880 1010
rect 1840 1000 1845 1005
rect 1190 985 1845 1000
rect 915 980 1845 985
rect 915 975 920 980
rect 880 970 920 975
rect 1840 975 1845 980
rect 1875 975 1880 1005
rect 1840 970 1880 975
rect -370 960 -330 965
rect -370 930 -365 960
rect -335 955 -330 960
rect -50 960 -10 965
rect -50 955 -45 960
rect -335 935 -45 955
rect -335 930 -330 935
rect -370 925 -330 930
rect -50 930 -45 935
rect -15 955 -10 960
rect 60 960 100 965
rect 60 955 65 960
rect -15 935 65 955
rect -15 930 -10 935
rect -50 925 -10 930
rect 60 930 65 935
rect 95 955 100 960
rect 170 960 210 965
rect 170 955 175 960
rect 95 935 175 955
rect 95 930 100 935
rect 60 925 100 930
rect 170 930 175 935
rect 205 955 210 960
rect 280 960 320 965
rect 280 955 285 960
rect 205 935 285 955
rect 205 930 210 935
rect 170 925 210 930
rect 280 930 285 935
rect 315 955 320 960
rect 390 960 430 965
rect 390 955 395 960
rect 315 935 395 955
rect 315 930 320 935
rect 280 925 320 930
rect 390 930 395 935
rect 425 955 430 960
rect 500 960 540 965
rect 500 955 505 960
rect 425 935 505 955
rect 425 930 430 935
rect 390 925 430 930
rect 500 930 505 935
rect 535 930 540 960
rect 500 925 540 930
rect 1150 960 1190 965
rect 1150 930 1155 960
rect 1185 955 1190 960
rect 1260 960 1300 965
rect 1260 955 1265 960
rect 1185 935 1265 955
rect 1185 930 1190 935
rect 1150 925 1190 930
rect 1260 930 1265 935
rect 1295 955 1300 960
rect 1370 960 1410 965
rect 1370 955 1375 960
rect 1295 935 1375 955
rect 1295 930 1300 935
rect 1260 925 1300 930
rect 1370 930 1375 935
rect 1405 955 1410 960
rect 1480 960 1520 965
rect 1480 955 1485 960
rect 1405 935 1485 955
rect 1405 930 1410 935
rect 1370 925 1410 930
rect 1480 930 1485 935
rect 1515 955 1520 960
rect 1590 960 1630 965
rect 1590 955 1595 960
rect 1515 935 1595 955
rect 1515 930 1520 935
rect 1480 925 1520 930
rect 1590 930 1595 935
rect 1625 955 1630 960
rect 1700 960 1740 965
rect 1700 955 1705 960
rect 1625 935 1705 955
rect 1625 930 1630 935
rect 1590 925 1630 930
rect 1700 930 1705 935
rect 1735 955 1740 960
rect 2020 960 2060 965
rect 2020 955 2025 960
rect 1735 935 2025 955
rect 1735 930 1740 935
rect 1700 925 1740 930
rect 2020 930 2025 935
rect 2055 930 2060 960
rect 2020 925 2060 930
rect -180 905 -140 910
rect -180 875 -175 905
rect -145 900 -140 905
rect 230 905 260 910
rect -145 880 230 900
rect -145 875 -140 880
rect -180 870 -140 875
rect 1430 905 1460 910
rect 260 880 1430 900
rect 230 870 260 875
rect 1430 870 1460 875
rect -1080 810 -1040 815
rect -1080 780 -1075 810
rect -1045 805 -1040 810
rect -970 810 -930 815
rect -970 805 -965 810
rect -1045 785 -965 805
rect -1045 780 -1040 785
rect -1080 775 -1040 780
rect -970 780 -965 785
rect -935 805 -930 810
rect -860 810 -820 815
rect -860 805 -855 810
rect -935 785 -855 805
rect -935 780 -930 785
rect -970 775 -930 780
rect -860 780 -855 785
rect -825 805 -820 810
rect -750 810 -710 815
rect -750 805 -745 810
rect -825 785 -745 805
rect -825 780 -820 785
rect -860 775 -820 780
rect -750 780 -745 785
rect -715 805 -710 810
rect -640 810 -600 815
rect -640 805 -635 810
rect -715 785 -635 805
rect -715 780 -710 785
rect -750 775 -710 780
rect -640 780 -635 785
rect -605 805 -600 810
rect -530 810 -490 815
rect -530 805 -525 810
rect -605 785 -525 805
rect -605 780 -600 785
rect -640 775 -600 780
rect -530 780 -525 785
rect -495 780 -490 810
rect -530 775 -490 780
rect 2180 810 2220 815
rect 2180 780 2185 810
rect 2215 805 2220 810
rect 2290 810 2330 815
rect 2290 805 2295 810
rect 2215 785 2295 805
rect 2215 780 2220 785
rect 2180 775 2220 780
rect 2290 780 2295 785
rect 2325 805 2330 810
rect 2400 810 2440 815
rect 2400 805 2405 810
rect 2325 785 2405 805
rect 2325 780 2330 785
rect 2290 775 2330 780
rect 2400 780 2405 785
rect 2435 805 2440 810
rect 2510 810 2550 815
rect 2510 805 2515 810
rect 2435 785 2515 805
rect 2435 780 2440 785
rect 2400 775 2440 780
rect 2510 780 2515 785
rect 2545 805 2550 810
rect 2620 810 2660 815
rect 2620 805 2625 810
rect 2545 785 2625 805
rect 2545 780 2550 785
rect 2510 775 2550 780
rect 2620 780 2625 785
rect 2655 805 2660 810
rect 2730 810 2770 815
rect 2730 805 2735 810
rect 2655 785 2735 805
rect 2655 780 2660 785
rect 2620 775 2660 780
rect 2730 780 2735 785
rect 2765 780 2770 810
rect 2730 775 2770 780
rect -280 770 -240 775
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 755 -1500 760
rect -970 755 -965 760
rect -1505 735 -965 755
rect -1505 730 -1500 735
rect -970 730 -965 735
rect -935 730 -930 760
rect -530 730 -525 760
rect -495 755 -490 760
rect -280 755 -275 770
rect -495 740 -275 755
rect -245 740 -240 770
rect -495 735 -240 740
rect 1930 770 1970 775
rect 1930 740 1935 770
rect 1965 755 1970 770
rect 3190 760 3230 765
rect 2180 755 2185 760
rect 1965 740 2185 755
rect 1930 735 2185 740
rect -495 730 -490 735
rect 2180 730 2185 735
rect 2215 730 2220 760
rect 2620 730 2625 760
rect 2655 755 2660 760
rect 3190 755 3195 760
rect 2655 735 3195 755
rect 2655 730 2660 735
rect 3190 730 3195 735
rect 3225 730 3230 760
rect -1540 725 -1500 730
rect 3190 725 3230 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 710 -1410 715
rect -805 715 -765 720
rect -805 710 -800 715
rect -1415 690 -800 710
rect -1415 685 -1410 690
rect -1450 680 -1410 685
rect -805 685 -800 690
rect -770 710 -765 715
rect -370 715 -330 720
rect -370 710 -365 715
rect -770 690 -365 710
rect -770 685 -765 690
rect -805 680 -765 685
rect -370 685 -365 690
rect -335 685 -330 715
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 710 2060 715
rect 2455 715 2495 720
rect 2455 710 2460 715
rect 2055 690 2460 710
rect 2055 685 2060 690
rect -370 680 -330 685
rect 5 680 45 685
rect -1145 670 -1105 675
rect -1145 640 -1140 670
rect -1110 640 -1105 670
rect -1145 635 -1105 640
rect -1080 670 -1040 675
rect -1080 640 -1075 670
rect -1045 665 -1040 670
rect -970 670 -930 675
rect -970 665 -965 670
rect -1045 645 -965 665
rect -1045 640 -1040 645
rect -1080 635 -1040 640
rect -970 640 -965 645
rect -935 665 -930 670
rect -860 670 -820 675
rect -860 665 -855 670
rect -935 645 -855 665
rect -935 640 -930 645
rect -970 635 -930 640
rect -860 640 -855 645
rect -825 665 -820 670
rect -750 670 -710 675
rect -750 665 -745 670
rect -825 645 -745 665
rect -825 640 -820 645
rect -860 635 -820 640
rect -750 640 -745 645
rect -715 665 -710 670
rect -640 670 -600 675
rect -640 665 -635 670
rect -715 645 -635 665
rect -715 640 -710 645
rect -750 635 -710 640
rect -640 640 -635 645
rect -605 665 -600 670
rect -530 670 -490 675
rect -530 665 -525 670
rect -605 645 -525 665
rect -605 640 -600 645
rect -640 635 -600 640
rect -530 640 -525 645
rect -495 640 -490 670
rect -530 635 -490 640
rect -465 670 -425 675
rect -465 640 -460 670
rect -430 665 -425 670
rect -235 670 -195 675
rect -235 665 -230 670
rect -430 645 -230 665
rect -430 640 -425 645
rect -465 635 -425 640
rect -235 640 -230 645
rect -200 640 -195 670
rect 5 650 10 680
rect 40 675 45 680
rect 115 680 155 685
rect 115 675 120 680
rect 40 655 120 675
rect 40 650 45 655
rect 5 645 45 650
rect 115 650 120 655
rect 150 675 155 680
rect 225 680 265 685
rect 225 675 230 680
rect 150 655 230 675
rect 150 650 155 655
rect 115 645 155 650
rect 225 650 230 655
rect 260 675 265 680
rect 335 680 375 685
rect 335 675 340 680
rect 260 655 340 675
rect 260 650 265 655
rect 225 645 265 650
rect 335 650 340 655
rect 370 675 375 680
rect 445 680 485 685
rect 445 675 450 680
rect 370 655 450 675
rect 370 650 375 655
rect 335 645 375 650
rect 445 650 450 655
rect 480 650 485 680
rect 445 645 485 650
rect 1205 680 1245 685
rect 1205 650 1210 680
rect 1240 675 1245 680
rect 1315 680 1355 685
rect 1315 675 1320 680
rect 1240 655 1320 675
rect 1240 650 1245 655
rect 1205 645 1245 650
rect 1315 650 1320 655
rect 1350 675 1355 680
rect 1425 680 1465 685
rect 1425 675 1430 680
rect 1350 655 1430 675
rect 1350 650 1355 655
rect 1315 645 1355 650
rect 1425 650 1430 655
rect 1460 675 1465 680
rect 1535 680 1575 685
rect 1535 675 1540 680
rect 1460 655 1540 675
rect 1460 650 1465 655
rect 1425 645 1465 650
rect 1535 650 1540 655
rect 1570 675 1575 680
rect 1645 680 1685 685
rect 2020 680 2060 685
rect 2455 685 2460 690
rect 2490 710 2495 715
rect 3100 715 3140 720
rect 3100 710 3105 715
rect 2490 690 3105 710
rect 2490 685 2495 690
rect 2455 680 2495 685
rect 3100 685 3105 690
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 1645 675 1650 680
rect 1570 655 1650 675
rect 1570 650 1575 655
rect 1535 645 1575 650
rect 1645 650 1650 655
rect 1680 650 1685 680
rect 1645 645 1685 650
rect 1885 670 1925 675
rect -235 635 -195 640
rect 1885 640 1890 670
rect 1920 665 1925 670
rect 2115 670 2155 675
rect 2115 665 2120 670
rect 1920 645 2120 665
rect 1920 640 1925 645
rect 1885 635 1925 640
rect 2115 640 2120 645
rect 2150 640 2155 670
rect 2115 635 2155 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 665 2220 670
rect 2290 670 2330 675
rect 2290 665 2295 670
rect 2215 645 2295 665
rect 2215 640 2220 645
rect 2180 635 2220 640
rect 2290 640 2295 645
rect 2325 665 2330 670
rect 2400 670 2440 675
rect 2400 665 2405 670
rect 2325 645 2405 665
rect 2325 640 2330 645
rect 2290 635 2330 640
rect 2400 640 2405 645
rect 2435 665 2440 670
rect 2510 670 2550 675
rect 2510 665 2515 670
rect 2435 645 2515 665
rect 2435 640 2440 645
rect 2400 635 2440 640
rect 2510 640 2515 645
rect 2545 665 2550 670
rect 2620 670 2660 675
rect 2620 665 2625 670
rect 2545 645 2625 665
rect 2545 640 2550 645
rect 2510 635 2550 640
rect 2620 640 2625 645
rect 2655 665 2660 670
rect 2730 670 2770 675
rect 2730 665 2735 670
rect 2655 645 2735 665
rect 2655 640 2660 645
rect 2620 635 2660 640
rect 2730 640 2735 645
rect 2765 640 2770 670
rect 2730 635 2770 640
rect 2795 670 2835 675
rect 2795 640 2800 670
rect 2830 640 2835 670
rect 2795 635 2835 640
rect -105 625 -65 630
rect -105 595 -100 625
rect -70 610 -65 625
rect 555 625 595 630
rect 555 610 560 625
rect -70 595 560 610
rect 590 610 595 625
rect 1095 625 1135 630
rect 1095 610 1100 625
rect 590 605 1100 610
rect 590 595 720 605
rect -105 590 720 595
rect 715 575 720 590
rect 750 590 830 605
rect 750 575 755 590
rect 715 570 755 575
rect 825 575 830 590
rect 860 590 940 605
rect 860 575 865 590
rect 825 570 865 575
rect 935 575 940 590
rect 970 595 1100 605
rect 1130 610 1135 625
rect 1755 625 1795 630
rect 1755 610 1760 625
rect 1130 595 1760 610
rect 1790 620 1795 625
rect 1790 615 1970 620
rect 1790 600 1935 615
rect 1790 595 1795 600
rect 970 590 1795 595
rect 970 575 975 590
rect 1930 585 1935 600
rect 1965 585 1970 615
rect 1930 580 1970 585
rect 935 570 975 575
rect 230 565 260 570
rect -50 555 -10 560
rect -50 525 -45 555
rect -15 550 -10 555
rect 60 555 100 560
rect 60 550 65 555
rect -15 530 65 550
rect -15 525 -10 530
rect -50 520 -10 525
rect 60 525 65 530
rect 95 550 100 555
rect 170 555 210 560
rect 170 550 175 555
rect 95 530 175 550
rect 95 525 100 530
rect 60 520 100 525
rect 170 525 175 530
rect 205 550 210 555
rect 205 535 230 550
rect 1430 565 1460 570
rect 280 555 320 560
rect 280 550 285 555
rect 260 535 285 550
rect 205 530 285 535
rect 205 525 210 530
rect 170 520 210 525
rect 280 525 285 530
rect 315 550 320 555
rect 390 555 430 560
rect 390 550 395 555
rect 315 530 395 550
rect 315 525 320 530
rect 280 520 320 525
rect 390 525 395 530
rect 425 550 430 555
rect 500 555 540 560
rect 500 550 505 555
rect 425 530 505 550
rect 425 525 430 530
rect 390 520 430 525
rect 500 525 505 530
rect 535 525 540 555
rect 500 520 540 525
rect 1150 555 1190 560
rect 1150 525 1155 555
rect 1185 550 1190 555
rect 1260 555 1300 560
rect 1260 550 1265 555
rect 1185 530 1265 550
rect 1185 525 1190 530
rect 1150 520 1190 525
rect 1260 525 1265 530
rect 1295 550 1300 555
rect 1370 555 1410 560
rect 1370 550 1375 555
rect 1295 530 1375 550
rect 1295 525 1300 530
rect 1260 520 1300 525
rect 1370 525 1375 530
rect 1405 550 1410 555
rect 1405 535 1430 550
rect 1480 555 1520 560
rect 1480 550 1485 555
rect 1460 535 1485 550
rect 1405 530 1485 535
rect 1405 525 1410 530
rect 1370 520 1410 525
rect 1480 525 1485 530
rect 1515 550 1520 555
rect 1590 555 1630 560
rect 1590 550 1595 555
rect 1515 530 1595 550
rect 1515 525 1520 530
rect 1480 520 1520 525
rect 1590 525 1595 530
rect 1625 550 1630 555
rect 1700 555 1740 560
rect 1700 550 1705 555
rect 1625 530 1705 550
rect 1625 525 1630 530
rect 1590 520 1630 525
rect 1700 525 1705 530
rect 1735 525 1740 555
rect 1700 520 1740 525
rect 230 505 260 510
rect -105 480 230 500
rect 795 505 825 510
rect 260 480 795 500
rect 230 470 260 475
rect 795 470 825 475
rect 865 505 895 510
rect 1430 505 1460 510
rect 895 480 1430 500
rect 865 470 895 475
rect 1460 480 1795 500
rect 1430 470 1460 475
rect -1270 395 -1230 400
rect -1270 365 -1265 395
rect -1235 390 -1230 395
rect -1025 395 -985 400
rect -1025 390 -1020 395
rect -1235 370 -1020 390
rect -1235 365 -1230 370
rect -1270 360 -1230 365
rect -1025 365 -1020 370
rect -990 390 -985 395
rect -915 395 -875 400
rect -915 390 -910 395
rect -990 370 -910 390
rect -990 365 -985 370
rect -1025 360 -985 365
rect -915 365 -910 370
rect -880 390 -875 395
rect -805 395 -765 400
rect -805 390 -800 395
rect -880 370 -800 390
rect -880 365 -875 370
rect -915 360 -875 365
rect -805 365 -800 370
rect -770 390 -765 395
rect -695 395 -655 400
rect -695 390 -690 395
rect -770 370 -690 390
rect -770 365 -765 370
rect -805 360 -765 365
rect -695 365 -690 370
rect -660 390 -655 395
rect -585 395 -545 400
rect -585 390 -580 395
rect -660 370 -580 390
rect -660 365 -655 370
rect -695 360 -655 365
rect -585 365 -580 370
rect -550 365 -545 395
rect -585 360 -545 365
rect 2235 395 2275 400
rect 2235 365 2240 395
rect 2270 390 2275 395
rect 2345 395 2385 400
rect 2345 390 2350 395
rect 2270 370 2350 390
rect 2270 365 2275 370
rect 2235 360 2275 365
rect 2345 365 2350 370
rect 2380 390 2385 395
rect 2455 395 2495 400
rect 2455 390 2460 395
rect 2380 370 2460 390
rect 2380 365 2385 370
rect 2345 360 2385 365
rect 2455 365 2460 370
rect 2490 390 2495 395
rect 2565 395 2605 400
rect 2565 390 2570 395
rect 2490 370 2570 390
rect 2490 365 2495 370
rect 2455 360 2495 365
rect 2565 365 2570 370
rect 2600 390 2605 395
rect 2675 395 2715 400
rect 2675 390 2680 395
rect 2600 370 2680 390
rect 2600 365 2605 370
rect 2565 360 2605 365
rect 2675 365 2680 370
rect 2710 390 2715 395
rect 2920 395 2960 400
rect 2920 390 2925 395
rect 2710 370 2925 390
rect 2710 365 2715 370
rect 2675 360 2715 365
rect 2920 365 2925 370
rect 2955 365 2960 395
rect 2920 360 2960 365
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect 3185 350 3235 360
rect -1545 310 -1495 320
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 335 -710 340
rect -370 340 -330 345
rect -370 335 -365 340
rect -715 315 -365 335
rect -715 310 -710 315
rect -750 305 -710 310
rect -370 310 -365 315
rect -335 310 -330 340
rect -370 305 -330 310
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 335 2060 340
rect 2400 340 2440 345
rect 2400 335 2405 340
rect 2055 315 2405 335
rect 2055 310 2060 315
rect 2020 305 2060 310
rect 2400 310 2405 315
rect 2435 310 2440 340
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2400 305 2440 310
rect -1225 285 -1185 290
rect -1225 255 -1220 285
rect -1190 280 -1185 285
rect -1025 285 -985 290
rect -1025 280 -1020 285
rect -1190 260 -1020 280
rect -1190 255 -1185 260
rect -1225 250 -1185 255
rect -1025 255 -1020 260
rect -990 280 -985 285
rect -915 285 -875 290
rect -915 280 -910 285
rect -990 260 -910 280
rect -990 255 -985 260
rect -1025 250 -985 255
rect -915 255 -910 260
rect -880 280 -875 285
rect -805 285 -765 290
rect -805 280 -800 285
rect -880 260 -800 280
rect -880 255 -875 260
rect -915 250 -875 255
rect -805 255 -800 260
rect -770 280 -765 285
rect -695 285 -655 290
rect -695 280 -690 285
rect -770 260 -690 280
rect -770 255 -765 260
rect -805 250 -765 255
rect -695 255 -690 260
rect -660 280 -655 285
rect -585 285 -545 290
rect -585 280 -580 285
rect -660 260 -580 280
rect -660 255 -655 260
rect -695 250 -655 255
rect -585 255 -580 260
rect -550 255 -545 285
rect -585 250 -545 255
rect 5 285 45 290
rect 5 255 10 285
rect 40 280 45 285
rect 115 285 155 290
rect 115 280 120 285
rect 40 260 120 280
rect 40 255 45 260
rect 5 250 45 255
rect 115 255 120 260
rect 150 280 155 285
rect 225 285 265 290
rect 225 280 230 285
rect 150 260 230 280
rect 150 255 155 260
rect 115 250 155 255
rect 225 255 230 260
rect 260 280 265 285
rect 335 285 375 290
rect 335 280 340 285
rect 260 260 340 280
rect 260 255 265 260
rect 225 250 265 255
rect 335 255 340 260
rect 370 280 375 285
rect 445 285 485 290
rect 445 280 450 285
rect 370 260 450 280
rect 370 255 375 260
rect 335 250 375 255
rect 445 255 450 260
rect 480 280 485 285
rect 1205 285 1245 290
rect 1205 280 1210 285
rect 480 260 1210 280
rect 480 255 485 260
rect 445 250 485 255
rect 1205 255 1210 260
rect 1240 280 1245 285
rect 1265 285 1295 290
rect 1240 260 1265 280
rect 1240 255 1245 260
rect 1205 250 1245 255
rect 1315 285 1355 290
rect 1315 280 1320 285
rect 1295 260 1320 280
rect 1265 250 1295 255
rect 1315 255 1320 260
rect 1350 280 1355 285
rect 1425 285 1465 290
rect 1425 280 1430 285
rect 1350 260 1430 280
rect 1350 255 1355 260
rect 1315 250 1355 255
rect 1425 255 1430 260
rect 1460 280 1465 285
rect 1535 285 1575 290
rect 1535 280 1540 285
rect 1460 260 1540 280
rect 1460 255 1465 260
rect 1425 250 1465 255
rect 1535 255 1540 260
rect 1570 280 1575 285
rect 1645 285 1685 290
rect 1645 280 1650 285
rect 1570 260 1650 280
rect 1570 255 1575 260
rect 1535 250 1575 255
rect 1645 255 1650 260
rect 1680 255 1685 285
rect 1645 250 1685 255
rect 2235 285 2275 290
rect 2235 255 2240 285
rect 2270 280 2275 285
rect 2345 285 2385 290
rect 2345 280 2350 285
rect 2270 260 2350 280
rect 2270 255 2275 260
rect 2235 250 2275 255
rect 2345 255 2350 260
rect 2380 280 2385 285
rect 2455 285 2495 290
rect 2455 280 2460 285
rect 2380 260 2460 280
rect 2380 255 2385 260
rect 2345 250 2385 255
rect 2455 255 2460 260
rect 2490 280 2495 285
rect 2565 285 2605 290
rect 2565 280 2570 285
rect 2490 260 2570 280
rect 2490 255 2495 260
rect 2455 250 2495 255
rect 2565 255 2570 260
rect 2600 280 2605 285
rect 2675 285 2715 290
rect 2675 280 2680 285
rect 2600 260 2680 280
rect 2600 255 2605 260
rect 2565 250 2605 255
rect 2675 255 2680 260
rect 2710 280 2715 285
rect 2875 285 2915 290
rect 2875 280 2880 285
rect 2710 260 2880 280
rect 2710 255 2715 260
rect 2675 250 2715 255
rect 2875 255 2880 260
rect 2910 255 2915 285
rect 2875 250 2915 255
rect 780 230 820 235
rect 780 200 785 230
rect 815 225 820 230
rect 870 230 910 235
rect 870 225 875 230
rect 815 205 875 225
rect 815 200 820 205
rect 780 195 820 200
rect 870 200 875 205
rect 905 200 910 230
rect 870 195 910 200
rect 855 175 895 180
rect 855 145 860 175
rect 890 145 895 175
rect 855 140 895 145
rect 795 120 835 125
rect 795 90 800 120
rect 830 90 835 120
rect 795 85 835 90
rect 780 65 820 70
rect 780 35 785 65
rect 815 60 820 65
rect 870 65 910 70
rect 870 60 875 65
rect 815 40 875 60
rect 815 35 820 40
rect 780 30 820 35
rect 870 35 875 40
rect 905 35 910 65
rect 870 30 910 35
rect 440 15 480 20
rect 440 -15 445 15
rect 475 10 480 15
rect 830 15 860 20
rect 475 -10 830 10
rect 475 -15 480 -10
rect 440 -20 480 -15
rect 830 -20 860 -15
rect -1490 -120 -1486 -85
rect -1459 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -95 -1275 -85
rect -1225 -90 -1185 -85
rect -1225 -95 -1220 -90
rect -1279 -115 -1220 -95
rect -1279 -120 -1275 -115
rect -1225 -120 -1220 -115
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -1080 -90 -1040 -85
rect -1080 -120 -1075 -90
rect -1045 -95 -1040 -90
rect -970 -90 -930 -85
rect -970 -95 -965 -90
rect -1045 -115 -965 -95
rect -1045 -120 -1040 -115
rect -1080 -125 -1040 -120
rect -970 -120 -965 -115
rect -935 -95 -930 -90
rect -860 -90 -820 -85
rect -860 -95 -855 -90
rect -935 -115 -855 -95
rect -935 -120 -930 -115
rect -970 -125 -930 -120
rect -860 -120 -855 -115
rect -825 -95 -820 -90
rect -750 -90 -710 -85
rect -750 -95 -745 -90
rect -825 -115 -745 -95
rect -825 -120 -820 -115
rect -860 -125 -820 -120
rect -750 -120 -745 -115
rect -715 -95 -710 -90
rect -640 -90 -600 -85
rect -640 -95 -635 -90
rect -715 -115 -635 -95
rect -715 -120 -710 -115
rect -750 -125 -710 -120
rect -640 -120 -635 -115
rect -605 -95 -600 -90
rect -530 -90 -490 -85
rect -530 -95 -525 -90
rect -605 -115 -525 -95
rect -605 -120 -600 -115
rect -640 -125 -600 -120
rect -530 -120 -525 -115
rect -495 -95 -490 -90
rect -235 -90 -195 -85
rect -235 -95 -230 -90
rect -495 -115 -230 -95
rect -495 -120 -490 -115
rect -530 -125 -490 -120
rect -235 -120 -230 -115
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -95 1925 -90
rect 2180 -90 2220 -85
rect 2180 -95 2185 -90
rect 1920 -115 2185 -95
rect 1920 -120 1925 -115
rect 1885 -125 1925 -120
rect 2180 -120 2185 -115
rect 2215 -95 2220 -90
rect 2290 -90 2330 -85
rect 2290 -95 2295 -90
rect 2215 -115 2295 -95
rect 2215 -120 2220 -115
rect 2180 -125 2220 -120
rect 2290 -120 2295 -115
rect 2325 -95 2330 -90
rect 2400 -90 2440 -85
rect 2400 -95 2405 -90
rect 2325 -115 2405 -95
rect 2325 -120 2330 -115
rect 2290 -125 2330 -120
rect 2400 -120 2405 -115
rect 2435 -95 2440 -90
rect 2510 -90 2550 -85
rect 2510 -95 2515 -90
rect 2435 -115 2515 -95
rect 2435 -120 2440 -115
rect 2400 -125 2440 -120
rect 2510 -120 2515 -115
rect 2545 -95 2550 -90
rect 2620 -90 2660 -85
rect 2620 -95 2625 -90
rect 2545 -115 2625 -95
rect 2545 -120 2550 -115
rect 2510 -125 2550 -120
rect 2620 -120 2625 -115
rect 2655 -95 2660 -90
rect 2730 -90 2770 -85
rect 2730 -95 2735 -90
rect 2655 -115 2735 -95
rect 2655 -120 2660 -115
rect 2620 -125 2660 -120
rect 2730 -120 2735 -115
rect 2765 -120 2770 -90
rect 2730 -125 2770 -120
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -95 2915 -90
rect 2965 -95 2969 -85
rect 2910 -115 2969 -95
rect 2910 -120 2915 -115
rect 2965 -120 2969 -115
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3149 -85
rect 3176 -120 3180 -85
rect 2875 -125 2915 -120
rect -1370 -145 -1335 -140
rect -1270 -145 -1230 -140
rect -1270 -150 -1265 -145
rect -1335 -170 -1265 -150
rect -1370 -180 -1335 -175
rect -1270 -175 -1265 -170
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1145 -145 -1105 -140
rect -1145 -175 -1140 -145
rect -1110 -150 -1105 -145
rect -465 -145 -425 -140
rect -465 -150 -460 -145
rect -1110 -170 -460 -150
rect -1110 -175 -1105 -170
rect -1145 -180 -1105 -175
rect -465 -175 -460 -170
rect -430 -150 -425 -145
rect -280 -145 -240 -140
rect -280 -150 -275 -145
rect -430 -170 -275 -150
rect -430 -175 -425 -170
rect -280 -175 -275 -170
rect -245 -175 -240 -145
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -150 1970 -145
rect 2115 -145 2155 -140
rect 2115 -150 2120 -145
rect 1965 -170 2120 -150
rect 1965 -175 1970 -170
rect 2115 -175 2120 -170
rect 2150 -150 2155 -145
rect 2795 -145 2835 -140
rect 2795 -150 2800 -145
rect 2150 -170 2800 -150
rect 2150 -175 2155 -170
rect -465 -180 -425 -175
rect 2115 -180 2155 -175
rect 2795 -175 2800 -170
rect 2830 -175 2835 -145
rect 2795 -180 2835 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -150 2960 -145
rect 3025 -145 3060 -140
rect 2955 -170 3025 -150
rect 2955 -175 2960 -170
rect 2920 -180 2960 -175
rect 3025 -180 3060 -175
rect -1490 -190 -1455 -185
rect 3145 -190 3180 -185
rect -325 -195 -320 -190
rect -1455 -215 -320 -195
rect -1490 -225 -1455 -220
rect -325 -220 -320 -215
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect 1975 -220 1980 -190
rect 2010 -195 2015 -190
rect 2010 -215 3145 -195
rect 2010 -220 2015 -215
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect -1210 -245 -1175 -240
rect -625 -245 -585 -240
rect -625 -250 -620 -245
rect -1175 -270 -620 -250
rect -1210 -280 -1175 -275
rect -625 -275 -620 -270
rect -590 -250 -585 -245
rect -235 -245 -195 -240
rect -235 -250 -230 -245
rect -590 -270 -230 -250
rect -590 -275 -585 -270
rect -625 -280 -585 -275
rect -235 -275 -230 -270
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -250 1925 -245
rect 2275 -245 2315 -240
rect 2275 -250 2280 -245
rect 1920 -270 2280 -250
rect 1920 -275 1925 -270
rect 1885 -280 1925 -275
rect 2275 -275 2280 -270
rect 2310 -250 2315 -245
rect 2865 -245 2900 -240
rect 2310 -270 2865 -250
rect 2310 -275 2315 -270
rect 2275 -280 2315 -275
rect 2865 -280 2900 -275
rect -1540 -300 -1500 -295
rect -1540 -330 -1535 -300
rect -1505 -305 -1500 -300
rect -1150 -300 -1115 -295
rect -1505 -325 -1150 -305
rect -1505 -330 -1500 -325
rect -1540 -335 -1500 -330
rect -925 -300 -885 -295
rect -925 -305 -920 -300
rect -1115 -325 -920 -305
rect -1150 -335 -1115 -330
rect -925 -330 -920 -325
rect -890 -305 -885 -300
rect -725 -300 -685 -295
rect -725 -305 -720 -300
rect -890 -325 -720 -305
rect -890 -330 -885 -325
rect -925 -335 -885 -330
rect -725 -330 -720 -325
rect -690 -305 -685 -300
rect -525 -300 -485 -295
rect -525 -305 -520 -300
rect -690 -325 -520 -305
rect -690 -330 -685 -325
rect -725 -335 -685 -330
rect -525 -330 -520 -325
rect -490 -330 -485 -300
rect 2175 -300 2215 -295
rect -525 -335 -485 -330
rect -105 -310 -65 -305
rect -105 -340 -100 -310
rect -70 -315 -65 -310
rect 595 -310 635 -305
rect 595 -315 600 -310
rect -70 -335 600 -315
rect -70 -340 -65 -335
rect -105 -345 -65 -340
rect 595 -340 600 -335
rect 630 -315 635 -310
rect 715 -310 755 -305
rect 715 -315 720 -310
rect 630 -335 720 -315
rect 630 -340 635 -335
rect 595 -345 635 -340
rect 715 -340 720 -335
rect 750 -315 755 -310
rect 825 -310 865 -305
rect 825 -315 830 -310
rect 750 -335 830 -315
rect 750 -340 755 -335
rect 715 -345 755 -340
rect 825 -340 830 -335
rect 860 -315 865 -310
rect 935 -310 975 -305
rect 935 -315 940 -310
rect 860 -335 940 -315
rect 860 -340 865 -335
rect 825 -345 865 -340
rect 935 -340 940 -335
rect 970 -315 975 -310
rect 1065 -310 1105 -305
rect 1065 -315 1070 -310
rect 970 -335 1070 -315
rect 970 -340 975 -335
rect 935 -345 975 -340
rect 1065 -340 1070 -335
rect 1100 -315 1105 -310
rect 1750 -310 1790 -305
rect 1750 -315 1755 -310
rect 1100 -335 1755 -315
rect 1100 -340 1105 -335
rect 1065 -345 1105 -340
rect 1750 -340 1755 -335
rect 1785 -315 1790 -310
rect 1940 -310 1980 -305
rect 1940 -315 1945 -310
rect 1785 -335 1945 -315
rect 1785 -340 1790 -335
rect 1750 -345 1790 -340
rect 1940 -340 1945 -335
rect 1975 -340 1980 -310
rect 2175 -330 2180 -300
rect 2210 -305 2215 -300
rect 2375 -300 2415 -295
rect 2375 -305 2380 -300
rect 2210 -325 2380 -305
rect 2210 -330 2215 -325
rect 2175 -335 2215 -330
rect 2375 -330 2380 -325
rect 2410 -305 2415 -300
rect 2575 -300 2615 -295
rect 2575 -305 2580 -300
rect 2410 -325 2580 -305
rect 2410 -330 2415 -325
rect 2375 -335 2415 -330
rect 2575 -330 2580 -325
rect 2610 -305 2615 -300
rect 2805 -300 2840 -295
rect 2610 -325 2805 -305
rect 2610 -330 2615 -325
rect 2575 -335 2615 -330
rect 3190 -300 3230 -295
rect 3190 -305 3195 -300
rect 2840 -325 3195 -305
rect 2805 -335 2840 -330
rect 3190 -330 3195 -325
rect 3225 -330 3230 -300
rect 3190 -335 3230 -330
rect 1940 -345 1980 -340
rect -235 -355 -195 -350
rect -1210 -415 -1206 -380
rect -1179 -415 -1175 -380
rect -1150 -415 -1146 -380
rect -1119 -415 -1115 -380
rect -235 -385 -230 -355
rect -200 -360 -195 -355
rect 1885 -355 1925 -350
rect 1885 -360 1890 -355
rect -200 -380 1890 -360
rect -200 -385 -195 -380
rect -235 -390 -195 -385
rect 1885 -385 1890 -380
rect 1920 -385 1925 -355
rect 1885 -390 1925 -385
rect 2805 -415 2809 -380
rect 2836 -415 2840 -380
rect 2865 -415 2869 -380
rect 2896 -415 2900 -380
rect 1335 -425 1375 -420
rect 1335 -455 1340 -425
rect 1370 -430 1375 -425
rect 1840 -425 1880 -420
rect 1840 -430 1845 -425
rect 1370 -450 1845 -430
rect 1370 -455 1375 -450
rect 1335 -460 1375 -455
rect 1840 -455 1845 -450
rect 1875 -455 1880 -425
rect 1840 -460 1880 -455
rect 190 -480 230 -475
rect 190 -510 195 -480
rect 225 -485 230 -480
rect 385 -480 425 -475
rect 385 -485 390 -480
rect 225 -505 390 -485
rect 225 -510 230 -505
rect 190 -515 230 -510
rect 385 -510 390 -505
rect 420 -485 425 -480
rect 495 -480 535 -475
rect 495 -485 500 -480
rect 420 -505 500 -485
rect 420 -510 425 -505
rect 385 -515 425 -510
rect 495 -510 500 -505
rect 530 -485 535 -480
rect 605 -480 645 -475
rect 605 -485 610 -480
rect 530 -505 610 -485
rect 530 -510 535 -505
rect 495 -515 535 -510
rect 605 -510 610 -505
rect 640 -485 645 -480
rect 715 -480 755 -475
rect 715 -485 720 -480
rect 640 -505 720 -485
rect 640 -510 645 -505
rect 605 -515 645 -510
rect 715 -510 720 -505
rect 750 -485 755 -480
rect 825 -480 865 -475
rect 825 -485 830 -480
rect 750 -505 830 -485
rect 750 -510 755 -505
rect 715 -515 755 -510
rect 825 -510 830 -505
rect 860 -485 865 -480
rect 935 -480 975 -475
rect 935 -485 940 -480
rect 860 -505 940 -485
rect 860 -510 865 -505
rect 825 -515 865 -510
rect 935 -510 940 -505
rect 970 -485 975 -480
rect 1045 -480 1085 -475
rect 1045 -485 1050 -480
rect 970 -505 1050 -485
rect 970 -510 975 -505
rect 935 -515 975 -510
rect 1045 -510 1050 -505
rect 1080 -485 1085 -480
rect 1155 -480 1195 -475
rect 1155 -485 1160 -480
rect 1080 -505 1160 -485
rect 1080 -510 1085 -505
rect 1045 -515 1085 -510
rect 1155 -510 1160 -505
rect 1190 -485 1195 -480
rect 1265 -480 1305 -475
rect 1265 -485 1270 -480
rect 1190 -505 1270 -485
rect 1190 -510 1195 -505
rect 1155 -515 1195 -510
rect 1265 -510 1270 -505
rect 1300 -485 1305 -480
rect 1390 -480 1430 -475
rect 1390 -485 1395 -480
rect 1300 -505 1395 -485
rect 1300 -510 1305 -505
rect 1265 -515 1305 -510
rect 1390 -510 1395 -505
rect 1425 -510 1430 -480
rect 1390 -515 1430 -510
rect 265 -805 305 -800
rect 265 -835 270 -805
rect 300 -810 305 -805
rect 330 -805 370 -800
rect 330 -810 335 -805
rect 300 -830 335 -810
rect 300 -835 305 -830
rect 265 -840 305 -835
rect 330 -835 335 -830
rect 365 -810 370 -805
rect 440 -805 480 -800
rect 440 -810 445 -805
rect 365 -830 445 -810
rect 365 -835 370 -830
rect 330 -840 370 -835
rect 440 -835 445 -830
rect 475 -810 480 -805
rect 550 -805 590 -800
rect 550 -810 555 -805
rect 475 -830 555 -810
rect 475 -835 480 -830
rect 440 -840 480 -835
rect 550 -835 555 -830
rect 585 -810 590 -805
rect 660 -805 700 -800
rect 660 -810 665 -805
rect 585 -830 665 -810
rect 585 -835 590 -830
rect 550 -840 590 -835
rect 660 -835 665 -830
rect 695 -810 700 -805
rect 770 -805 810 -800
rect 770 -810 775 -805
rect 695 -830 775 -810
rect 695 -835 700 -830
rect 660 -840 700 -835
rect 770 -835 775 -830
rect 805 -810 810 -805
rect 880 -805 920 -800
rect 880 -810 885 -805
rect 805 -830 885 -810
rect 805 -835 810 -830
rect 770 -840 810 -835
rect 880 -835 885 -830
rect 915 -810 920 -805
rect 990 -805 1030 -800
rect 990 -810 995 -805
rect 915 -830 995 -810
rect 915 -835 920 -830
rect 880 -840 920 -835
rect 990 -835 995 -830
rect 1025 -810 1030 -805
rect 1100 -805 1140 -800
rect 1100 -810 1105 -805
rect 1025 -830 1105 -810
rect 1025 -835 1030 -830
rect 990 -840 1030 -835
rect 1100 -835 1105 -830
rect 1135 -810 1140 -805
rect 1210 -805 1250 -800
rect 1210 -810 1215 -805
rect 1135 -830 1215 -810
rect 1135 -835 1140 -830
rect 1100 -840 1140 -835
rect 1210 -835 1215 -830
rect 1245 -810 1250 -805
rect 1320 -805 1360 -800
rect 1320 -810 1325 -805
rect 1245 -830 1325 -810
rect 1245 -835 1250 -830
rect 1210 -840 1250 -835
rect 1320 -835 1325 -830
rect 1355 -810 1360 -805
rect 1430 -805 1470 -800
rect 1430 -810 1435 -805
rect 1355 -830 1435 -810
rect 1355 -835 1360 -830
rect 1320 -840 1360 -835
rect 1430 -835 1435 -830
rect 1465 -810 1470 -805
rect 1930 -805 1970 -800
rect 1930 -810 1935 -805
rect 1465 -830 1935 -810
rect 1465 -835 1470 -830
rect 1430 -840 1470 -835
rect 1930 -835 1935 -830
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect 190 -855 230 -850
rect 190 -885 195 -855
rect 225 -860 230 -855
rect 225 -865 1355 -860
rect 225 -880 1320 -865
rect 225 -885 230 -880
rect 190 -890 230 -885
rect 1315 -895 1320 -880
rect 1350 -895 1355 -865
rect -190 -900 -150 -895
rect -190 -930 -185 -900
rect -155 -905 -150 -900
rect 550 -900 590 -895
rect 550 -905 555 -900
rect -155 -925 555 -905
rect -155 -930 -150 -925
rect -190 -935 -150 -930
rect 550 -930 555 -925
rect 585 -905 590 -900
rect 660 -900 700 -895
rect 660 -905 665 -900
rect 585 -925 665 -905
rect 585 -930 590 -925
rect 550 -935 590 -930
rect 660 -930 665 -925
rect 695 -905 700 -900
rect 770 -900 810 -895
rect 770 -905 775 -900
rect 695 -925 775 -905
rect 695 -930 700 -925
rect 660 -935 700 -930
rect 770 -930 775 -925
rect 805 -905 810 -900
rect 1005 -900 1045 -895
rect 1005 -905 1010 -900
rect 805 -925 1010 -905
rect 805 -930 810 -925
rect 770 -935 810 -930
rect 1005 -930 1010 -925
rect 1040 -905 1045 -900
rect 1125 -900 1165 -895
rect 1125 -905 1130 -900
rect 1040 -925 1130 -905
rect 1040 -930 1045 -925
rect 1005 -935 1045 -930
rect 1125 -930 1130 -925
rect 1160 -905 1165 -900
rect 1255 -900 1295 -895
rect 1315 -900 1355 -895
rect 1255 -905 1260 -900
rect 1160 -925 1260 -905
rect 1160 -930 1165 -925
rect 1125 -935 1165 -930
rect 1255 -930 1260 -925
rect 1290 -930 1295 -900
rect 1255 -935 1295 -930
rect 925 -1010 965 -1005
rect 925 -1040 930 -1010
rect 960 -1040 965 -1010
rect 925 -1045 965 -1040
rect -1025 -1075 -985 -1070
rect -1025 -1105 -1020 -1075
rect -990 -1080 -985 -1075
rect -825 -1075 -785 -1070
rect -825 -1080 -820 -1075
rect -990 -1100 -820 -1080
rect -990 -1105 -985 -1100
rect -1025 -1110 -985 -1105
rect -825 -1105 -820 -1100
rect -790 -1080 -785 -1075
rect -725 -1075 -685 -1070
rect -725 -1080 -720 -1075
rect -790 -1100 -720 -1080
rect -790 -1105 -785 -1100
rect -825 -1110 -785 -1105
rect -725 -1105 -720 -1100
rect -690 -1080 -685 -1075
rect -625 -1075 -585 -1070
rect -625 -1080 -620 -1075
rect -690 -1100 -620 -1080
rect -690 -1105 -685 -1100
rect -725 -1110 -685 -1105
rect -625 -1105 -620 -1100
rect -590 -1080 -585 -1075
rect -425 -1075 -385 -1070
rect -425 -1080 -420 -1075
rect -590 -1100 -420 -1080
rect -590 -1105 -585 -1100
rect -625 -1110 -585 -1105
rect -425 -1105 -420 -1100
rect -390 -1105 -385 -1075
rect -425 -1110 -385 -1105
rect 2075 -1075 2115 -1070
rect 2075 -1105 2080 -1075
rect 2110 -1080 2115 -1075
rect 2275 -1075 2315 -1070
rect 2275 -1080 2280 -1075
rect 2110 -1100 2280 -1080
rect 2110 -1105 2115 -1100
rect 2075 -1110 2115 -1105
rect 2275 -1105 2280 -1100
rect 2310 -1080 2315 -1075
rect 2375 -1075 2415 -1070
rect 2375 -1080 2380 -1075
rect 2310 -1100 2380 -1080
rect 2310 -1105 2315 -1100
rect 2275 -1110 2315 -1105
rect 2375 -1105 2380 -1100
rect 2410 -1080 2415 -1075
rect 2475 -1075 2515 -1070
rect 2475 -1080 2480 -1075
rect 2410 -1100 2480 -1080
rect 2410 -1105 2415 -1100
rect 2375 -1110 2415 -1105
rect 2475 -1105 2480 -1100
rect 2510 -1080 2515 -1075
rect 2675 -1075 2715 -1070
rect 2675 -1080 2680 -1075
rect 2510 -1100 2680 -1080
rect 2510 -1105 2515 -1100
rect 2475 -1110 2515 -1105
rect 2675 -1105 2680 -1100
rect 2710 -1105 2715 -1075
rect 2675 -1110 2715 -1105
rect 605 -1120 645 -1115
rect 605 -1150 610 -1120
rect 640 -1125 645 -1120
rect 715 -1120 755 -1115
rect 715 -1125 720 -1120
rect 640 -1145 720 -1125
rect 640 -1150 645 -1145
rect 605 -1155 645 -1150
rect 715 -1150 720 -1145
rect 750 -1125 755 -1120
rect 925 -1120 965 -1115
rect 925 -1125 930 -1120
rect 750 -1145 930 -1125
rect 750 -1150 755 -1145
rect 715 -1155 755 -1150
rect 925 -1150 930 -1145
rect 960 -1150 965 -1120
rect 925 -1155 965 -1150
rect -725 -1175 -685 -1170
rect -725 -1205 -720 -1175
rect -690 -1180 -685 -1175
rect -280 -1175 -240 -1170
rect -280 -1180 -275 -1175
rect -690 -1200 -275 -1180
rect -690 -1205 -685 -1200
rect -725 -1210 -685 -1205
rect -280 -1205 -275 -1200
rect -245 -1180 -240 -1175
rect 495 -1175 535 -1170
rect 495 -1180 500 -1175
rect -245 -1200 500 -1180
rect -245 -1205 -240 -1200
rect -280 -1210 -240 -1205
rect 495 -1205 500 -1200
rect 530 -1180 535 -1175
rect 825 -1175 865 -1170
rect 825 -1180 830 -1175
rect 530 -1200 830 -1180
rect 530 -1205 535 -1200
rect 495 -1210 535 -1205
rect 825 -1205 830 -1200
rect 860 -1180 865 -1175
rect 1930 -1175 1970 -1170
rect 1930 -1180 1935 -1175
rect 860 -1200 1935 -1180
rect 860 -1205 865 -1200
rect 825 -1210 865 -1205
rect 1930 -1205 1935 -1200
rect 1965 -1180 1970 -1175
rect 2375 -1175 2415 -1170
rect 2375 -1180 2380 -1175
rect 1965 -1200 2380 -1180
rect 1965 -1205 1970 -1200
rect 1930 -1210 1970 -1205
rect 2375 -1205 2380 -1200
rect 2410 -1205 2415 -1175
rect 2375 -1210 2415 -1205
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via2 >>
rect 830 4245 860 4275
rect -1445 1510 -1415 1540
rect 3105 1460 3135 1490
rect -1535 320 -1505 350
rect 3195 320 3225 350
rect 830 -2455 860 -2425
<< metal3 >>
rect 820 4280 870 4285
rect 820 4240 825 4280
rect 865 4240 870 4280
rect 820 4235 870 4240
rect -3295 3860 -3065 3945
rect -2945 3860 -2715 3945
rect -2595 3860 -2365 3945
rect -3295 3810 -2365 3860
rect -3295 3715 -3065 3810
rect -2945 3715 -2715 3810
rect -2595 3715 -2365 3810
rect -2245 3715 -2015 3945
rect -1895 3715 -1665 3945
rect -1545 3715 -1315 3945
rect -1195 3715 -965 3945
rect -845 3715 -615 3945
rect -495 3715 -265 3945
rect -145 3715 85 3945
rect 205 3715 435 3945
rect 555 3715 785 3945
rect 905 3715 1135 3945
rect 1255 3715 1485 3945
rect 1605 3715 1835 3945
rect 1955 3715 2185 3945
rect 2305 3715 2535 3945
rect 2655 3715 2885 3945
rect 3005 3715 3235 3945
rect 3355 3715 3585 3945
rect 3705 3715 3935 3945
rect 4055 3860 4285 3945
rect 4405 3860 4635 3945
rect 4755 3860 4985 3945
rect 4055 3810 4985 3860
rect 4055 3715 4285 3810
rect 4405 3715 4635 3810
rect 4755 3715 4985 3810
rect -2505 3595 -2455 3715
rect -2155 3595 -2105 3715
rect -1805 3595 -1755 3715
rect -1455 3595 -1405 3715
rect -1105 3595 -1055 3715
rect -755 3595 -705 3715
rect -405 3595 -355 3715
rect -55 3595 -5 3715
rect 295 3595 345 3715
rect 645 3595 695 3715
rect 995 3595 1045 3715
rect 1345 3595 1395 3715
rect 1695 3595 1745 3715
rect 2045 3595 2095 3715
rect 2395 3595 2445 3715
rect 2745 3595 2795 3715
rect 3095 3595 3145 3715
rect 3445 3595 3495 3715
rect 3795 3595 3845 3715
rect 4145 3595 4195 3715
rect -3295 3510 -3065 3595
rect -2945 3510 -2715 3595
rect -2595 3510 -2365 3595
rect -2245 3510 -2015 3595
rect -1895 3510 -1665 3595
rect -1545 3510 -1315 3595
rect -1195 3510 -965 3595
rect -845 3510 -615 3595
rect -495 3510 -265 3595
rect -145 3510 85 3595
rect 205 3510 435 3595
rect 555 3510 785 3595
rect -3295 3460 785 3510
rect -3295 3365 -3065 3460
rect -2945 3365 -2715 3460
rect -2595 3365 -2365 3460
rect -2245 3365 -2015 3460
rect -1895 3365 -1665 3460
rect -1545 3365 -1315 3460
rect -1195 3365 -965 3460
rect -845 3365 -615 3460
rect -495 3365 -265 3460
rect -145 3365 85 3460
rect 205 3365 435 3460
rect 555 3365 785 3460
rect 905 3510 1135 3595
rect 1255 3510 1485 3595
rect 1605 3510 1835 3595
rect 1955 3510 2185 3595
rect 2305 3510 2535 3595
rect 2655 3510 2885 3595
rect 3005 3510 3235 3595
rect 3355 3510 3585 3595
rect 3705 3510 3935 3595
rect 4055 3510 4285 3595
rect 4405 3510 4635 3595
rect 4755 3510 4985 3595
rect 905 3460 4985 3510
rect 905 3365 1135 3460
rect 1255 3365 1485 3460
rect 1605 3365 1835 3460
rect 1955 3365 2185 3460
rect 2305 3365 2535 3460
rect 2655 3365 2885 3460
rect 3005 3365 3235 3460
rect 3355 3365 3585 3460
rect 3705 3365 3935 3460
rect 4055 3365 4285 3460
rect 4405 3365 4635 3460
rect 4755 3365 4985 3460
rect -2505 3245 -2455 3365
rect -1805 3245 -1755 3365
rect -1455 3245 -1405 3365
rect -1105 3245 -1055 3365
rect -755 3245 -705 3365
rect -405 3245 -355 3365
rect -55 3245 -5 3365
rect 295 3245 345 3365
rect 645 3245 695 3365
rect 995 3245 1045 3365
rect 1345 3245 1395 3365
rect 1695 3245 1745 3365
rect 2045 3245 2095 3365
rect 2395 3245 2445 3365
rect 2745 3245 2795 3365
rect 3095 3245 3145 3365
rect 3445 3245 3495 3365
rect 4145 3245 4195 3365
rect -3295 3160 -3065 3245
rect -2945 3160 -2715 3245
rect -2595 3160 -2365 3245
rect -2245 3160 -2015 3245
rect -3295 3110 -2015 3160
rect -3295 3015 -3065 3110
rect -2945 3015 -2715 3110
rect -2595 3015 -2365 3110
rect -2245 3015 -2015 3110
rect -1895 3015 -1665 3245
rect -1545 3015 -1315 3245
rect -1195 3015 -965 3245
rect -845 3015 -615 3245
rect -495 3015 -265 3245
rect -145 3015 85 3245
rect 205 3015 435 3245
rect 555 3015 785 3245
rect 905 3015 1135 3245
rect 1255 3015 1485 3245
rect 1605 3015 1835 3245
rect 1955 3015 2185 3245
rect 2305 3015 2535 3245
rect 2655 3015 2885 3245
rect 3005 3015 3235 3245
rect 3355 3015 3585 3245
rect 3705 3160 3935 3245
rect 4055 3160 4285 3245
rect 4405 3160 4635 3245
rect 4755 3160 4985 3245
rect 3705 3110 4985 3160
rect 3705 3015 3935 3110
rect 4055 3015 4285 3110
rect 4405 3015 4635 3110
rect 4755 3015 4985 3110
rect -2505 2895 -2455 3015
rect -1805 2895 -1755 3015
rect -1455 2895 -1405 3015
rect -1105 2895 -1055 3015
rect -755 2895 -705 3015
rect 2395 2895 2445 3015
rect 2745 2895 2795 3015
rect 3095 2895 3145 3015
rect 3445 2895 3495 3015
rect 4145 2895 4195 3015
rect -3295 2810 -3065 2895
rect -2945 2810 -2715 2895
rect -2595 2810 -2365 2895
rect -2245 2810 -2015 2895
rect -3295 2760 -2015 2810
rect -3295 2665 -3065 2760
rect -2945 2665 -2715 2760
rect -2595 2665 -2365 2760
rect -2245 2665 -2015 2760
rect -1895 2665 -1665 2895
rect -1545 2665 -1315 2895
rect -1195 2665 -965 2895
rect -845 2665 -615 2895
rect 2305 2665 2535 2895
rect 2655 2665 2885 2895
rect 3005 2665 3235 2895
rect 3355 2665 3585 2895
rect 3705 2810 3935 2895
rect 4055 2810 4285 2895
rect 4405 2810 4635 2895
rect 4755 2810 4985 2895
rect 3705 2760 4985 2810
rect 3705 2665 3935 2760
rect 4055 2665 4285 2760
rect 4405 2665 4635 2760
rect 4755 2665 4985 2760
rect -2505 2545 -2455 2665
rect -1455 2545 -1405 2665
rect -1105 2545 -1055 2665
rect -755 2545 -705 2665
rect 2395 2545 2445 2665
rect 2745 2545 2795 2665
rect 3095 2545 3145 2665
rect 4145 2545 4195 2665
rect -3295 2460 -3065 2545
rect -2945 2460 -2715 2545
rect -2595 2460 -2365 2545
rect -2245 2460 -2015 2545
rect -1895 2460 -1665 2545
rect -3295 2410 -1665 2460
rect -3295 2315 -3065 2410
rect -2945 2315 -2715 2410
rect -2595 2315 -2365 2410
rect -2245 2315 -2015 2410
rect -1895 2315 -1665 2410
rect -1545 2315 -1315 2545
rect -1195 2315 -965 2545
rect -845 2315 -615 2545
rect 2305 2315 2535 2545
rect 2655 2315 2885 2545
rect 3005 2315 3235 2545
rect 3355 2460 3585 2545
rect 3705 2460 3935 2545
rect 4055 2460 4285 2545
rect 4405 2460 4635 2545
rect 4755 2460 4985 2545
rect 3355 2410 4985 2460
rect 3355 2315 3585 2410
rect 3705 2315 3935 2410
rect 4055 2315 4285 2410
rect 4405 2315 4635 2410
rect 4755 2315 4985 2410
rect -2505 2195 -2455 2315
rect -3295 2110 -3065 2195
rect -2945 2110 -2715 2195
rect -2595 2110 -2365 2195
rect -2245 2110 -2015 2195
rect -1895 2110 -1665 2195
rect -3295 2060 -1665 2110
rect -3295 1965 -3065 2060
rect -2945 1965 -2715 2060
rect -2595 1965 -2365 2060
rect -2245 1965 -2015 2060
rect -1895 1965 -1665 2060
rect -2505 1845 -2455 1965
rect -3295 1760 -3065 1845
rect -2945 1760 -2715 1845
rect -2595 1760 -2365 1845
rect -2245 1760 -2015 1845
rect -1895 1760 -1665 1845
rect -3295 1710 -1665 1760
rect -3295 1615 -3065 1710
rect -2945 1615 -2715 1710
rect -2595 1615 -2365 1710
rect -2245 1615 -2015 1710
rect -1895 1615 -1665 1710
rect -2505 1495 -2455 1615
rect -1450 1540 -1410 2315
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -3295 1410 -3065 1495
rect -2945 1410 -2715 1495
rect -2595 1410 -2365 1495
rect -2245 1410 -2015 1495
rect -1895 1410 -1665 1495
rect 3100 1490 3140 2315
rect 4145 2195 4195 2315
rect 3355 2110 3585 2195
rect 3705 2110 3935 2195
rect 4055 2110 4285 2195
rect 4405 2110 4635 2195
rect 4755 2110 4985 2195
rect 3355 2060 4985 2110
rect 3355 1965 3585 2060
rect 3705 1965 3935 2060
rect 4055 1965 4285 2060
rect 4405 1965 4635 2060
rect 4755 1965 4985 2060
rect 4145 1845 4195 1965
rect 3355 1760 3585 1845
rect 3705 1760 3935 1845
rect 4055 1760 4285 1845
rect 4405 1760 4635 1845
rect 4755 1760 4985 1845
rect 3355 1710 4985 1760
rect 3355 1615 3585 1710
rect 3705 1615 3935 1710
rect 4055 1615 4285 1710
rect 4405 1615 4635 1710
rect 4755 1615 4985 1710
rect 4145 1495 4195 1615
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect -3295 1360 -1665 1410
rect -3295 1265 -3065 1360
rect -2945 1265 -2715 1360
rect -2595 1265 -2365 1360
rect -2245 1265 -2015 1360
rect -1895 1265 -1665 1360
rect 3355 1410 3585 1495
rect 3705 1410 3935 1495
rect 4055 1410 4285 1495
rect 4405 1410 4635 1495
rect 4755 1410 4985 1495
rect 3355 1360 4985 1410
rect 3355 1265 3585 1360
rect 3705 1265 3935 1360
rect 4055 1265 4285 1360
rect 4405 1265 4635 1360
rect 4755 1265 4985 1360
rect -2505 1145 -2455 1265
rect 4145 1145 4195 1265
rect -3295 1060 -3065 1145
rect -2945 1060 -2715 1145
rect -2595 1060 -2365 1145
rect -2245 1060 -2015 1145
rect -1895 1060 -1665 1145
rect -3295 1010 -1665 1060
rect -3295 915 -3065 1010
rect -2945 915 -2715 1010
rect -2595 915 -2365 1010
rect -2245 915 -2015 1010
rect -1895 915 -1665 1010
rect 3355 1060 3585 1145
rect 3705 1060 3935 1145
rect 4055 1060 4285 1145
rect 4405 1060 4635 1145
rect 4755 1060 4985 1145
rect 3355 1010 4985 1060
rect 3355 915 3585 1010
rect 3705 915 3935 1010
rect 4055 915 4285 1010
rect 4405 915 4635 1010
rect 4755 915 4985 1010
rect -2505 795 -2455 915
rect 4145 795 4195 915
rect -3295 710 -3065 795
rect -2945 710 -2715 795
rect -2595 710 -2365 795
rect -2245 710 -2015 795
rect -1895 710 -1665 795
rect -3295 660 -1665 710
rect -3295 565 -3065 660
rect -2945 565 -2715 660
rect -2595 565 -2365 660
rect -2245 565 -2015 660
rect -1895 565 -1665 660
rect 3355 710 3585 795
rect 3705 710 3935 795
rect 4055 710 4285 795
rect 4405 710 4635 795
rect 4755 710 4985 795
rect 3355 660 4985 710
rect 3355 565 3585 660
rect 3705 565 3935 660
rect 4055 565 4285 660
rect 4405 565 4635 660
rect 4755 565 4985 660
rect -2505 445 -2455 565
rect 4145 445 4195 565
rect -3295 360 -3065 445
rect -2945 360 -2715 445
rect -2595 360 -2365 445
rect -2245 360 -2015 445
rect -1895 360 -1665 445
rect 3355 360 3585 445
rect 3705 360 3935 445
rect 4055 360 4285 445
rect 4405 360 4635 445
rect 4755 360 4985 445
rect -3295 310 -1665 360
rect -1545 355 -1495 360
rect -1545 315 -1540 355
rect -1500 315 -1495 355
rect -1545 310 -1495 315
rect 3185 355 3235 360
rect 3185 315 3190 355
rect 3230 315 3235 355
rect 3185 310 3235 315
rect 3355 310 4985 360
rect -3295 215 -3065 310
rect -2945 215 -2715 310
rect -2595 215 -2365 310
rect -2245 215 -2015 310
rect -1895 215 -1665 310
rect 3355 215 3585 310
rect 3705 215 3935 310
rect 4055 215 4285 310
rect 4405 215 4635 310
rect 4755 215 4985 310
rect -2505 95 -2455 215
rect 4145 95 4195 215
rect -3295 10 -3065 95
rect -2945 10 -2715 95
rect -2595 10 -2365 95
rect -2245 10 -2015 95
rect -1895 10 -1665 95
rect -3295 -40 -1665 10
rect -3295 -135 -3065 -40
rect -2945 -135 -2715 -40
rect -2595 -135 -2365 -40
rect -2245 -135 -2015 -40
rect -1895 -135 -1665 -40
rect 3355 10 3585 95
rect 3705 10 3935 95
rect 4055 10 4285 95
rect 4405 10 4635 95
rect 4755 10 4985 95
rect 3355 -40 4985 10
rect 3355 -135 3585 -40
rect 3705 -135 3935 -40
rect 4055 -135 4285 -40
rect 4405 -135 4635 -40
rect 4755 -135 4985 -40
rect -2505 -255 -2455 -135
rect 4145 -255 4195 -135
rect -3295 -340 -3065 -255
rect -2945 -340 -2715 -255
rect -2595 -340 -2365 -255
rect -2245 -340 -2015 -255
rect -1895 -340 -1665 -255
rect -3295 -390 -1665 -340
rect -3295 -485 -3065 -390
rect -2945 -485 -2715 -390
rect -2595 -485 -2365 -390
rect -2245 -485 -2015 -390
rect -1895 -485 -1665 -390
rect 3355 -340 3585 -255
rect 3705 -340 3935 -255
rect 4055 -340 4285 -255
rect 4405 -340 4635 -255
rect 4755 -340 4985 -255
rect 3355 -390 4985 -340
rect 3355 -485 3585 -390
rect 3705 -485 3935 -390
rect 4055 -485 4285 -390
rect 4405 -485 4635 -390
rect 4755 -485 4985 -390
rect -2505 -605 -2455 -485
rect 4145 -605 4195 -485
rect -3295 -690 -3065 -605
rect -2945 -690 -2715 -605
rect -2595 -690 -2365 -605
rect -2245 -690 -2015 -605
rect -1895 -690 -1665 -605
rect -3295 -740 -1665 -690
rect -3295 -835 -3065 -740
rect -2945 -835 -2715 -740
rect -2595 -835 -2365 -740
rect -2245 -835 -2015 -740
rect -1895 -835 -1665 -740
rect 3355 -690 3585 -605
rect 3705 -690 3935 -605
rect 4055 -690 4285 -605
rect 4405 -690 4635 -605
rect 4755 -690 4985 -605
rect 3355 -740 4985 -690
rect 3355 -835 3585 -740
rect 3705 -835 3935 -740
rect 4055 -835 4285 -740
rect 4405 -835 4635 -740
rect 4755 -835 4985 -740
rect -2505 -955 -2455 -835
rect 4145 -955 4195 -835
rect -3295 -1040 -3065 -955
rect -2945 -1040 -2715 -955
rect -2595 -1040 -2365 -955
rect -2245 -1040 -2015 -955
rect -1895 -1040 -1665 -955
rect -3295 -1090 -1665 -1040
rect -3295 -1185 -3065 -1090
rect -2945 -1185 -2715 -1090
rect -2595 -1185 -2365 -1090
rect -2245 -1185 -2015 -1090
rect -1895 -1185 -1665 -1090
rect 3355 -1040 3585 -955
rect 3705 -1040 3935 -955
rect 4055 -1040 4285 -955
rect 4405 -1040 4635 -955
rect 4755 -1040 4985 -955
rect 3355 -1090 4985 -1040
rect 3355 -1185 3585 -1090
rect 3705 -1185 3935 -1090
rect 4055 -1185 4285 -1090
rect 4405 -1185 4635 -1090
rect 4755 -1185 4985 -1090
rect -2505 -1305 -2455 -1185
rect 4145 -1305 4195 -1185
rect -3295 -1390 -3065 -1305
rect -2945 -1390 -2715 -1305
rect -2595 -1390 -2365 -1305
rect -2245 -1390 -2015 -1305
rect -1895 -1390 -1665 -1305
rect -3295 -1440 -1665 -1390
rect -3295 -1535 -3065 -1440
rect -2945 -1535 -2715 -1440
rect -2595 -1535 -2365 -1440
rect -2245 -1535 -2015 -1440
rect -1895 -1535 -1665 -1440
rect -1545 -1535 -1315 -1305
rect -1195 -1535 -965 -1305
rect -845 -1535 -615 -1305
rect -495 -1535 -265 -1305
rect -145 -1535 85 -1305
rect 205 -1535 435 -1305
rect 555 -1535 785 -1305
rect 905 -1535 1135 -1305
rect 1255 -1535 1485 -1305
rect 1605 -1535 1835 -1305
rect 1955 -1535 2185 -1305
rect 2305 -1535 2535 -1305
rect 2655 -1535 2885 -1305
rect 3005 -1535 3235 -1305
rect 3355 -1390 3585 -1305
rect 3705 -1390 3935 -1305
rect 4055 -1390 4285 -1305
rect 4405 -1390 4635 -1305
rect 4755 -1390 4985 -1305
rect 3355 -1440 4985 -1390
rect 3355 -1535 3585 -1440
rect 3705 -1535 3935 -1440
rect 4055 -1535 4285 -1440
rect 4405 -1535 4635 -1440
rect 4755 -1535 4985 -1440
rect -2505 -1655 -2455 -1535
rect -1455 -1655 -1405 -1535
rect -1105 -1655 -1055 -1535
rect -755 -1655 -705 -1535
rect -405 -1655 -355 -1535
rect -55 -1655 -5 -1535
rect 295 -1655 345 -1535
rect 645 -1655 695 -1535
rect 995 -1655 1045 -1535
rect 1345 -1655 1395 -1535
rect 1695 -1655 1745 -1535
rect 2045 -1655 2095 -1535
rect 2395 -1655 2445 -1535
rect 2745 -1655 2795 -1535
rect 3095 -1655 3145 -1535
rect 4145 -1655 4195 -1535
rect -3295 -1740 -3065 -1655
rect -2945 -1740 -2715 -1655
rect -2595 -1740 -2365 -1655
rect -2245 -1740 -2015 -1655
rect -1895 -1740 -1665 -1655
rect -1545 -1740 -1315 -1655
rect -1195 -1740 -965 -1655
rect -845 -1740 -615 -1655
rect -495 -1740 -265 -1655
rect -145 -1740 85 -1655
rect 205 -1740 435 -1655
rect 555 -1740 785 -1655
rect -3295 -1790 785 -1740
rect -3295 -1885 -3065 -1790
rect -2945 -1885 -2715 -1790
rect -2595 -1885 -2365 -1790
rect -2245 -1885 -2015 -1790
rect -1895 -1885 -1665 -1790
rect -1545 -1885 -1315 -1790
rect -1195 -1885 -965 -1790
rect -845 -1885 -615 -1790
rect -495 -1885 -265 -1790
rect -145 -1885 85 -1790
rect 205 -1885 435 -1790
rect 555 -1885 785 -1790
rect 905 -1740 1135 -1655
rect 1255 -1740 1485 -1655
rect 1605 -1740 1835 -1655
rect 1955 -1740 2185 -1655
rect 2305 -1740 2535 -1655
rect 2655 -1740 2885 -1655
rect 3005 -1740 3235 -1655
rect 3355 -1740 3585 -1655
rect 3705 -1740 3935 -1655
rect 4055 -1740 4285 -1655
rect 4405 -1740 4635 -1655
rect 4755 -1740 4985 -1655
rect 905 -1790 4985 -1740
rect 905 -1885 1135 -1790
rect 1255 -1885 1485 -1790
rect 1605 -1885 1835 -1790
rect 1955 -1885 2185 -1790
rect 2305 -1885 2535 -1790
rect 2655 -1885 2885 -1790
rect 3005 -1885 3235 -1790
rect 3355 -1885 3585 -1790
rect 3705 -1885 3935 -1790
rect 4055 -1885 4285 -1790
rect 4405 -1885 4635 -1790
rect 4755 -1885 4985 -1790
rect -2505 -2005 -2455 -1885
rect -2155 -2005 -2105 -1885
rect -1805 -2005 -1755 -1885
rect -1455 -2005 -1405 -1885
rect -1105 -2005 -1055 -1885
rect -755 -2005 -705 -1885
rect -405 -2005 -355 -1885
rect -55 -2005 -5 -1885
rect 295 -2005 345 -1885
rect 645 -2005 695 -1885
rect 995 -2005 1045 -1885
rect 1345 -2005 1395 -1885
rect 1695 -2005 1745 -1885
rect 2045 -2005 2095 -1885
rect 2395 -2005 2445 -1885
rect 2745 -2005 2795 -1885
rect 3095 -2005 3145 -1885
rect 3445 -2005 3495 -1885
rect 3795 -2005 3845 -1885
rect 4145 -2005 4195 -1885
rect -3295 -2090 -3065 -2005
rect -2945 -2090 -2715 -2005
rect -2595 -2090 -2365 -2005
rect -3295 -2140 -2365 -2090
rect -3295 -2235 -3065 -2140
rect -2945 -2235 -2715 -2140
rect -2595 -2235 -2365 -2140
rect -2245 -2235 -2015 -2005
rect -1895 -2235 -1665 -2005
rect -1545 -2235 -1315 -2005
rect -1195 -2235 -965 -2005
rect -845 -2235 -615 -2005
rect -495 -2235 -265 -2005
rect -145 -2235 85 -2005
rect 205 -2235 435 -2005
rect 555 -2235 785 -2005
rect 905 -2235 1135 -2005
rect 1255 -2235 1485 -2005
rect 1605 -2235 1835 -2005
rect 1955 -2235 2185 -2005
rect 2305 -2235 2535 -2005
rect 2655 -2235 2885 -2005
rect 3005 -2235 3235 -2005
rect 3355 -2235 3585 -2005
rect 3705 -2235 3935 -2005
rect 4055 -2090 4285 -2005
rect 4405 -2090 4635 -2005
rect 4755 -2090 4985 -2005
rect 4055 -2140 4985 -2090
rect 4055 -2235 4285 -2140
rect 4405 -2235 4635 -2140
rect 4755 -2235 4985 -2140
rect 820 -2420 870 -2415
rect 820 -2460 825 -2420
rect 865 -2460 870 -2420
rect 820 -2465 870 -2460
<< via3 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 830 4245 860 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect -1540 350 -1500 355
rect -1540 320 -1535 350
rect -1535 320 -1505 350
rect -1505 320 -1500 350
rect -1540 315 -1500 320
rect 3190 350 3230 355
rect 3190 320 3195 350
rect 3195 320 3225 350
rect 3225 320 3230 350
rect 3190 315 3230 320
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 830 -2455 860 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< mimcap >>
rect -3280 3855 -3080 3930
rect -3280 3815 -3200 3855
rect -3160 3815 -3080 3855
rect -3280 3730 -3080 3815
rect -2930 3855 -2730 3930
rect -2930 3815 -2850 3855
rect -2810 3815 -2730 3855
rect -2930 3730 -2730 3815
rect -2580 3855 -2380 3930
rect -2580 3815 -2500 3855
rect -2460 3815 -2380 3855
rect -2580 3730 -2380 3815
rect -2230 3855 -2030 3930
rect -2230 3815 -2150 3855
rect -2110 3815 -2030 3855
rect -2230 3730 -2030 3815
rect -1880 3855 -1680 3930
rect -1880 3815 -1800 3855
rect -1760 3815 -1680 3855
rect -1880 3730 -1680 3815
rect -1530 3855 -1330 3930
rect -1530 3815 -1450 3855
rect -1410 3815 -1330 3855
rect -1530 3730 -1330 3815
rect -1180 3855 -980 3930
rect -1180 3815 -1100 3855
rect -1060 3815 -980 3855
rect -1180 3730 -980 3815
rect -830 3855 -630 3930
rect -830 3815 -750 3855
rect -710 3815 -630 3855
rect -830 3730 -630 3815
rect -480 3855 -280 3930
rect -480 3815 -400 3855
rect -360 3815 -280 3855
rect -480 3730 -280 3815
rect -130 3855 70 3930
rect -130 3815 -50 3855
rect -10 3815 70 3855
rect -130 3730 70 3815
rect 220 3855 420 3930
rect 220 3815 300 3855
rect 340 3815 420 3855
rect 220 3730 420 3815
rect 570 3855 770 3930
rect 570 3815 650 3855
rect 690 3815 770 3855
rect 570 3730 770 3815
rect 920 3855 1120 3930
rect 920 3815 1000 3855
rect 1040 3815 1120 3855
rect 920 3730 1120 3815
rect 1270 3855 1470 3930
rect 1270 3815 1350 3855
rect 1390 3815 1470 3855
rect 1270 3730 1470 3815
rect 1620 3855 1820 3930
rect 1620 3815 1700 3855
rect 1740 3815 1820 3855
rect 1620 3730 1820 3815
rect 1970 3855 2170 3930
rect 1970 3815 2050 3855
rect 2090 3815 2170 3855
rect 1970 3730 2170 3815
rect 2320 3855 2520 3930
rect 2320 3815 2400 3855
rect 2440 3815 2520 3855
rect 2320 3730 2520 3815
rect 2670 3855 2870 3930
rect 2670 3815 2750 3855
rect 2790 3815 2870 3855
rect 2670 3730 2870 3815
rect 3020 3855 3220 3930
rect 3020 3815 3100 3855
rect 3140 3815 3220 3855
rect 3020 3730 3220 3815
rect 3370 3855 3570 3930
rect 3370 3815 3450 3855
rect 3490 3815 3570 3855
rect 3370 3730 3570 3815
rect 3720 3855 3920 3930
rect 3720 3815 3800 3855
rect 3840 3815 3920 3855
rect 3720 3730 3920 3815
rect 4070 3855 4270 3930
rect 4070 3815 4150 3855
rect 4190 3815 4270 3855
rect 4070 3730 4270 3815
rect 4420 3855 4620 3930
rect 4420 3815 4500 3855
rect 4540 3815 4620 3855
rect 4420 3730 4620 3815
rect 4770 3855 4970 3930
rect 4770 3815 4850 3855
rect 4890 3815 4970 3855
rect 4770 3730 4970 3815
rect -3280 3505 -3080 3580
rect -3280 3465 -3200 3505
rect -3160 3465 -3080 3505
rect -3280 3380 -3080 3465
rect -2930 3505 -2730 3580
rect -2930 3465 -2850 3505
rect -2810 3465 -2730 3505
rect -2930 3380 -2730 3465
rect -2580 3505 -2380 3580
rect -2580 3465 -2500 3505
rect -2460 3465 -2380 3505
rect -2580 3380 -2380 3465
rect -2230 3505 -2030 3580
rect -2230 3465 -2150 3505
rect -2110 3465 -2030 3505
rect -2230 3380 -2030 3465
rect -1880 3505 -1680 3580
rect -1880 3465 -1800 3505
rect -1760 3465 -1680 3505
rect -1880 3380 -1680 3465
rect -1530 3505 -1330 3580
rect -1530 3465 -1450 3505
rect -1410 3465 -1330 3505
rect -1530 3380 -1330 3465
rect -1180 3505 -980 3580
rect -1180 3465 -1100 3505
rect -1060 3465 -980 3505
rect -1180 3380 -980 3465
rect -830 3505 -630 3580
rect -830 3465 -750 3505
rect -710 3465 -630 3505
rect -830 3380 -630 3465
rect -480 3505 -280 3580
rect -480 3465 -400 3505
rect -360 3465 -280 3505
rect -480 3380 -280 3465
rect -130 3505 70 3580
rect -130 3465 -50 3505
rect -10 3465 70 3505
rect -130 3380 70 3465
rect 220 3505 420 3580
rect 220 3465 300 3505
rect 340 3465 420 3505
rect 220 3380 420 3465
rect 570 3505 770 3580
rect 570 3465 650 3505
rect 690 3465 770 3505
rect 570 3380 770 3465
rect 920 3505 1120 3580
rect 920 3465 1000 3505
rect 1040 3465 1120 3505
rect 920 3380 1120 3465
rect 1270 3505 1470 3580
rect 1270 3465 1350 3505
rect 1390 3465 1470 3505
rect 1270 3380 1470 3465
rect 1620 3505 1820 3580
rect 1620 3465 1700 3505
rect 1740 3465 1820 3505
rect 1620 3380 1820 3465
rect 1970 3505 2170 3580
rect 1970 3465 2050 3505
rect 2090 3465 2170 3505
rect 1970 3380 2170 3465
rect 2320 3505 2520 3580
rect 2320 3465 2400 3505
rect 2440 3465 2520 3505
rect 2320 3380 2520 3465
rect 2670 3505 2870 3580
rect 2670 3465 2750 3505
rect 2790 3465 2870 3505
rect 2670 3380 2870 3465
rect 3020 3505 3220 3580
rect 3020 3465 3100 3505
rect 3140 3465 3220 3505
rect 3020 3380 3220 3465
rect 3370 3505 3570 3580
rect 3370 3465 3450 3505
rect 3490 3465 3570 3505
rect 3370 3380 3570 3465
rect 3720 3505 3920 3580
rect 3720 3465 3800 3505
rect 3840 3465 3920 3505
rect 3720 3380 3920 3465
rect 4070 3505 4270 3580
rect 4070 3465 4150 3505
rect 4190 3465 4270 3505
rect 4070 3380 4270 3465
rect 4420 3505 4620 3580
rect 4420 3465 4500 3505
rect 4540 3465 4620 3505
rect 4420 3380 4620 3465
rect 4770 3505 4970 3580
rect 4770 3465 4850 3505
rect 4890 3465 4970 3505
rect 4770 3380 4970 3465
rect -3280 3155 -3080 3230
rect -3280 3115 -3200 3155
rect -3160 3115 -3080 3155
rect -3280 3030 -3080 3115
rect -2930 3155 -2730 3230
rect -2930 3115 -2850 3155
rect -2810 3115 -2730 3155
rect -2930 3030 -2730 3115
rect -2580 3155 -2380 3230
rect -2580 3115 -2500 3155
rect -2460 3115 -2380 3155
rect -2580 3030 -2380 3115
rect -2230 3155 -2030 3230
rect -2230 3115 -2150 3155
rect -2110 3115 -2030 3155
rect -2230 3030 -2030 3115
rect -1880 3155 -1680 3230
rect -1880 3115 -1800 3155
rect -1760 3115 -1680 3155
rect -1880 3030 -1680 3115
rect -1530 3155 -1330 3230
rect -1530 3115 -1450 3155
rect -1410 3115 -1330 3155
rect -1530 3030 -1330 3115
rect -1180 3155 -980 3230
rect -1180 3115 -1100 3155
rect -1060 3115 -980 3155
rect -1180 3030 -980 3115
rect -830 3155 -630 3230
rect -830 3115 -750 3155
rect -710 3115 -630 3155
rect -830 3030 -630 3115
rect -480 3155 -280 3230
rect -480 3115 -400 3155
rect -360 3115 -280 3155
rect -480 3030 -280 3115
rect -130 3145 70 3230
rect -130 3105 -50 3145
rect -10 3105 70 3145
rect -130 3030 70 3105
rect 220 3145 420 3230
rect 220 3105 300 3145
rect 340 3105 420 3145
rect 220 3030 420 3105
rect 570 3145 770 3230
rect 570 3105 650 3145
rect 690 3105 770 3145
rect 570 3030 770 3105
rect 920 3145 1120 3230
rect 920 3105 1000 3145
rect 1040 3105 1120 3145
rect 920 3030 1120 3105
rect 1270 3145 1470 3230
rect 1270 3105 1350 3145
rect 1390 3105 1470 3145
rect 1270 3030 1470 3105
rect 1620 3145 1820 3230
rect 1620 3105 1700 3145
rect 1740 3105 1820 3145
rect 1620 3030 1820 3105
rect 1970 3155 2170 3230
rect 1970 3115 2050 3155
rect 2090 3115 2170 3155
rect 1970 3030 2170 3115
rect 2320 3155 2520 3230
rect 2320 3115 2400 3155
rect 2440 3115 2520 3155
rect 2320 3030 2520 3115
rect 2670 3155 2870 3230
rect 2670 3115 2750 3155
rect 2790 3115 2870 3155
rect 2670 3030 2870 3115
rect 3020 3155 3220 3230
rect 3020 3115 3100 3155
rect 3140 3115 3220 3155
rect 3020 3030 3220 3115
rect 3370 3155 3570 3230
rect 3370 3115 3450 3155
rect 3490 3115 3570 3155
rect 3370 3030 3570 3115
rect 3720 3155 3920 3230
rect 3720 3115 3800 3155
rect 3840 3115 3920 3155
rect 3720 3030 3920 3115
rect 4070 3155 4270 3230
rect 4070 3115 4150 3155
rect 4190 3115 4270 3155
rect 4070 3030 4270 3115
rect 4420 3155 4620 3230
rect 4420 3115 4500 3155
rect 4540 3115 4620 3155
rect 4420 3030 4620 3115
rect 4770 3155 4970 3230
rect 4770 3115 4850 3155
rect 4890 3115 4970 3155
rect 4770 3030 4970 3115
rect -3280 2805 -3080 2880
rect -3280 2765 -3200 2805
rect -3160 2765 -3080 2805
rect -3280 2680 -3080 2765
rect -2930 2805 -2730 2880
rect -2930 2765 -2850 2805
rect -2810 2765 -2730 2805
rect -2930 2680 -2730 2765
rect -2580 2805 -2380 2880
rect -2580 2765 -2500 2805
rect -2460 2765 -2380 2805
rect -2580 2680 -2380 2765
rect -2230 2805 -2030 2880
rect -2230 2765 -2150 2805
rect -2110 2765 -2030 2805
rect -2230 2680 -2030 2765
rect -1880 2805 -1680 2880
rect -1880 2765 -1800 2805
rect -1760 2765 -1680 2805
rect -1880 2680 -1680 2765
rect -1530 2805 -1330 2880
rect -1530 2765 -1450 2805
rect -1410 2765 -1330 2805
rect -1530 2680 -1330 2765
rect -1180 2805 -980 2880
rect -1180 2765 -1100 2805
rect -1060 2765 -980 2805
rect -1180 2680 -980 2765
rect -830 2805 -630 2880
rect -830 2765 -750 2805
rect -710 2765 -630 2805
rect -830 2680 -630 2765
rect 2320 2805 2520 2880
rect 2320 2765 2400 2805
rect 2440 2765 2520 2805
rect 2320 2680 2520 2765
rect 2670 2805 2870 2880
rect 2670 2765 2750 2805
rect 2790 2765 2870 2805
rect 2670 2680 2870 2765
rect 3020 2805 3220 2880
rect 3020 2765 3100 2805
rect 3140 2765 3220 2805
rect 3020 2680 3220 2765
rect 3370 2805 3570 2880
rect 3370 2765 3450 2805
rect 3490 2765 3570 2805
rect 3370 2680 3570 2765
rect 3720 2805 3920 2880
rect 3720 2765 3800 2805
rect 3840 2765 3920 2805
rect 3720 2680 3920 2765
rect 4070 2805 4270 2880
rect 4070 2765 4150 2805
rect 4190 2765 4270 2805
rect 4070 2680 4270 2765
rect 4420 2805 4620 2880
rect 4420 2765 4500 2805
rect 4540 2765 4620 2805
rect 4420 2680 4620 2765
rect 4770 2805 4970 2880
rect 4770 2765 4850 2805
rect 4890 2765 4970 2805
rect 4770 2680 4970 2765
rect -3280 2455 -3080 2530
rect -3280 2415 -3200 2455
rect -3160 2415 -3080 2455
rect -3280 2330 -3080 2415
rect -2930 2455 -2730 2530
rect -2930 2415 -2850 2455
rect -2810 2415 -2730 2455
rect -2930 2330 -2730 2415
rect -2580 2455 -2380 2530
rect -2580 2415 -2500 2455
rect -2460 2415 -2380 2455
rect -2580 2330 -2380 2415
rect -2230 2455 -2030 2530
rect -2230 2415 -2150 2455
rect -2110 2415 -2030 2455
rect -2230 2330 -2030 2415
rect -1880 2455 -1680 2530
rect -1880 2415 -1800 2455
rect -1760 2415 -1680 2455
rect -1880 2330 -1680 2415
rect -1530 2455 -1330 2530
rect -1530 2415 -1450 2455
rect -1410 2415 -1330 2455
rect -1530 2330 -1330 2415
rect -1180 2455 -980 2530
rect -1180 2415 -1100 2455
rect -1060 2415 -980 2455
rect -1180 2330 -980 2415
rect -830 2455 -630 2530
rect -830 2415 -750 2455
rect -710 2415 -630 2455
rect -830 2330 -630 2415
rect 2320 2455 2520 2530
rect 2320 2415 2400 2455
rect 2440 2415 2520 2455
rect 2320 2330 2520 2415
rect 2670 2455 2870 2530
rect 2670 2415 2750 2455
rect 2790 2415 2870 2455
rect 2670 2330 2870 2415
rect 3020 2455 3220 2530
rect 3020 2415 3100 2455
rect 3140 2415 3220 2455
rect 3020 2330 3220 2415
rect 3370 2455 3570 2530
rect 3370 2415 3450 2455
rect 3490 2415 3570 2455
rect 3370 2330 3570 2415
rect 3720 2455 3920 2530
rect 3720 2415 3800 2455
rect 3840 2415 3920 2455
rect 3720 2330 3920 2415
rect 4070 2455 4270 2530
rect 4070 2415 4150 2455
rect 4190 2415 4270 2455
rect 4070 2330 4270 2415
rect 4420 2455 4620 2530
rect 4420 2415 4500 2455
rect 4540 2415 4620 2455
rect 4420 2330 4620 2415
rect 4770 2455 4970 2530
rect 4770 2415 4850 2455
rect 4890 2415 4970 2455
rect 4770 2330 4970 2415
rect -3280 2105 -3080 2180
rect -3280 2065 -3200 2105
rect -3160 2065 -3080 2105
rect -3280 1980 -3080 2065
rect -2930 2105 -2730 2180
rect -2930 2065 -2850 2105
rect -2810 2065 -2730 2105
rect -2930 1980 -2730 2065
rect -2580 2105 -2380 2180
rect -2580 2065 -2500 2105
rect -2460 2065 -2380 2105
rect -2580 1980 -2380 2065
rect -2230 2105 -2030 2180
rect -2230 2065 -2150 2105
rect -2110 2065 -2030 2105
rect -2230 1980 -2030 2065
rect -1880 2105 -1680 2180
rect -1880 2065 -1800 2105
rect -1760 2065 -1680 2105
rect -1880 1980 -1680 2065
rect 3370 2105 3570 2180
rect 3370 2065 3450 2105
rect 3490 2065 3570 2105
rect 3370 1980 3570 2065
rect 3720 2105 3920 2180
rect 3720 2065 3800 2105
rect 3840 2065 3920 2105
rect 3720 1980 3920 2065
rect 4070 2105 4270 2180
rect 4070 2065 4150 2105
rect 4190 2065 4270 2105
rect 4070 1980 4270 2065
rect 4420 2105 4620 2180
rect 4420 2065 4500 2105
rect 4540 2065 4620 2105
rect 4420 1980 4620 2065
rect 4770 2105 4970 2180
rect 4770 2065 4850 2105
rect 4890 2065 4970 2105
rect 4770 1980 4970 2065
rect -3280 1755 -3080 1830
rect -3280 1715 -3200 1755
rect -3160 1715 -3080 1755
rect -3280 1630 -3080 1715
rect -2930 1755 -2730 1830
rect -2930 1715 -2850 1755
rect -2810 1715 -2730 1755
rect -2930 1630 -2730 1715
rect -2580 1755 -2380 1830
rect -2580 1715 -2500 1755
rect -2460 1715 -2380 1755
rect -2580 1630 -2380 1715
rect -2230 1755 -2030 1830
rect -2230 1715 -2150 1755
rect -2110 1715 -2030 1755
rect -2230 1630 -2030 1715
rect -1880 1755 -1680 1830
rect -1880 1715 -1800 1755
rect -1760 1715 -1680 1755
rect -1880 1630 -1680 1715
rect 3370 1755 3570 1830
rect 3370 1715 3450 1755
rect 3490 1715 3570 1755
rect 3370 1630 3570 1715
rect 3720 1755 3920 1830
rect 3720 1715 3800 1755
rect 3840 1715 3920 1755
rect 3720 1630 3920 1715
rect 4070 1755 4270 1830
rect 4070 1715 4150 1755
rect 4190 1715 4270 1755
rect 4070 1630 4270 1715
rect 4420 1755 4620 1830
rect 4420 1715 4500 1755
rect 4540 1715 4620 1755
rect 4420 1630 4620 1715
rect 4770 1755 4970 1830
rect 4770 1715 4850 1755
rect 4890 1715 4970 1755
rect 4770 1630 4970 1715
rect -3280 1405 -3080 1480
rect -3280 1365 -3200 1405
rect -3160 1365 -3080 1405
rect -3280 1280 -3080 1365
rect -2930 1405 -2730 1480
rect -2930 1365 -2850 1405
rect -2810 1365 -2730 1405
rect -2930 1280 -2730 1365
rect -2580 1405 -2380 1480
rect -2580 1365 -2500 1405
rect -2460 1365 -2380 1405
rect -2580 1280 -2380 1365
rect -2230 1405 -2030 1480
rect -2230 1365 -2150 1405
rect -2110 1365 -2030 1405
rect -2230 1280 -2030 1365
rect -1880 1405 -1680 1480
rect -1880 1365 -1800 1405
rect -1760 1365 -1680 1405
rect -1880 1280 -1680 1365
rect 3370 1405 3570 1480
rect 3370 1365 3450 1405
rect 3490 1365 3570 1405
rect 3370 1280 3570 1365
rect 3720 1405 3920 1480
rect 3720 1365 3800 1405
rect 3840 1365 3920 1405
rect 3720 1280 3920 1365
rect 4070 1405 4270 1480
rect 4070 1365 4150 1405
rect 4190 1365 4270 1405
rect 4070 1280 4270 1365
rect 4420 1405 4620 1480
rect 4420 1365 4500 1405
rect 4540 1365 4620 1405
rect 4420 1280 4620 1365
rect 4770 1405 4970 1480
rect 4770 1365 4850 1405
rect 4890 1365 4970 1405
rect 4770 1280 4970 1365
rect -3280 1055 -3080 1130
rect -3280 1015 -3200 1055
rect -3160 1015 -3080 1055
rect -3280 930 -3080 1015
rect -2930 1055 -2730 1130
rect -2930 1015 -2850 1055
rect -2810 1015 -2730 1055
rect -2930 930 -2730 1015
rect -2580 1055 -2380 1130
rect -2580 1015 -2500 1055
rect -2460 1015 -2380 1055
rect -2580 930 -2380 1015
rect -2230 1055 -2030 1130
rect -2230 1015 -2150 1055
rect -2110 1015 -2030 1055
rect -2230 930 -2030 1015
rect -1880 1055 -1680 1130
rect -1880 1015 -1800 1055
rect -1760 1015 -1680 1055
rect -1880 930 -1680 1015
rect 3370 1055 3570 1130
rect 3370 1015 3450 1055
rect 3490 1015 3570 1055
rect 3370 930 3570 1015
rect 3720 1055 3920 1130
rect 3720 1015 3800 1055
rect 3840 1015 3920 1055
rect 3720 930 3920 1015
rect 4070 1055 4270 1130
rect 4070 1015 4150 1055
rect 4190 1015 4270 1055
rect 4070 930 4270 1015
rect 4420 1055 4620 1130
rect 4420 1015 4500 1055
rect 4540 1015 4620 1055
rect 4420 930 4620 1015
rect 4770 1055 4970 1130
rect 4770 1015 4850 1055
rect 4890 1015 4970 1055
rect 4770 930 4970 1015
rect -3280 705 -3080 780
rect -3280 665 -3200 705
rect -3160 665 -3080 705
rect -3280 580 -3080 665
rect -2930 705 -2730 780
rect -2930 665 -2850 705
rect -2810 665 -2730 705
rect -2930 580 -2730 665
rect -2580 705 -2380 780
rect -2580 665 -2500 705
rect -2460 665 -2380 705
rect -2580 580 -2380 665
rect -2230 705 -2030 780
rect -2230 665 -2150 705
rect -2110 665 -2030 705
rect -2230 580 -2030 665
rect -1880 705 -1680 780
rect -1880 665 -1800 705
rect -1760 665 -1680 705
rect -1880 580 -1680 665
rect 3370 705 3570 780
rect 3370 665 3450 705
rect 3490 665 3570 705
rect 3370 580 3570 665
rect 3720 705 3920 780
rect 3720 665 3800 705
rect 3840 665 3920 705
rect 3720 580 3920 665
rect 4070 705 4270 780
rect 4070 665 4150 705
rect 4190 665 4270 705
rect 4070 580 4270 665
rect 4420 705 4620 780
rect 4420 665 4500 705
rect 4540 665 4620 705
rect 4420 580 4620 665
rect 4770 705 4970 780
rect 4770 665 4850 705
rect 4890 665 4970 705
rect 4770 580 4970 665
rect -3280 355 -3080 430
rect -3280 315 -3200 355
rect -3160 315 -3080 355
rect -3280 230 -3080 315
rect -2930 355 -2730 430
rect -2930 315 -2850 355
rect -2810 315 -2730 355
rect -2930 230 -2730 315
rect -2580 355 -2380 430
rect -2580 315 -2500 355
rect -2460 315 -2380 355
rect -2580 230 -2380 315
rect -2230 355 -2030 430
rect -2230 315 -2150 355
rect -2110 315 -2030 355
rect -2230 230 -2030 315
rect -1880 355 -1680 430
rect -1880 315 -1800 355
rect -1760 315 -1680 355
rect -1880 230 -1680 315
rect 3370 355 3570 430
rect 3370 315 3450 355
rect 3490 315 3570 355
rect 3370 230 3570 315
rect 3720 355 3920 430
rect 3720 315 3800 355
rect 3840 315 3920 355
rect 3720 230 3920 315
rect 4070 355 4270 430
rect 4070 315 4150 355
rect 4190 315 4270 355
rect 4070 230 4270 315
rect 4420 355 4620 430
rect 4420 315 4500 355
rect 4540 315 4620 355
rect 4420 230 4620 315
rect 4770 355 4970 430
rect 4770 315 4850 355
rect 4890 315 4970 355
rect 4770 230 4970 315
rect -3280 5 -3080 80
rect -3280 -35 -3200 5
rect -3160 -35 -3080 5
rect -3280 -120 -3080 -35
rect -2930 5 -2730 80
rect -2930 -35 -2850 5
rect -2810 -35 -2730 5
rect -2930 -120 -2730 -35
rect -2580 5 -2380 80
rect -2580 -35 -2500 5
rect -2460 -35 -2380 5
rect -2580 -120 -2380 -35
rect -2230 5 -2030 80
rect -2230 -35 -2150 5
rect -2110 -35 -2030 5
rect -2230 -120 -2030 -35
rect -1880 5 -1680 80
rect -1880 -35 -1800 5
rect -1760 -35 -1680 5
rect -1880 -120 -1680 -35
rect 3370 5 3570 80
rect 3370 -35 3450 5
rect 3490 -35 3570 5
rect 3370 -120 3570 -35
rect 3720 5 3920 80
rect 3720 -35 3800 5
rect 3840 -35 3920 5
rect 3720 -120 3920 -35
rect 4070 5 4270 80
rect 4070 -35 4150 5
rect 4190 -35 4270 5
rect 4070 -120 4270 -35
rect 4420 5 4620 80
rect 4420 -35 4500 5
rect 4540 -35 4620 5
rect 4420 -120 4620 -35
rect 4770 5 4970 80
rect 4770 -35 4850 5
rect 4890 -35 4970 5
rect 4770 -120 4970 -35
rect -3280 -345 -3080 -270
rect -3280 -385 -3200 -345
rect -3160 -385 -3080 -345
rect -3280 -470 -3080 -385
rect -2930 -345 -2730 -270
rect -2930 -385 -2850 -345
rect -2810 -385 -2730 -345
rect -2930 -470 -2730 -385
rect -2580 -345 -2380 -270
rect -2580 -385 -2500 -345
rect -2460 -385 -2380 -345
rect -2580 -470 -2380 -385
rect -2230 -345 -2030 -270
rect -2230 -385 -2150 -345
rect -2110 -385 -2030 -345
rect -2230 -470 -2030 -385
rect -1880 -345 -1680 -270
rect -1880 -385 -1800 -345
rect -1760 -385 -1680 -345
rect -1880 -470 -1680 -385
rect 3370 -345 3570 -270
rect 3370 -385 3450 -345
rect 3490 -385 3570 -345
rect 3370 -470 3570 -385
rect 3720 -345 3920 -270
rect 3720 -385 3800 -345
rect 3840 -385 3920 -345
rect 3720 -470 3920 -385
rect 4070 -345 4270 -270
rect 4070 -385 4150 -345
rect 4190 -385 4270 -345
rect 4070 -470 4270 -385
rect 4420 -345 4620 -270
rect 4420 -385 4500 -345
rect 4540 -385 4620 -345
rect 4420 -470 4620 -385
rect 4770 -345 4970 -270
rect 4770 -385 4850 -345
rect 4890 -385 4970 -345
rect 4770 -470 4970 -385
rect -3280 -695 -3080 -620
rect -3280 -735 -3200 -695
rect -3160 -735 -3080 -695
rect -3280 -820 -3080 -735
rect -2930 -695 -2730 -620
rect -2930 -735 -2850 -695
rect -2810 -735 -2730 -695
rect -2930 -820 -2730 -735
rect -2580 -695 -2380 -620
rect -2580 -735 -2500 -695
rect -2460 -735 -2380 -695
rect -2580 -820 -2380 -735
rect -2230 -695 -2030 -620
rect -2230 -735 -2150 -695
rect -2110 -735 -2030 -695
rect -2230 -820 -2030 -735
rect -1880 -695 -1680 -620
rect -1880 -735 -1800 -695
rect -1760 -735 -1680 -695
rect -1880 -820 -1680 -735
rect 3370 -695 3570 -620
rect 3370 -735 3450 -695
rect 3490 -735 3570 -695
rect 3370 -820 3570 -735
rect 3720 -695 3920 -620
rect 3720 -735 3800 -695
rect 3840 -735 3920 -695
rect 3720 -820 3920 -735
rect 4070 -695 4270 -620
rect 4070 -735 4150 -695
rect 4190 -735 4270 -695
rect 4070 -820 4270 -735
rect 4420 -695 4620 -620
rect 4420 -735 4500 -695
rect 4540 -735 4620 -695
rect 4420 -820 4620 -735
rect 4770 -695 4970 -620
rect 4770 -735 4850 -695
rect 4890 -735 4970 -695
rect 4770 -820 4970 -735
rect -3280 -1045 -3080 -970
rect -3280 -1085 -3200 -1045
rect -3160 -1085 -3080 -1045
rect -3280 -1170 -3080 -1085
rect -2930 -1045 -2730 -970
rect -2930 -1085 -2850 -1045
rect -2810 -1085 -2730 -1045
rect -2930 -1170 -2730 -1085
rect -2580 -1045 -2380 -970
rect -2580 -1085 -2500 -1045
rect -2460 -1085 -2380 -1045
rect -2580 -1170 -2380 -1085
rect -2230 -1045 -2030 -970
rect -2230 -1085 -2150 -1045
rect -2110 -1085 -2030 -1045
rect -2230 -1170 -2030 -1085
rect -1880 -1045 -1680 -970
rect -1880 -1085 -1800 -1045
rect -1760 -1085 -1680 -1045
rect -1880 -1170 -1680 -1085
rect 3370 -1045 3570 -970
rect 3370 -1085 3450 -1045
rect 3490 -1085 3570 -1045
rect 3370 -1170 3570 -1085
rect 3720 -1045 3920 -970
rect 3720 -1085 3800 -1045
rect 3840 -1085 3920 -1045
rect 3720 -1170 3920 -1085
rect 4070 -1045 4270 -970
rect 4070 -1085 4150 -1045
rect 4190 -1085 4270 -1045
rect 4070 -1170 4270 -1085
rect 4420 -1045 4620 -970
rect 4420 -1085 4500 -1045
rect 4540 -1085 4620 -1045
rect 4420 -1170 4620 -1085
rect 4770 -1045 4970 -970
rect 4770 -1085 4850 -1045
rect 4890 -1085 4970 -1045
rect 4770 -1170 4970 -1085
rect -3280 -1395 -3080 -1320
rect -3280 -1435 -3200 -1395
rect -3160 -1435 -3080 -1395
rect -3280 -1520 -3080 -1435
rect -2930 -1395 -2730 -1320
rect -2930 -1435 -2850 -1395
rect -2810 -1435 -2730 -1395
rect -2930 -1520 -2730 -1435
rect -2580 -1395 -2380 -1320
rect -2580 -1435 -2500 -1395
rect -2460 -1435 -2380 -1395
rect -2580 -1520 -2380 -1435
rect -2230 -1395 -2030 -1320
rect -2230 -1435 -2150 -1395
rect -2110 -1435 -2030 -1395
rect -2230 -1520 -2030 -1435
rect -1880 -1395 -1680 -1320
rect -1880 -1435 -1800 -1395
rect -1760 -1435 -1680 -1395
rect -1880 -1520 -1680 -1435
rect -1530 -1395 -1330 -1320
rect -1530 -1435 -1450 -1395
rect -1410 -1435 -1330 -1395
rect -1530 -1520 -1330 -1435
rect -1180 -1395 -980 -1320
rect -1180 -1435 -1100 -1395
rect -1060 -1435 -980 -1395
rect -1180 -1520 -980 -1435
rect -830 -1395 -630 -1320
rect -830 -1435 -750 -1395
rect -710 -1435 -630 -1395
rect -830 -1520 -630 -1435
rect -480 -1395 -280 -1320
rect -480 -1435 -400 -1395
rect -360 -1435 -280 -1395
rect -480 -1520 -280 -1435
rect -130 -1395 70 -1320
rect -130 -1435 -50 -1395
rect -10 -1435 70 -1395
rect -130 -1520 70 -1435
rect 220 -1395 420 -1320
rect 220 -1435 300 -1395
rect 340 -1435 420 -1395
rect 220 -1520 420 -1435
rect 570 -1395 770 -1320
rect 570 -1435 650 -1395
rect 690 -1435 770 -1395
rect 570 -1520 770 -1435
rect 920 -1395 1120 -1320
rect 920 -1435 1000 -1395
rect 1040 -1435 1120 -1395
rect 920 -1520 1120 -1435
rect 1270 -1395 1470 -1320
rect 1270 -1435 1350 -1395
rect 1390 -1435 1470 -1395
rect 1270 -1520 1470 -1435
rect 1620 -1395 1820 -1320
rect 1620 -1435 1700 -1395
rect 1740 -1435 1820 -1395
rect 1620 -1520 1820 -1435
rect 1970 -1395 2170 -1320
rect 1970 -1435 2050 -1395
rect 2090 -1435 2170 -1395
rect 1970 -1520 2170 -1435
rect 2320 -1395 2520 -1320
rect 2320 -1435 2400 -1395
rect 2440 -1435 2520 -1395
rect 2320 -1520 2520 -1435
rect 2670 -1395 2870 -1320
rect 2670 -1435 2750 -1395
rect 2790 -1435 2870 -1395
rect 2670 -1520 2870 -1435
rect 3020 -1395 3220 -1320
rect 3020 -1435 3100 -1395
rect 3140 -1435 3220 -1395
rect 3020 -1520 3220 -1435
rect 3370 -1395 3570 -1320
rect 3370 -1435 3450 -1395
rect 3490 -1435 3570 -1395
rect 3370 -1520 3570 -1435
rect 3720 -1395 3920 -1320
rect 3720 -1435 3800 -1395
rect 3840 -1435 3920 -1395
rect 3720 -1520 3920 -1435
rect 4070 -1395 4270 -1320
rect 4070 -1435 4150 -1395
rect 4190 -1435 4270 -1395
rect 4070 -1520 4270 -1435
rect 4420 -1395 4620 -1320
rect 4420 -1435 4500 -1395
rect 4540 -1435 4620 -1395
rect 4420 -1520 4620 -1435
rect 4770 -1395 4970 -1320
rect 4770 -1435 4850 -1395
rect 4890 -1435 4970 -1395
rect 4770 -1520 4970 -1435
rect -3280 -1745 -3080 -1670
rect -3280 -1785 -3200 -1745
rect -3160 -1785 -3080 -1745
rect -3280 -1870 -3080 -1785
rect -2930 -1745 -2730 -1670
rect -2930 -1785 -2850 -1745
rect -2810 -1785 -2730 -1745
rect -2930 -1870 -2730 -1785
rect -2580 -1745 -2380 -1670
rect -2580 -1785 -2500 -1745
rect -2460 -1785 -2380 -1745
rect -2580 -1870 -2380 -1785
rect -2230 -1745 -2030 -1670
rect -2230 -1785 -2150 -1745
rect -2110 -1785 -2030 -1745
rect -2230 -1870 -2030 -1785
rect -1880 -1745 -1680 -1670
rect -1880 -1785 -1800 -1745
rect -1760 -1785 -1680 -1745
rect -1880 -1870 -1680 -1785
rect -1530 -1745 -1330 -1670
rect -1530 -1785 -1450 -1745
rect -1410 -1785 -1330 -1745
rect -1530 -1870 -1330 -1785
rect -1180 -1745 -980 -1670
rect -1180 -1785 -1100 -1745
rect -1060 -1785 -980 -1745
rect -1180 -1870 -980 -1785
rect -830 -1745 -630 -1670
rect -830 -1785 -750 -1745
rect -710 -1785 -630 -1745
rect -830 -1870 -630 -1785
rect -480 -1745 -280 -1670
rect -480 -1785 -400 -1745
rect -360 -1785 -280 -1745
rect -480 -1870 -280 -1785
rect -130 -1745 70 -1670
rect -130 -1785 -50 -1745
rect -10 -1785 70 -1745
rect -130 -1870 70 -1785
rect 220 -1745 420 -1670
rect 220 -1785 300 -1745
rect 340 -1785 420 -1745
rect 220 -1870 420 -1785
rect 570 -1745 770 -1670
rect 570 -1785 650 -1745
rect 690 -1785 770 -1745
rect 570 -1870 770 -1785
rect 920 -1745 1120 -1670
rect 920 -1785 1000 -1745
rect 1040 -1785 1120 -1745
rect 920 -1870 1120 -1785
rect 1270 -1745 1470 -1670
rect 1270 -1785 1350 -1745
rect 1390 -1785 1470 -1745
rect 1270 -1870 1470 -1785
rect 1620 -1745 1820 -1670
rect 1620 -1785 1700 -1745
rect 1740 -1785 1820 -1745
rect 1620 -1870 1820 -1785
rect 1970 -1745 2170 -1670
rect 1970 -1785 2050 -1745
rect 2090 -1785 2170 -1745
rect 1970 -1870 2170 -1785
rect 2320 -1745 2520 -1670
rect 2320 -1785 2400 -1745
rect 2440 -1785 2520 -1745
rect 2320 -1870 2520 -1785
rect 2670 -1745 2870 -1670
rect 2670 -1785 2750 -1745
rect 2790 -1785 2870 -1745
rect 2670 -1870 2870 -1785
rect 3020 -1745 3220 -1670
rect 3020 -1785 3100 -1745
rect 3140 -1785 3220 -1745
rect 3020 -1870 3220 -1785
rect 3370 -1745 3570 -1670
rect 3370 -1785 3450 -1745
rect 3490 -1785 3570 -1745
rect 3370 -1870 3570 -1785
rect 3720 -1745 3920 -1670
rect 3720 -1785 3800 -1745
rect 3840 -1785 3920 -1745
rect 3720 -1870 3920 -1785
rect 4070 -1745 4270 -1670
rect 4070 -1785 4150 -1745
rect 4190 -1785 4270 -1745
rect 4070 -1870 4270 -1785
rect 4420 -1745 4620 -1670
rect 4420 -1785 4500 -1745
rect 4540 -1785 4620 -1745
rect 4420 -1870 4620 -1785
rect 4770 -1745 4970 -1670
rect 4770 -1785 4850 -1745
rect 4890 -1785 4970 -1745
rect 4770 -1870 4970 -1785
rect -3280 -2095 -3080 -2020
rect -3280 -2135 -3200 -2095
rect -3160 -2135 -3080 -2095
rect -3280 -2220 -3080 -2135
rect -2930 -2095 -2730 -2020
rect -2930 -2135 -2850 -2095
rect -2810 -2135 -2730 -2095
rect -2930 -2220 -2730 -2135
rect -2580 -2095 -2380 -2020
rect -2580 -2135 -2500 -2095
rect -2460 -2135 -2380 -2095
rect -2580 -2220 -2380 -2135
rect -2230 -2095 -2030 -2020
rect -2230 -2135 -2150 -2095
rect -2110 -2135 -2030 -2095
rect -2230 -2220 -2030 -2135
rect -1880 -2095 -1680 -2020
rect -1880 -2135 -1800 -2095
rect -1760 -2135 -1680 -2095
rect -1880 -2220 -1680 -2135
rect -1530 -2095 -1330 -2020
rect -1530 -2135 -1450 -2095
rect -1410 -2135 -1330 -2095
rect -1530 -2220 -1330 -2135
rect -1180 -2095 -980 -2020
rect -1180 -2135 -1100 -2095
rect -1060 -2135 -980 -2095
rect -1180 -2220 -980 -2135
rect -830 -2095 -630 -2020
rect -830 -2135 -750 -2095
rect -710 -2135 -630 -2095
rect -830 -2220 -630 -2135
rect -480 -2095 -280 -2020
rect -480 -2135 -400 -2095
rect -360 -2135 -280 -2095
rect -480 -2220 -280 -2135
rect -130 -2095 70 -2020
rect -130 -2135 -50 -2095
rect -10 -2135 70 -2095
rect -130 -2220 70 -2135
rect 220 -2095 420 -2020
rect 220 -2135 300 -2095
rect 340 -2135 420 -2095
rect 220 -2220 420 -2135
rect 570 -2095 770 -2020
rect 570 -2135 650 -2095
rect 690 -2135 770 -2095
rect 570 -2220 770 -2135
rect 920 -2095 1120 -2020
rect 920 -2135 1000 -2095
rect 1040 -2135 1120 -2095
rect 920 -2220 1120 -2135
rect 1270 -2095 1470 -2020
rect 1270 -2135 1350 -2095
rect 1390 -2135 1470 -2095
rect 1270 -2220 1470 -2135
rect 1620 -2095 1820 -2020
rect 1620 -2135 1700 -2095
rect 1740 -2135 1820 -2095
rect 1620 -2220 1820 -2135
rect 1970 -2095 2170 -2020
rect 1970 -2135 2050 -2095
rect 2090 -2135 2170 -2095
rect 1970 -2220 2170 -2135
rect 2320 -2095 2520 -2020
rect 2320 -2135 2400 -2095
rect 2440 -2135 2520 -2095
rect 2320 -2220 2520 -2135
rect 2670 -2095 2870 -2020
rect 2670 -2135 2750 -2095
rect 2790 -2135 2870 -2095
rect 2670 -2220 2870 -2135
rect 3020 -2095 3220 -2020
rect 3020 -2135 3100 -2095
rect 3140 -2135 3220 -2095
rect 3020 -2220 3220 -2135
rect 3370 -2095 3570 -2020
rect 3370 -2135 3450 -2095
rect 3490 -2135 3570 -2095
rect 3370 -2220 3570 -2135
rect 3720 -2095 3920 -2020
rect 3720 -2135 3800 -2095
rect 3840 -2135 3920 -2095
rect 3720 -2220 3920 -2135
rect 4070 -2095 4270 -2020
rect 4070 -2135 4150 -2095
rect 4190 -2135 4270 -2095
rect 4070 -2220 4270 -2135
rect 4420 -2095 4620 -2020
rect 4420 -2135 4500 -2095
rect 4540 -2135 4620 -2095
rect 4420 -2220 4620 -2135
rect 4770 -2095 4970 -2020
rect 4770 -2135 4850 -2095
rect 4890 -2135 4970 -2095
rect 4770 -2220 4970 -2135
<< mimcapcontact >>
rect -3200 3815 -3160 3855
rect -2850 3815 -2810 3855
rect -2500 3815 -2460 3855
rect -2150 3815 -2110 3855
rect -1800 3815 -1760 3855
rect -1450 3815 -1410 3855
rect -1100 3815 -1060 3855
rect -750 3815 -710 3855
rect -400 3815 -360 3855
rect -50 3815 -10 3855
rect 300 3815 340 3855
rect 650 3815 690 3855
rect 1000 3815 1040 3855
rect 1350 3815 1390 3855
rect 1700 3815 1740 3855
rect 2050 3815 2090 3855
rect 2400 3815 2440 3855
rect 2750 3815 2790 3855
rect 3100 3815 3140 3855
rect 3450 3815 3490 3855
rect 3800 3815 3840 3855
rect 4150 3815 4190 3855
rect 4500 3815 4540 3855
rect 4850 3815 4890 3855
rect -3200 3465 -3160 3505
rect -2850 3465 -2810 3505
rect -2500 3465 -2460 3505
rect -2150 3465 -2110 3505
rect -1800 3465 -1760 3505
rect -1450 3465 -1410 3505
rect -1100 3465 -1060 3505
rect -750 3465 -710 3505
rect -400 3465 -360 3505
rect -50 3465 -10 3505
rect 300 3465 340 3505
rect 650 3465 690 3505
rect 1000 3465 1040 3505
rect 1350 3465 1390 3505
rect 1700 3465 1740 3505
rect 2050 3465 2090 3505
rect 2400 3465 2440 3505
rect 2750 3465 2790 3505
rect 3100 3465 3140 3505
rect 3450 3465 3490 3505
rect 3800 3465 3840 3505
rect 4150 3465 4190 3505
rect 4500 3465 4540 3505
rect 4850 3465 4890 3505
rect -3200 3115 -3160 3155
rect -2850 3115 -2810 3155
rect -2500 3115 -2460 3155
rect -2150 3115 -2110 3155
rect -1800 3115 -1760 3155
rect -1450 3115 -1410 3155
rect -1100 3115 -1060 3155
rect -750 3115 -710 3155
rect -400 3115 -360 3155
rect -50 3105 -10 3145
rect 300 3105 340 3145
rect 650 3105 690 3145
rect 1000 3105 1040 3145
rect 1350 3105 1390 3145
rect 1700 3105 1740 3145
rect 2050 3115 2090 3155
rect 2400 3115 2440 3155
rect 2750 3115 2790 3155
rect 3100 3115 3140 3155
rect 3450 3115 3490 3155
rect 3800 3115 3840 3155
rect 4150 3115 4190 3155
rect 4500 3115 4540 3155
rect 4850 3115 4890 3155
rect -3200 2765 -3160 2805
rect -2850 2765 -2810 2805
rect -2500 2765 -2460 2805
rect -2150 2765 -2110 2805
rect -1800 2765 -1760 2805
rect -1450 2765 -1410 2805
rect -1100 2765 -1060 2805
rect -750 2765 -710 2805
rect 2400 2765 2440 2805
rect 2750 2765 2790 2805
rect 3100 2765 3140 2805
rect 3450 2765 3490 2805
rect 3800 2765 3840 2805
rect 4150 2765 4190 2805
rect 4500 2765 4540 2805
rect 4850 2765 4890 2805
rect -3200 2415 -3160 2455
rect -2850 2415 -2810 2455
rect -2500 2415 -2460 2455
rect -2150 2415 -2110 2455
rect -1800 2415 -1760 2455
rect -1450 2415 -1410 2455
rect -1100 2415 -1060 2455
rect -750 2415 -710 2455
rect 2400 2415 2440 2455
rect 2750 2415 2790 2455
rect 3100 2415 3140 2455
rect 3450 2415 3490 2455
rect 3800 2415 3840 2455
rect 4150 2415 4190 2455
rect 4500 2415 4540 2455
rect 4850 2415 4890 2455
rect -3200 2065 -3160 2105
rect -2850 2065 -2810 2105
rect -2500 2065 -2460 2105
rect -2150 2065 -2110 2105
rect -1800 2065 -1760 2105
rect 3450 2065 3490 2105
rect 3800 2065 3840 2105
rect 4150 2065 4190 2105
rect 4500 2065 4540 2105
rect 4850 2065 4890 2105
rect -3200 1715 -3160 1755
rect -2850 1715 -2810 1755
rect -2500 1715 -2460 1755
rect -2150 1715 -2110 1755
rect -1800 1715 -1760 1755
rect 3450 1715 3490 1755
rect 3800 1715 3840 1755
rect 4150 1715 4190 1755
rect 4500 1715 4540 1755
rect 4850 1715 4890 1755
rect -3200 1365 -3160 1405
rect -2850 1365 -2810 1405
rect -2500 1365 -2460 1405
rect -2150 1365 -2110 1405
rect -1800 1365 -1760 1405
rect 3450 1365 3490 1405
rect 3800 1365 3840 1405
rect 4150 1365 4190 1405
rect 4500 1365 4540 1405
rect 4850 1365 4890 1405
rect -3200 1015 -3160 1055
rect -2850 1015 -2810 1055
rect -2500 1015 -2460 1055
rect -2150 1015 -2110 1055
rect -1800 1015 -1760 1055
rect 3450 1015 3490 1055
rect 3800 1015 3840 1055
rect 4150 1015 4190 1055
rect 4500 1015 4540 1055
rect 4850 1015 4890 1055
rect -3200 665 -3160 705
rect -2850 665 -2810 705
rect -2500 665 -2460 705
rect -2150 665 -2110 705
rect -1800 665 -1760 705
rect 3450 665 3490 705
rect 3800 665 3840 705
rect 4150 665 4190 705
rect 4500 665 4540 705
rect 4850 665 4890 705
rect -3200 315 -3160 355
rect -2850 315 -2810 355
rect -2500 315 -2460 355
rect -2150 315 -2110 355
rect -1800 315 -1760 355
rect 3450 315 3490 355
rect 3800 315 3840 355
rect 4150 315 4190 355
rect 4500 315 4540 355
rect 4850 315 4890 355
rect -3200 -35 -3160 5
rect -2850 -35 -2810 5
rect -2500 -35 -2460 5
rect -2150 -35 -2110 5
rect -1800 -35 -1760 5
rect 3450 -35 3490 5
rect 3800 -35 3840 5
rect 4150 -35 4190 5
rect 4500 -35 4540 5
rect 4850 -35 4890 5
rect -3200 -385 -3160 -345
rect -2850 -385 -2810 -345
rect -2500 -385 -2460 -345
rect -2150 -385 -2110 -345
rect -1800 -385 -1760 -345
rect 3450 -385 3490 -345
rect 3800 -385 3840 -345
rect 4150 -385 4190 -345
rect 4500 -385 4540 -345
rect 4850 -385 4890 -345
rect -3200 -735 -3160 -695
rect -2850 -735 -2810 -695
rect -2500 -735 -2460 -695
rect -2150 -735 -2110 -695
rect -1800 -735 -1760 -695
rect 3450 -735 3490 -695
rect 3800 -735 3840 -695
rect 4150 -735 4190 -695
rect 4500 -735 4540 -695
rect 4850 -735 4890 -695
rect -3200 -1085 -3160 -1045
rect -2850 -1085 -2810 -1045
rect -2500 -1085 -2460 -1045
rect -2150 -1085 -2110 -1045
rect -1800 -1085 -1760 -1045
rect 3450 -1085 3490 -1045
rect 3800 -1085 3840 -1045
rect 4150 -1085 4190 -1045
rect 4500 -1085 4540 -1045
rect 4850 -1085 4890 -1045
rect -3200 -1435 -3160 -1395
rect -2850 -1435 -2810 -1395
rect -2500 -1435 -2460 -1395
rect -2150 -1435 -2110 -1395
rect -1800 -1435 -1760 -1395
rect -1450 -1435 -1410 -1395
rect -1100 -1435 -1060 -1395
rect -750 -1435 -710 -1395
rect -400 -1435 -360 -1395
rect -50 -1435 -10 -1395
rect 300 -1435 340 -1395
rect 650 -1435 690 -1395
rect 1000 -1435 1040 -1395
rect 1350 -1435 1390 -1395
rect 1700 -1435 1740 -1395
rect 2050 -1435 2090 -1395
rect 2400 -1435 2440 -1395
rect 2750 -1435 2790 -1395
rect 3100 -1435 3140 -1395
rect 3450 -1435 3490 -1395
rect 3800 -1435 3840 -1395
rect 4150 -1435 4190 -1395
rect 4500 -1435 4540 -1395
rect 4850 -1435 4890 -1395
rect -3200 -1785 -3160 -1745
rect -2850 -1785 -2810 -1745
rect -2500 -1785 -2460 -1745
rect -2150 -1785 -2110 -1745
rect -1800 -1785 -1760 -1745
rect -1450 -1785 -1410 -1745
rect -1100 -1785 -1060 -1745
rect -750 -1785 -710 -1745
rect -400 -1785 -360 -1745
rect -50 -1785 -10 -1745
rect 300 -1785 340 -1745
rect 650 -1785 690 -1745
rect 1000 -1785 1040 -1745
rect 1350 -1785 1390 -1745
rect 1700 -1785 1740 -1745
rect 2050 -1785 2090 -1745
rect 2400 -1785 2440 -1745
rect 2750 -1785 2790 -1745
rect 3100 -1785 3140 -1745
rect 3450 -1785 3490 -1745
rect 3800 -1785 3840 -1745
rect 4150 -1785 4190 -1745
rect 4500 -1785 4540 -1745
rect 4850 -1785 4890 -1745
rect -3200 -2135 -3160 -2095
rect -2850 -2135 -2810 -2095
rect -2500 -2135 -2460 -2095
rect -2150 -2135 -2110 -2095
rect -1800 -2135 -1760 -2095
rect -1450 -2135 -1410 -2095
rect -1100 -2135 -1060 -2095
rect -750 -2135 -710 -2095
rect -400 -2135 -360 -2095
rect -50 -2135 -10 -2095
rect 300 -2135 340 -2095
rect 650 -2135 690 -2095
rect 1000 -2135 1040 -2095
rect 1350 -2135 1390 -2095
rect 1700 -2135 1740 -2095
rect 2050 -2135 2090 -2095
rect 2400 -2135 2440 -2095
rect 2750 -2135 2790 -2095
rect 3100 -2135 3140 -2095
rect 3450 -2135 3490 -2095
rect 3800 -2135 3840 -2095
rect 4150 -2135 4190 -2095
rect 4500 -2135 4540 -2095
rect 4850 -2135 4890 -2095
<< metal4 >>
rect -3850 4280 5140 4285
rect -3850 4240 825 4280
rect 865 4240 5140 4280
rect -3850 4235 5140 4240
rect -3205 3855 -2455 3860
rect -3205 3815 -3200 3855
rect -3160 3815 -2850 3855
rect -2810 3815 -2500 3855
rect -2460 3815 -2455 3855
rect -3205 3810 -2455 3815
rect -2505 3510 -2455 3810
rect -2155 3855 -2105 3860
rect -2155 3815 -2150 3855
rect -2110 3815 -2105 3855
rect -2155 3510 -2105 3815
rect -1805 3855 -1755 3860
rect -1805 3815 -1800 3855
rect -1760 3815 -1755 3855
rect -1805 3510 -1755 3815
rect -1455 3855 -1405 3860
rect -1455 3815 -1450 3855
rect -1410 3815 -1405 3855
rect -1455 3510 -1405 3815
rect -1105 3855 -1055 3860
rect -1105 3815 -1100 3855
rect -1060 3815 -1055 3855
rect -1105 3510 -1055 3815
rect -755 3855 -705 3860
rect -755 3815 -750 3855
rect -710 3815 -705 3855
rect -755 3510 -705 3815
rect -405 3855 -355 3860
rect -405 3815 -400 3855
rect -360 3815 -355 3855
rect -405 3510 -355 3815
rect -55 3855 -5 3860
rect -55 3815 -50 3855
rect -10 3815 -5 3855
rect -55 3510 -5 3815
rect 295 3855 345 3860
rect 295 3815 300 3855
rect 340 3815 345 3855
rect 295 3510 345 3815
rect 645 3855 695 3860
rect 645 3815 650 3855
rect 690 3815 695 3855
rect 645 3510 695 3815
rect -3205 3505 695 3510
rect -3205 3465 -3200 3505
rect -3160 3465 -2850 3505
rect -2810 3465 -2500 3505
rect -2460 3465 -2150 3505
rect -2110 3465 -1800 3505
rect -1760 3465 -1450 3505
rect -1410 3465 -1100 3505
rect -1060 3465 -750 3505
rect -710 3465 -400 3505
rect -360 3465 -50 3505
rect -10 3465 300 3505
rect 340 3465 650 3505
rect 690 3465 695 3505
rect -3205 3460 695 3465
rect -2505 3160 -2455 3460
rect -3205 3155 -2105 3160
rect -3205 3115 -3200 3155
rect -3160 3115 -2850 3155
rect -2810 3115 -2500 3155
rect -2460 3115 -2150 3155
rect -2110 3115 -2105 3155
rect -3205 3110 -2105 3115
rect -1805 3155 -1755 3460
rect -1805 3115 -1800 3155
rect -1760 3115 -1755 3155
rect -2505 2810 -2455 3110
rect -3205 2805 -2105 2810
rect -3205 2765 -3200 2805
rect -3160 2765 -2850 2805
rect -2810 2765 -2500 2805
rect -2460 2765 -2150 2805
rect -2110 2765 -2105 2805
rect -3205 2760 -2105 2765
rect -1805 2805 -1755 3115
rect -1805 2765 -1800 2805
rect -1760 2765 -1755 2805
rect -1805 2760 -1755 2765
rect -1455 3155 -1405 3460
rect -1455 3115 -1450 3155
rect -1410 3115 -1405 3155
rect -1455 2805 -1405 3115
rect -1455 2765 -1450 2805
rect -1410 2765 -1405 2805
rect -2505 2460 -2455 2760
rect -3205 2455 -1755 2460
rect -3205 2415 -3200 2455
rect -3160 2415 -2850 2455
rect -2810 2415 -2500 2455
rect -2460 2415 -2150 2455
rect -2110 2415 -1800 2455
rect -1760 2415 -1755 2455
rect -3205 2410 -1755 2415
rect -1455 2455 -1405 2765
rect -1455 2415 -1450 2455
rect -1410 2415 -1405 2455
rect -1455 2410 -1405 2415
rect -1105 3155 -1055 3460
rect -1105 3115 -1100 3155
rect -1060 3115 -1055 3155
rect -1105 2805 -1055 3115
rect -1105 2765 -1100 2805
rect -1060 2765 -1055 2805
rect -1105 2455 -1055 2765
rect -1105 2415 -1100 2455
rect -1060 2415 -1055 2455
rect -1105 2410 -1055 2415
rect -755 3155 -705 3460
rect -755 3115 -750 3155
rect -710 3115 -705 3155
rect -755 2805 -705 3115
rect -405 3155 -355 3460
rect -405 3115 -400 3155
rect -360 3115 -355 3155
rect -405 3110 -355 3115
rect -55 3145 -5 3460
rect -55 3105 -50 3145
rect -10 3105 -5 3145
rect -55 3100 -5 3105
rect 295 3145 345 3460
rect 295 3105 300 3145
rect 340 3105 345 3145
rect 295 3100 345 3105
rect 645 3145 695 3460
rect 645 3105 650 3145
rect 690 3105 695 3145
rect 645 3100 695 3105
rect 995 3855 1045 3860
rect 995 3815 1000 3855
rect 1040 3815 1045 3855
rect 995 3510 1045 3815
rect 1345 3855 1395 3860
rect 1345 3815 1350 3855
rect 1390 3815 1395 3855
rect 1345 3510 1395 3815
rect 1695 3855 1745 3860
rect 1695 3815 1700 3855
rect 1740 3815 1745 3855
rect 1695 3510 1745 3815
rect 2045 3855 2095 3860
rect 2045 3815 2050 3855
rect 2090 3815 2095 3855
rect 2045 3510 2095 3815
rect 2395 3855 2445 3860
rect 2395 3815 2400 3855
rect 2440 3815 2445 3855
rect 2395 3510 2445 3815
rect 2745 3855 2795 3860
rect 2745 3815 2750 3855
rect 2790 3815 2795 3855
rect 2745 3510 2795 3815
rect 3095 3855 3145 3860
rect 3095 3815 3100 3855
rect 3140 3815 3145 3855
rect 3095 3510 3145 3815
rect 3445 3855 3495 3860
rect 3445 3815 3450 3855
rect 3490 3815 3495 3855
rect 3445 3510 3495 3815
rect 3795 3855 3845 3860
rect 3795 3815 3800 3855
rect 3840 3815 3845 3855
rect 3795 3510 3845 3815
rect 4145 3855 4895 3860
rect 4145 3815 4150 3855
rect 4190 3815 4500 3855
rect 4540 3815 4850 3855
rect 4890 3815 4895 3855
rect 4145 3810 4895 3815
rect 4145 3510 4195 3810
rect 995 3505 4895 3510
rect 995 3465 1000 3505
rect 1040 3465 1350 3505
rect 1390 3465 1700 3505
rect 1740 3465 2050 3505
rect 2090 3465 2400 3505
rect 2440 3465 2750 3505
rect 2790 3465 3100 3505
rect 3140 3465 3450 3505
rect 3490 3465 3800 3505
rect 3840 3465 4150 3505
rect 4190 3465 4500 3505
rect 4540 3465 4850 3505
rect 4890 3465 4895 3505
rect 995 3460 4895 3465
rect 995 3145 1045 3460
rect 995 3105 1000 3145
rect 1040 3105 1045 3145
rect 995 3100 1045 3105
rect 1345 3145 1395 3460
rect 1345 3105 1350 3145
rect 1390 3105 1395 3145
rect 1345 3100 1395 3105
rect 1695 3145 1745 3460
rect 1695 3105 1700 3145
rect 1740 3105 1745 3145
rect 2045 3155 2095 3460
rect 2045 3115 2050 3155
rect 2090 3115 2095 3155
rect 2045 3110 2095 3115
rect 2395 3155 2445 3460
rect 2395 3115 2400 3155
rect 2440 3115 2445 3155
rect 1695 3100 1745 3105
rect -755 2765 -750 2805
rect -710 2765 -705 2805
rect -755 2455 -705 2765
rect -755 2415 -750 2455
rect -710 2415 -705 2455
rect -755 2410 -705 2415
rect 2395 2805 2445 3115
rect 2395 2765 2400 2805
rect 2440 2765 2445 2805
rect 2395 2455 2445 2765
rect 2395 2415 2400 2455
rect 2440 2415 2445 2455
rect 2395 2410 2445 2415
rect 2745 3155 2795 3460
rect 2745 3115 2750 3155
rect 2790 3115 2795 3155
rect 2745 2805 2795 3115
rect 2745 2765 2750 2805
rect 2790 2765 2795 2805
rect 2745 2455 2795 2765
rect 2745 2415 2750 2455
rect 2790 2415 2795 2455
rect 2745 2410 2795 2415
rect 3095 3155 3145 3460
rect 3095 3115 3100 3155
rect 3140 3115 3145 3155
rect 3095 2805 3145 3115
rect 3095 2765 3100 2805
rect 3140 2765 3145 2805
rect 3095 2455 3145 2765
rect 3445 3155 3495 3460
rect 4145 3160 4195 3460
rect 3445 3115 3450 3155
rect 3490 3115 3495 3155
rect 3445 2805 3495 3115
rect 3795 3155 4895 3160
rect 3795 3115 3800 3155
rect 3840 3115 4150 3155
rect 4190 3115 4500 3155
rect 4540 3115 4850 3155
rect 4890 3115 4895 3155
rect 3795 3110 4895 3115
rect 4145 2810 4195 3110
rect 3445 2765 3450 2805
rect 3490 2765 3495 2805
rect 3445 2760 3495 2765
rect 3795 2805 4895 2810
rect 3795 2765 3800 2805
rect 3840 2765 4150 2805
rect 4190 2765 4500 2805
rect 4540 2765 4850 2805
rect 4890 2765 4895 2805
rect 3795 2760 4895 2765
rect 4145 2460 4195 2760
rect 3095 2415 3100 2455
rect 3140 2415 3145 2455
rect 3095 2410 3145 2415
rect 3445 2455 4895 2460
rect 3445 2415 3450 2455
rect 3490 2415 3800 2455
rect 3840 2415 4150 2455
rect 4190 2415 4500 2455
rect 4540 2415 4850 2455
rect 4890 2415 4895 2455
rect 3445 2410 4895 2415
rect -2505 2110 -2455 2410
rect 4145 2110 4195 2410
rect -3205 2105 -1755 2110
rect -3205 2065 -3200 2105
rect -3160 2065 -2850 2105
rect -2810 2065 -2500 2105
rect -2460 2065 -2150 2105
rect -2110 2065 -1800 2105
rect -1760 2065 -1755 2105
rect -3205 2060 -1755 2065
rect 3445 2105 4895 2110
rect 3445 2065 3450 2105
rect 3490 2065 3800 2105
rect 3840 2065 4150 2105
rect 4190 2065 4500 2105
rect 4540 2065 4850 2105
rect 4890 2065 4895 2105
rect 3445 2060 4895 2065
rect -2505 1760 -2455 2060
rect 4145 1760 4195 2060
rect -3205 1755 -1755 1760
rect -3205 1715 -3200 1755
rect -3160 1715 -2850 1755
rect -2810 1715 -2500 1755
rect -2460 1715 -2150 1755
rect -2110 1715 -1800 1755
rect -1760 1715 -1755 1755
rect -3205 1710 -1755 1715
rect 3445 1755 4895 1760
rect 3445 1715 3450 1755
rect 3490 1715 3800 1755
rect 3840 1715 4150 1755
rect 4190 1715 4500 1755
rect 4540 1715 4850 1755
rect 4890 1715 4895 1755
rect 3445 1710 4895 1715
rect -2505 1410 -2455 1710
rect 4145 1410 4195 1710
rect -3205 1405 -1755 1410
rect -3205 1365 -3200 1405
rect -3160 1365 -2850 1405
rect -2810 1365 -2500 1405
rect -2460 1365 -2150 1405
rect -2110 1365 -1800 1405
rect -1760 1365 -1755 1405
rect -3205 1360 -1755 1365
rect 3445 1405 4895 1410
rect 3445 1365 3450 1405
rect 3490 1365 3800 1405
rect 3840 1365 4150 1405
rect 4190 1365 4500 1405
rect 4540 1365 4850 1405
rect 4890 1365 4895 1405
rect 3445 1360 4895 1365
rect -2505 1060 -2455 1360
rect 4145 1060 4195 1360
rect -3205 1055 -1755 1060
rect -3205 1015 -3200 1055
rect -3160 1015 -2850 1055
rect -2810 1015 -2500 1055
rect -2460 1015 -2150 1055
rect -2110 1015 -1800 1055
rect -1760 1015 -1755 1055
rect -3205 1010 -1755 1015
rect 3445 1055 4895 1060
rect 3445 1015 3450 1055
rect 3490 1015 3800 1055
rect 3840 1015 4150 1055
rect 4190 1015 4500 1055
rect 4540 1015 4850 1055
rect 4890 1015 4895 1055
rect 3445 1010 4895 1015
rect -2505 710 -2455 1010
rect 4145 710 4195 1010
rect -3205 705 -1755 710
rect -3205 665 -3200 705
rect -3160 665 -2850 705
rect -2810 665 -2500 705
rect -2460 665 -2150 705
rect -2110 665 -1800 705
rect -1760 665 -1755 705
rect -3205 660 -1755 665
rect 3445 705 4895 710
rect 3445 665 3450 705
rect 3490 665 3800 705
rect 3840 665 4150 705
rect 4190 665 4500 705
rect 4540 665 4850 705
rect 4890 665 4895 705
rect 3445 660 4895 665
rect -2505 360 -2455 660
rect 4145 360 4195 660
rect -3205 355 -1495 360
rect -3205 315 -3200 355
rect -3160 315 -2850 355
rect -2810 315 -2500 355
rect -2460 315 -2150 355
rect -2110 315 -1800 355
rect -1760 315 -1540 355
rect -1500 315 -1495 355
rect -3205 310 -1495 315
rect 3185 355 4895 360
rect 3185 315 3190 355
rect 3230 315 3450 355
rect 3490 315 3800 355
rect 3840 315 4150 355
rect 4190 315 4500 355
rect 4540 315 4850 355
rect 4890 315 4895 355
rect 3185 310 4895 315
rect -2505 10 -2455 310
rect 4145 10 4195 310
rect -3205 5 -1755 10
rect -3205 -35 -3200 5
rect -3160 -35 -2850 5
rect -2810 -35 -2500 5
rect -2460 -35 -2150 5
rect -2110 -35 -1800 5
rect -1760 -35 -1755 5
rect -3205 -40 -1755 -35
rect 3445 5 4895 10
rect 3445 -35 3450 5
rect 3490 -35 3800 5
rect 3840 -35 4150 5
rect 4190 -35 4500 5
rect 4540 -35 4850 5
rect 4890 -35 4895 5
rect 3445 -40 4895 -35
rect -2505 -340 -2455 -40
rect 4145 -340 4195 -40
rect -3205 -345 -1755 -340
rect -3205 -385 -3200 -345
rect -3160 -385 -2850 -345
rect -2810 -385 -2500 -345
rect -2460 -385 -2150 -345
rect -2110 -385 -1800 -345
rect -1760 -385 -1755 -345
rect -3205 -390 -1755 -385
rect 3445 -345 4895 -340
rect 3445 -385 3450 -345
rect 3490 -385 3800 -345
rect 3840 -385 4150 -345
rect 4190 -385 4500 -345
rect 4540 -385 4850 -345
rect 4890 -385 4895 -345
rect 3445 -390 4895 -385
rect -2505 -690 -2455 -390
rect 4145 -690 4195 -390
rect -3205 -695 -1755 -690
rect -3205 -735 -3200 -695
rect -3160 -735 -2850 -695
rect -2810 -735 -2500 -695
rect -2460 -735 -2150 -695
rect -2110 -735 -1800 -695
rect -1760 -735 -1755 -695
rect -3205 -740 -1755 -735
rect 3445 -695 4895 -690
rect 3445 -735 3450 -695
rect 3490 -735 3800 -695
rect 3840 -735 4150 -695
rect 4190 -735 4500 -695
rect 4540 -735 4850 -695
rect 4890 -735 4895 -695
rect 3445 -740 4895 -735
rect -2505 -1040 -2455 -740
rect 4145 -1040 4195 -740
rect -3205 -1045 -1755 -1040
rect -3205 -1085 -3200 -1045
rect -3160 -1085 -2850 -1045
rect -2810 -1085 -2500 -1045
rect -2460 -1085 -2150 -1045
rect -2110 -1085 -1800 -1045
rect -1760 -1085 -1755 -1045
rect -3205 -1090 -1755 -1085
rect 3445 -1045 4895 -1040
rect 3445 -1085 3450 -1045
rect 3490 -1085 3800 -1045
rect 3840 -1085 4150 -1045
rect 4190 -1085 4500 -1045
rect 4540 -1085 4850 -1045
rect 4890 -1085 4895 -1045
rect 3445 -1090 4895 -1085
rect -2505 -1390 -2455 -1090
rect 4145 -1390 4195 -1090
rect -3205 -1395 -1755 -1390
rect -3205 -1435 -3200 -1395
rect -3160 -1435 -2850 -1395
rect -2810 -1435 -2500 -1395
rect -2460 -1435 -2150 -1395
rect -2110 -1435 -1800 -1395
rect -1760 -1435 -1755 -1395
rect -3205 -1440 -1755 -1435
rect -1455 -1395 -1405 -1390
rect -1455 -1435 -1450 -1395
rect -1410 -1435 -1405 -1395
rect -2505 -1740 -2455 -1440
rect -1455 -1740 -1405 -1435
rect -1105 -1395 -1055 -1390
rect -1105 -1435 -1100 -1395
rect -1060 -1435 -1055 -1395
rect -1105 -1740 -1055 -1435
rect -755 -1395 -705 -1390
rect -755 -1435 -750 -1395
rect -710 -1435 -705 -1395
rect -755 -1740 -705 -1435
rect -405 -1395 -355 -1390
rect -405 -1435 -400 -1395
rect -360 -1435 -355 -1395
rect -405 -1740 -355 -1435
rect -55 -1395 -5 -1390
rect -55 -1435 -50 -1395
rect -10 -1435 -5 -1395
rect -55 -1740 -5 -1435
rect 295 -1395 345 -1390
rect 295 -1435 300 -1395
rect 340 -1435 345 -1395
rect 295 -1740 345 -1435
rect 645 -1395 695 -1390
rect 645 -1435 650 -1395
rect 690 -1435 695 -1395
rect 645 -1740 695 -1435
rect -3205 -1745 695 -1740
rect -3205 -1785 -3200 -1745
rect -3160 -1785 -2850 -1745
rect -2810 -1785 -2500 -1745
rect -2460 -1785 -2150 -1745
rect -2110 -1785 -1800 -1745
rect -1760 -1785 -1450 -1745
rect -1410 -1785 -1100 -1745
rect -1060 -1785 -750 -1745
rect -710 -1785 -400 -1745
rect -360 -1785 -50 -1745
rect -10 -1785 300 -1745
rect 340 -1785 650 -1745
rect 690 -1785 695 -1745
rect -3205 -1790 695 -1785
rect -2505 -2090 -2455 -1790
rect -3205 -2095 -2455 -2090
rect -3205 -2135 -3200 -2095
rect -3160 -2135 -2850 -2095
rect -2810 -2135 -2500 -2095
rect -2460 -2135 -2455 -2095
rect -3205 -2140 -2455 -2135
rect -2155 -2095 -2105 -1790
rect -2155 -2135 -2150 -2095
rect -2110 -2135 -2105 -2095
rect -2155 -2140 -2105 -2135
rect -1805 -2095 -1755 -1790
rect -1805 -2135 -1800 -2095
rect -1760 -2135 -1755 -2095
rect -1805 -2140 -1755 -2135
rect -1455 -2095 -1405 -1790
rect -1455 -2135 -1450 -2095
rect -1410 -2135 -1405 -2095
rect -1455 -2140 -1405 -2135
rect -1105 -2095 -1055 -1790
rect -1105 -2135 -1100 -2095
rect -1060 -2135 -1055 -2095
rect -1105 -2140 -1055 -2135
rect -755 -2095 -705 -1790
rect -755 -2135 -750 -2095
rect -710 -2135 -705 -2095
rect -755 -2140 -705 -2135
rect -405 -2095 -355 -1790
rect -405 -2135 -400 -2095
rect -360 -2135 -355 -2095
rect -405 -2140 -355 -2135
rect -55 -2095 -5 -1790
rect -55 -2135 -50 -2095
rect -10 -2135 -5 -2095
rect -55 -2140 -5 -2135
rect 295 -2095 345 -1790
rect 295 -2135 300 -2095
rect 340 -2135 345 -2095
rect 295 -2140 345 -2135
rect 645 -2095 695 -1790
rect 645 -2135 650 -2095
rect 690 -2135 695 -2095
rect 645 -2140 695 -2135
rect 995 -1395 1045 -1390
rect 995 -1435 1000 -1395
rect 1040 -1435 1045 -1395
rect 995 -1740 1045 -1435
rect 1345 -1395 1395 -1390
rect 1345 -1435 1350 -1395
rect 1390 -1435 1395 -1395
rect 1345 -1740 1395 -1435
rect 1695 -1395 1745 -1390
rect 1695 -1435 1700 -1395
rect 1740 -1435 1745 -1395
rect 1695 -1740 1745 -1435
rect 2045 -1395 2095 -1390
rect 2045 -1435 2050 -1395
rect 2090 -1435 2095 -1395
rect 2045 -1740 2095 -1435
rect 2395 -1395 2445 -1390
rect 2395 -1435 2400 -1395
rect 2440 -1435 2445 -1395
rect 2395 -1740 2445 -1435
rect 2745 -1395 2795 -1390
rect 2745 -1435 2750 -1395
rect 2790 -1435 2795 -1395
rect 2745 -1740 2795 -1435
rect 3095 -1395 3145 -1390
rect 3095 -1435 3100 -1395
rect 3140 -1435 3145 -1395
rect 3095 -1740 3145 -1435
rect 3445 -1395 4895 -1390
rect 3445 -1435 3450 -1395
rect 3490 -1435 3800 -1395
rect 3840 -1435 4150 -1395
rect 4190 -1435 4500 -1395
rect 4540 -1435 4850 -1395
rect 4890 -1435 4895 -1395
rect 3445 -1440 4895 -1435
rect 4145 -1740 4195 -1440
rect 995 -1745 4895 -1740
rect 995 -1785 1000 -1745
rect 1040 -1785 1350 -1745
rect 1390 -1785 1700 -1745
rect 1740 -1785 2050 -1745
rect 2090 -1785 2400 -1745
rect 2440 -1785 2750 -1745
rect 2790 -1785 3100 -1745
rect 3140 -1785 3450 -1745
rect 3490 -1785 3800 -1745
rect 3840 -1785 4150 -1745
rect 4190 -1785 4500 -1745
rect 4540 -1785 4850 -1745
rect 4890 -1785 4895 -1745
rect 995 -1790 4895 -1785
rect 995 -2095 1045 -1790
rect 995 -2135 1000 -2095
rect 1040 -2135 1045 -2095
rect 995 -2140 1045 -2135
rect 1345 -2095 1395 -1790
rect 1345 -2135 1350 -2095
rect 1390 -2135 1395 -2095
rect 1345 -2140 1395 -2135
rect 1695 -2095 1745 -1790
rect 1695 -2135 1700 -2095
rect 1740 -2135 1745 -2095
rect 1695 -2140 1745 -2135
rect 2045 -2095 2095 -1790
rect 2045 -2135 2050 -2095
rect 2090 -2135 2095 -2095
rect 2045 -2140 2095 -2135
rect 2395 -2095 2445 -1790
rect 2395 -2135 2400 -2095
rect 2440 -2135 2445 -2095
rect 2395 -2140 2445 -2135
rect 2745 -2095 2795 -1790
rect 2745 -2135 2750 -2095
rect 2790 -2135 2795 -2095
rect 2745 -2140 2795 -2135
rect 3095 -2095 3145 -1790
rect 3095 -2135 3100 -2095
rect 3140 -2135 3145 -2095
rect 3095 -2140 3145 -2135
rect 3445 -2095 3495 -1790
rect 3445 -2135 3450 -2095
rect 3490 -2135 3495 -2095
rect 3445 -2140 3495 -2135
rect 3795 -2095 3845 -1790
rect 3795 -2135 3800 -2095
rect 3840 -2135 3845 -2095
rect 3795 -2140 3845 -2135
rect 4145 -2090 4195 -1790
rect 4145 -2095 4895 -2090
rect 4145 -2135 4150 -2095
rect 4190 -2135 4500 -2095
rect 4540 -2135 4850 -2095
rect 4890 -2135 4895 -2095
rect 4145 -2140 4895 -2135
rect -3850 -2420 5140 -2415
rect -3850 -2460 825 -2420
rect 865 -2460 5140 -2420
rect -3850 -2465 5140 -2460
<< labels >>
flabel metal1 3210 -335 3210 -335 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal3 3100 1595 3100 1595 7 FreeSans 240 0 -80 0 cap_res_X
flabel metal1 -1520 -335 -1520 -335 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal3 -1410 1610 -1410 1610 3 FreeSans 240 0 80 0 cap_res_Y
flabel metal4 -3850 4260 -3850 4260 7 FreeSans 240 0 -80 0 VDDA
port 1 w
flabel metal4 -3850 -2440 -3850 -2440 7 FreeSans 240 0 -80 0 GNDA
port 16 w
flabel metal1 320 1655 320 1655 7 FreeSans 240 0 -80 0 Vb2
port 5 w
flabel metal2 1310 2775 1310 2775 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 400 2775 400 2775 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 1125 1520 1125 1520 3 FreeSans 240 0 80 0 V_err_p
flabel metal1 565 1520 565 1520 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal2 310 1140 310 1140 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 1525 1100 1525 1100 1 FreeSans 240 0 0 160 V_tot
flabel metal2 1070 1200 1070 1200 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 945 1045 945 1045 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal1 2940 400 2940 400 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 2895 290 2895 290 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal1 2040 305 2040 305 5 FreeSans 240 0 0 -80 X
flabel metal1 2495 1610 2495 1610 3 FreeSans 240 0 80 0 Vb3
port 4 e
flabel metal1 -1250 400 -1250 400 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 -1205 290 -1205 290 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 -350 305 -350 305 5 FreeSans 240 0 0 -80 Y
flabel metal2 845 900 845 900 1 FreeSans 240 0 0 80 Vb1
port 6 n
flabel metal2 1795 490 1795 490 3 FreeSans 240 0 80 0 VIN-
port 15 e
flabel metal1 1455 580 1455 580 3 FreeSans 240 0 80 0 VD1
flabel metal2 -105 490 -105 490 7 FreeSans 240 0 -80 0 VIN+
port 14 w
flabel metal1 235 580 235 580 7 FreeSans 240 0 -80 0 VD2
flabel metal1 910 50 910 50 3 FreeSans 240 0 80 0 V_p_mir
flabel metal1 1290 -140 1290 -140 3 FreeSans 240 0 80 0 V_source
flabel metal2 1570 -380 1570 -380 5 FreeSans 240 0 0 -80 V_b_2nd_stage
flabel metal1 -280 2135 -280 2135 7 FreeSans 240 0 -80 0 VD4
flabel metal1 1970 2135 1970 2135 3 FreeSans 240 0 80 0 VD3
flabel metal2 1470 1000 1470 1000 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 965 -1135 965 -1135 3 FreeSans 240 0 80 0 Vb1_2
flabel metal2 460 20 460 20 1 FreeSans 240 0 0 80 V_tail_gate
port 11 n
<< end >>
