magic
tech sky130A
timestamp 1752484787
<< nwell >>
rect 16180 1110 16560 1250
rect 16750 1110 17240 1250
rect 17555 1010 18045 1250
rect 18360 1110 18850 1250
rect 16375 545 16760 685
rect 16910 445 18690 785
rect 18895 495 19220 735
rect 16360 -45 17725 95
rect 17880 -45 19240 95
<< pwell >>
rect 17780 -4300 17820 -4120
<< nmos >>
rect 16890 -350 16910 -300
rect 16950 -350 16970 -300
rect 17010 -350 17030 -300
rect 17070 -350 17090 -300
rect 17130 -350 17150 -300
rect 17190 -350 17210 -300
rect 17250 -350 17270 -300
rect 17310 -350 17330 -300
rect 17370 -350 17390 -300
rect 17430 -350 17450 -300
rect 18150 -350 18170 -300
rect 18210 -350 18230 -300
rect 18270 -350 18290 -300
rect 18330 -350 18350 -300
rect 18390 -350 18410 -300
rect 18450 -350 18470 -300
rect 18510 -350 18530 -300
rect 18570 -350 18590 -300
rect 18630 -350 18650 -300
rect 18690 -350 18710 -300
rect 16570 -825 17070 -575
rect 17190 -825 17690 -575
rect 17910 -825 18410 -575
rect 18530 -825 19030 -575
rect 16780 -1145 17780 -1045
rect 17820 -1145 18820 -1045
rect 16930 -1420 16945 -1320
rect 16985 -1420 17000 -1320
rect 17040 -1420 17055 -1320
rect 17095 -1420 17110 -1320
rect 17150 -1420 17165 -1320
rect 17205 -1420 17220 -1320
rect 17260 -1420 17275 -1320
rect 17315 -1420 17330 -1320
rect 17545 -1420 17560 -1320
rect 17600 -1420 17615 -1320
rect 17655 -1420 17670 -1320
rect 17710 -1420 17725 -1320
rect 17765 -1420 17780 -1320
rect 17820 -1420 17835 -1320
rect 17875 -1420 17890 -1320
rect 17930 -1420 17945 -1320
rect 17985 -1420 18000 -1320
rect 18040 -1420 18055 -1320
rect 18270 -1420 18285 -1320
rect 18325 -1420 18340 -1320
rect 18380 -1420 18395 -1320
rect 18435 -1420 18450 -1320
rect 18490 -1420 18505 -1320
rect 18545 -1420 18560 -1320
rect 18600 -1420 18615 -1320
rect 18655 -1420 18670 -1320
<< pmos >>
rect 16280 1130 16295 1230
rect 16335 1130 16350 1230
rect 16390 1130 16405 1230
rect 16445 1130 16460 1230
rect 16850 1130 16865 1230
rect 16905 1130 16920 1230
rect 16960 1130 16975 1230
rect 17015 1130 17030 1230
rect 17070 1130 17085 1230
rect 17125 1130 17140 1230
rect 17655 1030 17670 1230
rect 17710 1030 17725 1230
rect 17765 1030 17780 1230
rect 17820 1030 17835 1230
rect 17875 1030 17890 1230
rect 17930 1030 17945 1230
rect 18460 1130 18475 1230
rect 18515 1130 18530 1230
rect 18570 1130 18585 1230
rect 18625 1130 18640 1230
rect 18680 1130 18695 1230
rect 18735 1130 18750 1230
rect 16475 565 16490 665
rect 16530 565 16545 665
rect 16585 565 16600 665
rect 16640 565 16655 665
rect 17010 465 17060 765
rect 17100 465 17150 765
rect 17190 465 17240 765
rect 17280 465 17330 765
rect 17370 465 17420 765
rect 17460 465 17510 765
rect 17550 465 17600 765
rect 17640 465 17690 765
rect 17730 465 17780 765
rect 17820 465 17870 765
rect 17910 465 17960 765
rect 18000 465 18050 765
rect 18090 465 18140 765
rect 18180 465 18230 765
rect 18270 465 18320 765
rect 18360 465 18410 765
rect 18450 465 18500 765
rect 18540 465 18590 765
rect 18995 515 19010 715
rect 19050 515 19065 715
rect 19105 515 19120 715
rect 16460 -25 16480 75
rect 16520 -25 16540 75
rect 16580 -25 16600 75
rect 16640 -25 16660 75
rect 16700 -25 16720 75
rect 16760 -25 16780 75
rect 16820 -25 16840 75
rect 16880 -25 16900 75
rect 16940 -25 16960 75
rect 17000 -25 17020 75
rect 17060 -25 17080 75
rect 17120 -25 17140 75
rect 17180 -25 17200 75
rect 17240 -25 17260 75
rect 17300 -25 17320 75
rect 17360 -25 17380 75
rect 17420 -25 17440 75
rect 17480 -25 17500 75
rect 17540 -25 17560 75
rect 17600 -25 17620 75
rect 17980 -25 18000 75
rect 18040 -25 18060 75
rect 18100 -25 18120 75
rect 18160 -25 18180 75
rect 18220 -25 18240 75
rect 18280 -25 18300 75
rect 18340 -25 18360 75
rect 18400 -25 18420 75
rect 18460 -25 18480 75
rect 18520 -25 18540 75
rect 18580 -25 18600 75
rect 18640 -25 18660 75
rect 18700 -25 18720 75
rect 18760 -25 18780 75
rect 18820 -25 18840 75
rect 18880 -25 18900 75
rect 18940 -25 18960 75
rect 19000 -25 19020 75
rect 19060 -25 19080 75
rect 19120 -25 19140 75
<< ndiff >>
rect 16850 -315 16890 -300
rect 16850 -335 16860 -315
rect 16880 -335 16890 -315
rect 16850 -350 16890 -335
rect 16910 -315 16950 -300
rect 16910 -335 16920 -315
rect 16940 -335 16950 -315
rect 16910 -350 16950 -335
rect 16970 -315 17010 -300
rect 16970 -335 16980 -315
rect 17000 -335 17010 -315
rect 16970 -350 17010 -335
rect 17030 -315 17070 -300
rect 17030 -335 17040 -315
rect 17060 -335 17070 -315
rect 17030 -350 17070 -335
rect 17090 -315 17130 -300
rect 17090 -335 17100 -315
rect 17120 -335 17130 -315
rect 17090 -350 17130 -335
rect 17150 -315 17190 -300
rect 17150 -335 17160 -315
rect 17180 -335 17190 -315
rect 17150 -350 17190 -335
rect 17210 -315 17250 -300
rect 17210 -335 17220 -315
rect 17240 -335 17250 -315
rect 17210 -350 17250 -335
rect 17270 -315 17310 -300
rect 17270 -335 17280 -315
rect 17300 -335 17310 -315
rect 17270 -350 17310 -335
rect 17330 -315 17370 -300
rect 17330 -335 17340 -315
rect 17360 -335 17370 -315
rect 17330 -350 17370 -335
rect 17390 -315 17430 -300
rect 17390 -335 17400 -315
rect 17420 -335 17430 -315
rect 17390 -350 17430 -335
rect 17450 -315 17490 -300
rect 17450 -335 17460 -315
rect 17480 -335 17490 -315
rect 17450 -350 17490 -335
rect 18110 -315 18150 -300
rect 18110 -335 18120 -315
rect 18140 -335 18150 -315
rect 18110 -350 18150 -335
rect 18170 -315 18210 -300
rect 18170 -335 18180 -315
rect 18200 -335 18210 -315
rect 18170 -350 18210 -335
rect 18230 -315 18270 -300
rect 18230 -335 18240 -315
rect 18260 -335 18270 -315
rect 18230 -350 18270 -335
rect 18290 -315 18330 -300
rect 18290 -335 18300 -315
rect 18320 -335 18330 -315
rect 18290 -350 18330 -335
rect 18350 -315 18390 -300
rect 18350 -335 18360 -315
rect 18380 -335 18390 -315
rect 18350 -350 18390 -335
rect 18410 -315 18450 -300
rect 18410 -335 18420 -315
rect 18440 -335 18450 -315
rect 18410 -350 18450 -335
rect 18470 -315 18510 -300
rect 18470 -335 18480 -315
rect 18500 -335 18510 -315
rect 18470 -350 18510 -335
rect 18530 -315 18570 -300
rect 18530 -335 18540 -315
rect 18560 -335 18570 -315
rect 18530 -350 18570 -335
rect 18590 -315 18630 -300
rect 18590 -335 18600 -315
rect 18620 -335 18630 -315
rect 18590 -350 18630 -335
rect 18650 -315 18690 -300
rect 18650 -335 18660 -315
rect 18680 -335 18690 -315
rect 18650 -350 18690 -335
rect 18710 -315 18750 -300
rect 18710 -335 18720 -315
rect 18740 -335 18750 -315
rect 18710 -350 18750 -335
rect 16530 -590 16570 -575
rect 16530 -610 16540 -590
rect 16560 -610 16570 -590
rect 16530 -640 16570 -610
rect 16530 -660 16540 -640
rect 16560 -660 16570 -640
rect 16530 -690 16570 -660
rect 16530 -710 16540 -690
rect 16560 -710 16570 -690
rect 16530 -740 16570 -710
rect 16530 -760 16540 -740
rect 16560 -760 16570 -740
rect 16530 -790 16570 -760
rect 16530 -810 16540 -790
rect 16560 -810 16570 -790
rect 16530 -825 16570 -810
rect 17070 -590 17110 -575
rect 17150 -590 17190 -575
rect 17070 -610 17080 -590
rect 17100 -610 17110 -590
rect 17150 -610 17160 -590
rect 17180 -610 17190 -590
rect 17070 -640 17110 -610
rect 17150 -640 17190 -610
rect 17070 -660 17080 -640
rect 17100 -660 17110 -640
rect 17150 -660 17160 -640
rect 17180 -660 17190 -640
rect 17070 -690 17110 -660
rect 17150 -690 17190 -660
rect 17070 -710 17080 -690
rect 17100 -710 17110 -690
rect 17150 -710 17160 -690
rect 17180 -710 17190 -690
rect 17070 -740 17110 -710
rect 17150 -740 17190 -710
rect 17070 -760 17080 -740
rect 17100 -760 17110 -740
rect 17150 -760 17160 -740
rect 17180 -760 17190 -740
rect 17070 -790 17110 -760
rect 17150 -790 17190 -760
rect 17070 -810 17080 -790
rect 17100 -810 17110 -790
rect 17150 -810 17160 -790
rect 17180 -810 17190 -790
rect 17070 -820 17110 -810
rect 17150 -820 17190 -810
rect 17070 -825 17190 -820
rect 17690 -590 17730 -575
rect 17690 -610 17700 -590
rect 17720 -610 17730 -590
rect 17690 -640 17730 -610
rect 17690 -660 17700 -640
rect 17720 -660 17730 -640
rect 17690 -690 17730 -660
rect 17690 -710 17700 -690
rect 17720 -710 17730 -690
rect 17690 -740 17730 -710
rect 17690 -760 17700 -740
rect 17720 -760 17730 -740
rect 17690 -790 17730 -760
rect 17690 -810 17700 -790
rect 17720 -810 17730 -790
rect 17690 -825 17730 -810
rect 17870 -590 17910 -575
rect 17870 -610 17880 -590
rect 17900 -610 17910 -590
rect 17870 -640 17910 -610
rect 17870 -660 17880 -640
rect 17900 -660 17910 -640
rect 17870 -690 17910 -660
rect 17870 -710 17880 -690
rect 17900 -710 17910 -690
rect 17870 -740 17910 -710
rect 17870 -760 17880 -740
rect 17900 -760 17910 -740
rect 17870 -790 17910 -760
rect 17870 -810 17880 -790
rect 17900 -810 17910 -790
rect 17870 -825 17910 -810
rect 18410 -590 18450 -575
rect 18490 -590 18530 -575
rect 18410 -610 18420 -590
rect 18440 -610 18450 -590
rect 18490 -610 18500 -590
rect 18520 -610 18530 -590
rect 18410 -640 18450 -610
rect 18490 -640 18530 -610
rect 18410 -660 18420 -640
rect 18440 -660 18450 -640
rect 18490 -660 18500 -640
rect 18520 -660 18530 -640
rect 18410 -690 18450 -660
rect 18490 -690 18530 -660
rect 18410 -710 18420 -690
rect 18440 -710 18450 -690
rect 18490 -710 18500 -690
rect 18520 -710 18530 -690
rect 18410 -740 18450 -710
rect 18490 -740 18530 -710
rect 18410 -760 18420 -740
rect 18440 -760 18450 -740
rect 18490 -760 18500 -740
rect 18520 -760 18530 -740
rect 18410 -790 18450 -760
rect 18490 -790 18530 -760
rect 18410 -810 18420 -790
rect 18440 -810 18450 -790
rect 18490 -810 18500 -790
rect 18520 -810 18530 -790
rect 18410 -825 18450 -810
rect 18490 -825 18530 -810
rect 19030 -590 19070 -575
rect 19030 -610 19040 -590
rect 19060 -610 19070 -590
rect 19030 -640 19070 -610
rect 19030 -660 19040 -640
rect 19060 -660 19070 -640
rect 19030 -690 19070 -660
rect 19030 -710 19040 -690
rect 19060 -710 19070 -690
rect 19030 -740 19070 -710
rect 19030 -760 19040 -740
rect 19060 -760 19070 -740
rect 19030 -790 19070 -760
rect 19030 -810 19040 -790
rect 19060 -810 19070 -790
rect 19030 -825 19070 -810
rect 16740 -1060 16780 -1045
rect 16740 -1080 16750 -1060
rect 16770 -1080 16780 -1060
rect 16740 -1110 16780 -1080
rect 16740 -1130 16750 -1110
rect 16770 -1130 16780 -1110
rect 16740 -1145 16780 -1130
rect 17780 -1060 17820 -1045
rect 17780 -1080 17790 -1060
rect 17810 -1080 17820 -1060
rect 17780 -1110 17820 -1080
rect 17780 -1130 17790 -1110
rect 17810 -1130 17820 -1110
rect 17780 -1145 17820 -1130
rect 18820 -1060 18860 -1045
rect 18820 -1080 18830 -1060
rect 18850 -1080 18860 -1060
rect 18820 -1110 18860 -1080
rect 18820 -1130 18830 -1110
rect 18850 -1130 18860 -1110
rect 18820 -1145 18860 -1130
rect 16890 -1335 16930 -1320
rect 16890 -1355 16900 -1335
rect 16920 -1355 16930 -1335
rect 16890 -1385 16930 -1355
rect 16890 -1405 16900 -1385
rect 16920 -1405 16930 -1385
rect 16890 -1420 16930 -1405
rect 16945 -1335 16985 -1320
rect 16945 -1355 16955 -1335
rect 16975 -1355 16985 -1335
rect 16945 -1385 16985 -1355
rect 16945 -1405 16955 -1385
rect 16975 -1405 16985 -1385
rect 16945 -1420 16985 -1405
rect 17000 -1335 17040 -1320
rect 17000 -1355 17010 -1335
rect 17030 -1355 17040 -1335
rect 17000 -1385 17040 -1355
rect 17000 -1405 17010 -1385
rect 17030 -1405 17040 -1385
rect 17000 -1420 17040 -1405
rect 17055 -1335 17095 -1320
rect 17055 -1355 17065 -1335
rect 17085 -1355 17095 -1335
rect 17055 -1385 17095 -1355
rect 17055 -1405 17065 -1385
rect 17085 -1405 17095 -1385
rect 17055 -1420 17095 -1405
rect 17110 -1335 17150 -1320
rect 17110 -1355 17120 -1335
rect 17140 -1355 17150 -1335
rect 17110 -1385 17150 -1355
rect 17110 -1405 17120 -1385
rect 17140 -1405 17150 -1385
rect 17110 -1420 17150 -1405
rect 17165 -1335 17205 -1320
rect 17165 -1355 17175 -1335
rect 17195 -1355 17205 -1335
rect 17165 -1385 17205 -1355
rect 17165 -1405 17175 -1385
rect 17195 -1405 17205 -1385
rect 17165 -1420 17205 -1405
rect 17220 -1335 17260 -1320
rect 17220 -1355 17230 -1335
rect 17250 -1355 17260 -1335
rect 17220 -1385 17260 -1355
rect 17220 -1405 17230 -1385
rect 17250 -1405 17260 -1385
rect 17220 -1420 17260 -1405
rect 17275 -1335 17315 -1320
rect 17275 -1355 17285 -1335
rect 17305 -1355 17315 -1335
rect 17275 -1385 17315 -1355
rect 17275 -1405 17285 -1385
rect 17305 -1405 17315 -1385
rect 17275 -1420 17315 -1405
rect 17330 -1335 17370 -1320
rect 17330 -1355 17340 -1335
rect 17360 -1355 17370 -1335
rect 17330 -1385 17370 -1355
rect 17330 -1405 17340 -1385
rect 17360 -1405 17370 -1385
rect 17330 -1420 17370 -1405
rect 17505 -1335 17545 -1320
rect 17505 -1355 17515 -1335
rect 17535 -1355 17545 -1335
rect 17505 -1385 17545 -1355
rect 17505 -1405 17515 -1385
rect 17535 -1405 17545 -1385
rect 17505 -1420 17545 -1405
rect 17560 -1335 17600 -1320
rect 17560 -1355 17570 -1335
rect 17590 -1355 17600 -1335
rect 17560 -1385 17600 -1355
rect 17560 -1405 17570 -1385
rect 17590 -1405 17600 -1385
rect 17560 -1420 17600 -1405
rect 17615 -1335 17655 -1320
rect 17615 -1355 17625 -1335
rect 17645 -1355 17655 -1335
rect 17615 -1385 17655 -1355
rect 17615 -1405 17625 -1385
rect 17645 -1405 17655 -1385
rect 17615 -1420 17655 -1405
rect 17670 -1335 17710 -1320
rect 17670 -1355 17680 -1335
rect 17700 -1355 17710 -1335
rect 17670 -1385 17710 -1355
rect 17670 -1405 17680 -1385
rect 17700 -1405 17710 -1385
rect 17670 -1420 17710 -1405
rect 17725 -1335 17765 -1320
rect 17725 -1355 17735 -1335
rect 17755 -1355 17765 -1335
rect 17725 -1385 17765 -1355
rect 17725 -1405 17735 -1385
rect 17755 -1405 17765 -1385
rect 17725 -1420 17765 -1405
rect 17780 -1335 17820 -1320
rect 17780 -1355 17790 -1335
rect 17810 -1355 17820 -1335
rect 17780 -1385 17820 -1355
rect 17780 -1405 17790 -1385
rect 17810 -1405 17820 -1385
rect 17780 -1420 17820 -1405
rect 17835 -1335 17875 -1320
rect 17835 -1355 17845 -1335
rect 17865 -1355 17875 -1335
rect 17835 -1385 17875 -1355
rect 17835 -1405 17845 -1385
rect 17865 -1405 17875 -1385
rect 17835 -1420 17875 -1405
rect 17890 -1335 17930 -1320
rect 17890 -1355 17900 -1335
rect 17920 -1355 17930 -1335
rect 17890 -1385 17930 -1355
rect 17890 -1405 17900 -1385
rect 17920 -1405 17930 -1385
rect 17890 -1420 17930 -1405
rect 17945 -1335 17985 -1320
rect 17945 -1355 17955 -1335
rect 17975 -1355 17985 -1335
rect 17945 -1385 17985 -1355
rect 17945 -1405 17955 -1385
rect 17975 -1405 17985 -1385
rect 17945 -1420 17985 -1405
rect 18000 -1335 18040 -1320
rect 18000 -1355 18010 -1335
rect 18030 -1355 18040 -1335
rect 18000 -1385 18040 -1355
rect 18000 -1405 18010 -1385
rect 18030 -1405 18040 -1385
rect 18000 -1420 18040 -1405
rect 18055 -1335 18095 -1320
rect 18055 -1355 18065 -1335
rect 18085 -1355 18095 -1335
rect 18055 -1385 18095 -1355
rect 18055 -1405 18065 -1385
rect 18085 -1405 18095 -1385
rect 18055 -1420 18095 -1405
rect 18230 -1335 18270 -1320
rect 18230 -1355 18240 -1335
rect 18260 -1355 18270 -1335
rect 18230 -1385 18270 -1355
rect 18230 -1405 18240 -1385
rect 18260 -1405 18270 -1385
rect 18230 -1420 18270 -1405
rect 18285 -1335 18325 -1320
rect 18285 -1355 18295 -1335
rect 18315 -1355 18325 -1335
rect 18285 -1385 18325 -1355
rect 18285 -1405 18295 -1385
rect 18315 -1405 18325 -1385
rect 18285 -1420 18325 -1405
rect 18340 -1335 18380 -1320
rect 18340 -1355 18350 -1335
rect 18370 -1355 18380 -1335
rect 18340 -1385 18380 -1355
rect 18340 -1405 18350 -1385
rect 18370 -1405 18380 -1385
rect 18340 -1420 18380 -1405
rect 18395 -1335 18435 -1320
rect 18395 -1355 18405 -1335
rect 18425 -1355 18435 -1335
rect 18395 -1385 18435 -1355
rect 18395 -1405 18405 -1385
rect 18425 -1405 18435 -1385
rect 18395 -1420 18435 -1405
rect 18450 -1335 18490 -1320
rect 18450 -1355 18460 -1335
rect 18480 -1355 18490 -1335
rect 18450 -1385 18490 -1355
rect 18450 -1405 18460 -1385
rect 18480 -1405 18490 -1385
rect 18450 -1420 18490 -1405
rect 18505 -1335 18545 -1320
rect 18505 -1355 18515 -1335
rect 18535 -1355 18545 -1335
rect 18505 -1385 18545 -1355
rect 18505 -1405 18515 -1385
rect 18535 -1405 18545 -1385
rect 18505 -1420 18545 -1405
rect 18560 -1335 18600 -1320
rect 18560 -1355 18570 -1335
rect 18590 -1355 18600 -1335
rect 18560 -1385 18600 -1355
rect 18560 -1405 18570 -1385
rect 18590 -1405 18600 -1385
rect 18560 -1420 18600 -1405
rect 18615 -1335 18655 -1320
rect 18615 -1355 18625 -1335
rect 18645 -1355 18655 -1335
rect 18615 -1385 18655 -1355
rect 18615 -1405 18625 -1385
rect 18645 -1405 18655 -1385
rect 18615 -1420 18655 -1405
rect 18670 -1335 18710 -1320
rect 18670 -1355 18680 -1335
rect 18700 -1355 18710 -1335
rect 18670 -1385 18710 -1355
rect 18670 -1405 18680 -1385
rect 18700 -1405 18710 -1385
rect 18670 -1420 18710 -1405
<< pdiff >>
rect 16240 1215 16280 1230
rect 16240 1143 16250 1215
rect 16270 1143 16280 1215
rect 16240 1130 16280 1143
rect 16295 1215 16335 1230
rect 16295 1143 16305 1215
rect 16325 1143 16335 1215
rect 16295 1130 16335 1143
rect 16350 1215 16390 1230
rect 16350 1143 16360 1215
rect 16380 1143 16390 1215
rect 16350 1130 16390 1143
rect 16405 1215 16445 1230
rect 16405 1143 16415 1215
rect 16435 1143 16445 1215
rect 16405 1130 16445 1143
rect 16460 1215 16500 1230
rect 16460 1143 16470 1215
rect 16490 1143 16500 1215
rect 16460 1130 16500 1143
rect 16810 1215 16850 1230
rect 16810 1143 16820 1215
rect 16840 1143 16850 1215
rect 16810 1130 16850 1143
rect 16865 1215 16905 1230
rect 16865 1143 16875 1215
rect 16895 1143 16905 1215
rect 16865 1130 16905 1143
rect 16920 1215 16960 1230
rect 16920 1143 16930 1215
rect 16950 1143 16960 1215
rect 16920 1130 16960 1143
rect 16975 1215 17015 1230
rect 16975 1143 16985 1215
rect 17005 1143 17015 1215
rect 16975 1130 17015 1143
rect 17030 1215 17070 1230
rect 17030 1143 17040 1215
rect 17060 1143 17070 1215
rect 17030 1130 17070 1143
rect 17085 1215 17125 1230
rect 17085 1143 17095 1215
rect 17115 1143 17125 1215
rect 17085 1130 17125 1143
rect 17140 1215 17180 1230
rect 17140 1143 17150 1215
rect 17170 1143 17180 1215
rect 17140 1130 17180 1143
rect 17615 1215 17655 1230
rect 17615 1195 17625 1215
rect 17645 1195 17655 1215
rect 17615 1165 17655 1195
rect 17615 1145 17625 1165
rect 17645 1145 17655 1165
rect 17615 1115 17655 1145
rect 17615 1095 17625 1115
rect 17645 1095 17655 1115
rect 17615 1065 17655 1095
rect 17615 1045 17625 1065
rect 17645 1045 17655 1065
rect 17615 1030 17655 1045
rect 17670 1215 17710 1230
rect 17670 1195 17680 1215
rect 17700 1195 17710 1215
rect 17670 1165 17710 1195
rect 17670 1145 17680 1165
rect 17700 1145 17710 1165
rect 17670 1115 17710 1145
rect 17670 1095 17680 1115
rect 17700 1095 17710 1115
rect 17670 1065 17710 1095
rect 17670 1045 17680 1065
rect 17700 1045 17710 1065
rect 17670 1030 17710 1045
rect 17725 1215 17765 1230
rect 17725 1195 17735 1215
rect 17755 1195 17765 1215
rect 17725 1165 17765 1195
rect 17725 1145 17735 1165
rect 17755 1145 17765 1165
rect 17725 1115 17765 1145
rect 17725 1095 17735 1115
rect 17755 1095 17765 1115
rect 17725 1065 17765 1095
rect 17725 1045 17735 1065
rect 17755 1045 17765 1065
rect 17725 1030 17765 1045
rect 17780 1215 17820 1230
rect 17780 1195 17790 1215
rect 17810 1195 17820 1215
rect 17780 1165 17820 1195
rect 17780 1145 17790 1165
rect 17810 1145 17820 1165
rect 17780 1115 17820 1145
rect 17780 1095 17790 1115
rect 17810 1095 17820 1115
rect 17780 1065 17820 1095
rect 17780 1045 17790 1065
rect 17810 1045 17820 1065
rect 17780 1030 17820 1045
rect 17835 1215 17875 1230
rect 17835 1195 17845 1215
rect 17865 1195 17875 1215
rect 17835 1165 17875 1195
rect 17835 1145 17845 1165
rect 17865 1145 17875 1165
rect 17835 1115 17875 1145
rect 17835 1095 17845 1115
rect 17865 1095 17875 1115
rect 17835 1065 17875 1095
rect 17835 1045 17845 1065
rect 17865 1045 17875 1065
rect 17835 1030 17875 1045
rect 17890 1215 17930 1230
rect 17890 1195 17900 1215
rect 17920 1195 17930 1215
rect 17890 1165 17930 1195
rect 17890 1145 17900 1165
rect 17920 1145 17930 1165
rect 17890 1115 17930 1145
rect 17890 1095 17900 1115
rect 17920 1095 17930 1115
rect 17890 1065 17930 1095
rect 17890 1045 17900 1065
rect 17920 1045 17930 1065
rect 17890 1030 17930 1045
rect 17945 1215 17985 1230
rect 17945 1195 17955 1215
rect 17975 1195 17985 1215
rect 17945 1165 17985 1195
rect 17945 1145 17955 1165
rect 17975 1145 17985 1165
rect 17945 1115 17985 1145
rect 18420 1215 18460 1230
rect 18420 1145 18430 1215
rect 18450 1145 18460 1215
rect 18420 1130 18460 1145
rect 18475 1215 18515 1230
rect 18475 1145 18485 1215
rect 18505 1145 18515 1215
rect 18475 1130 18515 1145
rect 18530 1215 18570 1230
rect 18530 1145 18540 1215
rect 18560 1145 18570 1215
rect 18530 1130 18570 1145
rect 18585 1215 18625 1230
rect 18585 1145 18595 1215
rect 18615 1145 18625 1215
rect 18585 1130 18625 1145
rect 18640 1215 18680 1230
rect 18640 1145 18650 1215
rect 18670 1145 18680 1215
rect 18640 1130 18680 1145
rect 18695 1215 18735 1230
rect 18695 1145 18705 1215
rect 18725 1145 18735 1215
rect 18695 1130 18735 1145
rect 18750 1215 18790 1230
rect 18750 1145 18760 1215
rect 18780 1145 18790 1215
rect 18750 1130 18790 1145
rect 17945 1095 17955 1115
rect 17975 1095 17985 1115
rect 17945 1065 17985 1095
rect 17945 1045 17955 1065
rect 17975 1045 17985 1065
rect 17945 1030 17985 1045
rect 16970 750 17010 765
rect 16970 730 16980 750
rect 17000 730 17010 750
rect 16970 700 17010 730
rect 16970 680 16980 700
rect 17000 680 17010 700
rect 16435 650 16475 665
rect 16435 630 16445 650
rect 16465 630 16475 650
rect 16435 600 16475 630
rect 16435 580 16445 600
rect 16465 580 16475 600
rect 16435 565 16475 580
rect 16490 650 16530 665
rect 16490 630 16500 650
rect 16520 630 16530 650
rect 16490 600 16530 630
rect 16490 580 16500 600
rect 16520 580 16530 600
rect 16490 565 16530 580
rect 16545 650 16585 665
rect 16545 630 16555 650
rect 16575 630 16585 650
rect 16545 600 16585 630
rect 16545 580 16555 600
rect 16575 580 16585 600
rect 16545 565 16585 580
rect 16600 650 16640 665
rect 16600 630 16610 650
rect 16630 630 16640 650
rect 16600 600 16640 630
rect 16600 580 16610 600
rect 16630 580 16640 600
rect 16600 565 16640 580
rect 16655 650 16700 665
rect 16655 630 16665 650
rect 16685 630 16700 650
rect 16655 600 16700 630
rect 16655 580 16665 600
rect 16685 580 16700 600
rect 16655 565 16700 580
rect 16970 650 17010 680
rect 16970 630 16980 650
rect 17000 630 17010 650
rect 16970 600 17010 630
rect 16970 580 16980 600
rect 17000 580 17010 600
rect 16970 550 17010 580
rect 16970 530 16980 550
rect 17000 530 17010 550
rect 16970 500 17010 530
rect 16970 480 16980 500
rect 17000 480 17010 500
rect 16970 465 17010 480
rect 17060 750 17100 765
rect 17060 730 17070 750
rect 17090 730 17100 750
rect 17060 700 17100 730
rect 17060 680 17070 700
rect 17090 680 17100 700
rect 17060 650 17100 680
rect 17060 630 17070 650
rect 17090 630 17100 650
rect 17060 600 17100 630
rect 17060 580 17070 600
rect 17090 580 17100 600
rect 17060 550 17100 580
rect 17060 530 17070 550
rect 17090 530 17100 550
rect 17060 500 17100 530
rect 17060 480 17070 500
rect 17090 480 17100 500
rect 17060 465 17100 480
rect 17150 750 17190 765
rect 17150 730 17160 750
rect 17180 730 17190 750
rect 17150 700 17190 730
rect 17150 680 17160 700
rect 17180 680 17190 700
rect 17150 650 17190 680
rect 17150 630 17160 650
rect 17180 630 17190 650
rect 17150 600 17190 630
rect 17150 580 17160 600
rect 17180 580 17190 600
rect 17150 550 17190 580
rect 17150 530 17160 550
rect 17180 530 17190 550
rect 17150 500 17190 530
rect 17150 480 17160 500
rect 17180 480 17190 500
rect 17150 465 17190 480
rect 17240 750 17280 765
rect 17240 730 17250 750
rect 17270 730 17280 750
rect 17240 700 17280 730
rect 17240 680 17250 700
rect 17270 680 17280 700
rect 17240 650 17280 680
rect 17240 630 17250 650
rect 17270 630 17280 650
rect 17240 600 17280 630
rect 17240 580 17250 600
rect 17270 580 17280 600
rect 17240 550 17280 580
rect 17240 530 17250 550
rect 17270 530 17280 550
rect 17240 500 17280 530
rect 17240 480 17250 500
rect 17270 480 17280 500
rect 17240 465 17280 480
rect 17330 750 17370 765
rect 17330 730 17340 750
rect 17360 730 17370 750
rect 17330 700 17370 730
rect 17330 680 17340 700
rect 17360 680 17370 700
rect 17330 650 17370 680
rect 17330 630 17340 650
rect 17360 630 17370 650
rect 17330 600 17370 630
rect 17330 580 17340 600
rect 17360 580 17370 600
rect 17330 550 17370 580
rect 17330 530 17340 550
rect 17360 530 17370 550
rect 17330 500 17370 530
rect 17330 480 17340 500
rect 17360 480 17370 500
rect 17330 465 17370 480
rect 17420 750 17460 765
rect 17420 730 17430 750
rect 17450 730 17460 750
rect 17420 700 17460 730
rect 17420 680 17430 700
rect 17450 680 17460 700
rect 17420 650 17460 680
rect 17420 630 17430 650
rect 17450 630 17460 650
rect 17420 600 17460 630
rect 17420 580 17430 600
rect 17450 580 17460 600
rect 17420 550 17460 580
rect 17420 530 17430 550
rect 17450 530 17460 550
rect 17420 500 17460 530
rect 17420 480 17430 500
rect 17450 480 17460 500
rect 17420 465 17460 480
rect 17510 750 17550 765
rect 17510 730 17520 750
rect 17540 730 17550 750
rect 17510 700 17550 730
rect 17510 680 17520 700
rect 17540 680 17550 700
rect 17510 650 17550 680
rect 17510 630 17520 650
rect 17540 630 17550 650
rect 17510 600 17550 630
rect 17510 580 17520 600
rect 17540 580 17550 600
rect 17510 550 17550 580
rect 17510 530 17520 550
rect 17540 530 17550 550
rect 17510 500 17550 530
rect 17510 480 17520 500
rect 17540 480 17550 500
rect 17510 465 17550 480
rect 17600 750 17640 765
rect 17600 730 17610 750
rect 17630 730 17640 750
rect 17600 700 17640 730
rect 17600 680 17610 700
rect 17630 680 17640 700
rect 17600 650 17640 680
rect 17600 630 17610 650
rect 17630 630 17640 650
rect 17600 600 17640 630
rect 17600 580 17610 600
rect 17630 580 17640 600
rect 17600 550 17640 580
rect 17600 530 17610 550
rect 17630 530 17640 550
rect 17600 500 17640 530
rect 17600 480 17610 500
rect 17630 480 17640 500
rect 17600 465 17640 480
rect 17690 750 17730 765
rect 17690 730 17700 750
rect 17720 730 17730 750
rect 17690 700 17730 730
rect 17690 680 17700 700
rect 17720 680 17730 700
rect 17690 650 17730 680
rect 17690 630 17700 650
rect 17720 630 17730 650
rect 17690 600 17730 630
rect 17690 580 17700 600
rect 17720 580 17730 600
rect 17690 550 17730 580
rect 17690 530 17700 550
rect 17720 530 17730 550
rect 17690 500 17730 530
rect 17690 480 17700 500
rect 17720 480 17730 500
rect 17690 465 17730 480
rect 17780 750 17820 765
rect 17780 730 17790 750
rect 17810 730 17820 750
rect 17780 700 17820 730
rect 17780 680 17790 700
rect 17810 680 17820 700
rect 17780 650 17820 680
rect 17780 630 17790 650
rect 17810 630 17820 650
rect 17780 600 17820 630
rect 17780 580 17790 600
rect 17810 580 17820 600
rect 17780 550 17820 580
rect 17780 530 17790 550
rect 17810 530 17820 550
rect 17780 500 17820 530
rect 17780 480 17790 500
rect 17810 480 17820 500
rect 17780 465 17820 480
rect 17870 750 17910 765
rect 17870 730 17880 750
rect 17900 730 17910 750
rect 17870 700 17910 730
rect 17870 680 17880 700
rect 17900 680 17910 700
rect 17870 650 17910 680
rect 17870 630 17880 650
rect 17900 630 17910 650
rect 17870 600 17910 630
rect 17870 580 17880 600
rect 17900 580 17910 600
rect 17870 550 17910 580
rect 17870 530 17880 550
rect 17900 530 17910 550
rect 17870 500 17910 530
rect 17870 480 17880 500
rect 17900 480 17910 500
rect 17870 465 17910 480
rect 17960 750 18000 765
rect 17960 730 17970 750
rect 17990 730 18000 750
rect 17960 700 18000 730
rect 17960 680 17970 700
rect 17990 680 18000 700
rect 17960 650 18000 680
rect 17960 630 17970 650
rect 17990 630 18000 650
rect 17960 600 18000 630
rect 17960 580 17970 600
rect 17990 580 18000 600
rect 17960 550 18000 580
rect 17960 530 17970 550
rect 17990 530 18000 550
rect 17960 500 18000 530
rect 17960 480 17970 500
rect 17990 480 18000 500
rect 17960 465 18000 480
rect 18050 750 18090 765
rect 18050 730 18060 750
rect 18080 730 18090 750
rect 18050 700 18090 730
rect 18050 680 18060 700
rect 18080 680 18090 700
rect 18050 650 18090 680
rect 18050 630 18060 650
rect 18080 630 18090 650
rect 18050 600 18090 630
rect 18050 580 18060 600
rect 18080 580 18090 600
rect 18050 550 18090 580
rect 18050 530 18060 550
rect 18080 530 18090 550
rect 18050 500 18090 530
rect 18050 480 18060 500
rect 18080 480 18090 500
rect 18050 465 18090 480
rect 18140 750 18180 765
rect 18140 730 18150 750
rect 18170 730 18180 750
rect 18140 700 18180 730
rect 18140 680 18150 700
rect 18170 680 18180 700
rect 18140 650 18180 680
rect 18140 630 18150 650
rect 18170 630 18180 650
rect 18140 600 18180 630
rect 18140 580 18150 600
rect 18170 580 18180 600
rect 18140 550 18180 580
rect 18140 530 18150 550
rect 18170 530 18180 550
rect 18140 500 18180 530
rect 18140 480 18150 500
rect 18170 480 18180 500
rect 18140 465 18180 480
rect 18230 750 18270 765
rect 18230 730 18240 750
rect 18260 730 18270 750
rect 18230 700 18270 730
rect 18230 680 18240 700
rect 18260 680 18270 700
rect 18230 650 18270 680
rect 18230 630 18240 650
rect 18260 630 18270 650
rect 18230 600 18270 630
rect 18230 580 18240 600
rect 18260 580 18270 600
rect 18230 550 18270 580
rect 18230 530 18240 550
rect 18260 530 18270 550
rect 18230 500 18270 530
rect 18230 480 18240 500
rect 18260 480 18270 500
rect 18230 465 18270 480
rect 18320 750 18360 765
rect 18320 730 18330 750
rect 18350 730 18360 750
rect 18320 700 18360 730
rect 18320 680 18330 700
rect 18350 680 18360 700
rect 18320 650 18360 680
rect 18320 630 18330 650
rect 18350 630 18360 650
rect 18320 600 18360 630
rect 18320 580 18330 600
rect 18350 580 18360 600
rect 18320 550 18360 580
rect 18320 530 18330 550
rect 18350 530 18360 550
rect 18320 500 18360 530
rect 18320 480 18330 500
rect 18350 480 18360 500
rect 18320 465 18360 480
rect 18410 750 18450 765
rect 18410 730 18420 750
rect 18440 730 18450 750
rect 18410 700 18450 730
rect 18410 680 18420 700
rect 18440 680 18450 700
rect 18410 650 18450 680
rect 18410 630 18420 650
rect 18440 630 18450 650
rect 18410 600 18450 630
rect 18410 580 18420 600
rect 18440 580 18450 600
rect 18410 550 18450 580
rect 18410 530 18420 550
rect 18440 530 18450 550
rect 18410 500 18450 530
rect 18410 480 18420 500
rect 18440 480 18450 500
rect 18410 465 18450 480
rect 18500 750 18540 765
rect 18500 730 18510 750
rect 18530 730 18540 750
rect 18500 700 18540 730
rect 18500 680 18510 700
rect 18530 680 18540 700
rect 18500 650 18540 680
rect 18500 630 18510 650
rect 18530 630 18540 650
rect 18500 600 18540 630
rect 18500 580 18510 600
rect 18530 580 18540 600
rect 18500 550 18540 580
rect 18500 530 18510 550
rect 18530 530 18540 550
rect 18500 500 18540 530
rect 18500 480 18510 500
rect 18530 480 18540 500
rect 18500 465 18540 480
rect 18590 750 18630 765
rect 18590 730 18600 750
rect 18620 730 18630 750
rect 18590 700 18630 730
rect 18590 680 18600 700
rect 18620 680 18630 700
rect 18590 650 18630 680
rect 18590 630 18600 650
rect 18620 630 18630 650
rect 18590 600 18630 630
rect 18590 580 18600 600
rect 18620 580 18630 600
rect 18590 550 18630 580
rect 18590 530 18600 550
rect 18620 530 18630 550
rect 18590 500 18630 530
rect 18955 700 18995 715
rect 18955 680 18965 700
rect 18985 680 18995 700
rect 18955 650 18995 680
rect 18955 630 18965 650
rect 18985 630 18995 650
rect 18955 600 18995 630
rect 18955 580 18965 600
rect 18985 580 18995 600
rect 18955 550 18995 580
rect 18955 530 18965 550
rect 18985 530 18995 550
rect 18955 515 18995 530
rect 19010 700 19050 715
rect 19010 680 19020 700
rect 19040 680 19050 700
rect 19010 650 19050 680
rect 19010 630 19020 650
rect 19040 630 19050 650
rect 19010 600 19050 630
rect 19010 580 19020 600
rect 19040 580 19050 600
rect 19010 550 19050 580
rect 19010 530 19020 550
rect 19040 530 19050 550
rect 19010 515 19050 530
rect 19065 700 19105 715
rect 19065 680 19075 700
rect 19095 680 19105 700
rect 19065 650 19105 680
rect 19065 630 19075 650
rect 19095 630 19105 650
rect 19065 600 19105 630
rect 19065 580 19075 600
rect 19095 580 19105 600
rect 19065 550 19105 580
rect 19065 530 19075 550
rect 19095 530 19105 550
rect 19065 515 19105 530
rect 19120 700 19160 715
rect 19120 680 19130 700
rect 19150 680 19160 700
rect 19120 650 19160 680
rect 19120 630 19130 650
rect 19150 630 19160 650
rect 19120 600 19160 630
rect 19120 580 19130 600
rect 19150 580 19160 600
rect 19120 550 19160 580
rect 19120 530 19130 550
rect 19150 530 19160 550
rect 19120 515 19160 530
rect 18590 480 18600 500
rect 18620 480 18630 500
rect 18590 465 18630 480
rect 16420 60 16460 75
rect 16420 40 16430 60
rect 16450 40 16460 60
rect 16420 10 16460 40
rect 16420 -10 16430 10
rect 16450 -10 16460 10
rect 16420 -25 16460 -10
rect 16480 60 16520 75
rect 16480 40 16490 60
rect 16510 40 16520 60
rect 16480 10 16520 40
rect 16480 -10 16490 10
rect 16510 -10 16520 10
rect 16480 -25 16520 -10
rect 16540 60 16580 75
rect 16540 40 16550 60
rect 16570 40 16580 60
rect 16540 10 16580 40
rect 16540 -10 16550 10
rect 16570 -10 16580 10
rect 16540 -25 16580 -10
rect 16600 60 16640 75
rect 16600 40 16610 60
rect 16630 40 16640 60
rect 16600 10 16640 40
rect 16600 -10 16610 10
rect 16630 -10 16640 10
rect 16600 -25 16640 -10
rect 16660 60 16700 75
rect 16660 40 16670 60
rect 16690 40 16700 60
rect 16660 10 16700 40
rect 16660 -10 16670 10
rect 16690 -10 16700 10
rect 16660 -25 16700 -10
rect 16720 60 16760 75
rect 16720 40 16730 60
rect 16750 40 16760 60
rect 16720 10 16760 40
rect 16720 -10 16730 10
rect 16750 -10 16760 10
rect 16720 -25 16760 -10
rect 16780 60 16820 75
rect 16780 40 16790 60
rect 16810 40 16820 60
rect 16780 10 16820 40
rect 16780 -10 16790 10
rect 16810 -10 16820 10
rect 16780 -25 16820 -10
rect 16840 60 16880 75
rect 16840 40 16850 60
rect 16870 40 16880 60
rect 16840 10 16880 40
rect 16840 -10 16850 10
rect 16870 -10 16880 10
rect 16840 -25 16880 -10
rect 16900 60 16940 75
rect 16900 40 16910 60
rect 16930 40 16940 60
rect 16900 10 16940 40
rect 16900 -10 16910 10
rect 16930 -10 16940 10
rect 16900 -25 16940 -10
rect 16960 60 17000 75
rect 16960 40 16970 60
rect 16990 40 17000 60
rect 16960 10 17000 40
rect 16960 -10 16970 10
rect 16990 -10 17000 10
rect 16960 -25 17000 -10
rect 17020 60 17060 75
rect 17020 40 17030 60
rect 17050 40 17060 60
rect 17020 10 17060 40
rect 17020 -10 17030 10
rect 17050 -10 17060 10
rect 17020 -25 17060 -10
rect 17080 60 17120 75
rect 17080 40 17090 60
rect 17110 40 17120 60
rect 17080 10 17120 40
rect 17080 -10 17090 10
rect 17110 -10 17120 10
rect 17080 -25 17120 -10
rect 17140 60 17180 75
rect 17140 40 17150 60
rect 17170 40 17180 60
rect 17140 10 17180 40
rect 17140 -10 17150 10
rect 17170 -10 17180 10
rect 17140 -25 17180 -10
rect 17200 60 17240 75
rect 17200 40 17210 60
rect 17230 40 17240 60
rect 17200 10 17240 40
rect 17200 -10 17210 10
rect 17230 -10 17240 10
rect 17200 -25 17240 -10
rect 17260 60 17300 75
rect 17260 40 17270 60
rect 17290 40 17300 60
rect 17260 10 17300 40
rect 17260 -10 17270 10
rect 17290 -10 17300 10
rect 17260 -25 17300 -10
rect 17320 60 17360 75
rect 17320 40 17330 60
rect 17350 40 17360 60
rect 17320 10 17360 40
rect 17320 -10 17330 10
rect 17350 -10 17360 10
rect 17320 -25 17360 -10
rect 17380 60 17420 75
rect 17380 40 17390 60
rect 17410 40 17420 60
rect 17380 10 17420 40
rect 17380 -10 17390 10
rect 17410 -10 17420 10
rect 17380 -25 17420 -10
rect 17440 60 17480 75
rect 17440 40 17450 60
rect 17470 40 17480 60
rect 17440 10 17480 40
rect 17440 -10 17450 10
rect 17470 -10 17480 10
rect 17440 -25 17480 -10
rect 17500 60 17540 75
rect 17500 40 17510 60
rect 17530 40 17540 60
rect 17500 10 17540 40
rect 17500 -10 17510 10
rect 17530 -10 17540 10
rect 17500 -25 17540 -10
rect 17560 60 17600 75
rect 17560 40 17570 60
rect 17590 40 17600 60
rect 17560 10 17600 40
rect 17560 -10 17570 10
rect 17590 -10 17600 10
rect 17560 -25 17600 -10
rect 17620 60 17660 75
rect 17620 40 17630 60
rect 17650 40 17660 60
rect 17620 10 17660 40
rect 17620 -10 17630 10
rect 17650 -10 17660 10
rect 17620 -25 17660 -10
rect 17940 60 17980 75
rect 17940 40 17950 60
rect 17970 40 17980 60
rect 17940 10 17980 40
rect 17940 -10 17950 10
rect 17970 -10 17980 10
rect 17940 -25 17980 -10
rect 18000 60 18040 75
rect 18000 40 18010 60
rect 18030 40 18040 60
rect 18000 10 18040 40
rect 18000 -10 18010 10
rect 18030 -10 18040 10
rect 18000 -25 18040 -10
rect 18060 60 18100 75
rect 18060 40 18070 60
rect 18090 40 18100 60
rect 18060 10 18100 40
rect 18060 -10 18070 10
rect 18090 -10 18100 10
rect 18060 -25 18100 -10
rect 18120 60 18160 75
rect 18120 40 18130 60
rect 18150 40 18160 60
rect 18120 10 18160 40
rect 18120 -10 18130 10
rect 18150 -10 18160 10
rect 18120 -25 18160 -10
rect 18180 60 18220 75
rect 18180 40 18190 60
rect 18210 40 18220 60
rect 18180 10 18220 40
rect 18180 -10 18190 10
rect 18210 -10 18220 10
rect 18180 -25 18220 -10
rect 18240 60 18280 75
rect 18240 40 18250 60
rect 18270 40 18280 60
rect 18240 10 18280 40
rect 18240 -10 18250 10
rect 18270 -10 18280 10
rect 18240 -25 18280 -10
rect 18300 60 18340 75
rect 18300 40 18310 60
rect 18330 40 18340 60
rect 18300 10 18340 40
rect 18300 -10 18310 10
rect 18330 -10 18340 10
rect 18300 -25 18340 -10
rect 18360 60 18400 75
rect 18360 40 18370 60
rect 18390 40 18400 60
rect 18360 10 18400 40
rect 18360 -10 18370 10
rect 18390 -10 18400 10
rect 18360 -25 18400 -10
rect 18420 60 18460 75
rect 18420 40 18430 60
rect 18450 40 18460 60
rect 18420 10 18460 40
rect 18420 -10 18430 10
rect 18450 -10 18460 10
rect 18420 -25 18460 -10
rect 18480 60 18520 75
rect 18480 40 18490 60
rect 18510 40 18520 60
rect 18480 10 18520 40
rect 18480 -10 18490 10
rect 18510 -10 18520 10
rect 18480 -25 18520 -10
rect 18540 60 18580 75
rect 18540 40 18550 60
rect 18570 40 18580 60
rect 18540 10 18580 40
rect 18540 -10 18550 10
rect 18570 -10 18580 10
rect 18540 -25 18580 -10
rect 18600 60 18640 75
rect 18600 40 18610 60
rect 18630 40 18640 60
rect 18600 10 18640 40
rect 18600 -10 18610 10
rect 18630 -10 18640 10
rect 18600 -25 18640 -10
rect 18660 60 18700 75
rect 18660 40 18670 60
rect 18690 40 18700 60
rect 18660 10 18700 40
rect 18660 -10 18670 10
rect 18690 -10 18700 10
rect 18660 -25 18700 -10
rect 18720 60 18760 75
rect 18720 40 18730 60
rect 18750 40 18760 60
rect 18720 10 18760 40
rect 18720 -10 18730 10
rect 18750 -10 18760 10
rect 18720 -25 18760 -10
rect 18780 60 18820 75
rect 18780 40 18790 60
rect 18810 40 18820 60
rect 18780 10 18820 40
rect 18780 -10 18790 10
rect 18810 -10 18820 10
rect 18780 -25 18820 -10
rect 18840 60 18880 75
rect 18840 40 18850 60
rect 18870 40 18880 60
rect 18840 10 18880 40
rect 18840 -10 18850 10
rect 18870 -10 18880 10
rect 18840 -25 18880 -10
rect 18900 60 18940 75
rect 18900 40 18910 60
rect 18930 40 18940 60
rect 18900 10 18940 40
rect 18900 -10 18910 10
rect 18930 -10 18940 10
rect 18900 -25 18940 -10
rect 18960 60 19000 75
rect 18960 40 18970 60
rect 18990 40 19000 60
rect 18960 10 19000 40
rect 18960 -10 18970 10
rect 18990 -10 19000 10
rect 18960 -25 19000 -10
rect 19020 60 19060 75
rect 19020 40 19030 60
rect 19050 40 19060 60
rect 19020 10 19060 40
rect 19020 -10 19030 10
rect 19050 -10 19060 10
rect 19020 -25 19060 -10
rect 19080 60 19120 75
rect 19080 40 19090 60
rect 19110 40 19120 60
rect 19080 10 19120 40
rect 19080 -10 19090 10
rect 19110 -10 19120 10
rect 19080 -25 19120 -10
rect 19140 60 19180 75
rect 19140 40 19150 60
rect 19170 40 19180 60
rect 19140 10 19180 40
rect 19140 -10 19150 10
rect 19170 -10 19180 10
rect 19140 -25 19180 -10
<< ndiffc >>
rect 16860 -335 16880 -315
rect 16920 -335 16940 -315
rect 16980 -335 17000 -315
rect 17040 -335 17060 -315
rect 17100 -335 17120 -315
rect 17160 -335 17180 -315
rect 17220 -335 17240 -315
rect 17280 -335 17300 -315
rect 17340 -335 17360 -315
rect 17400 -335 17420 -315
rect 17460 -335 17480 -315
rect 18120 -335 18140 -315
rect 18180 -335 18200 -315
rect 18240 -335 18260 -315
rect 18300 -335 18320 -315
rect 18360 -335 18380 -315
rect 18420 -335 18440 -315
rect 18480 -335 18500 -315
rect 18540 -335 18560 -315
rect 18600 -335 18620 -315
rect 18660 -335 18680 -315
rect 18720 -335 18740 -315
rect 16540 -610 16560 -590
rect 16540 -660 16560 -640
rect 16540 -710 16560 -690
rect 16540 -760 16560 -740
rect 16540 -810 16560 -790
rect 17080 -610 17100 -590
rect 17160 -610 17180 -590
rect 17080 -660 17100 -640
rect 17160 -660 17180 -640
rect 17080 -710 17100 -690
rect 17160 -710 17180 -690
rect 17080 -760 17100 -740
rect 17160 -760 17180 -740
rect 17080 -810 17100 -790
rect 17160 -810 17180 -790
rect 17700 -610 17720 -590
rect 17700 -660 17720 -640
rect 17700 -710 17720 -690
rect 17700 -760 17720 -740
rect 17700 -810 17720 -790
rect 17880 -610 17900 -590
rect 17880 -660 17900 -640
rect 17880 -710 17900 -690
rect 17880 -760 17900 -740
rect 17880 -810 17900 -790
rect 18420 -610 18440 -590
rect 18500 -610 18520 -590
rect 18420 -660 18440 -640
rect 18500 -660 18520 -640
rect 18420 -710 18440 -690
rect 18500 -710 18520 -690
rect 18420 -760 18440 -740
rect 18500 -760 18520 -740
rect 18420 -810 18440 -790
rect 18500 -810 18520 -790
rect 19040 -610 19060 -590
rect 19040 -660 19060 -640
rect 19040 -710 19060 -690
rect 19040 -760 19060 -740
rect 19040 -810 19060 -790
rect 16750 -1080 16770 -1060
rect 16750 -1130 16770 -1110
rect 17790 -1080 17810 -1060
rect 17790 -1130 17810 -1110
rect 18830 -1080 18850 -1060
rect 18830 -1130 18850 -1110
rect 16900 -1355 16920 -1335
rect 16900 -1405 16920 -1385
rect 16955 -1355 16975 -1335
rect 16955 -1405 16975 -1385
rect 17010 -1355 17030 -1335
rect 17010 -1405 17030 -1385
rect 17065 -1355 17085 -1335
rect 17065 -1405 17085 -1385
rect 17120 -1355 17140 -1335
rect 17120 -1405 17140 -1385
rect 17175 -1355 17195 -1335
rect 17175 -1405 17195 -1385
rect 17230 -1355 17250 -1335
rect 17230 -1405 17250 -1385
rect 17285 -1355 17305 -1335
rect 17285 -1405 17305 -1385
rect 17340 -1355 17360 -1335
rect 17340 -1405 17360 -1385
rect 17515 -1355 17535 -1335
rect 17515 -1405 17535 -1385
rect 17570 -1355 17590 -1335
rect 17570 -1405 17590 -1385
rect 17625 -1355 17645 -1335
rect 17625 -1405 17645 -1385
rect 17680 -1355 17700 -1335
rect 17680 -1405 17700 -1385
rect 17735 -1355 17755 -1335
rect 17735 -1405 17755 -1385
rect 17790 -1355 17810 -1335
rect 17790 -1405 17810 -1385
rect 17845 -1355 17865 -1335
rect 17845 -1405 17865 -1385
rect 17900 -1355 17920 -1335
rect 17900 -1405 17920 -1385
rect 17955 -1355 17975 -1335
rect 17955 -1405 17975 -1385
rect 18010 -1355 18030 -1335
rect 18010 -1405 18030 -1385
rect 18065 -1355 18085 -1335
rect 18065 -1405 18085 -1385
rect 18240 -1355 18260 -1335
rect 18240 -1405 18260 -1385
rect 18295 -1355 18315 -1335
rect 18295 -1405 18315 -1385
rect 18350 -1355 18370 -1335
rect 18350 -1405 18370 -1385
rect 18405 -1355 18425 -1335
rect 18405 -1405 18425 -1385
rect 18460 -1355 18480 -1335
rect 18460 -1405 18480 -1385
rect 18515 -1355 18535 -1335
rect 18515 -1405 18535 -1385
rect 18570 -1355 18590 -1335
rect 18570 -1405 18590 -1385
rect 18625 -1355 18645 -1335
rect 18625 -1405 18645 -1385
rect 18680 -1355 18700 -1335
rect 18680 -1405 18700 -1385
<< pdiffc >>
rect 16250 1143 16270 1215
rect 16305 1143 16325 1215
rect 16360 1143 16380 1215
rect 16415 1143 16435 1215
rect 16470 1143 16490 1215
rect 16820 1143 16840 1215
rect 16875 1143 16895 1215
rect 16930 1143 16950 1215
rect 16985 1143 17005 1215
rect 17040 1143 17060 1215
rect 17095 1143 17115 1215
rect 17150 1143 17170 1215
rect 17625 1195 17645 1215
rect 17625 1145 17645 1165
rect 17625 1095 17645 1115
rect 17625 1045 17645 1065
rect 17680 1195 17700 1215
rect 17680 1145 17700 1165
rect 17680 1095 17700 1115
rect 17680 1045 17700 1065
rect 17735 1195 17755 1215
rect 17735 1145 17755 1165
rect 17735 1095 17755 1115
rect 17735 1045 17755 1065
rect 17790 1195 17810 1215
rect 17790 1145 17810 1165
rect 17790 1095 17810 1115
rect 17790 1045 17810 1065
rect 17845 1195 17865 1215
rect 17845 1145 17865 1165
rect 17845 1095 17865 1115
rect 17845 1045 17865 1065
rect 17900 1195 17920 1215
rect 17900 1145 17920 1165
rect 17900 1095 17920 1115
rect 17900 1045 17920 1065
rect 17955 1195 17975 1215
rect 17955 1145 17975 1165
rect 18430 1145 18450 1215
rect 18485 1145 18505 1215
rect 18540 1145 18560 1215
rect 18595 1145 18615 1215
rect 18650 1145 18670 1215
rect 18705 1145 18725 1215
rect 18760 1145 18780 1215
rect 17955 1095 17975 1115
rect 17955 1045 17975 1065
rect 16980 730 17000 750
rect 16980 680 17000 700
rect 16445 630 16465 650
rect 16445 580 16465 600
rect 16500 630 16520 650
rect 16500 580 16520 600
rect 16555 630 16575 650
rect 16555 580 16575 600
rect 16610 630 16630 650
rect 16610 580 16630 600
rect 16665 630 16685 650
rect 16665 580 16685 600
rect 16980 630 17000 650
rect 16980 580 17000 600
rect 16980 530 17000 550
rect 16980 480 17000 500
rect 17070 730 17090 750
rect 17070 680 17090 700
rect 17070 630 17090 650
rect 17070 580 17090 600
rect 17070 530 17090 550
rect 17070 480 17090 500
rect 17160 730 17180 750
rect 17160 680 17180 700
rect 17160 630 17180 650
rect 17160 580 17180 600
rect 17160 530 17180 550
rect 17160 480 17180 500
rect 17250 730 17270 750
rect 17250 680 17270 700
rect 17250 630 17270 650
rect 17250 580 17270 600
rect 17250 530 17270 550
rect 17250 480 17270 500
rect 17340 730 17360 750
rect 17340 680 17360 700
rect 17340 630 17360 650
rect 17340 580 17360 600
rect 17340 530 17360 550
rect 17340 480 17360 500
rect 17430 730 17450 750
rect 17430 680 17450 700
rect 17430 630 17450 650
rect 17430 580 17450 600
rect 17430 530 17450 550
rect 17430 480 17450 500
rect 17520 730 17540 750
rect 17520 680 17540 700
rect 17520 630 17540 650
rect 17520 580 17540 600
rect 17520 530 17540 550
rect 17520 480 17540 500
rect 17610 730 17630 750
rect 17610 680 17630 700
rect 17610 630 17630 650
rect 17610 580 17630 600
rect 17610 530 17630 550
rect 17610 480 17630 500
rect 17700 730 17720 750
rect 17700 680 17720 700
rect 17700 630 17720 650
rect 17700 580 17720 600
rect 17700 530 17720 550
rect 17700 480 17720 500
rect 17790 730 17810 750
rect 17790 680 17810 700
rect 17790 630 17810 650
rect 17790 580 17810 600
rect 17790 530 17810 550
rect 17790 480 17810 500
rect 17880 730 17900 750
rect 17880 680 17900 700
rect 17880 630 17900 650
rect 17880 580 17900 600
rect 17880 530 17900 550
rect 17880 480 17900 500
rect 17970 730 17990 750
rect 17970 680 17990 700
rect 17970 630 17990 650
rect 17970 580 17990 600
rect 17970 530 17990 550
rect 17970 480 17990 500
rect 18060 730 18080 750
rect 18060 680 18080 700
rect 18060 630 18080 650
rect 18060 580 18080 600
rect 18060 530 18080 550
rect 18060 480 18080 500
rect 18150 730 18170 750
rect 18150 680 18170 700
rect 18150 630 18170 650
rect 18150 580 18170 600
rect 18150 530 18170 550
rect 18150 480 18170 500
rect 18240 730 18260 750
rect 18240 680 18260 700
rect 18240 630 18260 650
rect 18240 580 18260 600
rect 18240 530 18260 550
rect 18240 480 18260 500
rect 18330 730 18350 750
rect 18330 680 18350 700
rect 18330 630 18350 650
rect 18330 580 18350 600
rect 18330 530 18350 550
rect 18330 480 18350 500
rect 18420 730 18440 750
rect 18420 680 18440 700
rect 18420 630 18440 650
rect 18420 580 18440 600
rect 18420 530 18440 550
rect 18420 480 18440 500
rect 18510 730 18530 750
rect 18510 680 18530 700
rect 18510 630 18530 650
rect 18510 580 18530 600
rect 18510 530 18530 550
rect 18510 480 18530 500
rect 18600 730 18620 750
rect 18600 680 18620 700
rect 18600 630 18620 650
rect 18600 580 18620 600
rect 18600 530 18620 550
rect 18965 680 18985 700
rect 18965 630 18985 650
rect 18965 580 18985 600
rect 18965 530 18985 550
rect 19020 680 19040 700
rect 19020 630 19040 650
rect 19020 580 19040 600
rect 19020 530 19040 550
rect 19075 680 19095 700
rect 19075 630 19095 650
rect 19075 580 19095 600
rect 19075 530 19095 550
rect 19130 680 19150 700
rect 19130 630 19150 650
rect 19130 580 19150 600
rect 19130 530 19150 550
rect 18600 480 18620 500
rect 16430 40 16450 60
rect 16430 -10 16450 10
rect 16490 40 16510 60
rect 16490 -10 16510 10
rect 16550 40 16570 60
rect 16550 -10 16570 10
rect 16610 40 16630 60
rect 16610 -10 16630 10
rect 16670 40 16690 60
rect 16670 -10 16690 10
rect 16730 40 16750 60
rect 16730 -10 16750 10
rect 16790 40 16810 60
rect 16790 -10 16810 10
rect 16850 40 16870 60
rect 16850 -10 16870 10
rect 16910 40 16930 60
rect 16910 -10 16930 10
rect 16970 40 16990 60
rect 16970 -10 16990 10
rect 17030 40 17050 60
rect 17030 -10 17050 10
rect 17090 40 17110 60
rect 17090 -10 17110 10
rect 17150 40 17170 60
rect 17150 -10 17170 10
rect 17210 40 17230 60
rect 17210 -10 17230 10
rect 17270 40 17290 60
rect 17270 -10 17290 10
rect 17330 40 17350 60
rect 17330 -10 17350 10
rect 17390 40 17410 60
rect 17390 -10 17410 10
rect 17450 40 17470 60
rect 17450 -10 17470 10
rect 17510 40 17530 60
rect 17510 -10 17530 10
rect 17570 40 17590 60
rect 17570 -10 17590 10
rect 17630 40 17650 60
rect 17630 -10 17650 10
rect 17950 40 17970 60
rect 17950 -10 17970 10
rect 18010 40 18030 60
rect 18010 -10 18030 10
rect 18070 40 18090 60
rect 18070 -10 18090 10
rect 18130 40 18150 60
rect 18130 -10 18150 10
rect 18190 40 18210 60
rect 18190 -10 18210 10
rect 18250 40 18270 60
rect 18250 -10 18270 10
rect 18310 40 18330 60
rect 18310 -10 18330 10
rect 18370 40 18390 60
rect 18370 -10 18390 10
rect 18430 40 18450 60
rect 18430 -10 18450 10
rect 18490 40 18510 60
rect 18490 -10 18510 10
rect 18550 40 18570 60
rect 18550 -10 18570 10
rect 18610 40 18630 60
rect 18610 -10 18630 10
rect 18670 40 18690 60
rect 18670 -10 18690 10
rect 18730 40 18750 60
rect 18730 -10 18750 10
rect 18790 40 18810 60
rect 18790 -10 18810 10
rect 18850 40 18870 60
rect 18850 -10 18870 10
rect 18910 40 18930 60
rect 18910 -10 18930 10
rect 18970 40 18990 60
rect 18970 -10 18990 10
rect 19030 40 19050 60
rect 19030 -10 19050 10
rect 19090 40 19110 60
rect 19090 -10 19110 10
rect 19150 40 19170 60
rect 19150 -10 19170 10
<< psubdiff >>
rect 17560 -315 17600 -300
rect 17560 -335 17570 -315
rect 17590 -335 17600 -315
rect 17560 -350 17600 -335
rect 18000 -315 18040 -300
rect 18000 -335 18010 -315
rect 18030 -335 18040 -315
rect 18000 -350 18040 -335
rect 17110 -590 17150 -575
rect 17110 -610 17120 -590
rect 17140 -610 17150 -590
rect 17110 -640 17150 -610
rect 17110 -660 17120 -640
rect 17140 -660 17150 -640
rect 17110 -690 17150 -660
rect 17110 -710 17120 -690
rect 17140 -710 17150 -690
rect 17110 -740 17150 -710
rect 17110 -760 17120 -740
rect 17140 -760 17150 -740
rect 17110 -790 17150 -760
rect 17110 -810 17120 -790
rect 17140 -810 17150 -790
rect 17110 -820 17150 -810
rect 18450 -590 18490 -575
rect 18450 -610 18460 -590
rect 18480 -610 18490 -590
rect 18450 -640 18490 -610
rect 18450 -660 18460 -640
rect 18480 -660 18490 -640
rect 18450 -690 18490 -660
rect 18450 -710 18460 -690
rect 18480 -710 18490 -690
rect 18450 -740 18490 -710
rect 18450 -760 18460 -740
rect 18480 -760 18490 -740
rect 18450 -790 18490 -760
rect 18450 -810 18460 -790
rect 18480 -810 18490 -790
rect 18450 -825 18490 -810
rect 18860 -1060 18900 -1045
rect 18860 -1080 18870 -1060
rect 18890 -1080 18900 -1060
rect 18860 -1110 18900 -1080
rect 18860 -1130 18870 -1110
rect 18890 -1130 18900 -1110
rect 18860 -1145 18900 -1130
rect 16850 -1335 16890 -1320
rect 16850 -1355 16860 -1335
rect 16880 -1355 16890 -1335
rect 16850 -1385 16890 -1355
rect 16850 -1405 16860 -1385
rect 16880 -1405 16890 -1385
rect 16850 -1420 16890 -1405
rect 17370 -1335 17410 -1320
rect 17370 -1355 17380 -1335
rect 17400 -1355 17410 -1335
rect 17370 -1385 17410 -1355
rect 17370 -1405 17380 -1385
rect 17400 -1405 17410 -1385
rect 17370 -1420 17410 -1405
rect 17465 -1335 17505 -1320
rect 17465 -1355 17475 -1335
rect 17495 -1355 17505 -1335
rect 17465 -1385 17505 -1355
rect 17465 -1405 17475 -1385
rect 17495 -1405 17505 -1385
rect 17465 -1420 17505 -1405
rect 18095 -1335 18135 -1320
rect 18095 -1355 18105 -1335
rect 18125 -1355 18135 -1335
rect 18095 -1385 18135 -1355
rect 18095 -1405 18105 -1385
rect 18125 -1405 18135 -1385
rect 18095 -1420 18135 -1405
rect 18190 -1335 18230 -1320
rect 18190 -1355 18200 -1335
rect 18220 -1355 18230 -1335
rect 18190 -1385 18230 -1355
rect 18190 -1405 18200 -1385
rect 18220 -1405 18230 -1385
rect 18190 -1420 18230 -1405
rect 18710 -1335 18750 -1320
rect 18710 -1355 18720 -1335
rect 18740 -1355 18750 -1335
rect 18710 -1385 18750 -1355
rect 18710 -1405 18720 -1385
rect 18740 -1405 18750 -1385
rect 18710 -1420 18750 -1405
rect 17775 -4170 17825 -4155
rect 17775 -4190 17790 -4170
rect 17810 -4190 17825 -4170
rect 17775 -4220 17825 -4190
rect 17775 -4240 17790 -4220
rect 17810 -4240 17825 -4220
rect 17775 -4270 17825 -4240
rect 17775 -4290 17790 -4270
rect 17810 -4290 17825 -4270
rect 17775 -4305 17825 -4290
<< nsubdiff >>
rect 16200 1217 16240 1230
rect 16200 1145 16210 1217
rect 16230 1145 16240 1217
rect 16200 1130 16240 1145
rect 16500 1217 16540 1230
rect 16500 1145 16510 1217
rect 16530 1145 16540 1217
rect 16500 1130 16540 1145
rect 16770 1217 16810 1230
rect 16770 1145 16780 1217
rect 16800 1145 16810 1217
rect 16770 1130 16810 1145
rect 17180 1217 17220 1230
rect 17180 1145 17190 1217
rect 17210 1145 17220 1217
rect 17180 1130 17220 1145
rect 17575 1215 17615 1230
rect 17575 1195 17585 1215
rect 17605 1195 17615 1215
rect 17575 1165 17615 1195
rect 17575 1145 17585 1165
rect 17605 1145 17615 1165
rect 17575 1115 17615 1145
rect 17575 1095 17585 1115
rect 17605 1095 17615 1115
rect 17575 1065 17615 1095
rect 17575 1045 17585 1065
rect 17605 1045 17615 1065
rect 17575 1030 17615 1045
rect 17985 1215 18025 1230
rect 17985 1195 17995 1215
rect 18015 1195 18025 1215
rect 17985 1165 18025 1195
rect 17985 1145 17995 1165
rect 18015 1145 18025 1165
rect 17985 1115 18025 1145
rect 18380 1217 18420 1230
rect 18380 1145 18390 1217
rect 18410 1145 18420 1217
rect 18380 1130 18420 1145
rect 18790 1217 18830 1230
rect 18790 1145 18800 1217
rect 18820 1145 18830 1217
rect 18790 1130 18830 1145
rect 17985 1095 17995 1115
rect 18015 1095 18025 1115
rect 17985 1065 18025 1095
rect 17985 1045 17995 1065
rect 18015 1045 18025 1065
rect 17985 1030 18025 1045
rect 16930 750 16970 765
rect 16930 730 16940 750
rect 16960 730 16970 750
rect 16930 700 16970 730
rect 16930 680 16940 700
rect 16960 680 16970 700
rect 16395 650 16435 665
rect 16395 630 16405 650
rect 16425 630 16435 650
rect 16395 600 16435 630
rect 16395 580 16405 600
rect 16425 580 16435 600
rect 16395 565 16435 580
rect 16700 650 16740 665
rect 16700 630 16710 650
rect 16730 630 16740 650
rect 16700 600 16740 630
rect 16700 580 16710 600
rect 16730 580 16740 600
rect 16700 565 16740 580
rect 16930 650 16970 680
rect 16930 630 16940 650
rect 16960 630 16970 650
rect 16930 600 16970 630
rect 16930 580 16940 600
rect 16960 580 16970 600
rect 16930 550 16970 580
rect 16930 530 16940 550
rect 16960 530 16970 550
rect 16930 500 16970 530
rect 16930 480 16940 500
rect 16960 480 16970 500
rect 16930 465 16970 480
rect 18630 750 18670 765
rect 18630 730 18640 750
rect 18660 730 18670 750
rect 18630 700 18670 730
rect 18630 680 18640 700
rect 18660 680 18670 700
rect 18630 650 18670 680
rect 18630 630 18640 650
rect 18660 630 18670 650
rect 18630 600 18670 630
rect 18630 580 18640 600
rect 18660 580 18670 600
rect 18630 550 18670 580
rect 18630 530 18640 550
rect 18660 530 18670 550
rect 18630 500 18670 530
rect 18915 700 18955 715
rect 18915 680 18925 700
rect 18945 680 18955 700
rect 18915 650 18955 680
rect 18915 630 18925 650
rect 18945 630 18955 650
rect 18915 600 18955 630
rect 18915 580 18925 600
rect 18945 580 18955 600
rect 18915 550 18955 580
rect 18915 530 18925 550
rect 18945 530 18955 550
rect 18915 515 18955 530
rect 19160 700 19200 715
rect 19160 680 19170 700
rect 19190 680 19200 700
rect 19160 650 19200 680
rect 19160 630 19170 650
rect 19190 630 19200 650
rect 19160 600 19200 630
rect 19160 580 19170 600
rect 19190 580 19200 600
rect 19160 550 19200 580
rect 19160 530 19170 550
rect 19190 530 19200 550
rect 19160 515 19200 530
rect 18630 480 18640 500
rect 18660 480 18670 500
rect 18630 465 18670 480
rect 16380 60 16420 75
rect 16380 40 16390 60
rect 16410 40 16420 60
rect 16380 10 16420 40
rect 16380 -10 16390 10
rect 16410 -10 16420 10
rect 16380 -25 16420 -10
rect 17660 60 17700 75
rect 17660 40 17670 60
rect 17690 40 17700 60
rect 17660 10 17700 40
rect 17660 -10 17670 10
rect 17690 -10 17700 10
rect 17660 -25 17700 -10
rect 17900 60 17940 75
rect 17900 40 17910 60
rect 17930 40 17940 60
rect 17900 10 17940 40
rect 17900 -10 17910 10
rect 17930 -10 17940 10
rect 17900 -25 17940 -10
rect 19180 60 19220 75
rect 19180 40 19190 60
rect 19210 40 19220 60
rect 19180 10 19220 40
rect 19180 -10 19190 10
rect 19210 -10 19220 10
rect 19180 -25 19220 -10
<< psubdiffcont >>
rect 17570 -335 17590 -315
rect 18010 -335 18030 -315
rect 17120 -610 17140 -590
rect 17120 -660 17140 -640
rect 17120 -710 17140 -690
rect 17120 -760 17140 -740
rect 17120 -810 17140 -790
rect 18460 -610 18480 -590
rect 18460 -660 18480 -640
rect 18460 -710 18480 -690
rect 18460 -760 18480 -740
rect 18460 -810 18480 -790
rect 18870 -1080 18890 -1060
rect 18870 -1130 18890 -1110
rect 16860 -1355 16880 -1335
rect 16860 -1405 16880 -1385
rect 17380 -1355 17400 -1335
rect 17380 -1405 17400 -1385
rect 17475 -1355 17495 -1335
rect 17475 -1405 17495 -1385
rect 18105 -1355 18125 -1335
rect 18105 -1405 18125 -1385
rect 18200 -1355 18220 -1335
rect 18200 -1405 18220 -1385
rect 18720 -1355 18740 -1335
rect 18720 -1405 18740 -1385
rect 17790 -4190 17810 -4170
rect 17790 -4240 17810 -4220
rect 17790 -4290 17810 -4270
<< nsubdiffcont >>
rect 16210 1145 16230 1217
rect 16510 1145 16530 1217
rect 16780 1145 16800 1217
rect 17190 1145 17210 1217
rect 17585 1195 17605 1215
rect 17585 1145 17605 1165
rect 17585 1095 17605 1115
rect 17585 1045 17605 1065
rect 17995 1195 18015 1215
rect 17995 1145 18015 1165
rect 18390 1145 18410 1217
rect 18800 1145 18820 1217
rect 17995 1095 18015 1115
rect 17995 1045 18015 1065
rect 16940 730 16960 750
rect 16940 680 16960 700
rect 16405 630 16425 650
rect 16405 580 16425 600
rect 16710 630 16730 650
rect 16710 580 16730 600
rect 16940 630 16960 650
rect 16940 580 16960 600
rect 16940 530 16960 550
rect 16940 480 16960 500
rect 18640 730 18660 750
rect 18640 680 18660 700
rect 18640 630 18660 650
rect 18640 580 18660 600
rect 18640 530 18660 550
rect 18925 680 18945 700
rect 18925 630 18945 650
rect 18925 580 18945 600
rect 18925 530 18945 550
rect 19170 680 19190 700
rect 19170 630 19190 650
rect 19170 580 19190 600
rect 19170 530 19190 550
rect 18640 480 18660 500
rect 16390 40 16410 60
rect 16390 -10 16410 10
rect 17670 40 17690 60
rect 17670 -10 17690 10
rect 17910 40 17930 60
rect 17910 -10 17930 10
rect 19190 40 19210 60
rect 19190 -10 19210 10
<< poly >>
rect 16240 1275 16280 1285
rect 16240 1255 16250 1275
rect 16270 1260 16280 1275
rect 16394 1275 16424 1285
rect 16394 1260 16399 1275
rect 16270 1255 16295 1260
rect 16240 1245 16295 1255
rect 16280 1230 16295 1245
rect 16335 1255 16399 1260
rect 16419 1255 16424 1275
rect 16460 1275 16500 1285
rect 16460 1260 16470 1275
rect 16335 1245 16424 1255
rect 16445 1255 16470 1260
rect 16490 1255 16500 1275
rect 16445 1245 16500 1255
rect 16810 1275 16850 1285
rect 16810 1255 16820 1275
rect 16840 1260 16850 1275
rect 16980 1275 17010 1285
rect 16840 1255 16865 1260
rect 16980 1255 16985 1275
rect 17005 1255 17010 1275
rect 17140 1275 17180 1285
rect 17140 1255 17150 1275
rect 17170 1255 17180 1275
rect 16810 1245 16865 1255
rect 16335 1240 16405 1245
rect 16335 1230 16350 1240
rect 16390 1230 16405 1240
rect 16445 1230 16460 1245
rect 16850 1230 16865 1245
rect 16905 1240 17085 1255
rect 16905 1230 16920 1240
rect 16960 1230 16975 1240
rect 17015 1230 17030 1240
rect 17070 1230 17085 1240
rect 17125 1240 17180 1255
rect 17605 1275 17645 1285
rect 17605 1255 17615 1275
rect 17635 1260 17645 1275
rect 17840 1275 17870 1285
rect 17635 1255 17670 1260
rect 17840 1255 17845 1275
rect 17865 1255 17870 1275
rect 17955 1275 17995 1285
rect 17955 1260 17965 1275
rect 17930 1255 17965 1260
rect 17985 1255 17995 1275
rect 17605 1245 17670 1255
rect 17125 1230 17140 1240
rect 17655 1230 17670 1245
rect 17710 1240 17890 1255
rect 17710 1230 17725 1240
rect 17765 1230 17780 1240
rect 17820 1230 17835 1240
rect 17875 1230 17890 1240
rect 17930 1245 17995 1255
rect 18420 1275 18460 1285
rect 18420 1255 18430 1275
rect 18450 1260 18460 1275
rect 18590 1275 18620 1285
rect 18450 1255 18475 1260
rect 18590 1255 18595 1275
rect 18615 1255 18620 1275
rect 18750 1275 18790 1285
rect 18750 1260 18760 1275
rect 18735 1255 18760 1260
rect 18780 1255 18790 1275
rect 18420 1245 18475 1255
rect 17930 1230 17945 1245
rect 18460 1230 18475 1245
rect 18515 1240 18695 1255
rect 18515 1230 18530 1240
rect 18570 1230 18585 1240
rect 18625 1230 18640 1240
rect 18680 1230 18695 1240
rect 18735 1245 18790 1255
rect 18735 1230 18750 1245
rect 16280 1115 16295 1130
rect 16335 1115 16350 1130
rect 16390 1115 16405 1130
rect 16445 1115 16460 1130
rect 16850 1115 16865 1130
rect 16905 1115 16920 1130
rect 16960 1115 16975 1130
rect 17015 1115 17030 1130
rect 17070 1115 17085 1130
rect 17125 1115 17140 1130
rect 18460 1115 18475 1130
rect 18515 1115 18530 1130
rect 18570 1115 18585 1130
rect 18625 1115 18640 1130
rect 18680 1115 18695 1130
rect 18735 1115 18750 1130
rect 17655 1015 17670 1030
rect 17710 1015 17725 1030
rect 17765 1015 17780 1030
rect 17820 1015 17835 1030
rect 17875 1015 17890 1030
rect 17930 1015 17945 1030
rect 16970 810 17010 820
rect 16970 790 16980 810
rect 17000 795 17010 810
rect 18590 810 18630 820
rect 18590 795 18600 810
rect 17000 790 17060 795
rect 16970 780 17060 790
rect 18540 790 18600 795
rect 18620 790 18630 810
rect 18540 780 18630 790
rect 17010 765 17060 780
rect 17100 765 17150 780
rect 17190 765 17240 780
rect 17280 765 17330 780
rect 17370 765 17420 780
rect 17460 765 17510 780
rect 17550 765 17600 780
rect 17640 765 17690 780
rect 17730 765 17780 780
rect 17820 765 17870 780
rect 17910 765 17960 780
rect 18000 765 18050 780
rect 18090 765 18140 780
rect 18180 765 18230 780
rect 18270 765 18320 780
rect 18360 765 18410 780
rect 18450 765 18500 780
rect 18540 765 18590 780
rect 16440 710 16470 720
rect 16440 690 16445 710
rect 16465 690 16470 710
rect 16660 710 16690 720
rect 16660 690 16665 710
rect 16685 690 16690 710
rect 16440 675 16490 690
rect 16475 665 16490 675
rect 16530 665 16545 680
rect 16585 665 16600 680
rect 16640 675 16690 690
rect 16640 665 16655 675
rect 16475 550 16490 565
rect 16530 555 16545 565
rect 16585 555 16600 565
rect 16530 540 16600 555
rect 16640 550 16655 565
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 18950 760 18980 770
rect 18950 740 18955 760
rect 18975 745 18980 760
rect 19125 760 19155 770
rect 19125 745 19130 760
rect 18975 740 19010 745
rect 18950 730 19010 740
rect 19105 740 19130 745
rect 19150 740 19155 760
rect 19105 730 19155 740
rect 18995 715 19010 730
rect 19050 715 19065 730
rect 19105 715 19120 730
rect 18995 500 19010 515
rect 19050 500 19065 515
rect 19105 500 19120 515
rect 19031 490 19065 500
rect 19031 470 19036 490
rect 19056 480 19065 490
rect 19056 470 19061 480
rect 17010 450 17060 465
rect 17100 455 17150 465
rect 17190 455 17240 465
rect 17280 455 17330 465
rect 17370 455 17420 465
rect 17460 455 17510 465
rect 17550 455 17600 465
rect 17640 455 17690 465
rect 17730 455 17780 465
rect 17820 455 17870 465
rect 17910 455 17960 465
rect 18000 455 18050 465
rect 18090 455 18140 465
rect 18180 455 18230 465
rect 18270 455 18320 465
rect 18360 455 18410 465
rect 18450 455 18500 465
rect 17100 440 18500 455
rect 18540 450 18590 465
rect 19031 460 19061 470
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 16425 120 16455 130
rect 16425 100 16430 120
rect 16450 100 16455 120
rect 17625 120 17655 130
rect 17625 100 17630 120
rect 17650 100 17655 120
rect 16425 85 16480 100
rect 16460 75 16480 85
rect 16520 75 16540 90
rect 16580 75 16600 90
rect 16640 75 16660 90
rect 16700 75 16720 90
rect 16760 75 16780 90
rect 16820 75 16840 90
rect 16880 75 16900 90
rect 16940 75 16960 90
rect 17000 75 17020 90
rect 17060 75 17080 90
rect 17120 75 17140 90
rect 17180 75 17200 90
rect 17240 75 17260 90
rect 17300 75 17320 90
rect 17360 75 17380 90
rect 17420 75 17440 90
rect 17480 75 17500 90
rect 17540 75 17560 90
rect 17600 85 17655 100
rect 17945 120 17975 130
rect 17945 100 17950 120
rect 17970 100 17975 120
rect 19145 120 19175 130
rect 19145 100 19150 120
rect 19170 100 19175 120
rect 17945 85 18000 100
rect 17600 75 17620 85
rect 17980 75 18000 85
rect 18040 75 18060 90
rect 18100 75 18120 90
rect 18160 75 18180 90
rect 18220 75 18240 90
rect 18280 75 18300 90
rect 18340 75 18360 90
rect 18400 75 18420 90
rect 18460 75 18480 90
rect 18520 75 18540 90
rect 18580 75 18600 90
rect 18640 75 18660 90
rect 18700 75 18720 90
rect 18760 75 18780 90
rect 18820 75 18840 90
rect 18880 75 18900 90
rect 18940 75 18960 90
rect 19000 75 19020 90
rect 19060 75 19080 90
rect 19120 85 19175 100
rect 19120 75 19140 85
rect 16460 -35 16480 -25
rect 16425 -50 16480 -35
rect 16520 -40 16540 -25
rect 16580 -35 16600 -25
rect 16640 -35 16660 -25
rect 16700 -35 16720 -25
rect 16760 -35 16780 -25
rect 16510 -50 16550 -40
rect 16580 -50 16780 -35
rect 16820 -35 16840 -25
rect 16880 -35 16900 -25
rect 16820 -50 16900 -35
rect 16940 -35 16960 -25
rect 17000 -35 17020 -25
rect 17060 -35 17080 -25
rect 17120 -35 17140 -25
rect 16940 -50 17140 -35
rect 17180 -35 17200 -25
rect 17240 -35 17260 -25
rect 17180 -50 17260 -35
rect 17300 -35 17320 -25
rect 17360 -35 17380 -25
rect 17420 -35 17440 -25
rect 17480 -35 17500 -25
rect 17300 -50 17500 -35
rect 17540 -40 17560 -25
rect 17600 -40 17620 -25
rect 17980 -35 18000 -25
rect 17535 -50 17565 -40
rect 16425 -70 16430 -50
rect 16450 -70 16455 -50
rect 16425 -80 16455 -70
rect 16510 -70 16520 -50
rect 16540 -70 16550 -50
rect 16510 -80 16550 -70
rect 16600 -70 16610 -50
rect 16630 -70 16640 -50
rect 16600 -80 16640 -70
rect 16840 -70 16850 -50
rect 16870 -70 16880 -50
rect 16840 -80 16880 -70
rect 16960 -70 16970 -50
rect 16990 -70 17000 -50
rect 16960 -80 17000 -70
rect 17200 -70 17210 -50
rect 17230 -70 17240 -50
rect 17200 -80 17240 -70
rect 17320 -70 17330 -50
rect 17350 -70 17360 -50
rect 17320 -80 17360 -70
rect 17535 -70 17540 -50
rect 17560 -70 17565 -50
rect 17535 -80 17565 -70
rect 17945 -50 18000 -35
rect 18040 -40 18060 -25
rect 18100 -35 18120 -25
rect 18160 -35 18180 -25
rect 18220 -35 18240 -25
rect 18280 -35 18300 -25
rect 18035 -50 18065 -40
rect 18100 -50 18300 -35
rect 18340 -35 18360 -25
rect 18400 -35 18420 -25
rect 18340 -50 18420 -35
rect 18460 -35 18480 -25
rect 18520 -35 18540 -25
rect 18580 -35 18600 -25
rect 18640 -35 18660 -25
rect 18460 -50 18660 -35
rect 18700 -35 18720 -25
rect 18760 -35 18780 -25
rect 18700 -50 18780 -35
rect 18820 -35 18840 -25
rect 18880 -35 18900 -25
rect 18940 -35 18960 -25
rect 19000 -35 19020 -25
rect 18820 -50 19020 -35
rect 19060 -40 19080 -25
rect 19120 -35 19140 -25
rect 19050 -50 19090 -40
rect 19120 -50 19175 -35
rect 17945 -70 17950 -50
rect 17970 -70 17975 -50
rect 17945 -80 17975 -70
rect 18035 -70 18040 -50
rect 18060 -70 18065 -50
rect 18035 -80 18065 -70
rect 18240 -70 18250 -50
rect 18270 -70 18280 -50
rect 18240 -80 18280 -70
rect 18360 -70 18370 -50
rect 18390 -70 18400 -50
rect 18360 -80 18400 -70
rect 18600 -70 18610 -50
rect 18630 -70 18640 -50
rect 18600 -80 18640 -70
rect 18720 -70 18730 -50
rect 18750 -70 18760 -50
rect 18720 -80 18760 -70
rect 18960 -70 18970 -50
rect 18990 -70 19000 -50
rect 18960 -80 19000 -70
rect 19050 -70 19060 -50
rect 19080 -70 19090 -50
rect 19050 -80 19090 -70
rect 19145 -70 19150 -50
rect 19170 -70 19175 -50
rect 19145 -80 19175 -70
rect 16910 -210 16950 -200
rect 16910 -230 16920 -210
rect 16940 -230 16950 -210
rect 16910 -245 16950 -230
rect 18650 -210 18690 -200
rect 18650 -230 18660 -210
rect 18680 -230 18690 -210
rect 18650 -245 18690 -230
rect 16910 -260 17450 -245
rect 16890 -300 16910 -285
rect 16950 -300 16970 -260
rect 17010 -300 17030 -260
rect 17070 -300 17090 -285
rect 17130 -300 17150 -285
rect 17190 -300 17210 -260
rect 17250 -300 17270 -260
rect 17310 -300 17330 -285
rect 17370 -300 17390 -285
rect 17430 -300 17450 -260
rect 18150 -260 18690 -245
rect 18150 -300 18170 -260
rect 18210 -300 18230 -285
rect 18270 -300 18290 -285
rect 18330 -300 18350 -260
rect 18390 -300 18410 -260
rect 18450 -300 18470 -285
rect 18510 -300 18530 -285
rect 18570 -300 18590 -260
rect 18630 -300 18650 -260
rect 18690 -300 18710 -285
rect 16890 -365 16910 -350
rect 16950 -365 16970 -350
rect 17010 -365 17030 -350
rect 16850 -375 16910 -365
rect 16850 -395 16860 -375
rect 16880 -390 16910 -375
rect 17070 -390 17090 -350
rect 17130 -390 17150 -350
rect 17190 -365 17210 -350
rect 17250 -365 17270 -350
rect 17310 -390 17330 -350
rect 17370 -390 17390 -350
rect 17430 -365 17450 -350
rect 18150 -365 18170 -350
rect 16880 -395 17390 -390
rect 16850 -405 17390 -395
rect 18210 -390 18230 -350
rect 18270 -390 18290 -350
rect 18330 -365 18350 -350
rect 18390 -365 18410 -350
rect 18450 -390 18470 -350
rect 18510 -390 18530 -350
rect 18570 -365 18590 -350
rect 18630 -365 18650 -350
rect 18690 -365 18710 -350
rect 18690 -375 18750 -365
rect 18690 -390 18720 -375
rect 18210 -395 18720 -390
rect 18740 -395 18750 -375
rect 18210 -405 18750 -395
rect 16620 -535 16660 -525
rect 16620 -555 16630 -535
rect 16650 -555 16660 -535
rect 16620 -560 16660 -555
rect 16740 -535 16780 -525
rect 16740 -555 16750 -535
rect 16770 -555 16780 -535
rect 16740 -560 16780 -555
rect 16860 -535 16900 -525
rect 16860 -555 16870 -535
rect 16890 -555 16900 -535
rect 16860 -560 16900 -555
rect 16980 -535 17020 -525
rect 16980 -555 16990 -535
rect 17010 -555 17020 -535
rect 16980 -560 17020 -555
rect 17300 -535 17340 -525
rect 17300 -555 17310 -535
rect 17330 -555 17340 -535
rect 17300 -560 17340 -555
rect 17420 -535 17460 -525
rect 17420 -555 17430 -535
rect 17450 -555 17460 -535
rect 17420 -560 17460 -555
rect 17540 -535 17580 -525
rect 17540 -555 17550 -535
rect 17570 -555 17580 -535
rect 17540 -560 17580 -555
rect 18020 -535 18060 -525
rect 18020 -555 18030 -535
rect 18050 -555 18060 -535
rect 18020 -560 18060 -555
rect 18140 -535 18180 -525
rect 18140 -555 18150 -535
rect 18170 -555 18180 -535
rect 18140 -560 18180 -555
rect 18260 -535 18300 -525
rect 18260 -555 18270 -535
rect 18290 -555 18300 -535
rect 18260 -560 18300 -555
rect 18580 -535 18620 -525
rect 18580 -555 18590 -535
rect 18610 -555 18620 -535
rect 18580 -560 18620 -555
rect 18700 -535 18740 -525
rect 18700 -555 18710 -535
rect 18730 -555 18740 -535
rect 18700 -560 18740 -555
rect 18820 -535 18860 -525
rect 18820 -555 18830 -535
rect 18850 -555 18860 -535
rect 18820 -560 18860 -555
rect 18940 -535 18980 -525
rect 18940 -555 18950 -535
rect 18970 -555 18980 -535
rect 18940 -560 18980 -555
rect 16570 -575 17070 -560
rect 17190 -575 17690 -560
rect 17910 -575 18410 -560
rect 18530 -575 19030 -560
rect 16570 -840 17070 -825
rect 17190 -840 17690 -825
rect 17910 -840 18410 -825
rect 18530 -840 19030 -825
rect 16820 -1000 16860 -990
rect 16820 -1020 16830 -1000
rect 16850 -1020 16860 -1000
rect 16820 -1030 16860 -1020
rect 16900 -1000 16940 -990
rect 16900 -1020 16910 -1000
rect 16930 -1020 16940 -1000
rect 16900 -1030 16940 -1020
rect 16980 -1000 17020 -990
rect 16980 -1020 16990 -1000
rect 17010 -1020 17020 -1000
rect 16980 -1030 17020 -1020
rect 17060 -1000 17100 -990
rect 17060 -1020 17070 -1000
rect 17090 -1020 17100 -1000
rect 17060 -1030 17100 -1020
rect 17140 -1000 17180 -990
rect 17140 -1020 17150 -1000
rect 17170 -1020 17180 -1000
rect 17140 -1030 17180 -1020
rect 17220 -1000 17260 -990
rect 17220 -1020 17230 -1000
rect 17250 -1020 17260 -1000
rect 17220 -1030 17260 -1020
rect 17300 -1000 17340 -990
rect 17300 -1020 17310 -1000
rect 17330 -1020 17340 -1000
rect 17300 -1030 17340 -1020
rect 17380 -1000 17420 -990
rect 17380 -1020 17390 -1000
rect 17410 -1020 17420 -1000
rect 17380 -1030 17420 -1020
rect 17460 -1000 17500 -990
rect 17460 -1020 17470 -1000
rect 17490 -1020 17500 -1000
rect 17460 -1030 17500 -1020
rect 17540 -1000 17580 -990
rect 17540 -1020 17550 -1000
rect 17570 -1020 17580 -1000
rect 17540 -1030 17580 -1020
rect 17620 -1000 17660 -990
rect 17620 -1020 17630 -1000
rect 17650 -1020 17660 -1000
rect 17620 -1030 17660 -1020
rect 17700 -1000 17740 -990
rect 17700 -1020 17710 -1000
rect 17730 -1020 17740 -1000
rect 17700 -1030 17740 -1020
rect 17860 -1000 17900 -990
rect 17860 -1020 17870 -1000
rect 17890 -1020 17900 -1000
rect 17860 -1030 17900 -1020
rect 17940 -1000 17980 -990
rect 17940 -1020 17950 -1000
rect 17970 -1020 17980 -1000
rect 17940 -1030 17980 -1020
rect 18020 -1000 18060 -990
rect 18020 -1020 18030 -1000
rect 18050 -1020 18060 -1000
rect 18020 -1030 18060 -1020
rect 18100 -1000 18140 -990
rect 18100 -1020 18110 -1000
rect 18130 -1020 18140 -1000
rect 18100 -1030 18140 -1020
rect 18180 -1000 18220 -990
rect 18180 -1020 18190 -1000
rect 18210 -1020 18220 -1000
rect 18180 -1030 18220 -1020
rect 18260 -1000 18300 -990
rect 18260 -1020 18270 -1000
rect 18290 -1020 18300 -1000
rect 18260 -1030 18300 -1020
rect 18340 -1000 18380 -990
rect 18340 -1020 18350 -1000
rect 18370 -1020 18380 -1000
rect 18340 -1030 18380 -1020
rect 18420 -1000 18460 -990
rect 18420 -1020 18430 -1000
rect 18450 -1020 18460 -1000
rect 18420 -1030 18460 -1020
rect 18500 -1000 18540 -990
rect 18500 -1020 18510 -1000
rect 18530 -1020 18540 -1000
rect 18500 -1030 18540 -1020
rect 18580 -1000 18620 -990
rect 18580 -1020 18590 -1000
rect 18610 -1020 18620 -1000
rect 18580 -1030 18620 -1020
rect 18660 -1000 18700 -990
rect 18660 -1020 18670 -1000
rect 18690 -1020 18700 -1000
rect 18660 -1030 18700 -1020
rect 18740 -1000 18780 -990
rect 18740 -1020 18750 -1000
rect 18770 -1020 18780 -1000
rect 18740 -1030 18780 -1020
rect 16780 -1045 17780 -1030
rect 17820 -1045 18820 -1030
rect 16780 -1160 17780 -1145
rect 17820 -1160 18820 -1145
rect 16890 -1275 16930 -1265
rect 16890 -1295 16900 -1275
rect 16920 -1290 16930 -1275
rect 17170 -1275 17200 -1265
rect 16920 -1295 16945 -1290
rect 17170 -1295 17175 -1275
rect 17195 -1295 17200 -1275
rect 17330 -1275 17370 -1265
rect 17330 -1290 17340 -1275
rect 17315 -1295 17340 -1290
rect 17360 -1295 17370 -1275
rect 16890 -1305 16945 -1295
rect 16930 -1320 16945 -1305
rect 16985 -1310 17275 -1295
rect 16985 -1320 17000 -1310
rect 17040 -1320 17055 -1310
rect 17095 -1320 17110 -1310
rect 17150 -1320 17165 -1310
rect 17205 -1320 17220 -1310
rect 17260 -1320 17275 -1310
rect 17315 -1305 17370 -1295
rect 17505 -1275 17545 -1265
rect 17505 -1295 17515 -1275
rect 17535 -1290 17545 -1275
rect 17785 -1275 17815 -1265
rect 17535 -1295 17560 -1290
rect 17785 -1295 17790 -1275
rect 17810 -1295 17815 -1275
rect 18055 -1275 18095 -1265
rect 18055 -1290 18065 -1275
rect 18040 -1295 18065 -1290
rect 18085 -1295 18095 -1275
rect 17505 -1305 17560 -1295
rect 17315 -1320 17330 -1305
rect 17545 -1320 17560 -1305
rect 17600 -1310 18000 -1295
rect 17600 -1320 17615 -1310
rect 17655 -1320 17670 -1310
rect 17710 -1320 17725 -1310
rect 17765 -1320 17780 -1310
rect 17820 -1320 17835 -1310
rect 17875 -1320 17890 -1310
rect 17930 -1320 17945 -1310
rect 17985 -1320 18000 -1310
rect 18040 -1305 18095 -1295
rect 18230 -1275 18270 -1265
rect 18230 -1295 18240 -1275
rect 18260 -1290 18270 -1275
rect 18400 -1275 18430 -1265
rect 18260 -1295 18285 -1290
rect 18400 -1295 18405 -1275
rect 18425 -1295 18430 -1275
rect 18670 -1275 18710 -1265
rect 18670 -1290 18680 -1275
rect 18655 -1295 18680 -1290
rect 18700 -1295 18710 -1275
rect 18230 -1305 18285 -1295
rect 18040 -1320 18055 -1305
rect 18270 -1320 18285 -1305
rect 18325 -1310 18615 -1295
rect 18325 -1320 18340 -1310
rect 18380 -1320 18395 -1310
rect 18435 -1320 18450 -1310
rect 18490 -1320 18505 -1310
rect 18545 -1320 18560 -1310
rect 18600 -1320 18615 -1310
rect 18655 -1305 18710 -1295
rect 18655 -1320 18670 -1305
rect 16930 -1435 16945 -1420
rect 16985 -1435 17000 -1420
rect 17040 -1435 17055 -1420
rect 17095 -1435 17110 -1420
rect 17150 -1435 17165 -1420
rect 17205 -1435 17220 -1420
rect 17260 -1435 17275 -1420
rect 17315 -1435 17330 -1420
rect 17545 -1435 17560 -1420
rect 17600 -1435 17615 -1420
rect 17655 -1435 17670 -1420
rect 17710 -1435 17725 -1420
rect 17765 -1435 17780 -1420
rect 17820 -1435 17835 -1420
rect 17875 -1435 17890 -1420
rect 17930 -1435 17945 -1420
rect 17985 -1435 18000 -1420
rect 18040 -1435 18055 -1420
rect 18270 -1435 18285 -1420
rect 18325 -1435 18340 -1420
rect 18380 -1435 18395 -1420
rect 18435 -1435 18450 -1420
rect 18490 -1435 18505 -1420
rect 18545 -1435 18560 -1420
rect 18600 -1435 18615 -1420
rect 18655 -1435 18670 -1420
rect 17585 -1445 17625 -1435
rect 17585 -1465 17595 -1445
rect 17615 -1465 17625 -1445
rect 17585 -1475 17625 -1465
<< polycont >>
rect 16250 1255 16270 1275
rect 16399 1255 16419 1275
rect 16470 1255 16490 1275
rect 16820 1255 16840 1275
rect 16985 1255 17005 1275
rect 17150 1255 17170 1275
rect 17615 1255 17635 1275
rect 17845 1255 17865 1275
rect 17965 1255 17985 1275
rect 18430 1255 18450 1275
rect 18595 1255 18615 1275
rect 18760 1255 18780 1275
rect 16980 790 17000 810
rect 18600 790 18620 810
rect 16445 690 16465 710
rect 16665 690 16685 710
rect 16555 520 16575 540
rect 18955 740 18975 760
rect 19130 740 19150 760
rect 19036 470 19056 490
rect 17700 420 17720 440
rect 18420 420 18440 440
rect 16430 100 16450 120
rect 17630 100 17650 120
rect 17950 100 17970 120
rect 19150 100 19170 120
rect 16430 -70 16450 -50
rect 16520 -70 16540 -50
rect 16610 -70 16630 -50
rect 16850 -70 16870 -50
rect 16970 -70 16990 -50
rect 17210 -70 17230 -50
rect 17330 -70 17350 -50
rect 17540 -70 17560 -50
rect 17950 -70 17970 -50
rect 18040 -70 18060 -50
rect 18250 -70 18270 -50
rect 18370 -70 18390 -50
rect 18610 -70 18630 -50
rect 18730 -70 18750 -50
rect 18970 -70 18990 -50
rect 19060 -70 19080 -50
rect 19150 -70 19170 -50
rect 16920 -230 16940 -210
rect 18660 -230 18680 -210
rect 16860 -395 16880 -375
rect 18720 -395 18740 -375
rect 16630 -555 16650 -535
rect 16750 -555 16770 -535
rect 16870 -555 16890 -535
rect 16990 -555 17010 -535
rect 17310 -555 17330 -535
rect 17430 -555 17450 -535
rect 17550 -555 17570 -535
rect 18030 -555 18050 -535
rect 18150 -555 18170 -535
rect 18270 -555 18290 -535
rect 18590 -555 18610 -535
rect 18710 -555 18730 -535
rect 18830 -555 18850 -535
rect 18950 -555 18970 -535
rect 16830 -1020 16850 -1000
rect 16910 -1020 16930 -1000
rect 16990 -1020 17010 -1000
rect 17070 -1020 17090 -1000
rect 17150 -1020 17170 -1000
rect 17230 -1020 17250 -1000
rect 17310 -1020 17330 -1000
rect 17390 -1020 17410 -1000
rect 17470 -1020 17490 -1000
rect 17550 -1020 17570 -1000
rect 17630 -1020 17650 -1000
rect 17710 -1020 17730 -1000
rect 17870 -1020 17890 -1000
rect 17950 -1020 17970 -1000
rect 18030 -1020 18050 -1000
rect 18110 -1020 18130 -1000
rect 18190 -1020 18210 -1000
rect 18270 -1020 18290 -1000
rect 18350 -1020 18370 -1000
rect 18430 -1020 18450 -1000
rect 18510 -1020 18530 -1000
rect 18590 -1020 18610 -1000
rect 18670 -1020 18690 -1000
rect 18750 -1020 18770 -1000
rect 16900 -1295 16920 -1275
rect 17175 -1295 17195 -1275
rect 17340 -1295 17360 -1275
rect 17515 -1295 17535 -1275
rect 17790 -1295 17810 -1275
rect 18065 -1295 18085 -1275
rect 18240 -1295 18260 -1275
rect 18405 -1295 18425 -1275
rect 18680 -1295 18700 -1275
rect 17595 -1465 17615 -1445
<< xpolycontact >>
rect 17470 -1930 17690 -1895
rect 17904 -1930 18124 -1895
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3252 19320 -3032
rect 19285 -3889 19320 -3669
rect 19345 -3252 19380 -3032
rect 19345 -3889 19380 -3669
rect 19405 -3252 19440 -3032
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -1930 17904 -1895
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3252
rect 19345 -3669 19380 -3252
rect 19405 -3669 19440 -3252
<< locali >>
rect 16240 1275 16280 1285
rect 16240 1255 16250 1275
rect 16270 1255 16280 1275
rect 16240 1245 16280 1255
rect 16335 1275 16375 1285
rect 16335 1255 16345 1275
rect 16365 1255 16375 1275
rect 16335 1245 16375 1255
rect 16394 1275 16424 1285
rect 16394 1255 16399 1275
rect 16419 1255 16424 1275
rect 16394 1245 16424 1255
rect 16460 1275 16500 1285
rect 16460 1255 16470 1275
rect 16490 1255 16500 1275
rect 16460 1245 16500 1255
rect 16810 1275 16850 1285
rect 16810 1255 16820 1275
rect 16840 1255 16850 1275
rect 16810 1245 16850 1255
rect 16920 1275 16960 1285
rect 16920 1255 16930 1275
rect 16950 1255 16960 1275
rect 16920 1245 16960 1255
rect 16980 1275 17010 1285
rect 16980 1255 16985 1275
rect 17005 1255 17010 1275
rect 16980 1245 17010 1255
rect 17030 1275 17070 1285
rect 17030 1255 17040 1275
rect 17060 1255 17070 1275
rect 17030 1245 17070 1255
rect 17090 1275 17120 1285
rect 17090 1255 17095 1275
rect 17115 1255 17120 1275
rect 17090 1245 17120 1255
rect 17140 1275 17180 1285
rect 17140 1255 17150 1275
rect 17170 1255 17180 1275
rect 17140 1245 17180 1255
rect 17605 1275 17645 1285
rect 17605 1255 17615 1275
rect 17635 1255 17645 1275
rect 17605 1245 17645 1255
rect 17670 1275 17710 1285
rect 17670 1255 17680 1275
rect 17700 1255 17710 1275
rect 17670 1245 17710 1255
rect 17730 1275 17760 1285
rect 17730 1255 17735 1275
rect 17755 1255 17760 1275
rect 17730 1245 17760 1255
rect 17780 1275 17820 1285
rect 17780 1255 17790 1275
rect 17810 1255 17820 1275
rect 17780 1245 17820 1255
rect 17840 1275 17870 1285
rect 17840 1255 17845 1275
rect 17865 1255 17870 1275
rect 17840 1245 17870 1255
rect 17890 1275 17930 1285
rect 17890 1255 17900 1275
rect 17920 1255 17930 1275
rect 17890 1245 17930 1255
rect 17955 1275 17995 1285
rect 17955 1255 17965 1275
rect 17985 1255 17995 1275
rect 17955 1245 17995 1255
rect 18420 1275 18460 1285
rect 18420 1255 18430 1275
rect 18450 1255 18460 1275
rect 18420 1245 18460 1255
rect 18480 1275 18510 1285
rect 18480 1255 18485 1275
rect 18505 1255 18510 1275
rect 18480 1245 18510 1255
rect 18530 1275 18570 1285
rect 18530 1255 18540 1275
rect 18560 1255 18570 1275
rect 18530 1245 18570 1255
rect 18590 1275 18620 1285
rect 18590 1255 18595 1275
rect 18615 1255 18620 1275
rect 18590 1245 18620 1255
rect 18640 1275 18680 1285
rect 18640 1255 18650 1275
rect 18670 1255 18680 1275
rect 18640 1245 18680 1255
rect 18750 1275 18790 1285
rect 18750 1255 18760 1275
rect 18780 1255 18790 1275
rect 18750 1245 18790 1255
rect 16250 1225 16270 1245
rect 16355 1225 16375 1245
rect 16470 1225 16490 1245
rect 16820 1225 16840 1245
rect 16930 1225 16950 1245
rect 17040 1225 17060 1245
rect 17095 1225 17115 1245
rect 17150 1225 17170 1245
rect 17625 1225 17645 1245
rect 17680 1225 17700 1245
rect 17735 1225 17755 1245
rect 17790 1225 17810 1245
rect 17900 1225 17920 1245
rect 17955 1225 17975 1245
rect 18430 1225 18450 1245
rect 18485 1225 18505 1245
rect 18540 1225 18560 1245
rect 18650 1225 18670 1245
rect 18760 1225 18780 1245
rect 16205 1217 16275 1225
rect 16205 1145 16210 1217
rect 16230 1215 16275 1217
rect 16230 1145 16250 1215
rect 16205 1143 16250 1145
rect 16270 1143 16275 1215
rect 16205 1135 16275 1143
rect 16300 1215 16330 1225
rect 16300 1143 16305 1215
rect 16325 1143 16330 1215
rect 16300 1135 16330 1143
rect 16355 1215 16385 1225
rect 16355 1143 16360 1215
rect 16380 1143 16385 1215
rect 16355 1135 16385 1143
rect 16410 1215 16440 1225
rect 16410 1143 16415 1215
rect 16435 1143 16440 1215
rect 16410 1135 16440 1143
rect 16465 1217 16535 1225
rect 16465 1215 16510 1217
rect 16465 1143 16470 1215
rect 16490 1145 16510 1215
rect 16530 1145 16535 1217
rect 16490 1143 16535 1145
rect 16465 1135 16535 1143
rect 16775 1217 16845 1225
rect 16775 1145 16780 1217
rect 16800 1215 16845 1217
rect 16800 1145 16820 1215
rect 16775 1143 16820 1145
rect 16840 1143 16845 1215
rect 16775 1135 16845 1143
rect 16870 1215 16900 1225
rect 16870 1143 16875 1215
rect 16895 1143 16900 1215
rect 16870 1135 16900 1143
rect 16925 1215 16955 1225
rect 16925 1143 16930 1215
rect 16950 1143 16955 1215
rect 16925 1135 16955 1143
rect 16980 1215 17010 1225
rect 16980 1143 16985 1215
rect 17005 1143 17010 1215
rect 16980 1135 17010 1143
rect 17035 1215 17065 1225
rect 17035 1143 17040 1215
rect 17060 1143 17065 1215
rect 17035 1135 17065 1143
rect 17090 1215 17120 1225
rect 17090 1143 17095 1215
rect 17115 1143 17120 1215
rect 17090 1135 17120 1143
rect 17145 1217 17215 1225
rect 17145 1215 17190 1217
rect 17145 1143 17150 1215
rect 17170 1145 17190 1215
rect 17210 1145 17215 1217
rect 17170 1143 17215 1145
rect 17145 1135 17215 1143
rect 17580 1215 17650 1225
rect 17580 1195 17585 1215
rect 17605 1195 17625 1215
rect 17645 1195 17650 1215
rect 17580 1165 17650 1195
rect 17580 1145 17585 1165
rect 17605 1145 17625 1165
rect 17645 1145 17650 1165
rect 16305 1115 16325 1135
rect 16415 1115 16435 1135
rect 16875 1115 16895 1135
rect 16985 1115 17005 1135
rect 17095 1115 17115 1135
rect 17580 1115 17650 1145
rect 16300 1105 16330 1115
rect 16300 1085 16305 1105
rect 16325 1085 16330 1105
rect 16300 1075 16330 1085
rect 16410 1105 16440 1115
rect 16410 1085 16415 1105
rect 16435 1085 16440 1105
rect 16410 1075 16440 1085
rect 16865 1105 16905 1115
rect 16865 1085 16875 1105
rect 16895 1085 16905 1105
rect 16865 1075 16905 1085
rect 16975 1105 17015 1115
rect 16975 1085 16985 1105
rect 17005 1085 17015 1105
rect 16975 1075 17015 1085
rect 17085 1105 17125 1115
rect 17085 1085 17095 1105
rect 17115 1085 17125 1105
rect 17085 1075 17125 1085
rect 17580 1095 17585 1115
rect 17605 1095 17625 1115
rect 17645 1095 17650 1115
rect 17580 1065 17650 1095
rect 17580 1045 17585 1065
rect 17605 1045 17625 1065
rect 17645 1045 17650 1065
rect 17580 1035 17650 1045
rect 17675 1215 17705 1225
rect 17675 1195 17680 1215
rect 17700 1195 17705 1215
rect 17675 1165 17705 1195
rect 17675 1145 17680 1165
rect 17700 1145 17705 1165
rect 17675 1115 17705 1145
rect 17675 1095 17680 1115
rect 17700 1095 17705 1115
rect 17675 1065 17705 1095
rect 17675 1045 17680 1065
rect 17700 1045 17705 1065
rect 17675 1035 17705 1045
rect 17730 1215 17760 1225
rect 17730 1195 17735 1215
rect 17755 1195 17760 1215
rect 17730 1165 17760 1195
rect 17730 1145 17735 1165
rect 17755 1145 17760 1165
rect 17730 1115 17760 1145
rect 17730 1095 17735 1115
rect 17755 1095 17760 1115
rect 17730 1065 17760 1095
rect 17730 1045 17735 1065
rect 17755 1045 17760 1065
rect 17730 1035 17760 1045
rect 17785 1215 17815 1225
rect 17785 1195 17790 1215
rect 17810 1195 17815 1215
rect 17785 1165 17815 1195
rect 17785 1145 17790 1165
rect 17810 1145 17815 1165
rect 17785 1115 17815 1145
rect 17785 1095 17790 1115
rect 17810 1095 17815 1115
rect 17785 1065 17815 1095
rect 17785 1045 17790 1065
rect 17810 1045 17815 1065
rect 17785 1035 17815 1045
rect 17840 1215 17870 1225
rect 17840 1195 17845 1215
rect 17865 1195 17870 1215
rect 17840 1165 17870 1195
rect 17840 1145 17845 1165
rect 17865 1145 17870 1165
rect 17840 1115 17870 1145
rect 17840 1095 17845 1115
rect 17865 1095 17870 1115
rect 17840 1065 17870 1095
rect 17840 1045 17845 1065
rect 17865 1045 17870 1065
rect 17840 1035 17870 1045
rect 17895 1215 17925 1225
rect 17895 1195 17900 1215
rect 17920 1195 17925 1215
rect 17895 1165 17925 1195
rect 17895 1145 17900 1165
rect 17920 1145 17925 1165
rect 17895 1115 17925 1145
rect 17895 1095 17900 1115
rect 17920 1095 17925 1115
rect 17895 1065 17925 1095
rect 17895 1045 17900 1065
rect 17920 1045 17925 1065
rect 17895 1035 17925 1045
rect 17950 1215 18020 1225
rect 17950 1195 17955 1215
rect 17975 1195 17995 1215
rect 18015 1195 18020 1215
rect 17950 1165 18020 1195
rect 17950 1145 17955 1165
rect 17975 1145 17995 1165
rect 18015 1145 18020 1165
rect 17950 1115 18020 1145
rect 18385 1217 18455 1225
rect 18385 1145 18390 1217
rect 18410 1215 18455 1217
rect 18410 1145 18430 1215
rect 18450 1145 18455 1215
rect 18385 1135 18455 1145
rect 18480 1215 18510 1225
rect 18480 1145 18485 1215
rect 18505 1145 18510 1215
rect 18480 1135 18510 1145
rect 18535 1215 18565 1225
rect 18535 1145 18540 1215
rect 18560 1145 18565 1215
rect 18535 1135 18565 1145
rect 18590 1215 18620 1225
rect 18590 1145 18595 1215
rect 18615 1145 18620 1215
rect 18590 1135 18620 1145
rect 18645 1215 18675 1225
rect 18645 1145 18650 1215
rect 18670 1145 18675 1215
rect 18645 1135 18675 1145
rect 18700 1215 18730 1225
rect 18700 1145 18705 1215
rect 18725 1145 18730 1215
rect 18700 1135 18730 1145
rect 18755 1217 18825 1225
rect 18755 1215 18800 1217
rect 18755 1145 18760 1215
rect 18780 1145 18800 1215
rect 18820 1145 18825 1217
rect 18755 1135 18825 1145
rect 18485 1115 18505 1135
rect 18595 1115 18615 1135
rect 18705 1115 18725 1135
rect 17950 1095 17955 1115
rect 17975 1095 17995 1115
rect 18015 1095 18020 1115
rect 17950 1065 18020 1095
rect 18475 1105 18515 1115
rect 18475 1085 18485 1105
rect 18505 1085 18515 1105
rect 18475 1075 18515 1085
rect 18585 1105 18625 1115
rect 18585 1085 18595 1105
rect 18615 1085 18625 1105
rect 18585 1075 18625 1085
rect 18695 1105 18735 1115
rect 18695 1085 18705 1105
rect 18725 1085 18735 1105
rect 18695 1075 18735 1085
rect 17950 1045 17955 1065
rect 17975 1045 17995 1065
rect 18015 1045 18020 1065
rect 17950 1035 18020 1045
rect 17735 1015 17755 1035
rect 17845 1015 17865 1035
rect 17725 1005 17765 1015
rect 17725 985 17735 1005
rect 17755 985 17765 1005
rect 17725 975 17765 985
rect 17835 1005 17875 1015
rect 17835 985 17845 1005
rect 17865 985 17875 1005
rect 17835 975 17875 985
rect 16970 810 17010 820
rect 16970 790 16980 810
rect 17000 790 17010 810
rect 16970 780 17010 790
rect 17150 810 17190 820
rect 17150 790 17160 810
rect 17180 790 17190 810
rect 17150 780 17190 790
rect 17330 810 17370 820
rect 17330 790 17340 810
rect 17360 790 17370 810
rect 17330 780 17370 790
rect 17510 810 17550 820
rect 17510 790 17520 810
rect 17540 790 17550 810
rect 17510 780 17550 790
rect 17690 810 17730 820
rect 17690 790 17700 810
rect 17720 790 17730 810
rect 17690 780 17730 790
rect 17870 810 17910 820
rect 17870 790 17880 810
rect 17900 790 17910 810
rect 17870 780 17910 790
rect 18050 810 18090 820
rect 18050 790 18060 810
rect 18080 790 18090 810
rect 18050 780 18090 790
rect 18230 810 18270 820
rect 18230 790 18240 810
rect 18260 790 18270 810
rect 18230 780 18270 790
rect 18410 810 18450 820
rect 18410 790 18420 810
rect 18440 790 18450 810
rect 18410 780 18450 790
rect 18590 810 18630 820
rect 18590 790 18600 810
rect 18620 790 18630 810
rect 18590 780 18630 790
rect 16980 760 17000 780
rect 17160 760 17180 780
rect 17340 760 17360 780
rect 17520 760 17540 780
rect 17700 760 17720 780
rect 17880 760 17900 780
rect 18060 760 18080 780
rect 18240 760 18260 780
rect 18420 760 18440 780
rect 18600 760 18620 780
rect 18945 760 18985 770
rect 16935 750 17005 760
rect 16935 730 16940 750
rect 16960 730 16980 750
rect 17000 730 17005 750
rect 16440 710 16470 720
rect 16440 690 16445 710
rect 16465 690 16470 710
rect 16440 660 16470 690
rect 16545 710 16585 720
rect 16545 690 16555 710
rect 16575 690 16585 710
rect 16545 680 16585 690
rect 16655 710 16695 720
rect 16655 690 16665 710
rect 16685 690 16695 710
rect 16655 680 16695 690
rect 16935 700 17005 730
rect 16935 680 16940 700
rect 16960 680 16980 700
rect 17000 680 17005 700
rect 16555 660 16575 680
rect 16660 660 16690 680
rect 16400 650 16470 660
rect 16400 630 16405 650
rect 16425 630 16445 650
rect 16465 630 16470 650
rect 16400 600 16470 630
rect 16400 580 16405 600
rect 16425 580 16445 600
rect 16465 580 16470 600
rect 16400 570 16470 580
rect 16495 650 16525 660
rect 16495 630 16500 650
rect 16520 630 16525 650
rect 16495 600 16525 630
rect 16495 580 16500 600
rect 16520 580 16525 600
rect 16495 570 16525 580
rect 16550 650 16580 660
rect 16550 630 16555 650
rect 16575 630 16580 650
rect 16550 600 16580 630
rect 16550 580 16555 600
rect 16575 580 16580 600
rect 16550 570 16580 580
rect 16605 650 16635 660
rect 16605 630 16610 650
rect 16630 630 16635 650
rect 16605 600 16635 630
rect 16605 580 16610 600
rect 16630 580 16635 600
rect 16605 570 16635 580
rect 16660 650 16735 660
rect 16660 630 16665 650
rect 16685 630 16710 650
rect 16730 630 16735 650
rect 16660 600 16735 630
rect 16660 580 16665 600
rect 16685 580 16710 600
rect 16730 580 16735 600
rect 16660 570 16735 580
rect 16935 650 17005 680
rect 16935 630 16940 650
rect 16960 630 16980 650
rect 17000 630 17005 650
rect 16935 600 17005 630
rect 16935 580 16940 600
rect 16960 580 16980 600
rect 17000 580 17005 600
rect 16500 550 16520 570
rect 16610 550 16630 570
rect 16935 550 17005 580
rect 16480 540 16520 550
rect 16480 520 16490 540
rect 16510 520 16520 540
rect 16480 510 16520 520
rect 16545 540 16585 550
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 16610 540 16650 550
rect 16610 520 16620 540
rect 16640 520 16650 540
rect 16610 510 16650 520
rect 16935 530 16940 550
rect 16960 530 16980 550
rect 17000 530 17005 550
rect 16935 500 17005 530
rect 16935 480 16940 500
rect 16960 480 16980 500
rect 17000 480 17005 500
rect 16935 470 17005 480
rect 17065 750 17095 760
rect 17065 730 17070 750
rect 17090 730 17095 750
rect 17065 700 17095 730
rect 17065 680 17070 700
rect 17090 680 17095 700
rect 17065 650 17095 680
rect 17065 630 17070 650
rect 17090 630 17095 650
rect 17065 600 17095 630
rect 17065 580 17070 600
rect 17090 580 17095 600
rect 17065 550 17095 580
rect 17065 530 17070 550
rect 17090 530 17095 550
rect 17065 500 17095 530
rect 17065 480 17070 500
rect 17090 480 17095 500
rect 17065 470 17095 480
rect 17155 750 17185 760
rect 17155 730 17160 750
rect 17180 730 17185 750
rect 17155 700 17185 730
rect 17155 680 17160 700
rect 17180 680 17185 700
rect 17155 650 17185 680
rect 17155 630 17160 650
rect 17180 630 17185 650
rect 17155 600 17185 630
rect 17155 580 17160 600
rect 17180 580 17185 600
rect 17155 550 17185 580
rect 17155 530 17160 550
rect 17180 530 17185 550
rect 17155 500 17185 530
rect 17155 480 17160 500
rect 17180 480 17185 500
rect 17155 470 17185 480
rect 17245 750 17275 760
rect 17245 730 17250 750
rect 17270 730 17275 750
rect 17245 700 17275 730
rect 17245 680 17250 700
rect 17270 680 17275 700
rect 17245 650 17275 680
rect 17245 630 17250 650
rect 17270 630 17275 650
rect 17245 600 17275 630
rect 17245 580 17250 600
rect 17270 580 17275 600
rect 17245 550 17275 580
rect 17245 530 17250 550
rect 17270 530 17275 550
rect 17245 500 17275 530
rect 17245 480 17250 500
rect 17270 480 17275 500
rect 17245 470 17275 480
rect 17335 750 17365 760
rect 17335 730 17340 750
rect 17360 730 17365 750
rect 17335 700 17365 730
rect 17335 680 17340 700
rect 17360 680 17365 700
rect 17335 650 17365 680
rect 17335 630 17340 650
rect 17360 630 17365 650
rect 17335 600 17365 630
rect 17335 580 17340 600
rect 17360 580 17365 600
rect 17335 550 17365 580
rect 17335 530 17340 550
rect 17360 530 17365 550
rect 17335 500 17365 530
rect 17335 480 17340 500
rect 17360 480 17365 500
rect 17335 470 17365 480
rect 17425 750 17455 760
rect 17425 730 17430 750
rect 17450 730 17455 750
rect 17425 700 17455 730
rect 17425 680 17430 700
rect 17450 680 17455 700
rect 17425 650 17455 680
rect 17425 630 17430 650
rect 17450 630 17455 650
rect 17425 600 17455 630
rect 17425 580 17430 600
rect 17450 580 17455 600
rect 17425 550 17455 580
rect 17425 530 17430 550
rect 17450 530 17455 550
rect 17425 500 17455 530
rect 17425 480 17430 500
rect 17450 480 17455 500
rect 17425 470 17455 480
rect 17515 750 17545 760
rect 17515 730 17520 750
rect 17540 730 17545 750
rect 17515 700 17545 730
rect 17515 680 17520 700
rect 17540 680 17545 700
rect 17515 650 17545 680
rect 17515 630 17520 650
rect 17540 630 17545 650
rect 17515 600 17545 630
rect 17515 580 17520 600
rect 17540 580 17545 600
rect 17515 550 17545 580
rect 17515 530 17520 550
rect 17540 530 17545 550
rect 17515 500 17545 530
rect 17515 480 17520 500
rect 17540 480 17545 500
rect 17515 470 17545 480
rect 17605 750 17635 760
rect 17605 730 17610 750
rect 17630 730 17635 750
rect 17605 700 17635 730
rect 17605 680 17610 700
rect 17630 680 17635 700
rect 17605 650 17635 680
rect 17605 630 17610 650
rect 17630 630 17635 650
rect 17605 600 17635 630
rect 17605 580 17610 600
rect 17630 580 17635 600
rect 17605 550 17635 580
rect 17605 530 17610 550
rect 17630 530 17635 550
rect 17605 500 17635 530
rect 17605 480 17610 500
rect 17630 480 17635 500
rect 17605 470 17635 480
rect 17695 750 17725 760
rect 17695 730 17700 750
rect 17720 730 17725 750
rect 17695 700 17725 730
rect 17695 680 17700 700
rect 17720 680 17725 700
rect 17695 650 17725 680
rect 17695 630 17700 650
rect 17720 630 17725 650
rect 17695 600 17725 630
rect 17695 580 17700 600
rect 17720 580 17725 600
rect 17695 550 17725 580
rect 17695 530 17700 550
rect 17720 530 17725 550
rect 17695 500 17725 530
rect 17695 480 17700 500
rect 17720 480 17725 500
rect 17695 470 17725 480
rect 17785 750 17815 760
rect 17785 730 17790 750
rect 17810 730 17815 750
rect 17785 700 17815 730
rect 17785 680 17790 700
rect 17810 680 17815 700
rect 17785 650 17815 680
rect 17785 630 17790 650
rect 17810 630 17815 650
rect 17785 600 17815 630
rect 17785 580 17790 600
rect 17810 580 17815 600
rect 17785 550 17815 580
rect 17785 530 17790 550
rect 17810 530 17815 550
rect 17785 500 17815 530
rect 17785 480 17790 500
rect 17810 480 17815 500
rect 17785 470 17815 480
rect 17875 750 17905 760
rect 17875 730 17880 750
rect 17900 730 17905 750
rect 17875 700 17905 730
rect 17875 680 17880 700
rect 17900 680 17905 700
rect 17875 650 17905 680
rect 17875 630 17880 650
rect 17900 630 17905 650
rect 17875 600 17905 630
rect 17875 580 17880 600
rect 17900 580 17905 600
rect 17875 550 17905 580
rect 17875 530 17880 550
rect 17900 530 17905 550
rect 17875 500 17905 530
rect 17875 480 17880 500
rect 17900 480 17905 500
rect 17875 470 17905 480
rect 17965 750 17995 760
rect 17965 730 17970 750
rect 17990 730 17995 750
rect 17965 700 17995 730
rect 17965 680 17970 700
rect 17990 680 17995 700
rect 17965 650 17995 680
rect 17965 630 17970 650
rect 17990 630 17995 650
rect 17965 600 17995 630
rect 17965 580 17970 600
rect 17990 580 17995 600
rect 17965 550 17995 580
rect 17965 530 17970 550
rect 17990 530 17995 550
rect 17965 500 17995 530
rect 17965 480 17970 500
rect 17990 480 17995 500
rect 17965 470 17995 480
rect 18055 750 18085 760
rect 18055 730 18060 750
rect 18080 730 18085 750
rect 18055 700 18085 730
rect 18055 680 18060 700
rect 18080 680 18085 700
rect 18055 650 18085 680
rect 18055 630 18060 650
rect 18080 630 18085 650
rect 18055 600 18085 630
rect 18055 580 18060 600
rect 18080 580 18085 600
rect 18055 550 18085 580
rect 18055 530 18060 550
rect 18080 530 18085 550
rect 18055 500 18085 530
rect 18055 480 18060 500
rect 18080 480 18085 500
rect 18055 470 18085 480
rect 18145 750 18175 760
rect 18145 730 18150 750
rect 18170 730 18175 750
rect 18145 700 18175 730
rect 18145 680 18150 700
rect 18170 680 18175 700
rect 18145 650 18175 680
rect 18145 630 18150 650
rect 18170 630 18175 650
rect 18145 600 18175 630
rect 18145 580 18150 600
rect 18170 580 18175 600
rect 18145 550 18175 580
rect 18145 530 18150 550
rect 18170 530 18175 550
rect 18145 500 18175 530
rect 18145 480 18150 500
rect 18170 480 18175 500
rect 18145 470 18175 480
rect 18235 750 18265 760
rect 18235 730 18240 750
rect 18260 730 18265 750
rect 18235 700 18265 730
rect 18235 680 18240 700
rect 18260 680 18265 700
rect 18235 650 18265 680
rect 18235 630 18240 650
rect 18260 630 18265 650
rect 18235 600 18265 630
rect 18235 580 18240 600
rect 18260 580 18265 600
rect 18235 550 18265 580
rect 18235 530 18240 550
rect 18260 530 18265 550
rect 18235 500 18265 530
rect 18235 480 18240 500
rect 18260 480 18265 500
rect 18235 470 18265 480
rect 18325 750 18355 760
rect 18325 730 18330 750
rect 18350 730 18355 750
rect 18325 700 18355 730
rect 18325 680 18330 700
rect 18350 680 18355 700
rect 18325 650 18355 680
rect 18325 630 18330 650
rect 18350 630 18355 650
rect 18325 600 18355 630
rect 18325 580 18330 600
rect 18350 580 18355 600
rect 18325 550 18355 580
rect 18325 530 18330 550
rect 18350 530 18355 550
rect 18325 500 18355 530
rect 18325 480 18330 500
rect 18350 480 18355 500
rect 18325 470 18355 480
rect 18415 750 18445 760
rect 18415 730 18420 750
rect 18440 730 18445 750
rect 18415 700 18445 730
rect 18415 680 18420 700
rect 18440 680 18445 700
rect 18415 650 18445 680
rect 18415 630 18420 650
rect 18440 630 18445 650
rect 18415 600 18445 630
rect 18415 580 18420 600
rect 18440 580 18445 600
rect 18415 550 18445 580
rect 18415 530 18420 550
rect 18440 530 18445 550
rect 18415 500 18445 530
rect 18415 480 18420 500
rect 18440 480 18445 500
rect 18415 470 18445 480
rect 18505 750 18535 760
rect 18505 730 18510 750
rect 18530 730 18535 750
rect 18505 700 18535 730
rect 18505 680 18510 700
rect 18530 680 18535 700
rect 18505 650 18535 680
rect 18505 630 18510 650
rect 18530 630 18535 650
rect 18505 600 18535 630
rect 18505 580 18510 600
rect 18530 580 18535 600
rect 18505 550 18535 580
rect 18505 530 18510 550
rect 18530 530 18535 550
rect 18505 500 18535 530
rect 18505 480 18510 500
rect 18530 480 18535 500
rect 18505 470 18535 480
rect 18595 750 18665 760
rect 18595 730 18600 750
rect 18620 730 18640 750
rect 18660 730 18665 750
rect 18945 740 18955 760
rect 18975 740 18985 760
rect 18945 730 18985 740
rect 19010 760 19050 770
rect 19010 740 19020 760
rect 19040 740 19050 760
rect 19010 730 19050 740
rect 19120 760 19160 770
rect 19120 740 19130 760
rect 19150 740 19160 760
rect 19120 730 19160 740
rect 18595 700 18665 730
rect 18965 710 18985 730
rect 19020 710 19040 730
rect 19130 710 19150 730
rect 18595 680 18600 700
rect 18620 680 18640 700
rect 18660 680 18665 700
rect 18595 650 18665 680
rect 18595 630 18600 650
rect 18620 630 18640 650
rect 18660 630 18665 650
rect 18595 600 18665 630
rect 18595 580 18600 600
rect 18620 580 18640 600
rect 18660 580 18665 600
rect 18595 550 18665 580
rect 18595 530 18600 550
rect 18620 530 18640 550
rect 18660 530 18665 550
rect 18595 500 18665 530
rect 18920 700 18990 710
rect 18920 680 18925 700
rect 18945 680 18965 700
rect 18985 680 18990 700
rect 18920 650 18990 680
rect 18920 630 18925 650
rect 18945 630 18965 650
rect 18985 630 18990 650
rect 18920 600 18990 630
rect 18920 580 18925 600
rect 18945 580 18965 600
rect 18985 580 18990 600
rect 18920 550 18990 580
rect 18920 530 18925 550
rect 18945 530 18965 550
rect 18985 530 18990 550
rect 18920 520 18990 530
rect 19015 700 19045 710
rect 19015 680 19020 700
rect 19040 680 19045 700
rect 19015 650 19045 680
rect 19015 630 19020 650
rect 19040 630 19045 650
rect 19015 600 19045 630
rect 19015 580 19020 600
rect 19040 580 19045 600
rect 19015 550 19045 580
rect 19015 530 19020 550
rect 19040 530 19045 550
rect 19015 520 19045 530
rect 19070 700 19100 710
rect 19070 680 19075 700
rect 19095 680 19100 700
rect 19070 650 19100 680
rect 19070 630 19075 650
rect 19095 630 19100 650
rect 19070 600 19100 630
rect 19070 580 19075 600
rect 19095 580 19100 600
rect 19070 550 19100 580
rect 19070 530 19075 550
rect 19095 530 19100 550
rect 19070 520 19100 530
rect 19125 700 19195 710
rect 19125 680 19130 700
rect 19150 680 19170 700
rect 19190 680 19195 700
rect 19125 650 19195 680
rect 19125 630 19130 650
rect 19150 630 19170 650
rect 19190 630 19195 650
rect 19125 600 19195 630
rect 19125 580 19130 600
rect 19150 580 19170 600
rect 19190 580 19195 600
rect 19125 550 19195 580
rect 19125 530 19130 550
rect 19150 530 19170 550
rect 19190 530 19195 550
rect 19125 520 19195 530
rect 19080 500 19100 520
rect 18595 480 18600 500
rect 18620 480 18640 500
rect 18660 480 18665 500
rect 18595 470 18665 480
rect 19031 490 19061 500
rect 19031 470 19036 490
rect 19056 470 19061 490
rect 17070 450 17090 470
rect 17250 450 17270 470
rect 17430 450 17450 470
rect 17610 450 17630 470
rect 17790 450 17810 470
rect 17970 450 17990 470
rect 18150 450 18170 470
rect 18330 450 18350 470
rect 18510 450 18530 470
rect 19031 460 19061 470
rect 19080 490 19120 500
rect 19080 470 19090 490
rect 19110 470 19120 490
rect 19080 460 19120 470
rect 17060 440 17100 450
rect 17060 420 17070 440
rect 17090 420 17100 440
rect 17060 410 17100 420
rect 17240 440 17280 450
rect 17240 420 17250 440
rect 17270 420 17280 440
rect 17240 410 17280 420
rect 17420 440 17460 450
rect 17420 420 17430 440
rect 17450 420 17460 440
rect 17420 410 17460 420
rect 17600 440 17640 450
rect 17600 420 17610 440
rect 17630 420 17640 440
rect 17600 410 17640 420
rect 17690 440 17730 450
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 17780 440 17820 450
rect 17780 420 17790 440
rect 17810 420 17820 440
rect 17780 410 17820 420
rect 17960 440 18000 450
rect 17960 420 17970 440
rect 17990 420 18000 440
rect 17960 410 18000 420
rect 18140 440 18180 450
rect 18140 420 18150 440
rect 18170 420 18180 440
rect 18140 410 18180 420
rect 18320 440 18360 450
rect 18320 420 18330 440
rect 18350 420 18360 440
rect 18320 410 18360 420
rect 18410 440 18450 450
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 18500 440 18540 450
rect 18500 420 18510 440
rect 18530 420 18540 440
rect 18500 410 18540 420
rect 16425 120 16455 130
rect 16425 100 16430 120
rect 16450 100 16455 120
rect 16425 70 16455 100
rect 16480 120 16520 130
rect 16480 100 16490 120
rect 16510 100 16520 120
rect 16480 90 16520 100
rect 16545 120 16575 130
rect 16545 100 16550 120
rect 16570 100 16575 120
rect 16545 90 16575 100
rect 16665 120 16695 130
rect 16665 100 16670 120
rect 16690 100 16695 120
rect 16665 90 16695 100
rect 16785 120 16815 130
rect 16785 100 16790 120
rect 16810 100 16815 120
rect 16785 90 16815 100
rect 16840 120 16880 130
rect 16840 100 16850 120
rect 16870 100 16880 120
rect 16840 90 16880 100
rect 16905 120 16935 130
rect 16905 100 16910 120
rect 16930 100 16935 120
rect 16905 90 16935 100
rect 17025 120 17055 130
rect 17025 100 17030 120
rect 17050 100 17055 120
rect 17025 90 17055 100
rect 17145 120 17175 130
rect 17145 100 17150 120
rect 17170 100 17175 120
rect 17145 90 17175 100
rect 17200 120 17240 130
rect 17200 100 17210 120
rect 17230 100 17240 120
rect 17200 90 17240 100
rect 17265 120 17295 130
rect 17265 100 17270 120
rect 17290 100 17295 120
rect 17265 90 17295 100
rect 17385 120 17415 130
rect 17385 100 17390 120
rect 17410 100 17415 120
rect 17385 90 17415 100
rect 17505 120 17535 130
rect 17505 100 17510 120
rect 17530 100 17535 120
rect 17505 90 17535 100
rect 17560 120 17600 130
rect 17560 100 17570 120
rect 17590 100 17600 120
rect 17560 90 17600 100
rect 17625 120 17655 130
rect 17625 100 17630 120
rect 17650 100 17655 120
rect 16490 70 16510 90
rect 16550 70 16570 90
rect 16670 70 16690 90
rect 16790 70 16810 90
rect 16850 70 16870 90
rect 16910 70 16930 90
rect 17030 70 17050 90
rect 17150 70 17170 90
rect 17210 70 17230 90
rect 17270 70 17290 90
rect 17390 70 17410 90
rect 17510 70 17530 90
rect 17570 70 17590 90
rect 17625 70 17655 100
rect 17945 120 17975 130
rect 17945 100 17950 120
rect 17970 100 17975 120
rect 17945 70 17975 100
rect 18000 120 18040 130
rect 18000 100 18010 120
rect 18030 100 18040 120
rect 18000 90 18040 100
rect 18065 120 18095 130
rect 18065 100 18070 120
rect 18090 100 18095 120
rect 18065 90 18095 100
rect 18185 120 18215 130
rect 18185 100 18190 120
rect 18210 100 18215 120
rect 18185 90 18215 100
rect 18305 120 18335 130
rect 18305 100 18310 120
rect 18330 100 18335 120
rect 18305 90 18335 100
rect 18360 120 18400 130
rect 18360 100 18370 120
rect 18390 100 18400 120
rect 18360 90 18400 100
rect 18425 120 18455 130
rect 18425 100 18430 120
rect 18450 100 18455 120
rect 18425 90 18455 100
rect 18545 120 18575 130
rect 18545 100 18550 120
rect 18570 100 18575 120
rect 18545 90 18575 100
rect 18665 120 18695 130
rect 18665 100 18670 120
rect 18690 100 18695 120
rect 18665 90 18695 100
rect 18720 120 18760 130
rect 18720 100 18730 120
rect 18750 100 18760 120
rect 18720 90 18760 100
rect 18785 120 18815 130
rect 18785 100 18790 120
rect 18810 100 18815 120
rect 18785 90 18815 100
rect 18905 120 18935 130
rect 18905 100 18910 120
rect 18930 100 18935 120
rect 18905 90 18935 100
rect 19025 120 19055 130
rect 19025 100 19030 120
rect 19050 100 19055 120
rect 19025 90 19055 100
rect 19080 120 19120 130
rect 19080 100 19090 120
rect 19110 100 19120 120
rect 19080 90 19120 100
rect 19145 120 19175 130
rect 19145 100 19150 120
rect 19170 100 19175 120
rect 18010 70 18030 90
rect 18070 70 18090 90
rect 18190 70 18210 90
rect 18310 70 18330 90
rect 18370 70 18390 90
rect 18430 70 18450 90
rect 18550 70 18570 90
rect 18670 70 18690 90
rect 18730 70 18750 90
rect 18790 70 18810 90
rect 18910 70 18930 90
rect 19030 70 19050 90
rect 19090 70 19110 90
rect 19145 70 19175 100
rect 16385 60 16455 70
rect 16385 40 16390 60
rect 16410 40 16430 60
rect 16450 40 16455 60
rect 16385 10 16455 40
rect 16385 -10 16390 10
rect 16410 -10 16430 10
rect 16450 -10 16455 10
rect 16385 -20 16455 -10
rect 16485 60 16515 70
rect 16485 40 16490 60
rect 16510 40 16515 60
rect 16485 10 16515 40
rect 16485 -10 16490 10
rect 16510 -10 16515 10
rect 16485 -20 16515 -10
rect 16545 60 16575 70
rect 16545 40 16550 60
rect 16570 40 16575 60
rect 16545 10 16575 40
rect 16545 -10 16550 10
rect 16570 -10 16575 10
rect 16545 -20 16575 -10
rect 16605 60 16635 70
rect 16605 40 16610 60
rect 16630 40 16635 60
rect 16605 10 16635 40
rect 16605 -10 16610 10
rect 16630 -10 16635 10
rect 16605 -20 16635 -10
rect 16665 60 16695 70
rect 16665 40 16670 60
rect 16690 40 16695 60
rect 16665 10 16695 40
rect 16665 -10 16670 10
rect 16690 -10 16695 10
rect 16665 -20 16695 -10
rect 16725 60 16755 70
rect 16725 40 16730 60
rect 16750 40 16755 60
rect 16725 10 16755 40
rect 16725 -10 16730 10
rect 16750 -10 16755 10
rect 16725 -20 16755 -10
rect 16785 60 16815 70
rect 16785 40 16790 60
rect 16810 40 16815 60
rect 16785 10 16815 40
rect 16785 -10 16790 10
rect 16810 -10 16815 10
rect 16785 -20 16815 -10
rect 16845 60 16875 70
rect 16845 40 16850 60
rect 16870 40 16875 60
rect 16845 10 16875 40
rect 16845 -10 16850 10
rect 16870 -10 16875 10
rect 16845 -20 16875 -10
rect 16905 60 16935 70
rect 16905 40 16910 60
rect 16930 40 16935 60
rect 16905 10 16935 40
rect 16905 -10 16910 10
rect 16930 -10 16935 10
rect 16905 -20 16935 -10
rect 16965 60 16995 70
rect 16965 40 16970 60
rect 16990 40 16995 60
rect 16965 10 16995 40
rect 16965 -10 16970 10
rect 16990 -10 16995 10
rect 16965 -20 16995 -10
rect 17025 60 17055 70
rect 17025 40 17030 60
rect 17050 40 17055 60
rect 17025 10 17055 40
rect 17025 -10 17030 10
rect 17050 -10 17055 10
rect 17025 -20 17055 -10
rect 17085 60 17115 70
rect 17085 40 17090 60
rect 17110 40 17115 60
rect 17085 10 17115 40
rect 17085 -10 17090 10
rect 17110 -10 17115 10
rect 17085 -20 17115 -10
rect 17145 60 17175 70
rect 17145 40 17150 60
rect 17170 40 17175 60
rect 17145 10 17175 40
rect 17145 -10 17150 10
rect 17170 -10 17175 10
rect 17145 -20 17175 -10
rect 17205 60 17235 70
rect 17205 40 17210 60
rect 17230 40 17235 60
rect 17205 10 17235 40
rect 17205 -10 17210 10
rect 17230 -10 17235 10
rect 17205 -20 17235 -10
rect 17265 60 17295 70
rect 17265 40 17270 60
rect 17290 40 17295 60
rect 17265 10 17295 40
rect 17265 -10 17270 10
rect 17290 -10 17295 10
rect 17265 -20 17295 -10
rect 17325 60 17355 70
rect 17325 40 17330 60
rect 17350 40 17355 60
rect 17325 10 17355 40
rect 17325 -10 17330 10
rect 17350 -10 17355 10
rect 17325 -20 17355 -10
rect 17385 60 17415 70
rect 17385 40 17390 60
rect 17410 40 17415 60
rect 17385 10 17415 40
rect 17385 -10 17390 10
rect 17410 -10 17415 10
rect 17385 -20 17415 -10
rect 17445 60 17475 70
rect 17445 40 17450 60
rect 17470 40 17475 60
rect 17445 10 17475 40
rect 17445 -10 17450 10
rect 17470 -10 17475 10
rect 17445 -20 17475 -10
rect 17505 60 17535 70
rect 17505 40 17510 60
rect 17530 40 17535 60
rect 17505 10 17535 40
rect 17505 -10 17510 10
rect 17530 -10 17535 10
rect 17505 -20 17535 -10
rect 17565 60 17595 70
rect 17565 40 17570 60
rect 17590 40 17595 60
rect 17565 10 17595 40
rect 17565 -10 17570 10
rect 17590 -10 17595 10
rect 17565 -20 17595 -10
rect 17625 60 17695 70
rect 17625 40 17630 60
rect 17650 40 17670 60
rect 17690 40 17695 60
rect 17625 10 17695 40
rect 17625 -10 17630 10
rect 17650 -10 17670 10
rect 17690 -10 17695 10
rect 17625 -20 17695 -10
rect 17905 60 17975 70
rect 17905 40 17910 60
rect 17930 40 17950 60
rect 17970 40 17975 60
rect 17905 10 17975 40
rect 17905 -10 17910 10
rect 17930 -10 17950 10
rect 17970 -10 17975 10
rect 17905 -20 17975 -10
rect 18005 60 18035 70
rect 18005 40 18010 60
rect 18030 40 18035 60
rect 18005 10 18035 40
rect 18005 -10 18010 10
rect 18030 -10 18035 10
rect 18005 -20 18035 -10
rect 18065 60 18095 70
rect 18065 40 18070 60
rect 18090 40 18095 60
rect 18065 10 18095 40
rect 18065 -10 18070 10
rect 18090 -10 18095 10
rect 18065 -20 18095 -10
rect 18125 60 18155 70
rect 18125 40 18130 60
rect 18150 40 18155 60
rect 18125 10 18155 40
rect 18125 -10 18130 10
rect 18150 -10 18155 10
rect 18125 -20 18155 -10
rect 18185 60 18215 70
rect 18185 40 18190 60
rect 18210 40 18215 60
rect 18185 10 18215 40
rect 18185 -10 18190 10
rect 18210 -10 18215 10
rect 18185 -20 18215 -10
rect 18245 60 18275 70
rect 18245 40 18250 60
rect 18270 40 18275 60
rect 18245 10 18275 40
rect 18245 -10 18250 10
rect 18270 -10 18275 10
rect 18245 -20 18275 -10
rect 18305 60 18335 70
rect 18305 40 18310 60
rect 18330 40 18335 60
rect 18305 10 18335 40
rect 18305 -10 18310 10
rect 18330 -10 18335 10
rect 18305 -20 18335 -10
rect 18365 60 18395 70
rect 18365 40 18370 60
rect 18390 40 18395 60
rect 18365 10 18395 40
rect 18365 -10 18370 10
rect 18390 -10 18395 10
rect 18365 -20 18395 -10
rect 18425 60 18455 70
rect 18425 40 18430 60
rect 18450 40 18455 60
rect 18425 10 18455 40
rect 18425 -10 18430 10
rect 18450 -10 18455 10
rect 18425 -20 18455 -10
rect 18485 60 18515 70
rect 18485 40 18490 60
rect 18510 40 18515 60
rect 18485 10 18515 40
rect 18485 -10 18490 10
rect 18510 -10 18515 10
rect 18485 -20 18515 -10
rect 18545 60 18575 70
rect 18545 40 18550 60
rect 18570 40 18575 60
rect 18545 10 18575 40
rect 18545 -10 18550 10
rect 18570 -10 18575 10
rect 18545 -20 18575 -10
rect 18605 60 18635 70
rect 18605 40 18610 60
rect 18630 40 18635 60
rect 18605 10 18635 40
rect 18605 -10 18610 10
rect 18630 -10 18635 10
rect 18605 -20 18635 -10
rect 18665 60 18695 70
rect 18665 40 18670 60
rect 18690 40 18695 60
rect 18665 10 18695 40
rect 18665 -10 18670 10
rect 18690 -10 18695 10
rect 18665 -20 18695 -10
rect 18725 60 18755 70
rect 18725 40 18730 60
rect 18750 40 18755 60
rect 18725 10 18755 40
rect 18725 -10 18730 10
rect 18750 -10 18755 10
rect 18725 -20 18755 -10
rect 18785 60 18815 70
rect 18785 40 18790 60
rect 18810 40 18815 60
rect 18785 10 18815 40
rect 18785 -10 18790 10
rect 18810 -10 18815 10
rect 18785 -20 18815 -10
rect 18845 60 18875 70
rect 18845 40 18850 60
rect 18870 40 18875 60
rect 18845 10 18875 40
rect 18845 -10 18850 10
rect 18870 -10 18875 10
rect 18845 -20 18875 -10
rect 18905 60 18935 70
rect 18905 40 18910 60
rect 18930 40 18935 60
rect 18905 10 18935 40
rect 18905 -10 18910 10
rect 18930 -10 18935 10
rect 18905 -20 18935 -10
rect 18965 60 18995 70
rect 18965 40 18970 60
rect 18990 40 18995 60
rect 18965 10 18995 40
rect 18965 -10 18970 10
rect 18990 -10 18995 10
rect 18965 -20 18995 -10
rect 19025 60 19055 70
rect 19025 40 19030 60
rect 19050 40 19055 60
rect 19025 10 19055 40
rect 19025 -10 19030 10
rect 19050 -10 19055 10
rect 19025 -20 19055 -10
rect 19085 60 19115 70
rect 19085 40 19090 60
rect 19110 40 19115 60
rect 19085 10 19115 40
rect 19085 -10 19090 10
rect 19110 -10 19115 10
rect 19085 -20 19115 -10
rect 19145 60 19215 70
rect 19145 40 19150 60
rect 19170 40 19190 60
rect 19210 40 19215 60
rect 19145 10 19215 40
rect 19145 -10 19150 10
rect 19170 -10 19190 10
rect 19210 -10 19215 10
rect 19145 -20 19215 -10
rect 16425 -50 16455 -20
rect 16610 -40 16630 -20
rect 16730 -40 16750 -20
rect 16970 -40 16990 -20
rect 17090 -40 17110 -20
rect 17330 -40 17350 -20
rect 17450 -40 17470 -20
rect 16425 -70 16430 -50
rect 16450 -70 16455 -50
rect 16425 -80 16455 -70
rect 16510 -50 16550 -40
rect 16510 -70 16520 -50
rect 16540 -70 16550 -50
rect 16510 -80 16550 -70
rect 16600 -50 16640 -40
rect 16600 -70 16610 -50
rect 16630 -70 16640 -50
rect 16600 -80 16640 -70
rect 16720 -50 16760 -40
rect 16720 -70 16730 -50
rect 16750 -70 16760 -50
rect 16720 -80 16760 -70
rect 16840 -50 16880 -40
rect 16840 -70 16850 -50
rect 16870 -70 16880 -50
rect 16840 -80 16880 -70
rect 16960 -50 17000 -40
rect 16960 -70 16970 -50
rect 16990 -70 17000 -50
rect 16960 -80 17000 -70
rect 17080 -50 17120 -40
rect 17080 -70 17090 -50
rect 17110 -70 17120 -50
rect 17080 -80 17120 -70
rect 17200 -50 17240 -40
rect 17200 -70 17210 -50
rect 17230 -70 17240 -50
rect 17200 -80 17240 -70
rect 17320 -50 17360 -40
rect 17320 -70 17330 -50
rect 17350 -70 17360 -50
rect 17320 -80 17360 -70
rect 17440 -50 17480 -40
rect 17440 -70 17450 -50
rect 17470 -70 17480 -50
rect 17440 -80 17480 -70
rect 17535 -50 17565 -40
rect 17535 -70 17540 -50
rect 17560 -70 17565 -50
rect 17535 -80 17565 -70
rect 17945 -50 17975 -20
rect 18130 -40 18150 -20
rect 18250 -40 18270 -20
rect 18490 -40 18510 -20
rect 18610 -40 18630 -20
rect 18850 -40 18870 -20
rect 18970 -40 18990 -20
rect 19145 -25 19180 -20
rect 17945 -70 17950 -50
rect 17970 -70 17975 -50
rect 17945 -80 17975 -70
rect 18035 -50 18065 -40
rect 18035 -70 18040 -50
rect 18060 -70 18065 -50
rect 18035 -80 18065 -70
rect 18120 -50 18160 -40
rect 18120 -70 18130 -50
rect 18150 -70 18160 -50
rect 18120 -80 18160 -70
rect 18240 -50 18280 -40
rect 18240 -70 18250 -50
rect 18270 -70 18280 -50
rect 18240 -80 18280 -70
rect 18360 -50 18400 -40
rect 18360 -70 18370 -50
rect 18390 -70 18400 -50
rect 18360 -80 18400 -70
rect 18480 -50 18520 -40
rect 18480 -70 18490 -50
rect 18510 -70 18520 -50
rect 18480 -80 18520 -70
rect 18600 -50 18640 -40
rect 18600 -70 18610 -50
rect 18630 -70 18640 -50
rect 18600 -80 18640 -70
rect 18720 -50 18760 -40
rect 18720 -70 18730 -50
rect 18750 -70 18760 -50
rect 18720 -80 18760 -70
rect 18840 -50 18880 -40
rect 18840 -70 18850 -50
rect 18870 -70 18880 -50
rect 18840 -80 18880 -70
rect 18960 -50 19000 -40
rect 18960 -70 18970 -50
rect 18990 -70 19000 -50
rect 18960 -80 19000 -70
rect 19050 -50 19090 -40
rect 19050 -70 19060 -50
rect 19080 -70 19090 -50
rect 19050 -80 19090 -70
rect 19145 -50 19175 -25
rect 19145 -70 19150 -50
rect 19170 -70 19175 -50
rect 19145 -80 19175 -70
rect 16910 -210 16950 -200
rect 16910 -230 16920 -210
rect 16940 -230 16950 -210
rect 16910 -240 16950 -230
rect 18650 -210 18690 -205
rect 18650 -230 18660 -210
rect 18680 -230 18690 -210
rect 18650 -240 18690 -230
rect 16850 -255 16890 -245
rect 16850 -275 16860 -255
rect 16880 -275 16890 -255
rect 16850 -285 16890 -275
rect 16975 -255 17005 -245
rect 16975 -275 16980 -255
rect 17000 -275 17005 -255
rect 16975 -285 17005 -275
rect 17090 -255 17130 -245
rect 17090 -275 17100 -255
rect 17120 -275 17130 -255
rect 17090 -285 17130 -275
rect 17215 -255 17245 -245
rect 17215 -275 17220 -255
rect 17240 -275 17245 -255
rect 17215 -285 17245 -275
rect 17330 -255 17370 -245
rect 17330 -275 17340 -255
rect 17360 -275 17370 -255
rect 17330 -285 17370 -275
rect 17455 -255 17485 -245
rect 17455 -275 17460 -255
rect 17480 -275 17485 -255
rect 17455 -285 17485 -275
rect 18115 -255 18145 -245
rect 18115 -275 18120 -255
rect 18140 -275 18145 -255
rect 18115 -285 18145 -275
rect 18230 -255 18270 -245
rect 18230 -275 18240 -255
rect 18260 -275 18270 -255
rect 18230 -285 18270 -275
rect 18355 -255 18385 -245
rect 18355 -275 18360 -255
rect 18380 -275 18385 -255
rect 18355 -285 18385 -275
rect 18470 -255 18510 -245
rect 18470 -275 18480 -255
rect 18500 -275 18510 -255
rect 18470 -285 18510 -275
rect 18595 -255 18625 -245
rect 18595 -275 18600 -255
rect 18620 -275 18625 -255
rect 18595 -285 18625 -275
rect 18710 -255 18750 -245
rect 18710 -275 18720 -255
rect 18740 -275 18750 -255
rect 18710 -285 18750 -275
rect 16860 -305 16880 -285
rect 16980 -305 17000 -285
rect 17100 -305 17120 -285
rect 17220 -305 17240 -285
rect 17340 -305 17360 -285
rect 17460 -305 17480 -285
rect 18120 -305 18140 -285
rect 18240 -305 18260 -285
rect 18360 -305 18380 -285
rect 18480 -305 18500 -285
rect 18600 -305 18620 -285
rect 18720 -305 18740 -285
rect 16855 -315 16885 -305
rect 16855 -335 16860 -315
rect 16880 -335 16885 -315
rect 16855 -345 16885 -335
rect 16915 -315 16945 -305
rect 16915 -335 16920 -315
rect 16940 -335 16945 -315
rect 16915 -345 16945 -335
rect 16975 -315 17005 -305
rect 16975 -335 16980 -315
rect 17000 -335 17005 -315
rect 16975 -345 17005 -335
rect 17035 -315 17065 -305
rect 17035 -335 17040 -315
rect 17060 -335 17065 -315
rect 17035 -345 17065 -335
rect 17095 -315 17125 -305
rect 17095 -335 17100 -315
rect 17120 -335 17125 -315
rect 17095 -345 17125 -335
rect 17155 -315 17185 -305
rect 17155 -335 17160 -315
rect 17180 -335 17185 -315
rect 17155 -345 17185 -335
rect 17215 -315 17245 -305
rect 17215 -335 17220 -315
rect 17240 -335 17245 -315
rect 17215 -345 17245 -335
rect 17275 -315 17305 -305
rect 17275 -335 17280 -315
rect 17300 -335 17305 -315
rect 17275 -345 17305 -335
rect 17335 -315 17365 -305
rect 17335 -335 17340 -315
rect 17360 -335 17365 -315
rect 17335 -345 17365 -335
rect 17395 -315 17425 -305
rect 17395 -335 17400 -315
rect 17420 -335 17425 -315
rect 17395 -345 17425 -335
rect 17455 -315 17485 -305
rect 17455 -335 17460 -315
rect 17480 -335 17485 -315
rect 17455 -345 17485 -335
rect 17565 -315 17595 -305
rect 17565 -335 17570 -315
rect 17590 -335 17595 -315
rect 17565 -345 17595 -335
rect 18005 -315 18035 -305
rect 18005 -335 18010 -315
rect 18030 -335 18035 -315
rect 18005 -345 18035 -335
rect 18115 -315 18145 -305
rect 18115 -335 18120 -315
rect 18140 -335 18145 -315
rect 18115 -345 18145 -335
rect 18175 -315 18205 -305
rect 18175 -335 18180 -315
rect 18200 -335 18205 -315
rect 18175 -345 18205 -335
rect 18235 -315 18265 -305
rect 18235 -335 18240 -315
rect 18260 -335 18265 -315
rect 18235 -345 18265 -335
rect 18295 -315 18325 -305
rect 18295 -335 18300 -315
rect 18320 -335 18325 -315
rect 18295 -345 18325 -335
rect 18355 -315 18385 -305
rect 18355 -335 18360 -315
rect 18380 -335 18385 -315
rect 18355 -345 18385 -335
rect 18415 -315 18445 -305
rect 18415 -335 18420 -315
rect 18440 -335 18445 -315
rect 18415 -345 18445 -335
rect 18475 -315 18505 -305
rect 18475 -335 18480 -315
rect 18500 -335 18505 -315
rect 18475 -345 18505 -335
rect 18535 -315 18565 -305
rect 18535 -335 18540 -315
rect 18560 -335 18565 -315
rect 18535 -345 18565 -335
rect 18595 -315 18625 -305
rect 18595 -335 18600 -315
rect 18620 -335 18625 -315
rect 18595 -345 18625 -335
rect 18655 -315 18685 -305
rect 18655 -335 18660 -315
rect 18680 -335 18685 -315
rect 18655 -345 18685 -335
rect 18715 -315 18745 -305
rect 18715 -335 18720 -315
rect 18740 -335 18745 -315
rect 18715 -345 18745 -335
rect 16920 -365 16940 -345
rect 17040 -365 17060 -345
rect 17160 -365 17180 -345
rect 17280 -365 17300 -345
rect 17400 -365 17420 -345
rect 18180 -365 18200 -345
rect 18300 -365 18320 -345
rect 18420 -365 18440 -345
rect 18540 -365 18560 -345
rect 18660 -365 18680 -345
rect 16850 -375 16890 -365
rect 16850 -395 16860 -375
rect 16880 -395 16890 -375
rect 16850 -405 16890 -395
rect 16915 -375 16945 -365
rect 16915 -395 16920 -375
rect 16940 -395 16945 -375
rect 16915 -405 16945 -395
rect 17035 -375 17065 -365
rect 17035 -395 17040 -375
rect 17060 -395 17065 -375
rect 17035 -405 17065 -395
rect 17155 -375 17185 -365
rect 17155 -395 17160 -375
rect 17180 -395 17185 -375
rect 17155 -405 17185 -395
rect 17275 -375 17305 -365
rect 17275 -395 17280 -375
rect 17300 -395 17305 -375
rect 17275 -405 17305 -395
rect 17395 -375 17425 -365
rect 17395 -395 17400 -375
rect 17420 -395 17425 -375
rect 17395 -405 17425 -395
rect 18175 -375 18205 -365
rect 18175 -395 18180 -375
rect 18200 -395 18205 -375
rect 18175 -405 18205 -395
rect 18295 -375 18325 -365
rect 18295 -395 18300 -375
rect 18320 -395 18325 -375
rect 18295 -405 18325 -395
rect 18415 -375 18445 -365
rect 18415 -395 18420 -375
rect 18440 -395 18445 -375
rect 18415 -405 18445 -395
rect 18535 -375 18565 -365
rect 18535 -395 18540 -375
rect 18560 -395 18565 -375
rect 18535 -405 18565 -395
rect 18655 -375 18685 -365
rect 18655 -395 18660 -375
rect 18680 -395 18685 -375
rect 18655 -405 18685 -395
rect 18710 -375 18750 -365
rect 18710 -395 18720 -375
rect 18740 -395 18750 -375
rect 18710 -405 18750 -395
rect 16620 -535 16660 -530
rect 16530 -550 16570 -540
rect 16530 -570 16540 -550
rect 16560 -570 16570 -550
rect 16620 -555 16630 -535
rect 16650 -555 16660 -535
rect 16620 -565 16660 -555
rect 16740 -535 16780 -530
rect 16740 -555 16750 -535
rect 16770 -555 16780 -535
rect 16740 -565 16780 -555
rect 16860 -535 16900 -530
rect 16860 -555 16870 -535
rect 16890 -555 16900 -535
rect 16860 -565 16900 -555
rect 16980 -535 17020 -530
rect 16980 -555 16990 -535
rect 17010 -555 17020 -535
rect 16980 -565 17020 -555
rect 17300 -535 17340 -530
rect 17300 -555 17310 -535
rect 17330 -555 17340 -535
rect 17300 -565 17340 -555
rect 17420 -535 17460 -530
rect 17420 -555 17430 -535
rect 17450 -555 17460 -535
rect 17420 -565 17460 -555
rect 17540 -535 17580 -530
rect 17540 -555 17550 -535
rect 17570 -555 17580 -535
rect 18020 -535 18060 -525
rect 17540 -565 17580 -555
rect 17690 -550 17730 -540
rect 16530 -580 16570 -570
rect 17690 -570 17700 -550
rect 17720 -570 17730 -550
rect 17690 -580 17730 -570
rect 17870 -550 17910 -540
rect 17870 -570 17880 -550
rect 17900 -570 17910 -550
rect 18020 -555 18030 -535
rect 18050 -555 18060 -535
rect 18020 -565 18060 -555
rect 18140 -535 18180 -525
rect 18140 -555 18150 -535
rect 18170 -555 18180 -535
rect 18140 -565 18180 -555
rect 18260 -535 18300 -525
rect 18260 -555 18270 -535
rect 18290 -555 18300 -535
rect 18260 -565 18300 -555
rect 18580 -535 18620 -525
rect 18580 -555 18590 -535
rect 18610 -555 18620 -535
rect 18580 -565 18620 -555
rect 18700 -535 18740 -525
rect 18700 -555 18710 -535
rect 18730 -555 18740 -535
rect 18700 -565 18740 -555
rect 18820 -535 18860 -525
rect 18820 -555 18830 -535
rect 18850 -555 18860 -535
rect 18820 -565 18860 -555
rect 18940 -535 18980 -525
rect 18940 -555 18950 -535
rect 18970 -555 18980 -535
rect 18940 -565 18980 -555
rect 19030 -550 19070 -540
rect 17870 -580 17910 -570
rect 19030 -570 19040 -550
rect 19060 -570 19070 -550
rect 19030 -580 19070 -570
rect 16535 -590 16565 -580
rect 16535 -610 16540 -590
rect 16560 -610 16565 -590
rect 16535 -640 16565 -610
rect 16535 -660 16540 -640
rect 16560 -660 16565 -640
rect 16535 -690 16565 -660
rect 16535 -710 16540 -690
rect 16560 -710 16565 -690
rect 16535 -740 16565 -710
rect 16535 -760 16540 -740
rect 16560 -760 16565 -740
rect 16535 -790 16565 -760
rect 16535 -810 16540 -790
rect 16560 -810 16565 -790
rect 16535 -820 16565 -810
rect 17075 -590 17185 -580
rect 17075 -610 17080 -590
rect 17100 -610 17120 -590
rect 17140 -610 17160 -590
rect 17180 -610 17185 -590
rect 17075 -640 17185 -610
rect 17075 -660 17080 -640
rect 17100 -660 17120 -640
rect 17140 -660 17160 -640
rect 17180 -660 17185 -640
rect 17075 -690 17185 -660
rect 17075 -710 17080 -690
rect 17100 -710 17120 -690
rect 17140 -710 17160 -690
rect 17180 -710 17185 -690
rect 17075 -740 17185 -710
rect 17075 -760 17080 -740
rect 17100 -760 17120 -740
rect 17140 -760 17160 -740
rect 17180 -760 17185 -740
rect 17075 -790 17185 -760
rect 17075 -810 17080 -790
rect 17100 -810 17120 -790
rect 17140 -810 17160 -790
rect 17180 -810 17185 -790
rect 17075 -820 17185 -810
rect 17695 -590 17725 -580
rect 17695 -610 17700 -590
rect 17720 -610 17725 -590
rect 17695 -640 17725 -610
rect 17695 -660 17700 -640
rect 17720 -660 17725 -640
rect 17695 -690 17725 -660
rect 17695 -710 17700 -690
rect 17720 -710 17725 -690
rect 17695 -740 17725 -710
rect 17695 -760 17700 -740
rect 17720 -760 17725 -740
rect 17695 -790 17725 -760
rect 17695 -810 17700 -790
rect 17720 -810 17725 -790
rect 17695 -820 17725 -810
rect 17875 -590 17905 -580
rect 17875 -610 17880 -590
rect 17900 -610 17905 -590
rect 17875 -640 17905 -610
rect 17875 -660 17880 -640
rect 17900 -660 17905 -640
rect 17875 -690 17905 -660
rect 17875 -710 17880 -690
rect 17900 -710 17905 -690
rect 17875 -740 17905 -710
rect 17875 -760 17880 -740
rect 17900 -760 17905 -740
rect 17875 -790 17905 -760
rect 17875 -810 17880 -790
rect 17900 -810 17905 -790
rect 17875 -820 17905 -810
rect 18415 -590 18525 -580
rect 18415 -610 18420 -590
rect 18440 -610 18460 -590
rect 18480 -610 18500 -590
rect 18520 -610 18525 -590
rect 18415 -640 18525 -610
rect 18415 -660 18420 -640
rect 18440 -660 18460 -640
rect 18480 -660 18500 -640
rect 18520 -660 18525 -640
rect 18415 -690 18525 -660
rect 18415 -710 18420 -690
rect 18440 -710 18460 -690
rect 18480 -710 18500 -690
rect 18520 -710 18525 -690
rect 18415 -740 18525 -710
rect 18415 -760 18420 -740
rect 18440 -760 18460 -740
rect 18480 -760 18500 -740
rect 18520 -760 18525 -740
rect 18415 -790 18525 -760
rect 18415 -810 18420 -790
rect 18440 -810 18460 -790
rect 18480 -810 18500 -790
rect 18520 -810 18525 -790
rect 18415 -820 18525 -810
rect 19035 -590 19065 -580
rect 19035 -610 19040 -590
rect 19060 -610 19065 -590
rect 19035 -640 19065 -610
rect 19035 -660 19040 -640
rect 19060 -660 19065 -640
rect 19035 -690 19065 -660
rect 19035 -710 19040 -690
rect 19060 -710 19065 -690
rect 19035 -740 19065 -710
rect 19035 -760 19040 -740
rect 19060 -760 19065 -740
rect 19035 -790 19065 -760
rect 19035 -810 19040 -790
rect 19060 -810 19065 -790
rect 19035 -820 19065 -810
rect 17120 -840 17140 -820
rect 18460 -840 18480 -820
rect 17110 -850 17150 -840
rect 17110 -870 17120 -850
rect 17140 -870 17150 -850
rect 17110 -880 17150 -870
rect 18450 -850 18490 -840
rect 18450 -870 18460 -850
rect 18480 -870 18490 -850
rect 18450 -880 18490 -870
rect 16740 -1000 16780 -990
rect 16740 -1020 16750 -1000
rect 16770 -1020 16780 -1000
rect 16740 -1030 16780 -1020
rect 16820 -1000 16860 -990
rect 16820 -1020 16830 -1000
rect 16850 -1020 16860 -1000
rect 16820 -1030 16860 -1020
rect 16900 -1000 16940 -990
rect 16900 -1020 16910 -1000
rect 16930 -1020 16940 -1000
rect 16900 -1030 16940 -1020
rect 16980 -1000 17020 -990
rect 16980 -1020 16990 -1000
rect 17010 -1020 17020 -1000
rect 16980 -1030 17020 -1020
rect 17060 -1000 17100 -990
rect 17060 -1020 17070 -1000
rect 17090 -1020 17100 -1000
rect 17060 -1030 17100 -1020
rect 17140 -1000 17180 -990
rect 17140 -1020 17150 -1000
rect 17170 -1020 17180 -1000
rect 17140 -1030 17180 -1020
rect 17220 -1000 17260 -990
rect 17220 -1020 17230 -1000
rect 17250 -1020 17260 -1000
rect 17220 -1030 17260 -1020
rect 17300 -1000 17340 -990
rect 17300 -1020 17310 -1000
rect 17330 -1020 17340 -1000
rect 17300 -1030 17340 -1020
rect 17380 -1000 17420 -990
rect 17380 -1020 17390 -1000
rect 17410 -1020 17420 -1000
rect 17380 -1030 17420 -1020
rect 17460 -1000 17500 -990
rect 17460 -1020 17470 -1000
rect 17490 -1020 17500 -1000
rect 17460 -1030 17500 -1020
rect 17540 -1000 17580 -990
rect 17540 -1020 17550 -1000
rect 17570 -1020 17580 -1000
rect 17540 -1030 17580 -1020
rect 17620 -1000 17660 -990
rect 17620 -1020 17630 -1000
rect 17650 -1020 17660 -1000
rect 17620 -1030 17660 -1020
rect 17700 -1000 17740 -990
rect 17700 -1020 17710 -1000
rect 17730 -1020 17740 -1000
rect 17700 -1030 17740 -1020
rect 17780 -1000 17820 -990
rect 17780 -1020 17790 -1000
rect 17810 -1020 17820 -1000
rect 17780 -1030 17820 -1020
rect 17860 -1000 17900 -990
rect 17860 -1020 17870 -1000
rect 17890 -1020 17900 -1000
rect 17860 -1030 17900 -1020
rect 17940 -1000 17980 -990
rect 17940 -1020 17950 -1000
rect 17970 -1020 17980 -1000
rect 17940 -1030 17980 -1020
rect 18020 -1000 18060 -990
rect 18020 -1020 18030 -1000
rect 18050 -1020 18060 -1000
rect 18020 -1030 18060 -1020
rect 18100 -1000 18140 -990
rect 18100 -1020 18110 -1000
rect 18130 -1020 18140 -1000
rect 18100 -1030 18140 -1020
rect 18180 -1000 18220 -990
rect 18180 -1020 18190 -1000
rect 18210 -1020 18220 -1000
rect 18180 -1030 18220 -1020
rect 18260 -1000 18300 -990
rect 18260 -1020 18270 -1000
rect 18290 -1020 18300 -1000
rect 18260 -1030 18300 -1020
rect 18340 -1000 18380 -990
rect 18340 -1020 18350 -1000
rect 18370 -1020 18380 -1000
rect 18340 -1030 18380 -1020
rect 18420 -1000 18460 -990
rect 18420 -1020 18430 -1000
rect 18450 -1020 18460 -1000
rect 18420 -1030 18460 -1020
rect 18500 -1000 18540 -990
rect 18500 -1020 18510 -1000
rect 18530 -1020 18540 -1000
rect 18500 -1030 18540 -1020
rect 18580 -1000 18620 -990
rect 18580 -1020 18590 -1000
rect 18610 -1020 18620 -1000
rect 18580 -1030 18620 -1020
rect 18660 -1000 18700 -990
rect 18660 -1020 18670 -1000
rect 18690 -1020 18700 -1000
rect 18660 -1030 18700 -1020
rect 18740 -1000 18780 -990
rect 18740 -1020 18750 -1000
rect 18770 -1020 18780 -1000
rect 18740 -1030 18780 -1020
rect 16750 -1050 16770 -1030
rect 17790 -1050 17810 -1030
rect 16745 -1060 16775 -1050
rect 16745 -1075 16750 -1060
rect 16700 -1080 16750 -1075
rect 16770 -1080 16775 -1060
rect 16700 -1085 16775 -1080
rect 16700 -1105 16710 -1085
rect 16730 -1105 16775 -1085
rect 16700 -1110 16775 -1105
rect 16700 -1115 16750 -1110
rect 16745 -1130 16750 -1115
rect 16770 -1130 16775 -1110
rect 16745 -1140 16775 -1130
rect 17785 -1060 17815 -1050
rect 17785 -1080 17790 -1060
rect 17810 -1080 17815 -1060
rect 17785 -1110 17815 -1080
rect 17785 -1130 17790 -1110
rect 17810 -1130 17815 -1110
rect 17785 -1140 17815 -1130
rect 18825 -1060 18895 -1050
rect 18825 -1080 18830 -1060
rect 18850 -1080 18870 -1060
rect 18890 -1075 18895 -1060
rect 18890 -1080 18935 -1075
rect 18825 -1085 18935 -1080
rect 18825 -1105 18905 -1085
rect 18925 -1105 18935 -1085
rect 18825 -1110 18935 -1105
rect 18825 -1130 18830 -1110
rect 18850 -1130 18870 -1110
rect 18890 -1115 18935 -1110
rect 18890 -1130 18895 -1115
rect 18825 -1140 18895 -1130
rect 16890 -1275 16930 -1265
rect 16890 -1295 16900 -1275
rect 16920 -1295 16930 -1275
rect 16890 -1305 16930 -1295
rect 17000 -1275 17040 -1265
rect 17000 -1295 17010 -1275
rect 17030 -1295 17040 -1275
rect 17000 -1305 17040 -1295
rect 17110 -1275 17150 -1265
rect 17110 -1295 17120 -1275
rect 17140 -1295 17150 -1275
rect 17110 -1305 17150 -1295
rect 17170 -1275 17200 -1265
rect 17170 -1295 17175 -1275
rect 17195 -1295 17200 -1275
rect 17170 -1305 17200 -1295
rect 17220 -1275 17260 -1265
rect 17220 -1295 17230 -1275
rect 17250 -1295 17260 -1275
rect 17220 -1305 17260 -1295
rect 17330 -1275 17370 -1265
rect 17330 -1295 17340 -1275
rect 17360 -1295 17370 -1275
rect 17330 -1305 17370 -1295
rect 17505 -1275 17545 -1265
rect 17505 -1295 17515 -1275
rect 17535 -1295 17545 -1275
rect 17505 -1305 17545 -1295
rect 17615 -1275 17655 -1265
rect 17615 -1295 17625 -1275
rect 17645 -1295 17655 -1275
rect 17615 -1305 17655 -1295
rect 17725 -1275 17765 -1265
rect 17725 -1295 17735 -1275
rect 17755 -1295 17765 -1275
rect 17725 -1305 17765 -1295
rect 17785 -1275 17815 -1265
rect 17785 -1295 17790 -1275
rect 17810 -1295 17815 -1275
rect 17785 -1305 17815 -1295
rect 17835 -1275 17875 -1265
rect 17835 -1295 17845 -1275
rect 17865 -1295 17875 -1275
rect 17835 -1305 17875 -1295
rect 17945 -1275 17985 -1265
rect 17945 -1295 17955 -1275
rect 17975 -1295 17985 -1275
rect 17945 -1305 17985 -1295
rect 18055 -1275 18095 -1265
rect 18055 -1295 18065 -1275
rect 18085 -1295 18095 -1275
rect 18055 -1305 18095 -1295
rect 18230 -1275 18270 -1265
rect 18230 -1295 18240 -1275
rect 18260 -1295 18270 -1275
rect 18230 -1305 18270 -1295
rect 18340 -1275 18380 -1265
rect 18340 -1295 18350 -1275
rect 18370 -1295 18380 -1275
rect 18340 -1305 18380 -1295
rect 18400 -1275 18430 -1265
rect 18400 -1295 18405 -1275
rect 18425 -1295 18430 -1275
rect 18400 -1305 18430 -1295
rect 18450 -1275 18490 -1265
rect 18450 -1295 18460 -1275
rect 18480 -1295 18490 -1275
rect 18450 -1305 18490 -1295
rect 18560 -1275 18600 -1265
rect 18560 -1295 18570 -1275
rect 18590 -1295 18600 -1275
rect 18560 -1305 18600 -1295
rect 18670 -1275 18710 -1265
rect 18670 -1295 18680 -1275
rect 18700 -1295 18710 -1275
rect 18670 -1305 18710 -1295
rect 16895 -1325 16925 -1305
rect 17010 -1325 17030 -1305
rect 17120 -1325 17140 -1305
rect 17230 -1325 17250 -1305
rect 17335 -1325 17365 -1305
rect 17510 -1325 17540 -1305
rect 17625 -1325 17645 -1305
rect 17735 -1325 17755 -1305
rect 17845 -1325 17865 -1305
rect 17955 -1325 17975 -1305
rect 18060 -1325 18090 -1305
rect 18235 -1325 18265 -1305
rect 18350 -1325 18370 -1305
rect 18460 -1325 18480 -1305
rect 18570 -1325 18590 -1305
rect 18675 -1325 18705 -1305
rect 16855 -1335 16925 -1325
rect 16855 -1355 16860 -1335
rect 16880 -1355 16900 -1335
rect 16920 -1355 16925 -1335
rect 16855 -1385 16925 -1355
rect 16855 -1405 16860 -1385
rect 16880 -1405 16900 -1385
rect 16920 -1405 16925 -1385
rect 16855 -1415 16925 -1405
rect 16950 -1335 16980 -1325
rect 16950 -1355 16955 -1335
rect 16975 -1355 16980 -1335
rect 16950 -1385 16980 -1355
rect 16950 -1405 16955 -1385
rect 16975 -1405 16980 -1385
rect 16950 -1415 16980 -1405
rect 17005 -1335 17035 -1325
rect 17005 -1355 17010 -1335
rect 17030 -1355 17035 -1335
rect 17005 -1385 17035 -1355
rect 17005 -1405 17010 -1385
rect 17030 -1405 17035 -1385
rect 17005 -1415 17035 -1405
rect 17060 -1335 17090 -1325
rect 17060 -1355 17065 -1335
rect 17085 -1355 17090 -1335
rect 17060 -1385 17090 -1355
rect 17060 -1405 17065 -1385
rect 17085 -1405 17090 -1385
rect 17060 -1415 17090 -1405
rect 17115 -1335 17145 -1325
rect 17115 -1355 17120 -1335
rect 17140 -1355 17145 -1335
rect 17115 -1385 17145 -1355
rect 17115 -1405 17120 -1385
rect 17140 -1405 17145 -1385
rect 17115 -1415 17145 -1405
rect 17170 -1335 17200 -1325
rect 17170 -1355 17175 -1335
rect 17195 -1355 17200 -1335
rect 17170 -1385 17200 -1355
rect 17170 -1405 17175 -1385
rect 17195 -1405 17200 -1385
rect 17170 -1415 17200 -1405
rect 17225 -1335 17255 -1325
rect 17225 -1355 17230 -1335
rect 17250 -1355 17255 -1335
rect 17225 -1385 17255 -1355
rect 17225 -1405 17230 -1385
rect 17250 -1405 17255 -1385
rect 17225 -1415 17255 -1405
rect 17280 -1335 17310 -1325
rect 17280 -1355 17285 -1335
rect 17305 -1355 17310 -1335
rect 17280 -1385 17310 -1355
rect 17280 -1405 17285 -1385
rect 17305 -1405 17310 -1385
rect 17280 -1415 17310 -1405
rect 17335 -1335 17405 -1325
rect 17335 -1355 17340 -1335
rect 17360 -1355 17380 -1335
rect 17400 -1355 17405 -1335
rect 17335 -1385 17405 -1355
rect 17335 -1405 17340 -1385
rect 17360 -1405 17380 -1385
rect 17400 -1405 17405 -1385
rect 17335 -1415 17405 -1405
rect 17470 -1335 17540 -1325
rect 17470 -1355 17475 -1335
rect 17495 -1355 17515 -1335
rect 17535 -1355 17540 -1335
rect 17470 -1385 17540 -1355
rect 17470 -1405 17475 -1385
rect 17495 -1405 17515 -1385
rect 17535 -1405 17540 -1385
rect 17470 -1415 17540 -1405
rect 17565 -1335 17595 -1325
rect 17565 -1355 17570 -1335
rect 17590 -1355 17595 -1335
rect 17565 -1385 17595 -1355
rect 17565 -1405 17570 -1385
rect 17590 -1405 17595 -1385
rect 17565 -1415 17595 -1405
rect 17620 -1335 17650 -1325
rect 17620 -1355 17625 -1335
rect 17645 -1355 17650 -1335
rect 17620 -1385 17650 -1355
rect 17620 -1405 17625 -1385
rect 17645 -1405 17650 -1385
rect 17620 -1415 17650 -1405
rect 17675 -1335 17705 -1325
rect 17675 -1355 17680 -1335
rect 17700 -1355 17705 -1335
rect 17675 -1385 17705 -1355
rect 17675 -1405 17680 -1385
rect 17700 -1405 17705 -1385
rect 17675 -1415 17705 -1405
rect 17730 -1335 17760 -1325
rect 17730 -1355 17735 -1335
rect 17755 -1355 17760 -1335
rect 17730 -1385 17760 -1355
rect 17730 -1405 17735 -1385
rect 17755 -1405 17760 -1385
rect 17730 -1415 17760 -1405
rect 17785 -1335 17815 -1325
rect 17785 -1355 17790 -1335
rect 17810 -1355 17815 -1335
rect 17785 -1385 17815 -1355
rect 17785 -1405 17790 -1385
rect 17810 -1405 17815 -1385
rect 17785 -1415 17815 -1405
rect 17840 -1335 17870 -1325
rect 17840 -1355 17845 -1335
rect 17865 -1355 17870 -1335
rect 17840 -1385 17870 -1355
rect 17840 -1405 17845 -1385
rect 17865 -1405 17870 -1385
rect 17840 -1415 17870 -1405
rect 17895 -1335 17925 -1325
rect 17895 -1355 17900 -1335
rect 17920 -1355 17925 -1335
rect 17895 -1385 17925 -1355
rect 17895 -1405 17900 -1385
rect 17920 -1405 17925 -1385
rect 17895 -1415 17925 -1405
rect 17950 -1335 17980 -1325
rect 17950 -1355 17955 -1335
rect 17975 -1355 17980 -1335
rect 17950 -1385 17980 -1355
rect 17950 -1405 17955 -1385
rect 17975 -1405 17980 -1385
rect 17950 -1415 17980 -1405
rect 18005 -1335 18035 -1325
rect 18005 -1355 18010 -1335
rect 18030 -1355 18035 -1335
rect 18005 -1385 18035 -1355
rect 18005 -1405 18010 -1385
rect 18030 -1405 18035 -1385
rect 18005 -1415 18035 -1405
rect 18060 -1335 18130 -1325
rect 18060 -1355 18065 -1335
rect 18085 -1355 18105 -1335
rect 18125 -1355 18130 -1335
rect 18060 -1385 18130 -1355
rect 18060 -1405 18065 -1385
rect 18085 -1405 18105 -1385
rect 18125 -1405 18130 -1385
rect 18060 -1415 18130 -1405
rect 18195 -1335 18265 -1325
rect 18195 -1355 18200 -1335
rect 18220 -1355 18240 -1335
rect 18260 -1355 18265 -1335
rect 18195 -1385 18265 -1355
rect 18195 -1405 18200 -1385
rect 18220 -1405 18240 -1385
rect 18260 -1405 18265 -1385
rect 18195 -1415 18265 -1405
rect 18290 -1335 18320 -1325
rect 18290 -1355 18295 -1335
rect 18315 -1355 18320 -1335
rect 18290 -1385 18320 -1355
rect 18290 -1405 18295 -1385
rect 18315 -1405 18320 -1385
rect 18290 -1415 18320 -1405
rect 18345 -1335 18375 -1325
rect 18345 -1355 18350 -1335
rect 18370 -1355 18375 -1335
rect 18345 -1385 18375 -1355
rect 18345 -1405 18350 -1385
rect 18370 -1405 18375 -1385
rect 18345 -1415 18375 -1405
rect 18400 -1335 18430 -1325
rect 18400 -1355 18405 -1335
rect 18425 -1355 18430 -1335
rect 18400 -1385 18430 -1355
rect 18400 -1405 18405 -1385
rect 18425 -1405 18430 -1385
rect 18400 -1415 18430 -1405
rect 18455 -1335 18485 -1325
rect 18455 -1355 18460 -1335
rect 18480 -1355 18485 -1335
rect 18455 -1385 18485 -1355
rect 18455 -1405 18460 -1385
rect 18480 -1405 18485 -1385
rect 18455 -1415 18485 -1405
rect 18510 -1335 18540 -1325
rect 18510 -1355 18515 -1335
rect 18535 -1355 18540 -1335
rect 18510 -1385 18540 -1355
rect 18510 -1405 18515 -1385
rect 18535 -1405 18540 -1385
rect 18510 -1415 18540 -1405
rect 18565 -1335 18595 -1325
rect 18565 -1355 18570 -1335
rect 18590 -1355 18595 -1335
rect 18565 -1385 18595 -1355
rect 18565 -1405 18570 -1385
rect 18590 -1405 18595 -1385
rect 18565 -1415 18595 -1405
rect 18620 -1335 18650 -1325
rect 18620 -1355 18625 -1335
rect 18645 -1355 18650 -1335
rect 18620 -1385 18650 -1355
rect 18620 -1405 18625 -1385
rect 18645 -1405 18650 -1385
rect 18620 -1415 18650 -1405
rect 18675 -1335 18745 -1325
rect 18675 -1355 18680 -1335
rect 18700 -1355 18720 -1335
rect 18740 -1355 18745 -1335
rect 18675 -1385 18745 -1355
rect 18675 -1405 18680 -1385
rect 18700 -1405 18720 -1385
rect 18740 -1405 18745 -1385
rect 18675 -1415 18745 -1405
rect 16955 -1435 16975 -1415
rect 17065 -1435 17085 -1415
rect 17175 -1435 17195 -1415
rect 17285 -1435 17305 -1415
rect 17570 -1435 17590 -1415
rect 17680 -1435 17700 -1415
rect 17790 -1435 17810 -1415
rect 17900 -1435 17920 -1415
rect 18010 -1435 18030 -1415
rect 18295 -1435 18315 -1415
rect 18405 -1435 18425 -1415
rect 18515 -1435 18535 -1415
rect 18625 -1435 18645 -1415
rect 16945 -1445 16985 -1435
rect 16945 -1465 16955 -1445
rect 16975 -1465 16985 -1445
rect 16945 -1475 16985 -1465
rect 17055 -1445 17095 -1435
rect 17055 -1465 17065 -1445
rect 17085 -1465 17095 -1445
rect 17055 -1475 17095 -1465
rect 17165 -1445 17205 -1435
rect 17165 -1465 17175 -1445
rect 17195 -1465 17205 -1445
rect 17165 -1475 17205 -1465
rect 17275 -1445 17315 -1435
rect 17275 -1465 17285 -1445
rect 17305 -1465 17315 -1445
rect 17275 -1475 17315 -1465
rect 17570 -1445 17625 -1435
rect 17570 -1465 17595 -1445
rect 17615 -1465 17625 -1445
rect 17570 -1475 17625 -1465
rect 17670 -1445 17710 -1435
rect 17670 -1465 17680 -1445
rect 17700 -1465 17710 -1445
rect 17670 -1475 17710 -1465
rect 17780 -1445 17820 -1435
rect 17780 -1465 17790 -1445
rect 17810 -1465 17820 -1445
rect 17780 -1475 17820 -1465
rect 17890 -1445 17930 -1435
rect 17890 -1465 17900 -1445
rect 17920 -1465 17930 -1445
rect 17890 -1475 17930 -1465
rect 18000 -1445 18040 -1435
rect 18000 -1465 18010 -1445
rect 18030 -1465 18040 -1445
rect 18000 -1475 18040 -1465
rect 18285 -1445 18325 -1435
rect 18285 -1465 18295 -1445
rect 18315 -1465 18325 -1445
rect 18285 -1475 18325 -1465
rect 18395 -1445 18435 -1435
rect 18395 -1465 18405 -1445
rect 18425 -1465 18435 -1445
rect 18395 -1475 18435 -1465
rect 18505 -1445 18545 -1435
rect 18505 -1465 18515 -1445
rect 18535 -1465 18545 -1445
rect 18505 -1475 18545 -1465
rect 18615 -1445 18655 -1435
rect 18615 -1465 18625 -1445
rect 18645 -1465 18655 -1445
rect 18615 -1475 18655 -1465
rect 17425 -1900 17470 -1895
rect 17425 -1925 17435 -1900
rect 17460 -1925 17470 -1900
rect 17425 -1930 17470 -1925
rect 18124 -1900 18169 -1895
rect 18124 -1925 18134 -1900
rect 18159 -1925 18169 -1900
rect 18124 -1930 18169 -1925
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3111
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -2997 19440 -2987
rect 19405 -3022 19410 -2997
rect 19435 -3022 19440 -2997
rect 19405 -3032 19440 -3022
rect 19320 -3067 19345 -3032
rect 19610 -3121 19645 -3111
rect 19610 -3146 19615 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3156 19645 -3146
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4170 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4190 17790 -4170
rect 17810 -4190 17820 -4170
rect 17780 -4220 17820 -4190
rect 17780 -4240 17790 -4220
rect 17810 -4240 17820 -4220
rect 17780 -4270 17820 -4240
rect 17780 -4290 17790 -4270
rect 17810 -4290 17820 -4270
rect 17780 -4300 17820 -4290
<< viali >>
rect 16250 1255 16270 1275
rect 16345 1255 16365 1275
rect 16399 1255 16419 1275
rect 16470 1255 16490 1275
rect 16820 1255 16840 1275
rect 16930 1255 16950 1275
rect 16985 1255 17005 1275
rect 17040 1255 17060 1275
rect 17095 1255 17115 1275
rect 17150 1255 17170 1275
rect 17615 1255 17635 1275
rect 17680 1255 17700 1275
rect 17735 1255 17755 1275
rect 17790 1255 17810 1275
rect 17845 1255 17865 1275
rect 17900 1255 17920 1275
rect 17965 1255 17985 1275
rect 18430 1255 18450 1275
rect 18485 1255 18505 1275
rect 18540 1255 18560 1275
rect 18595 1255 18615 1275
rect 18650 1255 18670 1275
rect 18760 1255 18780 1275
rect 16305 1085 16325 1105
rect 16415 1085 16435 1105
rect 16875 1085 16895 1105
rect 16985 1085 17005 1105
rect 17095 1085 17115 1105
rect 18485 1085 18505 1105
rect 18595 1085 18615 1105
rect 18705 1085 18725 1105
rect 17735 985 17755 1005
rect 17845 985 17865 1005
rect 16980 790 17000 810
rect 17160 790 17180 810
rect 17340 790 17360 810
rect 17520 790 17540 810
rect 17700 790 17720 810
rect 17880 790 17900 810
rect 18060 790 18080 810
rect 18240 790 18260 810
rect 18420 790 18440 810
rect 18600 790 18620 810
rect 16445 690 16465 710
rect 16555 690 16575 710
rect 16665 690 16685 710
rect 16490 520 16510 540
rect 16555 520 16575 540
rect 16620 520 16640 540
rect 18955 740 18975 760
rect 19020 740 19040 760
rect 19130 740 19150 760
rect 19036 470 19056 490
rect 19090 470 19110 490
rect 17070 420 17090 440
rect 17250 420 17270 440
rect 17430 420 17450 440
rect 17610 420 17630 440
rect 17700 420 17720 440
rect 17790 420 17810 440
rect 17970 420 17990 440
rect 18150 420 18170 440
rect 18330 420 18350 440
rect 18420 420 18440 440
rect 18510 420 18530 440
rect 16430 100 16450 120
rect 16490 100 16510 120
rect 16550 100 16570 120
rect 16670 100 16690 120
rect 16790 100 16810 120
rect 16850 100 16870 120
rect 16910 100 16930 120
rect 17030 100 17050 120
rect 17150 100 17170 120
rect 17210 100 17230 120
rect 17270 100 17290 120
rect 17390 100 17410 120
rect 17510 100 17530 120
rect 17570 100 17590 120
rect 17630 100 17650 120
rect 17950 100 17970 120
rect 18010 100 18030 120
rect 18070 100 18090 120
rect 18190 100 18210 120
rect 18310 100 18330 120
rect 18370 100 18390 120
rect 18430 100 18450 120
rect 18550 100 18570 120
rect 18670 100 18690 120
rect 18730 100 18750 120
rect 18790 100 18810 120
rect 18910 100 18930 120
rect 19030 100 19050 120
rect 19090 100 19110 120
rect 19150 100 19170 120
rect 16520 -70 16540 -50
rect 16610 -70 16630 -50
rect 16730 -70 16750 -50
rect 16850 -70 16870 -50
rect 16970 -70 16990 -50
rect 17090 -70 17110 -50
rect 17210 -70 17230 -50
rect 17330 -70 17350 -50
rect 17450 -70 17470 -50
rect 17540 -70 17560 -50
rect 18040 -70 18060 -50
rect 18130 -70 18150 -50
rect 18250 -70 18270 -50
rect 18370 -70 18390 -50
rect 18490 -70 18510 -50
rect 18610 -70 18630 -50
rect 18730 -70 18750 -50
rect 18850 -70 18870 -50
rect 18970 -70 18990 -50
rect 19060 -70 19080 -50
rect 16920 -230 16940 -210
rect 18660 -230 18680 -210
rect 16860 -275 16880 -255
rect 16980 -275 17000 -255
rect 17100 -275 17120 -255
rect 17220 -275 17240 -255
rect 17340 -275 17360 -255
rect 17460 -275 17480 -255
rect 18120 -275 18140 -255
rect 18240 -275 18260 -255
rect 18360 -275 18380 -255
rect 18480 -275 18500 -255
rect 18600 -275 18620 -255
rect 18720 -275 18740 -255
rect 17570 -335 17590 -315
rect 18010 -335 18030 -315
rect 16860 -395 16880 -375
rect 16920 -395 16940 -375
rect 17040 -395 17060 -375
rect 17160 -395 17180 -375
rect 17280 -395 17300 -375
rect 17400 -395 17420 -375
rect 18180 -395 18200 -375
rect 18300 -395 18320 -375
rect 18420 -395 18440 -375
rect 18540 -395 18560 -375
rect 18660 -395 18680 -375
rect 18720 -395 18740 -375
rect 16540 -570 16560 -550
rect 16630 -555 16650 -535
rect 16750 -555 16770 -535
rect 16870 -555 16890 -535
rect 16990 -555 17010 -535
rect 17310 -555 17330 -535
rect 17430 -555 17450 -535
rect 17550 -555 17570 -535
rect 17700 -570 17720 -550
rect 17880 -570 17900 -550
rect 18030 -555 18050 -535
rect 18150 -555 18170 -535
rect 18270 -555 18290 -535
rect 18590 -555 18610 -535
rect 18710 -555 18730 -535
rect 18830 -555 18850 -535
rect 18950 -555 18970 -535
rect 19040 -570 19060 -550
rect 17120 -870 17140 -850
rect 18460 -870 18480 -850
rect 16750 -1020 16770 -1000
rect 16830 -1020 16850 -1000
rect 16910 -1020 16930 -1000
rect 16990 -1020 17010 -1000
rect 17070 -1020 17090 -1000
rect 17150 -1020 17170 -1000
rect 17230 -1020 17250 -1000
rect 17310 -1020 17330 -1000
rect 17390 -1020 17410 -1000
rect 17470 -1020 17490 -1000
rect 17550 -1020 17570 -1000
rect 17630 -1020 17650 -1000
rect 17710 -1020 17730 -1000
rect 17790 -1020 17810 -1000
rect 17870 -1020 17890 -1000
rect 17950 -1020 17970 -1000
rect 18030 -1020 18050 -1000
rect 18110 -1020 18130 -1000
rect 18190 -1020 18210 -1000
rect 18270 -1020 18290 -1000
rect 18350 -1020 18370 -1000
rect 18430 -1020 18450 -1000
rect 18510 -1020 18530 -1000
rect 18590 -1020 18610 -1000
rect 18670 -1020 18690 -1000
rect 18750 -1020 18770 -1000
rect 16710 -1105 16730 -1085
rect 18905 -1105 18925 -1085
rect 16900 -1295 16920 -1275
rect 17010 -1295 17030 -1275
rect 17120 -1295 17140 -1275
rect 17175 -1295 17195 -1275
rect 17230 -1295 17250 -1275
rect 17340 -1295 17360 -1275
rect 17515 -1295 17535 -1275
rect 17625 -1295 17645 -1275
rect 17735 -1295 17755 -1275
rect 17790 -1295 17810 -1275
rect 17845 -1295 17865 -1275
rect 17955 -1295 17975 -1275
rect 18065 -1295 18085 -1275
rect 18240 -1295 18260 -1275
rect 18350 -1295 18370 -1275
rect 18405 -1295 18425 -1275
rect 18460 -1295 18480 -1275
rect 18570 -1295 18590 -1275
rect 18680 -1295 18700 -1275
rect 16955 -1465 16975 -1445
rect 17065 -1465 17085 -1445
rect 17175 -1465 17195 -1445
rect 17285 -1465 17305 -1445
rect 17595 -1465 17615 -1445
rect 17680 -1465 17700 -1445
rect 17790 -1465 17810 -1445
rect 17900 -1465 17920 -1445
rect 18010 -1465 18030 -1445
rect 18295 -1465 18315 -1445
rect 18405 -1465 18425 -1445
rect 18515 -1465 18535 -1445
rect 18625 -1465 18645 -1445
rect 17435 -1925 17460 -1900
rect 18134 -1925 18159 -1900
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3022 19435 -2997
rect 19615 -3146 19640 -3121
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4290 17810 -4270
<< metal1 >>
rect 15725 -105 15765 -100
rect 15725 -135 15730 -105
rect 15760 -135 15765 -105
rect 15725 -140 15765 -135
rect 15735 -4310 15755 -140
rect 15795 -1585 15815 1595
rect 15950 125 15990 130
rect 15950 95 15955 125
rect 15985 95 15990 125
rect 15950 90 15990 95
rect 15785 -1590 15825 -1585
rect 15785 -1620 15790 -1590
rect 15820 -1620 15825 -1590
rect 15785 -1625 15825 -1620
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 90
rect 16040 -1540 16060 1595
rect 16030 -1545 16070 -1540
rect 16030 -1575 16035 -1545
rect 16065 -1575 16070 -1545
rect 16030 -1580 16070 -1575
rect 16115 -1680 16135 1595
rect 17095 1390 17115 1595
rect 17085 1385 17125 1390
rect 17085 1355 17090 1385
rect 17120 1355 17125 1385
rect 17085 1350 17125 1355
rect 16390 1340 16430 1345
rect 16390 1310 16395 1340
rect 16425 1310 16430 1340
rect 16390 1305 16430 1310
rect 16975 1340 17015 1345
rect 16975 1310 16980 1340
rect 17010 1310 17015 1340
rect 16975 1305 17015 1310
rect 16400 1285 16420 1305
rect 16985 1285 17005 1305
rect 17095 1285 17115 1350
rect 17740 1285 17760 1595
rect 18485 1390 18505 1595
rect 18475 1385 18515 1390
rect 18475 1355 18480 1385
rect 18510 1355 18515 1385
rect 18475 1350 18515 1355
rect 17835 1340 17875 1345
rect 17835 1310 17840 1340
rect 17870 1310 17875 1340
rect 17835 1305 17875 1310
rect 18230 1340 18270 1345
rect 18230 1310 18235 1340
rect 18265 1310 18270 1340
rect 18230 1305 18270 1310
rect 17845 1285 17865 1305
rect 16240 1280 16280 1285
rect 16240 1250 16245 1280
rect 16275 1250 16280 1280
rect 16240 1245 16280 1250
rect 16335 1280 16375 1285
rect 16335 1250 16340 1280
rect 16370 1250 16375 1280
rect 16335 1245 16375 1250
rect 16394 1275 16424 1285
rect 16394 1255 16399 1275
rect 16419 1255 16424 1275
rect 16394 1245 16424 1255
rect 16460 1280 16500 1285
rect 16460 1250 16465 1280
rect 16495 1250 16500 1280
rect 16460 1245 16500 1250
rect 16810 1280 16850 1285
rect 16810 1250 16815 1280
rect 16845 1250 16850 1280
rect 16810 1245 16850 1250
rect 16920 1280 16960 1285
rect 16920 1250 16925 1280
rect 16955 1250 16960 1280
rect 16920 1245 16960 1250
rect 16980 1275 17010 1285
rect 16980 1255 16985 1275
rect 17005 1255 17010 1275
rect 16980 1245 17010 1255
rect 17030 1280 17070 1285
rect 17030 1250 17035 1280
rect 17065 1250 17070 1280
rect 17030 1245 17070 1250
rect 17090 1275 17120 1285
rect 17090 1255 17095 1275
rect 17115 1255 17120 1275
rect 17090 1245 17120 1255
rect 17140 1280 17180 1285
rect 17140 1250 17145 1280
rect 17175 1250 17180 1280
rect 17140 1245 17180 1250
rect 17605 1280 17645 1285
rect 17605 1250 17610 1280
rect 17640 1250 17645 1280
rect 17605 1245 17645 1250
rect 17670 1280 17710 1285
rect 17670 1250 17675 1280
rect 17705 1250 17710 1280
rect 17670 1245 17710 1250
rect 17730 1275 17760 1285
rect 17730 1255 17735 1275
rect 17755 1255 17760 1275
rect 17730 1245 17760 1255
rect 17780 1280 17820 1285
rect 17780 1250 17785 1280
rect 17815 1250 17820 1280
rect 17780 1245 17820 1250
rect 17840 1275 17870 1285
rect 17840 1255 17845 1275
rect 17865 1255 17870 1275
rect 17840 1245 17870 1255
rect 17890 1280 17930 1285
rect 17890 1250 17895 1280
rect 17925 1250 17930 1280
rect 17890 1245 17930 1250
rect 17955 1280 17995 1285
rect 17955 1250 17960 1280
rect 17990 1250 17995 1280
rect 17955 1245 17995 1250
rect 16300 1105 16330 1115
rect 16300 1085 16305 1105
rect 16325 1085 16330 1105
rect 16300 1075 16330 1085
rect 16410 1105 16440 1115
rect 16410 1085 16415 1105
rect 16435 1085 16440 1105
rect 16410 1075 16440 1085
rect 16865 1110 16905 1115
rect 16865 1080 16870 1110
rect 16900 1080 16905 1110
rect 16865 1075 16905 1080
rect 16975 1110 17015 1115
rect 16975 1080 16980 1110
rect 17010 1080 17015 1110
rect 16975 1075 17015 1080
rect 17085 1110 17125 1115
rect 17085 1080 17090 1110
rect 17120 1080 17125 1110
rect 17085 1075 17125 1080
rect 16305 920 16325 1075
rect 16415 920 16435 1075
rect 17725 1010 17765 1015
rect 17725 980 17730 1010
rect 17760 980 17765 1010
rect 17725 975 17765 980
rect 17835 1010 17875 1015
rect 17835 980 17840 1010
rect 17870 980 17875 1010
rect 18240 1000 18260 1305
rect 18485 1285 18505 1350
rect 18585 1340 18625 1345
rect 18585 1310 18590 1340
rect 18620 1310 18625 1340
rect 18585 1305 18625 1310
rect 18595 1285 18615 1305
rect 18420 1280 18460 1285
rect 18420 1250 18425 1280
rect 18455 1250 18460 1280
rect 18420 1245 18460 1250
rect 18480 1275 18510 1285
rect 18480 1255 18485 1275
rect 18505 1255 18510 1275
rect 18480 1245 18510 1255
rect 18530 1280 18570 1285
rect 18530 1250 18535 1280
rect 18565 1250 18570 1280
rect 18530 1245 18570 1250
rect 18590 1275 18620 1285
rect 18590 1255 18595 1275
rect 18615 1255 18620 1275
rect 18590 1245 18620 1255
rect 18640 1280 18680 1285
rect 18640 1250 18645 1280
rect 18675 1250 18680 1280
rect 18640 1245 18680 1250
rect 18750 1280 18790 1285
rect 18750 1250 18755 1280
rect 18785 1250 18790 1280
rect 18750 1245 18790 1250
rect 18475 1110 18515 1115
rect 18475 1080 18480 1110
rect 18510 1080 18515 1110
rect 18475 1075 18515 1080
rect 18585 1110 18625 1115
rect 18585 1080 18590 1110
rect 18620 1080 18625 1110
rect 18585 1075 18625 1080
rect 18695 1110 18735 1115
rect 18695 1080 18700 1110
rect 18730 1080 18735 1110
rect 18695 1075 18735 1080
rect 17835 975 17875 980
rect 18230 995 18270 1000
rect 18230 965 18235 995
rect 18265 965 18270 995
rect 18230 960 18270 965
rect 18720 995 18760 1000
rect 18720 965 18725 995
rect 18755 965 18760 995
rect 18720 960 18760 965
rect 16160 915 16200 920
rect 16160 885 16165 915
rect 16195 885 16200 915
rect 16160 880 16200 885
rect 16295 915 16335 920
rect 16295 885 16300 915
rect 16330 885 16335 915
rect 16295 880 16335 885
rect 16405 915 16445 920
rect 16405 885 16410 915
rect 16440 885 16445 915
rect 16405 880 16445 885
rect 16170 -1635 16190 880
rect 16970 815 17010 820
rect 16435 805 16475 810
rect 16435 775 16440 805
rect 16470 775 16475 805
rect 16435 770 16475 775
rect 16655 805 16695 810
rect 16655 775 16660 805
rect 16690 775 16695 805
rect 16970 785 16975 815
rect 17005 785 17010 815
rect 16970 780 17010 785
rect 17150 815 17190 820
rect 17150 785 17155 815
rect 17185 785 17190 815
rect 17150 780 17190 785
rect 17330 815 17370 820
rect 17330 785 17335 815
rect 17365 785 17370 815
rect 17330 780 17370 785
rect 17510 815 17550 820
rect 17510 785 17515 815
rect 17545 785 17550 815
rect 17510 780 17550 785
rect 17690 815 17730 820
rect 17690 785 17695 815
rect 17725 785 17730 815
rect 17690 780 17730 785
rect 17870 815 17910 820
rect 17870 785 17875 815
rect 17905 785 17910 815
rect 17870 780 17910 785
rect 18050 815 18090 820
rect 18050 785 18055 815
rect 18085 785 18090 815
rect 18050 780 18090 785
rect 18230 815 18270 820
rect 18230 785 18235 815
rect 18265 785 18270 815
rect 18230 780 18270 785
rect 18410 815 18450 820
rect 18410 785 18415 815
rect 18445 785 18450 815
rect 18410 780 18450 785
rect 18590 815 18630 820
rect 18590 785 18595 815
rect 18625 785 18630 815
rect 18590 780 18630 785
rect 16655 770 16695 775
rect 16445 720 16465 770
rect 16665 720 16685 770
rect 16435 710 16475 720
rect 16435 690 16445 710
rect 16465 690 16475 710
rect 16435 680 16475 690
rect 16545 715 16585 720
rect 16545 685 16550 715
rect 16580 685 16585 715
rect 16545 680 16585 685
rect 16655 710 16695 720
rect 16655 690 16665 710
rect 16685 690 16695 710
rect 16655 680 16695 690
rect 16780 715 16820 720
rect 16780 685 16785 715
rect 16815 685 16820 715
rect 16780 680 16820 685
rect 16480 545 16520 550
rect 16480 515 16485 545
rect 16515 515 16520 545
rect 16480 510 16520 515
rect 16545 540 16585 550
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 16610 545 16650 550
rect 16610 515 16615 545
rect 16645 515 16650 545
rect 16610 510 16650 515
rect 16305 445 16345 450
rect 16305 415 16310 445
rect 16340 415 16345 445
rect 16305 410 16345 415
rect 16260 390 16300 395
rect 16260 360 16265 390
rect 16295 360 16300 390
rect 16260 355 16300 360
rect 16205 345 16245 350
rect 16205 315 16210 345
rect 16240 315 16245 345
rect 16205 310 16245 315
rect 16215 -1075 16235 310
rect 16270 -200 16290 355
rect 16260 -205 16300 -200
rect 16260 -235 16265 -205
rect 16295 -235 16300 -205
rect 16260 -240 16300 -235
rect 16205 -1080 16245 -1075
rect 16205 -1110 16210 -1080
rect 16240 -1110 16245 -1080
rect 16205 -1115 16245 -1110
rect 16160 -1640 16200 -1635
rect 16160 -1670 16165 -1640
rect 16195 -1670 16200 -1640
rect 16160 -1675 16200 -1670
rect 16105 -1685 16145 -1680
rect 16105 -1715 16110 -1685
rect 16140 -1715 16145 -1685
rect 16105 -1720 16145 -1715
rect 16155 -1760 16195 -1755
rect 16155 -1790 16160 -1760
rect 16190 -1790 16195 -1760
rect 16155 -1795 16195 -1790
rect 16165 -3020 16185 -1795
rect 16270 -1890 16290 -240
rect 16315 -365 16335 410
rect 16555 350 16575 510
rect 16790 395 16810 680
rect 16840 545 16880 550
rect 16840 515 16845 545
rect 16875 515 16880 545
rect 16840 510 16880 515
rect 16780 390 16820 395
rect 16780 360 16785 390
rect 16815 360 16820 390
rect 16780 355 16820 360
rect 16545 345 16585 350
rect 16545 315 16550 345
rect 16580 315 16585 345
rect 16545 310 16585 315
rect 16420 185 16460 190
rect 16420 155 16425 185
rect 16455 155 16460 185
rect 16420 150 16460 155
rect 16540 185 16580 190
rect 16540 155 16545 185
rect 16575 155 16580 185
rect 16540 150 16580 155
rect 16660 185 16700 190
rect 16660 155 16665 185
rect 16695 155 16700 185
rect 16660 150 16700 155
rect 16780 185 16820 190
rect 16780 155 16785 185
rect 16815 155 16820 185
rect 16780 150 16820 155
rect 16430 130 16450 150
rect 16550 130 16570 150
rect 16670 130 16690 150
rect 16790 130 16810 150
rect 16850 130 16870 510
rect 17060 440 17100 450
rect 17060 420 17070 440
rect 17090 420 17100 440
rect 17060 410 17100 420
rect 17240 440 17280 450
rect 17240 420 17250 440
rect 17270 420 17280 440
rect 17240 410 17280 420
rect 17420 440 17460 450
rect 17420 420 17430 440
rect 17450 420 17460 440
rect 17420 410 17460 420
rect 17600 445 17640 450
rect 17600 415 17605 445
rect 17635 415 17640 445
rect 17600 410 17640 415
rect 17690 440 17730 450
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 17780 440 17820 450
rect 17780 420 17790 440
rect 17810 420 17820 440
rect 17780 410 17820 420
rect 17960 445 18000 450
rect 17960 415 17965 445
rect 17995 415 18000 445
rect 17960 410 18000 415
rect 18140 440 18180 450
rect 18140 420 18150 440
rect 18170 420 18180 440
rect 18140 410 18180 420
rect 18320 440 18360 450
rect 18320 420 18330 440
rect 18350 420 18360 440
rect 18320 410 18360 420
rect 18410 440 18450 450
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 18500 440 18540 450
rect 18500 420 18510 440
rect 18530 420 18540 440
rect 18500 410 18540 420
rect 17070 305 17090 410
rect 17250 350 17270 410
rect 17430 395 17450 410
rect 17420 390 17460 395
rect 17420 360 17425 390
rect 17455 360 17460 390
rect 17420 355 17460 360
rect 17240 345 17280 350
rect 17240 315 17245 345
rect 17275 315 17280 345
rect 17240 310 17280 315
rect 17060 300 17100 305
rect 17060 270 17065 300
rect 17095 270 17100 300
rect 17060 265 17100 270
rect 16900 185 16940 190
rect 16900 155 16905 185
rect 16935 155 16940 185
rect 16900 150 16940 155
rect 17020 185 17060 190
rect 17020 155 17025 185
rect 17055 155 17060 185
rect 17020 150 17060 155
rect 17140 185 17180 190
rect 17140 155 17145 185
rect 17175 155 17180 185
rect 17140 150 17180 155
rect 17260 185 17300 190
rect 17260 155 17265 185
rect 17295 155 17300 185
rect 17260 150 17300 155
rect 17380 185 17420 190
rect 17380 155 17385 185
rect 17415 155 17420 185
rect 17380 150 17420 155
rect 17500 185 17540 190
rect 17500 155 17505 185
rect 17535 155 17540 185
rect 17500 150 17540 155
rect 17620 185 17660 190
rect 17620 155 17625 185
rect 17655 155 17660 185
rect 17620 150 17660 155
rect 16910 130 16930 150
rect 17030 130 17050 150
rect 17150 130 17170 150
rect 17270 130 17290 150
rect 17390 130 17410 150
rect 17510 130 17530 150
rect 17630 130 17650 150
rect 17700 130 17720 410
rect 17790 305 17810 410
rect 18150 395 18170 410
rect 18140 390 18180 395
rect 18140 360 18145 390
rect 18175 360 18180 390
rect 18140 355 18180 360
rect 18330 350 18350 410
rect 18420 405 18440 410
rect 18320 345 18360 350
rect 18320 315 18325 345
rect 18355 315 18360 345
rect 18320 310 18360 315
rect 18510 305 18530 410
rect 17780 300 17820 305
rect 17780 270 17785 300
rect 17815 270 17820 300
rect 17780 265 17820 270
rect 18500 300 18540 305
rect 18500 270 18505 300
rect 18535 270 18540 300
rect 18500 265 18540 270
rect 18730 255 18750 960
rect 19010 825 19050 830
rect 19010 795 19015 825
rect 19045 795 19050 825
rect 19010 790 19050 795
rect 19020 770 19040 790
rect 18945 765 18985 770
rect 18945 735 18950 765
rect 18980 735 18985 765
rect 18945 730 18985 735
rect 19010 765 19050 770
rect 19010 735 19015 765
rect 19045 735 19050 765
rect 19010 730 19050 735
rect 19120 765 19160 770
rect 19120 735 19125 765
rect 19155 735 19160 765
rect 19120 730 19160 735
rect 19270 500 19290 1595
rect 19325 915 19365 920
rect 19325 885 19330 915
rect 19360 885 19365 915
rect 19325 880 19365 885
rect 19031 490 19061 500
rect 19031 470 19036 490
rect 19056 470 19061 490
rect 19031 460 19061 470
rect 19080 495 19120 500
rect 19080 465 19085 495
rect 19115 465 19120 495
rect 19080 460 19120 465
rect 19260 495 19300 500
rect 19260 465 19265 495
rect 19295 465 19300 495
rect 19260 460 19300 465
rect 19035 255 19055 460
rect 18000 250 18040 255
rect 18000 220 18005 250
rect 18035 220 18040 250
rect 18000 215 18040 220
rect 18720 250 18760 255
rect 18720 220 18725 250
rect 18755 220 18760 250
rect 18720 215 18760 220
rect 19025 250 19065 255
rect 19025 220 19030 250
rect 19060 220 19065 250
rect 19025 215 19065 220
rect 17940 185 17980 190
rect 17940 155 17945 185
rect 17975 155 17980 185
rect 17940 150 17980 155
rect 17950 130 17970 150
rect 18010 130 18030 215
rect 18060 185 18100 190
rect 18060 155 18065 185
rect 18095 155 18100 185
rect 18060 150 18100 155
rect 18180 185 18220 190
rect 18180 155 18185 185
rect 18215 155 18220 185
rect 18180 150 18220 155
rect 18300 185 18340 190
rect 18300 155 18305 185
rect 18335 155 18340 185
rect 18300 150 18340 155
rect 18420 185 18460 190
rect 18420 155 18425 185
rect 18455 155 18460 185
rect 18420 150 18460 155
rect 18540 185 18580 190
rect 18540 155 18545 185
rect 18575 155 18580 185
rect 18540 150 18580 155
rect 18660 185 18700 190
rect 18660 155 18665 185
rect 18695 155 18700 185
rect 18660 150 18700 155
rect 18780 185 18820 190
rect 18780 155 18785 185
rect 18815 155 18820 185
rect 18780 150 18820 155
rect 18900 185 18940 190
rect 18900 155 18905 185
rect 18935 155 18940 185
rect 18900 150 18940 155
rect 19020 185 19060 190
rect 19020 155 19025 185
rect 19055 155 19060 185
rect 19020 150 19060 155
rect 19140 185 19180 190
rect 19140 155 19145 185
rect 19175 155 19180 185
rect 19140 150 19180 155
rect 18070 130 18090 150
rect 18190 130 18210 150
rect 18310 130 18330 150
rect 18430 130 18450 150
rect 18550 130 18570 150
rect 18670 130 18690 150
rect 18790 130 18810 150
rect 18910 130 18930 150
rect 19030 130 19050 150
rect 19150 130 19170 150
rect 16425 120 16455 130
rect 16425 100 16430 120
rect 16450 100 16455 120
rect 16425 85 16455 100
rect 16480 125 16520 130
rect 16480 95 16485 125
rect 16515 95 16520 125
rect 16480 90 16520 95
rect 16545 120 16575 130
rect 16545 100 16550 120
rect 16570 100 16575 120
rect 16545 90 16575 100
rect 16665 120 16695 130
rect 16665 100 16670 120
rect 16690 100 16695 120
rect 16665 90 16695 100
rect 16785 120 16815 130
rect 16785 100 16790 120
rect 16810 100 16815 120
rect 16785 90 16815 100
rect 16840 125 16880 130
rect 16840 95 16845 125
rect 16875 95 16880 125
rect 16840 90 16880 95
rect 16905 120 16935 130
rect 16905 100 16910 120
rect 16930 100 16935 120
rect 16905 90 16935 100
rect 17025 120 17055 130
rect 17025 100 17030 120
rect 17050 100 17055 120
rect 17025 90 17055 100
rect 17145 120 17175 130
rect 17145 100 17150 120
rect 17170 100 17175 120
rect 17145 90 17175 100
rect 17200 125 17240 130
rect 17200 95 17205 125
rect 17235 95 17240 125
rect 17200 90 17240 95
rect 17265 120 17295 130
rect 17265 100 17270 120
rect 17290 100 17295 120
rect 17265 90 17295 100
rect 17385 120 17415 130
rect 17385 100 17390 120
rect 17410 100 17415 120
rect 17385 90 17415 100
rect 17505 120 17535 130
rect 17505 100 17510 120
rect 17530 100 17535 120
rect 17505 90 17535 100
rect 17560 125 17600 130
rect 17560 95 17565 125
rect 17595 95 17600 125
rect 17560 90 17600 95
rect 17625 120 17655 130
rect 17625 100 17630 120
rect 17650 100 17655 120
rect 17625 85 17655 100
rect 17690 125 17730 130
rect 17690 95 17695 125
rect 17725 95 17730 125
rect 17690 90 17730 95
rect 17870 125 17910 130
rect 17870 95 17875 125
rect 17905 95 17910 125
rect 17870 90 17910 95
rect 17945 120 17975 130
rect 17945 100 17950 120
rect 17970 100 17975 120
rect 16510 -50 16550 -40
rect 16510 -70 16520 -50
rect 16540 -70 16550 -50
rect 16510 -80 16550 -70
rect 16600 -45 16640 -40
rect 16600 -75 16605 -45
rect 16635 -75 16640 -45
rect 16600 -80 16640 -75
rect 16720 -50 16760 -40
rect 16720 -70 16730 -50
rect 16750 -70 16760 -50
rect 16720 -80 16760 -70
rect 16840 -50 16880 -40
rect 16840 -70 16850 -50
rect 16870 -70 16880 -50
rect 16840 -80 16880 -70
rect 16960 -45 17000 -40
rect 16960 -75 16965 -45
rect 16995 -75 17000 -45
rect 16960 -80 17000 -75
rect 17080 -50 17120 -40
rect 17080 -70 17090 -50
rect 17110 -70 17120 -50
rect 17080 -80 17120 -70
rect 17200 -50 17240 -40
rect 17200 -70 17210 -50
rect 17230 -70 17240 -50
rect 17200 -80 17240 -70
rect 17320 -45 17360 -40
rect 17320 -75 17325 -45
rect 17355 -75 17360 -45
rect 17320 -80 17360 -75
rect 17440 -50 17480 -40
rect 17440 -70 17450 -50
rect 17470 -70 17480 -50
rect 17440 -80 17480 -70
rect 17535 -50 17565 -40
rect 17535 -70 17540 -50
rect 17560 -70 17565 -50
rect 17535 -80 17565 -70
rect 16520 -100 16540 -80
rect 16730 -100 16750 -80
rect 16850 -100 16870 -80
rect 16510 -105 16550 -100
rect 16510 -135 16515 -105
rect 16545 -135 16550 -105
rect 16510 -140 16550 -135
rect 16720 -105 16760 -100
rect 16720 -135 16725 -105
rect 16755 -135 16760 -105
rect 16720 -140 16760 -135
rect 16840 -105 16880 -100
rect 16840 -135 16845 -105
rect 16875 -135 16880 -105
rect 16840 -140 16880 -135
rect 16980 -185 17000 -80
rect 17090 -100 17110 -80
rect 17210 -100 17230 -80
rect 17450 -100 17470 -80
rect 17540 -100 17560 -80
rect 17080 -105 17120 -100
rect 17080 -135 17085 -105
rect 17115 -135 17120 -105
rect 17080 -140 17120 -135
rect 17200 -105 17240 -100
rect 17200 -135 17205 -105
rect 17235 -135 17240 -105
rect 17200 -140 17240 -135
rect 17440 -105 17480 -100
rect 17440 -135 17445 -105
rect 17475 -135 17480 -105
rect 17440 -140 17480 -135
rect 17530 -105 17570 -100
rect 17530 -135 17535 -105
rect 17565 -135 17570 -105
rect 17530 -140 17570 -135
rect 16970 -190 17010 -185
rect 16910 -205 16950 -200
rect 16910 -235 16915 -205
rect 16945 -235 16950 -205
rect 16970 -220 16975 -190
rect 17005 -220 17010 -190
rect 16970 -225 17010 -220
rect 16910 -240 16950 -235
rect 16980 -245 17000 -225
rect 17090 -245 17110 -140
rect 17210 -190 17250 -185
rect 17210 -220 17215 -190
rect 17245 -220 17250 -190
rect 17210 -225 17250 -220
rect 17450 -190 17490 -185
rect 17450 -220 17455 -190
rect 17485 -220 17490 -190
rect 17450 -225 17490 -220
rect 17220 -245 17240 -225
rect 17460 -245 17480 -225
rect 16850 -250 16890 -245
rect 16850 -280 16855 -250
rect 16885 -280 16890 -250
rect 16850 -285 16890 -280
rect 16975 -255 17005 -245
rect 16975 -275 16980 -255
rect 17000 -275 17005 -255
rect 16975 -285 17005 -275
rect 17090 -250 17130 -245
rect 17090 -280 17095 -250
rect 17125 -280 17130 -250
rect 17090 -285 17130 -280
rect 17215 -255 17245 -245
rect 17215 -275 17220 -255
rect 17240 -275 17245 -255
rect 17215 -285 17245 -275
rect 17330 -250 17370 -245
rect 17330 -280 17335 -250
rect 17365 -280 17370 -250
rect 17330 -285 17370 -280
rect 17455 -255 17485 -245
rect 17455 -275 17460 -255
rect 17480 -275 17485 -255
rect 17455 -285 17485 -275
rect 17565 -310 17595 -305
rect 17565 -345 17595 -340
rect 16305 -370 16345 -365
rect 16305 -400 16310 -370
rect 16340 -400 16345 -370
rect 16305 -405 16345 -400
rect 16850 -370 16890 -365
rect 16850 -400 16855 -370
rect 16885 -400 16890 -370
rect 16850 -405 16890 -400
rect 16915 -375 16945 -365
rect 16915 -395 16920 -375
rect 16940 -395 16945 -375
rect 16915 -405 16945 -395
rect 17035 -375 17065 -365
rect 17035 -395 17040 -375
rect 17060 -395 17065 -375
rect 17035 -405 17065 -395
rect 17155 -375 17185 -365
rect 17155 -395 17160 -375
rect 17180 -395 17185 -375
rect 17155 -405 17185 -395
rect 17275 -375 17305 -365
rect 17275 -395 17280 -375
rect 17300 -395 17305 -375
rect 17275 -405 17305 -395
rect 17395 -375 17425 -365
rect 17395 -395 17400 -375
rect 17420 -395 17425 -375
rect 17395 -405 17425 -395
rect 16920 -425 16940 -405
rect 17040 -425 17060 -405
rect 17160 -425 17180 -405
rect 17280 -425 17300 -405
rect 17400 -425 17420 -405
rect 16530 -430 16570 -425
rect 16530 -460 16535 -430
rect 16565 -460 16570 -430
rect 16530 -465 16570 -460
rect 16910 -430 16950 -425
rect 16910 -460 16915 -430
rect 16945 -460 16950 -430
rect 16910 -465 16950 -460
rect 17030 -430 17070 -425
rect 17030 -460 17035 -430
rect 17065 -460 17070 -430
rect 17030 -465 17070 -460
rect 17150 -430 17190 -425
rect 17150 -460 17155 -430
rect 17185 -460 17190 -430
rect 17150 -465 17190 -460
rect 17270 -430 17310 -425
rect 17270 -460 17275 -430
rect 17305 -460 17310 -430
rect 17270 -465 17310 -460
rect 17390 -430 17430 -425
rect 17390 -460 17395 -430
rect 17425 -460 17430 -430
rect 17390 -465 17430 -460
rect 16540 -540 16560 -465
rect 16620 -530 16660 -525
rect 16530 -550 16570 -540
rect 16530 -570 16540 -550
rect 16560 -570 16570 -550
rect 16620 -560 16625 -530
rect 16655 -560 16660 -530
rect 16620 -565 16660 -560
rect 16740 -530 16780 -525
rect 16740 -560 16745 -530
rect 16775 -560 16780 -530
rect 16740 -565 16780 -560
rect 16860 -530 16900 -525
rect 16860 -560 16865 -530
rect 16895 -560 16900 -530
rect 16860 -565 16900 -560
rect 16980 -530 17020 -525
rect 16980 -560 16985 -530
rect 17015 -560 17020 -530
rect 16980 -565 17020 -560
rect 17300 -530 17340 -525
rect 17300 -560 17305 -530
rect 17335 -560 17340 -530
rect 17300 -565 17340 -560
rect 17420 -530 17460 -525
rect 17420 -560 17425 -530
rect 17455 -560 17460 -530
rect 17420 -565 17460 -560
rect 17540 -530 17580 -525
rect 17540 -560 17545 -530
rect 17575 -560 17580 -530
rect 17700 -540 17720 90
rect 17780 -310 17820 -305
rect 17780 -340 17785 -310
rect 17815 -340 17820 -310
rect 17780 -345 17820 -340
rect 17540 -565 17580 -560
rect 17690 -550 17730 -540
rect 16530 -580 16570 -570
rect 17690 -570 17700 -550
rect 17720 -570 17730 -550
rect 17690 -580 17730 -570
rect 17790 -840 17810 -345
rect 17880 -540 17900 90
rect 17945 85 17975 100
rect 18000 125 18040 130
rect 18000 95 18005 125
rect 18035 95 18040 125
rect 18000 90 18040 95
rect 18065 120 18095 130
rect 18065 100 18070 120
rect 18090 100 18095 120
rect 18065 90 18095 100
rect 18185 120 18215 130
rect 18185 100 18190 120
rect 18210 100 18215 120
rect 18185 90 18215 100
rect 18305 120 18335 130
rect 18305 100 18310 120
rect 18330 100 18335 120
rect 18305 90 18335 100
rect 18360 125 18400 130
rect 18360 95 18365 125
rect 18395 95 18400 125
rect 18360 90 18400 95
rect 18425 120 18455 130
rect 18425 100 18430 120
rect 18450 100 18455 120
rect 18425 90 18455 100
rect 18545 120 18575 130
rect 18545 100 18550 120
rect 18570 100 18575 120
rect 18545 90 18575 100
rect 18665 120 18695 130
rect 18665 100 18670 120
rect 18690 100 18695 120
rect 18665 90 18695 100
rect 18720 125 18760 130
rect 18720 95 18725 125
rect 18755 95 18760 125
rect 18720 90 18760 95
rect 18785 120 18815 130
rect 18785 100 18790 120
rect 18810 100 18815 120
rect 18785 90 18815 100
rect 18905 120 18935 130
rect 18905 100 18910 120
rect 18930 100 18935 120
rect 18905 90 18935 100
rect 19025 120 19055 130
rect 19025 100 19030 120
rect 19050 100 19055 120
rect 19025 90 19055 100
rect 19080 125 19120 130
rect 19080 95 19085 125
rect 19115 95 19120 125
rect 19080 90 19120 95
rect 19145 120 19175 130
rect 19145 100 19150 120
rect 19170 100 19175 120
rect 19145 85 19175 100
rect 18035 -50 18065 -40
rect 18035 -70 18040 -50
rect 18060 -70 18065 -50
rect 18035 -80 18065 -70
rect 18120 -50 18160 -40
rect 18120 -70 18130 -50
rect 18150 -70 18160 -50
rect 18120 -80 18160 -70
rect 18240 -45 18280 -40
rect 18240 -75 18245 -45
rect 18275 -75 18280 -45
rect 18240 -80 18280 -75
rect 18360 -50 18400 -40
rect 18360 -70 18370 -50
rect 18390 -70 18400 -50
rect 18360 -80 18400 -70
rect 18480 -50 18520 -40
rect 18480 -70 18490 -50
rect 18510 -70 18520 -50
rect 18480 -80 18520 -70
rect 18600 -45 18640 -40
rect 18600 -75 18605 -45
rect 18635 -75 18640 -45
rect 18600 -80 18640 -75
rect 18720 -50 18760 -40
rect 18720 -70 18730 -50
rect 18750 -70 18760 -50
rect 18720 -80 18760 -70
rect 18840 -50 18880 -40
rect 18840 -70 18850 -50
rect 18870 -70 18880 -50
rect 18840 -80 18880 -70
rect 18960 -45 19000 -40
rect 18960 -75 18965 -45
rect 18995 -75 19000 -45
rect 18960 -80 19000 -75
rect 19050 -50 19090 -40
rect 19050 -70 19060 -50
rect 19080 -70 19090 -50
rect 19050 -80 19090 -70
rect 18040 -100 18060 -80
rect 18130 -100 18150 -80
rect 18370 -100 18390 -80
rect 18490 -100 18510 -80
rect 18030 -105 18070 -100
rect 18030 -135 18035 -105
rect 18065 -135 18070 -105
rect 18030 -140 18070 -135
rect 18120 -105 18160 -100
rect 18120 -135 18125 -105
rect 18155 -135 18160 -105
rect 18120 -140 18160 -135
rect 18360 -105 18400 -100
rect 18360 -135 18365 -105
rect 18395 -135 18400 -105
rect 18360 -140 18400 -135
rect 18480 -105 18520 -100
rect 18480 -135 18485 -105
rect 18515 -135 18520 -105
rect 18480 -140 18520 -135
rect 18110 -190 18150 -185
rect 18110 -220 18115 -190
rect 18145 -220 18150 -190
rect 18110 -225 18150 -220
rect 18350 -190 18390 -185
rect 18350 -220 18355 -190
rect 18385 -220 18390 -190
rect 18350 -225 18390 -220
rect 18120 -245 18140 -225
rect 18360 -245 18380 -225
rect 18480 -245 18500 -140
rect 18600 -185 18620 -80
rect 18730 -100 18750 -80
rect 18850 -100 18870 -80
rect 19060 -100 19080 -80
rect 18720 -105 18760 -100
rect 18720 -135 18725 -105
rect 18755 -135 18760 -105
rect 18720 -140 18760 -135
rect 18840 -105 18880 -100
rect 18840 -135 18845 -105
rect 18875 -135 18880 -105
rect 18840 -140 18880 -135
rect 19050 -105 19090 -100
rect 19050 -135 19055 -105
rect 19085 -135 19090 -105
rect 19050 -140 19090 -135
rect 18590 -190 18630 -185
rect 18590 -220 18595 -190
rect 18625 -220 18630 -190
rect 18590 -225 18630 -220
rect 18650 -205 18690 -200
rect 18600 -245 18620 -225
rect 18650 -235 18655 -205
rect 18685 -235 18690 -205
rect 18650 -240 18690 -235
rect 18115 -255 18145 -245
rect 18115 -275 18120 -255
rect 18140 -275 18145 -255
rect 18115 -285 18145 -275
rect 18230 -250 18270 -245
rect 18230 -280 18235 -250
rect 18265 -280 18270 -250
rect 18230 -285 18270 -280
rect 18355 -255 18385 -245
rect 18355 -275 18360 -255
rect 18380 -275 18385 -255
rect 18355 -285 18385 -275
rect 18470 -250 18510 -245
rect 18470 -280 18475 -250
rect 18505 -280 18510 -250
rect 18470 -285 18510 -280
rect 18595 -255 18625 -245
rect 18595 -275 18600 -255
rect 18620 -275 18625 -255
rect 18595 -285 18625 -275
rect 18710 -250 18750 -245
rect 18710 -280 18715 -250
rect 18745 -280 18750 -250
rect 18710 -285 18750 -280
rect 18005 -310 18035 -305
rect 18005 -345 18035 -340
rect 19335 -365 19355 880
rect 19415 305 19435 1600
rect 19460 445 19500 450
rect 19460 415 19465 445
rect 19495 415 19500 445
rect 19460 410 19500 415
rect 19405 300 19445 305
rect 19405 270 19410 300
rect 19440 270 19445 300
rect 19405 265 19445 270
rect 19415 -200 19435 265
rect 19405 -205 19445 -200
rect 19405 -235 19410 -205
rect 19440 -235 19445 -205
rect 19405 -240 19445 -235
rect 18175 -375 18205 -365
rect 18175 -395 18180 -375
rect 18200 -395 18205 -375
rect 18175 -405 18205 -395
rect 18295 -375 18325 -365
rect 18295 -395 18300 -375
rect 18320 -395 18325 -375
rect 18295 -405 18325 -395
rect 18415 -375 18445 -365
rect 18415 -395 18420 -375
rect 18440 -395 18445 -375
rect 18415 -405 18445 -395
rect 18535 -375 18565 -365
rect 18535 -395 18540 -375
rect 18560 -395 18565 -375
rect 18535 -405 18565 -395
rect 18655 -375 18685 -365
rect 18655 -395 18660 -375
rect 18680 -395 18685 -375
rect 18655 -405 18685 -395
rect 18710 -370 18750 -365
rect 18710 -400 18715 -370
rect 18745 -400 18750 -370
rect 18710 -405 18750 -400
rect 19325 -370 19365 -365
rect 19325 -400 19330 -370
rect 19360 -400 19365 -370
rect 19325 -405 19365 -400
rect 18180 -425 18200 -405
rect 18300 -425 18320 -405
rect 18420 -425 18440 -405
rect 18540 -425 18560 -405
rect 18660 -425 18680 -405
rect 18170 -430 18210 -425
rect 18170 -460 18175 -430
rect 18205 -460 18210 -430
rect 18170 -465 18210 -460
rect 18290 -430 18330 -425
rect 18290 -460 18295 -430
rect 18325 -460 18330 -430
rect 18290 -465 18330 -460
rect 18410 -430 18450 -425
rect 18410 -460 18415 -430
rect 18445 -460 18450 -430
rect 18410 -465 18450 -460
rect 18530 -430 18570 -425
rect 18530 -460 18535 -430
rect 18565 -460 18570 -430
rect 18530 -465 18570 -460
rect 18650 -430 18690 -425
rect 18650 -460 18655 -430
rect 18685 -460 18690 -430
rect 18650 -465 18690 -460
rect 19030 -430 19070 -425
rect 19030 -460 19035 -430
rect 19065 -460 19070 -430
rect 19030 -465 19070 -460
rect 18020 -530 18060 -525
rect 17870 -550 17910 -540
rect 17870 -570 17880 -550
rect 17900 -570 17910 -550
rect 18020 -560 18025 -530
rect 18055 -560 18060 -530
rect 18020 -565 18060 -560
rect 18140 -530 18180 -525
rect 18140 -560 18145 -530
rect 18175 -560 18180 -530
rect 18140 -565 18180 -560
rect 18260 -530 18300 -525
rect 18260 -560 18265 -530
rect 18295 -560 18300 -530
rect 18260 -565 18300 -560
rect 18580 -530 18620 -525
rect 18580 -560 18585 -530
rect 18615 -560 18620 -530
rect 18580 -565 18620 -560
rect 18700 -530 18740 -525
rect 18700 -560 18705 -530
rect 18735 -560 18740 -530
rect 18700 -565 18740 -560
rect 18820 -530 18860 -525
rect 18820 -560 18825 -530
rect 18855 -560 18860 -530
rect 18820 -565 18860 -560
rect 18940 -530 18980 -525
rect 18940 -560 18945 -530
rect 18975 -560 18980 -530
rect 19040 -540 19060 -465
rect 18940 -565 18980 -560
rect 19030 -550 19070 -540
rect 17870 -580 17910 -570
rect 19030 -570 19040 -550
rect 19060 -570 19070 -550
rect 19030 -580 19070 -570
rect 17110 -845 17150 -840
rect 17110 -875 17115 -845
rect 17145 -875 17150 -845
rect 17110 -880 17150 -875
rect 17780 -845 17820 -840
rect 17780 -875 17785 -845
rect 17815 -875 17820 -845
rect 17780 -880 17820 -875
rect 18450 -845 18490 -840
rect 18450 -875 18455 -845
rect 18485 -875 18490 -845
rect 18450 -880 18490 -875
rect 16740 -995 16780 -990
rect 16740 -1025 16745 -995
rect 16775 -1025 16780 -995
rect 16740 -1030 16780 -1025
rect 16820 -995 16860 -990
rect 16820 -1025 16825 -995
rect 16855 -1025 16860 -995
rect 16820 -1030 16860 -1025
rect 16900 -995 16940 -990
rect 16900 -1025 16905 -995
rect 16935 -1025 16940 -995
rect 16900 -1030 16940 -1025
rect 16980 -995 17020 -990
rect 16980 -1025 16985 -995
rect 17015 -1025 17020 -995
rect 16980 -1030 17020 -1025
rect 17060 -995 17100 -990
rect 17060 -1025 17065 -995
rect 17095 -1025 17100 -995
rect 17060 -1030 17100 -1025
rect 17140 -995 17180 -990
rect 17140 -1025 17145 -995
rect 17175 -1025 17180 -995
rect 17140 -1030 17180 -1025
rect 17220 -995 17260 -990
rect 17220 -1025 17225 -995
rect 17255 -1025 17260 -995
rect 17220 -1030 17260 -1025
rect 17300 -995 17340 -990
rect 17300 -1025 17305 -995
rect 17335 -1025 17340 -995
rect 17300 -1030 17340 -1025
rect 17380 -995 17420 -990
rect 17380 -1025 17385 -995
rect 17415 -1025 17420 -995
rect 17380 -1030 17420 -1025
rect 17460 -995 17500 -990
rect 17460 -1025 17465 -995
rect 17495 -1025 17500 -995
rect 17460 -1030 17500 -1025
rect 17540 -995 17580 -990
rect 17540 -1025 17545 -995
rect 17575 -1025 17580 -995
rect 17540 -1030 17580 -1025
rect 17620 -995 17660 -990
rect 17620 -1025 17625 -995
rect 17655 -1025 17660 -995
rect 17620 -1030 17660 -1025
rect 17700 -995 17740 -990
rect 17700 -1025 17705 -995
rect 17735 -1025 17740 -995
rect 17700 -1030 17740 -1025
rect 17780 -995 17820 -990
rect 17780 -1025 17785 -995
rect 17815 -1025 17820 -995
rect 17780 -1030 17820 -1025
rect 17860 -995 17900 -990
rect 17860 -1025 17865 -995
rect 17895 -1025 17900 -995
rect 17860 -1030 17900 -1025
rect 17940 -995 17980 -990
rect 17940 -1025 17945 -995
rect 17975 -1025 17980 -995
rect 17940 -1030 17980 -1025
rect 18020 -995 18060 -990
rect 18020 -1025 18025 -995
rect 18055 -1025 18060 -995
rect 18020 -1030 18060 -1025
rect 18100 -995 18140 -990
rect 18100 -1025 18105 -995
rect 18135 -1025 18140 -995
rect 18100 -1030 18140 -1025
rect 18180 -995 18220 -990
rect 18180 -1025 18185 -995
rect 18215 -1025 18220 -995
rect 18180 -1030 18220 -1025
rect 18260 -995 18300 -990
rect 18260 -1025 18265 -995
rect 18295 -1025 18300 -995
rect 18260 -1030 18300 -1025
rect 18340 -995 18380 -990
rect 18340 -1025 18345 -995
rect 18375 -1025 18380 -995
rect 18340 -1030 18380 -1025
rect 18420 -995 18460 -990
rect 18420 -1025 18425 -995
rect 18455 -1025 18460 -995
rect 18420 -1030 18460 -1025
rect 18500 -995 18540 -990
rect 18500 -1025 18505 -995
rect 18535 -1025 18540 -995
rect 18500 -1030 18540 -1025
rect 18580 -995 18620 -990
rect 18580 -1025 18585 -995
rect 18615 -1025 18620 -995
rect 18580 -1030 18620 -1025
rect 18660 -995 18700 -990
rect 18660 -1025 18665 -995
rect 18695 -1025 18700 -995
rect 18660 -1030 18700 -1025
rect 18740 -995 18780 -990
rect 18740 -1025 18745 -995
rect 18775 -1025 18780 -995
rect 18740 -1030 18780 -1025
rect 16700 -1080 16740 -1075
rect 16700 -1110 16705 -1080
rect 16735 -1110 16740 -1080
rect 16700 -1115 16740 -1110
rect 18895 -1080 18935 -1075
rect 18895 -1110 18900 -1080
rect 18930 -1110 18935 -1080
rect 18895 -1115 18935 -1110
rect 17165 -1200 17205 -1195
rect 17165 -1230 17170 -1200
rect 17200 -1230 17205 -1200
rect 17165 -1235 17205 -1230
rect 17780 -1200 17820 -1195
rect 17780 -1230 17785 -1200
rect 17815 -1230 17820 -1200
rect 17780 -1235 17820 -1230
rect 18395 -1200 18435 -1195
rect 18395 -1230 18400 -1200
rect 18430 -1230 18435 -1200
rect 18395 -1235 18435 -1230
rect 17175 -1265 17195 -1235
rect 17790 -1265 17810 -1235
rect 18405 -1265 18425 -1235
rect 16890 -1270 16930 -1265
rect 16890 -1300 16895 -1270
rect 16925 -1300 16930 -1270
rect 16890 -1305 16930 -1300
rect 17000 -1270 17040 -1265
rect 17000 -1300 17005 -1270
rect 17035 -1300 17040 -1270
rect 17000 -1305 17040 -1300
rect 17110 -1270 17150 -1265
rect 17110 -1300 17115 -1270
rect 17145 -1300 17150 -1270
rect 17110 -1305 17150 -1300
rect 17170 -1275 17200 -1265
rect 17170 -1295 17175 -1275
rect 17195 -1295 17200 -1275
rect 17170 -1305 17200 -1295
rect 17220 -1270 17260 -1265
rect 17220 -1300 17225 -1270
rect 17255 -1300 17260 -1270
rect 17220 -1305 17260 -1300
rect 17330 -1270 17370 -1265
rect 17330 -1300 17335 -1270
rect 17365 -1300 17370 -1270
rect 17330 -1305 17370 -1300
rect 17505 -1270 17545 -1265
rect 17505 -1300 17510 -1270
rect 17540 -1300 17545 -1270
rect 17505 -1305 17545 -1300
rect 17615 -1270 17655 -1265
rect 17615 -1300 17620 -1270
rect 17650 -1300 17655 -1270
rect 17615 -1305 17655 -1300
rect 17725 -1270 17765 -1265
rect 17725 -1300 17730 -1270
rect 17760 -1300 17765 -1270
rect 17725 -1305 17765 -1300
rect 17785 -1275 17815 -1265
rect 17785 -1295 17790 -1275
rect 17810 -1295 17815 -1275
rect 17785 -1305 17815 -1295
rect 17835 -1270 17875 -1265
rect 17835 -1300 17840 -1270
rect 17870 -1300 17875 -1270
rect 17835 -1305 17875 -1300
rect 17945 -1270 17985 -1265
rect 17945 -1300 17950 -1270
rect 17980 -1300 17985 -1270
rect 17945 -1305 17985 -1300
rect 18055 -1270 18095 -1265
rect 18055 -1300 18060 -1270
rect 18090 -1300 18095 -1270
rect 18055 -1305 18095 -1300
rect 18230 -1270 18270 -1265
rect 18230 -1300 18235 -1270
rect 18265 -1300 18270 -1270
rect 18230 -1305 18270 -1300
rect 18340 -1270 18380 -1265
rect 18340 -1300 18345 -1270
rect 18375 -1300 18380 -1270
rect 18340 -1305 18380 -1300
rect 18400 -1275 18430 -1265
rect 18400 -1295 18405 -1275
rect 18425 -1295 18430 -1275
rect 18400 -1305 18430 -1295
rect 18450 -1270 18490 -1265
rect 18450 -1300 18455 -1270
rect 18485 -1300 18490 -1270
rect 18450 -1305 18490 -1300
rect 18560 -1270 18600 -1265
rect 18560 -1300 18565 -1270
rect 18595 -1300 18600 -1270
rect 18560 -1305 18600 -1300
rect 18670 -1270 18710 -1265
rect 18670 -1300 18675 -1270
rect 18705 -1300 18710 -1270
rect 18670 -1305 18710 -1300
rect 16945 -1445 16985 -1435
rect 16945 -1465 16955 -1445
rect 16975 -1465 16985 -1445
rect 16945 -1475 16985 -1465
rect 17055 -1440 17095 -1435
rect 17055 -1470 17060 -1440
rect 17090 -1470 17095 -1440
rect 17055 -1475 17095 -1470
rect 17165 -1445 17205 -1435
rect 17165 -1465 17175 -1445
rect 17195 -1465 17205 -1445
rect 17165 -1475 17205 -1465
rect 17275 -1440 17315 -1435
rect 17275 -1470 17280 -1440
rect 17310 -1470 17315 -1440
rect 17275 -1475 17315 -1470
rect 17585 -1445 17625 -1435
rect 17585 -1465 17595 -1445
rect 17615 -1465 17625 -1445
rect 17585 -1475 17625 -1465
rect 17670 -1445 17710 -1435
rect 17670 -1465 17680 -1445
rect 17700 -1465 17710 -1445
rect 17670 -1475 17710 -1465
rect 17780 -1440 17820 -1435
rect 17780 -1470 17785 -1440
rect 17815 -1470 17820 -1440
rect 17780 -1475 17820 -1470
rect 17890 -1440 17930 -1435
rect 17890 -1470 17895 -1440
rect 17925 -1470 17930 -1440
rect 17890 -1475 17930 -1470
rect 18000 -1440 18040 -1435
rect 18000 -1470 18005 -1440
rect 18035 -1470 18040 -1440
rect 18000 -1475 18040 -1470
rect 18285 -1440 18325 -1435
rect 18285 -1470 18290 -1440
rect 18320 -1470 18325 -1440
rect 18285 -1475 18325 -1470
rect 18395 -1445 18435 -1435
rect 18395 -1465 18405 -1445
rect 18425 -1465 18435 -1445
rect 18395 -1475 18435 -1465
rect 18505 -1440 18545 -1435
rect 18505 -1470 18510 -1440
rect 18540 -1470 18545 -1440
rect 18505 -1475 18545 -1470
rect 18615 -1445 18655 -1435
rect 18615 -1465 18625 -1445
rect 18645 -1465 18655 -1445
rect 18615 -1475 18655 -1465
rect 16955 -1540 16975 -1475
rect 16945 -1545 16985 -1540
rect 16945 -1575 16950 -1545
rect 16980 -1575 16985 -1545
rect 16945 -1580 16985 -1575
rect 17065 -1585 17085 -1475
rect 17175 -1540 17195 -1475
rect 17165 -1545 17205 -1540
rect 17165 -1575 17170 -1545
rect 17200 -1575 17205 -1545
rect 17165 -1580 17205 -1575
rect 17055 -1590 17095 -1585
rect 17055 -1620 17060 -1590
rect 17090 -1620 17095 -1590
rect 17055 -1625 17095 -1620
rect 17595 -1635 17615 -1475
rect 17585 -1640 17625 -1635
rect 17585 -1670 17590 -1640
rect 17620 -1670 17625 -1640
rect 17585 -1675 17625 -1670
rect 17680 -1680 17700 -1475
rect 17780 -1500 17820 -1495
rect 17780 -1530 17785 -1500
rect 17815 -1530 17820 -1500
rect 17780 -1535 17820 -1530
rect 17670 -1685 17710 -1680
rect 17670 -1715 17675 -1685
rect 17705 -1715 17710 -1685
rect 17670 -1720 17710 -1715
rect 17790 -1805 17810 -1535
rect 17900 -1680 17920 -1475
rect 18405 -1540 18425 -1475
rect 18395 -1545 18435 -1540
rect 18395 -1575 18400 -1545
rect 18430 -1575 18435 -1545
rect 18395 -1580 18435 -1575
rect 18515 -1585 18535 -1475
rect 18625 -1540 18645 -1475
rect 18615 -1545 18655 -1540
rect 18615 -1575 18620 -1545
rect 18650 -1575 18655 -1545
rect 18615 -1580 18655 -1575
rect 18505 -1590 18545 -1585
rect 18505 -1620 18510 -1590
rect 18540 -1620 18545 -1590
rect 18505 -1625 18545 -1620
rect 17890 -1685 17930 -1680
rect 17890 -1715 17895 -1685
rect 17925 -1715 17930 -1685
rect 17890 -1720 17930 -1715
rect 19335 -1755 19355 -405
rect 19325 -1760 19365 -1755
rect 19325 -1790 19330 -1760
rect 19360 -1790 19365 -1760
rect 19325 -1795 19365 -1790
rect 17780 -1810 17820 -1805
rect 17780 -1840 17785 -1810
rect 17815 -1840 17820 -1810
rect 17780 -1845 17820 -1840
rect 16260 -1895 16300 -1890
rect 16260 -1925 16265 -1895
rect 16295 -1925 16300 -1895
rect 16260 -1930 16300 -1925
rect 16480 -1895 16520 -1890
rect 16480 -1925 16485 -1895
rect 16515 -1925 16520 -1895
rect 16480 -1930 16520 -1925
rect 16730 -1895 16770 -1890
rect 16730 -1925 16735 -1895
rect 16765 -1925 16770 -1895
rect 16730 -1930 16770 -1925
rect 17195 -1895 17235 -1890
rect 17195 -1925 17200 -1895
rect 17230 -1925 17235 -1895
rect 17195 -1930 17235 -1925
rect 17425 -1930 17430 -1895
rect 17465 -1930 17470 -1895
rect 18124 -1930 18129 -1895
rect 18164 -1930 18169 -1895
rect 19080 -1900 19120 -1895
rect 19080 -1930 19085 -1900
rect 19115 -1930 19120 -1900
rect 16490 -2895 16510 -1930
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16740 -3100 16760 -1930
rect 17205 -2010 17225 -1930
rect 19080 -1935 19120 -1930
rect 17195 -2015 17235 -2010
rect 17195 -2045 17200 -2015
rect 17230 -2045 17235 -2015
rect 17195 -2050 17235 -2045
rect 18830 -2015 18870 -2010
rect 18830 -2045 18835 -2015
rect 18865 -2045 18870 -2015
rect 18830 -2050 18870 -2045
rect 16945 -2615 18655 -2265
rect 16730 -3105 16770 -3100
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -3150 15860 -3145
rect 15950 -3116 15985 -3111
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 15830 -4260 15850 -3150
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18840 -3100 18860 -2050
rect 19090 -2895 19110 -1935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19415 -2987 19435 -240
rect 19470 -1895 19490 410
rect 19545 -1680 19565 1600
rect 19610 250 19650 255
rect 19610 220 19615 250
rect 19645 220 19650 250
rect 19610 215 19650 220
rect 19535 -1685 19575 -1680
rect 19535 -1715 19540 -1685
rect 19570 -1715 19575 -1685
rect 19535 -1720 19575 -1715
rect 19460 -1900 19500 -1895
rect 19460 -1930 19465 -1900
rect 19495 -1930 19500 -1900
rect 19460 -1935 19500 -1930
rect 19405 -2992 19440 -2987
rect 19405 -3032 19440 -3027
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -3100
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 19620 -3111 19640 215
rect 19730 -105 19770 -100
rect 19730 -135 19735 -105
rect 19765 -135 19770 -105
rect 19730 -140 19770 -135
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4295 15860 -4265
rect 15820 -4300 15860 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4345 15765 -4315
rect 15725 -4350 15765 -4345
rect 15960 -4355 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4185 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 16605 -4009 16640 -4004
rect 18960 -4009 18995 -4004
rect 16540 -4035 16580 -4030
rect 16540 -4065 16545 -4035
rect 16575 -4065 16580 -4035
rect 16540 -4070 16580 -4065
rect 16550 -4185 16570 -4070
rect 16615 -4185 16635 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16540 -4190 16580 -4185
rect 16540 -4220 16545 -4190
rect 16575 -4220 16580 -4190
rect 16540 -4225 16580 -4220
rect 16605 -4190 16645 -4185
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17250 -4265 17300 -4255
rect 18965 -4260 18985 -4009
rect 19290 -4260 19310 -3934
rect 17250 -4295 17260 -4265
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4295 17820 -4265
rect 17780 -4300 17820 -4295
rect 18955 -4265 18995 -4260
rect 18955 -4295 18960 -4265
rect 18990 -4295 18995 -4265
rect 18955 -4300 18995 -4295
rect 19280 -4265 19320 -4260
rect 19280 -4295 19285 -4265
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 16900 -4315 16950 -4305
rect 16900 -4345 16910 -4315
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4345 18700 -4315
rect 18650 -4355 18700 -4345
rect 19620 -4355 19640 -3829
rect 19740 -4310 19760 -140
rect 19785 -1585 19805 1595
rect 19775 -1590 19815 -1585
rect 19775 -1620 19780 -1590
rect 19810 -1620 19815 -1590
rect 19775 -1625 19815 -1620
rect 19730 -4315 19770 -4310
rect 19730 -4345 19735 -4315
rect 19765 -4345 19770 -4315
rect 19730 -4350 19770 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4390 15990 -4360
rect 15950 -4395 15990 -4390
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 19355 -4395 19395 -4390
rect 19610 -4360 19650 -4355
rect 19610 -4390 19615 -4360
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4445 17995 -4440
<< via1 >>
rect 15730 -135 15760 -105
rect 15955 95 15985 125
rect 15790 -1620 15820 -1590
rect 16035 -1575 16065 -1545
rect 17090 1355 17120 1385
rect 16395 1310 16425 1340
rect 16980 1310 17010 1340
rect 18480 1355 18510 1385
rect 17840 1310 17870 1340
rect 18235 1310 18265 1340
rect 16245 1275 16275 1280
rect 16245 1255 16250 1275
rect 16250 1255 16270 1275
rect 16270 1255 16275 1275
rect 16245 1250 16275 1255
rect 16340 1275 16370 1280
rect 16340 1255 16345 1275
rect 16345 1255 16365 1275
rect 16365 1255 16370 1275
rect 16340 1250 16370 1255
rect 16465 1275 16495 1280
rect 16465 1255 16470 1275
rect 16470 1255 16490 1275
rect 16490 1255 16495 1275
rect 16465 1250 16495 1255
rect 16815 1275 16845 1280
rect 16815 1255 16820 1275
rect 16820 1255 16840 1275
rect 16840 1255 16845 1275
rect 16815 1250 16845 1255
rect 16925 1275 16955 1280
rect 16925 1255 16930 1275
rect 16930 1255 16950 1275
rect 16950 1255 16955 1275
rect 16925 1250 16955 1255
rect 17035 1275 17065 1280
rect 17035 1255 17040 1275
rect 17040 1255 17060 1275
rect 17060 1255 17065 1275
rect 17035 1250 17065 1255
rect 17145 1275 17175 1280
rect 17145 1255 17150 1275
rect 17150 1255 17170 1275
rect 17170 1255 17175 1275
rect 17145 1250 17175 1255
rect 17610 1275 17640 1280
rect 17610 1255 17615 1275
rect 17615 1255 17635 1275
rect 17635 1255 17640 1275
rect 17610 1250 17640 1255
rect 17675 1275 17705 1280
rect 17675 1255 17680 1275
rect 17680 1255 17700 1275
rect 17700 1255 17705 1275
rect 17675 1250 17705 1255
rect 17785 1275 17815 1280
rect 17785 1255 17790 1275
rect 17790 1255 17810 1275
rect 17810 1255 17815 1275
rect 17785 1250 17815 1255
rect 17895 1275 17925 1280
rect 17895 1255 17900 1275
rect 17900 1255 17920 1275
rect 17920 1255 17925 1275
rect 17895 1250 17925 1255
rect 17960 1275 17990 1280
rect 17960 1255 17965 1275
rect 17965 1255 17985 1275
rect 17985 1255 17990 1275
rect 17960 1250 17990 1255
rect 16870 1105 16900 1110
rect 16870 1085 16875 1105
rect 16875 1085 16895 1105
rect 16895 1085 16900 1105
rect 16870 1080 16900 1085
rect 16980 1105 17010 1110
rect 16980 1085 16985 1105
rect 16985 1085 17005 1105
rect 17005 1085 17010 1105
rect 16980 1080 17010 1085
rect 17090 1105 17120 1110
rect 17090 1085 17095 1105
rect 17095 1085 17115 1105
rect 17115 1085 17120 1105
rect 17090 1080 17120 1085
rect 17730 1005 17760 1010
rect 17730 985 17735 1005
rect 17735 985 17755 1005
rect 17755 985 17760 1005
rect 17730 980 17760 985
rect 17840 1005 17870 1010
rect 17840 985 17845 1005
rect 17845 985 17865 1005
rect 17865 985 17870 1005
rect 17840 980 17870 985
rect 18590 1310 18620 1340
rect 18425 1275 18455 1280
rect 18425 1255 18430 1275
rect 18430 1255 18450 1275
rect 18450 1255 18455 1275
rect 18425 1250 18455 1255
rect 18535 1275 18565 1280
rect 18535 1255 18540 1275
rect 18540 1255 18560 1275
rect 18560 1255 18565 1275
rect 18535 1250 18565 1255
rect 18645 1275 18675 1280
rect 18645 1255 18650 1275
rect 18650 1255 18670 1275
rect 18670 1255 18675 1275
rect 18645 1250 18675 1255
rect 18755 1275 18785 1280
rect 18755 1255 18760 1275
rect 18760 1255 18780 1275
rect 18780 1255 18785 1275
rect 18755 1250 18785 1255
rect 18480 1105 18510 1110
rect 18480 1085 18485 1105
rect 18485 1085 18505 1105
rect 18505 1085 18510 1105
rect 18480 1080 18510 1085
rect 18590 1105 18620 1110
rect 18590 1085 18595 1105
rect 18595 1085 18615 1105
rect 18615 1085 18620 1105
rect 18590 1080 18620 1085
rect 18700 1105 18730 1110
rect 18700 1085 18705 1105
rect 18705 1085 18725 1105
rect 18725 1085 18730 1105
rect 18700 1080 18730 1085
rect 18235 965 18265 995
rect 18725 965 18755 995
rect 16165 885 16195 915
rect 16300 885 16330 915
rect 16410 885 16440 915
rect 16440 775 16470 805
rect 16660 775 16690 805
rect 16975 810 17005 815
rect 16975 790 16980 810
rect 16980 790 17000 810
rect 17000 790 17005 810
rect 16975 785 17005 790
rect 17155 810 17185 815
rect 17155 790 17160 810
rect 17160 790 17180 810
rect 17180 790 17185 810
rect 17155 785 17185 790
rect 17335 810 17365 815
rect 17335 790 17340 810
rect 17340 790 17360 810
rect 17360 790 17365 810
rect 17335 785 17365 790
rect 17515 810 17545 815
rect 17515 790 17520 810
rect 17520 790 17540 810
rect 17540 790 17545 810
rect 17515 785 17545 790
rect 17695 810 17725 815
rect 17695 790 17700 810
rect 17700 790 17720 810
rect 17720 790 17725 810
rect 17695 785 17725 790
rect 17875 810 17905 815
rect 17875 790 17880 810
rect 17880 790 17900 810
rect 17900 790 17905 810
rect 17875 785 17905 790
rect 18055 810 18085 815
rect 18055 790 18060 810
rect 18060 790 18080 810
rect 18080 790 18085 810
rect 18055 785 18085 790
rect 18235 810 18265 815
rect 18235 790 18240 810
rect 18240 790 18260 810
rect 18260 790 18265 810
rect 18235 785 18265 790
rect 18415 810 18445 815
rect 18415 790 18420 810
rect 18420 790 18440 810
rect 18440 790 18445 810
rect 18415 785 18445 790
rect 18595 810 18625 815
rect 18595 790 18600 810
rect 18600 790 18620 810
rect 18620 790 18625 810
rect 18595 785 18625 790
rect 16550 710 16580 715
rect 16550 690 16555 710
rect 16555 690 16575 710
rect 16575 690 16580 710
rect 16550 685 16580 690
rect 16785 685 16815 715
rect 16485 540 16515 545
rect 16485 520 16490 540
rect 16490 520 16510 540
rect 16510 520 16515 540
rect 16485 515 16515 520
rect 16615 540 16645 545
rect 16615 520 16620 540
rect 16620 520 16640 540
rect 16640 520 16645 540
rect 16615 515 16645 520
rect 16310 415 16340 445
rect 16265 360 16295 390
rect 16210 315 16240 345
rect 16265 -235 16295 -205
rect 16210 -1110 16240 -1080
rect 16165 -1670 16195 -1640
rect 16110 -1715 16140 -1685
rect 16160 -1790 16190 -1760
rect 16845 515 16875 545
rect 16785 360 16815 390
rect 16550 315 16580 345
rect 16425 155 16455 185
rect 16545 155 16575 185
rect 16665 155 16695 185
rect 16785 155 16815 185
rect 17605 440 17635 445
rect 17605 420 17610 440
rect 17610 420 17630 440
rect 17630 420 17635 440
rect 17605 415 17635 420
rect 17965 440 17995 445
rect 17965 420 17970 440
rect 17970 420 17990 440
rect 17990 420 17995 440
rect 17965 415 17995 420
rect 17425 360 17455 390
rect 17245 315 17275 345
rect 17065 270 17095 300
rect 16905 155 16935 185
rect 17025 155 17055 185
rect 17145 155 17175 185
rect 17265 155 17295 185
rect 17385 155 17415 185
rect 17505 155 17535 185
rect 17625 155 17655 185
rect 18145 360 18175 390
rect 18325 315 18355 345
rect 17785 270 17815 300
rect 18505 270 18535 300
rect 19015 795 19045 825
rect 18950 760 18980 765
rect 18950 740 18955 760
rect 18955 740 18975 760
rect 18975 740 18980 760
rect 18950 735 18980 740
rect 19015 760 19045 765
rect 19015 740 19020 760
rect 19020 740 19040 760
rect 19040 740 19045 760
rect 19015 735 19045 740
rect 19125 760 19155 765
rect 19125 740 19130 760
rect 19130 740 19150 760
rect 19150 740 19155 760
rect 19125 735 19155 740
rect 19330 885 19360 915
rect 19085 490 19115 495
rect 19085 470 19090 490
rect 19090 470 19110 490
rect 19110 470 19115 490
rect 19085 465 19115 470
rect 19265 465 19295 495
rect 18005 220 18035 250
rect 18725 220 18755 250
rect 19030 220 19060 250
rect 17945 155 17975 185
rect 18065 155 18095 185
rect 18185 155 18215 185
rect 18305 155 18335 185
rect 18425 155 18455 185
rect 18545 155 18575 185
rect 18665 155 18695 185
rect 18785 155 18815 185
rect 18905 155 18935 185
rect 19025 155 19055 185
rect 19145 155 19175 185
rect 16485 120 16515 125
rect 16485 100 16490 120
rect 16490 100 16510 120
rect 16510 100 16515 120
rect 16485 95 16515 100
rect 16845 120 16875 125
rect 16845 100 16850 120
rect 16850 100 16870 120
rect 16870 100 16875 120
rect 16845 95 16875 100
rect 17205 120 17235 125
rect 17205 100 17210 120
rect 17210 100 17230 120
rect 17230 100 17235 120
rect 17205 95 17235 100
rect 17565 120 17595 125
rect 17565 100 17570 120
rect 17570 100 17590 120
rect 17590 100 17595 120
rect 17565 95 17595 100
rect 17695 95 17725 125
rect 17875 95 17905 125
rect 16605 -50 16635 -45
rect 16605 -70 16610 -50
rect 16610 -70 16630 -50
rect 16630 -70 16635 -50
rect 16605 -75 16635 -70
rect 16965 -50 16995 -45
rect 16965 -70 16970 -50
rect 16970 -70 16990 -50
rect 16990 -70 16995 -50
rect 16965 -75 16995 -70
rect 17325 -50 17355 -45
rect 17325 -70 17330 -50
rect 17330 -70 17350 -50
rect 17350 -70 17355 -50
rect 17325 -75 17355 -70
rect 16515 -135 16545 -105
rect 16725 -135 16755 -105
rect 16845 -135 16875 -105
rect 17085 -135 17115 -105
rect 17205 -135 17235 -105
rect 17445 -135 17475 -105
rect 17535 -135 17565 -105
rect 16915 -210 16945 -205
rect 16915 -230 16920 -210
rect 16920 -230 16940 -210
rect 16940 -230 16945 -210
rect 16915 -235 16945 -230
rect 16975 -220 17005 -190
rect 17215 -220 17245 -190
rect 17455 -220 17485 -190
rect 16855 -255 16885 -250
rect 16855 -275 16860 -255
rect 16860 -275 16880 -255
rect 16880 -275 16885 -255
rect 16855 -280 16885 -275
rect 17095 -255 17125 -250
rect 17095 -275 17100 -255
rect 17100 -275 17120 -255
rect 17120 -275 17125 -255
rect 17095 -280 17125 -275
rect 17335 -255 17365 -250
rect 17335 -275 17340 -255
rect 17340 -275 17360 -255
rect 17360 -275 17365 -255
rect 17335 -280 17365 -275
rect 17565 -315 17595 -310
rect 17565 -335 17570 -315
rect 17570 -335 17590 -315
rect 17590 -335 17595 -315
rect 17565 -340 17595 -335
rect 16310 -400 16340 -370
rect 16855 -375 16885 -370
rect 16855 -395 16860 -375
rect 16860 -395 16880 -375
rect 16880 -395 16885 -375
rect 16855 -400 16885 -395
rect 16535 -460 16565 -430
rect 16915 -460 16945 -430
rect 17035 -460 17065 -430
rect 17155 -460 17185 -430
rect 17275 -460 17305 -430
rect 17395 -460 17425 -430
rect 16625 -535 16655 -530
rect 16625 -555 16630 -535
rect 16630 -555 16650 -535
rect 16650 -555 16655 -535
rect 16625 -560 16655 -555
rect 16745 -535 16775 -530
rect 16745 -555 16750 -535
rect 16750 -555 16770 -535
rect 16770 -555 16775 -535
rect 16745 -560 16775 -555
rect 16865 -535 16895 -530
rect 16865 -555 16870 -535
rect 16870 -555 16890 -535
rect 16890 -555 16895 -535
rect 16865 -560 16895 -555
rect 16985 -535 17015 -530
rect 16985 -555 16990 -535
rect 16990 -555 17010 -535
rect 17010 -555 17015 -535
rect 16985 -560 17015 -555
rect 17305 -535 17335 -530
rect 17305 -555 17310 -535
rect 17310 -555 17330 -535
rect 17330 -555 17335 -535
rect 17305 -560 17335 -555
rect 17425 -535 17455 -530
rect 17425 -555 17430 -535
rect 17430 -555 17450 -535
rect 17450 -555 17455 -535
rect 17425 -560 17455 -555
rect 17545 -535 17575 -530
rect 17545 -555 17550 -535
rect 17550 -555 17570 -535
rect 17570 -555 17575 -535
rect 17545 -560 17575 -555
rect 17785 -340 17815 -310
rect 18005 120 18035 125
rect 18005 100 18010 120
rect 18010 100 18030 120
rect 18030 100 18035 120
rect 18005 95 18035 100
rect 18365 120 18395 125
rect 18365 100 18370 120
rect 18370 100 18390 120
rect 18390 100 18395 120
rect 18365 95 18395 100
rect 18725 120 18755 125
rect 18725 100 18730 120
rect 18730 100 18750 120
rect 18750 100 18755 120
rect 18725 95 18755 100
rect 19085 120 19115 125
rect 19085 100 19090 120
rect 19090 100 19110 120
rect 19110 100 19115 120
rect 19085 95 19115 100
rect 18245 -50 18275 -45
rect 18245 -70 18250 -50
rect 18250 -70 18270 -50
rect 18270 -70 18275 -50
rect 18245 -75 18275 -70
rect 18605 -50 18635 -45
rect 18605 -70 18610 -50
rect 18610 -70 18630 -50
rect 18630 -70 18635 -50
rect 18605 -75 18635 -70
rect 18965 -50 18995 -45
rect 18965 -70 18970 -50
rect 18970 -70 18990 -50
rect 18990 -70 18995 -50
rect 18965 -75 18995 -70
rect 18035 -135 18065 -105
rect 18125 -135 18155 -105
rect 18365 -135 18395 -105
rect 18485 -135 18515 -105
rect 18115 -220 18145 -190
rect 18355 -220 18385 -190
rect 18725 -135 18755 -105
rect 18845 -135 18875 -105
rect 19055 -135 19085 -105
rect 18595 -220 18625 -190
rect 18655 -210 18685 -205
rect 18655 -230 18660 -210
rect 18660 -230 18680 -210
rect 18680 -230 18685 -210
rect 18655 -235 18685 -230
rect 18235 -255 18265 -250
rect 18235 -275 18240 -255
rect 18240 -275 18260 -255
rect 18260 -275 18265 -255
rect 18235 -280 18265 -275
rect 18475 -255 18505 -250
rect 18475 -275 18480 -255
rect 18480 -275 18500 -255
rect 18500 -275 18505 -255
rect 18475 -280 18505 -275
rect 18715 -255 18745 -250
rect 18715 -275 18720 -255
rect 18720 -275 18740 -255
rect 18740 -275 18745 -255
rect 18715 -280 18745 -275
rect 18005 -315 18035 -310
rect 18005 -335 18010 -315
rect 18010 -335 18030 -315
rect 18030 -335 18035 -315
rect 18005 -340 18035 -335
rect 19465 415 19495 445
rect 19410 270 19440 300
rect 19410 -235 19440 -205
rect 18715 -375 18745 -370
rect 18715 -395 18720 -375
rect 18720 -395 18740 -375
rect 18740 -395 18745 -375
rect 18715 -400 18745 -395
rect 19330 -400 19360 -370
rect 18175 -460 18205 -430
rect 18295 -460 18325 -430
rect 18415 -460 18445 -430
rect 18535 -460 18565 -430
rect 18655 -460 18685 -430
rect 19035 -460 19065 -430
rect 18025 -535 18055 -530
rect 18025 -555 18030 -535
rect 18030 -555 18050 -535
rect 18050 -555 18055 -535
rect 18025 -560 18055 -555
rect 18145 -535 18175 -530
rect 18145 -555 18150 -535
rect 18150 -555 18170 -535
rect 18170 -555 18175 -535
rect 18145 -560 18175 -555
rect 18265 -535 18295 -530
rect 18265 -555 18270 -535
rect 18270 -555 18290 -535
rect 18290 -555 18295 -535
rect 18265 -560 18295 -555
rect 18585 -535 18615 -530
rect 18585 -555 18590 -535
rect 18590 -555 18610 -535
rect 18610 -555 18615 -535
rect 18585 -560 18615 -555
rect 18705 -535 18735 -530
rect 18705 -555 18710 -535
rect 18710 -555 18730 -535
rect 18730 -555 18735 -535
rect 18705 -560 18735 -555
rect 18825 -535 18855 -530
rect 18825 -555 18830 -535
rect 18830 -555 18850 -535
rect 18850 -555 18855 -535
rect 18825 -560 18855 -555
rect 18945 -535 18975 -530
rect 18945 -555 18950 -535
rect 18950 -555 18970 -535
rect 18970 -555 18975 -535
rect 18945 -560 18975 -555
rect 17115 -850 17145 -845
rect 17115 -870 17120 -850
rect 17120 -870 17140 -850
rect 17140 -870 17145 -850
rect 17115 -875 17145 -870
rect 17785 -875 17815 -845
rect 18455 -850 18485 -845
rect 18455 -870 18460 -850
rect 18460 -870 18480 -850
rect 18480 -870 18485 -850
rect 18455 -875 18485 -870
rect 16745 -1000 16775 -995
rect 16745 -1020 16750 -1000
rect 16750 -1020 16770 -1000
rect 16770 -1020 16775 -1000
rect 16745 -1025 16775 -1020
rect 16825 -1000 16855 -995
rect 16825 -1020 16830 -1000
rect 16830 -1020 16850 -1000
rect 16850 -1020 16855 -1000
rect 16825 -1025 16855 -1020
rect 16905 -1000 16935 -995
rect 16905 -1020 16910 -1000
rect 16910 -1020 16930 -1000
rect 16930 -1020 16935 -1000
rect 16905 -1025 16935 -1020
rect 16985 -1000 17015 -995
rect 16985 -1020 16990 -1000
rect 16990 -1020 17010 -1000
rect 17010 -1020 17015 -1000
rect 16985 -1025 17015 -1020
rect 17065 -1000 17095 -995
rect 17065 -1020 17070 -1000
rect 17070 -1020 17090 -1000
rect 17090 -1020 17095 -1000
rect 17065 -1025 17095 -1020
rect 17145 -1000 17175 -995
rect 17145 -1020 17150 -1000
rect 17150 -1020 17170 -1000
rect 17170 -1020 17175 -1000
rect 17145 -1025 17175 -1020
rect 17225 -1000 17255 -995
rect 17225 -1020 17230 -1000
rect 17230 -1020 17250 -1000
rect 17250 -1020 17255 -1000
rect 17225 -1025 17255 -1020
rect 17305 -1000 17335 -995
rect 17305 -1020 17310 -1000
rect 17310 -1020 17330 -1000
rect 17330 -1020 17335 -1000
rect 17305 -1025 17335 -1020
rect 17385 -1000 17415 -995
rect 17385 -1020 17390 -1000
rect 17390 -1020 17410 -1000
rect 17410 -1020 17415 -1000
rect 17385 -1025 17415 -1020
rect 17465 -1000 17495 -995
rect 17465 -1020 17470 -1000
rect 17470 -1020 17490 -1000
rect 17490 -1020 17495 -1000
rect 17465 -1025 17495 -1020
rect 17545 -1000 17575 -995
rect 17545 -1020 17550 -1000
rect 17550 -1020 17570 -1000
rect 17570 -1020 17575 -1000
rect 17545 -1025 17575 -1020
rect 17625 -1000 17655 -995
rect 17625 -1020 17630 -1000
rect 17630 -1020 17650 -1000
rect 17650 -1020 17655 -1000
rect 17625 -1025 17655 -1020
rect 17705 -1000 17735 -995
rect 17705 -1020 17710 -1000
rect 17710 -1020 17730 -1000
rect 17730 -1020 17735 -1000
rect 17705 -1025 17735 -1020
rect 17785 -1000 17815 -995
rect 17785 -1020 17790 -1000
rect 17790 -1020 17810 -1000
rect 17810 -1020 17815 -1000
rect 17785 -1025 17815 -1020
rect 17865 -1000 17895 -995
rect 17865 -1020 17870 -1000
rect 17870 -1020 17890 -1000
rect 17890 -1020 17895 -1000
rect 17865 -1025 17895 -1020
rect 17945 -1000 17975 -995
rect 17945 -1020 17950 -1000
rect 17950 -1020 17970 -1000
rect 17970 -1020 17975 -1000
rect 17945 -1025 17975 -1020
rect 18025 -1000 18055 -995
rect 18025 -1020 18030 -1000
rect 18030 -1020 18050 -1000
rect 18050 -1020 18055 -1000
rect 18025 -1025 18055 -1020
rect 18105 -1000 18135 -995
rect 18105 -1020 18110 -1000
rect 18110 -1020 18130 -1000
rect 18130 -1020 18135 -1000
rect 18105 -1025 18135 -1020
rect 18185 -1000 18215 -995
rect 18185 -1020 18190 -1000
rect 18190 -1020 18210 -1000
rect 18210 -1020 18215 -1000
rect 18185 -1025 18215 -1020
rect 18265 -1000 18295 -995
rect 18265 -1020 18270 -1000
rect 18270 -1020 18290 -1000
rect 18290 -1020 18295 -1000
rect 18265 -1025 18295 -1020
rect 18345 -1000 18375 -995
rect 18345 -1020 18350 -1000
rect 18350 -1020 18370 -1000
rect 18370 -1020 18375 -1000
rect 18345 -1025 18375 -1020
rect 18425 -1000 18455 -995
rect 18425 -1020 18430 -1000
rect 18430 -1020 18450 -1000
rect 18450 -1020 18455 -1000
rect 18425 -1025 18455 -1020
rect 18505 -1000 18535 -995
rect 18505 -1020 18510 -1000
rect 18510 -1020 18530 -1000
rect 18530 -1020 18535 -1000
rect 18505 -1025 18535 -1020
rect 18585 -1000 18615 -995
rect 18585 -1020 18590 -1000
rect 18590 -1020 18610 -1000
rect 18610 -1020 18615 -1000
rect 18585 -1025 18615 -1020
rect 18665 -1000 18695 -995
rect 18665 -1020 18670 -1000
rect 18670 -1020 18690 -1000
rect 18690 -1020 18695 -1000
rect 18665 -1025 18695 -1020
rect 18745 -1000 18775 -995
rect 18745 -1020 18750 -1000
rect 18750 -1020 18770 -1000
rect 18770 -1020 18775 -1000
rect 18745 -1025 18775 -1020
rect 16705 -1085 16735 -1080
rect 16705 -1105 16710 -1085
rect 16710 -1105 16730 -1085
rect 16730 -1105 16735 -1085
rect 16705 -1110 16735 -1105
rect 18900 -1085 18930 -1080
rect 18900 -1105 18905 -1085
rect 18905 -1105 18925 -1085
rect 18925 -1105 18930 -1085
rect 18900 -1110 18930 -1105
rect 17170 -1230 17200 -1200
rect 17785 -1230 17815 -1200
rect 18400 -1230 18430 -1200
rect 16895 -1275 16925 -1270
rect 16895 -1295 16900 -1275
rect 16900 -1295 16920 -1275
rect 16920 -1295 16925 -1275
rect 16895 -1300 16925 -1295
rect 17005 -1275 17035 -1270
rect 17005 -1295 17010 -1275
rect 17010 -1295 17030 -1275
rect 17030 -1295 17035 -1275
rect 17005 -1300 17035 -1295
rect 17115 -1275 17145 -1270
rect 17115 -1295 17120 -1275
rect 17120 -1295 17140 -1275
rect 17140 -1295 17145 -1275
rect 17115 -1300 17145 -1295
rect 17225 -1275 17255 -1270
rect 17225 -1295 17230 -1275
rect 17230 -1295 17250 -1275
rect 17250 -1295 17255 -1275
rect 17225 -1300 17255 -1295
rect 17335 -1275 17365 -1270
rect 17335 -1295 17340 -1275
rect 17340 -1295 17360 -1275
rect 17360 -1295 17365 -1275
rect 17335 -1300 17365 -1295
rect 17510 -1275 17540 -1270
rect 17510 -1295 17515 -1275
rect 17515 -1295 17535 -1275
rect 17535 -1295 17540 -1275
rect 17510 -1300 17540 -1295
rect 17620 -1275 17650 -1270
rect 17620 -1295 17625 -1275
rect 17625 -1295 17645 -1275
rect 17645 -1295 17650 -1275
rect 17620 -1300 17650 -1295
rect 17730 -1275 17760 -1270
rect 17730 -1295 17735 -1275
rect 17735 -1295 17755 -1275
rect 17755 -1295 17760 -1275
rect 17730 -1300 17760 -1295
rect 17840 -1275 17870 -1270
rect 17840 -1295 17845 -1275
rect 17845 -1295 17865 -1275
rect 17865 -1295 17870 -1275
rect 17840 -1300 17870 -1295
rect 17950 -1275 17980 -1270
rect 17950 -1295 17955 -1275
rect 17955 -1295 17975 -1275
rect 17975 -1295 17980 -1275
rect 17950 -1300 17980 -1295
rect 18060 -1275 18090 -1270
rect 18060 -1295 18065 -1275
rect 18065 -1295 18085 -1275
rect 18085 -1295 18090 -1275
rect 18060 -1300 18090 -1295
rect 18235 -1275 18265 -1270
rect 18235 -1295 18240 -1275
rect 18240 -1295 18260 -1275
rect 18260 -1295 18265 -1275
rect 18235 -1300 18265 -1295
rect 18345 -1275 18375 -1270
rect 18345 -1295 18350 -1275
rect 18350 -1295 18370 -1275
rect 18370 -1295 18375 -1275
rect 18345 -1300 18375 -1295
rect 18455 -1275 18485 -1270
rect 18455 -1295 18460 -1275
rect 18460 -1295 18480 -1275
rect 18480 -1295 18485 -1275
rect 18455 -1300 18485 -1295
rect 18565 -1275 18595 -1270
rect 18565 -1295 18570 -1275
rect 18570 -1295 18590 -1275
rect 18590 -1295 18595 -1275
rect 18565 -1300 18595 -1295
rect 18675 -1275 18705 -1270
rect 18675 -1295 18680 -1275
rect 18680 -1295 18700 -1275
rect 18700 -1295 18705 -1275
rect 18675 -1300 18705 -1295
rect 17060 -1445 17090 -1440
rect 17060 -1465 17065 -1445
rect 17065 -1465 17085 -1445
rect 17085 -1465 17090 -1445
rect 17060 -1470 17090 -1465
rect 17280 -1445 17310 -1440
rect 17280 -1465 17285 -1445
rect 17285 -1465 17305 -1445
rect 17305 -1465 17310 -1445
rect 17280 -1470 17310 -1465
rect 17785 -1445 17815 -1440
rect 17785 -1465 17790 -1445
rect 17790 -1465 17810 -1445
rect 17810 -1465 17815 -1445
rect 17785 -1470 17815 -1465
rect 17895 -1445 17925 -1440
rect 17895 -1465 17900 -1445
rect 17900 -1465 17920 -1445
rect 17920 -1465 17925 -1445
rect 17895 -1470 17925 -1465
rect 18005 -1445 18035 -1440
rect 18005 -1465 18010 -1445
rect 18010 -1465 18030 -1445
rect 18030 -1465 18035 -1445
rect 18005 -1470 18035 -1465
rect 18290 -1445 18320 -1440
rect 18290 -1465 18295 -1445
rect 18295 -1465 18315 -1445
rect 18315 -1465 18320 -1445
rect 18290 -1470 18320 -1465
rect 18510 -1445 18540 -1440
rect 18510 -1465 18515 -1445
rect 18515 -1465 18535 -1445
rect 18535 -1465 18540 -1445
rect 18510 -1470 18540 -1465
rect 16950 -1575 16980 -1545
rect 17170 -1575 17200 -1545
rect 17060 -1620 17090 -1590
rect 17590 -1670 17620 -1640
rect 17785 -1530 17815 -1500
rect 17675 -1715 17705 -1685
rect 18400 -1575 18430 -1545
rect 18620 -1575 18650 -1545
rect 18510 -1620 18540 -1590
rect 17895 -1715 17925 -1685
rect 19330 -1790 19360 -1760
rect 17785 -1840 17815 -1810
rect 16265 -1925 16295 -1895
rect 16485 -1925 16515 -1895
rect 16735 -1925 16765 -1895
rect 17200 -1925 17230 -1895
rect 17430 -1900 17465 -1895
rect 17430 -1925 17435 -1900
rect 17435 -1925 17460 -1900
rect 17460 -1925 17465 -1900
rect 17430 -1930 17465 -1925
rect 18129 -1900 18164 -1895
rect 18129 -1925 18134 -1900
rect 18134 -1925 18159 -1900
rect 18159 -1925 18164 -1900
rect 18129 -1930 18164 -1925
rect 19085 -1930 19115 -1900
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 17200 -2045 17230 -2015
rect 18835 -2045 18865 -2015
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 220 19645 250
rect 19540 -1715 19570 -1685
rect 19465 -1930 19495 -1900
rect 19405 -2997 19440 -2992
rect 19405 -3022 19410 -2997
rect 19410 -3022 19435 -2997
rect 19435 -3022 19440 -2997
rect 19405 -3027 19440 -3022
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 19735 -135 19765 -105
rect 19610 -3121 19645 -3116
rect 19610 -3146 19615 -3121
rect 19615 -3146 19640 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3151 19645 -3146
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4295 15855 -4265
rect 15730 -4345 15760 -4315
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 16605 -4004 16640 -3999
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 16545 -4065 16575 -4035
rect 16285 -4220 16315 -4190
rect 16545 -4220 16575 -4190
rect 16610 -4220 16640 -4190
rect 17260 -4295 17290 -4265
rect 17785 -4270 17815 -4265
rect 17785 -4290 17790 -4270
rect 17790 -4290 17810 -4270
rect 17810 -4290 17815 -4270
rect 17785 -4295 17815 -4290
rect 18960 -4295 18990 -4265
rect 19285 -4295 19315 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 19780 -1620 19810 -1590
rect 19735 -4345 19765 -4315
rect 15955 -4390 15985 -4360
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 19615 -4390 19645 -4360
rect 17960 -4440 17990 -4410
<< metal2 >>
rect 17085 1385 17125 1390
rect 17085 1355 17090 1385
rect 17120 1355 17125 1385
rect 17085 1350 17125 1355
rect 18475 1385 18515 1390
rect 18475 1355 18480 1385
rect 18510 1355 18515 1385
rect 18475 1350 18515 1355
rect 16390 1340 16430 1345
rect 16390 1310 16395 1340
rect 16425 1335 16430 1340
rect 16975 1340 17015 1345
rect 16975 1335 16980 1340
rect 16425 1315 16980 1335
rect 16425 1310 16430 1315
rect 16390 1305 16430 1310
rect 16975 1310 16980 1315
rect 17010 1335 17015 1340
rect 17835 1340 17875 1345
rect 17835 1335 17840 1340
rect 17010 1315 17840 1335
rect 17010 1310 17015 1315
rect 16975 1305 17015 1310
rect 17835 1310 17840 1315
rect 17870 1335 17875 1340
rect 18230 1340 18270 1345
rect 18230 1335 18235 1340
rect 17870 1315 18235 1335
rect 17870 1310 17875 1315
rect 17835 1305 17875 1310
rect 18230 1310 18235 1315
rect 18265 1335 18270 1340
rect 18585 1340 18625 1345
rect 18585 1335 18590 1340
rect 18265 1315 18590 1335
rect 18265 1310 18270 1315
rect 18230 1305 18270 1310
rect 18585 1310 18590 1315
rect 18620 1310 18625 1340
rect 18585 1305 18625 1310
rect 16240 1280 16280 1285
rect 16240 1250 16245 1280
rect 16275 1275 16280 1280
rect 16335 1280 16375 1285
rect 16335 1275 16340 1280
rect 16275 1255 16340 1275
rect 16275 1250 16280 1255
rect 16240 1245 16280 1250
rect 16335 1250 16340 1255
rect 16370 1275 16375 1280
rect 16460 1280 16500 1285
rect 16460 1275 16465 1280
rect 16370 1255 16465 1275
rect 16370 1250 16375 1255
rect 16335 1245 16375 1250
rect 16460 1250 16465 1255
rect 16495 1275 16500 1280
rect 16810 1280 16850 1285
rect 16810 1275 16815 1280
rect 16495 1255 16815 1275
rect 16495 1250 16500 1255
rect 16460 1245 16500 1250
rect 16810 1250 16815 1255
rect 16845 1275 16850 1280
rect 16920 1280 16960 1285
rect 16920 1275 16925 1280
rect 16845 1255 16925 1275
rect 16845 1250 16850 1255
rect 16810 1245 16850 1250
rect 16920 1250 16925 1255
rect 16955 1275 16960 1280
rect 17030 1280 17070 1285
rect 17030 1275 17035 1280
rect 16955 1255 17035 1275
rect 16955 1250 16960 1255
rect 16920 1245 16960 1250
rect 17030 1250 17035 1255
rect 17065 1275 17070 1280
rect 17140 1280 17180 1285
rect 17140 1275 17145 1280
rect 17065 1255 17145 1275
rect 17065 1250 17070 1255
rect 17030 1245 17070 1250
rect 17140 1250 17145 1255
rect 17175 1275 17180 1280
rect 17605 1280 17645 1285
rect 17605 1275 17610 1280
rect 17175 1255 17610 1275
rect 17175 1250 17180 1255
rect 17140 1245 17180 1250
rect 17605 1250 17610 1255
rect 17640 1275 17645 1280
rect 17670 1280 17710 1285
rect 17670 1275 17675 1280
rect 17640 1255 17675 1275
rect 17640 1250 17645 1255
rect 17605 1245 17645 1250
rect 17670 1250 17675 1255
rect 17705 1275 17710 1280
rect 17780 1280 17820 1285
rect 17780 1275 17785 1280
rect 17705 1255 17785 1275
rect 17705 1250 17710 1255
rect 17670 1245 17710 1250
rect 17780 1250 17785 1255
rect 17815 1275 17820 1280
rect 17890 1280 17930 1285
rect 17890 1275 17895 1280
rect 17815 1255 17895 1275
rect 17815 1250 17820 1255
rect 17780 1245 17820 1250
rect 17890 1250 17895 1255
rect 17925 1275 17930 1280
rect 17955 1280 17995 1285
rect 17955 1275 17960 1280
rect 17925 1255 17960 1275
rect 17925 1250 17930 1255
rect 17890 1245 17930 1250
rect 17955 1250 17960 1255
rect 17990 1275 17995 1280
rect 18420 1280 18460 1285
rect 18420 1275 18425 1280
rect 17990 1255 18425 1275
rect 17990 1250 17995 1255
rect 17955 1245 17995 1250
rect 18420 1250 18425 1255
rect 18455 1275 18460 1280
rect 18530 1280 18570 1285
rect 18530 1275 18535 1280
rect 18455 1255 18535 1275
rect 18455 1250 18460 1255
rect 18420 1245 18460 1250
rect 18530 1250 18535 1255
rect 18565 1275 18570 1280
rect 18640 1280 18680 1285
rect 18640 1275 18645 1280
rect 18565 1255 18645 1275
rect 18565 1250 18570 1255
rect 18530 1245 18570 1250
rect 18640 1250 18645 1255
rect 18675 1275 18680 1280
rect 18750 1280 18790 1285
rect 18750 1275 18755 1280
rect 18675 1255 18755 1275
rect 18675 1250 18680 1255
rect 18640 1245 18680 1250
rect 18750 1250 18755 1255
rect 18785 1275 18790 1280
rect 20050 1280 20090 1285
rect 20050 1275 20055 1280
rect 18785 1255 20055 1275
rect 18785 1250 18790 1255
rect 18750 1245 18790 1250
rect 20050 1250 20055 1255
rect 20085 1250 20090 1280
rect 20050 1245 20090 1250
rect 16865 1110 16905 1115
rect 16865 1080 16870 1110
rect 16900 1105 16905 1110
rect 16975 1110 17015 1115
rect 16975 1105 16980 1110
rect 16900 1085 16980 1105
rect 16900 1080 16905 1085
rect 16865 1075 16905 1080
rect 16975 1080 16980 1085
rect 17010 1105 17015 1110
rect 17085 1110 17125 1115
rect 17085 1105 17090 1110
rect 17010 1085 17090 1105
rect 17010 1080 17015 1085
rect 16975 1075 17015 1080
rect 17085 1080 17090 1085
rect 17120 1080 17125 1110
rect 17085 1075 17125 1080
rect 18475 1110 18515 1115
rect 18475 1080 18480 1110
rect 18510 1105 18515 1110
rect 18585 1110 18625 1115
rect 18585 1105 18590 1110
rect 18510 1085 18590 1105
rect 18510 1080 18515 1085
rect 18475 1075 18515 1080
rect 18585 1080 18590 1085
rect 18620 1105 18625 1110
rect 18695 1110 18735 1115
rect 18695 1105 18700 1110
rect 18620 1085 18700 1105
rect 18620 1080 18625 1085
rect 18585 1075 18625 1080
rect 18695 1080 18700 1085
rect 18730 1080 18735 1110
rect 18695 1075 18735 1080
rect 17725 1010 17765 1015
rect 17725 980 17730 1010
rect 17760 1005 17765 1010
rect 17835 1010 17875 1015
rect 17835 1005 17840 1010
rect 17760 985 17840 1005
rect 17760 980 17765 985
rect 17725 975 17765 980
rect 17835 980 17840 985
rect 17870 980 17875 1010
rect 17835 975 17875 980
rect 18230 995 18270 1000
rect 18230 965 18235 995
rect 18265 990 18270 995
rect 18720 995 18760 1000
rect 18720 990 18725 995
rect 18265 970 18725 990
rect 18265 965 18270 970
rect 18230 960 18270 965
rect 18720 965 18725 970
rect 18755 965 18760 995
rect 18720 960 18760 965
rect 16160 915 16200 920
rect 16160 885 16165 915
rect 16195 910 16200 915
rect 16295 915 16335 920
rect 16295 910 16300 915
rect 16195 890 16300 910
rect 16195 885 16200 890
rect 16160 880 16200 885
rect 16295 885 16300 890
rect 16330 885 16335 915
rect 16295 880 16335 885
rect 16405 915 16445 920
rect 16405 885 16410 915
rect 16440 910 16445 915
rect 19325 915 19365 920
rect 19325 910 19330 915
rect 16440 890 19330 910
rect 16440 885 16445 890
rect 16405 880 16445 885
rect 19325 885 19330 890
rect 19360 885 19365 915
rect 19325 880 19365 885
rect 19010 825 19050 830
rect 16970 815 17010 820
rect 16435 805 16475 810
rect 16435 775 16440 805
rect 16470 800 16475 805
rect 16655 805 16695 810
rect 16655 800 16660 805
rect 16470 780 16660 800
rect 16470 775 16475 780
rect 16435 770 16475 775
rect 16655 775 16660 780
rect 16690 800 16695 805
rect 16970 800 16975 815
rect 16690 785 16975 800
rect 17005 810 17010 815
rect 17150 815 17190 820
rect 17150 810 17155 815
rect 17005 790 17155 810
rect 17005 785 17010 790
rect 16690 780 17010 785
rect 17150 785 17155 790
rect 17185 810 17190 815
rect 17330 815 17370 820
rect 17330 810 17335 815
rect 17185 790 17335 810
rect 17185 785 17190 790
rect 17150 780 17190 785
rect 17330 785 17335 790
rect 17365 810 17370 815
rect 17510 815 17550 820
rect 17510 810 17515 815
rect 17365 790 17515 810
rect 17365 785 17370 790
rect 17330 780 17370 785
rect 17510 785 17515 790
rect 17545 810 17550 815
rect 17690 815 17730 820
rect 17690 810 17695 815
rect 17545 790 17695 810
rect 17545 785 17550 790
rect 17510 780 17550 785
rect 17690 785 17695 790
rect 17725 810 17730 815
rect 17870 815 17910 820
rect 17870 810 17875 815
rect 17725 790 17875 810
rect 17725 785 17730 790
rect 17690 780 17730 785
rect 17870 785 17875 790
rect 17905 810 17910 815
rect 18050 815 18090 820
rect 18050 810 18055 815
rect 17905 790 18055 810
rect 17905 785 17910 790
rect 17870 780 17910 785
rect 18050 785 18055 790
rect 18085 810 18090 815
rect 18230 815 18270 820
rect 18230 810 18235 815
rect 18085 790 18235 810
rect 18085 785 18090 790
rect 18050 780 18090 785
rect 18230 785 18235 790
rect 18265 810 18270 815
rect 18410 815 18450 820
rect 18410 810 18415 815
rect 18265 790 18415 810
rect 18265 785 18270 790
rect 18230 780 18270 785
rect 18410 785 18415 790
rect 18445 810 18450 815
rect 18590 815 18630 820
rect 18590 810 18595 815
rect 18445 790 18595 810
rect 18445 785 18450 790
rect 18410 780 18450 785
rect 18590 785 18595 790
rect 18625 810 18630 815
rect 19010 810 19015 825
rect 18625 795 19015 810
rect 19045 810 19050 825
rect 20050 815 20090 820
rect 20050 810 20055 815
rect 19045 795 20055 810
rect 18625 790 20055 795
rect 18625 785 18630 790
rect 18590 780 18630 785
rect 20050 785 20055 790
rect 20085 785 20090 815
rect 20050 780 20090 785
rect 16690 775 16695 780
rect 16655 770 16695 775
rect 18945 765 18985 770
rect 18945 735 18950 765
rect 18980 760 18985 765
rect 19010 765 19050 770
rect 19010 760 19015 765
rect 18980 740 19015 760
rect 18980 735 18985 740
rect 18945 730 18985 735
rect 19010 735 19015 740
rect 19045 760 19050 765
rect 19120 765 19160 770
rect 19120 760 19125 765
rect 19045 740 19125 760
rect 19045 735 19050 740
rect 19010 730 19050 735
rect 19120 735 19125 740
rect 19155 735 19160 765
rect 19120 730 19160 735
rect 16545 715 16585 720
rect 16545 685 16550 715
rect 16580 710 16585 715
rect 16780 715 16820 720
rect 16780 710 16785 715
rect 16580 690 16785 710
rect 16580 685 16585 690
rect 16545 680 16585 685
rect 16780 685 16785 690
rect 16815 685 16820 715
rect 16780 680 16820 685
rect 16480 545 16520 550
rect 16480 515 16485 545
rect 16515 540 16520 545
rect 16610 545 16650 550
rect 16610 540 16615 545
rect 16515 520 16615 540
rect 16515 515 16520 520
rect 16480 510 16520 515
rect 16610 515 16615 520
rect 16645 540 16650 545
rect 16840 545 16880 550
rect 16840 540 16845 545
rect 16645 520 16845 540
rect 16645 515 16650 520
rect 16610 510 16650 515
rect 16840 515 16845 520
rect 16875 515 16880 545
rect 16840 510 16880 515
rect 19080 495 19120 500
rect 19080 465 19085 495
rect 19115 490 19120 495
rect 19260 495 19300 500
rect 19260 490 19265 495
rect 19115 470 19265 490
rect 19115 465 19120 470
rect 19080 460 19120 465
rect 19260 465 19265 470
rect 19295 465 19300 495
rect 19260 460 19300 465
rect 16305 445 16345 450
rect 16305 415 16310 445
rect 16340 440 16345 445
rect 17600 445 17640 450
rect 17600 440 17605 445
rect 16340 420 17605 440
rect 16340 415 16345 420
rect 16305 410 16345 415
rect 17600 415 17605 420
rect 17635 440 17640 445
rect 17960 445 18000 450
rect 17960 440 17965 445
rect 17635 420 17965 440
rect 17635 415 17640 420
rect 17600 410 17640 415
rect 17960 415 17965 420
rect 17995 440 18000 445
rect 19460 445 19500 450
rect 19460 440 19465 445
rect 17995 420 19465 440
rect 17995 415 18000 420
rect 17960 410 18000 415
rect 19460 415 19465 420
rect 19495 415 19500 445
rect 19460 410 19500 415
rect 16260 390 16300 395
rect 16260 360 16265 390
rect 16295 385 16300 390
rect 16780 390 16820 395
rect 16780 385 16785 390
rect 16295 365 16785 385
rect 16295 360 16300 365
rect 16260 355 16300 360
rect 16780 360 16785 365
rect 16815 385 16820 390
rect 17420 390 17460 395
rect 17420 385 17425 390
rect 16815 365 17425 385
rect 16815 360 16820 365
rect 16780 355 16820 360
rect 17420 360 17425 365
rect 17455 385 17460 390
rect 18140 390 18180 395
rect 18140 385 18145 390
rect 17455 365 18145 385
rect 17455 360 17460 365
rect 17420 355 17460 360
rect 18140 360 18145 365
rect 18175 360 18180 390
rect 18140 355 18180 360
rect 16205 345 16245 350
rect 16205 315 16210 345
rect 16240 340 16245 345
rect 16545 345 16585 350
rect 16545 340 16550 345
rect 16240 320 16550 340
rect 16240 315 16245 320
rect 16205 310 16245 315
rect 16545 315 16550 320
rect 16580 340 16585 345
rect 17240 345 17280 350
rect 17240 340 17245 345
rect 16580 320 17245 340
rect 16580 315 16585 320
rect 16545 310 16585 315
rect 17240 315 17245 320
rect 17275 340 17280 345
rect 18320 345 18360 350
rect 18320 340 18325 345
rect 17275 320 18325 340
rect 17275 315 17280 320
rect 17240 310 17280 315
rect 18320 315 18325 320
rect 18355 315 18360 345
rect 18320 310 18360 315
rect 17060 300 17100 305
rect 17060 270 17065 300
rect 17095 295 17100 300
rect 17780 300 17820 305
rect 17780 295 17785 300
rect 17095 275 17785 295
rect 17095 270 17100 275
rect 17060 265 17100 270
rect 17780 270 17785 275
rect 17815 295 17820 300
rect 18500 300 18540 305
rect 18500 295 18505 300
rect 17815 275 18505 295
rect 17815 270 17820 275
rect 17780 265 17820 270
rect 18500 270 18505 275
rect 18535 295 18540 300
rect 19405 300 19445 305
rect 19405 295 19410 300
rect 18535 275 19410 295
rect 18535 270 18540 275
rect 18500 265 18540 270
rect 19405 270 19410 275
rect 19440 270 19445 300
rect 19405 265 19445 270
rect 18000 250 18040 255
rect 18000 220 18005 250
rect 18035 245 18040 250
rect 18720 250 18760 255
rect 18720 245 18725 250
rect 18035 225 18725 245
rect 18035 220 18040 225
rect 18000 215 18040 220
rect 18720 220 18725 225
rect 18755 245 18760 250
rect 19025 250 19065 255
rect 19025 245 19030 250
rect 18755 225 19030 245
rect 18755 220 18760 225
rect 18720 215 18760 220
rect 19025 220 19030 225
rect 19060 245 19065 250
rect 19610 250 19650 255
rect 19610 245 19615 250
rect 19060 225 19615 245
rect 19060 220 19065 225
rect 19025 215 19065 220
rect 19610 220 19615 225
rect 19645 220 19650 250
rect 19610 215 19650 220
rect 16420 185 16460 190
rect 16420 155 16425 185
rect 16455 180 16460 185
rect 16540 185 16580 190
rect 16540 180 16545 185
rect 16455 160 16545 180
rect 16455 155 16460 160
rect 16420 150 16460 155
rect 16540 155 16545 160
rect 16575 180 16580 185
rect 16660 185 16700 190
rect 16660 180 16665 185
rect 16575 160 16665 180
rect 16575 155 16580 160
rect 16540 150 16580 155
rect 16660 155 16665 160
rect 16695 180 16700 185
rect 16780 185 16820 190
rect 16780 180 16785 185
rect 16695 160 16785 180
rect 16695 155 16700 160
rect 16660 150 16700 155
rect 16780 155 16785 160
rect 16815 180 16820 185
rect 16900 185 16940 190
rect 16900 180 16905 185
rect 16815 160 16905 180
rect 16815 155 16820 160
rect 16780 150 16820 155
rect 16900 155 16905 160
rect 16935 180 16940 185
rect 17020 185 17060 190
rect 17020 180 17025 185
rect 16935 160 17025 180
rect 16935 155 16940 160
rect 16900 150 16940 155
rect 17020 155 17025 160
rect 17055 180 17060 185
rect 17140 185 17180 190
rect 17140 180 17145 185
rect 17055 160 17145 180
rect 17055 155 17060 160
rect 17020 150 17060 155
rect 17140 155 17145 160
rect 17175 180 17180 185
rect 17260 185 17300 190
rect 17260 180 17265 185
rect 17175 160 17265 180
rect 17175 155 17180 160
rect 17140 150 17180 155
rect 17260 155 17265 160
rect 17295 180 17300 185
rect 17380 185 17420 190
rect 17380 180 17385 185
rect 17295 160 17385 180
rect 17295 155 17300 160
rect 17260 150 17300 155
rect 17380 155 17385 160
rect 17415 180 17420 185
rect 17500 185 17540 190
rect 17500 180 17505 185
rect 17415 160 17505 180
rect 17415 155 17420 160
rect 17380 150 17420 155
rect 17500 155 17505 160
rect 17535 180 17540 185
rect 17620 185 17660 190
rect 17620 180 17625 185
rect 17535 160 17625 180
rect 17535 155 17540 160
rect 17500 150 17540 155
rect 17620 155 17625 160
rect 17655 180 17660 185
rect 17940 185 17980 190
rect 17940 180 17945 185
rect 17655 160 17945 180
rect 17655 155 17660 160
rect 17620 150 17660 155
rect 17940 155 17945 160
rect 17975 180 17980 185
rect 18060 185 18100 190
rect 18060 180 18065 185
rect 17975 160 18065 180
rect 17975 155 17980 160
rect 17940 150 17980 155
rect 18060 155 18065 160
rect 18095 180 18100 185
rect 18180 185 18220 190
rect 18180 180 18185 185
rect 18095 160 18185 180
rect 18095 155 18100 160
rect 18060 150 18100 155
rect 18180 155 18185 160
rect 18215 180 18220 185
rect 18300 185 18340 190
rect 18300 180 18305 185
rect 18215 160 18305 180
rect 18215 155 18220 160
rect 18180 150 18220 155
rect 18300 155 18305 160
rect 18335 180 18340 185
rect 18420 185 18460 190
rect 18420 180 18425 185
rect 18335 160 18425 180
rect 18335 155 18340 160
rect 18300 150 18340 155
rect 18420 155 18425 160
rect 18455 180 18460 185
rect 18540 185 18580 190
rect 18540 180 18545 185
rect 18455 160 18545 180
rect 18455 155 18460 160
rect 18420 150 18460 155
rect 18540 155 18545 160
rect 18575 180 18580 185
rect 18660 185 18700 190
rect 18660 180 18665 185
rect 18575 160 18665 180
rect 18575 155 18580 160
rect 18540 150 18580 155
rect 18660 155 18665 160
rect 18695 180 18700 185
rect 18780 185 18820 190
rect 18780 180 18785 185
rect 18695 160 18785 180
rect 18695 155 18700 160
rect 18660 150 18700 155
rect 18780 155 18785 160
rect 18815 180 18820 185
rect 18900 185 18940 190
rect 18900 180 18905 185
rect 18815 160 18905 180
rect 18815 155 18820 160
rect 18780 150 18820 155
rect 18900 155 18905 160
rect 18935 180 18940 185
rect 19020 185 19060 190
rect 19020 180 19025 185
rect 18935 160 19025 180
rect 18935 155 18940 160
rect 18900 150 18940 155
rect 19020 155 19025 160
rect 19055 180 19060 185
rect 19140 185 19180 190
rect 19140 180 19145 185
rect 19055 160 19145 180
rect 19055 155 19060 160
rect 19020 150 19060 155
rect 19140 155 19145 160
rect 19175 180 19180 185
rect 20050 185 20090 190
rect 20050 180 20055 185
rect 19175 160 20055 180
rect 19175 155 19180 160
rect 19140 150 19180 155
rect 20050 155 20055 160
rect 20085 155 20090 185
rect 20050 150 20090 155
rect 15950 125 15990 130
rect 15950 95 15955 125
rect 15985 120 15990 125
rect 16480 125 16520 130
rect 16480 120 16485 125
rect 15985 100 16485 120
rect 15985 95 15990 100
rect 15950 90 15990 95
rect 16480 95 16485 100
rect 16515 120 16520 125
rect 16840 125 16880 130
rect 16840 120 16845 125
rect 16515 100 16845 120
rect 16515 95 16520 100
rect 16480 90 16520 95
rect 16840 95 16845 100
rect 16875 120 16880 125
rect 17200 125 17240 130
rect 17200 120 17205 125
rect 16875 100 17205 120
rect 16875 95 16880 100
rect 16840 90 16880 95
rect 17200 95 17205 100
rect 17235 120 17240 125
rect 17560 125 17600 130
rect 17560 120 17565 125
rect 17235 100 17565 120
rect 17235 95 17240 100
rect 17200 90 17240 95
rect 17560 95 17565 100
rect 17595 120 17600 125
rect 17690 125 17730 130
rect 17690 120 17695 125
rect 17595 100 17695 120
rect 17595 95 17600 100
rect 17560 90 17600 95
rect 17690 95 17695 100
rect 17725 95 17730 125
rect 17690 90 17730 95
rect 17870 125 17910 130
rect 17870 95 17875 125
rect 17905 120 17910 125
rect 18000 125 18040 130
rect 18000 120 18005 125
rect 17905 100 18005 120
rect 17905 95 17910 100
rect 17870 90 17910 95
rect 18000 95 18005 100
rect 18035 120 18040 125
rect 18360 125 18400 130
rect 18360 120 18365 125
rect 18035 100 18365 120
rect 18035 95 18040 100
rect 18000 90 18040 95
rect 18360 95 18365 100
rect 18395 120 18400 125
rect 18720 125 18760 130
rect 18720 120 18725 125
rect 18395 100 18725 120
rect 18395 95 18400 100
rect 18360 90 18400 95
rect 18720 95 18725 100
rect 18755 120 18760 125
rect 19080 125 19120 130
rect 19080 120 19085 125
rect 18755 100 19085 120
rect 18755 95 18760 100
rect 18720 90 18760 95
rect 19080 95 19085 100
rect 19115 95 19120 125
rect 19080 90 19120 95
rect 16600 -45 16640 -40
rect 16600 -75 16605 -45
rect 16635 -50 16640 -45
rect 16720 -50 16760 -40
rect 16960 -45 17000 -40
rect 16960 -50 16965 -45
rect 16635 -70 16965 -50
rect 16635 -75 16640 -70
rect 16600 -80 16640 -75
rect 16720 -80 16760 -70
rect 16960 -75 16965 -70
rect 16995 -50 17000 -45
rect 17080 -50 17120 -40
rect 17320 -45 17360 -40
rect 17320 -50 17325 -45
rect 16995 -70 17325 -50
rect 16995 -75 17000 -70
rect 16960 -80 17000 -75
rect 17080 -80 17120 -70
rect 17320 -75 17325 -70
rect 17355 -75 17360 -45
rect 17320 -80 17360 -75
rect 17440 -80 17480 -40
rect 18120 -80 18160 -40
rect 18240 -45 18280 -40
rect 18240 -75 18245 -45
rect 18275 -50 18280 -45
rect 18480 -50 18520 -40
rect 18600 -45 18640 -40
rect 18600 -50 18605 -45
rect 18275 -70 18605 -50
rect 18275 -75 18280 -70
rect 18240 -80 18280 -75
rect 18480 -80 18520 -70
rect 18600 -75 18605 -70
rect 18635 -50 18640 -45
rect 18840 -50 18880 -40
rect 18960 -45 19000 -40
rect 18960 -50 18965 -45
rect 18635 -70 18965 -50
rect 18635 -75 18640 -70
rect 18600 -80 18640 -75
rect 18840 -80 18880 -70
rect 18960 -75 18965 -70
rect 18995 -75 19000 -45
rect 18960 -80 19000 -75
rect 15725 -105 15765 -100
rect 15725 -135 15730 -105
rect 15760 -110 15765 -105
rect 16510 -105 16550 -100
rect 16510 -110 16515 -105
rect 15760 -130 16515 -110
rect 15760 -135 15765 -130
rect 15725 -140 15765 -135
rect 16510 -135 16515 -130
rect 16545 -110 16550 -105
rect 16720 -105 16760 -100
rect 16720 -110 16725 -105
rect 16545 -130 16725 -110
rect 16545 -135 16550 -130
rect 16510 -140 16550 -135
rect 16720 -135 16725 -130
rect 16755 -110 16760 -105
rect 16840 -105 16880 -100
rect 16840 -110 16845 -105
rect 16755 -130 16845 -110
rect 16755 -135 16760 -130
rect 16720 -140 16760 -135
rect 16840 -135 16845 -130
rect 16875 -110 16880 -105
rect 17080 -105 17120 -100
rect 17080 -110 17085 -105
rect 16875 -130 17085 -110
rect 16875 -135 16880 -130
rect 16840 -140 16880 -135
rect 17080 -135 17085 -130
rect 17115 -110 17120 -105
rect 17200 -105 17240 -100
rect 17200 -110 17205 -105
rect 17115 -130 17205 -110
rect 17115 -135 17120 -130
rect 17080 -140 17120 -135
rect 17200 -135 17205 -130
rect 17235 -110 17240 -105
rect 17440 -105 17480 -100
rect 17440 -110 17445 -105
rect 17235 -130 17445 -110
rect 17235 -135 17240 -130
rect 17200 -140 17240 -135
rect 17440 -135 17445 -130
rect 17475 -110 17480 -105
rect 17530 -105 17570 -100
rect 17530 -110 17535 -105
rect 17475 -130 17535 -110
rect 17475 -135 17480 -130
rect 17440 -140 17480 -135
rect 17530 -135 17535 -130
rect 17565 -135 17570 -105
rect 17530 -140 17570 -135
rect 18030 -105 18070 -100
rect 18030 -135 18035 -105
rect 18065 -110 18070 -105
rect 18120 -105 18160 -100
rect 18120 -110 18125 -105
rect 18065 -130 18125 -110
rect 18065 -135 18070 -130
rect 18030 -140 18070 -135
rect 18120 -135 18125 -130
rect 18155 -110 18160 -105
rect 18360 -105 18400 -100
rect 18360 -110 18365 -105
rect 18155 -130 18365 -110
rect 18155 -135 18160 -130
rect 18120 -140 18160 -135
rect 18360 -135 18365 -130
rect 18395 -110 18400 -105
rect 18480 -105 18520 -100
rect 18480 -110 18485 -105
rect 18395 -130 18485 -110
rect 18395 -135 18400 -130
rect 18360 -140 18400 -135
rect 18480 -135 18485 -130
rect 18515 -110 18520 -105
rect 18720 -105 18760 -100
rect 18720 -110 18725 -105
rect 18515 -130 18725 -110
rect 18515 -135 18520 -130
rect 18480 -140 18520 -135
rect 18720 -135 18725 -130
rect 18755 -110 18760 -105
rect 18840 -105 18880 -100
rect 18840 -110 18845 -105
rect 18755 -130 18845 -110
rect 18755 -135 18760 -130
rect 18720 -140 18760 -135
rect 18840 -135 18845 -130
rect 18875 -110 18880 -105
rect 19050 -105 19090 -100
rect 19050 -110 19055 -105
rect 18875 -130 19055 -110
rect 18875 -135 18880 -130
rect 18840 -140 18880 -135
rect 19050 -135 19055 -130
rect 19085 -110 19090 -105
rect 19730 -105 19770 -100
rect 19730 -110 19735 -105
rect 19085 -130 19735 -110
rect 19085 -135 19090 -130
rect 19050 -140 19090 -135
rect 19730 -135 19735 -130
rect 19765 -135 19770 -105
rect 19730 -140 19770 -135
rect 16970 -190 17010 -185
rect 16260 -205 16300 -200
rect 16260 -235 16265 -205
rect 16295 -210 16300 -205
rect 16910 -205 16950 -200
rect 16910 -210 16915 -205
rect 16295 -230 16915 -210
rect 16295 -235 16300 -230
rect 16260 -240 16300 -235
rect 16910 -235 16915 -230
rect 16945 -235 16950 -205
rect 16970 -220 16975 -190
rect 17005 -195 17010 -190
rect 17210 -190 17250 -185
rect 17210 -195 17215 -190
rect 17005 -215 17215 -195
rect 17005 -220 17010 -215
rect 16970 -225 17010 -220
rect 17210 -220 17215 -215
rect 17245 -195 17250 -190
rect 17450 -190 17490 -185
rect 17450 -195 17455 -190
rect 17245 -215 17455 -195
rect 17245 -220 17250 -215
rect 17210 -225 17250 -220
rect 17450 -220 17455 -215
rect 17485 -220 17490 -190
rect 17450 -225 17490 -220
rect 18110 -190 18150 -185
rect 18110 -220 18115 -190
rect 18145 -195 18150 -190
rect 18350 -190 18390 -185
rect 18350 -195 18355 -190
rect 18145 -215 18355 -195
rect 18145 -220 18150 -215
rect 18110 -225 18150 -220
rect 18350 -220 18355 -215
rect 18385 -195 18390 -190
rect 18590 -190 18630 -185
rect 18590 -195 18595 -190
rect 18385 -215 18595 -195
rect 18385 -220 18390 -215
rect 18350 -225 18390 -220
rect 18590 -220 18595 -215
rect 18625 -220 18630 -190
rect 18590 -225 18630 -220
rect 18650 -205 18690 -200
rect 16910 -240 16950 -235
rect 18650 -235 18655 -205
rect 18685 -210 18690 -205
rect 19405 -205 19445 -200
rect 19405 -210 19410 -205
rect 18685 -230 19410 -210
rect 18685 -235 18690 -230
rect 18650 -240 18690 -235
rect 19405 -235 19410 -230
rect 19440 -235 19445 -205
rect 19405 -240 19445 -235
rect 16850 -250 16890 -245
rect 16850 -280 16855 -250
rect 16885 -255 16890 -250
rect 17090 -250 17130 -245
rect 17090 -255 17095 -250
rect 16885 -275 17095 -255
rect 16885 -280 16890 -275
rect 16850 -285 16890 -280
rect 17090 -280 17095 -275
rect 17125 -255 17130 -250
rect 17330 -250 17370 -245
rect 17330 -255 17335 -250
rect 17125 -275 17335 -255
rect 17125 -280 17130 -275
rect 17090 -285 17130 -280
rect 17330 -280 17335 -275
rect 17365 -280 17370 -250
rect 17330 -285 17370 -280
rect 18230 -250 18270 -245
rect 18230 -280 18235 -250
rect 18265 -255 18270 -250
rect 18470 -250 18510 -245
rect 18470 -255 18475 -250
rect 18265 -275 18475 -255
rect 18265 -280 18270 -275
rect 18230 -285 18270 -280
rect 18470 -280 18475 -275
rect 18505 -255 18510 -250
rect 18710 -250 18750 -245
rect 18710 -255 18715 -250
rect 18505 -275 18715 -255
rect 18505 -280 18510 -275
rect 18470 -285 18510 -280
rect 18710 -280 18715 -275
rect 18745 -280 18750 -250
rect 18710 -285 18750 -280
rect 17565 -310 17595 -305
rect 17780 -310 17820 -305
rect 17780 -315 17785 -310
rect 17595 -335 17785 -315
rect 17565 -345 17595 -340
rect 17780 -340 17785 -335
rect 17815 -315 17820 -310
rect 18005 -310 18035 -305
rect 17815 -335 18005 -315
rect 17815 -340 17820 -335
rect 17780 -345 17820 -340
rect 18005 -345 18035 -340
rect 16305 -370 16345 -365
rect 16305 -400 16310 -370
rect 16340 -375 16345 -370
rect 16850 -370 16890 -365
rect 16850 -375 16855 -370
rect 16340 -395 16855 -375
rect 16340 -400 16345 -395
rect 16305 -405 16345 -400
rect 16850 -400 16855 -395
rect 16885 -400 16890 -370
rect 16850 -405 16890 -400
rect 18710 -370 18750 -365
rect 18710 -400 18715 -370
rect 18745 -375 18750 -370
rect 19325 -370 19365 -365
rect 19325 -375 19330 -370
rect 18745 -395 19330 -375
rect 18745 -400 18750 -395
rect 18710 -405 18750 -400
rect 19325 -400 19330 -395
rect 19360 -400 19365 -370
rect 19325 -405 19365 -400
rect 16530 -430 16570 -425
rect 16530 -460 16535 -430
rect 16565 -435 16570 -430
rect 16910 -430 16950 -425
rect 16910 -435 16915 -430
rect 16565 -455 16915 -435
rect 16565 -460 16570 -455
rect 16530 -465 16570 -460
rect 16910 -460 16915 -455
rect 16945 -435 16950 -430
rect 17030 -430 17070 -425
rect 17030 -435 17035 -430
rect 16945 -455 17035 -435
rect 16945 -460 16950 -455
rect 16910 -465 16950 -460
rect 17030 -460 17035 -455
rect 17065 -435 17070 -430
rect 17150 -430 17190 -425
rect 17150 -435 17155 -430
rect 17065 -455 17155 -435
rect 17065 -460 17070 -455
rect 17030 -465 17070 -460
rect 17150 -460 17155 -455
rect 17185 -435 17190 -430
rect 17270 -430 17310 -425
rect 17270 -435 17275 -430
rect 17185 -455 17275 -435
rect 17185 -460 17190 -455
rect 17150 -465 17190 -460
rect 17270 -460 17275 -455
rect 17305 -435 17310 -430
rect 17390 -430 17430 -425
rect 17390 -435 17395 -430
rect 17305 -455 17395 -435
rect 17305 -460 17310 -455
rect 17270 -465 17310 -460
rect 17390 -460 17395 -455
rect 17425 -460 17430 -430
rect 17390 -465 17430 -460
rect 18170 -430 18210 -425
rect 18170 -460 18175 -430
rect 18205 -435 18210 -430
rect 18290 -430 18330 -425
rect 18290 -435 18295 -430
rect 18205 -455 18295 -435
rect 18205 -460 18210 -455
rect 18170 -465 18210 -460
rect 18290 -460 18295 -455
rect 18325 -435 18330 -430
rect 18410 -430 18450 -425
rect 18410 -435 18415 -430
rect 18325 -455 18415 -435
rect 18325 -460 18330 -455
rect 18290 -465 18330 -460
rect 18410 -460 18415 -455
rect 18445 -435 18450 -430
rect 18530 -430 18570 -425
rect 18530 -435 18535 -430
rect 18445 -455 18535 -435
rect 18445 -460 18450 -455
rect 18410 -465 18450 -460
rect 18530 -460 18535 -455
rect 18565 -435 18570 -430
rect 18650 -430 18690 -425
rect 18650 -435 18655 -430
rect 18565 -455 18655 -435
rect 18565 -460 18570 -455
rect 18530 -465 18570 -460
rect 18650 -460 18655 -455
rect 18685 -435 18690 -430
rect 19030 -430 19070 -425
rect 19030 -435 19035 -430
rect 18685 -455 19035 -435
rect 18685 -460 18690 -455
rect 18650 -465 18690 -460
rect 19030 -460 19035 -455
rect 19065 -460 19070 -430
rect 19030 -465 19070 -460
rect 16620 -530 16660 -525
rect 16620 -560 16625 -530
rect 16655 -535 16660 -530
rect 16740 -530 16780 -525
rect 16740 -535 16745 -530
rect 16655 -555 16745 -535
rect 16655 -560 16660 -555
rect 16620 -565 16660 -560
rect 16740 -560 16745 -555
rect 16775 -535 16780 -530
rect 16860 -530 16900 -525
rect 16860 -535 16865 -530
rect 16775 -555 16865 -535
rect 16775 -560 16780 -555
rect 16740 -565 16780 -560
rect 16860 -560 16865 -555
rect 16895 -535 16900 -530
rect 16980 -530 17020 -525
rect 16980 -535 16985 -530
rect 16895 -555 16985 -535
rect 16895 -560 16900 -555
rect 16860 -565 16900 -560
rect 16980 -560 16985 -555
rect 17015 -535 17020 -530
rect 17300 -530 17340 -525
rect 17300 -535 17305 -530
rect 17015 -555 17305 -535
rect 17015 -560 17020 -555
rect 16980 -565 17020 -560
rect 17300 -560 17305 -555
rect 17335 -535 17340 -530
rect 17420 -530 17460 -525
rect 17420 -535 17425 -530
rect 17335 -555 17425 -535
rect 17335 -560 17340 -555
rect 17300 -565 17340 -560
rect 17420 -560 17425 -555
rect 17455 -535 17460 -530
rect 17540 -530 17580 -525
rect 17540 -535 17545 -530
rect 17455 -555 17545 -535
rect 17455 -560 17460 -555
rect 17420 -565 17460 -560
rect 17540 -560 17545 -555
rect 17575 -535 17580 -530
rect 18020 -530 18060 -525
rect 18020 -535 18025 -530
rect 17575 -555 18025 -535
rect 17575 -560 17580 -555
rect 17540 -565 17580 -560
rect 18020 -560 18025 -555
rect 18055 -535 18060 -530
rect 18140 -530 18180 -525
rect 18140 -535 18145 -530
rect 18055 -555 18145 -535
rect 18055 -560 18060 -555
rect 18020 -565 18060 -560
rect 18140 -560 18145 -555
rect 18175 -535 18180 -530
rect 18260 -530 18300 -525
rect 18260 -535 18265 -530
rect 18175 -555 18265 -535
rect 18175 -560 18180 -555
rect 18140 -565 18180 -560
rect 18260 -560 18265 -555
rect 18295 -535 18300 -530
rect 18580 -530 18620 -525
rect 18580 -535 18585 -530
rect 18295 -555 18585 -535
rect 18295 -560 18300 -555
rect 18260 -565 18300 -560
rect 18580 -560 18585 -555
rect 18615 -535 18620 -530
rect 18700 -530 18740 -525
rect 18700 -535 18705 -530
rect 18615 -555 18705 -535
rect 18615 -560 18620 -555
rect 18580 -565 18620 -560
rect 18700 -560 18705 -555
rect 18735 -535 18740 -530
rect 18820 -530 18860 -525
rect 18820 -535 18825 -530
rect 18735 -555 18825 -535
rect 18735 -560 18740 -555
rect 18700 -565 18740 -560
rect 18820 -560 18825 -555
rect 18855 -535 18860 -530
rect 18940 -530 18980 -525
rect 18940 -535 18945 -530
rect 18855 -555 18945 -535
rect 18855 -560 18860 -555
rect 18820 -565 18860 -560
rect 18940 -560 18945 -555
rect 18975 -535 18980 -530
rect 20050 -530 20090 -525
rect 20050 -535 20055 -530
rect 18975 -555 20055 -535
rect 18975 -560 18980 -555
rect 18940 -565 18980 -560
rect 20050 -560 20055 -555
rect 20085 -560 20090 -530
rect 20050 -565 20090 -560
rect 17110 -845 17150 -840
rect 17110 -875 17115 -845
rect 17145 -850 17150 -845
rect 17780 -845 17820 -840
rect 17780 -850 17785 -845
rect 17145 -870 17785 -850
rect 17145 -875 17150 -870
rect 17110 -880 17150 -875
rect 17780 -875 17785 -870
rect 17815 -850 17820 -845
rect 18450 -845 18490 -840
rect 18450 -850 18455 -845
rect 17815 -870 18455 -850
rect 17815 -875 17820 -870
rect 17780 -880 17820 -875
rect 18450 -875 18455 -870
rect 18485 -850 18490 -845
rect 19965 -845 20005 -840
rect 19965 -850 19970 -845
rect 18485 -870 19970 -850
rect 18485 -875 18490 -870
rect 18450 -880 18490 -875
rect 19965 -875 19970 -870
rect 20000 -875 20005 -845
rect 19965 -880 20005 -875
rect 16740 -995 16780 -990
rect 16740 -1025 16745 -995
rect 16775 -1000 16780 -995
rect 16820 -995 16860 -990
rect 16820 -1000 16825 -995
rect 16775 -1020 16825 -1000
rect 16775 -1025 16780 -1020
rect 16740 -1030 16780 -1025
rect 16820 -1025 16825 -1020
rect 16855 -1000 16860 -995
rect 16900 -995 16940 -990
rect 16900 -1000 16905 -995
rect 16855 -1020 16905 -1000
rect 16855 -1025 16860 -1020
rect 16820 -1030 16860 -1025
rect 16900 -1025 16905 -1020
rect 16935 -1000 16940 -995
rect 16980 -995 17020 -990
rect 16980 -1000 16985 -995
rect 16935 -1020 16985 -1000
rect 16935 -1025 16940 -1020
rect 16900 -1030 16940 -1025
rect 16980 -1025 16985 -1020
rect 17015 -1000 17020 -995
rect 17060 -995 17100 -990
rect 17060 -1000 17065 -995
rect 17015 -1020 17065 -1000
rect 17015 -1025 17020 -1020
rect 16980 -1030 17020 -1025
rect 17060 -1025 17065 -1020
rect 17095 -1000 17100 -995
rect 17140 -995 17180 -990
rect 17140 -1000 17145 -995
rect 17095 -1020 17145 -1000
rect 17095 -1025 17100 -1020
rect 17060 -1030 17100 -1025
rect 17140 -1025 17145 -1020
rect 17175 -1000 17180 -995
rect 17220 -995 17260 -990
rect 17220 -1000 17225 -995
rect 17175 -1020 17225 -1000
rect 17175 -1025 17180 -1020
rect 17140 -1030 17180 -1025
rect 17220 -1025 17225 -1020
rect 17255 -1000 17260 -995
rect 17300 -995 17340 -990
rect 17300 -1000 17305 -995
rect 17255 -1020 17305 -1000
rect 17255 -1025 17260 -1020
rect 17220 -1030 17260 -1025
rect 17300 -1025 17305 -1020
rect 17335 -1000 17340 -995
rect 17380 -995 17420 -990
rect 17380 -1000 17385 -995
rect 17335 -1020 17385 -1000
rect 17335 -1025 17340 -1020
rect 17300 -1030 17340 -1025
rect 17380 -1025 17385 -1020
rect 17415 -1000 17420 -995
rect 17460 -995 17500 -990
rect 17460 -1000 17465 -995
rect 17415 -1020 17465 -1000
rect 17415 -1025 17420 -1020
rect 17380 -1030 17420 -1025
rect 17460 -1025 17465 -1020
rect 17495 -1000 17500 -995
rect 17540 -995 17580 -990
rect 17540 -1000 17545 -995
rect 17495 -1020 17545 -1000
rect 17495 -1025 17500 -1020
rect 17460 -1030 17500 -1025
rect 17540 -1025 17545 -1020
rect 17575 -1000 17580 -995
rect 17620 -995 17660 -990
rect 17620 -1000 17625 -995
rect 17575 -1020 17625 -1000
rect 17575 -1025 17580 -1020
rect 17540 -1030 17580 -1025
rect 17620 -1025 17625 -1020
rect 17655 -1000 17660 -995
rect 17700 -995 17740 -990
rect 17700 -1000 17705 -995
rect 17655 -1020 17705 -1000
rect 17655 -1025 17660 -1020
rect 17620 -1030 17660 -1025
rect 17700 -1025 17705 -1020
rect 17735 -1025 17740 -995
rect 17700 -1030 17740 -1025
rect 17780 -995 17820 -990
rect 17780 -1025 17785 -995
rect 17815 -1000 17820 -995
rect 17860 -995 17900 -990
rect 17860 -1000 17865 -995
rect 17815 -1020 17865 -1000
rect 17815 -1025 17820 -1020
rect 17780 -1030 17820 -1025
rect 17860 -1025 17865 -1020
rect 17895 -1000 17900 -995
rect 17940 -995 17980 -990
rect 17940 -1000 17945 -995
rect 17895 -1020 17945 -1000
rect 17895 -1025 17900 -1020
rect 17860 -1030 17900 -1025
rect 17940 -1025 17945 -1020
rect 17975 -1000 17980 -995
rect 18020 -995 18060 -990
rect 18020 -1000 18025 -995
rect 17975 -1020 18025 -1000
rect 17975 -1025 17980 -1020
rect 17940 -1030 17980 -1025
rect 18020 -1025 18025 -1020
rect 18055 -1000 18060 -995
rect 18100 -995 18140 -990
rect 18100 -1000 18105 -995
rect 18055 -1020 18105 -1000
rect 18055 -1025 18060 -1020
rect 18020 -1030 18060 -1025
rect 18100 -1025 18105 -1020
rect 18135 -1000 18140 -995
rect 18180 -995 18220 -990
rect 18180 -1000 18185 -995
rect 18135 -1020 18185 -1000
rect 18135 -1025 18140 -1020
rect 18100 -1030 18140 -1025
rect 18180 -1025 18185 -1020
rect 18215 -1000 18220 -995
rect 18260 -995 18300 -990
rect 18260 -1000 18265 -995
rect 18215 -1020 18265 -1000
rect 18215 -1025 18220 -1020
rect 18180 -1030 18220 -1025
rect 18260 -1025 18265 -1020
rect 18295 -1000 18300 -995
rect 18340 -995 18380 -990
rect 18340 -1000 18345 -995
rect 18295 -1020 18345 -1000
rect 18295 -1025 18300 -1020
rect 18260 -1030 18300 -1025
rect 18340 -1025 18345 -1020
rect 18375 -1000 18380 -995
rect 18420 -995 18460 -990
rect 18420 -1000 18425 -995
rect 18375 -1020 18425 -1000
rect 18375 -1025 18380 -1020
rect 18340 -1030 18380 -1025
rect 18420 -1025 18425 -1020
rect 18455 -1000 18460 -995
rect 18500 -995 18540 -990
rect 18500 -1000 18505 -995
rect 18455 -1020 18505 -1000
rect 18455 -1025 18460 -1020
rect 18420 -1030 18460 -1025
rect 18500 -1025 18505 -1020
rect 18535 -1000 18540 -995
rect 18580 -995 18620 -990
rect 18580 -1000 18585 -995
rect 18535 -1020 18585 -1000
rect 18535 -1025 18540 -1020
rect 18500 -1030 18540 -1025
rect 18580 -1025 18585 -1020
rect 18615 -1000 18620 -995
rect 18660 -995 18700 -990
rect 18660 -1000 18665 -995
rect 18615 -1020 18665 -1000
rect 18615 -1025 18620 -1020
rect 18580 -1030 18620 -1025
rect 18660 -1025 18665 -1020
rect 18695 -1000 18700 -995
rect 18740 -995 18780 -990
rect 18740 -1000 18745 -995
rect 18695 -1020 18745 -1000
rect 18695 -1025 18700 -1020
rect 18660 -1030 18700 -1025
rect 18740 -1025 18745 -1020
rect 18775 -1025 18780 -995
rect 18740 -1030 18780 -1025
rect 16205 -1080 16245 -1075
rect 16205 -1110 16210 -1080
rect 16240 -1085 16245 -1080
rect 16700 -1080 16740 -1075
rect 16700 -1085 16705 -1080
rect 16240 -1105 16705 -1085
rect 16240 -1110 16245 -1105
rect 16205 -1115 16245 -1110
rect 16700 -1110 16705 -1105
rect 16735 -1110 16740 -1080
rect 16700 -1115 16740 -1110
rect 18895 -1080 18935 -1075
rect 18895 -1110 18900 -1080
rect 18930 -1085 18935 -1080
rect 19965 -1080 20005 -1075
rect 19965 -1085 19970 -1080
rect 18930 -1105 19970 -1085
rect 18930 -1110 18935 -1105
rect 18895 -1115 18935 -1110
rect 19965 -1110 19970 -1105
rect 20000 -1110 20005 -1080
rect 19965 -1115 20005 -1110
rect 17165 -1200 17205 -1195
rect 17165 -1230 17170 -1200
rect 17200 -1205 17205 -1200
rect 17780 -1200 17820 -1195
rect 17780 -1205 17785 -1200
rect 17200 -1225 17785 -1205
rect 17200 -1230 17205 -1225
rect 17165 -1235 17205 -1230
rect 17780 -1230 17785 -1225
rect 17815 -1205 17820 -1200
rect 18395 -1200 18435 -1195
rect 18395 -1205 18400 -1200
rect 17815 -1225 18400 -1205
rect 17815 -1230 17820 -1225
rect 17780 -1235 17820 -1230
rect 18395 -1230 18400 -1225
rect 18430 -1230 18435 -1200
rect 18395 -1235 18435 -1230
rect 16890 -1270 16930 -1265
rect 16890 -1300 16895 -1270
rect 16925 -1275 16930 -1270
rect 17000 -1270 17040 -1265
rect 17000 -1275 17005 -1270
rect 16925 -1295 17005 -1275
rect 16925 -1300 16930 -1295
rect 16890 -1305 16930 -1300
rect 17000 -1300 17005 -1295
rect 17035 -1275 17040 -1270
rect 17110 -1270 17150 -1265
rect 17110 -1275 17115 -1270
rect 17035 -1295 17115 -1275
rect 17035 -1300 17040 -1295
rect 17000 -1305 17040 -1300
rect 17110 -1300 17115 -1295
rect 17145 -1275 17150 -1270
rect 17220 -1270 17260 -1265
rect 17220 -1275 17225 -1270
rect 17145 -1295 17225 -1275
rect 17145 -1300 17150 -1295
rect 17110 -1305 17150 -1300
rect 17220 -1300 17225 -1295
rect 17255 -1275 17260 -1270
rect 17330 -1270 17370 -1265
rect 17330 -1275 17335 -1270
rect 17255 -1295 17335 -1275
rect 17255 -1300 17260 -1295
rect 17220 -1305 17260 -1300
rect 17330 -1300 17335 -1295
rect 17365 -1275 17370 -1270
rect 17505 -1270 17545 -1265
rect 17505 -1275 17510 -1270
rect 17365 -1295 17510 -1275
rect 17365 -1300 17370 -1295
rect 17330 -1305 17370 -1300
rect 17505 -1300 17510 -1295
rect 17540 -1275 17545 -1270
rect 17615 -1270 17655 -1265
rect 17615 -1275 17620 -1270
rect 17540 -1295 17620 -1275
rect 17540 -1300 17545 -1295
rect 17505 -1305 17545 -1300
rect 17615 -1300 17620 -1295
rect 17650 -1275 17655 -1270
rect 17725 -1270 17765 -1265
rect 17725 -1275 17730 -1270
rect 17650 -1295 17730 -1275
rect 17650 -1300 17655 -1295
rect 17615 -1305 17655 -1300
rect 17725 -1300 17730 -1295
rect 17760 -1275 17765 -1270
rect 17835 -1270 17875 -1265
rect 17835 -1275 17840 -1270
rect 17760 -1295 17840 -1275
rect 17760 -1300 17765 -1295
rect 17725 -1305 17765 -1300
rect 17835 -1300 17840 -1295
rect 17870 -1275 17875 -1270
rect 17945 -1270 17985 -1265
rect 17945 -1275 17950 -1270
rect 17870 -1295 17950 -1275
rect 17870 -1300 17875 -1295
rect 17835 -1305 17875 -1300
rect 17945 -1300 17950 -1295
rect 17980 -1275 17985 -1270
rect 18055 -1270 18095 -1265
rect 18055 -1275 18060 -1270
rect 17980 -1295 18060 -1275
rect 17980 -1300 17985 -1295
rect 17945 -1305 17985 -1300
rect 18055 -1300 18060 -1295
rect 18090 -1275 18095 -1270
rect 18230 -1270 18270 -1265
rect 18230 -1275 18235 -1270
rect 18090 -1295 18235 -1275
rect 18090 -1300 18095 -1295
rect 18055 -1305 18095 -1300
rect 18230 -1300 18235 -1295
rect 18265 -1275 18270 -1270
rect 18340 -1270 18380 -1265
rect 18340 -1275 18345 -1270
rect 18265 -1295 18345 -1275
rect 18265 -1300 18270 -1295
rect 18230 -1305 18270 -1300
rect 18340 -1300 18345 -1295
rect 18375 -1275 18380 -1270
rect 18450 -1270 18490 -1265
rect 18450 -1275 18455 -1270
rect 18375 -1295 18455 -1275
rect 18375 -1300 18380 -1295
rect 18340 -1305 18380 -1300
rect 18450 -1300 18455 -1295
rect 18485 -1275 18490 -1270
rect 18560 -1270 18600 -1265
rect 18560 -1275 18565 -1270
rect 18485 -1295 18565 -1275
rect 18485 -1300 18490 -1295
rect 18450 -1305 18490 -1300
rect 18560 -1300 18565 -1295
rect 18595 -1275 18600 -1270
rect 18670 -1270 18710 -1265
rect 18670 -1275 18675 -1270
rect 18595 -1295 18675 -1275
rect 18595 -1300 18600 -1295
rect 18560 -1305 18600 -1300
rect 18670 -1300 18675 -1295
rect 18705 -1275 18710 -1270
rect 19965 -1270 20005 -1265
rect 19965 -1275 19970 -1270
rect 18705 -1295 19970 -1275
rect 18705 -1300 18710 -1295
rect 18670 -1305 18710 -1300
rect 19965 -1300 19970 -1295
rect 20000 -1300 20005 -1270
rect 19965 -1305 20005 -1300
rect 17055 -1440 17095 -1435
rect 17055 -1470 17060 -1440
rect 17090 -1445 17095 -1440
rect 17275 -1440 17315 -1435
rect 17275 -1445 17280 -1440
rect 17090 -1465 17280 -1445
rect 17090 -1470 17095 -1465
rect 17055 -1475 17095 -1470
rect 17275 -1470 17280 -1465
rect 17310 -1470 17315 -1440
rect 17275 -1475 17315 -1470
rect 17780 -1440 17820 -1435
rect 17780 -1470 17785 -1440
rect 17815 -1445 17820 -1440
rect 17890 -1440 17930 -1435
rect 17890 -1445 17895 -1440
rect 17815 -1465 17895 -1445
rect 17815 -1470 17820 -1465
rect 17780 -1475 17820 -1470
rect 17890 -1470 17895 -1465
rect 17925 -1445 17930 -1440
rect 18000 -1440 18040 -1435
rect 18000 -1445 18005 -1440
rect 17925 -1465 18005 -1445
rect 17925 -1470 17930 -1465
rect 17890 -1475 17930 -1470
rect 18000 -1470 18005 -1465
rect 18035 -1470 18040 -1440
rect 18000 -1475 18040 -1470
rect 18285 -1440 18325 -1435
rect 18285 -1470 18290 -1440
rect 18320 -1445 18325 -1440
rect 18505 -1440 18545 -1435
rect 18505 -1445 18510 -1440
rect 18320 -1465 18510 -1445
rect 18320 -1470 18325 -1465
rect 18285 -1475 18325 -1470
rect 18505 -1470 18510 -1465
rect 18540 -1470 18545 -1440
rect 18505 -1475 18545 -1470
rect 17780 -1500 17820 -1495
rect 17780 -1530 17785 -1500
rect 17815 -1530 17820 -1500
rect 17780 -1535 17820 -1530
rect 16030 -1545 16070 -1540
rect 16030 -1575 16035 -1545
rect 16065 -1550 16070 -1545
rect 16945 -1545 16985 -1540
rect 16945 -1550 16950 -1545
rect 16065 -1570 16950 -1550
rect 16065 -1575 16070 -1570
rect 16030 -1580 16070 -1575
rect 16945 -1575 16950 -1570
rect 16980 -1550 16985 -1545
rect 17165 -1545 17205 -1540
rect 17165 -1550 17170 -1545
rect 16980 -1570 17170 -1550
rect 16980 -1575 16985 -1570
rect 16945 -1580 16985 -1575
rect 17165 -1575 17170 -1570
rect 17200 -1550 17205 -1545
rect 18395 -1545 18435 -1540
rect 18395 -1550 18400 -1545
rect 17200 -1570 18400 -1550
rect 17200 -1575 17205 -1570
rect 17165 -1580 17205 -1575
rect 18395 -1575 18400 -1570
rect 18430 -1550 18435 -1545
rect 18615 -1545 18655 -1540
rect 18615 -1550 18620 -1545
rect 18430 -1570 18620 -1550
rect 18430 -1575 18435 -1570
rect 18395 -1580 18435 -1575
rect 18615 -1575 18620 -1570
rect 18650 -1575 18655 -1545
rect 18615 -1580 18655 -1575
rect 15785 -1590 15825 -1585
rect 15785 -1620 15790 -1590
rect 15820 -1595 15825 -1590
rect 17055 -1590 17095 -1585
rect 17055 -1595 17060 -1590
rect 15820 -1615 17060 -1595
rect 15820 -1620 15825 -1615
rect 15785 -1625 15825 -1620
rect 17055 -1620 17060 -1615
rect 17090 -1620 17095 -1590
rect 17055 -1625 17095 -1620
rect 18505 -1590 18545 -1585
rect 18505 -1620 18510 -1590
rect 18540 -1595 18545 -1590
rect 19775 -1590 19815 -1585
rect 19775 -1595 19780 -1590
rect 18540 -1615 19780 -1595
rect 18540 -1620 18545 -1615
rect 18505 -1625 18545 -1620
rect 19775 -1620 19780 -1615
rect 19810 -1620 19815 -1590
rect 19775 -1625 19815 -1620
rect 16160 -1640 16200 -1635
rect 16160 -1670 16165 -1640
rect 16195 -1645 16200 -1640
rect 17585 -1640 17625 -1635
rect 17585 -1645 17590 -1640
rect 16195 -1665 17590 -1645
rect 16195 -1670 16200 -1665
rect 16160 -1675 16200 -1670
rect 17585 -1670 17590 -1665
rect 17620 -1670 17625 -1640
rect 17585 -1675 17625 -1670
rect 16105 -1685 16145 -1680
rect 16105 -1715 16110 -1685
rect 16140 -1690 16145 -1685
rect 17670 -1685 17710 -1680
rect 17670 -1690 17675 -1685
rect 16140 -1710 17675 -1690
rect 16140 -1715 16145 -1710
rect 16105 -1720 16145 -1715
rect 17670 -1715 17675 -1710
rect 17705 -1715 17710 -1685
rect 17670 -1720 17710 -1715
rect 17890 -1685 17930 -1680
rect 17890 -1715 17895 -1685
rect 17925 -1690 17930 -1685
rect 19535 -1685 19575 -1680
rect 19535 -1690 19540 -1685
rect 17925 -1710 19540 -1690
rect 17925 -1715 17930 -1710
rect 17890 -1720 17930 -1715
rect 19535 -1715 19540 -1710
rect 19570 -1715 19575 -1685
rect 19535 -1720 19575 -1715
rect 16155 -1760 16195 -1755
rect 16155 -1790 16160 -1760
rect 16190 -1765 16195 -1760
rect 19325 -1760 19365 -1755
rect 19325 -1765 19330 -1760
rect 16190 -1785 19330 -1765
rect 16190 -1790 16195 -1785
rect 16155 -1795 16195 -1790
rect 19325 -1790 19330 -1785
rect 19360 -1790 19365 -1760
rect 19325 -1795 19365 -1790
rect 17780 -1810 17820 -1805
rect 17780 -1840 17785 -1810
rect 17815 -1840 17820 -1810
rect 17780 -1845 17820 -1840
rect 16260 -1895 16300 -1890
rect 16260 -1925 16265 -1895
rect 16295 -1900 16300 -1895
rect 16480 -1895 16520 -1890
rect 16480 -1900 16485 -1895
rect 16295 -1920 16485 -1900
rect 16295 -1925 16300 -1920
rect 16260 -1930 16300 -1925
rect 16480 -1925 16485 -1920
rect 16515 -1900 16520 -1895
rect 16730 -1895 16770 -1890
rect 16730 -1900 16735 -1895
rect 16515 -1920 16735 -1900
rect 16515 -1925 16520 -1920
rect 16480 -1930 16520 -1925
rect 16730 -1925 16735 -1920
rect 16765 -1925 16770 -1895
rect 16730 -1930 16770 -1925
rect 17195 -1895 17235 -1890
rect 17195 -1925 17200 -1895
rect 17230 -1900 17235 -1895
rect 17425 -1900 17430 -1895
rect 17230 -1920 17430 -1900
rect 17230 -1925 17235 -1920
rect 17195 -1930 17235 -1925
rect 17425 -1930 17430 -1920
rect 17465 -1930 17470 -1895
rect 18124 -1930 18129 -1895
rect 18164 -1905 18169 -1895
rect 19080 -1900 19120 -1895
rect 19080 -1905 19085 -1900
rect 18164 -1925 19085 -1905
rect 18164 -1930 18169 -1925
rect 19080 -1930 19085 -1925
rect 19115 -1905 19120 -1900
rect 19460 -1900 19500 -1895
rect 19460 -1905 19465 -1900
rect 19115 -1925 19465 -1905
rect 19115 -1930 19120 -1925
rect 19080 -1935 19120 -1930
rect 19460 -1930 19465 -1925
rect 19495 -1930 19500 -1900
rect 19460 -1935 19500 -1930
rect 17195 -2015 17235 -2010
rect 17195 -2045 17200 -2015
rect 17230 -2020 17235 -2015
rect 18830 -2015 18870 -2010
rect 18830 -2020 18835 -2015
rect 17230 -2040 18835 -2020
rect 17230 -2045 17235 -2040
rect 17195 -2050 17235 -2045
rect 18830 -2045 18835 -2040
rect 18865 -2045 18870 -2015
rect 18830 -2050 18870 -2045
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2992 19440 -2987
rect 16160 -3025 16195 -3020
rect 19405 -3032 19440 -3027
rect 16160 -3065 16195 -3060
rect 16730 -3105 16770 -3100
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3120 15860 -3115
rect 15950 -3116 15985 -3111
rect 15855 -3140 15950 -3120
rect 15855 -3145 15860 -3140
rect 15820 -3150 15860 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3110 16770 -3105
rect 17780 -3105 17820 -3100
rect 17780 -3110 17785 -3105
rect 16765 -3130 17785 -3110
rect 16765 -3135 16770 -3130
rect 16730 -3140 16770 -3135
rect 17780 -3135 17785 -3130
rect 17815 -3135 17820 -3105
rect 17780 -3140 17820 -3135
rect 18615 -3105 18655 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3110 18655 -3105
rect 18830 -3105 18870 -3100
rect 18830 -3110 18835 -3105
rect 18650 -3130 18835 -3110
rect 18650 -3135 18655 -3130
rect 18615 -3140 18655 -3135
rect 18830 -3135 18835 -3130
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 15950 -3156 15985 -3151
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 16540 -4035 16580 -4030
rect 16540 -4065 16545 -4035
rect 16575 -4065 16580 -4035
rect 16540 -4070 16580 -4065
rect 15595 -4190 15635 -4185
rect 15595 -4220 15600 -4190
rect 15630 -4195 15635 -4190
rect 16280 -4190 16320 -4185
rect 16280 -4195 16285 -4190
rect 15630 -4215 16285 -4195
rect 15630 -4220 15635 -4215
rect 15595 -4225 15635 -4220
rect 16280 -4220 16285 -4215
rect 16315 -4195 16320 -4190
rect 16540 -4190 16580 -4185
rect 16540 -4195 16545 -4190
rect 16315 -4215 16545 -4195
rect 16315 -4220 16320 -4215
rect 16280 -4225 16320 -4220
rect 16540 -4220 16545 -4215
rect 16575 -4195 16580 -4190
rect 16605 -4190 16645 -4185
rect 16605 -4195 16610 -4190
rect 16575 -4215 16610 -4195
rect 16575 -4220 16580 -4215
rect 16540 -4225 16580 -4220
rect 16605 -4220 16610 -4215
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4270 15860 -4265
rect 17250 -4265 17300 -4255
rect 17250 -4270 17260 -4265
rect 15855 -4290 17260 -4270
rect 15855 -4295 15860 -4290
rect 15820 -4300 15860 -4295
rect 17250 -4295 17260 -4290
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4270 17820 -4265
rect 18955 -4265 18995 -4260
rect 18955 -4270 18960 -4265
rect 17815 -4290 18960 -4270
rect 17815 -4295 17820 -4290
rect 17780 -4300 17820 -4295
rect 18955 -4295 18960 -4290
rect 18990 -4270 18995 -4265
rect 19280 -4265 19320 -4260
rect 19280 -4270 19285 -4265
rect 18990 -4290 19285 -4270
rect 18990 -4295 18995 -4290
rect 18955 -4300 18995 -4295
rect 19280 -4295 19285 -4290
rect 19315 -4270 19320 -4265
rect 19965 -4265 20005 -4260
rect 19965 -4270 19970 -4265
rect 19315 -4290 19970 -4270
rect 19315 -4295 19320 -4290
rect 19280 -4300 19320 -4295
rect 19965 -4295 19970 -4290
rect 20000 -4295 20005 -4265
rect 19965 -4300 20005 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4320 15765 -4315
rect 16900 -4315 16950 -4305
rect 16900 -4320 16910 -4315
rect 15760 -4340 16910 -4320
rect 15760 -4345 15765 -4340
rect 15725 -4350 15765 -4345
rect 16900 -4345 16910 -4340
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4320 18700 -4315
rect 19730 -4315 19770 -4310
rect 19730 -4320 19735 -4315
rect 18690 -4340 19735 -4320
rect 18690 -4345 18700 -4340
rect 18650 -4355 18700 -4345
rect 19730 -4345 19735 -4340
rect 19765 -4345 19770 -4315
rect 19730 -4350 19770 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4365 15990 -4360
rect 16205 -4360 16245 -4355
rect 16205 -4365 16210 -4360
rect 15985 -4385 16210 -4365
rect 15985 -4390 15990 -4385
rect 15950 -4395 15990 -4390
rect 16205 -4390 16210 -4385
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4365 19395 -4360
rect 19610 -4360 19650 -4355
rect 19610 -4365 19615 -4360
rect 19390 -4385 19615 -4365
rect 19390 -4390 19395 -4385
rect 19355 -4395 19395 -4390
rect 19610 -4390 19615 -4385
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4415 17995 -4410
rect 20050 -4410 20090 -4405
rect 20050 -4415 20055 -4410
rect 17990 -4435 20055 -4415
rect 17990 -4440 17995 -4435
rect 17955 -4445 17995 -4440
rect 20050 -4440 20055 -4435
rect 20085 -4440 20090 -4410
rect 20050 -4445 20090 -4440
<< via2 >>
rect 20055 1250 20085 1280
rect 20055 785 20085 815
rect 20055 155 20085 185
rect 20055 -560 20085 -530
rect 19970 -875 20000 -845
rect 19970 -1110 20000 -1080
rect 19970 -1300 20000 -1270
rect 15600 -4220 15630 -4190
rect 17260 -4295 17290 -4265
rect 19970 -4295 20000 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 17960 -4440 17990 -4410
rect 20055 -4440 20085 -4410
<< metal3 >>
rect 15505 1545 15555 1550
rect 15505 1505 15510 1545
rect 15550 1505 15555 1545
rect 15505 1500 15555 1505
rect 20045 1545 20095 1550
rect 20045 1505 20050 1545
rect 20090 1505 20095 1545
rect 20045 1500 20095 1505
rect 15510 -6245 15550 1500
rect 15590 1460 15640 1465
rect 15590 1420 15595 1460
rect 15635 1420 15640 1460
rect 15590 1415 15640 1420
rect 19960 1460 20010 1465
rect 19960 1420 19965 1460
rect 20005 1420 20010 1460
rect 19960 1415 20010 1420
rect 15595 -4190 15635 1415
rect 15595 -4220 15600 -4190
rect 15630 -4220 15635 -4190
rect 15595 -6165 15635 -4220
rect 19965 -845 20005 1415
rect 19965 -875 19970 -845
rect 20000 -875 20005 -845
rect 19965 -1080 20005 -875
rect 19965 -1110 19970 -1080
rect 20000 -1110 20005 -1080
rect 19965 -1270 20005 -1110
rect 19965 -1300 19970 -1270
rect 20000 -1300 20005 -1270
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 17250 -4305 17300 -4300
rect 19965 -4265 20005 -1300
rect 19965 -4295 19970 -4265
rect 20000 -4295 20005 -4265
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4355 16950 -4350
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4355 18700 -4350
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4520 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4520 17995 -4440
rect 19355 -4520 19395 -4390
rect 15760 -4615 15990 -4520
rect 16110 -4615 16340 -4520
rect 16460 -4615 16690 -4520
rect 16810 -4615 17040 -4520
rect 15760 -4665 17040 -4615
rect 15760 -4750 15990 -4665
rect 16110 -4750 16340 -4665
rect 16460 -4750 16690 -4665
rect 16810 -4750 17040 -4665
rect 17160 -4615 17390 -4520
rect 17510 -4615 17740 -4520
rect 17860 -4615 18090 -4520
rect 18210 -4615 18440 -4520
rect 17160 -4665 18440 -4615
rect 17160 -4750 17390 -4665
rect 17510 -4750 17740 -4665
rect 17860 -4750 18090 -4665
rect 18210 -4750 18440 -4665
rect 18560 -4615 18790 -4520
rect 18910 -4615 19140 -4520
rect 19260 -4615 19490 -4520
rect 19610 -4615 19840 -4520
rect 18560 -4665 19840 -4615
rect 18560 -4750 18790 -4665
rect 18910 -4750 19140 -4665
rect 19260 -4750 19490 -4665
rect 19610 -4750 19840 -4665
rect 16200 -4870 16250 -4750
rect 17950 -4870 18000 -4750
rect 19350 -4870 19400 -4750
rect 15760 -4965 15990 -4870
rect 16110 -4965 16340 -4870
rect 16460 -4965 16690 -4870
rect 16810 -4965 17040 -4870
rect 15760 -5015 17040 -4965
rect 15760 -5100 15990 -5015
rect 16110 -5100 16340 -5015
rect 16460 -5100 16690 -5015
rect 16810 -5100 17040 -5015
rect 17160 -4965 17390 -4870
rect 17510 -4965 17740 -4870
rect 17860 -4965 18090 -4870
rect 18210 -4965 18440 -4870
rect 17160 -5015 18440 -4965
rect 17160 -5100 17390 -5015
rect 17510 -5100 17740 -5015
rect 17860 -5100 18090 -5015
rect 18210 -5100 18440 -5015
rect 18560 -4965 18790 -4870
rect 18910 -4965 19140 -4870
rect 19260 -4965 19490 -4870
rect 19610 -4965 19840 -4870
rect 18560 -5015 19840 -4965
rect 18560 -5100 18790 -5015
rect 18910 -5100 19140 -5015
rect 19260 -5100 19490 -5015
rect 19610 -5100 19840 -5015
rect 16200 -5220 16250 -5100
rect 17950 -5220 18000 -5100
rect 19350 -5220 19400 -5100
rect 15760 -5315 15990 -5220
rect 16110 -5315 16340 -5220
rect 16460 -5315 16690 -5220
rect 16810 -5315 17040 -5220
rect 15760 -5365 17040 -5315
rect 15760 -5450 15990 -5365
rect 16110 -5450 16340 -5365
rect 16460 -5450 16690 -5365
rect 16810 -5450 17040 -5365
rect 17160 -5315 17390 -5220
rect 17510 -5315 17740 -5220
rect 17860 -5315 18090 -5220
rect 18210 -5315 18440 -5220
rect 17160 -5365 18440 -5315
rect 17160 -5450 17390 -5365
rect 17510 -5450 17740 -5365
rect 17860 -5450 18090 -5365
rect 18210 -5450 18440 -5365
rect 18560 -5315 18790 -5220
rect 18910 -5315 19140 -5220
rect 19260 -5315 19490 -5220
rect 19610 -5315 19840 -5220
rect 18560 -5365 19840 -5315
rect 18560 -5450 18790 -5365
rect 18910 -5450 19140 -5365
rect 19260 -5450 19490 -5365
rect 19610 -5450 19840 -5365
rect 16200 -5570 16250 -5450
rect 17950 -5570 18000 -5450
rect 19350 -5570 19400 -5450
rect 15760 -5665 15990 -5570
rect 16110 -5665 16340 -5570
rect 16460 -5665 16690 -5570
rect 16810 -5665 17040 -5570
rect 15760 -5715 17040 -5665
rect 15760 -5800 15990 -5715
rect 16110 -5800 16340 -5715
rect 16460 -5800 16690 -5715
rect 16810 -5800 17040 -5715
rect 17160 -5665 17390 -5570
rect 17510 -5665 17740 -5570
rect 17860 -5665 18090 -5570
rect 18210 -5665 18440 -5570
rect 17160 -5715 18440 -5665
rect 17160 -5800 17390 -5715
rect 17510 -5800 17740 -5715
rect 17860 -5800 18090 -5715
rect 18210 -5800 18440 -5715
rect 18560 -5665 18790 -5570
rect 18910 -5665 19140 -5570
rect 19260 -5665 19490 -5570
rect 19610 -5665 19840 -5570
rect 18560 -5715 19840 -5665
rect 18560 -5800 18790 -5715
rect 18910 -5800 19140 -5715
rect 19260 -5800 19490 -5715
rect 19610 -5800 19840 -5715
rect 16200 -5920 16250 -5800
rect 17950 -5920 18000 -5800
rect 19350 -5920 19400 -5800
rect 15760 -6015 15990 -5920
rect 16110 -6015 16340 -5920
rect 16460 -6015 16690 -5920
rect 16810 -6015 17040 -5920
rect 15760 -6065 17040 -6015
rect 15760 -6150 15990 -6065
rect 16110 -6150 16340 -6065
rect 16460 -6150 16690 -6065
rect 16810 -6150 17040 -6065
rect 17160 -6015 17390 -5920
rect 17510 -6015 17740 -5920
rect 17860 -6015 18090 -5920
rect 18210 -6015 18440 -5920
rect 17160 -6065 18440 -6015
rect 17160 -6150 17390 -6065
rect 17510 -6150 17740 -6065
rect 17860 -6150 18090 -6065
rect 18210 -6150 18440 -6065
rect 18560 -6015 18790 -5920
rect 18910 -6015 19140 -5920
rect 19260 -6015 19490 -5920
rect 19610 -6015 19840 -5920
rect 18560 -6065 19840 -6015
rect 18560 -6150 18790 -6065
rect 18910 -6150 19140 -6065
rect 19260 -6150 19490 -6065
rect 19610 -6150 19840 -6065
rect 19965 -6165 20005 -4295
rect 20050 1280 20090 1500
rect 20050 1250 20055 1280
rect 20085 1250 20090 1280
rect 20050 815 20090 1250
rect 20050 785 20055 815
rect 20085 785 20090 815
rect 20050 185 20090 785
rect 20050 155 20055 185
rect 20085 155 20090 185
rect 20050 -530 20090 155
rect 20050 -560 20055 -530
rect 20085 -560 20090 -530
rect 20050 -4410 20090 -560
rect 20050 -4440 20055 -4410
rect 20085 -4440 20090 -4410
rect 15590 -6170 15640 -6165
rect 15590 -6210 15595 -6170
rect 15635 -6210 15640 -6170
rect 15590 -6215 15640 -6210
rect 19960 -6170 20010 -6165
rect 19960 -6210 19965 -6170
rect 20005 -6210 20010 -6170
rect 19960 -6215 20010 -6210
rect 20050 -6245 20090 -4440
rect 15505 -6250 15555 -6245
rect 15505 -6290 15510 -6250
rect 15550 -6290 15555 -6250
rect 15505 -6295 15555 -6290
rect 20045 -6250 20095 -6245
rect 20045 -6290 20050 -6250
rect 20090 -6290 20095 -6250
rect 20045 -6295 20095 -6290
<< via3 >>
rect 15510 1505 15550 1545
rect 20050 1505 20090 1545
rect 15595 1420 15635 1460
rect 19965 1420 20005 1460
rect 17255 -4265 17295 -4260
rect 17255 -4295 17260 -4265
rect 17260 -4295 17290 -4265
rect 17290 -4295 17295 -4265
rect 17255 -4300 17295 -4295
rect 16905 -4315 16945 -4310
rect 16905 -4345 16910 -4315
rect 16910 -4345 16940 -4315
rect 16940 -4345 16945 -4315
rect 16905 -4350 16945 -4345
rect 18655 -4315 18695 -4310
rect 18655 -4345 18660 -4315
rect 18660 -4345 18690 -4315
rect 18690 -4345 18695 -4315
rect 18655 -4350 18695 -4345
rect 15595 -6210 15635 -6170
rect 19965 -6210 20005 -6170
rect 15510 -6290 15550 -6250
rect 20050 -6290 20090 -6250
<< mimcap >>
rect 15775 -4620 15975 -4535
rect 15775 -4660 15855 -4620
rect 15895 -4660 15975 -4620
rect 15775 -4735 15975 -4660
rect 16125 -4620 16325 -4535
rect 16125 -4660 16205 -4620
rect 16245 -4660 16325 -4620
rect 16125 -4735 16325 -4660
rect 16475 -4620 16675 -4535
rect 16475 -4660 16555 -4620
rect 16595 -4660 16675 -4620
rect 16475 -4735 16675 -4660
rect 16825 -4620 17025 -4535
rect 16825 -4660 16905 -4620
rect 16945 -4660 17025 -4620
rect 16825 -4735 17025 -4660
rect 17175 -4620 17375 -4535
rect 17175 -4660 17255 -4620
rect 17295 -4660 17375 -4620
rect 17175 -4735 17375 -4660
rect 17525 -4620 17725 -4535
rect 17525 -4660 17605 -4620
rect 17645 -4660 17725 -4620
rect 17525 -4735 17725 -4660
rect 17875 -4620 18075 -4535
rect 17875 -4660 17955 -4620
rect 17995 -4660 18075 -4620
rect 17875 -4735 18075 -4660
rect 18225 -4620 18425 -4535
rect 18225 -4660 18305 -4620
rect 18345 -4660 18425 -4620
rect 18225 -4735 18425 -4660
rect 18575 -4620 18775 -4535
rect 18575 -4660 18655 -4620
rect 18695 -4660 18775 -4620
rect 18575 -4735 18775 -4660
rect 18925 -4620 19125 -4535
rect 18925 -4660 19005 -4620
rect 19045 -4660 19125 -4620
rect 18925 -4735 19125 -4660
rect 19275 -4620 19475 -4535
rect 19275 -4660 19355 -4620
rect 19395 -4660 19475 -4620
rect 19275 -4735 19475 -4660
rect 19625 -4620 19825 -4535
rect 19625 -4660 19705 -4620
rect 19745 -4660 19825 -4620
rect 19625 -4735 19825 -4660
rect 15775 -4970 15975 -4885
rect 15775 -5010 15855 -4970
rect 15895 -5010 15975 -4970
rect 15775 -5085 15975 -5010
rect 16125 -4970 16325 -4885
rect 16125 -5010 16205 -4970
rect 16245 -5010 16325 -4970
rect 16125 -5085 16325 -5010
rect 16475 -4970 16675 -4885
rect 16475 -5010 16555 -4970
rect 16595 -5010 16675 -4970
rect 16475 -5085 16675 -5010
rect 16825 -4970 17025 -4885
rect 16825 -5010 16905 -4970
rect 16945 -5010 17025 -4970
rect 16825 -5085 17025 -5010
rect 17175 -4970 17375 -4885
rect 17175 -5010 17255 -4970
rect 17295 -5010 17375 -4970
rect 17175 -5085 17375 -5010
rect 17525 -4970 17725 -4885
rect 17525 -5010 17605 -4970
rect 17645 -5010 17725 -4970
rect 17525 -5085 17725 -5010
rect 17875 -4970 18075 -4885
rect 17875 -5010 17955 -4970
rect 17995 -5010 18075 -4970
rect 17875 -5085 18075 -5010
rect 18225 -4970 18425 -4885
rect 18225 -5010 18305 -4970
rect 18345 -5010 18425 -4970
rect 18225 -5085 18425 -5010
rect 18575 -4970 18775 -4885
rect 18575 -5010 18655 -4970
rect 18695 -5010 18775 -4970
rect 18575 -5085 18775 -5010
rect 18925 -4970 19125 -4885
rect 18925 -5010 19005 -4970
rect 19045 -5010 19125 -4970
rect 18925 -5085 19125 -5010
rect 19275 -4970 19475 -4885
rect 19275 -5010 19355 -4970
rect 19395 -5010 19475 -4970
rect 19275 -5085 19475 -5010
rect 19625 -4970 19825 -4885
rect 19625 -5010 19705 -4970
rect 19745 -5010 19825 -4970
rect 19625 -5085 19825 -5010
rect 15775 -5320 15975 -5235
rect 15775 -5360 15855 -5320
rect 15895 -5360 15975 -5320
rect 15775 -5435 15975 -5360
rect 16125 -5320 16325 -5235
rect 16125 -5360 16205 -5320
rect 16245 -5360 16325 -5320
rect 16125 -5435 16325 -5360
rect 16475 -5320 16675 -5235
rect 16475 -5360 16555 -5320
rect 16595 -5360 16675 -5320
rect 16475 -5435 16675 -5360
rect 16825 -5320 17025 -5235
rect 16825 -5360 16905 -5320
rect 16945 -5360 17025 -5320
rect 16825 -5435 17025 -5360
rect 17175 -5320 17375 -5235
rect 17175 -5360 17255 -5320
rect 17295 -5360 17375 -5320
rect 17175 -5435 17375 -5360
rect 17525 -5320 17725 -5235
rect 17525 -5360 17605 -5320
rect 17645 -5360 17725 -5320
rect 17525 -5435 17725 -5360
rect 17875 -5320 18075 -5235
rect 17875 -5360 17955 -5320
rect 17995 -5360 18075 -5320
rect 17875 -5435 18075 -5360
rect 18225 -5320 18425 -5235
rect 18225 -5360 18305 -5320
rect 18345 -5360 18425 -5320
rect 18225 -5435 18425 -5360
rect 18575 -5320 18775 -5235
rect 18575 -5360 18655 -5320
rect 18695 -5360 18775 -5320
rect 18575 -5435 18775 -5360
rect 18925 -5320 19125 -5235
rect 18925 -5360 19005 -5320
rect 19045 -5360 19125 -5320
rect 18925 -5435 19125 -5360
rect 19275 -5320 19475 -5235
rect 19275 -5360 19355 -5320
rect 19395 -5360 19475 -5320
rect 19275 -5435 19475 -5360
rect 19625 -5320 19825 -5235
rect 19625 -5360 19705 -5320
rect 19745 -5360 19825 -5320
rect 19625 -5435 19825 -5360
rect 15775 -5670 15975 -5585
rect 15775 -5710 15855 -5670
rect 15895 -5710 15975 -5670
rect 15775 -5785 15975 -5710
rect 16125 -5670 16325 -5585
rect 16125 -5710 16205 -5670
rect 16245 -5710 16325 -5670
rect 16125 -5785 16325 -5710
rect 16475 -5670 16675 -5585
rect 16475 -5710 16555 -5670
rect 16595 -5710 16675 -5670
rect 16475 -5785 16675 -5710
rect 16825 -5670 17025 -5585
rect 16825 -5710 16905 -5670
rect 16945 -5710 17025 -5670
rect 16825 -5785 17025 -5710
rect 17175 -5670 17375 -5585
rect 17175 -5710 17255 -5670
rect 17295 -5710 17375 -5670
rect 17175 -5785 17375 -5710
rect 17525 -5670 17725 -5585
rect 17525 -5710 17605 -5670
rect 17645 -5710 17725 -5670
rect 17525 -5785 17725 -5710
rect 17875 -5670 18075 -5585
rect 17875 -5710 17955 -5670
rect 17995 -5710 18075 -5670
rect 17875 -5785 18075 -5710
rect 18225 -5670 18425 -5585
rect 18225 -5710 18305 -5670
rect 18345 -5710 18425 -5670
rect 18225 -5785 18425 -5710
rect 18575 -5670 18775 -5585
rect 18575 -5710 18655 -5670
rect 18695 -5710 18775 -5670
rect 18575 -5785 18775 -5710
rect 18925 -5670 19125 -5585
rect 18925 -5710 19005 -5670
rect 19045 -5710 19125 -5670
rect 18925 -5785 19125 -5710
rect 19275 -5670 19475 -5585
rect 19275 -5710 19355 -5670
rect 19395 -5710 19475 -5670
rect 19275 -5785 19475 -5710
rect 19625 -5670 19825 -5585
rect 19625 -5710 19705 -5670
rect 19745 -5710 19825 -5670
rect 19625 -5785 19825 -5710
rect 15775 -6020 15975 -5935
rect 15775 -6060 15855 -6020
rect 15895 -6060 15975 -6020
rect 15775 -6135 15975 -6060
rect 16125 -6020 16325 -5935
rect 16125 -6060 16205 -6020
rect 16245 -6060 16325 -6020
rect 16125 -6135 16325 -6060
rect 16475 -6020 16675 -5935
rect 16475 -6060 16555 -6020
rect 16595 -6060 16675 -6020
rect 16475 -6135 16675 -6060
rect 16825 -6020 17025 -5935
rect 16825 -6060 16905 -6020
rect 16945 -6060 17025 -6020
rect 16825 -6135 17025 -6060
rect 17175 -6020 17375 -5935
rect 17175 -6060 17255 -6020
rect 17295 -6060 17375 -6020
rect 17175 -6135 17375 -6060
rect 17525 -6020 17725 -5935
rect 17525 -6060 17605 -6020
rect 17645 -6060 17725 -6020
rect 17525 -6135 17725 -6060
rect 17875 -6020 18075 -5935
rect 17875 -6060 17955 -6020
rect 17995 -6060 18075 -6020
rect 17875 -6135 18075 -6060
rect 18225 -6020 18425 -5935
rect 18225 -6060 18305 -6020
rect 18345 -6060 18425 -6020
rect 18225 -6135 18425 -6060
rect 18575 -6020 18775 -5935
rect 18575 -6060 18655 -6020
rect 18695 -6060 18775 -6020
rect 18575 -6135 18775 -6060
rect 18925 -6020 19125 -5935
rect 18925 -6060 19005 -6020
rect 19045 -6060 19125 -6020
rect 18925 -6135 19125 -6060
rect 19275 -6020 19475 -5935
rect 19275 -6060 19355 -6020
rect 19395 -6060 19475 -6020
rect 19275 -6135 19475 -6060
rect 19625 -6020 19825 -5935
rect 19625 -6060 19705 -6020
rect 19745 -6060 19825 -6020
rect 19625 -6135 19825 -6060
<< mimcapcontact >>
rect 15855 -4660 15895 -4620
rect 16205 -4660 16245 -4620
rect 16555 -4660 16595 -4620
rect 16905 -4660 16945 -4620
rect 17255 -4660 17295 -4620
rect 17605 -4660 17645 -4620
rect 17955 -4660 17995 -4620
rect 18305 -4660 18345 -4620
rect 18655 -4660 18695 -4620
rect 19005 -4660 19045 -4620
rect 19355 -4660 19395 -4620
rect 19705 -4660 19745 -4620
rect 15855 -5010 15895 -4970
rect 16205 -5010 16245 -4970
rect 16555 -5010 16595 -4970
rect 16905 -5010 16945 -4970
rect 17255 -5010 17295 -4970
rect 17605 -5010 17645 -4970
rect 17955 -5010 17995 -4970
rect 18305 -5010 18345 -4970
rect 18655 -5010 18695 -4970
rect 19005 -5010 19045 -4970
rect 19355 -5010 19395 -4970
rect 19705 -5010 19745 -4970
rect 15855 -5360 15895 -5320
rect 16205 -5360 16245 -5320
rect 16555 -5360 16595 -5320
rect 16905 -5360 16945 -5320
rect 17255 -5360 17295 -5320
rect 17605 -5360 17645 -5320
rect 17955 -5360 17995 -5320
rect 18305 -5360 18345 -5320
rect 18655 -5360 18695 -5320
rect 19005 -5360 19045 -5320
rect 19355 -5360 19395 -5320
rect 19705 -5360 19745 -5320
rect 15855 -5710 15895 -5670
rect 16205 -5710 16245 -5670
rect 16555 -5710 16595 -5670
rect 16905 -5710 16945 -5670
rect 17255 -5710 17295 -5670
rect 17605 -5710 17645 -5670
rect 17955 -5710 17995 -5670
rect 18305 -5710 18345 -5670
rect 18655 -5710 18695 -5670
rect 19005 -5710 19045 -5670
rect 19355 -5710 19395 -5670
rect 19705 -5710 19745 -5670
rect 15855 -6060 15895 -6020
rect 16205 -6060 16245 -6020
rect 16555 -6060 16595 -6020
rect 16905 -6060 16945 -6020
rect 17255 -6060 17295 -6020
rect 17605 -6060 17645 -6020
rect 17955 -6060 17995 -6020
rect 18305 -6060 18345 -6020
rect 18655 -6060 18695 -6020
rect 19005 -6060 19045 -6020
rect 19355 -6060 19395 -6020
rect 19705 -6060 19745 -6020
<< metal4 >>
rect 15505 1545 20095 1550
rect 15505 1505 15510 1545
rect 15550 1505 20050 1545
rect 20090 1505 20095 1545
rect 15505 1500 20095 1505
rect 15590 1460 20010 1465
rect 15590 1420 15595 1460
rect 15635 1420 19965 1460
rect 20005 1420 20010 1460
rect 15590 1415 20010 1420
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4615 16950 -4350
rect 15850 -4620 16950 -4615
rect 15850 -4660 15855 -4620
rect 15895 -4660 16205 -4620
rect 16245 -4660 16555 -4620
rect 16595 -4660 16905 -4620
rect 16945 -4660 16950 -4620
rect 15850 -4665 16950 -4660
rect 17250 -4615 17300 -4300
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4615 18700 -4350
rect 17250 -4620 18350 -4615
rect 17250 -4660 17255 -4620
rect 17295 -4660 17605 -4620
rect 17645 -4660 17955 -4620
rect 17995 -4660 18305 -4620
rect 18345 -4660 18350 -4620
rect 17250 -4665 18350 -4660
rect 18650 -4620 19750 -4615
rect 18650 -4660 18655 -4620
rect 18695 -4660 19005 -4620
rect 19045 -4660 19355 -4620
rect 19395 -4660 19705 -4620
rect 19745 -4660 19750 -4620
rect 18650 -4665 19750 -4660
rect 16200 -4965 16250 -4665
rect 17950 -4965 18000 -4665
rect 19350 -4965 19400 -4665
rect 15850 -4970 16950 -4965
rect 15850 -5010 15855 -4970
rect 15895 -5010 16205 -4970
rect 16245 -5010 16555 -4970
rect 16595 -5010 16905 -4970
rect 16945 -5010 16950 -4970
rect 15850 -5015 16950 -5010
rect 17250 -4970 18350 -4965
rect 17250 -5010 17255 -4970
rect 17295 -5010 17605 -4970
rect 17645 -5010 17955 -4970
rect 17995 -5010 18305 -4970
rect 18345 -5010 18350 -4970
rect 17250 -5015 18350 -5010
rect 18650 -4970 19750 -4965
rect 18650 -5010 18655 -4970
rect 18695 -5010 19005 -4970
rect 19045 -5010 19355 -4970
rect 19395 -5010 19705 -4970
rect 19745 -5010 19750 -4970
rect 18650 -5015 19750 -5010
rect 16200 -5315 16250 -5015
rect 17950 -5315 18000 -5015
rect 19350 -5315 19400 -5015
rect 15850 -5320 16950 -5315
rect 15850 -5360 15855 -5320
rect 15895 -5360 16205 -5320
rect 16245 -5360 16555 -5320
rect 16595 -5360 16905 -5320
rect 16945 -5360 16950 -5320
rect 15850 -5365 16950 -5360
rect 17250 -5320 18350 -5315
rect 17250 -5360 17255 -5320
rect 17295 -5360 17605 -5320
rect 17645 -5360 17955 -5320
rect 17995 -5360 18305 -5320
rect 18345 -5360 18350 -5320
rect 17250 -5365 18350 -5360
rect 18650 -5320 19750 -5315
rect 18650 -5360 18655 -5320
rect 18695 -5360 19005 -5320
rect 19045 -5360 19355 -5320
rect 19395 -5360 19705 -5320
rect 19745 -5360 19750 -5320
rect 18650 -5365 19750 -5360
rect 16200 -5665 16250 -5365
rect 17950 -5665 18000 -5365
rect 19350 -5665 19400 -5365
rect 15850 -5670 16950 -5665
rect 15850 -5710 15855 -5670
rect 15895 -5710 16205 -5670
rect 16245 -5710 16555 -5670
rect 16595 -5710 16905 -5670
rect 16945 -5710 16950 -5670
rect 15850 -5715 16950 -5710
rect 17250 -5670 18350 -5665
rect 17250 -5710 17255 -5670
rect 17295 -5710 17605 -5670
rect 17645 -5710 17955 -5670
rect 17995 -5710 18305 -5670
rect 18345 -5710 18350 -5670
rect 17250 -5715 18350 -5710
rect 18650 -5670 19750 -5665
rect 18650 -5710 18655 -5670
rect 18695 -5710 19005 -5670
rect 19045 -5710 19355 -5670
rect 19395 -5710 19705 -5670
rect 19745 -5710 19750 -5670
rect 18650 -5715 19750 -5710
rect 16200 -6015 16250 -5715
rect 17950 -6015 18000 -5715
rect 19350 -6015 19400 -5715
rect 15850 -6020 16950 -6015
rect 15850 -6060 15855 -6020
rect 15895 -6060 16205 -6020
rect 16245 -6060 16555 -6020
rect 16595 -6060 16905 -6020
rect 16945 -6060 16950 -6020
rect 15850 -6065 16950 -6060
rect 17250 -6020 18350 -6015
rect 17250 -6060 17255 -6020
rect 17295 -6060 17605 -6020
rect 17645 -6060 17955 -6020
rect 17995 -6060 18305 -6020
rect 18345 -6060 18350 -6020
rect 17250 -6065 18350 -6060
rect 18650 -6020 19750 -6015
rect 18650 -6060 18655 -6020
rect 18695 -6060 19005 -6020
rect 19045 -6060 19355 -6020
rect 19395 -6060 19705 -6020
rect 19745 -6060 19750 -6020
rect 18650 -6065 19750 -6060
rect 15590 -6170 20010 -6165
rect 15590 -6210 15595 -6170
rect 15635 -6210 19965 -6170
rect 20005 -6210 20010 -6170
rect 15590 -6215 20010 -6210
rect 15505 -6250 20095 -6245
rect 15505 -6290 15510 -6250
rect 15550 -6290 20050 -6250
rect 20090 -6290 20095 -6250
rect 15505 -6295 20095 -6290
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel poly 18430 440 18430 440 5 FreeSans 400 0 0 -40 V_TOP
flabel metal1 18780 -1010 18780 -1010 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 18930 -375 18930 -375 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 18980 -80 18980 -80 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 16670 -375 16670 -375 1 FreeSans 400 0 0 80 Vin+
flabel metal2 16665 -230 16665 -230 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 18030 -120 18030 -120 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 18170 -465 18170 -465 7 FreeSans 400 0 -200 0 V_p_2
flabel metal2 17430 -465 17430 -465 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 16620 -80 16620 -80 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 17570 -120 17570 -120 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal1 16190 -1255 16190 -1255 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal1 16235 -795 16235 -795 3 FreeSans 400 0 200 0 START_UP
flabel metal2 15995 -4385 15995 -4385 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19355 -4375 19355 -4375 7 FreeSans 400 180 -40 0 cap_res2
flabel metal3 20005 925 20005 925 3 FreeSans 400 0 200 0 GNDA
port 12 e
flabel metal1 16125 1595 16125 1595 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 19280 1595 19280 1595 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
flabel metal1 19795 1595 19795 1595 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16040 1585 16040 1585 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 19415 1590 19415 1590 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 19565 1590 19565 1590 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel metal1 15805 1595 15805 1595 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal1 17750 1595 17750 1595 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 17105 1595 17105 1595 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
flabel metal1 18495 1595 18495 1595 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal3 20090 1150 20090 1150 3 FreeSans 400 0 200 0 VDDA
port 1 e
flabel via1 17855 1335 17855 1335 1 FreeSans 400 0 0 200 PFET_GATE_10uA
<< end >>
