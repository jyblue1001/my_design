** sch_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/tb_buck_converter.sch
**.subckt tb_buck_converter
V1 net2 GND 25
R48 vout GND 1 m=1
D1 GND net1 D1N914 area=1
L1 vout net1 30u m=1
C1 net3 GND 250u m=1
R1 vout net3 0.05 m=1
V2 net4 GND pulse(0 1.8 0ns 10ps 10ps 19.2ns 50ns)
S1 net2 net1 net4 GND SW1
**** begin user architecture code



.options method=gear
.options wnflag=1
* .options savecurrents


.model D1N914 D(Is=168.1E-21 N=1 Rs=.1 Ikf=1 Xti=3 Eg=1.11 Cjo=4p M=.3333 Vj=.75 Fc=.5 Bv=100 Ibv=100u Tt=11.54n)


.control
  * save all
  save v(vout)
  * dc V1 0.0 2.0 0.005
  tran 100us 2ms
  remzerovec
  write tb_buck_converter.raw
  set appendwrite

.endc




**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code
.MODEL SW1 SW( VT=0.9 VH=0.01 RON=0.01 ROFF=10G )
**** end user architecture code
.end
