magic
tech sky130A
timestamp 1738174613
<< nwell >>
rect -3570 220 -1745 460
rect -1550 230 460 370
<< pwell >>
rect -3030 5 -2825 115
rect -2575 5 -2370 115
rect -2115 5 -1910 115
<< nmos >>
rect -3500 10 -3485 110
rect -3350 10 -3335 110
rect -3200 10 -3185 110
rect -2975 10 -2960 110
rect -2750 10 -2735 110
rect -2520 10 -2505 110
rect -2290 10 -2275 110
rect -2060 10 -2045 110
rect -1830 10 -1815 110
rect -1430 0 -1370 100
rect -1320 0 -1260 100
rect -1210 0 -1150 100
rect -1100 0 -1040 100
rect -770 0 -710 100
rect -660 0 -600 100
rect -550 0 -490 100
rect -440 0 -380 100
rect 0 0 60 100
rect 110 0 170 100
rect 220 0 280 100
rect 330 0 390 100
<< pmos >>
rect -3500 240 -3485 440
rect -3350 240 -3335 440
rect -3200 240 -3185 440
rect -2975 240 -2960 440
rect -2750 240 -2735 440
rect -2520 240 -2505 440
rect -2290 240 -2275 440
rect -2060 240 -2045 440
rect -1830 240 -1815 440
rect -1480 250 -1420 350
rect -1370 250 -1310 350
rect -1260 250 -1200 350
rect -1150 250 -1090 350
rect -1040 250 -980 350
rect -930 250 -870 350
rect -820 250 -760 350
rect -710 250 -650 350
rect -440 250 -380 350
rect -330 250 -270 350
rect -220 250 -160 350
rect -110 250 -50 350
rect 0 250 60 350
rect 110 250 170 350
rect 220 250 280 350
rect 330 250 390 350
<< ndiff >>
rect -3550 95 -3500 110
rect -3550 25 -3535 95
rect -3515 25 -3500 95
rect -3550 10 -3500 25
rect -3485 95 -3435 110
rect -3485 25 -3470 95
rect -3450 25 -3435 95
rect -3485 10 -3435 25
rect -3400 95 -3350 110
rect -3400 25 -3385 95
rect -3365 25 -3350 95
rect -3400 10 -3350 25
rect -3335 95 -3285 110
rect -3335 25 -3320 95
rect -3300 25 -3285 95
rect -3335 10 -3285 25
rect -3250 95 -3200 110
rect -3250 25 -3235 95
rect -3215 25 -3200 95
rect -3250 10 -3200 25
rect -3185 95 -3135 110
rect -3185 25 -3170 95
rect -3150 25 -3135 95
rect -3025 95 -2975 110
rect -3185 10 -3135 25
rect -3025 25 -3010 95
rect -2990 25 -2975 95
rect -3025 10 -2975 25
rect -2960 95 -2910 110
rect -2960 25 -2945 95
rect -2925 25 -2910 95
rect -2960 10 -2910 25
rect -2800 95 -2750 110
rect -2800 25 -2785 95
rect -2765 25 -2750 95
rect -2800 10 -2750 25
rect -2735 95 -2685 110
rect -2735 25 -2720 95
rect -2700 25 -2685 95
rect -2570 95 -2520 110
rect -2735 10 -2685 25
rect -2570 25 -2555 95
rect -2535 25 -2520 95
rect -2570 10 -2520 25
rect -2505 95 -2455 110
rect -2505 25 -2490 95
rect -2470 25 -2455 95
rect -2505 10 -2455 25
rect -2340 95 -2290 110
rect -2340 25 -2325 95
rect -2305 25 -2290 95
rect -2340 10 -2290 25
rect -2275 95 -2225 110
rect -2275 25 -2260 95
rect -2240 25 -2225 95
rect -2110 95 -2060 110
rect -2275 10 -2225 25
rect -2110 25 -2095 95
rect -2075 25 -2060 95
rect -2110 10 -2060 25
rect -2045 95 -1995 110
rect -2045 25 -2030 95
rect -2010 25 -1995 95
rect -2045 10 -1995 25
rect -1880 95 -1830 110
rect -1880 25 -1865 95
rect -1845 25 -1830 95
rect -1880 10 -1830 25
rect -1815 95 -1765 110
rect -1815 25 -1800 95
rect -1780 25 -1765 95
rect -1815 10 -1765 25
rect -1480 85 -1430 100
rect -1480 15 -1465 85
rect -1445 15 -1430 85
rect -1480 0 -1430 15
rect -1370 85 -1320 100
rect -1370 15 -1355 85
rect -1335 15 -1320 85
rect -1370 0 -1320 15
rect -1260 85 -1210 100
rect -1260 15 -1245 85
rect -1225 15 -1210 85
rect -1260 0 -1210 15
rect -1150 85 -1100 100
rect -1150 15 -1135 85
rect -1115 15 -1100 85
rect -1150 0 -1100 15
rect -1040 85 -990 100
rect -1040 15 -1025 85
rect -1005 15 -990 85
rect -1040 0 -990 15
rect -820 85 -770 100
rect -820 15 -805 85
rect -785 15 -770 85
rect -820 0 -770 15
rect -710 85 -660 100
rect -710 15 -695 85
rect -675 15 -660 85
rect -710 0 -660 15
rect -600 85 -550 100
rect -600 15 -585 85
rect -565 15 -550 85
rect -600 0 -550 15
rect -490 85 -440 100
rect -490 15 -475 85
rect -455 15 -440 85
rect -490 0 -440 15
rect -380 85 -330 100
rect -380 15 -365 85
rect -345 15 -330 85
rect -380 0 -330 15
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 60 85 110 100
rect 60 15 75 85
rect 95 15 110 85
rect 60 0 110 15
rect 170 85 220 100
rect 170 15 185 85
rect 205 15 220 85
rect 170 0 220 15
rect 280 85 330 100
rect 280 15 295 85
rect 315 15 330 85
rect 280 0 330 15
rect 390 85 440 100
rect 390 15 405 85
rect 425 15 440 85
rect 390 0 440 15
<< pdiff >>
rect -3550 425 -3500 440
rect -3550 255 -3535 425
rect -3515 255 -3500 425
rect -3550 240 -3500 255
rect -3485 425 -3435 440
rect -3485 255 -3470 425
rect -3450 255 -3435 425
rect -3485 240 -3435 255
rect -3400 425 -3350 440
rect -3400 255 -3385 425
rect -3365 255 -3350 425
rect -3400 240 -3350 255
rect -3335 425 -3285 440
rect -3335 255 -3320 425
rect -3300 255 -3285 425
rect -3335 240 -3285 255
rect -3250 425 -3200 440
rect -3250 255 -3235 425
rect -3215 255 -3200 425
rect -3250 240 -3200 255
rect -3185 425 -3135 440
rect -3185 255 -3170 425
rect -3150 255 -3135 425
rect -3185 240 -3135 255
rect -3025 425 -2975 440
rect -3025 255 -3010 425
rect -2990 255 -2975 425
rect -3025 240 -2975 255
rect -2960 425 -2910 440
rect -2960 255 -2945 425
rect -2925 255 -2910 425
rect -2800 425 -2750 440
rect -2960 240 -2910 255
rect -2800 255 -2785 425
rect -2765 255 -2750 425
rect -2800 240 -2750 255
rect -2735 425 -2685 440
rect -2735 255 -2720 425
rect -2700 255 -2685 425
rect -2735 240 -2685 255
rect -2570 425 -2520 440
rect -2570 255 -2555 425
rect -2535 255 -2520 425
rect -2570 240 -2520 255
rect -2505 425 -2455 440
rect -2505 255 -2490 425
rect -2470 255 -2455 425
rect -2340 425 -2290 440
rect -2505 240 -2455 255
rect -2340 255 -2325 425
rect -2305 255 -2290 425
rect -2340 240 -2290 255
rect -2275 425 -2225 440
rect -2275 255 -2260 425
rect -2240 255 -2225 425
rect -2275 240 -2225 255
rect -2110 425 -2060 440
rect -2110 255 -2095 425
rect -2075 255 -2060 425
rect -2110 240 -2060 255
rect -2045 425 -1995 440
rect -2045 255 -2030 425
rect -2010 255 -1995 425
rect -1880 425 -1830 440
rect -2045 240 -1995 255
rect -1880 255 -1865 425
rect -1845 255 -1830 425
rect -1880 240 -1830 255
rect -1815 425 -1765 440
rect -1815 255 -1800 425
rect -1780 255 -1765 425
rect -1815 240 -1765 255
rect -1530 335 -1480 350
rect -1530 265 -1515 335
rect -1495 265 -1480 335
rect -1530 250 -1480 265
rect -1420 335 -1370 350
rect -1420 265 -1405 335
rect -1385 265 -1370 335
rect -1420 250 -1370 265
rect -1310 335 -1260 350
rect -1310 265 -1295 335
rect -1275 265 -1260 335
rect -1310 250 -1260 265
rect -1200 335 -1150 350
rect -1200 265 -1185 335
rect -1165 265 -1150 335
rect -1200 250 -1150 265
rect -1090 335 -1040 350
rect -1090 265 -1075 335
rect -1055 265 -1040 335
rect -1090 250 -1040 265
rect -980 335 -930 350
rect -980 265 -965 335
rect -945 265 -930 335
rect -980 250 -930 265
rect -870 335 -820 350
rect -870 265 -855 335
rect -835 265 -820 335
rect -870 250 -820 265
rect -760 335 -710 350
rect -760 265 -745 335
rect -725 265 -710 335
rect -760 250 -710 265
rect -650 335 -600 350
rect -650 265 -635 335
rect -615 265 -600 335
rect -650 250 -600 265
rect -490 335 -440 350
rect -490 265 -475 335
rect -455 265 -440 335
rect -490 250 -440 265
rect -380 335 -330 350
rect -380 265 -365 335
rect -345 265 -330 335
rect -380 250 -330 265
rect -270 335 -220 350
rect -270 265 -255 335
rect -235 265 -220 335
rect -270 250 -220 265
rect -160 335 -110 350
rect -160 265 -145 335
rect -125 265 -110 335
rect -160 250 -110 265
rect -50 335 0 350
rect -50 265 -35 335
rect -15 265 0 335
rect -50 250 0 265
rect 60 335 110 350
rect 60 265 75 335
rect 95 265 110 335
rect 60 250 110 265
rect 170 335 220 350
rect 170 265 185 335
rect 205 265 220 335
rect 170 250 220 265
rect 280 335 330 350
rect 280 265 295 335
rect 315 265 330 335
rect 280 250 330 265
rect 390 335 440 350
rect 390 265 405 335
rect 425 265 440 335
rect 390 250 440 265
<< ndiffc >>
rect -3535 25 -3515 95
rect -3470 25 -3450 95
rect -3385 25 -3365 95
rect -3320 25 -3300 95
rect -3235 25 -3215 95
rect -3170 25 -3150 95
rect -3010 25 -2990 95
rect -2945 25 -2925 95
rect -2785 25 -2765 95
rect -2720 25 -2700 95
rect -2555 25 -2535 95
rect -2490 25 -2470 95
rect -2325 25 -2305 95
rect -2260 25 -2240 95
rect -2095 25 -2075 95
rect -2030 25 -2010 95
rect -1865 25 -1845 95
rect -1800 25 -1780 95
rect -1465 15 -1445 85
rect -1355 15 -1335 85
rect -1245 15 -1225 85
rect -1135 15 -1115 85
rect -1025 15 -1005 85
rect -805 15 -785 85
rect -695 15 -675 85
rect -585 15 -565 85
rect -475 15 -455 85
rect -365 15 -345 85
rect -35 15 -15 85
rect 75 15 95 85
rect 185 15 205 85
rect 295 15 315 85
rect 405 15 425 85
<< pdiffc >>
rect -3535 255 -3515 425
rect -3470 255 -3450 425
rect -3385 255 -3365 425
rect -3320 255 -3300 425
rect -3235 255 -3215 425
rect -3170 255 -3150 425
rect -3010 255 -2990 425
rect -2945 255 -2925 425
rect -2785 255 -2765 425
rect -2720 255 -2700 425
rect -2555 255 -2535 425
rect -2490 255 -2470 425
rect -2325 255 -2305 425
rect -2260 255 -2240 425
rect -2095 255 -2075 425
rect -2030 255 -2010 425
rect -1865 255 -1845 425
rect -1800 255 -1780 425
rect -1515 265 -1495 335
rect -1405 265 -1385 335
rect -1295 265 -1275 335
rect -1185 265 -1165 335
rect -1075 265 -1055 335
rect -965 265 -945 335
rect -855 265 -835 335
rect -745 265 -725 335
rect -635 265 -615 335
rect -475 265 -455 335
rect -365 265 -345 335
rect -255 265 -235 335
rect -145 265 -125 335
rect -35 265 -15 335
rect 75 265 95 335
rect 185 265 205 335
rect 295 265 315 335
rect 405 265 425 335
<< psubdiff >>
rect -2880 95 -2830 110
rect -2880 25 -2865 95
rect -2845 25 -2830 95
rect -2880 10 -2830 25
rect -2425 95 -2375 110
rect -2425 25 -2410 95
rect -2390 25 -2375 95
rect -2425 10 -2375 25
rect -1965 95 -1915 110
rect -1965 25 -1950 95
rect -1930 25 -1915 95
rect -1965 10 -1915 25
rect -955 85 -905 100
rect -955 15 -940 85
rect -920 15 -905 85
rect -955 0 -905 15
rect -300 85 -250 100
rect -300 15 -285 85
rect -265 15 -250 85
rect -300 0 -250 15
<< nsubdiff >>
rect -3105 425 -3055 440
rect -3105 255 -3090 425
rect -3070 255 -3055 425
rect -3105 240 -3055 255
rect -2650 425 -2600 440
rect -2650 255 -2635 425
rect -2615 255 -2600 425
rect -2650 240 -2600 255
rect -2190 425 -2140 440
rect -2190 255 -2175 425
rect -2155 255 -2140 425
rect -2190 240 -2140 255
rect -570 335 -520 350
rect -570 265 -555 335
rect -535 265 -520 335
rect -570 250 -520 265
<< psubdiffcont >>
rect -2865 25 -2845 95
rect -2410 25 -2390 95
rect -1950 25 -1930 95
rect -940 15 -920 85
rect -285 15 -265 85
<< nsubdiffcont >>
rect -3090 255 -3070 425
rect -2635 255 -2615 425
rect -2175 255 -2155 425
rect -555 265 -535 335
<< poly >>
rect -3160 860 590 875
rect -3160 740 -3145 860
rect -1695 740 -1680 860
rect -3160 730 -3120 740
rect -3160 710 -3150 730
rect -3130 710 -3120 730
rect -3160 700 -3120 710
rect -3020 730 -1680 740
rect -3020 710 -3010 730
rect -2990 725 -1680 730
rect -2990 710 -2980 725
rect -3020 700 -2980 710
rect -2940 690 -1720 700
rect -2940 670 -2930 690
rect -2910 685 -1720 690
rect -2910 670 -2900 685
rect -2940 660 -2900 670
rect -3200 620 -1815 635
rect -3500 440 -3485 455
rect -3350 440 -3335 455
rect -3200 440 -3185 620
rect -3160 585 -3120 595
rect -3160 565 -3150 585
rect -3130 570 -3120 585
rect -3130 565 -2960 570
rect -3160 555 -2960 565
rect -2975 440 -2960 555
rect -2520 455 -2415 470
rect -2750 440 -2735 455
rect -2520 440 -2505 455
rect -2430 445 -2415 455
rect -2885 430 -2845 440
rect -2885 410 -2875 430
rect -2855 410 -2845 430
rect -2885 400 -2845 410
rect -2430 435 -2390 445
rect -2290 440 -2275 455
rect -2060 440 -2045 455
rect -1830 440 -1815 620
rect -2430 415 -2420 435
rect -2400 415 -2390 435
rect -2430 405 -2390 415
rect -1970 425 -1930 435
rect -1970 405 -1960 425
rect -1940 405 -1930 425
rect -1970 395 -1930 405
rect -3500 185 -3485 240
rect -3350 200 -3335 240
rect -3200 200 -3185 240
rect -2975 225 -2960 240
rect -3565 170 -3485 185
rect -3500 110 -3485 170
rect -3375 190 -3335 200
rect -3375 170 -3365 190
rect -3345 170 -3335 190
rect -3375 160 -3335 170
rect -3225 190 -3185 200
rect -3225 170 -3215 190
rect -3195 170 -3185 190
rect -3225 160 -3185 170
rect -3020 190 -2980 200
rect -3020 170 -3010 190
rect -2990 170 -2980 190
rect -3020 160 -2980 170
rect -2955 190 -2915 200
rect -2955 170 -2945 190
rect -2925 170 -2915 190
rect -2955 160 -2915 170
rect -3350 110 -3335 160
rect -3200 135 -3185 160
rect -3200 120 -2960 135
rect -3200 110 -3185 120
rect -2975 110 -2960 120
rect -2750 110 -2735 240
rect -2520 225 -2505 240
rect -2290 215 -2275 240
rect -2060 215 -2045 240
rect -1830 225 -1815 240
rect -2290 200 -1850 215
rect -2710 190 -2670 200
rect -2710 170 -2700 190
rect -2680 185 -2670 190
rect -2565 190 -2525 200
rect -2565 185 -2555 190
rect -2680 170 -2555 185
rect -2535 170 -2525 190
rect -2710 160 -2670 170
rect -2565 160 -2525 170
rect -2500 190 -2460 200
rect -2500 170 -2490 190
rect -2470 185 -2460 190
rect -2315 190 -2275 200
rect -2315 185 -2305 190
rect -2470 170 -2305 185
rect -2285 170 -2275 190
rect -2500 160 -2460 170
rect -2315 160 -2275 170
rect -2520 110 -2505 125
rect -2290 110 -2275 160
rect -1865 135 -1850 200
rect -1735 200 -1720 685
rect -1480 350 -1420 365
rect -1370 350 -1310 365
rect -1260 350 -1200 365
rect -1150 350 -1090 365
rect -1040 350 -980 365
rect -930 350 -870 365
rect -820 350 -760 365
rect -710 350 -650 365
rect -440 350 -380 365
rect -330 350 -270 365
rect -220 350 -160 365
rect -110 350 -50 365
rect 0 350 60 365
rect 110 350 170 365
rect 220 350 280 365
rect 330 350 390 365
rect -1480 240 -1420 250
rect -1370 240 -1310 250
rect -1260 240 -1200 250
rect -1150 240 -1090 250
rect -1040 240 -980 250
rect -930 240 -870 250
rect -820 240 -760 250
rect -710 240 -650 250
rect -1480 225 -650 240
rect -440 240 -380 250
rect -330 240 -270 250
rect -220 240 -160 250
rect -110 240 -50 250
rect 0 240 60 250
rect 110 240 170 250
rect 220 240 280 250
rect 330 240 390 250
rect 590 240 605 250
rect -440 225 605 240
rect -440 200 -425 225
rect -1735 185 -425 200
rect -1475 145 -1435 155
rect -1475 135 -1465 145
rect -2060 110 -2045 125
rect -1865 120 -1815 135
rect -1830 110 -1815 120
rect -1680 125 -1465 135
rect -1445 135 -1435 145
rect -1255 145 -1215 155
rect -1255 135 -1245 145
rect -1445 125 -1245 135
rect -1225 135 -1215 145
rect -1035 145 -995 155
rect -1035 135 -1025 145
rect -1225 125 -1025 135
rect -1005 135 -995 145
rect -1005 125 -380 135
rect -1680 110 -380 125
rect -3090 40 -3050 50
rect -3090 20 -3080 40
rect -3060 20 -3050 40
rect -3090 10 -3050 20
rect -2635 40 -2595 50
rect -2635 20 -2625 40
rect -2605 20 -2595 40
rect -2635 10 -2595 20
rect -2175 40 -2135 50
rect -2175 20 -2165 40
rect -2145 20 -2135 40
rect -2175 10 -2135 20
rect -3500 -5 -3485 10
rect -3350 -5 -3335 10
rect -3200 -5 -3185 10
rect -2975 -5 -2960 10
rect -2750 -120 -2735 10
rect -2610 0 -2595 10
rect -2520 0 -2505 10
rect -2610 -15 -2505 0
rect -2290 -5 -2275 10
rect -2250 -15 -2210 -10
rect -2060 -15 -2045 10
rect -1830 -5 -1815 10
rect -3565 -135 -2735 -120
rect -2250 -20 -2045 -15
rect -2250 -40 -2240 -20
rect -2220 -30 -2045 -20
rect -2020 -15 -1980 -5
rect -2220 -40 -2210 -30
rect -2250 -50 -2210 -40
rect -2020 -35 -2010 -15
rect -1990 -30 -1980 -15
rect -1680 -30 -1665 110
rect -1430 100 -1370 110
rect -1320 100 -1260 110
rect -1210 100 -1150 110
rect -1100 100 -1040 110
rect -770 100 -710 110
rect -660 100 -600 110
rect -550 100 -490 110
rect -440 100 -380 110
rect 0 110 605 125
rect 0 100 60 110
rect 110 100 170 110
rect 220 100 280 110
rect 330 100 390 110
rect 590 100 605 110
rect -1430 -15 -1370 0
rect -1320 -15 -1260 0
rect -1210 -15 -1150 0
rect -1100 -15 -1040 0
rect -770 -15 -710 0
rect -660 -15 -600 0
rect -550 -15 -490 0
rect -440 -15 -380 0
rect 0 -15 60 0
rect 110 -15 170 0
rect 220 -15 280 0
rect 330 -15 390 0
rect -1990 -35 -1665 -30
rect -2020 -45 -1665 -35
rect -2250 -160 -2235 -50
rect -2105 -105 -2065 -95
rect -2105 -125 -2095 -105
rect -2075 -120 -2065 -105
rect -1885 -105 -1845 -95
rect -1885 -120 -1875 -105
rect -2075 -125 -1875 -120
rect -1855 -120 -1845 -105
rect -1855 -125 -1640 -120
rect -2105 -135 -1640 -125
rect -1655 -160 -1640 -135
rect -2250 -175 590 -160
<< polycont >>
rect -3150 710 -3130 730
rect -3010 710 -2990 730
rect -2930 670 -2910 690
rect -3150 565 -3130 585
rect -2875 410 -2855 430
rect -2420 415 -2400 435
rect -1960 405 -1940 425
rect -3365 170 -3345 190
rect -3215 170 -3195 190
rect -3010 170 -2990 190
rect -2945 170 -2925 190
rect -2700 170 -2680 190
rect -2555 170 -2535 190
rect -2490 170 -2470 190
rect -2305 170 -2285 190
rect -1465 125 -1445 145
rect -1245 125 -1225 145
rect -1025 125 -1005 145
rect -3080 20 -3060 40
rect -2625 20 -2605 40
rect -2165 20 -2145 40
rect -2240 -40 -2220 -20
rect -2010 -35 -1990 -15
rect -2095 -125 -2075 -105
rect -1875 -125 -1855 -105
<< locali >>
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect -3310 760 -1855 780
rect -3310 435 -3290 760
rect -3160 730 -3120 740
rect -3160 710 -3150 730
rect -3130 710 -3120 730
rect -3160 700 -3120 710
rect -3020 730 -2980 740
rect -3020 710 -3010 730
rect -2990 710 -2980 730
rect -3020 700 -2980 710
rect -3160 595 -3140 700
rect -3160 585 -3120 595
rect -3160 565 -3150 585
rect -3130 565 -3120 585
rect -3160 555 -3120 565
rect -3160 435 -3140 555
rect -3020 435 -3000 700
rect -2940 690 -2900 700
rect -2940 670 -2930 690
rect -2910 670 -2900 690
rect -2940 660 -2900 670
rect -2940 435 -2920 660
rect -3545 425 -3505 435
rect -3545 255 -3535 425
rect -3515 255 -3505 425
rect -3545 245 -3505 255
rect -3480 425 -3440 435
rect -3480 255 -3470 425
rect -3450 255 -3440 425
rect -3480 245 -3440 255
rect -3395 425 -3355 435
rect -3395 255 -3385 425
rect -3365 255 -3355 425
rect -3395 245 -3355 255
rect -3330 425 -3290 435
rect -3330 255 -3320 425
rect -3300 255 -3290 425
rect -3330 245 -3290 255
rect -3245 425 -3205 435
rect -3245 255 -3235 425
rect -3215 255 -3205 425
rect -3245 245 -3205 255
rect -3180 425 -3140 435
rect -3180 255 -3170 425
rect -3150 255 -3140 425
rect -3180 245 -3140 255
rect -3100 425 -3060 435
rect -3100 255 -3090 425
rect -3070 255 -3060 425
rect -3100 245 -3060 255
rect -3020 425 -2980 435
rect -3020 255 -3010 425
rect -2990 255 -2980 425
rect -3020 245 -2980 255
rect -2955 425 -2915 435
rect -2955 255 -2945 425
rect -2925 255 -2915 425
rect -2885 430 -2845 440
rect -2430 435 -2390 445
rect -1875 435 -1855 760
rect -2885 410 -2875 430
rect -2855 410 -2845 430
rect -2885 400 -2845 410
rect -2955 245 -2915 255
rect -3460 190 -3440 245
rect -3375 190 -3335 200
rect -3460 170 -3365 190
rect -3345 170 -3335 190
rect -3460 105 -3440 170
rect -3375 160 -3335 170
rect -3310 190 -3290 245
rect -3225 190 -3185 200
rect -3310 170 -3215 190
rect -3195 170 -3185 190
rect -3310 105 -3290 170
rect -3225 160 -3185 170
rect -3160 105 -3140 245
rect -3545 95 -3505 105
rect -3545 25 -3535 95
rect -3515 25 -3505 95
rect -3545 15 -3505 25
rect -3480 95 -3440 105
rect -3480 25 -3470 95
rect -3450 25 -3440 95
rect -3480 15 -3440 25
rect -3395 95 -3355 105
rect -3395 25 -3385 95
rect -3365 25 -3355 95
rect -3395 15 -3355 25
rect -3330 95 -3290 105
rect -3330 25 -3320 95
rect -3300 25 -3290 95
rect -3330 15 -3290 25
rect -3245 95 -3205 105
rect -3245 25 -3235 95
rect -3215 25 -3205 95
rect -3245 15 -3205 25
rect -3180 95 -3140 105
rect -3180 25 -3170 95
rect -3150 25 -3140 95
rect -3180 15 -3140 25
rect -3090 50 -3070 245
rect -3010 200 -2990 245
rect -2945 200 -2925 245
rect -3020 190 -2980 200
rect -3020 170 -3010 190
rect -2990 170 -2980 190
rect -3020 160 -2980 170
rect -2955 190 -2915 200
rect -2955 170 -2945 190
rect -2925 170 -2915 190
rect -2955 160 -2915 170
rect -3010 105 -2990 160
rect -2945 105 -2925 160
rect -2865 105 -2845 400
rect -2795 425 -2755 435
rect -2795 255 -2785 425
rect -2765 255 -2755 425
rect -2795 245 -2755 255
rect -2730 425 -2690 435
rect -2730 255 -2720 425
rect -2700 255 -2690 425
rect -2730 245 -2690 255
rect -2645 425 -2605 435
rect -2645 255 -2635 425
rect -2615 255 -2605 425
rect -2645 245 -2605 255
rect -2565 425 -2525 435
rect -2565 255 -2555 425
rect -2535 255 -2525 425
rect -2565 245 -2525 255
rect -2500 425 -2460 435
rect -2500 255 -2490 425
rect -2470 255 -2460 425
rect -2430 415 -2420 435
rect -2400 415 -2390 435
rect -2430 405 -2390 415
rect -2500 245 -2460 255
rect -2710 200 -2690 245
rect -2710 190 -2670 200
rect -2710 170 -2700 190
rect -2680 170 -2670 190
rect -2710 160 -2670 170
rect -2710 105 -2690 160
rect -3020 95 -2980 105
rect -3090 40 -3050 50
rect -3090 20 -3080 40
rect -3060 20 -3050 40
rect -3090 10 -3050 20
rect -3020 25 -3010 95
rect -2990 25 -2980 95
rect -3020 15 -2980 25
rect -2955 95 -2915 105
rect -2955 25 -2945 95
rect -2925 25 -2915 95
rect -2955 15 -2915 25
rect -2875 95 -2835 105
rect -2875 25 -2865 95
rect -2845 25 -2835 95
rect -2875 15 -2835 25
rect -2795 95 -2755 105
rect -2795 25 -2785 95
rect -2765 25 -2755 95
rect -2795 15 -2755 25
rect -2730 95 -2690 105
rect -2730 25 -2720 95
rect -2700 25 -2690 95
rect -2730 15 -2690 25
rect -2635 50 -2615 245
rect -2555 200 -2535 245
rect -2490 200 -2470 245
rect -2565 190 -2525 200
rect -2565 170 -2555 190
rect -2535 170 -2525 190
rect -2565 160 -2525 170
rect -2500 190 -2460 200
rect -2500 170 -2490 190
rect -2470 170 -2460 190
rect -2500 160 -2460 170
rect -2555 105 -2535 160
rect -2490 105 -2470 160
rect -2410 105 -2390 405
rect -2335 425 -2295 435
rect -2335 255 -2325 425
rect -2305 255 -2295 425
rect -2335 245 -2295 255
rect -2270 425 -2230 435
rect -2270 255 -2260 425
rect -2240 255 -2230 425
rect -2270 245 -2230 255
rect -2185 425 -2145 435
rect -2185 255 -2175 425
rect -2155 255 -2145 425
rect -2185 245 -2145 255
rect -2105 425 -2065 435
rect -2105 255 -2095 425
rect -2075 255 -2065 425
rect -2105 245 -2065 255
rect -2040 425 -2000 435
rect -2040 255 -2030 425
rect -2010 255 -2000 425
rect -1970 425 -1930 435
rect -1970 405 -1960 425
rect -1940 405 -1930 425
rect -1970 395 -1930 405
rect -2040 245 -2000 255
rect -2315 190 -2275 200
rect -2315 170 -2305 190
rect -2285 170 -2275 190
rect -2315 160 -2275 170
rect -2250 105 -2230 245
rect -2565 95 -2525 105
rect -2635 40 -2595 50
rect -2635 20 -2625 40
rect -2605 20 -2595 40
rect -2635 10 -2595 20
rect -2565 25 -2555 95
rect -2535 25 -2525 95
rect -2565 15 -2525 25
rect -2500 95 -2460 105
rect -2500 25 -2490 95
rect -2470 25 -2460 95
rect -2500 15 -2460 25
rect -2420 95 -2380 105
rect -2420 25 -2410 95
rect -2390 25 -2380 95
rect -2420 15 -2380 25
rect -2335 95 -2295 105
rect -2335 25 -2325 95
rect -2305 25 -2295 95
rect -2335 15 -2295 25
rect -2270 95 -2230 105
rect -2270 25 -2260 95
rect -2240 25 -2230 95
rect -2270 15 -2230 25
rect -2250 -10 -2230 15
rect -2175 50 -2155 245
rect -2095 105 -2075 245
rect -2030 105 -2010 245
rect -1950 105 -1930 395
rect -1875 425 -1835 435
rect -1875 255 -1865 425
rect -1845 255 -1835 425
rect -1875 245 -1835 255
rect -1810 425 -1770 435
rect -1810 255 -1800 425
rect -1780 255 -1770 425
rect -1515 365 -615 385
rect -1515 345 -1495 365
rect -1295 345 -1275 365
rect -1075 345 -1055 365
rect -855 345 -835 365
rect -635 345 -615 365
rect -475 365 425 385
rect -475 345 -455 365
rect -255 345 -235 365
rect -35 345 -15 365
rect 185 345 205 365
rect 405 345 425 365
rect -1525 335 -1485 345
rect -1525 265 -1515 335
rect -1495 265 -1485 335
rect -1525 255 -1485 265
rect -1415 335 -1375 345
rect -1415 265 -1405 335
rect -1385 265 -1375 335
rect -1415 255 -1375 265
rect -1305 335 -1265 345
rect -1305 265 -1295 335
rect -1275 265 -1265 335
rect -1305 255 -1265 265
rect -1195 335 -1155 345
rect -1195 265 -1185 335
rect -1165 265 -1155 335
rect -1195 255 -1155 265
rect -1085 335 -1045 345
rect -1085 265 -1075 335
rect -1055 265 -1045 335
rect -1085 255 -1045 265
rect -975 335 -935 345
rect -975 265 -965 335
rect -945 265 -935 335
rect -975 255 -935 265
rect -865 335 -825 345
rect -865 265 -855 335
rect -835 265 -825 335
rect -865 255 -825 265
rect -755 335 -715 345
rect -755 265 -745 335
rect -725 265 -715 335
rect -755 255 -715 265
rect -645 335 -605 345
rect -645 265 -635 335
rect -615 265 -605 335
rect -645 255 -605 265
rect -565 335 -525 345
rect -565 265 -555 335
rect -535 265 -525 335
rect -565 255 -525 265
rect -485 335 -445 345
rect -485 265 -475 335
rect -455 265 -445 335
rect -485 255 -445 265
rect -375 335 -335 345
rect -375 265 -365 335
rect -345 265 -335 335
rect -375 255 -335 265
rect -265 335 -225 345
rect -265 265 -255 335
rect -235 265 -225 335
rect -265 255 -225 265
rect -155 335 -115 345
rect -155 265 -145 335
rect -125 265 -115 335
rect -155 255 -115 265
rect -45 335 -5 345
rect -45 265 -35 335
rect -15 265 -5 335
rect -45 255 -5 265
rect 65 335 105 345
rect 65 265 75 335
rect 95 265 105 335
rect 65 255 105 265
rect 175 335 215 345
rect 175 265 185 335
rect 205 265 215 335
rect 175 255 215 265
rect 285 335 325 345
rect 285 265 295 335
rect 315 265 325 335
rect 285 255 325 265
rect 395 335 435 345
rect 395 265 405 335
rect 425 265 435 335
rect 395 255 435 265
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect -1810 245 -1770 255
rect -635 220 -615 255
rect -635 200 -565 220
rect -1475 145 -1435 155
rect -1475 125 -1465 145
rect -1445 125 -1435 145
rect -1475 115 -1435 125
rect -1255 145 -1215 155
rect -1255 125 -1245 145
rect -1225 125 -1215 145
rect -1255 115 -1215 125
rect -1035 145 -995 155
rect -1035 125 -1025 145
rect -1005 125 -995 145
rect -1035 115 -995 125
rect -2105 95 -2065 105
rect -2175 40 -2135 50
rect -2175 20 -2165 40
rect -2145 20 -2135 40
rect -2175 10 -2135 20
rect -2105 25 -2095 95
rect -2075 25 -2065 95
rect -2105 15 -2065 25
rect -2040 95 -1995 105
rect -2040 25 -2030 95
rect -2010 25 -1995 95
rect -2040 15 -1995 25
rect -1965 95 -1920 105
rect -1965 25 -1950 95
rect -1930 25 -1920 95
rect -1965 15 -1920 25
rect -1875 95 -1835 105
rect -1875 25 -1865 95
rect -1845 25 -1835 95
rect -1875 15 -1835 25
rect -1810 95 -1770 105
rect -1465 95 -1445 115
rect -1245 95 -1225 115
rect -1025 95 -1005 115
rect -585 95 -565 200
rect 405 185 425 255
rect 590 250 645 260
rect 405 165 1325 185
rect 405 95 425 165
rect -1810 25 -1800 95
rect -1780 25 -1770 95
rect -1810 15 -1770 25
rect -1475 85 -1435 95
rect -1475 15 -1465 85
rect -1445 15 -1435 85
rect -2250 -20 -2210 -10
rect -2250 -40 -2240 -20
rect -2220 -40 -2210 -20
rect -2250 -50 -2210 -40
rect -2095 -95 -2075 15
rect -2020 -5 -2000 15
rect -2020 -15 -1980 -5
rect -2020 -35 -2010 -15
rect -1990 -35 -1980 -15
rect -2020 -45 -1980 -35
rect -1865 -95 -1845 15
rect -1475 5 -1435 15
rect -1365 85 -1325 95
rect -1365 15 -1355 85
rect -1335 15 -1325 85
rect -1365 5 -1325 15
rect -1255 85 -1215 95
rect -1255 15 -1245 85
rect -1225 15 -1215 85
rect -1255 5 -1215 15
rect -1145 85 -1105 95
rect -1145 15 -1135 85
rect -1115 15 -1105 85
rect -1145 5 -1105 15
rect -1035 85 -995 95
rect -1035 15 -1025 85
rect -1005 15 -995 85
rect -1035 5 -995 15
rect -950 85 -910 95
rect -950 15 -940 85
rect -920 15 -910 85
rect -950 5 -910 15
rect -815 85 -775 95
rect -815 15 -805 85
rect -785 15 -775 85
rect -815 5 -775 15
rect -705 85 -665 95
rect -705 15 -695 85
rect -675 15 -665 85
rect -705 5 -665 15
rect -595 85 -555 95
rect -595 15 -585 85
rect -565 15 -555 85
rect -595 5 -555 15
rect -485 85 -445 95
rect -485 15 -475 85
rect -455 15 -445 85
rect -485 5 -445 15
rect -375 85 -335 95
rect -375 15 -365 85
rect -345 15 -335 85
rect -375 5 -335 15
rect -295 85 -255 95
rect -295 15 -285 85
rect -265 15 -255 85
rect -295 5 -255 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 65 85 105 95
rect 65 15 75 85
rect 95 15 105 85
rect 65 5 105 15
rect 175 85 215 95
rect 175 15 185 85
rect 205 15 215 85
rect 175 5 215 15
rect 285 85 325 95
rect 285 15 295 85
rect 315 15 325 85
rect 285 5 325 15
rect 395 85 435 95
rect 395 15 405 85
rect 425 15 435 85
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 395 5 435 15
rect -1465 -15 -1445 5
rect -1245 -15 -1225 5
rect -1025 -15 -1005 5
rect -2105 -105 -2065 -95
rect -2105 -125 -2095 -105
rect -2075 -125 -2065 -105
rect -2105 -135 -2065 -125
rect -1885 -105 -1845 -95
rect -1885 -125 -1875 -105
rect -1855 -125 -1845 -105
rect -1885 -135 -1845 -125
rect -1630 -35 -1005 -15
rect -805 -15 -785 5
rect -585 -15 -565 5
rect -365 -15 -345 5
rect -805 -35 -345 -15
rect -35 -15 -15 5
rect 185 -15 205 5
rect 405 -15 425 5
rect -35 -35 425 -15
rect -1630 -210 -1610 -35
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
rect -3565 -230 -1610 -210
<< viali >>
rect 600 855 635 890
rect -3535 255 -3515 425
rect -3385 255 -3365 425
rect -3235 255 -3215 425
rect -2875 410 -2855 430
rect -3535 25 -3515 95
rect -3385 25 -3365 95
rect -3235 25 -3215 95
rect -2785 255 -2765 425
rect -2420 415 -2400 435
rect -3080 20 -3060 40
rect -2785 25 -2765 95
rect -2325 255 -2305 425
rect -1960 405 -1940 425
rect -2625 20 -2605 40
rect -2325 25 -2305 95
rect -1800 255 -1780 425
rect -1405 265 -1385 335
rect -1185 265 -1165 335
rect -965 265 -945 335
rect -745 265 -725 335
rect -555 265 -535 335
rect -365 265 -345 335
rect -145 265 -125 335
rect 75 265 95 335
rect 295 265 315 335
rect 600 260 635 295
rect -2165 20 -2145 40
rect -1800 25 -1780 95
rect -1355 15 -1335 85
rect -1135 15 -1115 85
rect -940 15 -920 85
rect -695 15 -675 85
rect -475 15 -455 85
rect -285 15 -265 85
rect 75 15 95 85
rect 295 15 315 85
rect 600 55 635 90
rect 600 -165 635 -130
<< metal1 >>
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect -3600 435 440 440
rect -3600 430 -2420 435
rect -3600 425 -2875 430
rect -3600 255 -3535 425
rect -3515 255 -3385 425
rect -3365 255 -3235 425
rect -3215 410 -2875 425
rect -2855 425 -2420 430
rect -2855 410 -2785 425
rect -3215 255 -2785 410
rect -2765 415 -2420 425
rect -2400 425 440 435
rect -2400 415 -2325 425
rect -2765 255 -2325 415
rect -2305 405 -1960 425
rect -1940 405 -1800 425
rect -2305 255 -1800 405
rect -1780 335 440 425
rect -1780 265 -1405 335
rect -1385 265 -1185 335
rect -1165 265 -965 335
rect -945 265 -745 335
rect -725 265 -555 335
rect -535 265 -365 335
rect -345 265 -145 335
rect -125 265 75 335
rect 95 265 295 335
rect 315 265 440 335
rect -1780 255 440 265
rect -3600 240 440 255
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect -3600 95 440 110
rect -3600 25 -3535 95
rect -3515 25 -3385 95
rect -3365 25 -3235 95
rect -3215 40 -2785 95
rect -3215 25 -3080 40
rect -3600 20 -3080 25
rect -3060 25 -2785 40
rect -2765 40 -2325 95
rect -2765 25 -2625 40
rect -3060 20 -2625 25
rect -2605 25 -2325 40
rect -2305 40 -1800 95
rect -2305 25 -2165 40
rect -2605 20 -2165 25
rect -2145 25 -1800 40
rect -1780 85 440 95
rect -1780 25 -1355 85
rect -2145 20 -1355 25
rect -3600 15 -1355 20
rect -1335 15 -1135 85
rect -1115 15 -940 85
rect -920 15 -695 85
rect -675 15 -475 85
rect -455 15 -285 85
rect -265 15 75 85
rect 95 15 295 85
rect 315 15 440 85
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect -3600 0 440 15
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
<< via1 >>
rect 600 855 635 890
rect 600 260 635 295
rect 600 55 635 90
rect 600 -165 635 -130
<< metal2 >>
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
<< via2 >>
rect 600 855 635 890
rect 600 260 635 295
rect 600 55 635 90
rect 600 -165 635 -130
<< metal3 >>
rect 765 900 1215 925
rect 590 890 1215 900
rect 590 855 600 890
rect 635 855 1215 890
rect 590 845 1215 855
rect 765 305 1215 845
rect 590 295 1215 305
rect 590 260 600 295
rect 635 260 1215 295
rect 590 250 1215 260
rect 765 235 1215 250
rect 765 100 1055 115
rect 590 90 1055 100
rect 590 55 600 90
rect 635 55 1055 90
rect 590 45 1055 55
rect 765 -120 1055 45
rect 590 -130 1055 -120
rect 590 -165 600 -130
rect 635 -165 1055 -130
rect 590 -175 1055 -165
<< via3 >>
rect 600 260 635 295
rect 600 55 635 90
<< mimcap >>
rect 780 295 1200 910
rect 780 260 790 295
rect 825 260 1200 295
rect 780 250 1200 260
rect 780 90 1040 100
rect 780 55 790 90
rect 825 55 1040 90
rect 780 -160 1040 55
<< mimcapcontact >>
rect 790 260 825 295
rect 790 55 825 90
<< metal4 >>
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect 780 295 835 305
rect 780 260 790 295
rect 825 260 835 295
rect 780 250 835 260
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 780 90 835 100
rect 780 55 790 90
rect 825 55 835 90
rect 780 45 835 55
<< labels >>
flabel locali 1325 175 1325 175 3 FreeSans 400 0 80 0 VOUT
flabel locali -3565 -220 -3565 -220 7 FreeSans 400 0 -200 0 I_IN
flabel poly -3565 -125 -3565 -125 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel poly -3565 175 -3565 175 7 FreeSans 400 0 -200 0 UP_PFD
flabel metal1 -3600 340 -3600 340 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 -3600 60 -3600 60 7 FreeSans 400 0 -200 0 GNDA
<< end >>
