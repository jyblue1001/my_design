magic
tech sky130A
timestamp 1750039422
<< nwell >>
rect 31150 4635 31940 4950
rect 32120 4635 32790 4925
rect 31180 4225 32570 4505
rect 31130 3810 32715 4095
rect 29885 2950 30725 3780
rect 31150 3090 32650 3670
rect 29885 2390 30725 2820
rect 30935 2380 31835 2960
rect 31965 2380 32865 2960
rect 33075 2950 33915 3780
rect 33075 2390 33915 2820
<< pwell >>
rect 29480 3700 29770 3705
rect 29480 3680 29585 3700
rect 29665 3680 29770 3700
rect 29480 2970 29770 3680
rect 29395 1900 29760 2674
rect 34030 3700 34320 3705
rect 34030 3680 34135 3700
rect 34215 3680 34320 3700
rect 34030 2970 34320 3680
rect 29900 1845 30710 2345
rect 31090 1930 32710 2280
rect 31890 1925 31910 1930
rect 33090 1845 33900 2345
rect 34040 1900 34405 2674
rect 29650 833 29905 1720
rect 29980 855 30730 1765
rect 30935 1460 32865 1810
rect 31135 835 32585 1320
rect 33070 845 33820 1765
rect 33425 840 33465 845
rect 33900 833 34150 1720
rect 31200 530 31595 795
rect 31810 535 32640 795
<< nmos >>
rect 29995 1945 30010 2245
rect 30050 1945 30065 2245
rect 30105 1945 30120 2245
rect 30160 1945 30175 2245
rect 30215 1945 30230 2245
rect 30270 1945 30285 2245
rect 30325 1945 30340 2245
rect 30380 1945 30395 2245
rect 30435 1945 30450 2245
rect 30490 1945 30505 2245
rect 30545 1945 30560 2245
rect 30600 1945 30615 2245
rect 31225 2030 31240 2180
rect 31280 2030 31295 2180
rect 31335 2030 31350 2180
rect 31390 2030 31405 2180
rect 31445 2030 31460 2180
rect 31500 2030 31515 2180
rect 31555 2030 31570 2180
rect 31610 2030 31625 2180
rect 31665 2030 31680 2180
rect 31720 2030 31735 2180
rect 31775 2030 31790 2180
rect 31830 2030 31845 2180
rect 31955 2030 31970 2180
rect 32010 2030 32025 2180
rect 32065 2030 32080 2180
rect 32120 2030 32135 2180
rect 32175 2030 32190 2180
rect 32230 2030 32245 2180
rect 32285 2030 32300 2180
rect 32340 2030 32355 2180
rect 32395 2030 32410 2180
rect 32450 2030 32465 2180
rect 32505 2030 32520 2180
rect 32560 2030 32575 2180
rect 33185 1945 33200 2245
rect 33240 1945 33255 2245
rect 33295 1945 33310 2245
rect 33350 1945 33365 2245
rect 33405 1945 33420 2245
rect 33460 1945 33475 2245
rect 33515 1945 33530 2245
rect 33570 1945 33585 2245
rect 33625 1945 33640 2245
rect 33680 1945 33695 2245
rect 33735 1945 33750 2245
rect 33790 1945 33805 2245
rect 30075 955 30135 1655
rect 30175 955 30235 1655
rect 30275 955 30335 1655
rect 30375 955 30435 1655
rect 30475 955 30535 1655
rect 30575 955 30635 1655
rect 31070 1560 31085 1710
rect 31125 1560 31140 1710
rect 31180 1560 31195 1710
rect 31235 1560 31250 1710
rect 31290 1560 31305 1710
rect 31345 1560 31360 1710
rect 31400 1560 31415 1710
rect 31455 1560 31470 1710
rect 31510 1560 31525 1710
rect 31565 1560 31580 1710
rect 31620 1560 31635 1710
rect 31675 1560 31690 1710
rect 31810 1560 31825 1710
rect 31865 1560 31880 1710
rect 31920 1560 31935 1710
rect 31975 1560 31990 1710
rect 32110 1560 32125 1710
rect 32165 1560 32180 1710
rect 32220 1560 32235 1710
rect 32275 1560 32290 1710
rect 32330 1560 32345 1710
rect 32385 1560 32400 1710
rect 32440 1560 32455 1710
rect 32495 1560 32510 1710
rect 32550 1560 32565 1710
rect 32605 1560 32620 1710
rect 32660 1560 32675 1710
rect 32715 1560 32730 1710
rect 31245 955 31260 1205
rect 31300 955 31315 1205
rect 31355 955 31370 1205
rect 31410 955 31425 1205
rect 31465 955 31480 1205
rect 31520 955 31535 1205
rect 31575 955 31590 1205
rect 31630 955 31645 1205
rect 31685 955 31700 1205
rect 31740 955 31755 1205
rect 31795 955 31810 1205
rect 31850 955 31865 1205
rect 31905 955 31920 1205
rect 31960 955 31975 1205
rect 32015 955 32030 1205
rect 32070 955 32085 1205
rect 32125 955 32140 1205
rect 32180 955 32195 1205
rect 32235 955 32250 1205
rect 32290 955 32305 1205
rect 32345 955 32360 1205
rect 32400 955 32415 1205
rect 32455 955 32470 1205
rect 33165 955 33225 1655
rect 33265 955 33325 1655
rect 33365 955 33425 1655
rect 33465 955 33525 1655
rect 33565 955 33625 1655
rect 33665 955 33725 1655
rect 31300 590 31490 690
rect 31920 635 31935 685
rect 31975 635 31990 685
rect 32030 635 32045 685
rect 32085 635 32100 685
rect 32140 635 32155 685
rect 32195 635 32210 685
rect 32250 635 32265 685
rect 32305 635 32320 685
rect 32360 635 32375 685
rect 32415 635 32430 685
rect 32470 635 32485 685
rect 32525 635 32540 685
<< pmos >>
rect 31260 4755 31280 4818
rect 31320 4755 31340 4818
rect 31380 4755 31400 4818
rect 31510 4755 31530 4835
rect 31570 4755 31590 4835
rect 31630 4755 31650 4835
rect 31690 4755 31710 4835
rect 31750 4755 31770 4835
rect 31810 4755 31830 4835
rect 32240 4750 32260 4810
rect 32300 4750 32320 4810
rect 32360 4750 32380 4810
rect 32420 4750 32440 4810
rect 32480 4750 32500 4810
rect 32540 4750 32560 4810
rect 32600 4750 32620 4810
rect 32660 4750 32680 4810
rect 31290 4340 31305 4390
rect 31345 4340 31360 4390
rect 31400 4340 31415 4390
rect 31455 4340 31470 4390
rect 31510 4340 31525 4390
rect 31565 4340 31580 4390
rect 31620 4340 31635 4390
rect 31675 4340 31690 4390
rect 31730 4340 31745 4390
rect 31785 4340 31800 4390
rect 31840 4340 31855 4390
rect 31895 4340 31910 4390
rect 31950 4340 31965 4390
rect 32005 4340 32020 4390
rect 32060 4340 32075 4390
rect 32115 4340 32130 4390
rect 32170 4340 32185 4390
rect 32225 4340 32240 4390
rect 32280 4340 32295 4390
rect 32335 4340 32350 4390
rect 32390 4340 32405 4390
rect 32445 4340 32460 4390
rect 31240 3930 31255 3980
rect 31295 3930 31310 3980
rect 31350 3930 31365 3980
rect 31405 3930 31420 3980
rect 31460 3930 31475 3980
rect 31515 3930 31530 3980
rect 31570 3930 31585 3980
rect 31625 3930 31640 3980
rect 31680 3930 31695 3980
rect 31735 3930 31750 3980
rect 31790 3930 31805 3980
rect 31845 3930 31860 3980
rect 31970 3930 31985 3980
rect 32025 3930 32040 3980
rect 32080 3930 32095 3980
rect 32135 3930 32150 3980
rect 32190 3930 32205 3980
rect 32245 3930 32260 3980
rect 32300 3930 32315 3980
rect 32355 3930 32370 3980
rect 32410 3930 32425 3980
rect 32465 3930 32480 3980
rect 32520 3930 32535 3980
rect 32575 3930 32590 3980
rect 29995 3065 30010 3665
rect 30050 3065 30065 3665
rect 30105 3065 30120 3665
rect 30160 3065 30175 3665
rect 30215 3065 30230 3665
rect 30270 3065 30285 3665
rect 30325 3065 30340 3665
rect 30380 3065 30395 3665
rect 30435 3065 30450 3665
rect 30490 3065 30505 3665
rect 30545 3065 30560 3665
rect 30600 3065 30615 3665
rect 31260 3205 31280 3555
rect 31320 3205 31340 3555
rect 31380 3205 31400 3555
rect 31440 3205 31460 3555
rect 31500 3205 31520 3555
rect 31560 3205 31580 3555
rect 31620 3205 31640 3555
rect 31680 3205 31700 3555
rect 31740 3205 31760 3555
rect 31800 3205 31820 3555
rect 31860 3205 31880 3555
rect 31920 3205 31940 3555
rect 31980 3205 32000 3555
rect 32040 3205 32060 3555
rect 32100 3205 32120 3555
rect 32160 3205 32180 3555
rect 32220 3205 32240 3555
rect 32280 3205 32300 3555
rect 32340 3205 32360 3555
rect 32400 3205 32420 3555
rect 32460 3205 32480 3555
rect 32520 3205 32540 3555
rect 33185 3065 33200 3665
rect 33240 3065 33255 3665
rect 33295 3065 33310 3665
rect 33350 3065 33365 3665
rect 33405 3065 33420 3665
rect 33460 3065 33475 3665
rect 33515 3065 33530 3665
rect 33570 3065 33585 3665
rect 33625 3065 33640 3665
rect 33680 3065 33695 3665
rect 33735 3065 33750 3665
rect 33790 3065 33805 3665
rect 29995 2505 30010 2705
rect 30050 2505 30065 2705
rect 30105 2505 30120 2705
rect 30160 2505 30175 2705
rect 30215 2505 30230 2705
rect 30270 2505 30285 2705
rect 30325 2505 30340 2705
rect 30380 2505 30395 2705
rect 30435 2505 30450 2705
rect 30490 2505 30505 2705
rect 30545 2505 30560 2705
rect 30600 2505 30615 2705
rect 31045 2495 31065 2845
rect 31105 2495 31125 2845
rect 31165 2495 31185 2845
rect 31225 2495 31245 2845
rect 31285 2495 31305 2845
rect 31345 2495 31365 2845
rect 31405 2495 31425 2845
rect 31465 2495 31485 2845
rect 31525 2495 31545 2845
rect 31585 2495 31605 2845
rect 31645 2495 31665 2845
rect 31705 2495 31725 2845
rect 32075 2495 32095 2845
rect 32135 2495 32155 2845
rect 32195 2495 32215 2845
rect 32255 2495 32275 2845
rect 32315 2495 32335 2845
rect 32375 2495 32395 2845
rect 32435 2495 32455 2845
rect 32495 2495 32515 2845
rect 32555 2495 32575 2845
rect 32615 2495 32635 2845
rect 32675 2495 32695 2845
rect 32735 2495 32755 2845
rect 33185 2505 33200 2705
rect 33240 2505 33255 2705
rect 33295 2505 33310 2705
rect 33350 2505 33365 2705
rect 33405 2505 33420 2705
rect 33460 2505 33475 2705
rect 33515 2505 33530 2705
rect 33570 2505 33585 2705
rect 33625 2505 33640 2705
rect 33680 2505 33695 2705
rect 33735 2505 33750 2705
rect 33790 2505 33805 2705
<< ndiff >>
rect 29955 2230 29995 2245
rect 29955 2210 29965 2230
rect 29985 2210 29995 2230
rect 29955 2180 29995 2210
rect 29955 2160 29965 2180
rect 29985 2160 29995 2180
rect 29955 2130 29995 2160
rect 29955 2110 29965 2130
rect 29985 2110 29995 2130
rect 29955 2080 29995 2110
rect 29955 2060 29965 2080
rect 29985 2060 29995 2080
rect 29955 2030 29995 2060
rect 29955 2010 29965 2030
rect 29985 2010 29995 2030
rect 29955 1980 29995 2010
rect 29955 1960 29965 1980
rect 29985 1960 29995 1980
rect 29955 1945 29995 1960
rect 30010 2230 30050 2245
rect 30010 2210 30020 2230
rect 30040 2210 30050 2230
rect 30010 2180 30050 2210
rect 30010 2160 30020 2180
rect 30040 2160 30050 2180
rect 30010 2130 30050 2160
rect 30010 2110 30020 2130
rect 30040 2110 30050 2130
rect 30010 2080 30050 2110
rect 30010 2060 30020 2080
rect 30040 2060 30050 2080
rect 30010 2030 30050 2060
rect 30010 2010 30020 2030
rect 30040 2010 30050 2030
rect 30010 1980 30050 2010
rect 30010 1960 30020 1980
rect 30040 1960 30050 1980
rect 30010 1945 30050 1960
rect 30065 2230 30105 2245
rect 30065 2210 30075 2230
rect 30095 2210 30105 2230
rect 30065 2180 30105 2210
rect 30065 2160 30075 2180
rect 30095 2160 30105 2180
rect 30065 2130 30105 2160
rect 30065 2110 30075 2130
rect 30095 2110 30105 2130
rect 30065 2080 30105 2110
rect 30065 2060 30075 2080
rect 30095 2060 30105 2080
rect 30065 2030 30105 2060
rect 30065 2010 30075 2030
rect 30095 2010 30105 2030
rect 30065 1980 30105 2010
rect 30065 1960 30075 1980
rect 30095 1960 30105 1980
rect 30065 1945 30105 1960
rect 30120 2230 30160 2245
rect 30120 2210 30130 2230
rect 30150 2210 30160 2230
rect 30120 2180 30160 2210
rect 30120 2160 30130 2180
rect 30150 2160 30160 2180
rect 30120 2130 30160 2160
rect 30120 2110 30130 2130
rect 30150 2110 30160 2130
rect 30120 2080 30160 2110
rect 30120 2060 30130 2080
rect 30150 2060 30160 2080
rect 30120 2030 30160 2060
rect 30120 2010 30130 2030
rect 30150 2010 30160 2030
rect 30120 1980 30160 2010
rect 30120 1960 30130 1980
rect 30150 1960 30160 1980
rect 30120 1945 30160 1960
rect 30175 2230 30215 2245
rect 30175 2210 30185 2230
rect 30205 2210 30215 2230
rect 30175 2180 30215 2210
rect 30175 2160 30185 2180
rect 30205 2160 30215 2180
rect 30175 2130 30215 2160
rect 30175 2110 30185 2130
rect 30205 2110 30215 2130
rect 30175 2080 30215 2110
rect 30175 2060 30185 2080
rect 30205 2060 30215 2080
rect 30175 2030 30215 2060
rect 30175 2010 30185 2030
rect 30205 2010 30215 2030
rect 30175 1980 30215 2010
rect 30175 1960 30185 1980
rect 30205 1960 30215 1980
rect 30175 1945 30215 1960
rect 30230 2230 30270 2245
rect 30230 2210 30240 2230
rect 30260 2210 30270 2230
rect 30230 2180 30270 2210
rect 30230 2160 30240 2180
rect 30260 2160 30270 2180
rect 30230 2130 30270 2160
rect 30230 2110 30240 2130
rect 30260 2110 30270 2130
rect 30230 2080 30270 2110
rect 30230 2060 30240 2080
rect 30260 2060 30270 2080
rect 30230 2030 30270 2060
rect 30230 2010 30240 2030
rect 30260 2010 30270 2030
rect 30230 1980 30270 2010
rect 30230 1960 30240 1980
rect 30260 1960 30270 1980
rect 30230 1945 30270 1960
rect 30285 2230 30325 2245
rect 30285 2210 30295 2230
rect 30315 2210 30325 2230
rect 30285 2180 30325 2210
rect 30285 2160 30295 2180
rect 30315 2160 30325 2180
rect 30285 2130 30325 2160
rect 30285 2110 30295 2130
rect 30315 2110 30325 2130
rect 30285 2080 30325 2110
rect 30285 2060 30295 2080
rect 30315 2060 30325 2080
rect 30285 2030 30325 2060
rect 30285 2010 30295 2030
rect 30315 2010 30325 2030
rect 30285 1980 30325 2010
rect 30285 1960 30295 1980
rect 30315 1960 30325 1980
rect 30285 1945 30325 1960
rect 30340 2230 30380 2245
rect 30340 2210 30350 2230
rect 30370 2210 30380 2230
rect 30340 2180 30380 2210
rect 30340 2160 30350 2180
rect 30370 2160 30380 2180
rect 30340 2130 30380 2160
rect 30340 2110 30350 2130
rect 30370 2110 30380 2130
rect 30340 2080 30380 2110
rect 30340 2060 30350 2080
rect 30370 2060 30380 2080
rect 30340 2030 30380 2060
rect 30340 2010 30350 2030
rect 30370 2010 30380 2030
rect 30340 1980 30380 2010
rect 30340 1960 30350 1980
rect 30370 1960 30380 1980
rect 30340 1945 30380 1960
rect 30395 2230 30435 2245
rect 30395 2210 30405 2230
rect 30425 2210 30435 2230
rect 30395 2180 30435 2210
rect 30395 2160 30405 2180
rect 30425 2160 30435 2180
rect 30395 2130 30435 2160
rect 30395 2110 30405 2130
rect 30425 2110 30435 2130
rect 30395 2080 30435 2110
rect 30395 2060 30405 2080
rect 30425 2060 30435 2080
rect 30395 2030 30435 2060
rect 30395 2010 30405 2030
rect 30425 2010 30435 2030
rect 30395 1980 30435 2010
rect 30395 1960 30405 1980
rect 30425 1960 30435 1980
rect 30395 1945 30435 1960
rect 30450 2230 30490 2245
rect 30450 2210 30460 2230
rect 30480 2210 30490 2230
rect 30450 2180 30490 2210
rect 30450 2160 30460 2180
rect 30480 2160 30490 2180
rect 30450 2130 30490 2160
rect 30450 2110 30460 2130
rect 30480 2110 30490 2130
rect 30450 2080 30490 2110
rect 30450 2060 30460 2080
rect 30480 2060 30490 2080
rect 30450 2030 30490 2060
rect 30450 2010 30460 2030
rect 30480 2010 30490 2030
rect 30450 1980 30490 2010
rect 30450 1960 30460 1980
rect 30480 1960 30490 1980
rect 30450 1945 30490 1960
rect 30505 2230 30545 2245
rect 30505 2210 30515 2230
rect 30535 2210 30545 2230
rect 30505 2180 30545 2210
rect 30505 2160 30515 2180
rect 30535 2160 30545 2180
rect 30505 2130 30545 2160
rect 30505 2110 30515 2130
rect 30535 2110 30545 2130
rect 30505 2080 30545 2110
rect 30505 2060 30515 2080
rect 30535 2060 30545 2080
rect 30505 2030 30545 2060
rect 30505 2010 30515 2030
rect 30535 2010 30545 2030
rect 30505 1980 30545 2010
rect 30505 1960 30515 1980
rect 30535 1960 30545 1980
rect 30505 1945 30545 1960
rect 30560 2230 30600 2245
rect 30560 2210 30570 2230
rect 30590 2210 30600 2230
rect 30560 2180 30600 2210
rect 30560 2160 30570 2180
rect 30590 2160 30600 2180
rect 30560 2130 30600 2160
rect 30560 2110 30570 2130
rect 30590 2110 30600 2130
rect 30560 2080 30600 2110
rect 30560 2060 30570 2080
rect 30590 2060 30600 2080
rect 30560 2030 30600 2060
rect 30560 2010 30570 2030
rect 30590 2010 30600 2030
rect 30560 1980 30600 2010
rect 30560 1960 30570 1980
rect 30590 1960 30600 1980
rect 30560 1945 30600 1960
rect 30615 2230 30655 2245
rect 30615 2210 30625 2230
rect 30645 2210 30655 2230
rect 30615 2180 30655 2210
rect 30615 2160 30625 2180
rect 30645 2160 30655 2180
rect 30615 2130 30655 2160
rect 30615 2110 30625 2130
rect 30645 2110 30655 2130
rect 30615 2080 30655 2110
rect 30615 2060 30625 2080
rect 30645 2060 30655 2080
rect 30615 2030 30655 2060
rect 30615 2010 30625 2030
rect 30645 2010 30655 2030
rect 30615 1980 30655 2010
rect 30615 1960 30625 1980
rect 30645 1960 30655 1980
rect 30615 1945 30655 1960
rect 31185 2165 31225 2180
rect 31185 2145 31195 2165
rect 31215 2145 31225 2165
rect 31185 2115 31225 2145
rect 31185 2095 31195 2115
rect 31215 2095 31225 2115
rect 31185 2065 31225 2095
rect 31185 2045 31195 2065
rect 31215 2045 31225 2065
rect 31185 2030 31225 2045
rect 31240 2165 31280 2180
rect 31240 2145 31250 2165
rect 31270 2145 31280 2165
rect 31240 2115 31280 2145
rect 31240 2095 31250 2115
rect 31270 2095 31280 2115
rect 31240 2065 31280 2095
rect 31240 2045 31250 2065
rect 31270 2045 31280 2065
rect 31240 2030 31280 2045
rect 31295 2165 31335 2180
rect 31295 2145 31305 2165
rect 31325 2145 31335 2165
rect 31295 2115 31335 2145
rect 31295 2095 31305 2115
rect 31325 2095 31335 2115
rect 31295 2065 31335 2095
rect 31295 2045 31305 2065
rect 31325 2045 31335 2065
rect 31295 2030 31335 2045
rect 31350 2165 31390 2180
rect 31350 2145 31360 2165
rect 31380 2145 31390 2165
rect 31350 2115 31390 2145
rect 31350 2095 31360 2115
rect 31380 2095 31390 2115
rect 31350 2065 31390 2095
rect 31350 2045 31360 2065
rect 31380 2045 31390 2065
rect 31350 2030 31390 2045
rect 31405 2165 31445 2180
rect 31405 2145 31415 2165
rect 31435 2145 31445 2165
rect 31405 2115 31445 2145
rect 31405 2095 31415 2115
rect 31435 2095 31445 2115
rect 31405 2065 31445 2095
rect 31405 2045 31415 2065
rect 31435 2045 31445 2065
rect 31405 2030 31445 2045
rect 31460 2165 31500 2180
rect 31460 2145 31470 2165
rect 31490 2145 31500 2165
rect 31460 2115 31500 2145
rect 31460 2095 31470 2115
rect 31490 2095 31500 2115
rect 31460 2065 31500 2095
rect 31460 2045 31470 2065
rect 31490 2045 31500 2065
rect 31460 2030 31500 2045
rect 31515 2165 31555 2180
rect 31515 2145 31525 2165
rect 31545 2145 31555 2165
rect 31515 2115 31555 2145
rect 31515 2095 31525 2115
rect 31545 2095 31555 2115
rect 31515 2065 31555 2095
rect 31515 2045 31525 2065
rect 31545 2045 31555 2065
rect 31515 2030 31555 2045
rect 31570 2165 31610 2180
rect 31570 2145 31580 2165
rect 31600 2145 31610 2165
rect 31570 2115 31610 2145
rect 31570 2095 31580 2115
rect 31600 2095 31610 2115
rect 31570 2065 31610 2095
rect 31570 2045 31580 2065
rect 31600 2045 31610 2065
rect 31570 2030 31610 2045
rect 31625 2165 31665 2180
rect 31625 2145 31635 2165
rect 31655 2145 31665 2165
rect 31625 2115 31665 2145
rect 31625 2095 31635 2115
rect 31655 2095 31665 2115
rect 31625 2065 31665 2095
rect 31625 2045 31635 2065
rect 31655 2045 31665 2065
rect 31625 2030 31665 2045
rect 31680 2165 31720 2180
rect 31680 2145 31690 2165
rect 31710 2145 31720 2165
rect 31680 2115 31720 2145
rect 31680 2095 31690 2115
rect 31710 2095 31720 2115
rect 31680 2065 31720 2095
rect 31680 2045 31690 2065
rect 31710 2045 31720 2065
rect 31680 2030 31720 2045
rect 31735 2165 31775 2180
rect 31735 2145 31745 2165
rect 31765 2145 31775 2165
rect 31735 2115 31775 2145
rect 31735 2095 31745 2115
rect 31765 2095 31775 2115
rect 31735 2065 31775 2095
rect 31735 2045 31745 2065
rect 31765 2045 31775 2065
rect 31735 2030 31775 2045
rect 31790 2165 31830 2180
rect 31790 2145 31800 2165
rect 31820 2145 31830 2165
rect 31790 2115 31830 2145
rect 31790 2095 31800 2115
rect 31820 2095 31830 2115
rect 31790 2065 31830 2095
rect 31790 2045 31800 2065
rect 31820 2045 31830 2065
rect 31790 2030 31830 2045
rect 31845 2165 31885 2180
rect 31845 2145 31855 2165
rect 31875 2145 31885 2165
rect 31845 2115 31885 2145
rect 31845 2095 31855 2115
rect 31875 2095 31885 2115
rect 31845 2065 31885 2095
rect 31845 2045 31855 2065
rect 31875 2045 31885 2065
rect 31845 2030 31885 2045
rect 31915 2165 31955 2180
rect 31915 2145 31925 2165
rect 31945 2145 31955 2165
rect 31915 2115 31955 2145
rect 31915 2095 31925 2115
rect 31945 2095 31955 2115
rect 31915 2065 31955 2095
rect 31915 2045 31925 2065
rect 31945 2045 31955 2065
rect 31915 2030 31955 2045
rect 31970 2165 32010 2180
rect 31970 2145 31980 2165
rect 32000 2145 32010 2165
rect 31970 2115 32010 2145
rect 31970 2095 31980 2115
rect 32000 2095 32010 2115
rect 31970 2065 32010 2095
rect 31970 2045 31980 2065
rect 32000 2045 32010 2065
rect 31970 2030 32010 2045
rect 32025 2165 32065 2180
rect 32025 2145 32035 2165
rect 32055 2145 32065 2165
rect 32025 2115 32065 2145
rect 32025 2095 32035 2115
rect 32055 2095 32065 2115
rect 32025 2065 32065 2095
rect 32025 2045 32035 2065
rect 32055 2045 32065 2065
rect 32025 2030 32065 2045
rect 32080 2165 32120 2180
rect 32080 2145 32090 2165
rect 32110 2145 32120 2165
rect 32080 2115 32120 2145
rect 32080 2095 32090 2115
rect 32110 2095 32120 2115
rect 32080 2065 32120 2095
rect 32080 2045 32090 2065
rect 32110 2045 32120 2065
rect 32080 2030 32120 2045
rect 32135 2165 32175 2180
rect 32135 2145 32145 2165
rect 32165 2145 32175 2165
rect 32135 2115 32175 2145
rect 32135 2095 32145 2115
rect 32165 2095 32175 2115
rect 32135 2065 32175 2095
rect 32135 2045 32145 2065
rect 32165 2045 32175 2065
rect 32135 2030 32175 2045
rect 32190 2165 32230 2180
rect 32190 2145 32200 2165
rect 32220 2145 32230 2165
rect 32190 2115 32230 2145
rect 32190 2095 32200 2115
rect 32220 2095 32230 2115
rect 32190 2065 32230 2095
rect 32190 2045 32200 2065
rect 32220 2045 32230 2065
rect 32190 2030 32230 2045
rect 32245 2165 32285 2180
rect 32245 2145 32255 2165
rect 32275 2145 32285 2165
rect 32245 2115 32285 2145
rect 32245 2095 32255 2115
rect 32275 2095 32285 2115
rect 32245 2065 32285 2095
rect 32245 2045 32255 2065
rect 32275 2045 32285 2065
rect 32245 2030 32285 2045
rect 32300 2165 32340 2180
rect 32300 2145 32310 2165
rect 32330 2145 32340 2165
rect 32300 2115 32340 2145
rect 32300 2095 32310 2115
rect 32330 2095 32340 2115
rect 32300 2065 32340 2095
rect 32300 2045 32310 2065
rect 32330 2045 32340 2065
rect 32300 2030 32340 2045
rect 32355 2165 32395 2180
rect 32355 2145 32365 2165
rect 32385 2145 32395 2165
rect 32355 2115 32395 2145
rect 32355 2095 32365 2115
rect 32385 2095 32395 2115
rect 32355 2065 32395 2095
rect 32355 2045 32365 2065
rect 32385 2045 32395 2065
rect 32355 2030 32395 2045
rect 32410 2165 32450 2180
rect 32410 2145 32420 2165
rect 32440 2145 32450 2165
rect 32410 2115 32450 2145
rect 32410 2095 32420 2115
rect 32440 2095 32450 2115
rect 32410 2065 32450 2095
rect 32410 2045 32420 2065
rect 32440 2045 32450 2065
rect 32410 2030 32450 2045
rect 32465 2165 32505 2180
rect 32465 2145 32475 2165
rect 32495 2145 32505 2165
rect 32465 2115 32505 2145
rect 32465 2095 32475 2115
rect 32495 2095 32505 2115
rect 32465 2065 32505 2095
rect 32465 2045 32475 2065
rect 32495 2045 32505 2065
rect 32465 2030 32505 2045
rect 32520 2165 32560 2180
rect 32520 2145 32530 2165
rect 32550 2145 32560 2165
rect 32520 2115 32560 2145
rect 32520 2095 32530 2115
rect 32550 2095 32560 2115
rect 32520 2065 32560 2095
rect 32520 2045 32530 2065
rect 32550 2045 32560 2065
rect 32520 2030 32560 2045
rect 32575 2165 32615 2180
rect 32575 2145 32585 2165
rect 32605 2145 32615 2165
rect 32575 2115 32615 2145
rect 32575 2095 32585 2115
rect 32605 2095 32615 2115
rect 32575 2065 32615 2095
rect 32575 2045 32585 2065
rect 32605 2045 32615 2065
rect 32575 2030 32615 2045
rect 33145 2230 33185 2245
rect 33145 2210 33155 2230
rect 33175 2210 33185 2230
rect 33145 2180 33185 2210
rect 33145 2160 33155 2180
rect 33175 2160 33185 2180
rect 33145 2130 33185 2160
rect 33145 2110 33155 2130
rect 33175 2110 33185 2130
rect 33145 2080 33185 2110
rect 33145 2060 33155 2080
rect 33175 2060 33185 2080
rect 33145 2030 33185 2060
rect 33145 2010 33155 2030
rect 33175 2010 33185 2030
rect 33145 1980 33185 2010
rect 33145 1960 33155 1980
rect 33175 1960 33185 1980
rect 33145 1945 33185 1960
rect 33200 2230 33240 2245
rect 33200 2210 33210 2230
rect 33230 2210 33240 2230
rect 33200 2180 33240 2210
rect 33200 2160 33210 2180
rect 33230 2160 33240 2180
rect 33200 2130 33240 2160
rect 33200 2110 33210 2130
rect 33230 2110 33240 2130
rect 33200 2080 33240 2110
rect 33200 2060 33210 2080
rect 33230 2060 33240 2080
rect 33200 2030 33240 2060
rect 33200 2010 33210 2030
rect 33230 2010 33240 2030
rect 33200 1980 33240 2010
rect 33200 1960 33210 1980
rect 33230 1960 33240 1980
rect 33200 1945 33240 1960
rect 33255 2230 33295 2245
rect 33255 2210 33265 2230
rect 33285 2210 33295 2230
rect 33255 2180 33295 2210
rect 33255 2160 33265 2180
rect 33285 2160 33295 2180
rect 33255 2130 33295 2160
rect 33255 2110 33265 2130
rect 33285 2110 33295 2130
rect 33255 2080 33295 2110
rect 33255 2060 33265 2080
rect 33285 2060 33295 2080
rect 33255 2030 33295 2060
rect 33255 2010 33265 2030
rect 33285 2010 33295 2030
rect 33255 1980 33295 2010
rect 33255 1960 33265 1980
rect 33285 1960 33295 1980
rect 33255 1945 33295 1960
rect 33310 2230 33350 2245
rect 33310 2210 33320 2230
rect 33340 2210 33350 2230
rect 33310 2180 33350 2210
rect 33310 2160 33320 2180
rect 33340 2160 33350 2180
rect 33310 2130 33350 2160
rect 33310 2110 33320 2130
rect 33340 2110 33350 2130
rect 33310 2080 33350 2110
rect 33310 2060 33320 2080
rect 33340 2060 33350 2080
rect 33310 2030 33350 2060
rect 33310 2010 33320 2030
rect 33340 2010 33350 2030
rect 33310 1980 33350 2010
rect 33310 1960 33320 1980
rect 33340 1960 33350 1980
rect 33310 1945 33350 1960
rect 33365 2230 33405 2245
rect 33365 2210 33375 2230
rect 33395 2210 33405 2230
rect 33365 2180 33405 2210
rect 33365 2160 33375 2180
rect 33395 2160 33405 2180
rect 33365 2130 33405 2160
rect 33365 2110 33375 2130
rect 33395 2110 33405 2130
rect 33365 2080 33405 2110
rect 33365 2060 33375 2080
rect 33395 2060 33405 2080
rect 33365 2030 33405 2060
rect 33365 2010 33375 2030
rect 33395 2010 33405 2030
rect 33365 1980 33405 2010
rect 33365 1960 33375 1980
rect 33395 1960 33405 1980
rect 33365 1945 33405 1960
rect 33420 2230 33460 2245
rect 33420 2210 33430 2230
rect 33450 2210 33460 2230
rect 33420 2180 33460 2210
rect 33420 2160 33430 2180
rect 33450 2160 33460 2180
rect 33420 2130 33460 2160
rect 33420 2110 33430 2130
rect 33450 2110 33460 2130
rect 33420 2080 33460 2110
rect 33420 2060 33430 2080
rect 33450 2060 33460 2080
rect 33420 2030 33460 2060
rect 33420 2010 33430 2030
rect 33450 2010 33460 2030
rect 33420 1980 33460 2010
rect 33420 1960 33430 1980
rect 33450 1960 33460 1980
rect 33420 1945 33460 1960
rect 33475 2230 33515 2245
rect 33475 2210 33485 2230
rect 33505 2210 33515 2230
rect 33475 2180 33515 2210
rect 33475 2160 33485 2180
rect 33505 2160 33515 2180
rect 33475 2130 33515 2160
rect 33475 2110 33485 2130
rect 33505 2110 33515 2130
rect 33475 2080 33515 2110
rect 33475 2060 33485 2080
rect 33505 2060 33515 2080
rect 33475 2030 33515 2060
rect 33475 2010 33485 2030
rect 33505 2010 33515 2030
rect 33475 1980 33515 2010
rect 33475 1960 33485 1980
rect 33505 1960 33515 1980
rect 33475 1945 33515 1960
rect 33530 2230 33570 2245
rect 33530 2210 33540 2230
rect 33560 2210 33570 2230
rect 33530 2180 33570 2210
rect 33530 2160 33540 2180
rect 33560 2160 33570 2180
rect 33530 2130 33570 2160
rect 33530 2110 33540 2130
rect 33560 2110 33570 2130
rect 33530 2080 33570 2110
rect 33530 2060 33540 2080
rect 33560 2060 33570 2080
rect 33530 2030 33570 2060
rect 33530 2010 33540 2030
rect 33560 2010 33570 2030
rect 33530 1980 33570 2010
rect 33530 1960 33540 1980
rect 33560 1960 33570 1980
rect 33530 1945 33570 1960
rect 33585 2230 33625 2245
rect 33585 2210 33595 2230
rect 33615 2210 33625 2230
rect 33585 2180 33625 2210
rect 33585 2160 33595 2180
rect 33615 2160 33625 2180
rect 33585 2130 33625 2160
rect 33585 2110 33595 2130
rect 33615 2110 33625 2130
rect 33585 2080 33625 2110
rect 33585 2060 33595 2080
rect 33615 2060 33625 2080
rect 33585 2030 33625 2060
rect 33585 2010 33595 2030
rect 33615 2010 33625 2030
rect 33585 1980 33625 2010
rect 33585 1960 33595 1980
rect 33615 1960 33625 1980
rect 33585 1945 33625 1960
rect 33640 2230 33680 2245
rect 33640 2210 33650 2230
rect 33670 2210 33680 2230
rect 33640 2180 33680 2210
rect 33640 2160 33650 2180
rect 33670 2160 33680 2180
rect 33640 2130 33680 2160
rect 33640 2110 33650 2130
rect 33670 2110 33680 2130
rect 33640 2080 33680 2110
rect 33640 2060 33650 2080
rect 33670 2060 33680 2080
rect 33640 2030 33680 2060
rect 33640 2010 33650 2030
rect 33670 2010 33680 2030
rect 33640 1980 33680 2010
rect 33640 1960 33650 1980
rect 33670 1960 33680 1980
rect 33640 1945 33680 1960
rect 33695 2230 33735 2245
rect 33695 2210 33705 2230
rect 33725 2210 33735 2230
rect 33695 2180 33735 2210
rect 33695 2160 33705 2180
rect 33725 2160 33735 2180
rect 33695 2130 33735 2160
rect 33695 2110 33705 2130
rect 33725 2110 33735 2130
rect 33695 2080 33735 2110
rect 33695 2060 33705 2080
rect 33725 2060 33735 2080
rect 33695 2030 33735 2060
rect 33695 2010 33705 2030
rect 33725 2010 33735 2030
rect 33695 1980 33735 2010
rect 33695 1960 33705 1980
rect 33725 1960 33735 1980
rect 33695 1945 33735 1960
rect 33750 2230 33790 2245
rect 33750 2210 33760 2230
rect 33780 2210 33790 2230
rect 33750 2180 33790 2210
rect 33750 2160 33760 2180
rect 33780 2160 33790 2180
rect 33750 2130 33790 2160
rect 33750 2110 33760 2130
rect 33780 2110 33790 2130
rect 33750 2080 33790 2110
rect 33750 2060 33760 2080
rect 33780 2060 33790 2080
rect 33750 2030 33790 2060
rect 33750 2010 33760 2030
rect 33780 2010 33790 2030
rect 33750 1980 33790 2010
rect 33750 1960 33760 1980
rect 33780 1960 33790 1980
rect 33750 1945 33790 1960
rect 33805 2230 33845 2245
rect 33805 2210 33815 2230
rect 33835 2210 33845 2230
rect 33805 2180 33845 2210
rect 33805 2160 33815 2180
rect 33835 2160 33845 2180
rect 33805 2130 33845 2160
rect 33805 2110 33815 2130
rect 33835 2110 33845 2130
rect 33805 2080 33845 2110
rect 33805 2060 33815 2080
rect 33835 2060 33845 2080
rect 33805 2030 33845 2060
rect 33805 2010 33815 2030
rect 33835 2010 33845 2030
rect 33805 1980 33845 2010
rect 33805 1960 33815 1980
rect 33835 1960 33845 1980
rect 33805 1945 33845 1960
rect 30035 1640 30075 1655
rect 30035 1620 30045 1640
rect 30065 1620 30075 1640
rect 30035 1590 30075 1620
rect 30035 1570 30045 1590
rect 30065 1570 30075 1590
rect 30035 1540 30075 1570
rect 30035 1520 30045 1540
rect 30065 1520 30075 1540
rect 30035 1490 30075 1520
rect 30035 1470 30045 1490
rect 30065 1470 30075 1490
rect 30035 1440 30075 1470
rect 30035 1420 30045 1440
rect 30065 1420 30075 1440
rect 30035 1390 30075 1420
rect 30035 1370 30045 1390
rect 30065 1370 30075 1390
rect 30035 1340 30075 1370
rect 30035 1320 30045 1340
rect 30065 1320 30075 1340
rect 30035 1290 30075 1320
rect 30035 1270 30045 1290
rect 30065 1270 30075 1290
rect 30035 1240 30075 1270
rect 30035 1220 30045 1240
rect 30065 1220 30075 1240
rect 30035 1190 30075 1220
rect 30035 1170 30045 1190
rect 30065 1170 30075 1190
rect 30035 1140 30075 1170
rect 30035 1120 30045 1140
rect 30065 1120 30075 1140
rect 30035 1090 30075 1120
rect 30035 1070 30045 1090
rect 30065 1070 30075 1090
rect 30035 1040 30075 1070
rect 30035 1020 30045 1040
rect 30065 1020 30075 1040
rect 30035 990 30075 1020
rect 30035 970 30045 990
rect 30065 970 30075 990
rect 30035 955 30075 970
rect 30135 1640 30175 1655
rect 30135 1620 30145 1640
rect 30165 1620 30175 1640
rect 30135 1590 30175 1620
rect 30135 1570 30145 1590
rect 30165 1570 30175 1590
rect 30135 1540 30175 1570
rect 30135 1520 30145 1540
rect 30165 1520 30175 1540
rect 30135 1490 30175 1520
rect 30135 1470 30145 1490
rect 30165 1470 30175 1490
rect 30135 1440 30175 1470
rect 30135 1420 30145 1440
rect 30165 1420 30175 1440
rect 30135 1390 30175 1420
rect 30135 1370 30145 1390
rect 30165 1370 30175 1390
rect 30135 1340 30175 1370
rect 30135 1320 30145 1340
rect 30165 1320 30175 1340
rect 30135 1290 30175 1320
rect 30135 1270 30145 1290
rect 30165 1270 30175 1290
rect 30135 1240 30175 1270
rect 30135 1220 30145 1240
rect 30165 1220 30175 1240
rect 30135 1190 30175 1220
rect 30135 1170 30145 1190
rect 30165 1170 30175 1190
rect 30135 1140 30175 1170
rect 30135 1120 30145 1140
rect 30165 1120 30175 1140
rect 30135 1090 30175 1120
rect 30135 1070 30145 1090
rect 30165 1070 30175 1090
rect 30135 1040 30175 1070
rect 30135 1020 30145 1040
rect 30165 1020 30175 1040
rect 30135 990 30175 1020
rect 30135 970 30145 990
rect 30165 970 30175 990
rect 30135 955 30175 970
rect 30235 1640 30275 1655
rect 30235 1620 30245 1640
rect 30265 1620 30275 1640
rect 30235 1590 30275 1620
rect 30235 1570 30245 1590
rect 30265 1570 30275 1590
rect 30235 1540 30275 1570
rect 30235 1520 30245 1540
rect 30265 1520 30275 1540
rect 30235 1490 30275 1520
rect 30235 1470 30245 1490
rect 30265 1470 30275 1490
rect 30235 1440 30275 1470
rect 30235 1420 30245 1440
rect 30265 1420 30275 1440
rect 30235 1390 30275 1420
rect 30235 1370 30245 1390
rect 30265 1370 30275 1390
rect 30235 1340 30275 1370
rect 30235 1320 30245 1340
rect 30265 1320 30275 1340
rect 30235 1290 30275 1320
rect 30235 1270 30245 1290
rect 30265 1270 30275 1290
rect 30235 1240 30275 1270
rect 30235 1220 30245 1240
rect 30265 1220 30275 1240
rect 30235 1190 30275 1220
rect 30235 1170 30245 1190
rect 30265 1170 30275 1190
rect 30235 1140 30275 1170
rect 30235 1120 30245 1140
rect 30265 1120 30275 1140
rect 30235 1090 30275 1120
rect 30235 1070 30245 1090
rect 30265 1070 30275 1090
rect 30235 1040 30275 1070
rect 30235 1020 30245 1040
rect 30265 1020 30275 1040
rect 30235 990 30275 1020
rect 30235 970 30245 990
rect 30265 970 30275 990
rect 30235 955 30275 970
rect 30335 1640 30375 1655
rect 30335 1620 30345 1640
rect 30365 1620 30375 1640
rect 30335 1590 30375 1620
rect 30335 1570 30345 1590
rect 30365 1570 30375 1590
rect 30335 1540 30375 1570
rect 30335 1520 30345 1540
rect 30365 1520 30375 1540
rect 30335 1490 30375 1520
rect 30335 1470 30345 1490
rect 30365 1470 30375 1490
rect 30335 1440 30375 1470
rect 30335 1420 30345 1440
rect 30365 1420 30375 1440
rect 30335 1390 30375 1420
rect 30335 1370 30345 1390
rect 30365 1370 30375 1390
rect 30335 1340 30375 1370
rect 30335 1320 30345 1340
rect 30365 1320 30375 1340
rect 30335 1290 30375 1320
rect 30335 1270 30345 1290
rect 30365 1270 30375 1290
rect 30335 1240 30375 1270
rect 30335 1220 30345 1240
rect 30365 1220 30375 1240
rect 30335 1190 30375 1220
rect 30335 1170 30345 1190
rect 30365 1170 30375 1190
rect 30335 1140 30375 1170
rect 30335 1120 30345 1140
rect 30365 1120 30375 1140
rect 30335 1090 30375 1120
rect 30335 1070 30345 1090
rect 30365 1070 30375 1090
rect 30335 1040 30375 1070
rect 30335 1020 30345 1040
rect 30365 1020 30375 1040
rect 30335 990 30375 1020
rect 30335 970 30345 990
rect 30365 970 30375 990
rect 30335 955 30375 970
rect 30435 1640 30475 1655
rect 30435 1620 30445 1640
rect 30465 1620 30475 1640
rect 30435 1590 30475 1620
rect 30435 1570 30445 1590
rect 30465 1570 30475 1590
rect 30435 1540 30475 1570
rect 30435 1520 30445 1540
rect 30465 1520 30475 1540
rect 30435 1490 30475 1520
rect 30435 1470 30445 1490
rect 30465 1470 30475 1490
rect 30435 1440 30475 1470
rect 30435 1420 30445 1440
rect 30465 1420 30475 1440
rect 30435 1390 30475 1420
rect 30435 1370 30445 1390
rect 30465 1370 30475 1390
rect 30435 1340 30475 1370
rect 30435 1320 30445 1340
rect 30465 1320 30475 1340
rect 30435 1290 30475 1320
rect 30435 1270 30445 1290
rect 30465 1270 30475 1290
rect 30435 1240 30475 1270
rect 30435 1220 30445 1240
rect 30465 1220 30475 1240
rect 30435 1190 30475 1220
rect 30435 1170 30445 1190
rect 30465 1170 30475 1190
rect 30435 1140 30475 1170
rect 30435 1120 30445 1140
rect 30465 1120 30475 1140
rect 30435 1090 30475 1120
rect 30435 1070 30445 1090
rect 30465 1070 30475 1090
rect 30435 1040 30475 1070
rect 30435 1020 30445 1040
rect 30465 1020 30475 1040
rect 30435 990 30475 1020
rect 30435 970 30445 990
rect 30465 970 30475 990
rect 30435 955 30475 970
rect 30535 1640 30575 1655
rect 30535 1620 30545 1640
rect 30565 1620 30575 1640
rect 30535 1590 30575 1620
rect 30535 1570 30545 1590
rect 30565 1570 30575 1590
rect 30535 1540 30575 1570
rect 30535 1520 30545 1540
rect 30565 1520 30575 1540
rect 30535 1490 30575 1520
rect 30535 1470 30545 1490
rect 30565 1470 30575 1490
rect 30535 1440 30575 1470
rect 30535 1420 30545 1440
rect 30565 1420 30575 1440
rect 30535 1390 30575 1420
rect 30535 1370 30545 1390
rect 30565 1370 30575 1390
rect 30535 1340 30575 1370
rect 30535 1320 30545 1340
rect 30565 1320 30575 1340
rect 30535 1290 30575 1320
rect 30535 1270 30545 1290
rect 30565 1270 30575 1290
rect 30535 1240 30575 1270
rect 30535 1220 30545 1240
rect 30565 1220 30575 1240
rect 30535 1190 30575 1220
rect 30535 1170 30545 1190
rect 30565 1170 30575 1190
rect 30535 1140 30575 1170
rect 30535 1120 30545 1140
rect 30565 1120 30575 1140
rect 30535 1090 30575 1120
rect 30535 1070 30545 1090
rect 30565 1070 30575 1090
rect 30535 1040 30575 1070
rect 30535 1020 30545 1040
rect 30565 1020 30575 1040
rect 30535 990 30575 1020
rect 30535 970 30545 990
rect 30565 970 30575 990
rect 30535 955 30575 970
rect 30635 1640 30675 1655
rect 30635 1620 30645 1640
rect 30665 1620 30675 1640
rect 30635 1590 30675 1620
rect 30635 1570 30645 1590
rect 30665 1570 30675 1590
rect 30635 1540 30675 1570
rect 30635 1520 30645 1540
rect 30665 1520 30675 1540
rect 30635 1490 30675 1520
rect 30635 1470 30645 1490
rect 30665 1470 30675 1490
rect 30635 1440 30675 1470
rect 30635 1420 30645 1440
rect 30665 1420 30675 1440
rect 30635 1390 30675 1420
rect 30635 1370 30645 1390
rect 30665 1370 30675 1390
rect 30635 1340 30675 1370
rect 30635 1320 30645 1340
rect 30665 1320 30675 1340
rect 30635 1290 30675 1320
rect 30635 1270 30645 1290
rect 30665 1270 30675 1290
rect 30635 1240 30675 1270
rect 30635 1220 30645 1240
rect 30665 1220 30675 1240
rect 30635 1190 30675 1220
rect 30635 1170 30645 1190
rect 30665 1170 30675 1190
rect 30635 1140 30675 1170
rect 30635 1120 30645 1140
rect 30665 1120 30675 1140
rect 30635 1090 30675 1120
rect 30635 1070 30645 1090
rect 30665 1070 30675 1090
rect 30635 1040 30675 1070
rect 30635 1020 30645 1040
rect 30665 1020 30675 1040
rect 30635 990 30675 1020
rect 30635 970 30645 990
rect 30665 970 30675 990
rect 30635 955 30675 970
rect 31030 1695 31070 1710
rect 31030 1675 31040 1695
rect 31060 1675 31070 1695
rect 31030 1645 31070 1675
rect 31030 1625 31040 1645
rect 31060 1625 31070 1645
rect 31030 1595 31070 1625
rect 31030 1575 31040 1595
rect 31060 1575 31070 1595
rect 31030 1560 31070 1575
rect 31085 1695 31125 1710
rect 31085 1675 31095 1695
rect 31115 1675 31125 1695
rect 31085 1645 31125 1675
rect 31085 1625 31095 1645
rect 31115 1625 31125 1645
rect 31085 1595 31125 1625
rect 31085 1575 31095 1595
rect 31115 1575 31125 1595
rect 31085 1560 31125 1575
rect 31140 1695 31180 1710
rect 31140 1675 31150 1695
rect 31170 1675 31180 1695
rect 31140 1645 31180 1675
rect 31140 1625 31150 1645
rect 31170 1625 31180 1645
rect 31140 1595 31180 1625
rect 31140 1575 31150 1595
rect 31170 1575 31180 1595
rect 31140 1560 31180 1575
rect 31195 1695 31235 1710
rect 31195 1675 31205 1695
rect 31225 1675 31235 1695
rect 31195 1645 31235 1675
rect 31195 1625 31205 1645
rect 31225 1625 31235 1645
rect 31195 1595 31235 1625
rect 31195 1575 31205 1595
rect 31225 1575 31235 1595
rect 31195 1560 31235 1575
rect 31250 1695 31290 1710
rect 31250 1675 31260 1695
rect 31280 1675 31290 1695
rect 31250 1645 31290 1675
rect 31250 1625 31260 1645
rect 31280 1625 31290 1645
rect 31250 1595 31290 1625
rect 31250 1575 31260 1595
rect 31280 1575 31290 1595
rect 31250 1560 31290 1575
rect 31305 1695 31345 1710
rect 31305 1675 31315 1695
rect 31335 1675 31345 1695
rect 31305 1645 31345 1675
rect 31305 1625 31315 1645
rect 31335 1625 31345 1645
rect 31305 1595 31345 1625
rect 31305 1575 31315 1595
rect 31335 1575 31345 1595
rect 31305 1560 31345 1575
rect 31360 1695 31400 1710
rect 31360 1675 31370 1695
rect 31390 1675 31400 1695
rect 31360 1645 31400 1675
rect 31360 1625 31370 1645
rect 31390 1625 31400 1645
rect 31360 1595 31400 1625
rect 31360 1575 31370 1595
rect 31390 1575 31400 1595
rect 31360 1560 31400 1575
rect 31415 1695 31455 1710
rect 31415 1675 31425 1695
rect 31445 1675 31455 1695
rect 31415 1645 31455 1675
rect 31415 1625 31425 1645
rect 31445 1625 31455 1645
rect 31415 1595 31455 1625
rect 31415 1575 31425 1595
rect 31445 1575 31455 1595
rect 31415 1560 31455 1575
rect 31470 1695 31510 1710
rect 31470 1675 31480 1695
rect 31500 1675 31510 1695
rect 31470 1645 31510 1675
rect 31470 1625 31480 1645
rect 31500 1625 31510 1645
rect 31470 1595 31510 1625
rect 31470 1575 31480 1595
rect 31500 1575 31510 1595
rect 31470 1560 31510 1575
rect 31525 1695 31565 1710
rect 31525 1675 31535 1695
rect 31555 1675 31565 1695
rect 31525 1645 31565 1675
rect 31525 1625 31535 1645
rect 31555 1625 31565 1645
rect 31525 1595 31565 1625
rect 31525 1575 31535 1595
rect 31555 1575 31565 1595
rect 31525 1560 31565 1575
rect 31580 1695 31620 1710
rect 31580 1675 31590 1695
rect 31610 1675 31620 1695
rect 31580 1645 31620 1675
rect 31580 1625 31590 1645
rect 31610 1625 31620 1645
rect 31580 1595 31620 1625
rect 31580 1575 31590 1595
rect 31610 1575 31620 1595
rect 31580 1560 31620 1575
rect 31635 1695 31675 1710
rect 31635 1675 31645 1695
rect 31665 1675 31675 1695
rect 31635 1645 31675 1675
rect 31635 1625 31645 1645
rect 31665 1625 31675 1645
rect 31635 1595 31675 1625
rect 31635 1575 31645 1595
rect 31665 1575 31675 1595
rect 31635 1560 31675 1575
rect 31690 1695 31730 1710
rect 31690 1675 31700 1695
rect 31720 1675 31730 1695
rect 31690 1645 31730 1675
rect 31690 1625 31700 1645
rect 31720 1625 31730 1645
rect 31690 1595 31730 1625
rect 31690 1575 31700 1595
rect 31720 1575 31730 1595
rect 31690 1560 31730 1575
rect 31770 1695 31810 1710
rect 31770 1675 31780 1695
rect 31800 1675 31810 1695
rect 31770 1645 31810 1675
rect 31770 1625 31780 1645
rect 31800 1625 31810 1645
rect 31770 1595 31810 1625
rect 31770 1575 31780 1595
rect 31800 1575 31810 1595
rect 31770 1560 31810 1575
rect 31825 1695 31865 1710
rect 31825 1675 31835 1695
rect 31855 1675 31865 1695
rect 31825 1645 31865 1675
rect 31825 1625 31835 1645
rect 31855 1625 31865 1645
rect 31825 1595 31865 1625
rect 31825 1575 31835 1595
rect 31855 1575 31865 1595
rect 31825 1560 31865 1575
rect 31880 1695 31920 1710
rect 31880 1675 31890 1695
rect 31910 1675 31920 1695
rect 31880 1645 31920 1675
rect 31880 1625 31890 1645
rect 31910 1625 31920 1645
rect 31880 1595 31920 1625
rect 31880 1575 31890 1595
rect 31910 1575 31920 1595
rect 31880 1560 31920 1575
rect 31935 1695 31975 1710
rect 31935 1675 31945 1695
rect 31965 1675 31975 1695
rect 31935 1645 31975 1675
rect 31935 1625 31945 1645
rect 31965 1625 31975 1645
rect 31935 1595 31975 1625
rect 31935 1575 31945 1595
rect 31965 1575 31975 1595
rect 31935 1560 31975 1575
rect 31990 1695 32030 1710
rect 31990 1675 32000 1695
rect 32020 1675 32030 1695
rect 31990 1645 32030 1675
rect 31990 1625 32000 1645
rect 32020 1625 32030 1645
rect 31990 1595 32030 1625
rect 31990 1575 32000 1595
rect 32020 1575 32030 1595
rect 31990 1560 32030 1575
rect 32070 1695 32110 1710
rect 32070 1675 32080 1695
rect 32100 1675 32110 1695
rect 32070 1645 32110 1675
rect 32070 1625 32080 1645
rect 32100 1625 32110 1645
rect 32070 1595 32110 1625
rect 32070 1575 32080 1595
rect 32100 1575 32110 1595
rect 32070 1560 32110 1575
rect 32125 1695 32165 1710
rect 32125 1675 32135 1695
rect 32155 1675 32165 1695
rect 32125 1645 32165 1675
rect 32125 1625 32135 1645
rect 32155 1625 32165 1645
rect 32125 1595 32165 1625
rect 32125 1575 32135 1595
rect 32155 1575 32165 1595
rect 32125 1560 32165 1575
rect 32180 1695 32220 1710
rect 32180 1675 32190 1695
rect 32210 1675 32220 1695
rect 32180 1645 32220 1675
rect 32180 1625 32190 1645
rect 32210 1625 32220 1645
rect 32180 1595 32220 1625
rect 32180 1575 32190 1595
rect 32210 1575 32220 1595
rect 32180 1560 32220 1575
rect 32235 1695 32275 1710
rect 32235 1675 32245 1695
rect 32265 1675 32275 1695
rect 32235 1645 32275 1675
rect 32235 1625 32245 1645
rect 32265 1625 32275 1645
rect 32235 1595 32275 1625
rect 32235 1575 32245 1595
rect 32265 1575 32275 1595
rect 32235 1560 32275 1575
rect 32290 1695 32330 1710
rect 32290 1675 32300 1695
rect 32320 1675 32330 1695
rect 32290 1645 32330 1675
rect 32290 1625 32300 1645
rect 32320 1625 32330 1645
rect 32290 1595 32330 1625
rect 32290 1575 32300 1595
rect 32320 1575 32330 1595
rect 32290 1560 32330 1575
rect 32345 1695 32385 1710
rect 32345 1675 32355 1695
rect 32375 1675 32385 1695
rect 32345 1645 32385 1675
rect 32345 1625 32355 1645
rect 32375 1625 32385 1645
rect 32345 1595 32385 1625
rect 32345 1575 32355 1595
rect 32375 1575 32385 1595
rect 32345 1560 32385 1575
rect 32400 1695 32440 1710
rect 32400 1675 32410 1695
rect 32430 1675 32440 1695
rect 32400 1645 32440 1675
rect 32400 1625 32410 1645
rect 32430 1625 32440 1645
rect 32400 1595 32440 1625
rect 32400 1575 32410 1595
rect 32430 1575 32440 1595
rect 32400 1560 32440 1575
rect 32455 1695 32495 1710
rect 32455 1675 32465 1695
rect 32485 1675 32495 1695
rect 32455 1645 32495 1675
rect 32455 1625 32465 1645
rect 32485 1625 32495 1645
rect 32455 1595 32495 1625
rect 32455 1575 32465 1595
rect 32485 1575 32495 1595
rect 32455 1560 32495 1575
rect 32510 1695 32550 1710
rect 32510 1675 32520 1695
rect 32540 1675 32550 1695
rect 32510 1645 32550 1675
rect 32510 1625 32520 1645
rect 32540 1625 32550 1645
rect 32510 1595 32550 1625
rect 32510 1575 32520 1595
rect 32540 1575 32550 1595
rect 32510 1560 32550 1575
rect 32565 1695 32605 1710
rect 32565 1675 32575 1695
rect 32595 1675 32605 1695
rect 32565 1645 32605 1675
rect 32565 1625 32575 1645
rect 32595 1625 32605 1645
rect 32565 1595 32605 1625
rect 32565 1575 32575 1595
rect 32595 1575 32605 1595
rect 32565 1560 32605 1575
rect 32620 1695 32660 1710
rect 32620 1675 32630 1695
rect 32650 1675 32660 1695
rect 32620 1645 32660 1675
rect 32620 1625 32630 1645
rect 32650 1625 32660 1645
rect 32620 1595 32660 1625
rect 32620 1575 32630 1595
rect 32650 1575 32660 1595
rect 32620 1560 32660 1575
rect 32675 1695 32715 1710
rect 32675 1675 32685 1695
rect 32705 1675 32715 1695
rect 32675 1645 32715 1675
rect 32675 1625 32685 1645
rect 32705 1625 32715 1645
rect 32675 1595 32715 1625
rect 32675 1575 32685 1595
rect 32705 1575 32715 1595
rect 32675 1560 32715 1575
rect 32730 1695 32770 1710
rect 32730 1675 32740 1695
rect 32760 1675 32770 1695
rect 32730 1645 32770 1675
rect 32730 1625 32740 1645
rect 32760 1625 32770 1645
rect 32730 1595 32770 1625
rect 32730 1575 32740 1595
rect 32760 1575 32770 1595
rect 32730 1560 32770 1575
rect 31205 1190 31245 1205
rect 31205 1170 31215 1190
rect 31235 1170 31245 1190
rect 31205 1140 31245 1170
rect 31205 1120 31215 1140
rect 31235 1120 31245 1140
rect 31205 1090 31245 1120
rect 31205 1070 31215 1090
rect 31235 1070 31245 1090
rect 31205 1040 31245 1070
rect 31205 1020 31215 1040
rect 31235 1020 31245 1040
rect 31205 990 31245 1020
rect 31205 970 31215 990
rect 31235 970 31245 990
rect 31205 955 31245 970
rect 31260 1190 31300 1205
rect 31260 1170 31270 1190
rect 31290 1170 31300 1190
rect 31260 1140 31300 1170
rect 31260 1120 31270 1140
rect 31290 1120 31300 1140
rect 31260 1090 31300 1120
rect 31260 1070 31270 1090
rect 31290 1070 31300 1090
rect 31260 1040 31300 1070
rect 31260 1020 31270 1040
rect 31290 1020 31300 1040
rect 31260 990 31300 1020
rect 31260 970 31270 990
rect 31290 970 31300 990
rect 31260 955 31300 970
rect 31315 1190 31355 1205
rect 31315 1170 31325 1190
rect 31345 1170 31355 1190
rect 31315 1140 31355 1170
rect 31315 1120 31325 1140
rect 31345 1120 31355 1140
rect 31315 1090 31355 1120
rect 31315 1070 31325 1090
rect 31345 1070 31355 1090
rect 31315 1040 31355 1070
rect 31315 1020 31325 1040
rect 31345 1020 31355 1040
rect 31315 990 31355 1020
rect 31315 970 31325 990
rect 31345 970 31355 990
rect 31315 955 31355 970
rect 31370 1190 31410 1205
rect 31370 1170 31380 1190
rect 31400 1170 31410 1190
rect 31370 1140 31410 1170
rect 31370 1120 31380 1140
rect 31400 1120 31410 1140
rect 31370 1090 31410 1120
rect 31370 1070 31380 1090
rect 31400 1070 31410 1090
rect 31370 1040 31410 1070
rect 31370 1020 31380 1040
rect 31400 1020 31410 1040
rect 31370 990 31410 1020
rect 31370 970 31380 990
rect 31400 970 31410 990
rect 31370 955 31410 970
rect 31425 1190 31465 1205
rect 31425 1170 31435 1190
rect 31455 1170 31465 1190
rect 31425 1140 31465 1170
rect 31425 1120 31435 1140
rect 31455 1120 31465 1140
rect 31425 1090 31465 1120
rect 31425 1070 31435 1090
rect 31455 1070 31465 1090
rect 31425 1040 31465 1070
rect 31425 1020 31435 1040
rect 31455 1020 31465 1040
rect 31425 990 31465 1020
rect 31425 970 31435 990
rect 31455 970 31465 990
rect 31425 955 31465 970
rect 31480 1190 31520 1205
rect 31480 1170 31490 1190
rect 31510 1170 31520 1190
rect 31480 1140 31520 1170
rect 31480 1120 31490 1140
rect 31510 1120 31520 1140
rect 31480 1090 31520 1120
rect 31480 1070 31490 1090
rect 31510 1070 31520 1090
rect 31480 1040 31520 1070
rect 31480 1020 31490 1040
rect 31510 1020 31520 1040
rect 31480 990 31520 1020
rect 31480 970 31490 990
rect 31510 970 31520 990
rect 31480 955 31520 970
rect 31535 1190 31575 1205
rect 31535 1170 31545 1190
rect 31565 1170 31575 1190
rect 31535 1140 31575 1170
rect 31535 1120 31545 1140
rect 31565 1120 31575 1140
rect 31535 1090 31575 1120
rect 31535 1070 31545 1090
rect 31565 1070 31575 1090
rect 31535 1040 31575 1070
rect 31535 1020 31545 1040
rect 31565 1020 31575 1040
rect 31535 990 31575 1020
rect 31535 970 31545 990
rect 31565 970 31575 990
rect 31535 955 31575 970
rect 31590 1190 31630 1205
rect 31590 1170 31600 1190
rect 31620 1170 31630 1190
rect 31590 1140 31630 1170
rect 31590 1120 31600 1140
rect 31620 1120 31630 1140
rect 31590 1090 31630 1120
rect 31590 1070 31600 1090
rect 31620 1070 31630 1090
rect 31590 1040 31630 1070
rect 31590 1020 31600 1040
rect 31620 1020 31630 1040
rect 31590 990 31630 1020
rect 31590 970 31600 990
rect 31620 970 31630 990
rect 31590 955 31630 970
rect 31645 1190 31685 1205
rect 31645 1170 31655 1190
rect 31675 1170 31685 1190
rect 31645 1140 31685 1170
rect 31645 1120 31655 1140
rect 31675 1120 31685 1140
rect 31645 1090 31685 1120
rect 31645 1070 31655 1090
rect 31675 1070 31685 1090
rect 31645 1040 31685 1070
rect 31645 1020 31655 1040
rect 31675 1020 31685 1040
rect 31645 990 31685 1020
rect 31645 970 31655 990
rect 31675 970 31685 990
rect 31645 955 31685 970
rect 31700 1190 31740 1205
rect 31700 1170 31710 1190
rect 31730 1170 31740 1190
rect 31700 1140 31740 1170
rect 31700 1120 31710 1140
rect 31730 1120 31740 1140
rect 31700 1090 31740 1120
rect 31700 1070 31710 1090
rect 31730 1070 31740 1090
rect 31700 1040 31740 1070
rect 31700 1020 31710 1040
rect 31730 1020 31740 1040
rect 31700 990 31740 1020
rect 31700 970 31710 990
rect 31730 970 31740 990
rect 31700 955 31740 970
rect 31755 1190 31795 1205
rect 31755 1170 31765 1190
rect 31785 1170 31795 1190
rect 31755 1140 31795 1170
rect 31755 1120 31765 1140
rect 31785 1120 31795 1140
rect 31755 1090 31795 1120
rect 31755 1070 31765 1090
rect 31785 1070 31795 1090
rect 31755 1040 31795 1070
rect 31755 1020 31765 1040
rect 31785 1020 31795 1040
rect 31755 990 31795 1020
rect 31755 970 31765 990
rect 31785 970 31795 990
rect 31755 955 31795 970
rect 31810 1190 31850 1205
rect 31810 1170 31820 1190
rect 31840 1170 31850 1190
rect 31810 1140 31850 1170
rect 31810 1120 31820 1140
rect 31840 1120 31850 1140
rect 31810 1090 31850 1120
rect 31810 1070 31820 1090
rect 31840 1070 31850 1090
rect 31810 1040 31850 1070
rect 31810 1020 31820 1040
rect 31840 1020 31850 1040
rect 31810 990 31850 1020
rect 31810 970 31820 990
rect 31840 970 31850 990
rect 31810 955 31850 970
rect 31865 1190 31905 1205
rect 31865 1170 31875 1190
rect 31895 1170 31905 1190
rect 31865 1140 31905 1170
rect 31865 1120 31875 1140
rect 31895 1120 31905 1140
rect 31865 1090 31905 1120
rect 31865 1070 31875 1090
rect 31895 1070 31905 1090
rect 31865 1040 31905 1070
rect 31865 1020 31875 1040
rect 31895 1020 31905 1040
rect 31865 990 31905 1020
rect 31865 970 31875 990
rect 31895 970 31905 990
rect 31865 955 31905 970
rect 31920 1190 31960 1205
rect 31920 1170 31930 1190
rect 31950 1170 31960 1190
rect 31920 1140 31960 1170
rect 31920 1120 31930 1140
rect 31950 1120 31960 1140
rect 31920 1090 31960 1120
rect 31920 1070 31930 1090
rect 31950 1070 31960 1090
rect 31920 1040 31960 1070
rect 31920 1020 31930 1040
rect 31950 1020 31960 1040
rect 31920 990 31960 1020
rect 31920 970 31930 990
rect 31950 970 31960 990
rect 31920 955 31960 970
rect 31975 1190 32015 1205
rect 31975 1170 31985 1190
rect 32005 1170 32015 1190
rect 31975 1140 32015 1170
rect 31975 1120 31985 1140
rect 32005 1120 32015 1140
rect 31975 1090 32015 1120
rect 31975 1070 31985 1090
rect 32005 1070 32015 1090
rect 31975 1040 32015 1070
rect 31975 1020 31985 1040
rect 32005 1020 32015 1040
rect 31975 990 32015 1020
rect 31975 970 31985 990
rect 32005 970 32015 990
rect 31975 955 32015 970
rect 32030 1190 32070 1205
rect 32030 1170 32040 1190
rect 32060 1170 32070 1190
rect 32030 1140 32070 1170
rect 32030 1120 32040 1140
rect 32060 1120 32070 1140
rect 32030 1090 32070 1120
rect 32030 1070 32040 1090
rect 32060 1070 32070 1090
rect 32030 1040 32070 1070
rect 32030 1020 32040 1040
rect 32060 1020 32070 1040
rect 32030 990 32070 1020
rect 32030 970 32040 990
rect 32060 970 32070 990
rect 32030 955 32070 970
rect 32085 1190 32125 1205
rect 32085 1170 32095 1190
rect 32115 1170 32125 1190
rect 32085 1140 32125 1170
rect 32085 1120 32095 1140
rect 32115 1120 32125 1140
rect 32085 1090 32125 1120
rect 32085 1070 32095 1090
rect 32115 1070 32125 1090
rect 32085 1040 32125 1070
rect 32085 1020 32095 1040
rect 32115 1020 32125 1040
rect 32085 990 32125 1020
rect 32085 970 32095 990
rect 32115 970 32125 990
rect 32085 955 32125 970
rect 32140 1190 32180 1205
rect 32140 1170 32150 1190
rect 32170 1170 32180 1190
rect 32140 1140 32180 1170
rect 32140 1120 32150 1140
rect 32170 1120 32180 1140
rect 32140 1090 32180 1120
rect 32140 1070 32150 1090
rect 32170 1070 32180 1090
rect 32140 1040 32180 1070
rect 32140 1020 32150 1040
rect 32170 1020 32180 1040
rect 32140 990 32180 1020
rect 32140 970 32150 990
rect 32170 970 32180 990
rect 32140 955 32180 970
rect 32195 1190 32235 1205
rect 32195 1170 32205 1190
rect 32225 1170 32235 1190
rect 32195 1140 32235 1170
rect 32195 1120 32205 1140
rect 32225 1120 32235 1140
rect 32195 1090 32235 1120
rect 32195 1070 32205 1090
rect 32225 1070 32235 1090
rect 32195 1040 32235 1070
rect 32195 1020 32205 1040
rect 32225 1020 32235 1040
rect 32195 990 32235 1020
rect 32195 970 32205 990
rect 32225 970 32235 990
rect 32195 955 32235 970
rect 32250 1190 32290 1205
rect 32250 1170 32260 1190
rect 32280 1170 32290 1190
rect 32250 1140 32290 1170
rect 32250 1120 32260 1140
rect 32280 1120 32290 1140
rect 32250 1090 32290 1120
rect 32250 1070 32260 1090
rect 32280 1070 32290 1090
rect 32250 1040 32290 1070
rect 32250 1020 32260 1040
rect 32280 1020 32290 1040
rect 32250 990 32290 1020
rect 32250 970 32260 990
rect 32280 970 32290 990
rect 32250 955 32290 970
rect 32305 1190 32345 1205
rect 32305 1170 32315 1190
rect 32335 1170 32345 1190
rect 32305 1140 32345 1170
rect 32305 1120 32315 1140
rect 32335 1120 32345 1140
rect 32305 1090 32345 1120
rect 32305 1070 32315 1090
rect 32335 1070 32345 1090
rect 32305 1040 32345 1070
rect 32305 1020 32315 1040
rect 32335 1020 32345 1040
rect 32305 990 32345 1020
rect 32305 970 32315 990
rect 32335 970 32345 990
rect 32305 955 32345 970
rect 32360 1190 32400 1205
rect 32360 1170 32370 1190
rect 32390 1170 32400 1190
rect 32360 1140 32400 1170
rect 32360 1120 32370 1140
rect 32390 1120 32400 1140
rect 32360 1090 32400 1120
rect 32360 1070 32370 1090
rect 32390 1070 32400 1090
rect 32360 1040 32400 1070
rect 32360 1020 32370 1040
rect 32390 1020 32400 1040
rect 32360 990 32400 1020
rect 32360 970 32370 990
rect 32390 970 32400 990
rect 32360 955 32400 970
rect 32415 1190 32455 1205
rect 32415 1170 32425 1190
rect 32445 1170 32455 1190
rect 32415 1140 32455 1170
rect 32415 1120 32425 1140
rect 32445 1120 32455 1140
rect 32415 1090 32455 1120
rect 32415 1070 32425 1090
rect 32445 1070 32455 1090
rect 32415 1040 32455 1070
rect 32415 1020 32425 1040
rect 32445 1020 32455 1040
rect 32415 990 32455 1020
rect 32415 970 32425 990
rect 32445 970 32455 990
rect 32415 955 32455 970
rect 32470 1190 32510 1205
rect 32470 1170 32480 1190
rect 32500 1170 32510 1190
rect 32470 1140 32510 1170
rect 32470 1120 32480 1140
rect 32500 1120 32510 1140
rect 32470 1090 32510 1120
rect 32470 1070 32480 1090
rect 32500 1070 32510 1090
rect 32470 1040 32510 1070
rect 32470 1020 32480 1040
rect 32500 1020 32510 1040
rect 32470 990 32510 1020
rect 32470 970 32480 990
rect 32500 970 32510 990
rect 32470 955 32510 970
rect 33125 1640 33165 1655
rect 33125 1620 33135 1640
rect 33155 1620 33165 1640
rect 33125 1590 33165 1620
rect 33125 1570 33135 1590
rect 33155 1570 33165 1590
rect 33125 1540 33165 1570
rect 33125 1520 33135 1540
rect 33155 1520 33165 1540
rect 33125 1490 33165 1520
rect 33125 1470 33135 1490
rect 33155 1470 33165 1490
rect 33125 1440 33165 1470
rect 33125 1420 33135 1440
rect 33155 1420 33165 1440
rect 33125 1390 33165 1420
rect 33125 1370 33135 1390
rect 33155 1370 33165 1390
rect 33125 1340 33165 1370
rect 33125 1320 33135 1340
rect 33155 1320 33165 1340
rect 33125 1290 33165 1320
rect 33125 1270 33135 1290
rect 33155 1270 33165 1290
rect 33125 1240 33165 1270
rect 33125 1220 33135 1240
rect 33155 1220 33165 1240
rect 33125 1190 33165 1220
rect 33125 1170 33135 1190
rect 33155 1170 33165 1190
rect 33125 1140 33165 1170
rect 33125 1120 33135 1140
rect 33155 1120 33165 1140
rect 33125 1090 33165 1120
rect 33125 1070 33135 1090
rect 33155 1070 33165 1090
rect 33125 1040 33165 1070
rect 33125 1020 33135 1040
rect 33155 1020 33165 1040
rect 33125 990 33165 1020
rect 33125 970 33135 990
rect 33155 970 33165 990
rect 33125 955 33165 970
rect 33225 1640 33265 1655
rect 33225 1620 33235 1640
rect 33255 1620 33265 1640
rect 33225 1590 33265 1620
rect 33225 1570 33235 1590
rect 33255 1570 33265 1590
rect 33225 1540 33265 1570
rect 33225 1520 33235 1540
rect 33255 1520 33265 1540
rect 33225 1490 33265 1520
rect 33225 1470 33235 1490
rect 33255 1470 33265 1490
rect 33225 1440 33265 1470
rect 33225 1420 33235 1440
rect 33255 1420 33265 1440
rect 33225 1390 33265 1420
rect 33225 1370 33235 1390
rect 33255 1370 33265 1390
rect 33225 1340 33265 1370
rect 33225 1320 33235 1340
rect 33255 1320 33265 1340
rect 33225 1290 33265 1320
rect 33225 1270 33235 1290
rect 33255 1270 33265 1290
rect 33225 1240 33265 1270
rect 33225 1220 33235 1240
rect 33255 1220 33265 1240
rect 33225 1190 33265 1220
rect 33225 1170 33235 1190
rect 33255 1170 33265 1190
rect 33225 1140 33265 1170
rect 33225 1120 33235 1140
rect 33255 1120 33265 1140
rect 33225 1090 33265 1120
rect 33225 1070 33235 1090
rect 33255 1070 33265 1090
rect 33225 1040 33265 1070
rect 33225 1020 33235 1040
rect 33255 1020 33265 1040
rect 33225 990 33265 1020
rect 33225 970 33235 990
rect 33255 970 33265 990
rect 33225 955 33265 970
rect 33325 1640 33365 1655
rect 33325 1620 33335 1640
rect 33355 1620 33365 1640
rect 33325 1590 33365 1620
rect 33325 1570 33335 1590
rect 33355 1570 33365 1590
rect 33325 1540 33365 1570
rect 33325 1520 33335 1540
rect 33355 1520 33365 1540
rect 33325 1490 33365 1520
rect 33325 1470 33335 1490
rect 33355 1470 33365 1490
rect 33325 1440 33365 1470
rect 33325 1420 33335 1440
rect 33355 1420 33365 1440
rect 33325 1390 33365 1420
rect 33325 1370 33335 1390
rect 33355 1370 33365 1390
rect 33325 1340 33365 1370
rect 33325 1320 33335 1340
rect 33355 1320 33365 1340
rect 33325 1290 33365 1320
rect 33325 1270 33335 1290
rect 33355 1270 33365 1290
rect 33325 1240 33365 1270
rect 33325 1220 33335 1240
rect 33355 1220 33365 1240
rect 33325 1190 33365 1220
rect 33325 1170 33335 1190
rect 33355 1170 33365 1190
rect 33325 1140 33365 1170
rect 33325 1120 33335 1140
rect 33355 1120 33365 1140
rect 33325 1090 33365 1120
rect 33325 1070 33335 1090
rect 33355 1070 33365 1090
rect 33325 1040 33365 1070
rect 33325 1020 33335 1040
rect 33355 1020 33365 1040
rect 33325 990 33365 1020
rect 33325 970 33335 990
rect 33355 970 33365 990
rect 33325 955 33365 970
rect 33425 1640 33465 1655
rect 33425 1620 33435 1640
rect 33455 1620 33465 1640
rect 33425 1590 33465 1620
rect 33425 1570 33435 1590
rect 33455 1570 33465 1590
rect 33425 1540 33465 1570
rect 33425 1520 33435 1540
rect 33455 1520 33465 1540
rect 33425 1490 33465 1520
rect 33425 1470 33435 1490
rect 33455 1470 33465 1490
rect 33425 1440 33465 1470
rect 33425 1420 33435 1440
rect 33455 1420 33465 1440
rect 33425 1390 33465 1420
rect 33425 1370 33435 1390
rect 33455 1370 33465 1390
rect 33425 1340 33465 1370
rect 33425 1320 33435 1340
rect 33455 1320 33465 1340
rect 33425 1290 33465 1320
rect 33425 1270 33435 1290
rect 33455 1270 33465 1290
rect 33425 1240 33465 1270
rect 33425 1220 33435 1240
rect 33455 1220 33465 1240
rect 33425 1190 33465 1220
rect 33425 1170 33435 1190
rect 33455 1170 33465 1190
rect 33425 1140 33465 1170
rect 33425 1120 33435 1140
rect 33455 1120 33465 1140
rect 33425 1090 33465 1120
rect 33425 1070 33435 1090
rect 33455 1070 33465 1090
rect 33425 1040 33465 1070
rect 33425 1020 33435 1040
rect 33455 1020 33465 1040
rect 33425 990 33465 1020
rect 33425 970 33435 990
rect 33455 970 33465 990
rect 33425 955 33465 970
rect 33525 1640 33565 1655
rect 33525 1620 33535 1640
rect 33555 1620 33565 1640
rect 33525 1590 33565 1620
rect 33525 1570 33535 1590
rect 33555 1570 33565 1590
rect 33525 1540 33565 1570
rect 33525 1520 33535 1540
rect 33555 1520 33565 1540
rect 33525 1490 33565 1520
rect 33525 1470 33535 1490
rect 33555 1470 33565 1490
rect 33525 1440 33565 1470
rect 33525 1420 33535 1440
rect 33555 1420 33565 1440
rect 33525 1390 33565 1420
rect 33525 1370 33535 1390
rect 33555 1370 33565 1390
rect 33525 1340 33565 1370
rect 33525 1320 33535 1340
rect 33555 1320 33565 1340
rect 33525 1290 33565 1320
rect 33525 1270 33535 1290
rect 33555 1270 33565 1290
rect 33525 1240 33565 1270
rect 33525 1220 33535 1240
rect 33555 1220 33565 1240
rect 33525 1190 33565 1220
rect 33525 1170 33535 1190
rect 33555 1170 33565 1190
rect 33525 1140 33565 1170
rect 33525 1120 33535 1140
rect 33555 1120 33565 1140
rect 33525 1090 33565 1120
rect 33525 1070 33535 1090
rect 33555 1070 33565 1090
rect 33525 1040 33565 1070
rect 33525 1020 33535 1040
rect 33555 1020 33565 1040
rect 33525 990 33565 1020
rect 33525 970 33535 990
rect 33555 970 33565 990
rect 33525 955 33565 970
rect 33625 1640 33665 1655
rect 33625 1620 33635 1640
rect 33655 1620 33665 1640
rect 33625 1590 33665 1620
rect 33625 1570 33635 1590
rect 33655 1570 33665 1590
rect 33625 1540 33665 1570
rect 33625 1520 33635 1540
rect 33655 1520 33665 1540
rect 33625 1490 33665 1520
rect 33625 1470 33635 1490
rect 33655 1470 33665 1490
rect 33625 1440 33665 1470
rect 33625 1420 33635 1440
rect 33655 1420 33665 1440
rect 33625 1390 33665 1420
rect 33625 1370 33635 1390
rect 33655 1370 33665 1390
rect 33625 1340 33665 1370
rect 33625 1320 33635 1340
rect 33655 1320 33665 1340
rect 33625 1290 33665 1320
rect 33625 1270 33635 1290
rect 33655 1270 33665 1290
rect 33625 1240 33665 1270
rect 33625 1220 33635 1240
rect 33655 1220 33665 1240
rect 33625 1190 33665 1220
rect 33625 1170 33635 1190
rect 33655 1170 33665 1190
rect 33625 1140 33665 1170
rect 33625 1120 33635 1140
rect 33655 1120 33665 1140
rect 33625 1090 33665 1120
rect 33625 1070 33635 1090
rect 33655 1070 33665 1090
rect 33625 1040 33665 1070
rect 33625 1020 33635 1040
rect 33655 1020 33665 1040
rect 33625 990 33665 1020
rect 33625 970 33635 990
rect 33655 970 33665 990
rect 33625 955 33665 970
rect 33725 1640 33765 1655
rect 33725 1620 33735 1640
rect 33755 1620 33765 1640
rect 33725 1590 33765 1620
rect 33725 1570 33735 1590
rect 33755 1570 33765 1590
rect 33725 1540 33765 1570
rect 33725 1520 33735 1540
rect 33755 1520 33765 1540
rect 33725 1490 33765 1520
rect 33725 1470 33735 1490
rect 33755 1470 33765 1490
rect 33725 1440 33765 1470
rect 33725 1420 33735 1440
rect 33755 1420 33765 1440
rect 33725 1390 33765 1420
rect 33725 1370 33735 1390
rect 33755 1370 33765 1390
rect 33725 1340 33765 1370
rect 33725 1320 33735 1340
rect 33755 1320 33765 1340
rect 33725 1290 33765 1320
rect 33725 1270 33735 1290
rect 33755 1270 33765 1290
rect 33725 1240 33765 1270
rect 33725 1220 33735 1240
rect 33755 1220 33765 1240
rect 33725 1190 33765 1220
rect 33725 1170 33735 1190
rect 33755 1170 33765 1190
rect 33725 1140 33765 1170
rect 33725 1120 33735 1140
rect 33755 1120 33765 1140
rect 33725 1090 33765 1120
rect 33725 1070 33735 1090
rect 33755 1070 33765 1090
rect 33725 1040 33765 1070
rect 33725 1020 33735 1040
rect 33755 1020 33765 1040
rect 33725 990 33765 1020
rect 33725 970 33735 990
rect 33755 970 33765 990
rect 33725 955 33765 970
rect 31260 675 31300 690
rect 31260 655 31270 675
rect 31290 655 31300 675
rect 31260 625 31300 655
rect 31260 605 31270 625
rect 31290 605 31300 625
rect 31260 590 31300 605
rect 31490 675 31530 690
rect 31490 655 31500 675
rect 31520 655 31530 675
rect 31490 625 31530 655
rect 31490 605 31500 625
rect 31520 605 31530 625
rect 31490 590 31530 605
rect 31880 670 31920 685
rect 31880 650 31890 670
rect 31910 650 31920 670
rect 31880 635 31920 650
rect 31935 670 31975 685
rect 31935 650 31945 670
rect 31965 650 31975 670
rect 31935 635 31975 650
rect 31990 670 32030 685
rect 31990 650 32000 670
rect 32020 650 32030 670
rect 31990 635 32030 650
rect 32045 670 32085 685
rect 32045 650 32055 670
rect 32075 650 32085 670
rect 32045 635 32085 650
rect 32100 670 32140 685
rect 32100 650 32110 670
rect 32130 650 32140 670
rect 32100 635 32140 650
rect 32155 670 32195 685
rect 32155 650 32165 670
rect 32185 650 32195 670
rect 32155 635 32195 650
rect 32210 670 32250 685
rect 32210 650 32220 670
rect 32240 650 32250 670
rect 32210 635 32250 650
rect 32265 670 32305 685
rect 32265 650 32275 670
rect 32295 650 32305 670
rect 32265 635 32305 650
rect 32320 670 32360 685
rect 32320 650 32330 670
rect 32350 650 32360 670
rect 32320 635 32360 650
rect 32375 670 32415 685
rect 32375 650 32385 670
rect 32405 650 32415 670
rect 32375 635 32415 650
rect 32430 670 32470 685
rect 32430 650 32440 670
rect 32460 650 32470 670
rect 32430 635 32470 650
rect 32485 670 32525 685
rect 32485 650 32495 670
rect 32515 650 32525 670
rect 32485 635 32525 650
rect 32540 670 32580 685
rect 32540 650 32550 670
rect 32570 650 32580 670
rect 32540 635 32580 650
<< pdiff >>
rect 31220 4795 31260 4818
rect 31220 4775 31230 4795
rect 31250 4775 31260 4795
rect 31220 4755 31260 4775
rect 31280 4795 31320 4818
rect 31280 4775 31290 4795
rect 31310 4775 31320 4795
rect 31280 4755 31320 4775
rect 31340 4795 31380 4818
rect 31340 4775 31350 4795
rect 31370 4775 31380 4795
rect 31340 4755 31380 4775
rect 31400 4795 31440 4818
rect 31400 4775 31410 4795
rect 31430 4775 31440 4795
rect 31400 4755 31440 4775
rect 31470 4805 31510 4835
rect 31470 4785 31480 4805
rect 31500 4785 31510 4805
rect 31470 4755 31510 4785
rect 31530 4805 31570 4835
rect 31530 4785 31540 4805
rect 31560 4785 31570 4805
rect 31530 4755 31570 4785
rect 31590 4805 31630 4835
rect 31590 4785 31600 4805
rect 31620 4785 31630 4805
rect 31590 4755 31630 4785
rect 31650 4805 31690 4835
rect 31650 4785 31660 4805
rect 31680 4785 31690 4805
rect 31650 4755 31690 4785
rect 31710 4805 31750 4835
rect 31710 4785 31720 4805
rect 31740 4785 31750 4805
rect 31710 4755 31750 4785
rect 31770 4805 31810 4835
rect 31770 4785 31780 4805
rect 31800 4785 31810 4805
rect 31770 4755 31810 4785
rect 31830 4805 31870 4835
rect 31830 4785 31840 4805
rect 31860 4785 31870 4805
rect 31830 4755 31870 4785
rect 32200 4790 32240 4810
rect 32200 4770 32210 4790
rect 32230 4770 32240 4790
rect 32200 4750 32240 4770
rect 32260 4790 32300 4810
rect 32260 4770 32270 4790
rect 32290 4770 32300 4790
rect 32260 4750 32300 4770
rect 32320 4790 32360 4810
rect 32320 4770 32330 4790
rect 32350 4770 32360 4790
rect 32320 4750 32360 4770
rect 32380 4790 32420 4810
rect 32380 4770 32390 4790
rect 32410 4770 32420 4790
rect 32380 4750 32420 4770
rect 32440 4790 32480 4810
rect 32440 4770 32450 4790
rect 32470 4770 32480 4790
rect 32440 4750 32480 4770
rect 32500 4790 32540 4810
rect 32500 4770 32510 4790
rect 32530 4770 32540 4790
rect 32500 4750 32540 4770
rect 32560 4790 32600 4810
rect 32560 4770 32570 4790
rect 32590 4770 32600 4790
rect 32560 4750 32600 4770
rect 32620 4790 32660 4810
rect 32620 4770 32630 4790
rect 32650 4770 32660 4790
rect 32620 4750 32660 4770
rect 32680 4790 32720 4810
rect 32680 4770 32690 4790
rect 32710 4770 32720 4790
rect 32680 4750 32720 4770
rect 31250 4375 31290 4390
rect 31250 4355 31260 4375
rect 31280 4355 31290 4375
rect 31250 4340 31290 4355
rect 31305 4375 31345 4390
rect 31305 4355 31315 4375
rect 31335 4355 31345 4375
rect 31305 4340 31345 4355
rect 31360 4375 31400 4390
rect 31360 4355 31370 4375
rect 31390 4355 31400 4375
rect 31360 4340 31400 4355
rect 31415 4375 31455 4390
rect 31415 4355 31425 4375
rect 31445 4355 31455 4375
rect 31415 4340 31455 4355
rect 31470 4375 31510 4390
rect 31470 4355 31480 4375
rect 31500 4355 31510 4375
rect 31470 4340 31510 4355
rect 31525 4375 31565 4390
rect 31525 4355 31535 4375
rect 31555 4355 31565 4375
rect 31525 4340 31565 4355
rect 31580 4375 31620 4390
rect 31580 4355 31590 4375
rect 31610 4355 31620 4375
rect 31580 4340 31620 4355
rect 31635 4375 31675 4390
rect 31635 4355 31645 4375
rect 31665 4355 31675 4375
rect 31635 4340 31675 4355
rect 31690 4375 31730 4390
rect 31690 4355 31700 4375
rect 31720 4355 31730 4375
rect 31690 4340 31730 4355
rect 31745 4375 31785 4390
rect 31745 4355 31755 4375
rect 31775 4355 31785 4375
rect 31745 4340 31785 4355
rect 31800 4375 31840 4390
rect 31800 4355 31810 4375
rect 31830 4355 31840 4375
rect 31800 4340 31840 4355
rect 31855 4375 31895 4390
rect 31855 4355 31865 4375
rect 31885 4355 31895 4375
rect 31855 4340 31895 4355
rect 31910 4375 31950 4390
rect 31910 4355 31920 4375
rect 31940 4355 31950 4375
rect 31910 4340 31950 4355
rect 31965 4375 32005 4390
rect 31965 4355 31975 4375
rect 31995 4355 32005 4375
rect 31965 4340 32005 4355
rect 32020 4375 32060 4390
rect 32020 4355 32030 4375
rect 32050 4355 32060 4375
rect 32020 4340 32060 4355
rect 32075 4375 32115 4390
rect 32075 4355 32085 4375
rect 32105 4355 32115 4375
rect 32075 4340 32115 4355
rect 32130 4375 32170 4390
rect 32130 4355 32140 4375
rect 32160 4355 32170 4375
rect 32130 4340 32170 4355
rect 32185 4375 32225 4390
rect 32185 4355 32195 4375
rect 32215 4355 32225 4375
rect 32185 4340 32225 4355
rect 32240 4375 32280 4390
rect 32240 4355 32250 4375
rect 32270 4355 32280 4375
rect 32240 4340 32280 4355
rect 32295 4375 32335 4390
rect 32295 4355 32305 4375
rect 32325 4355 32335 4375
rect 32295 4340 32335 4355
rect 32350 4375 32390 4390
rect 32350 4355 32360 4375
rect 32380 4355 32390 4375
rect 32350 4340 32390 4355
rect 32405 4375 32445 4390
rect 32405 4355 32415 4375
rect 32435 4355 32445 4375
rect 32405 4340 32445 4355
rect 32460 4375 32500 4390
rect 32460 4355 32470 4375
rect 32490 4355 32500 4375
rect 32460 4340 32500 4355
rect 31200 3965 31240 3980
rect 31200 3945 31210 3965
rect 31230 3945 31240 3965
rect 31200 3930 31240 3945
rect 31255 3965 31295 3980
rect 31255 3945 31265 3965
rect 31285 3945 31295 3965
rect 31255 3930 31295 3945
rect 31310 3965 31350 3980
rect 31310 3945 31320 3965
rect 31340 3945 31350 3965
rect 31310 3930 31350 3945
rect 31365 3965 31405 3980
rect 31365 3945 31375 3965
rect 31395 3945 31405 3965
rect 31365 3930 31405 3945
rect 31420 3965 31460 3980
rect 31420 3945 31430 3965
rect 31450 3945 31460 3965
rect 31420 3930 31460 3945
rect 31475 3965 31515 3980
rect 31475 3945 31485 3965
rect 31505 3945 31515 3965
rect 31475 3930 31515 3945
rect 31530 3965 31570 3980
rect 31530 3945 31540 3965
rect 31560 3945 31570 3965
rect 31530 3930 31570 3945
rect 31585 3965 31625 3980
rect 31585 3945 31595 3965
rect 31615 3945 31625 3965
rect 31585 3930 31625 3945
rect 31640 3965 31680 3980
rect 31640 3945 31650 3965
rect 31670 3945 31680 3965
rect 31640 3930 31680 3945
rect 31695 3965 31735 3980
rect 31695 3945 31705 3965
rect 31725 3945 31735 3965
rect 31695 3930 31735 3945
rect 31750 3965 31790 3980
rect 31750 3945 31760 3965
rect 31780 3945 31790 3965
rect 31750 3930 31790 3945
rect 31805 3965 31845 3980
rect 31805 3945 31815 3965
rect 31835 3945 31845 3965
rect 31805 3930 31845 3945
rect 31860 3965 31900 3980
rect 31860 3945 31870 3965
rect 31890 3945 31900 3965
rect 31860 3930 31900 3945
rect 31930 3965 31970 3980
rect 31930 3945 31940 3965
rect 31960 3945 31970 3965
rect 31930 3930 31970 3945
rect 31985 3965 32025 3980
rect 31985 3945 31995 3965
rect 32015 3945 32025 3965
rect 31985 3930 32025 3945
rect 32040 3965 32080 3980
rect 32040 3945 32050 3965
rect 32070 3945 32080 3965
rect 32040 3930 32080 3945
rect 32095 3965 32135 3980
rect 32095 3945 32105 3965
rect 32125 3945 32135 3965
rect 32095 3930 32135 3945
rect 32150 3965 32190 3980
rect 32150 3945 32160 3965
rect 32180 3945 32190 3965
rect 32150 3930 32190 3945
rect 32205 3965 32245 3980
rect 32205 3945 32215 3965
rect 32235 3945 32245 3965
rect 32205 3930 32245 3945
rect 32260 3965 32300 3980
rect 32260 3945 32270 3965
rect 32290 3945 32300 3965
rect 32260 3930 32300 3945
rect 32315 3965 32355 3980
rect 32315 3945 32325 3965
rect 32345 3945 32355 3965
rect 32315 3930 32355 3945
rect 32370 3965 32410 3980
rect 32370 3945 32380 3965
rect 32400 3945 32410 3965
rect 32370 3930 32410 3945
rect 32425 3965 32465 3980
rect 32425 3945 32435 3965
rect 32455 3945 32465 3965
rect 32425 3930 32465 3945
rect 32480 3965 32520 3980
rect 32480 3945 32490 3965
rect 32510 3945 32520 3965
rect 32480 3930 32520 3945
rect 32535 3965 32575 3980
rect 32535 3945 32545 3965
rect 32565 3945 32575 3965
rect 32535 3930 32575 3945
rect 32590 3965 32630 3980
rect 32590 3945 32600 3965
rect 32620 3945 32630 3965
rect 32590 3930 32630 3945
rect 29955 3650 29995 3665
rect 29955 3630 29965 3650
rect 29985 3630 29995 3650
rect 29955 3600 29995 3630
rect 29955 3580 29965 3600
rect 29985 3580 29995 3600
rect 29955 3550 29995 3580
rect 29955 3530 29965 3550
rect 29985 3530 29995 3550
rect 29955 3500 29995 3530
rect 29955 3480 29965 3500
rect 29985 3480 29995 3500
rect 29955 3450 29995 3480
rect 29955 3430 29965 3450
rect 29985 3430 29995 3450
rect 29955 3400 29995 3430
rect 29955 3380 29965 3400
rect 29985 3380 29995 3400
rect 29955 3350 29995 3380
rect 29955 3330 29965 3350
rect 29985 3330 29995 3350
rect 29955 3300 29995 3330
rect 29955 3280 29965 3300
rect 29985 3280 29995 3300
rect 29955 3250 29995 3280
rect 29955 3230 29965 3250
rect 29985 3230 29995 3250
rect 29955 3200 29995 3230
rect 29955 3180 29965 3200
rect 29985 3180 29995 3200
rect 29955 3150 29995 3180
rect 29955 3130 29965 3150
rect 29985 3130 29995 3150
rect 29955 3100 29995 3130
rect 29955 3080 29965 3100
rect 29985 3080 29995 3100
rect 29955 3065 29995 3080
rect 30010 3650 30050 3665
rect 30010 3630 30020 3650
rect 30040 3630 30050 3650
rect 30010 3600 30050 3630
rect 30010 3580 30020 3600
rect 30040 3580 30050 3600
rect 30010 3550 30050 3580
rect 30010 3530 30020 3550
rect 30040 3530 30050 3550
rect 30010 3500 30050 3530
rect 30010 3480 30020 3500
rect 30040 3480 30050 3500
rect 30010 3450 30050 3480
rect 30010 3430 30020 3450
rect 30040 3430 30050 3450
rect 30010 3400 30050 3430
rect 30010 3380 30020 3400
rect 30040 3380 30050 3400
rect 30010 3350 30050 3380
rect 30010 3330 30020 3350
rect 30040 3330 30050 3350
rect 30010 3300 30050 3330
rect 30010 3280 30020 3300
rect 30040 3280 30050 3300
rect 30010 3250 30050 3280
rect 30010 3230 30020 3250
rect 30040 3230 30050 3250
rect 30010 3200 30050 3230
rect 30010 3180 30020 3200
rect 30040 3180 30050 3200
rect 30010 3150 30050 3180
rect 30010 3130 30020 3150
rect 30040 3130 30050 3150
rect 30010 3100 30050 3130
rect 30010 3080 30020 3100
rect 30040 3080 30050 3100
rect 30010 3065 30050 3080
rect 30065 3650 30105 3665
rect 30065 3630 30075 3650
rect 30095 3630 30105 3650
rect 30065 3600 30105 3630
rect 30065 3580 30075 3600
rect 30095 3580 30105 3600
rect 30065 3550 30105 3580
rect 30065 3530 30075 3550
rect 30095 3530 30105 3550
rect 30065 3500 30105 3530
rect 30065 3480 30075 3500
rect 30095 3480 30105 3500
rect 30065 3450 30105 3480
rect 30065 3430 30075 3450
rect 30095 3430 30105 3450
rect 30065 3400 30105 3430
rect 30065 3380 30075 3400
rect 30095 3380 30105 3400
rect 30065 3350 30105 3380
rect 30065 3330 30075 3350
rect 30095 3330 30105 3350
rect 30065 3300 30105 3330
rect 30065 3280 30075 3300
rect 30095 3280 30105 3300
rect 30065 3250 30105 3280
rect 30065 3230 30075 3250
rect 30095 3230 30105 3250
rect 30065 3200 30105 3230
rect 30065 3180 30075 3200
rect 30095 3180 30105 3200
rect 30065 3150 30105 3180
rect 30065 3130 30075 3150
rect 30095 3130 30105 3150
rect 30065 3100 30105 3130
rect 30065 3080 30075 3100
rect 30095 3080 30105 3100
rect 30065 3065 30105 3080
rect 30120 3650 30160 3665
rect 30120 3630 30130 3650
rect 30150 3630 30160 3650
rect 30120 3600 30160 3630
rect 30120 3580 30130 3600
rect 30150 3580 30160 3600
rect 30120 3550 30160 3580
rect 30120 3530 30130 3550
rect 30150 3530 30160 3550
rect 30120 3500 30160 3530
rect 30120 3480 30130 3500
rect 30150 3480 30160 3500
rect 30120 3450 30160 3480
rect 30120 3430 30130 3450
rect 30150 3430 30160 3450
rect 30120 3400 30160 3430
rect 30120 3380 30130 3400
rect 30150 3380 30160 3400
rect 30120 3350 30160 3380
rect 30120 3330 30130 3350
rect 30150 3330 30160 3350
rect 30120 3300 30160 3330
rect 30120 3280 30130 3300
rect 30150 3280 30160 3300
rect 30120 3250 30160 3280
rect 30120 3230 30130 3250
rect 30150 3230 30160 3250
rect 30120 3200 30160 3230
rect 30120 3180 30130 3200
rect 30150 3180 30160 3200
rect 30120 3150 30160 3180
rect 30120 3130 30130 3150
rect 30150 3130 30160 3150
rect 30120 3100 30160 3130
rect 30120 3080 30130 3100
rect 30150 3080 30160 3100
rect 30120 3065 30160 3080
rect 30175 3650 30215 3665
rect 30175 3630 30185 3650
rect 30205 3630 30215 3650
rect 30175 3600 30215 3630
rect 30175 3580 30185 3600
rect 30205 3580 30215 3600
rect 30175 3550 30215 3580
rect 30175 3530 30185 3550
rect 30205 3530 30215 3550
rect 30175 3500 30215 3530
rect 30175 3480 30185 3500
rect 30205 3480 30215 3500
rect 30175 3450 30215 3480
rect 30175 3430 30185 3450
rect 30205 3430 30215 3450
rect 30175 3400 30215 3430
rect 30175 3380 30185 3400
rect 30205 3380 30215 3400
rect 30175 3350 30215 3380
rect 30175 3330 30185 3350
rect 30205 3330 30215 3350
rect 30175 3300 30215 3330
rect 30175 3280 30185 3300
rect 30205 3280 30215 3300
rect 30175 3250 30215 3280
rect 30175 3230 30185 3250
rect 30205 3230 30215 3250
rect 30175 3200 30215 3230
rect 30175 3180 30185 3200
rect 30205 3180 30215 3200
rect 30175 3150 30215 3180
rect 30175 3130 30185 3150
rect 30205 3130 30215 3150
rect 30175 3100 30215 3130
rect 30175 3080 30185 3100
rect 30205 3080 30215 3100
rect 30175 3065 30215 3080
rect 30230 3650 30270 3665
rect 30230 3630 30240 3650
rect 30260 3630 30270 3650
rect 30230 3600 30270 3630
rect 30230 3580 30240 3600
rect 30260 3580 30270 3600
rect 30230 3550 30270 3580
rect 30230 3530 30240 3550
rect 30260 3530 30270 3550
rect 30230 3500 30270 3530
rect 30230 3480 30240 3500
rect 30260 3480 30270 3500
rect 30230 3450 30270 3480
rect 30230 3430 30240 3450
rect 30260 3430 30270 3450
rect 30230 3400 30270 3430
rect 30230 3380 30240 3400
rect 30260 3380 30270 3400
rect 30230 3350 30270 3380
rect 30230 3330 30240 3350
rect 30260 3330 30270 3350
rect 30230 3300 30270 3330
rect 30230 3280 30240 3300
rect 30260 3280 30270 3300
rect 30230 3250 30270 3280
rect 30230 3230 30240 3250
rect 30260 3230 30270 3250
rect 30230 3200 30270 3230
rect 30230 3180 30240 3200
rect 30260 3180 30270 3200
rect 30230 3150 30270 3180
rect 30230 3130 30240 3150
rect 30260 3130 30270 3150
rect 30230 3100 30270 3130
rect 30230 3080 30240 3100
rect 30260 3080 30270 3100
rect 30230 3065 30270 3080
rect 30285 3650 30325 3665
rect 30285 3630 30295 3650
rect 30315 3630 30325 3650
rect 30285 3600 30325 3630
rect 30285 3580 30295 3600
rect 30315 3580 30325 3600
rect 30285 3550 30325 3580
rect 30285 3530 30295 3550
rect 30315 3530 30325 3550
rect 30285 3500 30325 3530
rect 30285 3480 30295 3500
rect 30315 3480 30325 3500
rect 30285 3450 30325 3480
rect 30285 3430 30295 3450
rect 30315 3430 30325 3450
rect 30285 3400 30325 3430
rect 30285 3380 30295 3400
rect 30315 3380 30325 3400
rect 30285 3350 30325 3380
rect 30285 3330 30295 3350
rect 30315 3330 30325 3350
rect 30285 3300 30325 3330
rect 30285 3280 30295 3300
rect 30315 3280 30325 3300
rect 30285 3250 30325 3280
rect 30285 3230 30295 3250
rect 30315 3230 30325 3250
rect 30285 3200 30325 3230
rect 30285 3180 30295 3200
rect 30315 3180 30325 3200
rect 30285 3150 30325 3180
rect 30285 3130 30295 3150
rect 30315 3130 30325 3150
rect 30285 3100 30325 3130
rect 30285 3080 30295 3100
rect 30315 3080 30325 3100
rect 30285 3065 30325 3080
rect 30340 3650 30380 3665
rect 30340 3630 30350 3650
rect 30370 3630 30380 3650
rect 30340 3600 30380 3630
rect 30340 3580 30350 3600
rect 30370 3580 30380 3600
rect 30340 3550 30380 3580
rect 30340 3530 30350 3550
rect 30370 3530 30380 3550
rect 30340 3500 30380 3530
rect 30340 3480 30350 3500
rect 30370 3480 30380 3500
rect 30340 3450 30380 3480
rect 30340 3430 30350 3450
rect 30370 3430 30380 3450
rect 30340 3400 30380 3430
rect 30340 3380 30350 3400
rect 30370 3380 30380 3400
rect 30340 3350 30380 3380
rect 30340 3330 30350 3350
rect 30370 3330 30380 3350
rect 30340 3300 30380 3330
rect 30340 3280 30350 3300
rect 30370 3280 30380 3300
rect 30340 3250 30380 3280
rect 30340 3230 30350 3250
rect 30370 3230 30380 3250
rect 30340 3200 30380 3230
rect 30340 3180 30350 3200
rect 30370 3180 30380 3200
rect 30340 3150 30380 3180
rect 30340 3130 30350 3150
rect 30370 3130 30380 3150
rect 30340 3100 30380 3130
rect 30340 3080 30350 3100
rect 30370 3080 30380 3100
rect 30340 3065 30380 3080
rect 30395 3650 30435 3665
rect 30395 3630 30405 3650
rect 30425 3630 30435 3650
rect 30395 3600 30435 3630
rect 30395 3580 30405 3600
rect 30425 3580 30435 3600
rect 30395 3550 30435 3580
rect 30395 3530 30405 3550
rect 30425 3530 30435 3550
rect 30395 3500 30435 3530
rect 30395 3480 30405 3500
rect 30425 3480 30435 3500
rect 30395 3450 30435 3480
rect 30395 3430 30405 3450
rect 30425 3430 30435 3450
rect 30395 3400 30435 3430
rect 30395 3380 30405 3400
rect 30425 3380 30435 3400
rect 30395 3350 30435 3380
rect 30395 3330 30405 3350
rect 30425 3330 30435 3350
rect 30395 3300 30435 3330
rect 30395 3280 30405 3300
rect 30425 3280 30435 3300
rect 30395 3250 30435 3280
rect 30395 3230 30405 3250
rect 30425 3230 30435 3250
rect 30395 3200 30435 3230
rect 30395 3180 30405 3200
rect 30425 3180 30435 3200
rect 30395 3150 30435 3180
rect 30395 3130 30405 3150
rect 30425 3130 30435 3150
rect 30395 3100 30435 3130
rect 30395 3080 30405 3100
rect 30425 3080 30435 3100
rect 30395 3065 30435 3080
rect 30450 3650 30490 3665
rect 30450 3630 30460 3650
rect 30480 3630 30490 3650
rect 30450 3600 30490 3630
rect 30450 3580 30460 3600
rect 30480 3580 30490 3600
rect 30450 3550 30490 3580
rect 30450 3530 30460 3550
rect 30480 3530 30490 3550
rect 30450 3500 30490 3530
rect 30450 3480 30460 3500
rect 30480 3480 30490 3500
rect 30450 3450 30490 3480
rect 30450 3430 30460 3450
rect 30480 3430 30490 3450
rect 30450 3400 30490 3430
rect 30450 3380 30460 3400
rect 30480 3380 30490 3400
rect 30450 3350 30490 3380
rect 30450 3330 30460 3350
rect 30480 3330 30490 3350
rect 30450 3300 30490 3330
rect 30450 3280 30460 3300
rect 30480 3280 30490 3300
rect 30450 3250 30490 3280
rect 30450 3230 30460 3250
rect 30480 3230 30490 3250
rect 30450 3200 30490 3230
rect 30450 3180 30460 3200
rect 30480 3180 30490 3200
rect 30450 3150 30490 3180
rect 30450 3130 30460 3150
rect 30480 3130 30490 3150
rect 30450 3100 30490 3130
rect 30450 3080 30460 3100
rect 30480 3080 30490 3100
rect 30450 3065 30490 3080
rect 30505 3650 30545 3665
rect 30505 3630 30515 3650
rect 30535 3630 30545 3650
rect 30505 3600 30545 3630
rect 30505 3580 30515 3600
rect 30535 3580 30545 3600
rect 30505 3550 30545 3580
rect 30505 3530 30515 3550
rect 30535 3530 30545 3550
rect 30505 3500 30545 3530
rect 30505 3480 30515 3500
rect 30535 3480 30545 3500
rect 30505 3450 30545 3480
rect 30505 3430 30515 3450
rect 30535 3430 30545 3450
rect 30505 3400 30545 3430
rect 30505 3380 30515 3400
rect 30535 3380 30545 3400
rect 30505 3350 30545 3380
rect 30505 3330 30515 3350
rect 30535 3330 30545 3350
rect 30505 3300 30545 3330
rect 30505 3280 30515 3300
rect 30535 3280 30545 3300
rect 30505 3250 30545 3280
rect 30505 3230 30515 3250
rect 30535 3230 30545 3250
rect 30505 3200 30545 3230
rect 30505 3180 30515 3200
rect 30535 3180 30545 3200
rect 30505 3150 30545 3180
rect 30505 3130 30515 3150
rect 30535 3130 30545 3150
rect 30505 3100 30545 3130
rect 30505 3080 30515 3100
rect 30535 3080 30545 3100
rect 30505 3065 30545 3080
rect 30560 3650 30600 3665
rect 30560 3630 30570 3650
rect 30590 3630 30600 3650
rect 30560 3600 30600 3630
rect 30560 3580 30570 3600
rect 30590 3580 30600 3600
rect 30560 3550 30600 3580
rect 30560 3530 30570 3550
rect 30590 3530 30600 3550
rect 30560 3500 30600 3530
rect 30560 3480 30570 3500
rect 30590 3480 30600 3500
rect 30560 3450 30600 3480
rect 30560 3430 30570 3450
rect 30590 3430 30600 3450
rect 30560 3400 30600 3430
rect 30560 3380 30570 3400
rect 30590 3380 30600 3400
rect 30560 3350 30600 3380
rect 30560 3330 30570 3350
rect 30590 3330 30600 3350
rect 30560 3300 30600 3330
rect 30560 3280 30570 3300
rect 30590 3280 30600 3300
rect 30560 3250 30600 3280
rect 30560 3230 30570 3250
rect 30590 3230 30600 3250
rect 30560 3200 30600 3230
rect 30560 3180 30570 3200
rect 30590 3180 30600 3200
rect 30560 3150 30600 3180
rect 30560 3130 30570 3150
rect 30590 3130 30600 3150
rect 30560 3100 30600 3130
rect 30560 3080 30570 3100
rect 30590 3080 30600 3100
rect 30560 3065 30600 3080
rect 30615 3650 30655 3665
rect 30615 3630 30625 3650
rect 30645 3630 30655 3650
rect 30615 3600 30655 3630
rect 30615 3580 30625 3600
rect 30645 3580 30655 3600
rect 30615 3550 30655 3580
rect 30615 3530 30625 3550
rect 30645 3530 30655 3550
rect 30615 3500 30655 3530
rect 30615 3480 30625 3500
rect 30645 3480 30655 3500
rect 30615 3450 30655 3480
rect 30615 3430 30625 3450
rect 30645 3430 30655 3450
rect 30615 3400 30655 3430
rect 30615 3380 30625 3400
rect 30645 3380 30655 3400
rect 30615 3350 30655 3380
rect 30615 3330 30625 3350
rect 30645 3330 30655 3350
rect 30615 3300 30655 3330
rect 30615 3280 30625 3300
rect 30645 3280 30655 3300
rect 30615 3250 30655 3280
rect 30615 3230 30625 3250
rect 30645 3230 30655 3250
rect 30615 3200 30655 3230
rect 30615 3180 30625 3200
rect 30645 3180 30655 3200
rect 30615 3150 30655 3180
rect 30615 3130 30625 3150
rect 30645 3130 30655 3150
rect 30615 3100 30655 3130
rect 30615 3080 30625 3100
rect 30645 3080 30655 3100
rect 30615 3065 30655 3080
rect 31220 3540 31260 3555
rect 31220 3520 31230 3540
rect 31250 3520 31260 3540
rect 31220 3490 31260 3520
rect 31220 3470 31230 3490
rect 31250 3470 31260 3490
rect 31220 3440 31260 3470
rect 31220 3420 31230 3440
rect 31250 3420 31260 3440
rect 31220 3390 31260 3420
rect 31220 3370 31230 3390
rect 31250 3370 31260 3390
rect 31220 3340 31260 3370
rect 31220 3320 31230 3340
rect 31250 3320 31260 3340
rect 31220 3290 31260 3320
rect 31220 3270 31230 3290
rect 31250 3270 31260 3290
rect 31220 3240 31260 3270
rect 31220 3220 31230 3240
rect 31250 3220 31260 3240
rect 31220 3205 31260 3220
rect 31280 3540 31320 3555
rect 31280 3520 31290 3540
rect 31310 3520 31320 3540
rect 31280 3490 31320 3520
rect 31280 3470 31290 3490
rect 31310 3470 31320 3490
rect 31280 3440 31320 3470
rect 31280 3420 31290 3440
rect 31310 3420 31320 3440
rect 31280 3390 31320 3420
rect 31280 3370 31290 3390
rect 31310 3370 31320 3390
rect 31280 3340 31320 3370
rect 31280 3320 31290 3340
rect 31310 3320 31320 3340
rect 31280 3290 31320 3320
rect 31280 3270 31290 3290
rect 31310 3270 31320 3290
rect 31280 3240 31320 3270
rect 31280 3220 31290 3240
rect 31310 3220 31320 3240
rect 31280 3205 31320 3220
rect 31340 3540 31380 3555
rect 31340 3520 31350 3540
rect 31370 3520 31380 3540
rect 31340 3490 31380 3520
rect 31340 3470 31350 3490
rect 31370 3470 31380 3490
rect 31340 3440 31380 3470
rect 31340 3420 31350 3440
rect 31370 3420 31380 3440
rect 31340 3390 31380 3420
rect 31340 3370 31350 3390
rect 31370 3370 31380 3390
rect 31340 3340 31380 3370
rect 31340 3320 31350 3340
rect 31370 3320 31380 3340
rect 31340 3290 31380 3320
rect 31340 3270 31350 3290
rect 31370 3270 31380 3290
rect 31340 3240 31380 3270
rect 31340 3220 31350 3240
rect 31370 3220 31380 3240
rect 31340 3205 31380 3220
rect 31400 3540 31440 3555
rect 31400 3520 31410 3540
rect 31430 3520 31440 3540
rect 31400 3490 31440 3520
rect 31400 3470 31410 3490
rect 31430 3470 31440 3490
rect 31400 3440 31440 3470
rect 31400 3420 31410 3440
rect 31430 3420 31440 3440
rect 31400 3390 31440 3420
rect 31400 3370 31410 3390
rect 31430 3370 31440 3390
rect 31400 3340 31440 3370
rect 31400 3320 31410 3340
rect 31430 3320 31440 3340
rect 31400 3290 31440 3320
rect 31400 3270 31410 3290
rect 31430 3270 31440 3290
rect 31400 3240 31440 3270
rect 31400 3220 31410 3240
rect 31430 3220 31440 3240
rect 31400 3205 31440 3220
rect 31460 3540 31500 3555
rect 31460 3520 31470 3540
rect 31490 3520 31500 3540
rect 31460 3490 31500 3520
rect 31460 3470 31470 3490
rect 31490 3470 31500 3490
rect 31460 3440 31500 3470
rect 31460 3420 31470 3440
rect 31490 3420 31500 3440
rect 31460 3390 31500 3420
rect 31460 3370 31470 3390
rect 31490 3370 31500 3390
rect 31460 3340 31500 3370
rect 31460 3320 31470 3340
rect 31490 3320 31500 3340
rect 31460 3290 31500 3320
rect 31460 3270 31470 3290
rect 31490 3270 31500 3290
rect 31460 3240 31500 3270
rect 31460 3220 31470 3240
rect 31490 3220 31500 3240
rect 31460 3205 31500 3220
rect 31520 3540 31560 3555
rect 31520 3520 31530 3540
rect 31550 3520 31560 3540
rect 31520 3490 31560 3520
rect 31520 3470 31530 3490
rect 31550 3470 31560 3490
rect 31520 3440 31560 3470
rect 31520 3420 31530 3440
rect 31550 3420 31560 3440
rect 31520 3390 31560 3420
rect 31520 3370 31530 3390
rect 31550 3370 31560 3390
rect 31520 3340 31560 3370
rect 31520 3320 31530 3340
rect 31550 3320 31560 3340
rect 31520 3290 31560 3320
rect 31520 3270 31530 3290
rect 31550 3270 31560 3290
rect 31520 3240 31560 3270
rect 31520 3220 31530 3240
rect 31550 3220 31560 3240
rect 31520 3205 31560 3220
rect 31580 3540 31620 3555
rect 31580 3520 31590 3540
rect 31610 3520 31620 3540
rect 31580 3490 31620 3520
rect 31580 3470 31590 3490
rect 31610 3470 31620 3490
rect 31580 3440 31620 3470
rect 31580 3420 31590 3440
rect 31610 3420 31620 3440
rect 31580 3390 31620 3420
rect 31580 3370 31590 3390
rect 31610 3370 31620 3390
rect 31580 3340 31620 3370
rect 31580 3320 31590 3340
rect 31610 3320 31620 3340
rect 31580 3290 31620 3320
rect 31580 3270 31590 3290
rect 31610 3270 31620 3290
rect 31580 3240 31620 3270
rect 31580 3220 31590 3240
rect 31610 3220 31620 3240
rect 31580 3205 31620 3220
rect 31640 3540 31680 3555
rect 31640 3520 31650 3540
rect 31670 3520 31680 3540
rect 31640 3490 31680 3520
rect 31640 3470 31650 3490
rect 31670 3470 31680 3490
rect 31640 3440 31680 3470
rect 31640 3420 31650 3440
rect 31670 3420 31680 3440
rect 31640 3390 31680 3420
rect 31640 3370 31650 3390
rect 31670 3370 31680 3390
rect 31640 3340 31680 3370
rect 31640 3320 31650 3340
rect 31670 3320 31680 3340
rect 31640 3290 31680 3320
rect 31640 3270 31650 3290
rect 31670 3270 31680 3290
rect 31640 3240 31680 3270
rect 31640 3220 31650 3240
rect 31670 3220 31680 3240
rect 31640 3205 31680 3220
rect 31700 3540 31740 3555
rect 31700 3520 31710 3540
rect 31730 3520 31740 3540
rect 31700 3490 31740 3520
rect 31700 3470 31710 3490
rect 31730 3470 31740 3490
rect 31700 3440 31740 3470
rect 31700 3420 31710 3440
rect 31730 3420 31740 3440
rect 31700 3390 31740 3420
rect 31700 3370 31710 3390
rect 31730 3370 31740 3390
rect 31700 3340 31740 3370
rect 31700 3320 31710 3340
rect 31730 3320 31740 3340
rect 31700 3290 31740 3320
rect 31700 3270 31710 3290
rect 31730 3270 31740 3290
rect 31700 3240 31740 3270
rect 31700 3220 31710 3240
rect 31730 3220 31740 3240
rect 31700 3205 31740 3220
rect 31760 3540 31800 3555
rect 31760 3520 31770 3540
rect 31790 3520 31800 3540
rect 31760 3490 31800 3520
rect 31760 3470 31770 3490
rect 31790 3470 31800 3490
rect 31760 3440 31800 3470
rect 31760 3420 31770 3440
rect 31790 3420 31800 3440
rect 31760 3390 31800 3420
rect 31760 3370 31770 3390
rect 31790 3370 31800 3390
rect 31760 3340 31800 3370
rect 31760 3320 31770 3340
rect 31790 3320 31800 3340
rect 31760 3290 31800 3320
rect 31760 3270 31770 3290
rect 31790 3270 31800 3290
rect 31760 3240 31800 3270
rect 31760 3220 31770 3240
rect 31790 3220 31800 3240
rect 31760 3205 31800 3220
rect 31820 3540 31860 3555
rect 31820 3520 31830 3540
rect 31850 3520 31860 3540
rect 31820 3490 31860 3520
rect 31820 3470 31830 3490
rect 31850 3470 31860 3490
rect 31820 3440 31860 3470
rect 31820 3420 31830 3440
rect 31850 3420 31860 3440
rect 31820 3390 31860 3420
rect 31820 3370 31830 3390
rect 31850 3370 31860 3390
rect 31820 3340 31860 3370
rect 31820 3320 31830 3340
rect 31850 3320 31860 3340
rect 31820 3290 31860 3320
rect 31820 3270 31830 3290
rect 31850 3270 31860 3290
rect 31820 3240 31860 3270
rect 31820 3220 31830 3240
rect 31850 3220 31860 3240
rect 31820 3205 31860 3220
rect 31880 3540 31920 3555
rect 31880 3520 31890 3540
rect 31910 3520 31920 3540
rect 31880 3490 31920 3520
rect 31880 3470 31890 3490
rect 31910 3470 31920 3490
rect 31880 3440 31920 3470
rect 31880 3420 31890 3440
rect 31910 3420 31920 3440
rect 31880 3390 31920 3420
rect 31880 3370 31890 3390
rect 31910 3370 31920 3390
rect 31880 3340 31920 3370
rect 31880 3320 31890 3340
rect 31910 3320 31920 3340
rect 31880 3290 31920 3320
rect 31880 3270 31890 3290
rect 31910 3270 31920 3290
rect 31880 3240 31920 3270
rect 31880 3220 31890 3240
rect 31910 3220 31920 3240
rect 31880 3205 31920 3220
rect 31940 3540 31980 3555
rect 31940 3520 31950 3540
rect 31970 3520 31980 3540
rect 31940 3490 31980 3520
rect 31940 3470 31950 3490
rect 31970 3470 31980 3490
rect 31940 3440 31980 3470
rect 31940 3420 31950 3440
rect 31970 3420 31980 3440
rect 31940 3390 31980 3420
rect 31940 3370 31950 3390
rect 31970 3370 31980 3390
rect 31940 3340 31980 3370
rect 31940 3320 31950 3340
rect 31970 3320 31980 3340
rect 31940 3290 31980 3320
rect 31940 3270 31950 3290
rect 31970 3270 31980 3290
rect 31940 3240 31980 3270
rect 31940 3220 31950 3240
rect 31970 3220 31980 3240
rect 31940 3205 31980 3220
rect 32000 3540 32040 3555
rect 32000 3520 32010 3540
rect 32030 3520 32040 3540
rect 32000 3490 32040 3520
rect 32000 3470 32010 3490
rect 32030 3470 32040 3490
rect 32000 3440 32040 3470
rect 32000 3420 32010 3440
rect 32030 3420 32040 3440
rect 32000 3390 32040 3420
rect 32000 3370 32010 3390
rect 32030 3370 32040 3390
rect 32000 3340 32040 3370
rect 32000 3320 32010 3340
rect 32030 3320 32040 3340
rect 32000 3290 32040 3320
rect 32000 3270 32010 3290
rect 32030 3270 32040 3290
rect 32000 3240 32040 3270
rect 32000 3220 32010 3240
rect 32030 3220 32040 3240
rect 32000 3205 32040 3220
rect 32060 3540 32100 3555
rect 32060 3520 32070 3540
rect 32090 3520 32100 3540
rect 32060 3490 32100 3520
rect 32060 3470 32070 3490
rect 32090 3470 32100 3490
rect 32060 3440 32100 3470
rect 32060 3420 32070 3440
rect 32090 3420 32100 3440
rect 32060 3390 32100 3420
rect 32060 3370 32070 3390
rect 32090 3370 32100 3390
rect 32060 3340 32100 3370
rect 32060 3320 32070 3340
rect 32090 3320 32100 3340
rect 32060 3290 32100 3320
rect 32060 3270 32070 3290
rect 32090 3270 32100 3290
rect 32060 3240 32100 3270
rect 32060 3220 32070 3240
rect 32090 3220 32100 3240
rect 32060 3205 32100 3220
rect 32120 3540 32160 3555
rect 32120 3520 32130 3540
rect 32150 3520 32160 3540
rect 32120 3490 32160 3520
rect 32120 3470 32130 3490
rect 32150 3470 32160 3490
rect 32120 3440 32160 3470
rect 32120 3420 32130 3440
rect 32150 3420 32160 3440
rect 32120 3390 32160 3420
rect 32120 3370 32130 3390
rect 32150 3370 32160 3390
rect 32120 3340 32160 3370
rect 32120 3320 32130 3340
rect 32150 3320 32160 3340
rect 32120 3290 32160 3320
rect 32120 3270 32130 3290
rect 32150 3270 32160 3290
rect 32120 3240 32160 3270
rect 32120 3220 32130 3240
rect 32150 3220 32160 3240
rect 32120 3205 32160 3220
rect 32180 3540 32220 3555
rect 32180 3520 32190 3540
rect 32210 3520 32220 3540
rect 32180 3490 32220 3520
rect 32180 3470 32190 3490
rect 32210 3470 32220 3490
rect 32180 3440 32220 3470
rect 32180 3420 32190 3440
rect 32210 3420 32220 3440
rect 32180 3390 32220 3420
rect 32180 3370 32190 3390
rect 32210 3370 32220 3390
rect 32180 3340 32220 3370
rect 32180 3320 32190 3340
rect 32210 3320 32220 3340
rect 32180 3290 32220 3320
rect 32180 3270 32190 3290
rect 32210 3270 32220 3290
rect 32180 3240 32220 3270
rect 32180 3220 32190 3240
rect 32210 3220 32220 3240
rect 32180 3205 32220 3220
rect 32240 3540 32280 3555
rect 32240 3520 32250 3540
rect 32270 3520 32280 3540
rect 32240 3490 32280 3520
rect 32240 3470 32250 3490
rect 32270 3470 32280 3490
rect 32240 3440 32280 3470
rect 32240 3420 32250 3440
rect 32270 3420 32280 3440
rect 32240 3390 32280 3420
rect 32240 3370 32250 3390
rect 32270 3370 32280 3390
rect 32240 3340 32280 3370
rect 32240 3320 32250 3340
rect 32270 3320 32280 3340
rect 32240 3290 32280 3320
rect 32240 3270 32250 3290
rect 32270 3270 32280 3290
rect 32240 3240 32280 3270
rect 32240 3220 32250 3240
rect 32270 3220 32280 3240
rect 32240 3205 32280 3220
rect 32300 3540 32340 3555
rect 32300 3520 32310 3540
rect 32330 3520 32340 3540
rect 32300 3490 32340 3520
rect 32300 3470 32310 3490
rect 32330 3470 32340 3490
rect 32300 3440 32340 3470
rect 32300 3420 32310 3440
rect 32330 3420 32340 3440
rect 32300 3390 32340 3420
rect 32300 3370 32310 3390
rect 32330 3370 32340 3390
rect 32300 3340 32340 3370
rect 32300 3320 32310 3340
rect 32330 3320 32340 3340
rect 32300 3290 32340 3320
rect 32300 3270 32310 3290
rect 32330 3270 32340 3290
rect 32300 3240 32340 3270
rect 32300 3220 32310 3240
rect 32330 3220 32340 3240
rect 32300 3205 32340 3220
rect 32360 3540 32400 3555
rect 32360 3520 32370 3540
rect 32390 3520 32400 3540
rect 32360 3490 32400 3520
rect 32360 3470 32370 3490
rect 32390 3470 32400 3490
rect 32360 3440 32400 3470
rect 32360 3420 32370 3440
rect 32390 3420 32400 3440
rect 32360 3390 32400 3420
rect 32360 3370 32370 3390
rect 32390 3370 32400 3390
rect 32360 3340 32400 3370
rect 32360 3320 32370 3340
rect 32390 3320 32400 3340
rect 32360 3290 32400 3320
rect 32360 3270 32370 3290
rect 32390 3270 32400 3290
rect 32360 3240 32400 3270
rect 32360 3220 32370 3240
rect 32390 3220 32400 3240
rect 32360 3205 32400 3220
rect 32420 3540 32460 3555
rect 32420 3520 32430 3540
rect 32450 3520 32460 3540
rect 32420 3490 32460 3520
rect 32420 3470 32430 3490
rect 32450 3470 32460 3490
rect 32420 3440 32460 3470
rect 32420 3420 32430 3440
rect 32450 3420 32460 3440
rect 32420 3390 32460 3420
rect 32420 3370 32430 3390
rect 32450 3370 32460 3390
rect 32420 3340 32460 3370
rect 32420 3320 32430 3340
rect 32450 3320 32460 3340
rect 32420 3290 32460 3320
rect 32420 3270 32430 3290
rect 32450 3270 32460 3290
rect 32420 3240 32460 3270
rect 32420 3220 32430 3240
rect 32450 3220 32460 3240
rect 32420 3205 32460 3220
rect 32480 3540 32520 3555
rect 32480 3520 32490 3540
rect 32510 3520 32520 3540
rect 32480 3490 32520 3520
rect 32480 3470 32490 3490
rect 32510 3470 32520 3490
rect 32480 3440 32520 3470
rect 32480 3420 32490 3440
rect 32510 3420 32520 3440
rect 32480 3390 32520 3420
rect 32480 3370 32490 3390
rect 32510 3370 32520 3390
rect 32480 3340 32520 3370
rect 32480 3320 32490 3340
rect 32510 3320 32520 3340
rect 32480 3290 32520 3320
rect 32480 3270 32490 3290
rect 32510 3270 32520 3290
rect 32480 3240 32520 3270
rect 32480 3220 32490 3240
rect 32510 3220 32520 3240
rect 32480 3205 32520 3220
rect 32540 3540 32580 3555
rect 32540 3520 32550 3540
rect 32570 3520 32580 3540
rect 32540 3490 32580 3520
rect 32540 3470 32550 3490
rect 32570 3470 32580 3490
rect 32540 3440 32580 3470
rect 32540 3420 32550 3440
rect 32570 3420 32580 3440
rect 32540 3390 32580 3420
rect 32540 3370 32550 3390
rect 32570 3370 32580 3390
rect 32540 3340 32580 3370
rect 32540 3320 32550 3340
rect 32570 3320 32580 3340
rect 32540 3290 32580 3320
rect 32540 3270 32550 3290
rect 32570 3270 32580 3290
rect 32540 3240 32580 3270
rect 32540 3220 32550 3240
rect 32570 3220 32580 3240
rect 32540 3205 32580 3220
rect 33145 3650 33185 3665
rect 33145 3630 33155 3650
rect 33175 3630 33185 3650
rect 33145 3600 33185 3630
rect 33145 3580 33155 3600
rect 33175 3580 33185 3600
rect 33145 3550 33185 3580
rect 33145 3530 33155 3550
rect 33175 3530 33185 3550
rect 33145 3500 33185 3530
rect 33145 3480 33155 3500
rect 33175 3480 33185 3500
rect 33145 3450 33185 3480
rect 33145 3430 33155 3450
rect 33175 3430 33185 3450
rect 33145 3400 33185 3430
rect 33145 3380 33155 3400
rect 33175 3380 33185 3400
rect 33145 3350 33185 3380
rect 33145 3330 33155 3350
rect 33175 3330 33185 3350
rect 33145 3300 33185 3330
rect 33145 3280 33155 3300
rect 33175 3280 33185 3300
rect 33145 3250 33185 3280
rect 33145 3230 33155 3250
rect 33175 3230 33185 3250
rect 33145 3200 33185 3230
rect 33145 3180 33155 3200
rect 33175 3180 33185 3200
rect 33145 3150 33185 3180
rect 33145 3130 33155 3150
rect 33175 3130 33185 3150
rect 33145 3100 33185 3130
rect 33145 3080 33155 3100
rect 33175 3080 33185 3100
rect 33145 3065 33185 3080
rect 33200 3650 33240 3665
rect 33200 3630 33210 3650
rect 33230 3630 33240 3650
rect 33200 3600 33240 3630
rect 33200 3580 33210 3600
rect 33230 3580 33240 3600
rect 33200 3550 33240 3580
rect 33200 3530 33210 3550
rect 33230 3530 33240 3550
rect 33200 3500 33240 3530
rect 33200 3480 33210 3500
rect 33230 3480 33240 3500
rect 33200 3450 33240 3480
rect 33200 3430 33210 3450
rect 33230 3430 33240 3450
rect 33200 3400 33240 3430
rect 33200 3380 33210 3400
rect 33230 3380 33240 3400
rect 33200 3350 33240 3380
rect 33200 3330 33210 3350
rect 33230 3330 33240 3350
rect 33200 3300 33240 3330
rect 33200 3280 33210 3300
rect 33230 3280 33240 3300
rect 33200 3250 33240 3280
rect 33200 3230 33210 3250
rect 33230 3230 33240 3250
rect 33200 3200 33240 3230
rect 33200 3180 33210 3200
rect 33230 3180 33240 3200
rect 33200 3150 33240 3180
rect 33200 3130 33210 3150
rect 33230 3130 33240 3150
rect 33200 3100 33240 3130
rect 33200 3080 33210 3100
rect 33230 3080 33240 3100
rect 33200 3065 33240 3080
rect 33255 3650 33295 3665
rect 33255 3630 33265 3650
rect 33285 3630 33295 3650
rect 33255 3600 33295 3630
rect 33255 3580 33265 3600
rect 33285 3580 33295 3600
rect 33255 3550 33295 3580
rect 33255 3530 33265 3550
rect 33285 3530 33295 3550
rect 33255 3500 33295 3530
rect 33255 3480 33265 3500
rect 33285 3480 33295 3500
rect 33255 3450 33295 3480
rect 33255 3430 33265 3450
rect 33285 3430 33295 3450
rect 33255 3400 33295 3430
rect 33255 3380 33265 3400
rect 33285 3380 33295 3400
rect 33255 3350 33295 3380
rect 33255 3330 33265 3350
rect 33285 3330 33295 3350
rect 33255 3300 33295 3330
rect 33255 3280 33265 3300
rect 33285 3280 33295 3300
rect 33255 3250 33295 3280
rect 33255 3230 33265 3250
rect 33285 3230 33295 3250
rect 33255 3200 33295 3230
rect 33255 3180 33265 3200
rect 33285 3180 33295 3200
rect 33255 3150 33295 3180
rect 33255 3130 33265 3150
rect 33285 3130 33295 3150
rect 33255 3100 33295 3130
rect 33255 3080 33265 3100
rect 33285 3080 33295 3100
rect 33255 3065 33295 3080
rect 33310 3650 33350 3665
rect 33310 3630 33320 3650
rect 33340 3630 33350 3650
rect 33310 3600 33350 3630
rect 33310 3580 33320 3600
rect 33340 3580 33350 3600
rect 33310 3550 33350 3580
rect 33310 3530 33320 3550
rect 33340 3530 33350 3550
rect 33310 3500 33350 3530
rect 33310 3480 33320 3500
rect 33340 3480 33350 3500
rect 33310 3450 33350 3480
rect 33310 3430 33320 3450
rect 33340 3430 33350 3450
rect 33310 3400 33350 3430
rect 33310 3380 33320 3400
rect 33340 3380 33350 3400
rect 33310 3350 33350 3380
rect 33310 3330 33320 3350
rect 33340 3330 33350 3350
rect 33310 3300 33350 3330
rect 33310 3280 33320 3300
rect 33340 3280 33350 3300
rect 33310 3250 33350 3280
rect 33310 3230 33320 3250
rect 33340 3230 33350 3250
rect 33310 3200 33350 3230
rect 33310 3180 33320 3200
rect 33340 3180 33350 3200
rect 33310 3150 33350 3180
rect 33310 3130 33320 3150
rect 33340 3130 33350 3150
rect 33310 3100 33350 3130
rect 33310 3080 33320 3100
rect 33340 3080 33350 3100
rect 33310 3065 33350 3080
rect 33365 3650 33405 3665
rect 33365 3630 33375 3650
rect 33395 3630 33405 3650
rect 33365 3600 33405 3630
rect 33365 3580 33375 3600
rect 33395 3580 33405 3600
rect 33365 3550 33405 3580
rect 33365 3530 33375 3550
rect 33395 3530 33405 3550
rect 33365 3500 33405 3530
rect 33365 3480 33375 3500
rect 33395 3480 33405 3500
rect 33365 3450 33405 3480
rect 33365 3430 33375 3450
rect 33395 3430 33405 3450
rect 33365 3400 33405 3430
rect 33365 3380 33375 3400
rect 33395 3380 33405 3400
rect 33365 3350 33405 3380
rect 33365 3330 33375 3350
rect 33395 3330 33405 3350
rect 33365 3300 33405 3330
rect 33365 3280 33375 3300
rect 33395 3280 33405 3300
rect 33365 3250 33405 3280
rect 33365 3230 33375 3250
rect 33395 3230 33405 3250
rect 33365 3200 33405 3230
rect 33365 3180 33375 3200
rect 33395 3180 33405 3200
rect 33365 3150 33405 3180
rect 33365 3130 33375 3150
rect 33395 3130 33405 3150
rect 33365 3100 33405 3130
rect 33365 3080 33375 3100
rect 33395 3080 33405 3100
rect 33365 3065 33405 3080
rect 33420 3650 33460 3665
rect 33420 3630 33430 3650
rect 33450 3630 33460 3650
rect 33420 3600 33460 3630
rect 33420 3580 33430 3600
rect 33450 3580 33460 3600
rect 33420 3550 33460 3580
rect 33420 3530 33430 3550
rect 33450 3530 33460 3550
rect 33420 3500 33460 3530
rect 33420 3480 33430 3500
rect 33450 3480 33460 3500
rect 33420 3450 33460 3480
rect 33420 3430 33430 3450
rect 33450 3430 33460 3450
rect 33420 3400 33460 3430
rect 33420 3380 33430 3400
rect 33450 3380 33460 3400
rect 33420 3350 33460 3380
rect 33420 3330 33430 3350
rect 33450 3330 33460 3350
rect 33420 3300 33460 3330
rect 33420 3280 33430 3300
rect 33450 3280 33460 3300
rect 33420 3250 33460 3280
rect 33420 3230 33430 3250
rect 33450 3230 33460 3250
rect 33420 3200 33460 3230
rect 33420 3180 33430 3200
rect 33450 3180 33460 3200
rect 33420 3150 33460 3180
rect 33420 3130 33430 3150
rect 33450 3130 33460 3150
rect 33420 3100 33460 3130
rect 33420 3080 33430 3100
rect 33450 3080 33460 3100
rect 33420 3065 33460 3080
rect 33475 3650 33515 3665
rect 33475 3630 33485 3650
rect 33505 3630 33515 3650
rect 33475 3600 33515 3630
rect 33475 3580 33485 3600
rect 33505 3580 33515 3600
rect 33475 3550 33515 3580
rect 33475 3530 33485 3550
rect 33505 3530 33515 3550
rect 33475 3500 33515 3530
rect 33475 3480 33485 3500
rect 33505 3480 33515 3500
rect 33475 3450 33515 3480
rect 33475 3430 33485 3450
rect 33505 3430 33515 3450
rect 33475 3400 33515 3430
rect 33475 3380 33485 3400
rect 33505 3380 33515 3400
rect 33475 3350 33515 3380
rect 33475 3330 33485 3350
rect 33505 3330 33515 3350
rect 33475 3300 33515 3330
rect 33475 3280 33485 3300
rect 33505 3280 33515 3300
rect 33475 3250 33515 3280
rect 33475 3230 33485 3250
rect 33505 3230 33515 3250
rect 33475 3200 33515 3230
rect 33475 3180 33485 3200
rect 33505 3180 33515 3200
rect 33475 3150 33515 3180
rect 33475 3130 33485 3150
rect 33505 3130 33515 3150
rect 33475 3100 33515 3130
rect 33475 3080 33485 3100
rect 33505 3080 33515 3100
rect 33475 3065 33515 3080
rect 33530 3650 33570 3665
rect 33530 3630 33540 3650
rect 33560 3630 33570 3650
rect 33530 3600 33570 3630
rect 33530 3580 33540 3600
rect 33560 3580 33570 3600
rect 33530 3550 33570 3580
rect 33530 3530 33540 3550
rect 33560 3530 33570 3550
rect 33530 3500 33570 3530
rect 33530 3480 33540 3500
rect 33560 3480 33570 3500
rect 33530 3450 33570 3480
rect 33530 3430 33540 3450
rect 33560 3430 33570 3450
rect 33530 3400 33570 3430
rect 33530 3380 33540 3400
rect 33560 3380 33570 3400
rect 33530 3350 33570 3380
rect 33530 3330 33540 3350
rect 33560 3330 33570 3350
rect 33530 3300 33570 3330
rect 33530 3280 33540 3300
rect 33560 3280 33570 3300
rect 33530 3250 33570 3280
rect 33530 3230 33540 3250
rect 33560 3230 33570 3250
rect 33530 3200 33570 3230
rect 33530 3180 33540 3200
rect 33560 3180 33570 3200
rect 33530 3150 33570 3180
rect 33530 3130 33540 3150
rect 33560 3130 33570 3150
rect 33530 3100 33570 3130
rect 33530 3080 33540 3100
rect 33560 3080 33570 3100
rect 33530 3065 33570 3080
rect 33585 3650 33625 3665
rect 33585 3630 33595 3650
rect 33615 3630 33625 3650
rect 33585 3600 33625 3630
rect 33585 3580 33595 3600
rect 33615 3580 33625 3600
rect 33585 3550 33625 3580
rect 33585 3530 33595 3550
rect 33615 3530 33625 3550
rect 33585 3500 33625 3530
rect 33585 3480 33595 3500
rect 33615 3480 33625 3500
rect 33585 3450 33625 3480
rect 33585 3430 33595 3450
rect 33615 3430 33625 3450
rect 33585 3400 33625 3430
rect 33585 3380 33595 3400
rect 33615 3380 33625 3400
rect 33585 3350 33625 3380
rect 33585 3330 33595 3350
rect 33615 3330 33625 3350
rect 33585 3300 33625 3330
rect 33585 3280 33595 3300
rect 33615 3280 33625 3300
rect 33585 3250 33625 3280
rect 33585 3230 33595 3250
rect 33615 3230 33625 3250
rect 33585 3200 33625 3230
rect 33585 3180 33595 3200
rect 33615 3180 33625 3200
rect 33585 3150 33625 3180
rect 33585 3130 33595 3150
rect 33615 3130 33625 3150
rect 33585 3100 33625 3130
rect 33585 3080 33595 3100
rect 33615 3080 33625 3100
rect 33585 3065 33625 3080
rect 33640 3650 33680 3665
rect 33640 3630 33650 3650
rect 33670 3630 33680 3650
rect 33640 3600 33680 3630
rect 33640 3580 33650 3600
rect 33670 3580 33680 3600
rect 33640 3550 33680 3580
rect 33640 3530 33650 3550
rect 33670 3530 33680 3550
rect 33640 3500 33680 3530
rect 33640 3480 33650 3500
rect 33670 3480 33680 3500
rect 33640 3450 33680 3480
rect 33640 3430 33650 3450
rect 33670 3430 33680 3450
rect 33640 3400 33680 3430
rect 33640 3380 33650 3400
rect 33670 3380 33680 3400
rect 33640 3350 33680 3380
rect 33640 3330 33650 3350
rect 33670 3330 33680 3350
rect 33640 3300 33680 3330
rect 33640 3280 33650 3300
rect 33670 3280 33680 3300
rect 33640 3250 33680 3280
rect 33640 3230 33650 3250
rect 33670 3230 33680 3250
rect 33640 3200 33680 3230
rect 33640 3180 33650 3200
rect 33670 3180 33680 3200
rect 33640 3150 33680 3180
rect 33640 3130 33650 3150
rect 33670 3130 33680 3150
rect 33640 3100 33680 3130
rect 33640 3080 33650 3100
rect 33670 3080 33680 3100
rect 33640 3065 33680 3080
rect 33695 3650 33735 3665
rect 33695 3630 33705 3650
rect 33725 3630 33735 3650
rect 33695 3600 33735 3630
rect 33695 3580 33705 3600
rect 33725 3580 33735 3600
rect 33695 3550 33735 3580
rect 33695 3530 33705 3550
rect 33725 3530 33735 3550
rect 33695 3500 33735 3530
rect 33695 3480 33705 3500
rect 33725 3480 33735 3500
rect 33695 3450 33735 3480
rect 33695 3430 33705 3450
rect 33725 3430 33735 3450
rect 33695 3400 33735 3430
rect 33695 3380 33705 3400
rect 33725 3380 33735 3400
rect 33695 3350 33735 3380
rect 33695 3330 33705 3350
rect 33725 3330 33735 3350
rect 33695 3300 33735 3330
rect 33695 3280 33705 3300
rect 33725 3280 33735 3300
rect 33695 3250 33735 3280
rect 33695 3230 33705 3250
rect 33725 3230 33735 3250
rect 33695 3200 33735 3230
rect 33695 3180 33705 3200
rect 33725 3180 33735 3200
rect 33695 3150 33735 3180
rect 33695 3130 33705 3150
rect 33725 3130 33735 3150
rect 33695 3100 33735 3130
rect 33695 3080 33705 3100
rect 33725 3080 33735 3100
rect 33695 3065 33735 3080
rect 33750 3650 33790 3665
rect 33750 3630 33760 3650
rect 33780 3630 33790 3650
rect 33750 3600 33790 3630
rect 33750 3580 33760 3600
rect 33780 3580 33790 3600
rect 33750 3550 33790 3580
rect 33750 3530 33760 3550
rect 33780 3530 33790 3550
rect 33750 3500 33790 3530
rect 33750 3480 33760 3500
rect 33780 3480 33790 3500
rect 33750 3450 33790 3480
rect 33750 3430 33760 3450
rect 33780 3430 33790 3450
rect 33750 3400 33790 3430
rect 33750 3380 33760 3400
rect 33780 3380 33790 3400
rect 33750 3350 33790 3380
rect 33750 3330 33760 3350
rect 33780 3330 33790 3350
rect 33750 3300 33790 3330
rect 33750 3280 33760 3300
rect 33780 3280 33790 3300
rect 33750 3250 33790 3280
rect 33750 3230 33760 3250
rect 33780 3230 33790 3250
rect 33750 3200 33790 3230
rect 33750 3180 33760 3200
rect 33780 3180 33790 3200
rect 33750 3150 33790 3180
rect 33750 3130 33760 3150
rect 33780 3130 33790 3150
rect 33750 3100 33790 3130
rect 33750 3080 33760 3100
rect 33780 3080 33790 3100
rect 33750 3065 33790 3080
rect 33805 3650 33845 3665
rect 33805 3630 33815 3650
rect 33835 3630 33845 3650
rect 33805 3600 33845 3630
rect 33805 3580 33815 3600
rect 33835 3580 33845 3600
rect 33805 3550 33845 3580
rect 33805 3530 33815 3550
rect 33835 3530 33845 3550
rect 33805 3500 33845 3530
rect 33805 3480 33815 3500
rect 33835 3480 33845 3500
rect 33805 3450 33845 3480
rect 33805 3430 33815 3450
rect 33835 3430 33845 3450
rect 33805 3400 33845 3430
rect 33805 3380 33815 3400
rect 33835 3380 33845 3400
rect 33805 3350 33845 3380
rect 33805 3330 33815 3350
rect 33835 3330 33845 3350
rect 33805 3300 33845 3330
rect 33805 3280 33815 3300
rect 33835 3280 33845 3300
rect 33805 3250 33845 3280
rect 33805 3230 33815 3250
rect 33835 3230 33845 3250
rect 33805 3200 33845 3230
rect 33805 3180 33815 3200
rect 33835 3180 33845 3200
rect 33805 3150 33845 3180
rect 33805 3130 33815 3150
rect 33835 3130 33845 3150
rect 33805 3100 33845 3130
rect 33805 3080 33815 3100
rect 33835 3080 33845 3100
rect 33805 3065 33845 3080
rect 29955 2690 29995 2705
rect 29955 2670 29965 2690
rect 29985 2670 29995 2690
rect 29955 2640 29995 2670
rect 29955 2620 29965 2640
rect 29985 2620 29995 2640
rect 29955 2590 29995 2620
rect 29955 2570 29965 2590
rect 29985 2570 29995 2590
rect 29955 2540 29995 2570
rect 29955 2520 29965 2540
rect 29985 2520 29995 2540
rect 29955 2505 29995 2520
rect 30010 2690 30050 2705
rect 30010 2670 30020 2690
rect 30040 2670 30050 2690
rect 30010 2640 30050 2670
rect 30010 2620 30020 2640
rect 30040 2620 30050 2640
rect 30010 2590 30050 2620
rect 30010 2570 30020 2590
rect 30040 2570 30050 2590
rect 30010 2540 30050 2570
rect 30010 2520 30020 2540
rect 30040 2520 30050 2540
rect 30010 2505 30050 2520
rect 30065 2690 30105 2705
rect 30065 2670 30075 2690
rect 30095 2670 30105 2690
rect 30065 2640 30105 2670
rect 30065 2620 30075 2640
rect 30095 2620 30105 2640
rect 30065 2590 30105 2620
rect 30065 2570 30075 2590
rect 30095 2570 30105 2590
rect 30065 2540 30105 2570
rect 30065 2520 30075 2540
rect 30095 2520 30105 2540
rect 30065 2505 30105 2520
rect 30120 2690 30160 2705
rect 30120 2670 30130 2690
rect 30150 2670 30160 2690
rect 30120 2640 30160 2670
rect 30120 2620 30130 2640
rect 30150 2620 30160 2640
rect 30120 2590 30160 2620
rect 30120 2570 30130 2590
rect 30150 2570 30160 2590
rect 30120 2540 30160 2570
rect 30120 2520 30130 2540
rect 30150 2520 30160 2540
rect 30120 2505 30160 2520
rect 30175 2690 30215 2705
rect 30175 2670 30185 2690
rect 30205 2670 30215 2690
rect 30175 2640 30215 2670
rect 30175 2620 30185 2640
rect 30205 2620 30215 2640
rect 30175 2590 30215 2620
rect 30175 2570 30185 2590
rect 30205 2570 30215 2590
rect 30175 2540 30215 2570
rect 30175 2520 30185 2540
rect 30205 2520 30215 2540
rect 30175 2505 30215 2520
rect 30230 2690 30270 2705
rect 30230 2670 30240 2690
rect 30260 2670 30270 2690
rect 30230 2640 30270 2670
rect 30230 2620 30240 2640
rect 30260 2620 30270 2640
rect 30230 2590 30270 2620
rect 30230 2570 30240 2590
rect 30260 2570 30270 2590
rect 30230 2540 30270 2570
rect 30230 2520 30240 2540
rect 30260 2520 30270 2540
rect 30230 2505 30270 2520
rect 30285 2690 30325 2705
rect 30285 2670 30295 2690
rect 30315 2670 30325 2690
rect 30285 2640 30325 2670
rect 30285 2620 30295 2640
rect 30315 2620 30325 2640
rect 30285 2590 30325 2620
rect 30285 2570 30295 2590
rect 30315 2570 30325 2590
rect 30285 2540 30325 2570
rect 30285 2520 30295 2540
rect 30315 2520 30325 2540
rect 30285 2505 30325 2520
rect 30340 2690 30380 2705
rect 30340 2670 30350 2690
rect 30370 2670 30380 2690
rect 30340 2640 30380 2670
rect 30340 2620 30350 2640
rect 30370 2620 30380 2640
rect 30340 2590 30380 2620
rect 30340 2570 30350 2590
rect 30370 2570 30380 2590
rect 30340 2540 30380 2570
rect 30340 2520 30350 2540
rect 30370 2520 30380 2540
rect 30340 2505 30380 2520
rect 30395 2690 30435 2705
rect 30395 2670 30405 2690
rect 30425 2670 30435 2690
rect 30395 2640 30435 2670
rect 30395 2620 30405 2640
rect 30425 2620 30435 2640
rect 30395 2590 30435 2620
rect 30395 2570 30405 2590
rect 30425 2570 30435 2590
rect 30395 2540 30435 2570
rect 30395 2520 30405 2540
rect 30425 2520 30435 2540
rect 30395 2505 30435 2520
rect 30450 2690 30490 2705
rect 30450 2670 30460 2690
rect 30480 2670 30490 2690
rect 30450 2640 30490 2670
rect 30450 2620 30460 2640
rect 30480 2620 30490 2640
rect 30450 2590 30490 2620
rect 30450 2570 30460 2590
rect 30480 2570 30490 2590
rect 30450 2540 30490 2570
rect 30450 2520 30460 2540
rect 30480 2520 30490 2540
rect 30450 2505 30490 2520
rect 30505 2690 30545 2705
rect 30505 2670 30515 2690
rect 30535 2670 30545 2690
rect 30505 2640 30545 2670
rect 30505 2620 30515 2640
rect 30535 2620 30545 2640
rect 30505 2590 30545 2620
rect 30505 2570 30515 2590
rect 30535 2570 30545 2590
rect 30505 2540 30545 2570
rect 30505 2520 30515 2540
rect 30535 2520 30545 2540
rect 30505 2505 30545 2520
rect 30560 2690 30600 2705
rect 30560 2670 30570 2690
rect 30590 2670 30600 2690
rect 30560 2640 30600 2670
rect 30560 2620 30570 2640
rect 30590 2620 30600 2640
rect 30560 2590 30600 2620
rect 30560 2570 30570 2590
rect 30590 2570 30600 2590
rect 30560 2540 30600 2570
rect 30560 2520 30570 2540
rect 30590 2520 30600 2540
rect 30560 2505 30600 2520
rect 30615 2690 30655 2705
rect 30615 2670 30625 2690
rect 30645 2670 30655 2690
rect 30615 2640 30655 2670
rect 30615 2620 30625 2640
rect 30645 2620 30655 2640
rect 30615 2590 30655 2620
rect 30615 2570 30625 2590
rect 30645 2570 30655 2590
rect 30615 2540 30655 2570
rect 30615 2520 30625 2540
rect 30645 2520 30655 2540
rect 30615 2505 30655 2520
rect 31005 2830 31045 2845
rect 31005 2810 31015 2830
rect 31035 2810 31045 2830
rect 31005 2780 31045 2810
rect 31005 2760 31015 2780
rect 31035 2760 31045 2780
rect 31005 2730 31045 2760
rect 31005 2710 31015 2730
rect 31035 2710 31045 2730
rect 31005 2680 31045 2710
rect 31005 2660 31015 2680
rect 31035 2660 31045 2680
rect 31005 2630 31045 2660
rect 31005 2610 31015 2630
rect 31035 2610 31045 2630
rect 31005 2580 31045 2610
rect 31005 2560 31015 2580
rect 31035 2560 31045 2580
rect 31005 2530 31045 2560
rect 31005 2510 31015 2530
rect 31035 2510 31045 2530
rect 31005 2495 31045 2510
rect 31065 2830 31105 2845
rect 31065 2810 31075 2830
rect 31095 2810 31105 2830
rect 31065 2780 31105 2810
rect 31065 2760 31075 2780
rect 31095 2760 31105 2780
rect 31065 2730 31105 2760
rect 31065 2710 31075 2730
rect 31095 2710 31105 2730
rect 31065 2680 31105 2710
rect 31065 2660 31075 2680
rect 31095 2660 31105 2680
rect 31065 2630 31105 2660
rect 31065 2610 31075 2630
rect 31095 2610 31105 2630
rect 31065 2580 31105 2610
rect 31065 2560 31075 2580
rect 31095 2560 31105 2580
rect 31065 2530 31105 2560
rect 31065 2510 31075 2530
rect 31095 2510 31105 2530
rect 31065 2495 31105 2510
rect 31125 2830 31165 2845
rect 31125 2810 31135 2830
rect 31155 2810 31165 2830
rect 31125 2780 31165 2810
rect 31125 2760 31135 2780
rect 31155 2760 31165 2780
rect 31125 2730 31165 2760
rect 31125 2710 31135 2730
rect 31155 2710 31165 2730
rect 31125 2680 31165 2710
rect 31125 2660 31135 2680
rect 31155 2660 31165 2680
rect 31125 2630 31165 2660
rect 31125 2610 31135 2630
rect 31155 2610 31165 2630
rect 31125 2580 31165 2610
rect 31125 2560 31135 2580
rect 31155 2560 31165 2580
rect 31125 2530 31165 2560
rect 31125 2510 31135 2530
rect 31155 2510 31165 2530
rect 31125 2495 31165 2510
rect 31185 2830 31225 2845
rect 31185 2810 31195 2830
rect 31215 2810 31225 2830
rect 31185 2780 31225 2810
rect 31185 2760 31195 2780
rect 31215 2760 31225 2780
rect 31185 2730 31225 2760
rect 31185 2710 31195 2730
rect 31215 2710 31225 2730
rect 31185 2680 31225 2710
rect 31185 2660 31195 2680
rect 31215 2660 31225 2680
rect 31185 2630 31225 2660
rect 31185 2610 31195 2630
rect 31215 2610 31225 2630
rect 31185 2580 31225 2610
rect 31185 2560 31195 2580
rect 31215 2560 31225 2580
rect 31185 2530 31225 2560
rect 31185 2510 31195 2530
rect 31215 2510 31225 2530
rect 31185 2495 31225 2510
rect 31245 2830 31285 2845
rect 31245 2810 31255 2830
rect 31275 2810 31285 2830
rect 31245 2780 31285 2810
rect 31245 2760 31255 2780
rect 31275 2760 31285 2780
rect 31245 2730 31285 2760
rect 31245 2710 31255 2730
rect 31275 2710 31285 2730
rect 31245 2680 31285 2710
rect 31245 2660 31255 2680
rect 31275 2660 31285 2680
rect 31245 2630 31285 2660
rect 31245 2610 31255 2630
rect 31275 2610 31285 2630
rect 31245 2580 31285 2610
rect 31245 2560 31255 2580
rect 31275 2560 31285 2580
rect 31245 2530 31285 2560
rect 31245 2510 31255 2530
rect 31275 2510 31285 2530
rect 31245 2495 31285 2510
rect 31305 2830 31345 2845
rect 31305 2810 31315 2830
rect 31335 2810 31345 2830
rect 31305 2780 31345 2810
rect 31305 2760 31315 2780
rect 31335 2760 31345 2780
rect 31305 2730 31345 2760
rect 31305 2710 31315 2730
rect 31335 2710 31345 2730
rect 31305 2680 31345 2710
rect 31305 2660 31315 2680
rect 31335 2660 31345 2680
rect 31305 2630 31345 2660
rect 31305 2610 31315 2630
rect 31335 2610 31345 2630
rect 31305 2580 31345 2610
rect 31305 2560 31315 2580
rect 31335 2560 31345 2580
rect 31305 2530 31345 2560
rect 31305 2510 31315 2530
rect 31335 2510 31345 2530
rect 31305 2495 31345 2510
rect 31365 2830 31405 2845
rect 31365 2810 31375 2830
rect 31395 2810 31405 2830
rect 31365 2780 31405 2810
rect 31365 2760 31375 2780
rect 31395 2760 31405 2780
rect 31365 2730 31405 2760
rect 31365 2710 31375 2730
rect 31395 2710 31405 2730
rect 31365 2680 31405 2710
rect 31365 2660 31375 2680
rect 31395 2660 31405 2680
rect 31365 2630 31405 2660
rect 31365 2610 31375 2630
rect 31395 2610 31405 2630
rect 31365 2580 31405 2610
rect 31365 2560 31375 2580
rect 31395 2560 31405 2580
rect 31365 2530 31405 2560
rect 31365 2510 31375 2530
rect 31395 2510 31405 2530
rect 31365 2495 31405 2510
rect 31425 2830 31465 2845
rect 31425 2810 31435 2830
rect 31455 2810 31465 2830
rect 31425 2780 31465 2810
rect 31425 2760 31435 2780
rect 31455 2760 31465 2780
rect 31425 2730 31465 2760
rect 31425 2710 31435 2730
rect 31455 2710 31465 2730
rect 31425 2680 31465 2710
rect 31425 2660 31435 2680
rect 31455 2660 31465 2680
rect 31425 2630 31465 2660
rect 31425 2610 31435 2630
rect 31455 2610 31465 2630
rect 31425 2580 31465 2610
rect 31425 2560 31435 2580
rect 31455 2560 31465 2580
rect 31425 2530 31465 2560
rect 31425 2510 31435 2530
rect 31455 2510 31465 2530
rect 31425 2495 31465 2510
rect 31485 2830 31525 2845
rect 31485 2810 31495 2830
rect 31515 2810 31525 2830
rect 31485 2780 31525 2810
rect 31485 2760 31495 2780
rect 31515 2760 31525 2780
rect 31485 2730 31525 2760
rect 31485 2710 31495 2730
rect 31515 2710 31525 2730
rect 31485 2680 31525 2710
rect 31485 2660 31495 2680
rect 31515 2660 31525 2680
rect 31485 2630 31525 2660
rect 31485 2610 31495 2630
rect 31515 2610 31525 2630
rect 31485 2580 31525 2610
rect 31485 2560 31495 2580
rect 31515 2560 31525 2580
rect 31485 2530 31525 2560
rect 31485 2510 31495 2530
rect 31515 2510 31525 2530
rect 31485 2495 31525 2510
rect 31545 2830 31585 2845
rect 31545 2810 31555 2830
rect 31575 2810 31585 2830
rect 31545 2780 31585 2810
rect 31545 2760 31555 2780
rect 31575 2760 31585 2780
rect 31545 2730 31585 2760
rect 31545 2710 31555 2730
rect 31575 2710 31585 2730
rect 31545 2680 31585 2710
rect 31545 2660 31555 2680
rect 31575 2660 31585 2680
rect 31545 2630 31585 2660
rect 31545 2610 31555 2630
rect 31575 2610 31585 2630
rect 31545 2580 31585 2610
rect 31545 2560 31555 2580
rect 31575 2560 31585 2580
rect 31545 2530 31585 2560
rect 31545 2510 31555 2530
rect 31575 2510 31585 2530
rect 31545 2495 31585 2510
rect 31605 2830 31645 2845
rect 31605 2810 31615 2830
rect 31635 2810 31645 2830
rect 31605 2780 31645 2810
rect 31605 2760 31615 2780
rect 31635 2760 31645 2780
rect 31605 2730 31645 2760
rect 31605 2710 31615 2730
rect 31635 2710 31645 2730
rect 31605 2680 31645 2710
rect 31605 2660 31615 2680
rect 31635 2660 31645 2680
rect 31605 2630 31645 2660
rect 31605 2610 31615 2630
rect 31635 2610 31645 2630
rect 31605 2580 31645 2610
rect 31605 2560 31615 2580
rect 31635 2560 31645 2580
rect 31605 2530 31645 2560
rect 31605 2510 31615 2530
rect 31635 2510 31645 2530
rect 31605 2495 31645 2510
rect 31665 2830 31705 2845
rect 31665 2810 31675 2830
rect 31695 2810 31705 2830
rect 31665 2780 31705 2810
rect 31665 2760 31675 2780
rect 31695 2760 31705 2780
rect 31665 2730 31705 2760
rect 31665 2710 31675 2730
rect 31695 2710 31705 2730
rect 31665 2680 31705 2710
rect 31665 2660 31675 2680
rect 31695 2660 31705 2680
rect 31665 2630 31705 2660
rect 31665 2610 31675 2630
rect 31695 2610 31705 2630
rect 31665 2580 31705 2610
rect 31665 2560 31675 2580
rect 31695 2560 31705 2580
rect 31665 2530 31705 2560
rect 31665 2510 31675 2530
rect 31695 2510 31705 2530
rect 31665 2495 31705 2510
rect 31725 2830 31765 2845
rect 31725 2810 31735 2830
rect 31755 2810 31765 2830
rect 31725 2780 31765 2810
rect 31725 2760 31735 2780
rect 31755 2760 31765 2780
rect 31725 2730 31765 2760
rect 31725 2710 31735 2730
rect 31755 2710 31765 2730
rect 31725 2680 31765 2710
rect 31725 2660 31735 2680
rect 31755 2660 31765 2680
rect 31725 2630 31765 2660
rect 31725 2610 31735 2630
rect 31755 2610 31765 2630
rect 31725 2580 31765 2610
rect 31725 2560 31735 2580
rect 31755 2560 31765 2580
rect 31725 2530 31765 2560
rect 31725 2510 31735 2530
rect 31755 2510 31765 2530
rect 31725 2495 31765 2510
rect 32035 2830 32075 2845
rect 32035 2810 32045 2830
rect 32065 2810 32075 2830
rect 32035 2780 32075 2810
rect 32035 2760 32045 2780
rect 32065 2760 32075 2780
rect 32035 2730 32075 2760
rect 32035 2710 32045 2730
rect 32065 2710 32075 2730
rect 32035 2680 32075 2710
rect 32035 2660 32045 2680
rect 32065 2660 32075 2680
rect 32035 2630 32075 2660
rect 32035 2610 32045 2630
rect 32065 2610 32075 2630
rect 32035 2580 32075 2610
rect 32035 2560 32045 2580
rect 32065 2560 32075 2580
rect 32035 2530 32075 2560
rect 32035 2510 32045 2530
rect 32065 2510 32075 2530
rect 32035 2495 32075 2510
rect 32095 2830 32135 2845
rect 32095 2810 32105 2830
rect 32125 2810 32135 2830
rect 32095 2780 32135 2810
rect 32095 2760 32105 2780
rect 32125 2760 32135 2780
rect 32095 2730 32135 2760
rect 32095 2710 32105 2730
rect 32125 2710 32135 2730
rect 32095 2680 32135 2710
rect 32095 2660 32105 2680
rect 32125 2660 32135 2680
rect 32095 2630 32135 2660
rect 32095 2610 32105 2630
rect 32125 2610 32135 2630
rect 32095 2580 32135 2610
rect 32095 2560 32105 2580
rect 32125 2560 32135 2580
rect 32095 2530 32135 2560
rect 32095 2510 32105 2530
rect 32125 2510 32135 2530
rect 32095 2495 32135 2510
rect 32155 2830 32195 2845
rect 32155 2810 32165 2830
rect 32185 2810 32195 2830
rect 32155 2780 32195 2810
rect 32155 2760 32165 2780
rect 32185 2760 32195 2780
rect 32155 2730 32195 2760
rect 32155 2710 32165 2730
rect 32185 2710 32195 2730
rect 32155 2680 32195 2710
rect 32155 2660 32165 2680
rect 32185 2660 32195 2680
rect 32155 2630 32195 2660
rect 32155 2610 32165 2630
rect 32185 2610 32195 2630
rect 32155 2580 32195 2610
rect 32155 2560 32165 2580
rect 32185 2560 32195 2580
rect 32155 2530 32195 2560
rect 32155 2510 32165 2530
rect 32185 2510 32195 2530
rect 32155 2495 32195 2510
rect 32215 2830 32255 2845
rect 32215 2810 32225 2830
rect 32245 2810 32255 2830
rect 32215 2780 32255 2810
rect 32215 2760 32225 2780
rect 32245 2760 32255 2780
rect 32215 2730 32255 2760
rect 32215 2710 32225 2730
rect 32245 2710 32255 2730
rect 32215 2680 32255 2710
rect 32215 2660 32225 2680
rect 32245 2660 32255 2680
rect 32215 2630 32255 2660
rect 32215 2610 32225 2630
rect 32245 2610 32255 2630
rect 32215 2580 32255 2610
rect 32215 2560 32225 2580
rect 32245 2560 32255 2580
rect 32215 2530 32255 2560
rect 32215 2510 32225 2530
rect 32245 2510 32255 2530
rect 32215 2495 32255 2510
rect 32275 2830 32315 2845
rect 32275 2810 32285 2830
rect 32305 2810 32315 2830
rect 32275 2780 32315 2810
rect 32275 2760 32285 2780
rect 32305 2760 32315 2780
rect 32275 2730 32315 2760
rect 32275 2710 32285 2730
rect 32305 2710 32315 2730
rect 32275 2680 32315 2710
rect 32275 2660 32285 2680
rect 32305 2660 32315 2680
rect 32275 2630 32315 2660
rect 32275 2610 32285 2630
rect 32305 2610 32315 2630
rect 32275 2580 32315 2610
rect 32275 2560 32285 2580
rect 32305 2560 32315 2580
rect 32275 2530 32315 2560
rect 32275 2510 32285 2530
rect 32305 2510 32315 2530
rect 32275 2495 32315 2510
rect 32335 2830 32375 2845
rect 32335 2810 32345 2830
rect 32365 2810 32375 2830
rect 32335 2780 32375 2810
rect 32335 2760 32345 2780
rect 32365 2760 32375 2780
rect 32335 2730 32375 2760
rect 32335 2710 32345 2730
rect 32365 2710 32375 2730
rect 32335 2680 32375 2710
rect 32335 2660 32345 2680
rect 32365 2660 32375 2680
rect 32335 2630 32375 2660
rect 32335 2610 32345 2630
rect 32365 2610 32375 2630
rect 32335 2580 32375 2610
rect 32335 2560 32345 2580
rect 32365 2560 32375 2580
rect 32335 2530 32375 2560
rect 32335 2510 32345 2530
rect 32365 2510 32375 2530
rect 32335 2495 32375 2510
rect 32395 2830 32435 2845
rect 32395 2810 32405 2830
rect 32425 2810 32435 2830
rect 32395 2780 32435 2810
rect 32395 2760 32405 2780
rect 32425 2760 32435 2780
rect 32395 2730 32435 2760
rect 32395 2710 32405 2730
rect 32425 2710 32435 2730
rect 32395 2680 32435 2710
rect 32395 2660 32405 2680
rect 32425 2660 32435 2680
rect 32395 2630 32435 2660
rect 32395 2610 32405 2630
rect 32425 2610 32435 2630
rect 32395 2580 32435 2610
rect 32395 2560 32405 2580
rect 32425 2560 32435 2580
rect 32395 2530 32435 2560
rect 32395 2510 32405 2530
rect 32425 2510 32435 2530
rect 32395 2495 32435 2510
rect 32455 2830 32495 2845
rect 32455 2810 32465 2830
rect 32485 2810 32495 2830
rect 32455 2780 32495 2810
rect 32455 2760 32465 2780
rect 32485 2760 32495 2780
rect 32455 2730 32495 2760
rect 32455 2710 32465 2730
rect 32485 2710 32495 2730
rect 32455 2680 32495 2710
rect 32455 2660 32465 2680
rect 32485 2660 32495 2680
rect 32455 2630 32495 2660
rect 32455 2610 32465 2630
rect 32485 2610 32495 2630
rect 32455 2580 32495 2610
rect 32455 2560 32465 2580
rect 32485 2560 32495 2580
rect 32455 2530 32495 2560
rect 32455 2510 32465 2530
rect 32485 2510 32495 2530
rect 32455 2495 32495 2510
rect 32515 2830 32555 2845
rect 32515 2810 32525 2830
rect 32545 2810 32555 2830
rect 32515 2780 32555 2810
rect 32515 2760 32525 2780
rect 32545 2760 32555 2780
rect 32515 2730 32555 2760
rect 32515 2710 32525 2730
rect 32545 2710 32555 2730
rect 32515 2680 32555 2710
rect 32515 2660 32525 2680
rect 32545 2660 32555 2680
rect 32515 2630 32555 2660
rect 32515 2610 32525 2630
rect 32545 2610 32555 2630
rect 32515 2580 32555 2610
rect 32515 2560 32525 2580
rect 32545 2560 32555 2580
rect 32515 2530 32555 2560
rect 32515 2510 32525 2530
rect 32545 2510 32555 2530
rect 32515 2495 32555 2510
rect 32575 2830 32615 2845
rect 32575 2810 32585 2830
rect 32605 2810 32615 2830
rect 32575 2780 32615 2810
rect 32575 2760 32585 2780
rect 32605 2760 32615 2780
rect 32575 2730 32615 2760
rect 32575 2710 32585 2730
rect 32605 2710 32615 2730
rect 32575 2680 32615 2710
rect 32575 2660 32585 2680
rect 32605 2660 32615 2680
rect 32575 2630 32615 2660
rect 32575 2610 32585 2630
rect 32605 2610 32615 2630
rect 32575 2580 32615 2610
rect 32575 2560 32585 2580
rect 32605 2560 32615 2580
rect 32575 2530 32615 2560
rect 32575 2510 32585 2530
rect 32605 2510 32615 2530
rect 32575 2495 32615 2510
rect 32635 2830 32675 2845
rect 32635 2810 32645 2830
rect 32665 2810 32675 2830
rect 32635 2780 32675 2810
rect 32635 2760 32645 2780
rect 32665 2760 32675 2780
rect 32635 2730 32675 2760
rect 32635 2710 32645 2730
rect 32665 2710 32675 2730
rect 32635 2680 32675 2710
rect 32635 2660 32645 2680
rect 32665 2660 32675 2680
rect 32635 2630 32675 2660
rect 32635 2610 32645 2630
rect 32665 2610 32675 2630
rect 32635 2580 32675 2610
rect 32635 2560 32645 2580
rect 32665 2560 32675 2580
rect 32635 2530 32675 2560
rect 32635 2510 32645 2530
rect 32665 2510 32675 2530
rect 32635 2495 32675 2510
rect 32695 2830 32735 2845
rect 32695 2810 32705 2830
rect 32725 2810 32735 2830
rect 32695 2780 32735 2810
rect 32695 2760 32705 2780
rect 32725 2760 32735 2780
rect 32695 2730 32735 2760
rect 32695 2710 32705 2730
rect 32725 2710 32735 2730
rect 32695 2680 32735 2710
rect 32695 2660 32705 2680
rect 32725 2660 32735 2680
rect 32695 2630 32735 2660
rect 32695 2610 32705 2630
rect 32725 2610 32735 2630
rect 32695 2580 32735 2610
rect 32695 2560 32705 2580
rect 32725 2560 32735 2580
rect 32695 2530 32735 2560
rect 32695 2510 32705 2530
rect 32725 2510 32735 2530
rect 32695 2495 32735 2510
rect 32755 2830 32795 2845
rect 32755 2810 32765 2830
rect 32785 2810 32795 2830
rect 32755 2780 32795 2810
rect 32755 2760 32765 2780
rect 32785 2760 32795 2780
rect 32755 2730 32795 2760
rect 32755 2710 32765 2730
rect 32785 2710 32795 2730
rect 32755 2680 32795 2710
rect 32755 2660 32765 2680
rect 32785 2660 32795 2680
rect 32755 2630 32795 2660
rect 32755 2610 32765 2630
rect 32785 2610 32795 2630
rect 32755 2580 32795 2610
rect 32755 2560 32765 2580
rect 32785 2560 32795 2580
rect 32755 2530 32795 2560
rect 32755 2510 32765 2530
rect 32785 2510 32795 2530
rect 32755 2495 32795 2510
rect 33145 2690 33185 2705
rect 33145 2670 33155 2690
rect 33175 2670 33185 2690
rect 33145 2640 33185 2670
rect 33145 2620 33155 2640
rect 33175 2620 33185 2640
rect 33145 2590 33185 2620
rect 33145 2570 33155 2590
rect 33175 2570 33185 2590
rect 33145 2540 33185 2570
rect 33145 2520 33155 2540
rect 33175 2520 33185 2540
rect 33145 2505 33185 2520
rect 33200 2690 33240 2705
rect 33200 2670 33210 2690
rect 33230 2670 33240 2690
rect 33200 2640 33240 2670
rect 33200 2620 33210 2640
rect 33230 2620 33240 2640
rect 33200 2590 33240 2620
rect 33200 2570 33210 2590
rect 33230 2570 33240 2590
rect 33200 2540 33240 2570
rect 33200 2520 33210 2540
rect 33230 2520 33240 2540
rect 33200 2505 33240 2520
rect 33255 2690 33295 2705
rect 33255 2670 33265 2690
rect 33285 2670 33295 2690
rect 33255 2640 33295 2670
rect 33255 2620 33265 2640
rect 33285 2620 33295 2640
rect 33255 2590 33295 2620
rect 33255 2570 33265 2590
rect 33285 2570 33295 2590
rect 33255 2540 33295 2570
rect 33255 2520 33265 2540
rect 33285 2520 33295 2540
rect 33255 2505 33295 2520
rect 33310 2690 33350 2705
rect 33310 2670 33320 2690
rect 33340 2670 33350 2690
rect 33310 2640 33350 2670
rect 33310 2620 33320 2640
rect 33340 2620 33350 2640
rect 33310 2590 33350 2620
rect 33310 2570 33320 2590
rect 33340 2570 33350 2590
rect 33310 2540 33350 2570
rect 33310 2520 33320 2540
rect 33340 2520 33350 2540
rect 33310 2505 33350 2520
rect 33365 2690 33405 2705
rect 33365 2670 33375 2690
rect 33395 2670 33405 2690
rect 33365 2640 33405 2670
rect 33365 2620 33375 2640
rect 33395 2620 33405 2640
rect 33365 2590 33405 2620
rect 33365 2570 33375 2590
rect 33395 2570 33405 2590
rect 33365 2540 33405 2570
rect 33365 2520 33375 2540
rect 33395 2520 33405 2540
rect 33365 2505 33405 2520
rect 33420 2690 33460 2705
rect 33420 2670 33430 2690
rect 33450 2670 33460 2690
rect 33420 2640 33460 2670
rect 33420 2620 33430 2640
rect 33450 2620 33460 2640
rect 33420 2590 33460 2620
rect 33420 2570 33430 2590
rect 33450 2570 33460 2590
rect 33420 2540 33460 2570
rect 33420 2520 33430 2540
rect 33450 2520 33460 2540
rect 33420 2505 33460 2520
rect 33475 2690 33515 2705
rect 33475 2670 33485 2690
rect 33505 2670 33515 2690
rect 33475 2640 33515 2670
rect 33475 2620 33485 2640
rect 33505 2620 33515 2640
rect 33475 2590 33515 2620
rect 33475 2570 33485 2590
rect 33505 2570 33515 2590
rect 33475 2540 33515 2570
rect 33475 2520 33485 2540
rect 33505 2520 33515 2540
rect 33475 2505 33515 2520
rect 33530 2690 33570 2705
rect 33530 2670 33540 2690
rect 33560 2670 33570 2690
rect 33530 2640 33570 2670
rect 33530 2620 33540 2640
rect 33560 2620 33570 2640
rect 33530 2590 33570 2620
rect 33530 2570 33540 2590
rect 33560 2570 33570 2590
rect 33530 2540 33570 2570
rect 33530 2520 33540 2540
rect 33560 2520 33570 2540
rect 33530 2505 33570 2520
rect 33585 2690 33625 2705
rect 33585 2670 33595 2690
rect 33615 2670 33625 2690
rect 33585 2640 33625 2670
rect 33585 2620 33595 2640
rect 33615 2620 33625 2640
rect 33585 2590 33625 2620
rect 33585 2570 33595 2590
rect 33615 2570 33625 2590
rect 33585 2540 33625 2570
rect 33585 2520 33595 2540
rect 33615 2520 33625 2540
rect 33585 2505 33625 2520
rect 33640 2690 33680 2705
rect 33640 2670 33650 2690
rect 33670 2670 33680 2690
rect 33640 2640 33680 2670
rect 33640 2620 33650 2640
rect 33670 2620 33680 2640
rect 33640 2590 33680 2620
rect 33640 2570 33650 2590
rect 33670 2570 33680 2590
rect 33640 2540 33680 2570
rect 33640 2520 33650 2540
rect 33670 2520 33680 2540
rect 33640 2505 33680 2520
rect 33695 2690 33735 2705
rect 33695 2670 33705 2690
rect 33725 2670 33735 2690
rect 33695 2640 33735 2670
rect 33695 2620 33705 2640
rect 33725 2620 33735 2640
rect 33695 2590 33735 2620
rect 33695 2570 33705 2590
rect 33725 2570 33735 2590
rect 33695 2540 33735 2570
rect 33695 2520 33705 2540
rect 33725 2520 33735 2540
rect 33695 2505 33735 2520
rect 33750 2690 33790 2705
rect 33750 2670 33760 2690
rect 33780 2670 33790 2690
rect 33750 2640 33790 2670
rect 33750 2620 33760 2640
rect 33780 2620 33790 2640
rect 33750 2590 33790 2620
rect 33750 2570 33760 2590
rect 33780 2570 33790 2590
rect 33750 2540 33790 2570
rect 33750 2520 33760 2540
rect 33780 2520 33790 2540
rect 33750 2505 33790 2520
rect 33805 2690 33845 2705
rect 33805 2670 33815 2690
rect 33835 2670 33845 2690
rect 33805 2640 33845 2670
rect 33805 2620 33815 2640
rect 33835 2620 33845 2640
rect 33805 2590 33845 2620
rect 33805 2570 33815 2590
rect 33835 2570 33845 2590
rect 33805 2540 33845 2570
rect 33805 2520 33815 2540
rect 33835 2520 33845 2540
rect 33805 2505 33845 2520
<< ndiffc >>
rect 29965 2210 29985 2230
rect 29965 2160 29985 2180
rect 29965 2110 29985 2130
rect 29965 2060 29985 2080
rect 29965 2010 29985 2030
rect 29965 1960 29985 1980
rect 30020 2210 30040 2230
rect 30020 2160 30040 2180
rect 30020 2110 30040 2130
rect 30020 2060 30040 2080
rect 30020 2010 30040 2030
rect 30020 1960 30040 1980
rect 30075 2210 30095 2230
rect 30075 2160 30095 2180
rect 30075 2110 30095 2130
rect 30075 2060 30095 2080
rect 30075 2010 30095 2030
rect 30075 1960 30095 1980
rect 30130 2210 30150 2230
rect 30130 2160 30150 2180
rect 30130 2110 30150 2130
rect 30130 2060 30150 2080
rect 30130 2010 30150 2030
rect 30130 1960 30150 1980
rect 30185 2210 30205 2230
rect 30185 2160 30205 2180
rect 30185 2110 30205 2130
rect 30185 2060 30205 2080
rect 30185 2010 30205 2030
rect 30185 1960 30205 1980
rect 30240 2210 30260 2230
rect 30240 2160 30260 2180
rect 30240 2110 30260 2130
rect 30240 2060 30260 2080
rect 30240 2010 30260 2030
rect 30240 1960 30260 1980
rect 30295 2210 30315 2230
rect 30295 2160 30315 2180
rect 30295 2110 30315 2130
rect 30295 2060 30315 2080
rect 30295 2010 30315 2030
rect 30295 1960 30315 1980
rect 30350 2210 30370 2230
rect 30350 2160 30370 2180
rect 30350 2110 30370 2130
rect 30350 2060 30370 2080
rect 30350 2010 30370 2030
rect 30350 1960 30370 1980
rect 30405 2210 30425 2230
rect 30405 2160 30425 2180
rect 30405 2110 30425 2130
rect 30405 2060 30425 2080
rect 30405 2010 30425 2030
rect 30405 1960 30425 1980
rect 30460 2210 30480 2230
rect 30460 2160 30480 2180
rect 30460 2110 30480 2130
rect 30460 2060 30480 2080
rect 30460 2010 30480 2030
rect 30460 1960 30480 1980
rect 30515 2210 30535 2230
rect 30515 2160 30535 2180
rect 30515 2110 30535 2130
rect 30515 2060 30535 2080
rect 30515 2010 30535 2030
rect 30515 1960 30535 1980
rect 30570 2210 30590 2230
rect 30570 2160 30590 2180
rect 30570 2110 30590 2130
rect 30570 2060 30590 2080
rect 30570 2010 30590 2030
rect 30570 1960 30590 1980
rect 30625 2210 30645 2230
rect 30625 2160 30645 2180
rect 30625 2110 30645 2130
rect 30625 2060 30645 2080
rect 30625 2010 30645 2030
rect 30625 1960 30645 1980
rect 31195 2145 31215 2165
rect 31195 2095 31215 2115
rect 31195 2045 31215 2065
rect 31250 2145 31270 2165
rect 31250 2095 31270 2115
rect 31250 2045 31270 2065
rect 31305 2145 31325 2165
rect 31305 2095 31325 2115
rect 31305 2045 31325 2065
rect 31360 2145 31380 2165
rect 31360 2095 31380 2115
rect 31360 2045 31380 2065
rect 31415 2145 31435 2165
rect 31415 2095 31435 2115
rect 31415 2045 31435 2065
rect 31470 2145 31490 2165
rect 31470 2095 31490 2115
rect 31470 2045 31490 2065
rect 31525 2145 31545 2165
rect 31525 2095 31545 2115
rect 31525 2045 31545 2065
rect 31580 2145 31600 2165
rect 31580 2095 31600 2115
rect 31580 2045 31600 2065
rect 31635 2145 31655 2165
rect 31635 2095 31655 2115
rect 31635 2045 31655 2065
rect 31690 2145 31710 2165
rect 31690 2095 31710 2115
rect 31690 2045 31710 2065
rect 31745 2145 31765 2165
rect 31745 2095 31765 2115
rect 31745 2045 31765 2065
rect 31800 2145 31820 2165
rect 31800 2095 31820 2115
rect 31800 2045 31820 2065
rect 31855 2145 31875 2165
rect 31855 2095 31875 2115
rect 31855 2045 31875 2065
rect 31925 2145 31945 2165
rect 31925 2095 31945 2115
rect 31925 2045 31945 2065
rect 31980 2145 32000 2165
rect 31980 2095 32000 2115
rect 31980 2045 32000 2065
rect 32035 2145 32055 2165
rect 32035 2095 32055 2115
rect 32035 2045 32055 2065
rect 32090 2145 32110 2165
rect 32090 2095 32110 2115
rect 32090 2045 32110 2065
rect 32145 2145 32165 2165
rect 32145 2095 32165 2115
rect 32145 2045 32165 2065
rect 32200 2145 32220 2165
rect 32200 2095 32220 2115
rect 32200 2045 32220 2065
rect 32255 2145 32275 2165
rect 32255 2095 32275 2115
rect 32255 2045 32275 2065
rect 32310 2145 32330 2165
rect 32310 2095 32330 2115
rect 32310 2045 32330 2065
rect 32365 2145 32385 2165
rect 32365 2095 32385 2115
rect 32365 2045 32385 2065
rect 32420 2145 32440 2165
rect 32420 2095 32440 2115
rect 32420 2045 32440 2065
rect 32475 2145 32495 2165
rect 32475 2095 32495 2115
rect 32475 2045 32495 2065
rect 32530 2145 32550 2165
rect 32530 2095 32550 2115
rect 32530 2045 32550 2065
rect 32585 2145 32605 2165
rect 32585 2095 32605 2115
rect 32585 2045 32605 2065
rect 33155 2210 33175 2230
rect 33155 2160 33175 2180
rect 33155 2110 33175 2130
rect 33155 2060 33175 2080
rect 33155 2010 33175 2030
rect 33155 1960 33175 1980
rect 33210 2210 33230 2230
rect 33210 2160 33230 2180
rect 33210 2110 33230 2130
rect 33210 2060 33230 2080
rect 33210 2010 33230 2030
rect 33210 1960 33230 1980
rect 33265 2210 33285 2230
rect 33265 2160 33285 2180
rect 33265 2110 33285 2130
rect 33265 2060 33285 2080
rect 33265 2010 33285 2030
rect 33265 1960 33285 1980
rect 33320 2210 33340 2230
rect 33320 2160 33340 2180
rect 33320 2110 33340 2130
rect 33320 2060 33340 2080
rect 33320 2010 33340 2030
rect 33320 1960 33340 1980
rect 33375 2210 33395 2230
rect 33375 2160 33395 2180
rect 33375 2110 33395 2130
rect 33375 2060 33395 2080
rect 33375 2010 33395 2030
rect 33375 1960 33395 1980
rect 33430 2210 33450 2230
rect 33430 2160 33450 2180
rect 33430 2110 33450 2130
rect 33430 2060 33450 2080
rect 33430 2010 33450 2030
rect 33430 1960 33450 1980
rect 33485 2210 33505 2230
rect 33485 2160 33505 2180
rect 33485 2110 33505 2130
rect 33485 2060 33505 2080
rect 33485 2010 33505 2030
rect 33485 1960 33505 1980
rect 33540 2210 33560 2230
rect 33540 2160 33560 2180
rect 33540 2110 33560 2130
rect 33540 2060 33560 2080
rect 33540 2010 33560 2030
rect 33540 1960 33560 1980
rect 33595 2210 33615 2230
rect 33595 2160 33615 2180
rect 33595 2110 33615 2130
rect 33595 2060 33615 2080
rect 33595 2010 33615 2030
rect 33595 1960 33615 1980
rect 33650 2210 33670 2230
rect 33650 2160 33670 2180
rect 33650 2110 33670 2130
rect 33650 2060 33670 2080
rect 33650 2010 33670 2030
rect 33650 1960 33670 1980
rect 33705 2210 33725 2230
rect 33705 2160 33725 2180
rect 33705 2110 33725 2130
rect 33705 2060 33725 2080
rect 33705 2010 33725 2030
rect 33705 1960 33725 1980
rect 33760 2210 33780 2230
rect 33760 2160 33780 2180
rect 33760 2110 33780 2130
rect 33760 2060 33780 2080
rect 33760 2010 33780 2030
rect 33760 1960 33780 1980
rect 33815 2210 33835 2230
rect 33815 2160 33835 2180
rect 33815 2110 33835 2130
rect 33815 2060 33835 2080
rect 33815 2010 33835 2030
rect 33815 1960 33835 1980
rect 30045 1620 30065 1640
rect 30045 1570 30065 1590
rect 30045 1520 30065 1540
rect 30045 1470 30065 1490
rect 30045 1420 30065 1440
rect 30045 1370 30065 1390
rect 30045 1320 30065 1340
rect 30045 1270 30065 1290
rect 30045 1220 30065 1240
rect 30045 1170 30065 1190
rect 30045 1120 30065 1140
rect 30045 1070 30065 1090
rect 30045 1020 30065 1040
rect 30045 970 30065 990
rect 30145 1620 30165 1640
rect 30145 1570 30165 1590
rect 30145 1520 30165 1540
rect 30145 1470 30165 1490
rect 30145 1420 30165 1440
rect 30145 1370 30165 1390
rect 30145 1320 30165 1340
rect 30145 1270 30165 1290
rect 30145 1220 30165 1240
rect 30145 1170 30165 1190
rect 30145 1120 30165 1140
rect 30145 1070 30165 1090
rect 30145 1020 30165 1040
rect 30145 970 30165 990
rect 30245 1620 30265 1640
rect 30245 1570 30265 1590
rect 30245 1520 30265 1540
rect 30245 1470 30265 1490
rect 30245 1420 30265 1440
rect 30245 1370 30265 1390
rect 30245 1320 30265 1340
rect 30245 1270 30265 1290
rect 30245 1220 30265 1240
rect 30245 1170 30265 1190
rect 30245 1120 30265 1140
rect 30245 1070 30265 1090
rect 30245 1020 30265 1040
rect 30245 970 30265 990
rect 30345 1620 30365 1640
rect 30345 1570 30365 1590
rect 30345 1520 30365 1540
rect 30345 1470 30365 1490
rect 30345 1420 30365 1440
rect 30345 1370 30365 1390
rect 30345 1320 30365 1340
rect 30345 1270 30365 1290
rect 30345 1220 30365 1240
rect 30345 1170 30365 1190
rect 30345 1120 30365 1140
rect 30345 1070 30365 1090
rect 30345 1020 30365 1040
rect 30345 970 30365 990
rect 30445 1620 30465 1640
rect 30445 1570 30465 1590
rect 30445 1520 30465 1540
rect 30445 1470 30465 1490
rect 30445 1420 30465 1440
rect 30445 1370 30465 1390
rect 30445 1320 30465 1340
rect 30445 1270 30465 1290
rect 30445 1220 30465 1240
rect 30445 1170 30465 1190
rect 30445 1120 30465 1140
rect 30445 1070 30465 1090
rect 30445 1020 30465 1040
rect 30445 970 30465 990
rect 30545 1620 30565 1640
rect 30545 1570 30565 1590
rect 30545 1520 30565 1540
rect 30545 1470 30565 1490
rect 30545 1420 30565 1440
rect 30545 1370 30565 1390
rect 30545 1320 30565 1340
rect 30545 1270 30565 1290
rect 30545 1220 30565 1240
rect 30545 1170 30565 1190
rect 30545 1120 30565 1140
rect 30545 1070 30565 1090
rect 30545 1020 30565 1040
rect 30545 970 30565 990
rect 30645 1620 30665 1640
rect 30645 1570 30665 1590
rect 30645 1520 30665 1540
rect 30645 1470 30665 1490
rect 30645 1420 30665 1440
rect 30645 1370 30665 1390
rect 30645 1320 30665 1340
rect 30645 1270 30665 1290
rect 30645 1220 30665 1240
rect 30645 1170 30665 1190
rect 30645 1120 30665 1140
rect 30645 1070 30665 1090
rect 30645 1020 30665 1040
rect 30645 970 30665 990
rect 31040 1675 31060 1695
rect 31040 1625 31060 1645
rect 31040 1575 31060 1595
rect 31095 1675 31115 1695
rect 31095 1625 31115 1645
rect 31095 1575 31115 1595
rect 31150 1675 31170 1695
rect 31150 1625 31170 1645
rect 31150 1575 31170 1595
rect 31205 1675 31225 1695
rect 31205 1625 31225 1645
rect 31205 1575 31225 1595
rect 31260 1675 31280 1695
rect 31260 1625 31280 1645
rect 31260 1575 31280 1595
rect 31315 1675 31335 1695
rect 31315 1625 31335 1645
rect 31315 1575 31335 1595
rect 31370 1675 31390 1695
rect 31370 1625 31390 1645
rect 31370 1575 31390 1595
rect 31425 1675 31445 1695
rect 31425 1625 31445 1645
rect 31425 1575 31445 1595
rect 31480 1675 31500 1695
rect 31480 1625 31500 1645
rect 31480 1575 31500 1595
rect 31535 1675 31555 1695
rect 31535 1625 31555 1645
rect 31535 1575 31555 1595
rect 31590 1675 31610 1695
rect 31590 1625 31610 1645
rect 31590 1575 31610 1595
rect 31645 1675 31665 1695
rect 31645 1625 31665 1645
rect 31645 1575 31665 1595
rect 31700 1675 31720 1695
rect 31700 1625 31720 1645
rect 31700 1575 31720 1595
rect 31780 1675 31800 1695
rect 31780 1625 31800 1645
rect 31780 1575 31800 1595
rect 31835 1675 31855 1695
rect 31835 1625 31855 1645
rect 31835 1575 31855 1595
rect 31890 1675 31910 1695
rect 31890 1625 31910 1645
rect 31890 1575 31910 1595
rect 31945 1675 31965 1695
rect 31945 1625 31965 1645
rect 31945 1575 31965 1595
rect 32000 1675 32020 1695
rect 32000 1625 32020 1645
rect 32000 1575 32020 1595
rect 32080 1675 32100 1695
rect 32080 1625 32100 1645
rect 32080 1575 32100 1595
rect 32135 1675 32155 1695
rect 32135 1625 32155 1645
rect 32135 1575 32155 1595
rect 32190 1675 32210 1695
rect 32190 1625 32210 1645
rect 32190 1575 32210 1595
rect 32245 1675 32265 1695
rect 32245 1625 32265 1645
rect 32245 1575 32265 1595
rect 32300 1675 32320 1695
rect 32300 1625 32320 1645
rect 32300 1575 32320 1595
rect 32355 1675 32375 1695
rect 32355 1625 32375 1645
rect 32355 1575 32375 1595
rect 32410 1675 32430 1695
rect 32410 1625 32430 1645
rect 32410 1575 32430 1595
rect 32465 1675 32485 1695
rect 32465 1625 32485 1645
rect 32465 1575 32485 1595
rect 32520 1675 32540 1695
rect 32520 1625 32540 1645
rect 32520 1575 32540 1595
rect 32575 1675 32595 1695
rect 32575 1625 32595 1645
rect 32575 1575 32595 1595
rect 32630 1675 32650 1695
rect 32630 1625 32650 1645
rect 32630 1575 32650 1595
rect 32685 1675 32705 1695
rect 32685 1625 32705 1645
rect 32685 1575 32705 1595
rect 32740 1675 32760 1695
rect 32740 1625 32760 1645
rect 32740 1575 32760 1595
rect 31215 1170 31235 1190
rect 31215 1120 31235 1140
rect 31215 1070 31235 1090
rect 31215 1020 31235 1040
rect 31215 970 31235 990
rect 31270 1170 31290 1190
rect 31270 1120 31290 1140
rect 31270 1070 31290 1090
rect 31270 1020 31290 1040
rect 31270 970 31290 990
rect 31325 1170 31345 1190
rect 31325 1120 31345 1140
rect 31325 1070 31345 1090
rect 31325 1020 31345 1040
rect 31325 970 31345 990
rect 31380 1170 31400 1190
rect 31380 1120 31400 1140
rect 31380 1070 31400 1090
rect 31380 1020 31400 1040
rect 31380 970 31400 990
rect 31435 1170 31455 1190
rect 31435 1120 31455 1140
rect 31435 1070 31455 1090
rect 31435 1020 31455 1040
rect 31435 970 31455 990
rect 31490 1170 31510 1190
rect 31490 1120 31510 1140
rect 31490 1070 31510 1090
rect 31490 1020 31510 1040
rect 31490 970 31510 990
rect 31545 1170 31565 1190
rect 31545 1120 31565 1140
rect 31545 1070 31565 1090
rect 31545 1020 31565 1040
rect 31545 970 31565 990
rect 31600 1170 31620 1190
rect 31600 1120 31620 1140
rect 31600 1070 31620 1090
rect 31600 1020 31620 1040
rect 31600 970 31620 990
rect 31655 1170 31675 1190
rect 31655 1120 31675 1140
rect 31655 1070 31675 1090
rect 31655 1020 31675 1040
rect 31655 970 31675 990
rect 31710 1170 31730 1190
rect 31710 1120 31730 1140
rect 31710 1070 31730 1090
rect 31710 1020 31730 1040
rect 31710 970 31730 990
rect 31765 1170 31785 1190
rect 31765 1120 31785 1140
rect 31765 1070 31785 1090
rect 31765 1020 31785 1040
rect 31765 970 31785 990
rect 31820 1170 31840 1190
rect 31820 1120 31840 1140
rect 31820 1070 31840 1090
rect 31820 1020 31840 1040
rect 31820 970 31840 990
rect 31875 1170 31895 1190
rect 31875 1120 31895 1140
rect 31875 1070 31895 1090
rect 31875 1020 31895 1040
rect 31875 970 31895 990
rect 31930 1170 31950 1190
rect 31930 1120 31950 1140
rect 31930 1070 31950 1090
rect 31930 1020 31950 1040
rect 31930 970 31950 990
rect 31985 1170 32005 1190
rect 31985 1120 32005 1140
rect 31985 1070 32005 1090
rect 31985 1020 32005 1040
rect 31985 970 32005 990
rect 32040 1170 32060 1190
rect 32040 1120 32060 1140
rect 32040 1070 32060 1090
rect 32040 1020 32060 1040
rect 32040 970 32060 990
rect 32095 1170 32115 1190
rect 32095 1120 32115 1140
rect 32095 1070 32115 1090
rect 32095 1020 32115 1040
rect 32095 970 32115 990
rect 32150 1170 32170 1190
rect 32150 1120 32170 1140
rect 32150 1070 32170 1090
rect 32150 1020 32170 1040
rect 32150 970 32170 990
rect 32205 1170 32225 1190
rect 32205 1120 32225 1140
rect 32205 1070 32225 1090
rect 32205 1020 32225 1040
rect 32205 970 32225 990
rect 32260 1170 32280 1190
rect 32260 1120 32280 1140
rect 32260 1070 32280 1090
rect 32260 1020 32280 1040
rect 32260 970 32280 990
rect 32315 1170 32335 1190
rect 32315 1120 32335 1140
rect 32315 1070 32335 1090
rect 32315 1020 32335 1040
rect 32315 970 32335 990
rect 32370 1170 32390 1190
rect 32370 1120 32390 1140
rect 32370 1070 32390 1090
rect 32370 1020 32390 1040
rect 32370 970 32390 990
rect 32425 1170 32445 1190
rect 32425 1120 32445 1140
rect 32425 1070 32445 1090
rect 32425 1020 32445 1040
rect 32425 970 32445 990
rect 32480 1170 32500 1190
rect 32480 1120 32500 1140
rect 32480 1070 32500 1090
rect 32480 1020 32500 1040
rect 32480 970 32500 990
rect 33135 1620 33155 1640
rect 33135 1570 33155 1590
rect 33135 1520 33155 1540
rect 33135 1470 33155 1490
rect 33135 1420 33155 1440
rect 33135 1370 33155 1390
rect 33135 1320 33155 1340
rect 33135 1270 33155 1290
rect 33135 1220 33155 1240
rect 33135 1170 33155 1190
rect 33135 1120 33155 1140
rect 33135 1070 33155 1090
rect 33135 1020 33155 1040
rect 33135 970 33155 990
rect 33235 1620 33255 1640
rect 33235 1570 33255 1590
rect 33235 1520 33255 1540
rect 33235 1470 33255 1490
rect 33235 1420 33255 1440
rect 33235 1370 33255 1390
rect 33235 1320 33255 1340
rect 33235 1270 33255 1290
rect 33235 1220 33255 1240
rect 33235 1170 33255 1190
rect 33235 1120 33255 1140
rect 33235 1070 33255 1090
rect 33235 1020 33255 1040
rect 33235 970 33255 990
rect 33335 1620 33355 1640
rect 33335 1570 33355 1590
rect 33335 1520 33355 1540
rect 33335 1470 33355 1490
rect 33335 1420 33355 1440
rect 33335 1370 33355 1390
rect 33335 1320 33355 1340
rect 33335 1270 33355 1290
rect 33335 1220 33355 1240
rect 33335 1170 33355 1190
rect 33335 1120 33355 1140
rect 33335 1070 33355 1090
rect 33335 1020 33355 1040
rect 33335 970 33355 990
rect 33435 1620 33455 1640
rect 33435 1570 33455 1590
rect 33435 1520 33455 1540
rect 33435 1470 33455 1490
rect 33435 1420 33455 1440
rect 33435 1370 33455 1390
rect 33435 1320 33455 1340
rect 33435 1270 33455 1290
rect 33435 1220 33455 1240
rect 33435 1170 33455 1190
rect 33435 1120 33455 1140
rect 33435 1070 33455 1090
rect 33435 1020 33455 1040
rect 33435 970 33455 990
rect 33535 1620 33555 1640
rect 33535 1570 33555 1590
rect 33535 1520 33555 1540
rect 33535 1470 33555 1490
rect 33535 1420 33555 1440
rect 33535 1370 33555 1390
rect 33535 1320 33555 1340
rect 33535 1270 33555 1290
rect 33535 1220 33555 1240
rect 33535 1170 33555 1190
rect 33535 1120 33555 1140
rect 33535 1070 33555 1090
rect 33535 1020 33555 1040
rect 33535 970 33555 990
rect 33635 1620 33655 1640
rect 33635 1570 33655 1590
rect 33635 1520 33655 1540
rect 33635 1470 33655 1490
rect 33635 1420 33655 1440
rect 33635 1370 33655 1390
rect 33635 1320 33655 1340
rect 33635 1270 33655 1290
rect 33635 1220 33655 1240
rect 33635 1170 33655 1190
rect 33635 1120 33655 1140
rect 33635 1070 33655 1090
rect 33635 1020 33655 1040
rect 33635 970 33655 990
rect 33735 1620 33755 1640
rect 33735 1570 33755 1590
rect 33735 1520 33755 1540
rect 33735 1470 33755 1490
rect 33735 1420 33755 1440
rect 33735 1370 33755 1390
rect 33735 1320 33755 1340
rect 33735 1270 33755 1290
rect 33735 1220 33755 1240
rect 33735 1170 33755 1190
rect 33735 1120 33755 1140
rect 33735 1070 33755 1090
rect 33735 1020 33755 1040
rect 33735 970 33755 990
rect 31270 655 31290 675
rect 31270 605 31290 625
rect 31500 655 31520 675
rect 31500 605 31520 625
rect 31890 650 31910 670
rect 31945 650 31965 670
rect 32000 650 32020 670
rect 32055 650 32075 670
rect 32110 650 32130 670
rect 32165 650 32185 670
rect 32220 650 32240 670
rect 32275 650 32295 670
rect 32330 650 32350 670
rect 32385 650 32405 670
rect 32440 650 32460 670
rect 32495 650 32515 670
rect 32550 650 32570 670
<< pdiffc >>
rect 31230 4775 31250 4795
rect 31290 4775 31310 4795
rect 31350 4775 31370 4795
rect 31410 4775 31430 4795
rect 31480 4785 31500 4805
rect 31540 4785 31560 4805
rect 31600 4785 31620 4805
rect 31660 4785 31680 4805
rect 31720 4785 31740 4805
rect 31780 4785 31800 4805
rect 31840 4785 31860 4805
rect 32210 4770 32230 4790
rect 32270 4770 32290 4790
rect 32330 4770 32350 4790
rect 32390 4770 32410 4790
rect 32450 4770 32470 4790
rect 32510 4770 32530 4790
rect 32570 4770 32590 4790
rect 32630 4770 32650 4790
rect 32690 4770 32710 4790
rect 31260 4355 31280 4375
rect 31315 4355 31335 4375
rect 31370 4355 31390 4375
rect 31425 4355 31445 4375
rect 31480 4355 31500 4375
rect 31535 4355 31555 4375
rect 31590 4355 31610 4375
rect 31645 4355 31665 4375
rect 31700 4355 31720 4375
rect 31755 4355 31775 4375
rect 31810 4355 31830 4375
rect 31865 4355 31885 4375
rect 31920 4355 31940 4375
rect 31975 4355 31995 4375
rect 32030 4355 32050 4375
rect 32085 4355 32105 4375
rect 32140 4355 32160 4375
rect 32195 4355 32215 4375
rect 32250 4355 32270 4375
rect 32305 4355 32325 4375
rect 32360 4355 32380 4375
rect 32415 4355 32435 4375
rect 32470 4355 32490 4375
rect 31210 3945 31230 3965
rect 31265 3945 31285 3965
rect 31320 3945 31340 3965
rect 31375 3945 31395 3965
rect 31430 3945 31450 3965
rect 31485 3945 31505 3965
rect 31540 3945 31560 3965
rect 31595 3945 31615 3965
rect 31650 3945 31670 3965
rect 31705 3945 31725 3965
rect 31760 3945 31780 3965
rect 31815 3945 31835 3965
rect 31870 3945 31890 3965
rect 31940 3945 31960 3965
rect 31995 3945 32015 3965
rect 32050 3945 32070 3965
rect 32105 3945 32125 3965
rect 32160 3945 32180 3965
rect 32215 3945 32235 3965
rect 32270 3945 32290 3965
rect 32325 3945 32345 3965
rect 32380 3945 32400 3965
rect 32435 3945 32455 3965
rect 32490 3945 32510 3965
rect 32545 3945 32565 3965
rect 32600 3945 32620 3965
rect 29965 3630 29985 3650
rect 29965 3580 29985 3600
rect 29965 3530 29985 3550
rect 29965 3480 29985 3500
rect 29965 3430 29985 3450
rect 29965 3380 29985 3400
rect 29965 3330 29985 3350
rect 29965 3280 29985 3300
rect 29965 3230 29985 3250
rect 29965 3180 29985 3200
rect 29965 3130 29985 3150
rect 29965 3080 29985 3100
rect 30020 3630 30040 3650
rect 30020 3580 30040 3600
rect 30020 3530 30040 3550
rect 30020 3480 30040 3500
rect 30020 3430 30040 3450
rect 30020 3380 30040 3400
rect 30020 3330 30040 3350
rect 30020 3280 30040 3300
rect 30020 3230 30040 3250
rect 30020 3180 30040 3200
rect 30020 3130 30040 3150
rect 30020 3080 30040 3100
rect 30075 3630 30095 3650
rect 30075 3580 30095 3600
rect 30075 3530 30095 3550
rect 30075 3480 30095 3500
rect 30075 3430 30095 3450
rect 30075 3380 30095 3400
rect 30075 3330 30095 3350
rect 30075 3280 30095 3300
rect 30075 3230 30095 3250
rect 30075 3180 30095 3200
rect 30075 3130 30095 3150
rect 30075 3080 30095 3100
rect 30130 3630 30150 3650
rect 30130 3580 30150 3600
rect 30130 3530 30150 3550
rect 30130 3480 30150 3500
rect 30130 3430 30150 3450
rect 30130 3380 30150 3400
rect 30130 3330 30150 3350
rect 30130 3280 30150 3300
rect 30130 3230 30150 3250
rect 30130 3180 30150 3200
rect 30130 3130 30150 3150
rect 30130 3080 30150 3100
rect 30185 3630 30205 3650
rect 30185 3580 30205 3600
rect 30185 3530 30205 3550
rect 30185 3480 30205 3500
rect 30185 3430 30205 3450
rect 30185 3380 30205 3400
rect 30185 3330 30205 3350
rect 30185 3280 30205 3300
rect 30185 3230 30205 3250
rect 30185 3180 30205 3200
rect 30185 3130 30205 3150
rect 30185 3080 30205 3100
rect 30240 3630 30260 3650
rect 30240 3580 30260 3600
rect 30240 3530 30260 3550
rect 30240 3480 30260 3500
rect 30240 3430 30260 3450
rect 30240 3380 30260 3400
rect 30240 3330 30260 3350
rect 30240 3280 30260 3300
rect 30240 3230 30260 3250
rect 30240 3180 30260 3200
rect 30240 3130 30260 3150
rect 30240 3080 30260 3100
rect 30295 3630 30315 3650
rect 30295 3580 30315 3600
rect 30295 3530 30315 3550
rect 30295 3480 30315 3500
rect 30295 3430 30315 3450
rect 30295 3380 30315 3400
rect 30295 3330 30315 3350
rect 30295 3280 30315 3300
rect 30295 3230 30315 3250
rect 30295 3180 30315 3200
rect 30295 3130 30315 3150
rect 30295 3080 30315 3100
rect 30350 3630 30370 3650
rect 30350 3580 30370 3600
rect 30350 3530 30370 3550
rect 30350 3480 30370 3500
rect 30350 3430 30370 3450
rect 30350 3380 30370 3400
rect 30350 3330 30370 3350
rect 30350 3280 30370 3300
rect 30350 3230 30370 3250
rect 30350 3180 30370 3200
rect 30350 3130 30370 3150
rect 30350 3080 30370 3100
rect 30405 3630 30425 3650
rect 30405 3580 30425 3600
rect 30405 3530 30425 3550
rect 30405 3480 30425 3500
rect 30405 3430 30425 3450
rect 30405 3380 30425 3400
rect 30405 3330 30425 3350
rect 30405 3280 30425 3300
rect 30405 3230 30425 3250
rect 30405 3180 30425 3200
rect 30405 3130 30425 3150
rect 30405 3080 30425 3100
rect 30460 3630 30480 3650
rect 30460 3580 30480 3600
rect 30460 3530 30480 3550
rect 30460 3480 30480 3500
rect 30460 3430 30480 3450
rect 30460 3380 30480 3400
rect 30460 3330 30480 3350
rect 30460 3280 30480 3300
rect 30460 3230 30480 3250
rect 30460 3180 30480 3200
rect 30460 3130 30480 3150
rect 30460 3080 30480 3100
rect 30515 3630 30535 3650
rect 30515 3580 30535 3600
rect 30515 3530 30535 3550
rect 30515 3480 30535 3500
rect 30515 3430 30535 3450
rect 30515 3380 30535 3400
rect 30515 3330 30535 3350
rect 30515 3280 30535 3300
rect 30515 3230 30535 3250
rect 30515 3180 30535 3200
rect 30515 3130 30535 3150
rect 30515 3080 30535 3100
rect 30570 3630 30590 3650
rect 30570 3580 30590 3600
rect 30570 3530 30590 3550
rect 30570 3480 30590 3500
rect 30570 3430 30590 3450
rect 30570 3380 30590 3400
rect 30570 3330 30590 3350
rect 30570 3280 30590 3300
rect 30570 3230 30590 3250
rect 30570 3180 30590 3200
rect 30570 3130 30590 3150
rect 30570 3080 30590 3100
rect 30625 3630 30645 3650
rect 30625 3580 30645 3600
rect 30625 3530 30645 3550
rect 30625 3480 30645 3500
rect 30625 3430 30645 3450
rect 30625 3380 30645 3400
rect 30625 3330 30645 3350
rect 30625 3280 30645 3300
rect 30625 3230 30645 3250
rect 30625 3180 30645 3200
rect 30625 3130 30645 3150
rect 30625 3080 30645 3100
rect 31230 3520 31250 3540
rect 31230 3470 31250 3490
rect 31230 3420 31250 3440
rect 31230 3370 31250 3390
rect 31230 3320 31250 3340
rect 31230 3270 31250 3290
rect 31230 3220 31250 3240
rect 31290 3520 31310 3540
rect 31290 3470 31310 3490
rect 31290 3420 31310 3440
rect 31290 3370 31310 3390
rect 31290 3320 31310 3340
rect 31290 3270 31310 3290
rect 31290 3220 31310 3240
rect 31350 3520 31370 3540
rect 31350 3470 31370 3490
rect 31350 3420 31370 3440
rect 31350 3370 31370 3390
rect 31350 3320 31370 3340
rect 31350 3270 31370 3290
rect 31350 3220 31370 3240
rect 31410 3520 31430 3540
rect 31410 3470 31430 3490
rect 31410 3420 31430 3440
rect 31410 3370 31430 3390
rect 31410 3320 31430 3340
rect 31410 3270 31430 3290
rect 31410 3220 31430 3240
rect 31470 3520 31490 3540
rect 31470 3470 31490 3490
rect 31470 3420 31490 3440
rect 31470 3370 31490 3390
rect 31470 3320 31490 3340
rect 31470 3270 31490 3290
rect 31470 3220 31490 3240
rect 31530 3520 31550 3540
rect 31530 3470 31550 3490
rect 31530 3420 31550 3440
rect 31530 3370 31550 3390
rect 31530 3320 31550 3340
rect 31530 3270 31550 3290
rect 31530 3220 31550 3240
rect 31590 3520 31610 3540
rect 31590 3470 31610 3490
rect 31590 3420 31610 3440
rect 31590 3370 31610 3390
rect 31590 3320 31610 3340
rect 31590 3270 31610 3290
rect 31590 3220 31610 3240
rect 31650 3520 31670 3540
rect 31650 3470 31670 3490
rect 31650 3420 31670 3440
rect 31650 3370 31670 3390
rect 31650 3320 31670 3340
rect 31650 3270 31670 3290
rect 31650 3220 31670 3240
rect 31710 3520 31730 3540
rect 31710 3470 31730 3490
rect 31710 3420 31730 3440
rect 31710 3370 31730 3390
rect 31710 3320 31730 3340
rect 31710 3270 31730 3290
rect 31710 3220 31730 3240
rect 31770 3520 31790 3540
rect 31770 3470 31790 3490
rect 31770 3420 31790 3440
rect 31770 3370 31790 3390
rect 31770 3320 31790 3340
rect 31770 3270 31790 3290
rect 31770 3220 31790 3240
rect 31830 3520 31850 3540
rect 31830 3470 31850 3490
rect 31830 3420 31850 3440
rect 31830 3370 31850 3390
rect 31830 3320 31850 3340
rect 31830 3270 31850 3290
rect 31830 3220 31850 3240
rect 31890 3520 31910 3540
rect 31890 3470 31910 3490
rect 31890 3420 31910 3440
rect 31890 3370 31910 3390
rect 31890 3320 31910 3340
rect 31890 3270 31910 3290
rect 31890 3220 31910 3240
rect 31950 3520 31970 3540
rect 31950 3470 31970 3490
rect 31950 3420 31970 3440
rect 31950 3370 31970 3390
rect 31950 3320 31970 3340
rect 31950 3270 31970 3290
rect 31950 3220 31970 3240
rect 32010 3520 32030 3540
rect 32010 3470 32030 3490
rect 32010 3420 32030 3440
rect 32010 3370 32030 3390
rect 32010 3320 32030 3340
rect 32010 3270 32030 3290
rect 32010 3220 32030 3240
rect 32070 3520 32090 3540
rect 32070 3470 32090 3490
rect 32070 3420 32090 3440
rect 32070 3370 32090 3390
rect 32070 3320 32090 3340
rect 32070 3270 32090 3290
rect 32070 3220 32090 3240
rect 32130 3520 32150 3540
rect 32130 3470 32150 3490
rect 32130 3420 32150 3440
rect 32130 3370 32150 3390
rect 32130 3320 32150 3340
rect 32130 3270 32150 3290
rect 32130 3220 32150 3240
rect 32190 3520 32210 3540
rect 32190 3470 32210 3490
rect 32190 3420 32210 3440
rect 32190 3370 32210 3390
rect 32190 3320 32210 3340
rect 32190 3270 32210 3290
rect 32190 3220 32210 3240
rect 32250 3520 32270 3540
rect 32250 3470 32270 3490
rect 32250 3420 32270 3440
rect 32250 3370 32270 3390
rect 32250 3320 32270 3340
rect 32250 3270 32270 3290
rect 32250 3220 32270 3240
rect 32310 3520 32330 3540
rect 32310 3470 32330 3490
rect 32310 3420 32330 3440
rect 32310 3370 32330 3390
rect 32310 3320 32330 3340
rect 32310 3270 32330 3290
rect 32310 3220 32330 3240
rect 32370 3520 32390 3540
rect 32370 3470 32390 3490
rect 32370 3420 32390 3440
rect 32370 3370 32390 3390
rect 32370 3320 32390 3340
rect 32370 3270 32390 3290
rect 32370 3220 32390 3240
rect 32430 3520 32450 3540
rect 32430 3470 32450 3490
rect 32430 3420 32450 3440
rect 32430 3370 32450 3390
rect 32430 3320 32450 3340
rect 32430 3270 32450 3290
rect 32430 3220 32450 3240
rect 32490 3520 32510 3540
rect 32490 3470 32510 3490
rect 32490 3420 32510 3440
rect 32490 3370 32510 3390
rect 32490 3320 32510 3340
rect 32490 3270 32510 3290
rect 32490 3220 32510 3240
rect 32550 3520 32570 3540
rect 32550 3470 32570 3490
rect 32550 3420 32570 3440
rect 32550 3370 32570 3390
rect 32550 3320 32570 3340
rect 32550 3270 32570 3290
rect 32550 3220 32570 3240
rect 33155 3630 33175 3650
rect 33155 3580 33175 3600
rect 33155 3530 33175 3550
rect 33155 3480 33175 3500
rect 33155 3430 33175 3450
rect 33155 3380 33175 3400
rect 33155 3330 33175 3350
rect 33155 3280 33175 3300
rect 33155 3230 33175 3250
rect 33155 3180 33175 3200
rect 33155 3130 33175 3150
rect 33155 3080 33175 3100
rect 33210 3630 33230 3650
rect 33210 3580 33230 3600
rect 33210 3530 33230 3550
rect 33210 3480 33230 3500
rect 33210 3430 33230 3450
rect 33210 3380 33230 3400
rect 33210 3330 33230 3350
rect 33210 3280 33230 3300
rect 33210 3230 33230 3250
rect 33210 3180 33230 3200
rect 33210 3130 33230 3150
rect 33210 3080 33230 3100
rect 33265 3630 33285 3650
rect 33265 3580 33285 3600
rect 33265 3530 33285 3550
rect 33265 3480 33285 3500
rect 33265 3430 33285 3450
rect 33265 3380 33285 3400
rect 33265 3330 33285 3350
rect 33265 3280 33285 3300
rect 33265 3230 33285 3250
rect 33265 3180 33285 3200
rect 33265 3130 33285 3150
rect 33265 3080 33285 3100
rect 33320 3630 33340 3650
rect 33320 3580 33340 3600
rect 33320 3530 33340 3550
rect 33320 3480 33340 3500
rect 33320 3430 33340 3450
rect 33320 3380 33340 3400
rect 33320 3330 33340 3350
rect 33320 3280 33340 3300
rect 33320 3230 33340 3250
rect 33320 3180 33340 3200
rect 33320 3130 33340 3150
rect 33320 3080 33340 3100
rect 33375 3630 33395 3650
rect 33375 3580 33395 3600
rect 33375 3530 33395 3550
rect 33375 3480 33395 3500
rect 33375 3430 33395 3450
rect 33375 3380 33395 3400
rect 33375 3330 33395 3350
rect 33375 3280 33395 3300
rect 33375 3230 33395 3250
rect 33375 3180 33395 3200
rect 33375 3130 33395 3150
rect 33375 3080 33395 3100
rect 33430 3630 33450 3650
rect 33430 3580 33450 3600
rect 33430 3530 33450 3550
rect 33430 3480 33450 3500
rect 33430 3430 33450 3450
rect 33430 3380 33450 3400
rect 33430 3330 33450 3350
rect 33430 3280 33450 3300
rect 33430 3230 33450 3250
rect 33430 3180 33450 3200
rect 33430 3130 33450 3150
rect 33430 3080 33450 3100
rect 33485 3630 33505 3650
rect 33485 3580 33505 3600
rect 33485 3530 33505 3550
rect 33485 3480 33505 3500
rect 33485 3430 33505 3450
rect 33485 3380 33505 3400
rect 33485 3330 33505 3350
rect 33485 3280 33505 3300
rect 33485 3230 33505 3250
rect 33485 3180 33505 3200
rect 33485 3130 33505 3150
rect 33485 3080 33505 3100
rect 33540 3630 33560 3650
rect 33540 3580 33560 3600
rect 33540 3530 33560 3550
rect 33540 3480 33560 3500
rect 33540 3430 33560 3450
rect 33540 3380 33560 3400
rect 33540 3330 33560 3350
rect 33540 3280 33560 3300
rect 33540 3230 33560 3250
rect 33540 3180 33560 3200
rect 33540 3130 33560 3150
rect 33540 3080 33560 3100
rect 33595 3630 33615 3650
rect 33595 3580 33615 3600
rect 33595 3530 33615 3550
rect 33595 3480 33615 3500
rect 33595 3430 33615 3450
rect 33595 3380 33615 3400
rect 33595 3330 33615 3350
rect 33595 3280 33615 3300
rect 33595 3230 33615 3250
rect 33595 3180 33615 3200
rect 33595 3130 33615 3150
rect 33595 3080 33615 3100
rect 33650 3630 33670 3650
rect 33650 3580 33670 3600
rect 33650 3530 33670 3550
rect 33650 3480 33670 3500
rect 33650 3430 33670 3450
rect 33650 3380 33670 3400
rect 33650 3330 33670 3350
rect 33650 3280 33670 3300
rect 33650 3230 33670 3250
rect 33650 3180 33670 3200
rect 33650 3130 33670 3150
rect 33650 3080 33670 3100
rect 33705 3630 33725 3650
rect 33705 3580 33725 3600
rect 33705 3530 33725 3550
rect 33705 3480 33725 3500
rect 33705 3430 33725 3450
rect 33705 3380 33725 3400
rect 33705 3330 33725 3350
rect 33705 3280 33725 3300
rect 33705 3230 33725 3250
rect 33705 3180 33725 3200
rect 33705 3130 33725 3150
rect 33705 3080 33725 3100
rect 33760 3630 33780 3650
rect 33760 3580 33780 3600
rect 33760 3530 33780 3550
rect 33760 3480 33780 3500
rect 33760 3430 33780 3450
rect 33760 3380 33780 3400
rect 33760 3330 33780 3350
rect 33760 3280 33780 3300
rect 33760 3230 33780 3250
rect 33760 3180 33780 3200
rect 33760 3130 33780 3150
rect 33760 3080 33780 3100
rect 33815 3630 33835 3650
rect 33815 3580 33835 3600
rect 33815 3530 33835 3550
rect 33815 3480 33835 3500
rect 33815 3430 33835 3450
rect 33815 3380 33835 3400
rect 33815 3330 33835 3350
rect 33815 3280 33835 3300
rect 33815 3230 33835 3250
rect 33815 3180 33835 3200
rect 33815 3130 33835 3150
rect 33815 3080 33835 3100
rect 29965 2670 29985 2690
rect 29965 2620 29985 2640
rect 29965 2570 29985 2590
rect 29965 2520 29985 2540
rect 30020 2670 30040 2690
rect 30020 2620 30040 2640
rect 30020 2570 30040 2590
rect 30020 2520 30040 2540
rect 30075 2670 30095 2690
rect 30075 2620 30095 2640
rect 30075 2570 30095 2590
rect 30075 2520 30095 2540
rect 30130 2670 30150 2690
rect 30130 2620 30150 2640
rect 30130 2570 30150 2590
rect 30130 2520 30150 2540
rect 30185 2670 30205 2690
rect 30185 2620 30205 2640
rect 30185 2570 30205 2590
rect 30185 2520 30205 2540
rect 30240 2670 30260 2690
rect 30240 2620 30260 2640
rect 30240 2570 30260 2590
rect 30240 2520 30260 2540
rect 30295 2670 30315 2690
rect 30295 2620 30315 2640
rect 30295 2570 30315 2590
rect 30295 2520 30315 2540
rect 30350 2670 30370 2690
rect 30350 2620 30370 2640
rect 30350 2570 30370 2590
rect 30350 2520 30370 2540
rect 30405 2670 30425 2690
rect 30405 2620 30425 2640
rect 30405 2570 30425 2590
rect 30405 2520 30425 2540
rect 30460 2670 30480 2690
rect 30460 2620 30480 2640
rect 30460 2570 30480 2590
rect 30460 2520 30480 2540
rect 30515 2670 30535 2690
rect 30515 2620 30535 2640
rect 30515 2570 30535 2590
rect 30515 2520 30535 2540
rect 30570 2670 30590 2690
rect 30570 2620 30590 2640
rect 30570 2570 30590 2590
rect 30570 2520 30590 2540
rect 30625 2670 30645 2690
rect 30625 2620 30645 2640
rect 30625 2570 30645 2590
rect 30625 2520 30645 2540
rect 31015 2810 31035 2830
rect 31015 2760 31035 2780
rect 31015 2710 31035 2730
rect 31015 2660 31035 2680
rect 31015 2610 31035 2630
rect 31015 2560 31035 2580
rect 31015 2510 31035 2530
rect 31075 2810 31095 2830
rect 31075 2760 31095 2780
rect 31075 2710 31095 2730
rect 31075 2660 31095 2680
rect 31075 2610 31095 2630
rect 31075 2560 31095 2580
rect 31075 2510 31095 2530
rect 31135 2810 31155 2830
rect 31135 2760 31155 2780
rect 31135 2710 31155 2730
rect 31135 2660 31155 2680
rect 31135 2610 31155 2630
rect 31135 2560 31155 2580
rect 31135 2510 31155 2530
rect 31195 2810 31215 2830
rect 31195 2760 31215 2780
rect 31195 2710 31215 2730
rect 31195 2660 31215 2680
rect 31195 2610 31215 2630
rect 31195 2560 31215 2580
rect 31195 2510 31215 2530
rect 31255 2810 31275 2830
rect 31255 2760 31275 2780
rect 31255 2710 31275 2730
rect 31255 2660 31275 2680
rect 31255 2610 31275 2630
rect 31255 2560 31275 2580
rect 31255 2510 31275 2530
rect 31315 2810 31335 2830
rect 31315 2760 31335 2780
rect 31315 2710 31335 2730
rect 31315 2660 31335 2680
rect 31315 2610 31335 2630
rect 31315 2560 31335 2580
rect 31315 2510 31335 2530
rect 31375 2810 31395 2830
rect 31375 2760 31395 2780
rect 31375 2710 31395 2730
rect 31375 2660 31395 2680
rect 31375 2610 31395 2630
rect 31375 2560 31395 2580
rect 31375 2510 31395 2530
rect 31435 2810 31455 2830
rect 31435 2760 31455 2780
rect 31435 2710 31455 2730
rect 31435 2660 31455 2680
rect 31435 2610 31455 2630
rect 31435 2560 31455 2580
rect 31435 2510 31455 2530
rect 31495 2810 31515 2830
rect 31495 2760 31515 2780
rect 31495 2710 31515 2730
rect 31495 2660 31515 2680
rect 31495 2610 31515 2630
rect 31495 2560 31515 2580
rect 31495 2510 31515 2530
rect 31555 2810 31575 2830
rect 31555 2760 31575 2780
rect 31555 2710 31575 2730
rect 31555 2660 31575 2680
rect 31555 2610 31575 2630
rect 31555 2560 31575 2580
rect 31555 2510 31575 2530
rect 31615 2810 31635 2830
rect 31615 2760 31635 2780
rect 31615 2710 31635 2730
rect 31615 2660 31635 2680
rect 31615 2610 31635 2630
rect 31615 2560 31635 2580
rect 31615 2510 31635 2530
rect 31675 2810 31695 2830
rect 31675 2760 31695 2780
rect 31675 2710 31695 2730
rect 31675 2660 31695 2680
rect 31675 2610 31695 2630
rect 31675 2560 31695 2580
rect 31675 2510 31695 2530
rect 31735 2810 31755 2830
rect 31735 2760 31755 2780
rect 31735 2710 31755 2730
rect 31735 2660 31755 2680
rect 31735 2610 31755 2630
rect 31735 2560 31755 2580
rect 31735 2510 31755 2530
rect 32045 2810 32065 2830
rect 32045 2760 32065 2780
rect 32045 2710 32065 2730
rect 32045 2660 32065 2680
rect 32045 2610 32065 2630
rect 32045 2560 32065 2580
rect 32045 2510 32065 2530
rect 32105 2810 32125 2830
rect 32105 2760 32125 2780
rect 32105 2710 32125 2730
rect 32105 2660 32125 2680
rect 32105 2610 32125 2630
rect 32105 2560 32125 2580
rect 32105 2510 32125 2530
rect 32165 2810 32185 2830
rect 32165 2760 32185 2780
rect 32165 2710 32185 2730
rect 32165 2660 32185 2680
rect 32165 2610 32185 2630
rect 32165 2560 32185 2580
rect 32165 2510 32185 2530
rect 32225 2810 32245 2830
rect 32225 2760 32245 2780
rect 32225 2710 32245 2730
rect 32225 2660 32245 2680
rect 32225 2610 32245 2630
rect 32225 2560 32245 2580
rect 32225 2510 32245 2530
rect 32285 2810 32305 2830
rect 32285 2760 32305 2780
rect 32285 2710 32305 2730
rect 32285 2660 32305 2680
rect 32285 2610 32305 2630
rect 32285 2560 32305 2580
rect 32285 2510 32305 2530
rect 32345 2810 32365 2830
rect 32345 2760 32365 2780
rect 32345 2710 32365 2730
rect 32345 2660 32365 2680
rect 32345 2610 32365 2630
rect 32345 2560 32365 2580
rect 32345 2510 32365 2530
rect 32405 2810 32425 2830
rect 32405 2760 32425 2780
rect 32405 2710 32425 2730
rect 32405 2660 32425 2680
rect 32405 2610 32425 2630
rect 32405 2560 32425 2580
rect 32405 2510 32425 2530
rect 32465 2810 32485 2830
rect 32465 2760 32485 2780
rect 32465 2710 32485 2730
rect 32465 2660 32485 2680
rect 32465 2610 32485 2630
rect 32465 2560 32485 2580
rect 32465 2510 32485 2530
rect 32525 2810 32545 2830
rect 32525 2760 32545 2780
rect 32525 2710 32545 2730
rect 32525 2660 32545 2680
rect 32525 2610 32545 2630
rect 32525 2560 32545 2580
rect 32525 2510 32545 2530
rect 32585 2810 32605 2830
rect 32585 2760 32605 2780
rect 32585 2710 32605 2730
rect 32585 2660 32605 2680
rect 32585 2610 32605 2630
rect 32585 2560 32605 2580
rect 32585 2510 32605 2530
rect 32645 2810 32665 2830
rect 32645 2760 32665 2780
rect 32645 2710 32665 2730
rect 32645 2660 32665 2680
rect 32645 2610 32665 2630
rect 32645 2560 32665 2580
rect 32645 2510 32665 2530
rect 32705 2810 32725 2830
rect 32705 2760 32725 2780
rect 32705 2710 32725 2730
rect 32705 2660 32725 2680
rect 32705 2610 32725 2630
rect 32705 2560 32725 2580
rect 32705 2510 32725 2530
rect 32765 2810 32785 2830
rect 32765 2760 32785 2780
rect 32765 2710 32785 2730
rect 32765 2660 32785 2680
rect 32765 2610 32785 2630
rect 32765 2560 32785 2580
rect 32765 2510 32785 2530
rect 33155 2670 33175 2690
rect 33155 2620 33175 2640
rect 33155 2570 33175 2590
rect 33155 2520 33175 2540
rect 33210 2670 33230 2690
rect 33210 2620 33230 2640
rect 33210 2570 33230 2590
rect 33210 2520 33230 2540
rect 33265 2670 33285 2690
rect 33265 2620 33285 2640
rect 33265 2570 33285 2590
rect 33265 2520 33285 2540
rect 33320 2670 33340 2690
rect 33320 2620 33340 2640
rect 33320 2570 33340 2590
rect 33320 2520 33340 2540
rect 33375 2670 33395 2690
rect 33375 2620 33395 2640
rect 33375 2570 33395 2590
rect 33375 2520 33395 2540
rect 33430 2670 33450 2690
rect 33430 2620 33450 2640
rect 33430 2570 33450 2590
rect 33430 2520 33450 2540
rect 33485 2670 33505 2690
rect 33485 2620 33505 2640
rect 33485 2570 33505 2590
rect 33485 2520 33505 2540
rect 33540 2670 33560 2690
rect 33540 2620 33560 2640
rect 33540 2570 33560 2590
rect 33540 2520 33560 2540
rect 33595 2670 33615 2690
rect 33595 2620 33615 2640
rect 33595 2570 33615 2590
rect 33595 2520 33615 2540
rect 33650 2670 33670 2690
rect 33650 2620 33670 2640
rect 33650 2570 33670 2590
rect 33650 2520 33670 2540
rect 33705 2670 33725 2690
rect 33705 2620 33725 2640
rect 33705 2570 33725 2590
rect 33705 2520 33725 2540
rect 33760 2670 33780 2690
rect 33760 2620 33780 2640
rect 33760 2570 33780 2590
rect 33760 2520 33780 2540
rect 33815 2670 33835 2690
rect 33815 2620 33835 2640
rect 33815 2570 33835 2590
rect 33815 2520 33835 2540
<< psubdiff >>
rect 29485 3680 29765 3700
rect 29485 3375 29505 3680
rect 29485 2995 29505 3280
rect 29745 3375 29765 3680
rect 29745 2995 29765 3280
rect 29485 2975 29585 2995
rect 29665 2975 29765 2995
rect 34035 3680 34315 3700
rect 34035 3375 34055 3680
rect 34035 2995 34055 3280
rect 34295 3375 34315 3680
rect 34295 2995 34315 3280
rect 34035 2975 34135 2995
rect 34215 2975 34315 2995
rect 29400 2649 29535 2669
rect 29615 2649 29755 2669
rect 29400 2335 29420 2649
rect 29400 1925 29420 2255
rect 29735 2335 29755 2649
rect 34045 2649 34185 2669
rect 34265 2649 34400 2669
rect 29735 1925 29755 2255
rect 29400 1905 29535 1925
rect 29615 1905 29755 1925
rect 29905 2320 30265 2340
rect 30345 2320 30705 2340
rect 29905 2135 29925 2320
rect 29905 1870 29925 2055
rect 30685 2135 30705 2320
rect 33095 2320 33455 2340
rect 33535 2320 33895 2340
rect 30685 1870 30705 2055
rect 31095 2255 31860 2275
rect 31940 2255 32705 2275
rect 31095 2145 31115 2255
rect 31095 1955 31115 2065
rect 32685 2145 32705 2255
rect 32685 1955 32705 2065
rect 31095 1935 31860 1955
rect 31940 1935 32705 1955
rect 33095 2135 33115 2320
rect 29905 1850 30265 1870
rect 30345 1850 30705 1870
rect 33095 1870 33115 2055
rect 33875 2135 33895 2320
rect 33875 1870 33895 2055
rect 34045 2335 34065 2649
rect 34045 1925 34065 2255
rect 34380 2335 34400 2649
rect 34380 1925 34400 2255
rect 34045 1905 34185 1925
rect 34265 1905 34400 1925
rect 33095 1850 33455 1870
rect 33535 1850 33895 1870
rect 30940 1785 31860 1805
rect 31940 1785 32860 1805
rect 29985 1730 30315 1750
rect 30395 1730 30725 1750
rect 29660 1675 29735 1695
rect 29815 1675 29895 1695
rect 29660 1300 29680 1675
rect 29660 868 29680 1220
rect 29875 1300 29895 1675
rect 29875 868 29895 1220
rect 29660 848 29735 868
rect 29815 848 29895 868
rect 29985 1345 30005 1730
rect 29985 880 30005 1265
rect 30705 1345 30725 1730
rect 30940 1675 30960 1785
rect 30940 1485 30960 1595
rect 32840 1675 32860 1785
rect 32840 1485 32860 1595
rect 30940 1465 31860 1485
rect 31940 1465 32860 1485
rect 33075 1730 33405 1750
rect 33485 1730 33815 1750
rect 33075 1345 33095 1730
rect 30705 880 30725 1265
rect 29985 860 30315 880
rect 30395 860 30725 880
rect 31155 1280 31845 1300
rect 31925 1280 32565 1300
rect 31155 1100 31175 1280
rect 31155 875 31175 1020
rect 32545 1100 32565 1280
rect 32545 875 32565 1020
rect 31155 855 31845 875
rect 31925 855 32565 875
rect 33075 880 33095 1265
rect 33795 1345 33815 1730
rect 33795 880 33815 1265
rect 33075 860 33405 880
rect 33485 860 33815 880
rect 33905 1675 33985 1695
rect 34065 1675 34140 1695
rect 33905 1300 33925 1675
rect 33905 868 33925 1220
rect 34120 1300 34140 1675
rect 34120 868 34140 1220
rect 33905 848 33985 868
rect 34065 848 34140 868
rect 31210 765 31355 785
rect 31435 765 31585 785
rect 31210 695 31230 765
rect 31565 695 31585 765
rect 31210 555 31230 615
rect 31565 555 31585 615
rect 31210 535 31355 555
rect 31435 535 31585 555
rect 31830 760 32190 780
rect 32270 760 32630 780
rect 31830 690 31850 760
rect 32610 690 32630 760
rect 31830 560 31850 610
rect 32610 560 32630 610
rect 31830 540 32190 560
rect 32270 540 32630 560
<< nsubdiff >>
rect 31170 4910 31485 4930
rect 31565 4910 31920 4930
rect 31170 4825 31190 4910
rect 31900 4825 31920 4910
rect 31170 4675 31190 4745
rect 31900 4675 31920 4745
rect 31170 4655 31485 4675
rect 31565 4655 31920 4675
rect 32150 4885 32420 4905
rect 32500 4885 32770 4905
rect 32150 4820 32170 4885
rect 32750 4825 32770 4885
rect 32150 4675 32170 4740
rect 32750 4675 32770 4740
rect 32150 4655 32420 4675
rect 32500 4655 32770 4675
rect 31200 4465 31835 4485
rect 31915 4465 32550 4485
rect 31200 4405 31220 4465
rect 32530 4405 32550 4465
rect 31200 4265 31220 4325
rect 32530 4265 32550 4325
rect 31200 4245 31835 4265
rect 31915 4245 32550 4265
rect 31150 4055 31875 4075
rect 31955 4055 32680 4075
rect 31150 3995 31170 4055
rect 32660 3995 32680 4055
rect 31150 3855 31170 3915
rect 32660 3855 32680 3915
rect 31150 3835 31875 3855
rect 31955 3835 32680 3855
rect 29905 3740 30265 3760
rect 30345 3740 30705 3760
rect 29905 3410 29925 3740
rect 29905 2990 29925 3315
rect 30685 3410 30705 3740
rect 33095 3740 33455 3760
rect 33535 3740 33895 3760
rect 30685 2990 30705 3315
rect 31170 3630 31860 3650
rect 31940 3630 32630 3650
rect 31170 3445 31190 3630
rect 31170 3130 31190 3365
rect 32610 3445 32630 3630
rect 32610 3130 32630 3365
rect 31170 3110 31860 3130
rect 31940 3110 32630 3130
rect 33095 3410 33115 3740
rect 29905 2970 30265 2990
rect 30345 2970 30705 2990
rect 33095 2990 33115 3315
rect 33875 3410 33895 3740
rect 33875 2990 33895 3315
rect 33095 2970 33455 2990
rect 33535 2970 33895 2990
rect 30955 2920 31345 2940
rect 31425 2920 31815 2940
rect 29905 2780 30265 2800
rect 30345 2780 30705 2800
rect 29905 2645 29925 2780
rect 29905 2430 29925 2565
rect 30685 2645 30705 2780
rect 30685 2430 30705 2565
rect 29905 2410 30265 2430
rect 30345 2410 30705 2430
rect 30955 2710 30975 2920
rect 30955 2420 30975 2630
rect 31795 2710 31815 2920
rect 31795 2420 31815 2630
rect 30955 2400 31345 2420
rect 31425 2400 31815 2420
rect 31985 2920 32375 2940
rect 32455 2920 32845 2940
rect 31985 2710 32005 2920
rect 31985 2420 32005 2630
rect 32825 2710 32845 2920
rect 32825 2420 32845 2630
rect 31985 2400 32375 2420
rect 32455 2400 32845 2420
rect 33095 2780 33455 2800
rect 33535 2780 33895 2800
rect 33095 2645 33115 2780
rect 33095 2430 33115 2565
rect 33875 2645 33895 2780
rect 33875 2430 33895 2565
rect 33095 2410 33455 2430
rect 33535 2410 33895 2430
<< psubdiffcont >>
rect 29485 3280 29505 3375
rect 29745 3280 29765 3375
rect 29585 2975 29665 2995
rect 34035 3280 34055 3375
rect 34295 3280 34315 3375
rect 34135 2975 34215 2995
rect 29535 2649 29615 2669
rect 29400 2255 29420 2335
rect 34185 2649 34265 2669
rect 29735 2255 29755 2335
rect 29535 1905 29615 1925
rect 30265 2320 30345 2340
rect 29905 2055 29925 2135
rect 33455 2320 33535 2340
rect 30685 2055 30705 2135
rect 31860 2255 31940 2275
rect 31095 2065 31115 2145
rect 32685 2065 32705 2145
rect 31860 1935 31940 1955
rect 33095 2055 33115 2135
rect 30265 1850 30345 1870
rect 33875 2055 33895 2135
rect 34045 2255 34065 2335
rect 34380 2255 34400 2335
rect 34185 1905 34265 1925
rect 33455 1850 33535 1870
rect 31860 1785 31940 1805
rect 30315 1730 30395 1750
rect 29735 1675 29815 1695
rect 29660 1220 29680 1300
rect 29875 1220 29895 1300
rect 29735 848 29815 868
rect 29985 1265 30005 1345
rect 30940 1595 30960 1675
rect 32840 1595 32860 1675
rect 31860 1465 31940 1485
rect 33405 1730 33485 1750
rect 30705 1265 30725 1345
rect 30315 860 30395 880
rect 31845 1280 31925 1300
rect 31155 1020 31175 1100
rect 32545 1020 32565 1100
rect 31845 855 31925 875
rect 33075 1265 33095 1345
rect 33795 1265 33815 1345
rect 33405 860 33485 880
rect 33985 1675 34065 1695
rect 33905 1220 33925 1300
rect 34120 1220 34140 1300
rect 33985 848 34065 868
rect 31355 765 31435 785
rect 31210 615 31230 695
rect 31565 615 31585 695
rect 31355 535 31435 555
rect 32190 760 32270 780
rect 31830 610 31850 690
rect 32610 610 32630 690
rect 32190 540 32270 560
<< nsubdiffcont >>
rect 31485 4910 31565 4930
rect 31170 4745 31190 4825
rect 31900 4745 31920 4825
rect 31485 4655 31565 4675
rect 32420 4885 32500 4905
rect 32150 4740 32170 4820
rect 32750 4740 32770 4825
rect 32420 4655 32500 4675
rect 31835 4465 31915 4485
rect 31200 4325 31220 4405
rect 32530 4325 32550 4405
rect 31835 4245 31915 4265
rect 31875 4055 31955 4075
rect 31150 3915 31170 3995
rect 32660 3915 32680 3995
rect 31875 3835 31955 3855
rect 30265 3740 30345 3760
rect 29905 3315 29925 3410
rect 33455 3740 33535 3760
rect 30685 3315 30705 3410
rect 31860 3630 31940 3650
rect 31170 3365 31190 3445
rect 32610 3365 32630 3445
rect 31860 3110 31940 3130
rect 33095 3315 33115 3410
rect 30265 2970 30345 2990
rect 33875 3315 33895 3410
rect 33455 2970 33535 2990
rect 31345 2920 31425 2940
rect 30265 2780 30345 2800
rect 29905 2565 29925 2645
rect 30685 2565 30705 2645
rect 30265 2410 30345 2430
rect 30955 2630 30975 2710
rect 31795 2630 31815 2710
rect 31345 2400 31425 2420
rect 32375 2920 32455 2940
rect 31985 2630 32005 2710
rect 32825 2630 32845 2710
rect 32375 2400 32455 2420
rect 33455 2780 33535 2800
rect 33095 2565 33115 2645
rect 33875 2565 33895 2645
rect 33455 2410 33535 2430
<< poly >>
rect 31830 4880 31870 4890
rect 31830 4865 31840 4880
rect 31810 4860 31840 4865
rect 31860 4860 31870 4880
rect 31810 4850 31870 4860
rect 31510 4835 31530 4850
rect 31570 4835 31590 4850
rect 31630 4835 31650 4850
rect 31690 4835 31710 4850
rect 31750 4835 31770 4850
rect 31810 4835 31830 4850
rect 31260 4818 31280 4835
rect 31320 4818 31340 4833
rect 31380 4818 31400 4833
rect 31260 4745 31280 4755
rect 31225 4730 31280 4745
rect 31320 4740 31340 4755
rect 31380 4745 31400 4755
rect 31510 4745 31530 4755
rect 31310 4730 31350 4740
rect 31380 4730 31435 4745
rect 31225 4710 31230 4730
rect 31250 4710 31255 4730
rect 31225 4700 31255 4710
rect 31310 4710 31320 4730
rect 31340 4710 31350 4730
rect 31310 4700 31350 4710
rect 31405 4710 31410 4730
rect 31430 4710 31435 4730
rect 31405 4700 31435 4710
rect 31475 4730 31530 4745
rect 31570 4745 31590 4755
rect 31630 4745 31650 4755
rect 31690 4745 31710 4755
rect 31750 4745 31770 4755
rect 31570 4730 31770 4745
rect 31810 4745 31830 4755
rect 31810 4730 31865 4745
rect 31475 4710 31480 4730
rect 31500 4710 31505 4730
rect 31475 4700 31505 4710
rect 31650 4725 31690 4730
rect 31650 4705 31660 4725
rect 31680 4705 31690 4725
rect 31650 4695 31690 4705
rect 31835 4710 31840 4730
rect 31860 4710 31865 4730
rect 31835 4700 31865 4710
rect 32240 4810 32260 4825
rect 32300 4810 32320 4825
rect 32360 4810 32380 4825
rect 32420 4810 32440 4825
rect 32480 4810 32500 4825
rect 32540 4810 32560 4825
rect 32600 4810 32620 4825
rect 32660 4810 32680 4825
rect 32240 4740 32260 4750
rect 32205 4725 32260 4740
rect 32300 4740 32320 4750
rect 32360 4740 32380 4750
rect 32420 4740 32440 4750
rect 32480 4740 32500 4750
rect 32540 4740 32560 4750
rect 32600 4740 32620 4750
rect 32300 4725 32620 4740
rect 32660 4740 32680 4750
rect 32660 4725 32715 4740
rect 32205 4705 32210 4725
rect 32230 4705 32235 4725
rect 32205 4695 32235 4705
rect 32323 4705 32331 4725
rect 32349 4705 32357 4725
rect 32323 4695 32357 4705
rect 32685 4705 32690 4725
rect 32710 4705 32715 4725
rect 32685 4695 32715 4705
rect 31290 4390 31305 4405
rect 31345 4390 31360 4405
rect 31400 4390 31415 4405
rect 31455 4390 31470 4405
rect 31510 4390 31525 4405
rect 31565 4390 31580 4405
rect 31620 4390 31635 4405
rect 31675 4390 31690 4405
rect 31730 4390 31745 4405
rect 31785 4390 31800 4405
rect 31840 4390 31855 4405
rect 31895 4390 31910 4405
rect 31950 4390 31965 4405
rect 32005 4390 32020 4405
rect 32060 4390 32075 4405
rect 32115 4390 32130 4405
rect 32170 4390 32185 4405
rect 32225 4390 32240 4405
rect 32280 4390 32295 4405
rect 32335 4390 32350 4405
rect 32390 4390 32405 4405
rect 32445 4390 32460 4405
rect 31290 4330 31305 4340
rect 31255 4315 31305 4330
rect 31345 4330 31360 4340
rect 31400 4330 31415 4340
rect 31455 4330 31470 4340
rect 31510 4330 31525 4340
rect 31565 4330 31580 4340
rect 31620 4330 31635 4340
rect 31675 4330 31690 4340
rect 31730 4330 31745 4340
rect 31785 4330 31800 4340
rect 31840 4330 31855 4340
rect 31895 4330 31910 4340
rect 31950 4330 31965 4340
rect 32005 4330 32020 4340
rect 32060 4330 32075 4340
rect 32115 4330 32130 4340
rect 32170 4330 32185 4340
rect 32225 4330 32240 4340
rect 32280 4330 32295 4340
rect 32335 4330 32350 4340
rect 32390 4330 32405 4340
rect 31345 4315 32405 4330
rect 32445 4330 32460 4340
rect 32445 4315 32495 4330
rect 31255 4295 31260 4315
rect 31280 4295 31285 4315
rect 31255 4285 31285 4295
rect 31362 4295 31370 4315
rect 31390 4295 31398 4315
rect 31362 4285 31398 4295
rect 32465 4295 32470 4315
rect 32490 4295 32495 4315
rect 32465 4285 32495 4295
rect 31280 4025 31310 4035
rect 31280 4005 31285 4025
rect 31305 4005 31310 4025
rect 31480 4025 31510 4035
rect 31480 4005 31485 4025
rect 31505 4005 31510 4025
rect 31695 4025 31735 4035
rect 31695 4005 31705 4025
rect 31725 4005 31735 4025
rect 32008 4025 32038 4035
rect 32008 4005 32013 4025
rect 32033 4005 32038 4025
rect 32205 4025 32245 4035
rect 32205 4005 32215 4025
rect 32235 4005 32245 4025
rect 32425 4025 32465 4035
rect 32425 4005 32435 4025
rect 32455 4005 32465 4025
rect 31280 3995 31310 4005
rect 31240 3980 31255 3995
rect 31295 3980 31310 3995
rect 31350 3980 31365 3995
rect 31405 3980 31420 3995
rect 31460 3990 31530 4005
rect 31460 3980 31475 3990
rect 31515 3980 31530 3990
rect 31570 3980 31585 3995
rect 31625 3980 31640 3995
rect 31680 3990 31750 4005
rect 32008 3995 32040 4005
rect 31680 3980 31695 3990
rect 31735 3980 31750 3990
rect 31790 3980 31805 3995
rect 31845 3980 31860 3995
rect 31970 3980 31985 3995
rect 32025 3980 32040 3995
rect 32080 3980 32095 3995
rect 32135 3980 32150 3995
rect 32190 3990 32260 4005
rect 32190 3980 32205 3990
rect 32245 3980 32260 3990
rect 32300 3980 32315 3995
rect 32355 3980 32370 3995
rect 32410 3990 32480 4005
rect 32410 3980 32425 3990
rect 32465 3980 32480 3990
rect 32520 3980 32535 3995
rect 32575 3980 32590 3995
rect 31240 3920 31255 3930
rect 31205 3905 31255 3920
rect 31295 3915 31310 3930
rect 31350 3920 31365 3930
rect 31405 3920 31420 3930
rect 31350 3915 31420 3920
rect 31460 3915 31475 3930
rect 31515 3915 31530 3930
rect 31570 3920 31585 3930
rect 31625 3920 31640 3930
rect 31570 3915 31640 3920
rect 31680 3915 31695 3930
rect 31735 3915 31750 3930
rect 31790 3915 31805 3930
rect 31350 3905 31439 3915
rect 31570 3905 31659 3915
rect 31205 3885 31210 3905
rect 31230 3885 31235 3905
rect 31205 3875 31235 3885
rect 31407 3885 31413 3905
rect 31430 3885 31439 3905
rect 31407 3875 31439 3885
rect 31627 3885 31633 3905
rect 31650 3885 31659 3905
rect 31627 3875 31659 3885
rect 31771 3905 31805 3915
rect 31845 3920 31860 3930
rect 31970 3920 31985 3930
rect 31845 3905 31895 3920
rect 31771 3885 31780 3905
rect 31797 3885 31805 3905
rect 31771 3875 31805 3885
rect 31865 3885 31870 3905
rect 31890 3885 31895 3905
rect 31865 3875 31895 3885
rect 31935 3905 31985 3920
rect 32025 3915 32040 3930
rect 32080 3920 32095 3930
rect 32135 3920 32150 3930
rect 32080 3915 32150 3920
rect 32190 3915 32205 3930
rect 32245 3915 32260 3930
rect 32300 3920 32315 3930
rect 32355 3920 32370 3930
rect 32300 3915 32370 3920
rect 32410 3915 32425 3930
rect 32465 3915 32480 3930
rect 32520 3915 32535 3930
rect 32080 3905 32169 3915
rect 32300 3905 32389 3915
rect 31935 3885 31940 3905
rect 31960 3885 31965 3905
rect 31935 3875 31965 3885
rect 32137 3885 32143 3905
rect 32160 3885 32169 3905
rect 32137 3875 32169 3885
rect 32357 3885 32363 3905
rect 32380 3885 32389 3905
rect 32357 3875 32389 3885
rect 32501 3905 32535 3915
rect 32575 3920 32590 3930
rect 32575 3905 32625 3920
rect 32501 3885 32510 3905
rect 32527 3885 32535 3905
rect 32501 3875 32535 3885
rect 32595 3885 32600 3905
rect 32620 3885 32625 3905
rect 32595 3875 32625 3885
rect 29995 3665 30010 3680
rect 30050 3665 30065 3680
rect 30105 3665 30120 3680
rect 30160 3665 30175 3680
rect 30215 3665 30230 3680
rect 30270 3665 30285 3680
rect 30325 3665 30340 3680
rect 30380 3665 30395 3680
rect 30435 3665 30450 3680
rect 30490 3665 30505 3680
rect 30545 3665 30560 3680
rect 30600 3665 30615 3680
rect 29995 3055 30010 3065
rect 29960 3040 30010 3055
rect 30050 3055 30065 3065
rect 30105 3055 30120 3065
rect 30160 3055 30175 3065
rect 30215 3055 30230 3065
rect 30270 3055 30285 3065
rect 30325 3055 30340 3065
rect 30380 3055 30395 3065
rect 30435 3055 30450 3065
rect 30490 3055 30505 3065
rect 30545 3055 30560 3065
rect 30050 3040 30560 3055
rect 30600 3055 30615 3065
rect 30600 3040 30650 3055
rect 29960 3020 29965 3040
rect 29985 3020 29990 3040
rect 29960 3010 29990 3020
rect 30178 3020 30186 3040
rect 30204 3020 30212 3040
rect 30178 3010 30212 3020
rect 30620 3020 30625 3040
rect 30645 3020 30650 3040
rect 30620 3010 30650 3020
rect 31260 3555 31280 3570
rect 31320 3555 31340 3570
rect 31380 3555 31400 3570
rect 31440 3555 31460 3570
rect 31500 3555 31520 3570
rect 31560 3555 31580 3570
rect 31620 3555 31640 3570
rect 31680 3555 31700 3570
rect 31740 3555 31760 3570
rect 31800 3555 31820 3570
rect 31860 3555 31880 3570
rect 31920 3555 31940 3570
rect 31980 3555 32000 3570
rect 32040 3555 32060 3570
rect 32100 3555 32120 3570
rect 32160 3555 32180 3570
rect 32220 3555 32240 3570
rect 32280 3555 32300 3570
rect 32340 3555 32360 3570
rect 32400 3555 32420 3570
rect 32460 3555 32480 3570
rect 32520 3555 32540 3570
rect 31260 3195 31280 3205
rect 31225 3180 31280 3195
rect 31320 3195 31340 3205
rect 31380 3195 31400 3205
rect 31440 3195 31460 3205
rect 31500 3195 31520 3205
rect 31560 3195 31580 3205
rect 31620 3195 31640 3205
rect 31680 3195 31700 3205
rect 31740 3195 31760 3205
rect 31800 3195 31820 3205
rect 31860 3195 31880 3205
rect 31920 3195 31940 3205
rect 31980 3195 32000 3205
rect 32040 3195 32060 3205
rect 32100 3195 32120 3205
rect 32160 3195 32180 3205
rect 32220 3195 32240 3205
rect 32280 3195 32300 3205
rect 32340 3195 32360 3205
rect 32400 3195 32420 3205
rect 32460 3195 32480 3205
rect 31320 3180 32480 3195
rect 32520 3195 32540 3205
rect 32520 3180 32575 3195
rect 31225 3160 31230 3180
rect 31250 3160 31255 3180
rect 31225 3150 31255 3160
rect 31823 3160 31831 3180
rect 31849 3160 31857 3180
rect 31823 3150 31857 3160
rect 32545 3160 32550 3180
rect 32570 3160 32575 3180
rect 32545 3150 32575 3160
rect 33185 3665 33200 3680
rect 33240 3665 33255 3680
rect 33295 3665 33310 3680
rect 33350 3665 33365 3680
rect 33405 3665 33420 3680
rect 33460 3665 33475 3680
rect 33515 3665 33530 3680
rect 33570 3665 33585 3680
rect 33625 3665 33640 3680
rect 33680 3665 33695 3680
rect 33735 3665 33750 3680
rect 33790 3665 33805 3680
rect 33185 3055 33200 3065
rect 33150 3040 33200 3055
rect 33240 3055 33255 3065
rect 33295 3055 33310 3065
rect 33350 3055 33365 3065
rect 33405 3055 33420 3065
rect 33460 3055 33475 3065
rect 33515 3055 33530 3065
rect 33570 3055 33585 3065
rect 33625 3055 33640 3065
rect 33680 3055 33695 3065
rect 33735 3055 33750 3065
rect 33240 3040 33750 3055
rect 33790 3055 33805 3065
rect 33790 3040 33840 3055
rect 33150 3020 33155 3040
rect 33175 3020 33180 3040
rect 33150 3010 33180 3020
rect 33588 3020 33596 3040
rect 33614 3020 33622 3040
rect 33588 3010 33622 3020
rect 33810 3020 33815 3040
rect 33835 3020 33840 3040
rect 33810 3010 33840 3020
rect 29995 2705 30010 2720
rect 30050 2705 30065 2720
rect 30105 2705 30120 2720
rect 30160 2705 30175 2720
rect 30215 2705 30230 2720
rect 30270 2705 30285 2720
rect 30325 2705 30340 2720
rect 30380 2705 30395 2720
rect 30435 2705 30450 2720
rect 30490 2705 30505 2720
rect 30545 2705 30560 2720
rect 30600 2705 30615 2720
rect 29995 2495 30010 2505
rect 29960 2480 30010 2495
rect 30050 2495 30065 2505
rect 30105 2495 30120 2505
rect 30160 2495 30175 2505
rect 30215 2495 30230 2505
rect 30270 2495 30285 2505
rect 30325 2495 30340 2505
rect 30380 2495 30395 2505
rect 30435 2495 30450 2505
rect 30490 2495 30505 2505
rect 30545 2495 30560 2505
rect 30050 2480 30560 2495
rect 30600 2495 30615 2505
rect 30600 2480 30650 2495
rect 29960 2460 29965 2480
rect 29985 2460 29990 2480
rect 29960 2450 29990 2460
rect 30453 2460 30461 2480
rect 30479 2460 30487 2480
rect 30453 2450 30487 2460
rect 30620 2460 30625 2480
rect 30645 2460 30650 2480
rect 30620 2450 30650 2460
rect 31045 2845 31065 2860
rect 31105 2845 31125 2860
rect 31165 2845 31185 2860
rect 31225 2845 31245 2860
rect 31285 2845 31305 2860
rect 31345 2845 31365 2860
rect 31405 2845 31425 2860
rect 31465 2845 31485 2860
rect 31525 2845 31545 2860
rect 31585 2845 31605 2860
rect 31645 2845 31665 2860
rect 31705 2845 31725 2860
rect 31045 2485 31065 2495
rect 31010 2470 31065 2485
rect 31105 2485 31125 2495
rect 31165 2485 31185 2495
rect 31225 2485 31245 2495
rect 31285 2485 31305 2495
rect 31345 2485 31365 2495
rect 31405 2485 31425 2495
rect 31465 2485 31485 2495
rect 31525 2485 31545 2495
rect 31585 2485 31605 2495
rect 31645 2485 31665 2495
rect 31105 2470 31665 2485
rect 31705 2485 31725 2495
rect 31705 2470 31760 2485
rect 31010 2450 31015 2470
rect 31035 2450 31040 2470
rect 31010 2440 31040 2450
rect 31368 2450 31376 2470
rect 31394 2450 31402 2470
rect 31368 2440 31402 2450
rect 31730 2450 31735 2470
rect 31755 2450 31760 2470
rect 31730 2440 31760 2450
rect 32075 2845 32095 2860
rect 32135 2845 32155 2860
rect 32195 2845 32215 2860
rect 32255 2845 32275 2860
rect 32315 2845 32335 2860
rect 32375 2845 32395 2860
rect 32435 2845 32455 2860
rect 32495 2845 32515 2860
rect 32555 2845 32575 2860
rect 32615 2845 32635 2860
rect 32675 2845 32695 2860
rect 32735 2845 32755 2860
rect 32075 2485 32095 2495
rect 32040 2470 32095 2485
rect 32135 2485 32155 2495
rect 32195 2485 32215 2495
rect 32255 2485 32275 2495
rect 32315 2485 32335 2495
rect 32375 2485 32395 2495
rect 32435 2485 32455 2495
rect 32495 2485 32515 2495
rect 32555 2485 32575 2495
rect 32615 2485 32635 2495
rect 32675 2485 32695 2495
rect 32135 2470 32695 2485
rect 32735 2485 32755 2495
rect 32735 2470 32790 2485
rect 32040 2450 32045 2470
rect 32065 2450 32070 2470
rect 32040 2440 32070 2450
rect 32398 2450 32406 2470
rect 32424 2450 32432 2470
rect 32398 2440 32432 2450
rect 32760 2450 32765 2470
rect 32785 2450 32790 2470
rect 32760 2440 32790 2450
rect 33185 2705 33200 2720
rect 33240 2705 33255 2720
rect 33295 2705 33310 2720
rect 33350 2705 33365 2720
rect 33405 2705 33420 2720
rect 33460 2705 33475 2720
rect 33515 2705 33530 2720
rect 33570 2705 33585 2720
rect 33625 2705 33640 2720
rect 33680 2705 33695 2720
rect 33735 2705 33750 2720
rect 33790 2705 33805 2720
rect 33185 2495 33200 2505
rect 33150 2480 33200 2495
rect 33240 2495 33255 2505
rect 33295 2495 33310 2505
rect 33350 2495 33365 2505
rect 33405 2495 33420 2505
rect 33460 2495 33475 2505
rect 33515 2495 33530 2505
rect 33570 2495 33585 2505
rect 33625 2495 33640 2505
rect 33680 2495 33695 2505
rect 33735 2495 33750 2505
rect 33240 2480 33750 2495
rect 33790 2495 33805 2505
rect 33790 2480 33840 2495
rect 33150 2460 33155 2480
rect 33175 2460 33180 2480
rect 33150 2450 33180 2460
rect 33313 2460 33321 2480
rect 33339 2460 33347 2480
rect 33313 2450 33347 2460
rect 33810 2460 33815 2480
rect 33835 2460 33840 2480
rect 33810 2450 33840 2460
rect 29960 2290 29990 2300
rect 29960 2270 29965 2290
rect 29985 2270 29990 2290
rect 30453 2290 30487 2300
rect 30453 2270 30461 2290
rect 30479 2270 30487 2290
rect 30620 2290 30650 2300
rect 30620 2270 30625 2290
rect 30645 2270 30650 2290
rect 29960 2255 30010 2270
rect 29995 2245 30010 2255
rect 30050 2255 30560 2270
rect 30050 2245 30065 2255
rect 30105 2245 30120 2255
rect 30160 2245 30175 2255
rect 30215 2245 30230 2255
rect 30270 2245 30285 2255
rect 30325 2245 30340 2255
rect 30380 2245 30395 2255
rect 30435 2245 30450 2255
rect 30490 2245 30505 2255
rect 30545 2245 30560 2255
rect 30600 2255 30650 2270
rect 30600 2245 30615 2255
rect 29995 1930 30010 1945
rect 30050 1930 30065 1945
rect 30105 1930 30120 1945
rect 30160 1930 30175 1945
rect 30215 1930 30230 1945
rect 30270 1930 30285 1945
rect 30325 1930 30340 1945
rect 30380 1930 30395 1945
rect 30435 1930 30450 1945
rect 30490 1930 30505 1945
rect 30545 1930 30560 1945
rect 30600 1930 30615 1945
rect 31190 2225 31220 2235
rect 31190 2205 31195 2225
rect 31215 2205 31220 2225
rect 31520 2225 31550 2235
rect 31520 2205 31525 2225
rect 31545 2205 31550 2225
rect 31850 2225 31880 2235
rect 31850 2205 31855 2225
rect 31875 2205 31880 2225
rect 31190 2190 31240 2205
rect 31225 2180 31240 2190
rect 31280 2190 31790 2205
rect 31280 2180 31295 2190
rect 31335 2180 31350 2190
rect 31390 2180 31405 2190
rect 31445 2180 31460 2190
rect 31500 2180 31515 2190
rect 31555 2180 31570 2190
rect 31610 2180 31625 2190
rect 31665 2180 31680 2190
rect 31720 2180 31735 2190
rect 31775 2180 31790 2190
rect 31830 2190 31880 2205
rect 31920 2225 31950 2235
rect 31920 2205 31925 2225
rect 31945 2205 31950 2225
rect 32250 2225 32280 2235
rect 32250 2205 32255 2225
rect 32275 2205 32280 2225
rect 32580 2225 32610 2235
rect 32580 2205 32585 2225
rect 32605 2205 32610 2225
rect 31920 2190 31970 2205
rect 31830 2180 31845 2190
rect 31955 2180 31970 2190
rect 32010 2190 32520 2205
rect 32010 2180 32025 2190
rect 32065 2180 32080 2190
rect 32120 2180 32135 2190
rect 32175 2180 32190 2190
rect 32230 2180 32245 2190
rect 32285 2180 32300 2190
rect 32340 2180 32355 2190
rect 32395 2180 32410 2190
rect 32450 2180 32465 2190
rect 32505 2180 32520 2190
rect 32560 2190 32610 2205
rect 32560 2180 32575 2190
rect 31225 2015 31240 2030
rect 31280 2015 31295 2030
rect 31335 2015 31350 2030
rect 31390 2015 31405 2030
rect 31445 2015 31460 2030
rect 31500 2015 31515 2030
rect 31555 2015 31570 2030
rect 31610 2015 31625 2030
rect 31665 2015 31680 2030
rect 31720 2015 31735 2030
rect 31775 2015 31790 2030
rect 31830 2015 31845 2030
rect 31955 2015 31970 2030
rect 32010 2015 32025 2030
rect 32065 2015 32080 2030
rect 32120 2015 32135 2030
rect 32175 2015 32190 2030
rect 32230 2015 32245 2030
rect 32285 2015 32300 2030
rect 32340 2015 32355 2030
rect 32395 2015 32410 2030
rect 32450 2015 32465 2030
rect 32505 2015 32520 2030
rect 32560 2015 32575 2030
rect 33150 2290 33180 2300
rect 33150 2270 33155 2290
rect 33175 2270 33180 2290
rect 33313 2290 33347 2300
rect 33313 2270 33321 2290
rect 33339 2270 33347 2290
rect 33810 2290 33840 2300
rect 33810 2270 33815 2290
rect 33835 2270 33840 2290
rect 33150 2255 33200 2270
rect 33185 2245 33200 2255
rect 33240 2255 33750 2270
rect 33240 2245 33255 2255
rect 33295 2245 33310 2255
rect 33350 2245 33365 2255
rect 33405 2245 33420 2255
rect 33460 2245 33475 2255
rect 33515 2245 33530 2255
rect 33570 2245 33585 2255
rect 33625 2245 33640 2255
rect 33680 2245 33695 2255
rect 33735 2245 33750 2255
rect 33790 2255 33840 2270
rect 33790 2245 33805 2255
rect 33185 1930 33200 1945
rect 33240 1930 33255 1945
rect 33295 1930 33310 1945
rect 33350 1930 33365 1945
rect 33405 1930 33420 1945
rect 33460 1930 33475 1945
rect 33515 1930 33530 1945
rect 33570 1930 33585 1945
rect 33625 1930 33640 1945
rect 33680 1930 33695 1945
rect 33735 1930 33750 1945
rect 33790 1930 33805 1945
rect 30040 1700 30070 1710
rect 30040 1680 30045 1700
rect 30065 1680 30070 1700
rect 30438 1700 30472 1710
rect 30438 1680 30446 1700
rect 30464 1680 30472 1700
rect 30640 1700 30670 1710
rect 30640 1680 30645 1700
rect 30665 1680 30670 1700
rect 30040 1665 30135 1680
rect 30075 1655 30135 1665
rect 30175 1665 30535 1680
rect 30175 1655 30235 1665
rect 30275 1655 30335 1665
rect 30375 1655 30435 1665
rect 30475 1655 30535 1665
rect 30575 1665 30670 1680
rect 30575 1655 30635 1665
rect 31035 1755 31065 1765
rect 31035 1735 31040 1755
rect 31060 1735 31065 1755
rect 31237 1755 31269 1765
rect 31237 1735 31243 1755
rect 31260 1735 31269 1755
rect 31457 1755 31489 1765
rect 31457 1735 31463 1755
rect 31480 1735 31489 1755
rect 31035 1720 31085 1735
rect 31180 1725 31269 1735
rect 31400 1725 31489 1735
rect 31601 1755 31635 1765
rect 31601 1735 31610 1755
rect 31627 1735 31635 1755
rect 31695 1755 31725 1765
rect 31695 1735 31700 1755
rect 31720 1735 31725 1755
rect 31601 1725 31635 1735
rect 31070 1710 31085 1720
rect 31125 1710 31140 1725
rect 31180 1720 31250 1725
rect 31180 1710 31195 1720
rect 31235 1710 31250 1720
rect 31290 1710 31305 1725
rect 31345 1710 31360 1725
rect 31400 1720 31470 1725
rect 31400 1710 31415 1720
rect 31455 1710 31470 1720
rect 31510 1710 31525 1725
rect 31565 1710 31580 1725
rect 31620 1710 31635 1725
rect 31675 1720 31725 1735
rect 31775 1755 31805 1765
rect 31775 1735 31780 1755
rect 31800 1735 31805 1755
rect 31867 1755 31899 1765
rect 31867 1740 31873 1755
rect 31865 1735 31873 1740
rect 31890 1735 31899 1755
rect 31995 1755 32025 1765
rect 31995 1735 32000 1755
rect 32020 1735 32025 1755
rect 31775 1720 31825 1735
rect 31675 1710 31690 1720
rect 31810 1710 31825 1720
rect 31865 1725 31899 1735
rect 31865 1710 31880 1725
rect 31920 1710 31935 1725
rect 31975 1720 32025 1735
rect 32075 1755 32105 1765
rect 32075 1735 32080 1755
rect 32100 1735 32105 1755
rect 32277 1755 32309 1765
rect 32277 1735 32283 1755
rect 32300 1735 32309 1755
rect 32497 1755 32529 1765
rect 32497 1735 32503 1755
rect 32520 1735 32529 1755
rect 32075 1720 32125 1735
rect 32220 1725 32309 1735
rect 32440 1725 32529 1735
rect 32641 1755 32675 1765
rect 32641 1735 32650 1755
rect 32667 1735 32675 1755
rect 32735 1755 32765 1765
rect 32735 1735 32740 1755
rect 32760 1735 32765 1755
rect 32641 1725 32675 1735
rect 31975 1710 31990 1720
rect 32110 1710 32125 1720
rect 32165 1710 32180 1725
rect 32220 1720 32290 1725
rect 32220 1710 32235 1720
rect 32275 1710 32290 1720
rect 32330 1710 32345 1725
rect 32385 1710 32400 1725
rect 32440 1720 32510 1725
rect 32440 1710 32455 1720
rect 32495 1710 32510 1720
rect 32550 1710 32565 1725
rect 32605 1710 32620 1725
rect 32660 1710 32675 1725
rect 32715 1720 32765 1735
rect 32715 1710 32730 1720
rect 31070 1545 31085 1560
rect 31125 1545 31140 1560
rect 31180 1545 31195 1560
rect 31235 1545 31250 1560
rect 31290 1550 31305 1560
rect 31345 1550 31360 1560
rect 31106 1535 31140 1545
rect 31290 1535 31360 1550
rect 31400 1545 31415 1560
rect 31455 1545 31470 1560
rect 31510 1550 31525 1560
rect 31565 1550 31580 1560
rect 31510 1535 31580 1550
rect 31620 1545 31635 1560
rect 31675 1545 31690 1560
rect 31810 1545 31825 1560
rect 31865 1545 31880 1560
rect 31920 1545 31935 1560
rect 31975 1545 31990 1560
rect 32110 1545 32125 1560
rect 32165 1545 32180 1560
rect 32220 1545 32235 1560
rect 32275 1545 32290 1560
rect 32330 1550 32345 1560
rect 32385 1550 32400 1560
rect 31920 1535 31954 1545
rect 31106 1515 31112 1535
rect 31129 1515 31138 1535
rect 31106 1505 31138 1515
rect 31305 1515 31315 1535
rect 31335 1515 31345 1535
rect 31305 1505 31345 1515
rect 31525 1515 31535 1535
rect 31555 1515 31565 1535
rect 31525 1505 31565 1515
rect 31922 1515 31928 1535
rect 31945 1515 31954 1535
rect 31922 1505 31954 1515
rect 32146 1535 32180 1545
rect 32330 1535 32400 1550
rect 32440 1545 32455 1560
rect 32495 1545 32510 1560
rect 32550 1550 32565 1560
rect 32605 1550 32620 1560
rect 32550 1535 32620 1550
rect 32660 1545 32675 1560
rect 32715 1545 32730 1560
rect 32146 1515 32152 1535
rect 32169 1515 32178 1535
rect 32146 1505 32178 1515
rect 32345 1515 32355 1535
rect 32375 1515 32385 1535
rect 32345 1505 32385 1515
rect 32565 1515 32575 1535
rect 32595 1515 32605 1535
rect 32565 1505 32605 1515
rect 33130 1700 33160 1710
rect 33130 1680 33135 1700
rect 33155 1680 33160 1700
rect 33328 1700 33362 1710
rect 33328 1680 33336 1700
rect 33354 1680 33362 1700
rect 33730 1700 33760 1710
rect 33730 1680 33735 1700
rect 33755 1680 33760 1700
rect 33130 1665 33225 1680
rect 33165 1655 33225 1665
rect 33265 1665 33625 1680
rect 33265 1655 33325 1665
rect 33365 1655 33425 1665
rect 33465 1655 33525 1665
rect 33565 1655 33625 1665
rect 33665 1665 33760 1680
rect 33665 1655 33725 1665
rect 30075 940 30135 955
rect 30175 940 30235 955
rect 30275 940 30335 955
rect 30375 940 30435 955
rect 30475 940 30535 955
rect 30575 940 30635 955
rect 31815 1250 31845 1260
rect 31815 1230 31820 1250
rect 31840 1230 31845 1250
rect 32381 1250 32411 1260
rect 32381 1230 32386 1250
rect 32406 1235 32411 1250
rect 32406 1230 32415 1235
rect 31245 1205 31260 1220
rect 31300 1215 32360 1230
rect 32381 1220 32415 1230
rect 31300 1205 31315 1215
rect 31355 1205 31370 1215
rect 31410 1205 31425 1215
rect 31465 1205 31480 1215
rect 31520 1205 31535 1215
rect 31575 1205 31590 1215
rect 31630 1205 31645 1215
rect 31685 1205 31700 1215
rect 31740 1205 31755 1215
rect 31795 1205 31810 1215
rect 31850 1205 31865 1215
rect 31905 1205 31920 1215
rect 31960 1205 31975 1215
rect 32015 1205 32030 1215
rect 32070 1205 32085 1215
rect 32125 1205 32140 1215
rect 32180 1205 32195 1215
rect 32235 1205 32250 1215
rect 32290 1205 32305 1215
rect 32345 1205 32360 1215
rect 32400 1205 32415 1220
rect 32455 1205 32470 1220
rect 31245 940 31260 955
rect 31300 940 31315 955
rect 31355 940 31370 955
rect 31410 940 31425 955
rect 31465 940 31480 955
rect 31520 940 31535 955
rect 31575 940 31590 955
rect 31630 940 31645 955
rect 31685 940 31700 955
rect 31740 940 31755 955
rect 31795 940 31810 955
rect 31850 940 31865 955
rect 31905 940 31920 955
rect 31960 940 31975 955
rect 32015 940 32030 955
rect 32070 940 32085 955
rect 32125 940 32140 955
rect 32180 940 32195 955
rect 32235 940 32250 955
rect 32290 940 32305 955
rect 32345 940 32360 955
rect 32400 940 32415 955
rect 32455 940 32470 955
rect 31195 930 31260 940
rect 31195 910 31205 930
rect 31225 925 31260 930
rect 32455 930 32515 940
rect 32455 925 32485 930
rect 31225 910 31235 925
rect 31195 900 31235 910
rect 32475 910 32485 925
rect 32505 910 32515 930
rect 32475 900 32515 910
rect 33165 940 33225 955
rect 33265 940 33325 955
rect 33365 940 33425 955
rect 33465 940 33525 955
rect 33565 940 33625 955
rect 33665 940 33725 955
rect 31305 735 31345 745
rect 31305 715 31315 735
rect 31335 715 31345 735
rect 31305 705 31345 715
rect 31375 735 31415 745
rect 31375 715 31385 735
rect 31405 715 31415 735
rect 31375 705 31415 715
rect 31445 735 31485 745
rect 31445 715 31455 735
rect 31475 715 31485 735
rect 31445 705 31485 715
rect 31300 690 31490 705
rect 31300 575 31490 590
rect 31885 730 31915 740
rect 31885 710 31890 730
rect 31910 710 31915 730
rect 32155 730 32195 740
rect 32155 710 32165 730
rect 32185 710 32195 730
rect 32375 730 32415 740
rect 32375 710 32385 730
rect 32405 710 32415 730
rect 32545 730 32575 740
rect 32545 710 32550 730
rect 32570 710 32575 730
rect 31885 695 31935 710
rect 31920 685 31935 695
rect 31975 695 32485 710
rect 31975 685 31990 695
rect 32030 685 32045 695
rect 32085 685 32100 695
rect 32140 685 32155 695
rect 32195 685 32210 695
rect 32250 685 32265 695
rect 32305 685 32320 695
rect 32360 685 32375 695
rect 32415 685 32430 695
rect 32470 685 32485 695
rect 32525 695 32575 710
rect 32525 685 32540 695
rect 31920 620 31935 635
rect 31975 620 31990 635
rect 32030 620 32045 635
rect 32085 620 32100 635
rect 32140 620 32155 635
rect 32195 620 32210 635
rect 32250 620 32265 635
rect 32305 620 32320 635
rect 32360 620 32375 635
rect 32415 620 32430 635
rect 32470 620 32485 635
rect 32525 620 32540 635
<< polycont >>
rect 31840 4860 31860 4880
rect 31230 4710 31250 4730
rect 31320 4710 31340 4730
rect 31410 4710 31430 4730
rect 31480 4710 31500 4730
rect 31660 4705 31680 4725
rect 31840 4710 31860 4730
rect 32210 4705 32230 4725
rect 32331 4705 32349 4725
rect 32690 4705 32710 4725
rect 31260 4295 31280 4315
rect 31370 4295 31390 4315
rect 32470 4295 32490 4315
rect 31285 4005 31305 4025
rect 31485 4005 31505 4025
rect 31705 4005 31725 4025
rect 32013 4005 32033 4025
rect 32215 4005 32235 4025
rect 32435 4005 32455 4025
rect 31210 3885 31230 3905
rect 31413 3885 31430 3905
rect 31633 3885 31650 3905
rect 31780 3885 31797 3905
rect 31870 3885 31890 3905
rect 31940 3885 31960 3905
rect 32143 3885 32160 3905
rect 32363 3885 32380 3905
rect 32510 3885 32527 3905
rect 32600 3885 32620 3905
rect 29965 3020 29985 3040
rect 30186 3020 30204 3040
rect 30625 3020 30645 3040
rect 31230 3160 31250 3180
rect 31831 3160 31849 3180
rect 32550 3160 32570 3180
rect 33155 3020 33175 3040
rect 33596 3020 33614 3040
rect 33815 3020 33835 3040
rect 29965 2460 29985 2480
rect 30461 2460 30479 2480
rect 30625 2460 30645 2480
rect 31015 2450 31035 2470
rect 31376 2450 31394 2470
rect 31735 2450 31755 2470
rect 32045 2450 32065 2470
rect 32406 2450 32424 2470
rect 32765 2450 32785 2470
rect 33155 2460 33175 2480
rect 33321 2460 33339 2480
rect 33815 2460 33835 2480
rect 29965 2270 29985 2290
rect 30461 2270 30479 2290
rect 30625 2270 30645 2290
rect 31195 2205 31215 2225
rect 31525 2205 31545 2225
rect 31855 2205 31875 2225
rect 31925 2205 31945 2225
rect 32255 2205 32275 2225
rect 32585 2205 32605 2225
rect 33155 2270 33175 2290
rect 33321 2270 33339 2290
rect 33815 2270 33835 2290
rect 30045 1680 30065 1700
rect 30446 1680 30464 1700
rect 30645 1680 30665 1700
rect 31040 1735 31060 1755
rect 31243 1735 31260 1755
rect 31463 1735 31480 1755
rect 31610 1735 31627 1755
rect 31700 1735 31720 1755
rect 31780 1735 31800 1755
rect 31873 1735 31890 1755
rect 32000 1735 32020 1755
rect 32080 1735 32100 1755
rect 32283 1735 32300 1755
rect 32503 1735 32520 1755
rect 32650 1735 32667 1755
rect 32740 1735 32760 1755
rect 31112 1515 31129 1535
rect 31315 1515 31335 1535
rect 31535 1515 31555 1535
rect 31928 1515 31945 1535
rect 32152 1515 32169 1535
rect 32355 1515 32375 1535
rect 32575 1515 32595 1535
rect 33135 1680 33155 1700
rect 33336 1680 33354 1700
rect 33735 1680 33755 1700
rect 31820 1230 31840 1250
rect 32386 1230 32406 1250
rect 31205 910 31225 930
rect 32485 910 32505 930
rect 31315 715 31335 735
rect 31385 715 31405 735
rect 31455 715 31475 735
rect 31890 710 31910 730
rect 32165 710 32185 730
rect 32385 710 32405 730
rect 32550 710 32570 730
<< xpolycontact >>
rect 29554 3400 29695 3620
rect 29554 3055 29695 3275
rect 34105 3400 34246 3620
rect 34105 3055 34246 3275
rect 29470 2369 29505 2589
rect 29470 1990 29505 2210
rect 29530 2369 29565 2589
rect 29530 1990 29565 2210
rect 29590 2369 29625 2589
rect 29590 1990 29625 2210
rect 29650 2369 29685 2589
rect 29650 1990 29685 2210
rect 34115 2369 34150 2589
rect 34115 1990 34150 2210
rect 34175 2369 34210 2589
rect 34175 1990 34210 2210
rect 34235 2369 34270 2589
rect 34235 1990 34270 2210
rect 34295 2369 34330 2589
rect 34295 1990 34330 2210
rect 29730 1385 29765 1605
rect 29730 918 29765 1138
rect 29790 1385 29825 1605
rect 29790 918 29825 1138
rect 33975 1385 34010 1605
rect 33975 918 34010 1138
rect 34035 1385 34070 1605
rect 34035 918 34070 1138
<< ppolyres >>
rect 29554 3275 29695 3400
rect 34105 3275 34246 3400
<< xpolyres >>
rect 29470 2210 29505 2369
rect 29530 2210 29565 2369
rect 29590 2210 29625 2369
rect 29650 2210 29685 2369
rect 34115 2210 34150 2369
rect 34175 2210 34210 2369
rect 34235 2210 34270 2369
rect 34295 2210 34330 2369
rect 29730 1138 29765 1385
rect 29790 1138 29825 1385
rect 33975 1138 34010 1385
rect 34035 1138 34070 1385
<< locali >>
rect 31170 4910 31485 4930
rect 31565 4910 31920 4930
rect 31170 4825 31190 4910
rect 31470 4880 31510 4890
rect 31280 4865 31320 4875
rect 31280 4845 31290 4865
rect 31310 4845 31320 4865
rect 31470 4860 31480 4880
rect 31500 4860 31510 4880
rect 31470 4850 31510 4860
rect 31537 4880 31563 4890
rect 31537 4860 31540 4880
rect 31560 4860 31563 4880
rect 31537 4850 31563 4860
rect 31590 4880 31630 4890
rect 31590 4860 31600 4880
rect 31620 4860 31630 4880
rect 31590 4850 31630 4860
rect 31657 4880 31683 4890
rect 31657 4860 31660 4880
rect 31680 4860 31683 4880
rect 31657 4850 31683 4860
rect 31710 4880 31750 4890
rect 31710 4860 31720 4880
rect 31740 4860 31750 4880
rect 31710 4850 31750 4860
rect 31777 4880 31803 4890
rect 31777 4860 31780 4880
rect 31800 4860 31803 4880
rect 31777 4850 31803 4860
rect 31830 4880 31870 4890
rect 31830 4860 31840 4880
rect 31860 4860 31870 4880
rect 31830 4850 31870 4860
rect 31280 4835 31320 4845
rect 31290 4813 31310 4835
rect 31480 4830 31500 4850
rect 31540 4830 31560 4850
rect 31600 4830 31620 4850
rect 31660 4830 31680 4850
rect 31720 4830 31740 4850
rect 31780 4830 31800 4850
rect 31840 4830 31860 4850
rect 31170 4675 31190 4745
rect 31225 4795 31255 4813
rect 31225 4775 31230 4795
rect 31250 4775 31255 4795
rect 31225 4730 31255 4775
rect 31285 4795 31315 4813
rect 31285 4775 31290 4795
rect 31310 4775 31315 4795
rect 31285 4760 31315 4775
rect 31345 4795 31375 4813
rect 31345 4775 31350 4795
rect 31370 4775 31375 4795
rect 31345 4760 31375 4775
rect 31405 4795 31435 4813
rect 31405 4775 31410 4795
rect 31430 4775 31435 4795
rect 31350 4740 31370 4760
rect 31225 4710 31230 4730
rect 31250 4710 31255 4730
rect 31225 4700 31255 4710
rect 31310 4730 31370 4740
rect 31310 4710 31320 4730
rect 31340 4720 31370 4730
rect 31405 4730 31435 4775
rect 31340 4710 31350 4720
rect 31310 4700 31350 4710
rect 31405 4710 31410 4730
rect 31430 4710 31435 4730
rect 31405 4700 31435 4710
rect 31475 4805 31505 4830
rect 31475 4785 31480 4805
rect 31500 4785 31505 4805
rect 31475 4730 31505 4785
rect 31535 4805 31565 4830
rect 31535 4785 31540 4805
rect 31560 4785 31565 4805
rect 31535 4760 31565 4785
rect 31595 4805 31625 4830
rect 31595 4785 31600 4805
rect 31620 4785 31625 4805
rect 31595 4760 31625 4785
rect 31655 4805 31685 4830
rect 31655 4785 31660 4805
rect 31680 4785 31685 4805
rect 31655 4760 31685 4785
rect 31715 4805 31745 4830
rect 31715 4785 31720 4805
rect 31740 4785 31745 4805
rect 31715 4760 31745 4785
rect 31775 4805 31805 4830
rect 31775 4785 31780 4805
rect 31800 4785 31805 4805
rect 31775 4760 31805 4785
rect 31835 4805 31865 4830
rect 31835 4785 31840 4805
rect 31860 4785 31865 4805
rect 31475 4710 31480 4730
rect 31500 4710 31505 4730
rect 31475 4700 31505 4710
rect 31650 4725 31690 4735
rect 31650 4705 31660 4725
rect 31680 4705 31690 4725
rect 31230 4675 31250 4700
rect 31410 4675 31430 4700
rect 31480 4675 31500 4700
rect 31650 4695 31690 4705
rect 31835 4730 31865 4785
rect 31835 4710 31840 4730
rect 31860 4710 31865 4730
rect 31835 4700 31865 4710
rect 31900 4825 31920 4910
rect 31840 4675 31860 4700
rect 31900 4675 31920 4745
rect 31170 4655 31485 4675
rect 31565 4655 31920 4675
rect 32150 4885 32420 4905
rect 32500 4885 32770 4905
rect 32150 4820 32170 4885
rect 32200 4855 32240 4865
rect 32200 4835 32210 4855
rect 32230 4835 32240 4855
rect 32200 4825 32240 4835
rect 32320 4855 32360 4865
rect 32320 4835 32330 4855
rect 32350 4835 32360 4855
rect 32320 4825 32360 4835
rect 32440 4855 32480 4865
rect 32440 4835 32450 4855
rect 32470 4835 32480 4855
rect 32440 4825 32480 4835
rect 32560 4855 32600 4865
rect 32560 4835 32570 4855
rect 32590 4835 32600 4855
rect 32560 4825 32600 4835
rect 32680 4855 32720 4865
rect 32680 4835 32690 4855
rect 32710 4835 32720 4855
rect 32680 4825 32720 4835
rect 32750 4825 32770 4885
rect 32210 4805 32230 4825
rect 32330 4805 32350 4825
rect 32450 4805 32470 4825
rect 32570 4805 32590 4825
rect 32690 4805 32710 4825
rect 32150 4675 32170 4740
rect 32205 4790 32235 4805
rect 32205 4770 32210 4790
rect 32230 4770 32235 4790
rect 32205 4725 32235 4770
rect 32265 4790 32295 4805
rect 32265 4770 32270 4790
rect 32290 4770 32295 4790
rect 32265 4755 32295 4770
rect 32325 4790 32355 4805
rect 32325 4770 32330 4790
rect 32350 4770 32355 4790
rect 32325 4755 32355 4770
rect 32385 4790 32415 4805
rect 32385 4770 32390 4790
rect 32410 4770 32415 4790
rect 32385 4755 32415 4770
rect 32445 4790 32475 4805
rect 32445 4770 32450 4790
rect 32470 4770 32475 4790
rect 32445 4755 32475 4770
rect 32505 4790 32535 4805
rect 32505 4770 32510 4790
rect 32530 4770 32535 4790
rect 32505 4755 32535 4770
rect 32565 4790 32595 4805
rect 32565 4770 32570 4790
rect 32590 4770 32595 4790
rect 32565 4755 32595 4770
rect 32625 4790 32655 4805
rect 32625 4770 32630 4790
rect 32650 4770 32655 4790
rect 32625 4755 32655 4770
rect 32685 4790 32715 4805
rect 32685 4770 32690 4790
rect 32710 4770 32715 4790
rect 32270 4735 32290 4755
rect 32390 4735 32410 4755
rect 32510 4735 32530 4755
rect 32630 4735 32650 4755
rect 32205 4705 32210 4725
rect 32230 4705 32235 4725
rect 32205 4695 32235 4705
rect 32260 4725 32300 4735
rect 32260 4705 32270 4725
rect 32290 4705 32300 4725
rect 32260 4695 32300 4705
rect 32323 4725 32357 4735
rect 32323 4705 32331 4725
rect 32349 4705 32357 4725
rect 32323 4695 32357 4705
rect 32380 4725 32420 4735
rect 32380 4705 32390 4725
rect 32410 4705 32420 4725
rect 32380 4695 32420 4705
rect 32500 4725 32540 4735
rect 32500 4705 32510 4725
rect 32530 4705 32540 4725
rect 32500 4695 32540 4705
rect 32620 4725 32660 4735
rect 32620 4705 32630 4725
rect 32650 4705 32660 4725
rect 32620 4695 32660 4705
rect 32685 4725 32715 4770
rect 32685 4705 32690 4725
rect 32710 4705 32715 4725
rect 32685 4695 32715 4705
rect 32210 4675 32230 4695
rect 32690 4675 32710 4695
rect 32750 4675 32770 4740
rect 32150 4655 32420 4675
rect 32500 4655 32770 4675
rect 31200 4465 31835 4485
rect 31915 4465 32550 4485
rect 31200 4405 31220 4465
rect 31250 4435 31290 4445
rect 31250 4415 31260 4435
rect 31280 4415 31290 4435
rect 31250 4405 31290 4415
rect 31360 4435 31400 4445
rect 31360 4415 31370 4435
rect 31390 4415 31400 4435
rect 31360 4405 31400 4415
rect 31470 4435 31510 4445
rect 31470 4415 31480 4435
rect 31500 4415 31510 4435
rect 31470 4405 31510 4415
rect 31580 4435 31620 4445
rect 31580 4415 31590 4435
rect 31610 4415 31620 4435
rect 31580 4405 31620 4415
rect 31690 4435 31730 4445
rect 31690 4415 31700 4435
rect 31720 4415 31730 4435
rect 31690 4405 31730 4415
rect 31800 4435 31840 4445
rect 31800 4415 31810 4435
rect 31830 4415 31840 4435
rect 31800 4405 31840 4415
rect 31910 4435 31950 4445
rect 31910 4415 31920 4435
rect 31940 4415 31950 4435
rect 31910 4405 31950 4415
rect 32020 4435 32060 4445
rect 32020 4415 32030 4435
rect 32050 4415 32060 4435
rect 32020 4405 32060 4415
rect 32130 4435 32170 4445
rect 32130 4415 32140 4435
rect 32160 4415 32170 4435
rect 32130 4405 32170 4415
rect 32240 4435 32280 4445
rect 32240 4415 32250 4435
rect 32270 4415 32280 4435
rect 32240 4405 32280 4415
rect 32350 4435 32390 4445
rect 32350 4415 32360 4435
rect 32380 4415 32390 4435
rect 32350 4405 32390 4415
rect 32460 4435 32500 4445
rect 32460 4415 32470 4435
rect 32490 4415 32500 4435
rect 32460 4405 32500 4415
rect 32530 4405 32550 4465
rect 31260 4385 31280 4405
rect 31370 4385 31390 4405
rect 31480 4385 31500 4405
rect 31590 4385 31610 4405
rect 31700 4385 31720 4405
rect 31810 4385 31830 4405
rect 31920 4385 31940 4405
rect 32030 4385 32050 4405
rect 32140 4385 32160 4405
rect 32250 4385 32270 4405
rect 32360 4385 32380 4405
rect 32470 4385 32490 4405
rect 31200 4265 31220 4325
rect 31255 4375 31285 4385
rect 31255 4355 31260 4375
rect 31280 4355 31285 4375
rect 31255 4315 31285 4355
rect 31310 4375 31340 4385
rect 31310 4355 31315 4375
rect 31335 4355 31340 4375
rect 31310 4345 31340 4355
rect 31365 4375 31395 4385
rect 31365 4355 31370 4375
rect 31390 4355 31395 4375
rect 31365 4345 31395 4355
rect 31420 4375 31450 4385
rect 31420 4355 31425 4375
rect 31445 4355 31450 4375
rect 31420 4345 31450 4355
rect 31475 4375 31505 4385
rect 31475 4355 31480 4375
rect 31500 4355 31505 4375
rect 31475 4345 31505 4355
rect 31530 4375 31560 4385
rect 31530 4355 31535 4375
rect 31555 4355 31560 4375
rect 31530 4345 31560 4355
rect 31585 4375 31615 4385
rect 31585 4355 31590 4375
rect 31610 4355 31615 4375
rect 31585 4345 31615 4355
rect 31640 4375 31670 4385
rect 31640 4355 31645 4375
rect 31665 4355 31670 4375
rect 31640 4345 31670 4355
rect 31695 4375 31725 4385
rect 31695 4355 31700 4375
rect 31720 4355 31725 4375
rect 31695 4345 31725 4355
rect 31750 4375 31780 4385
rect 31750 4355 31755 4375
rect 31775 4355 31780 4375
rect 31750 4345 31780 4355
rect 31805 4375 31835 4385
rect 31805 4355 31810 4375
rect 31830 4355 31835 4375
rect 31805 4345 31835 4355
rect 31860 4375 31890 4385
rect 31860 4355 31865 4375
rect 31885 4355 31890 4375
rect 31860 4345 31890 4355
rect 31915 4375 31945 4385
rect 31915 4355 31920 4375
rect 31940 4355 31945 4375
rect 31915 4345 31945 4355
rect 31970 4375 32000 4385
rect 31970 4355 31975 4375
rect 31995 4355 32000 4375
rect 31970 4345 32000 4355
rect 32025 4375 32055 4385
rect 32025 4355 32030 4375
rect 32050 4355 32055 4375
rect 32025 4345 32055 4355
rect 32080 4375 32110 4385
rect 32080 4355 32085 4375
rect 32105 4355 32110 4375
rect 32080 4345 32110 4355
rect 32135 4375 32165 4385
rect 32135 4355 32140 4375
rect 32160 4355 32165 4375
rect 32135 4345 32165 4355
rect 32190 4375 32220 4385
rect 32190 4355 32195 4375
rect 32215 4355 32220 4375
rect 32190 4345 32220 4355
rect 32245 4375 32275 4385
rect 32245 4355 32250 4375
rect 32270 4355 32275 4375
rect 32245 4345 32275 4355
rect 32300 4375 32330 4385
rect 32300 4355 32305 4375
rect 32325 4355 32330 4375
rect 32300 4345 32330 4355
rect 32355 4375 32385 4385
rect 32355 4355 32360 4375
rect 32380 4355 32385 4375
rect 32355 4345 32385 4355
rect 32410 4375 32440 4385
rect 32410 4355 32415 4375
rect 32435 4355 32440 4375
rect 32410 4345 32440 4355
rect 32465 4375 32495 4385
rect 32465 4355 32470 4375
rect 32490 4355 32495 4375
rect 31315 4325 31335 4345
rect 31425 4325 31445 4345
rect 31535 4325 31555 4345
rect 31645 4325 31665 4345
rect 31755 4325 31775 4345
rect 31865 4325 31885 4345
rect 31975 4325 31995 4345
rect 32085 4325 32105 4345
rect 32195 4325 32215 4345
rect 32305 4325 32325 4345
rect 32415 4325 32435 4345
rect 31255 4295 31260 4315
rect 31280 4295 31285 4315
rect 31255 4285 31285 4295
rect 31305 4315 31345 4325
rect 31305 4295 31315 4315
rect 31335 4295 31345 4315
rect 31305 4285 31345 4295
rect 31362 4315 31398 4325
rect 31362 4295 31370 4315
rect 31390 4295 31398 4315
rect 31362 4285 31398 4295
rect 31415 4315 31455 4325
rect 31415 4295 31425 4315
rect 31445 4295 31455 4315
rect 31415 4285 31455 4295
rect 31525 4315 31565 4325
rect 31525 4295 31535 4315
rect 31555 4295 31565 4315
rect 31525 4285 31565 4295
rect 31635 4315 31675 4325
rect 31635 4295 31645 4315
rect 31665 4295 31675 4315
rect 31635 4285 31675 4295
rect 31745 4315 31785 4325
rect 31745 4295 31755 4315
rect 31775 4295 31785 4315
rect 31745 4285 31785 4295
rect 31855 4315 31895 4325
rect 31855 4295 31865 4315
rect 31885 4295 31895 4315
rect 31855 4285 31895 4295
rect 31965 4315 32005 4325
rect 31965 4295 31975 4315
rect 31995 4295 32005 4315
rect 31965 4285 32005 4295
rect 32075 4315 32115 4325
rect 32075 4295 32085 4315
rect 32105 4295 32115 4315
rect 32075 4285 32115 4295
rect 32185 4315 32225 4325
rect 32185 4295 32195 4315
rect 32215 4295 32225 4315
rect 32185 4285 32225 4295
rect 32295 4315 32335 4325
rect 32295 4295 32305 4315
rect 32325 4295 32335 4315
rect 32295 4285 32335 4295
rect 32405 4315 32445 4325
rect 32405 4295 32415 4315
rect 32435 4295 32445 4315
rect 32405 4285 32445 4295
rect 32465 4315 32495 4355
rect 32465 4295 32470 4315
rect 32490 4295 32495 4315
rect 32465 4285 32495 4295
rect 31260 4265 31280 4285
rect 32470 4265 32490 4285
rect 32530 4265 32550 4325
rect 31200 4245 31835 4265
rect 31915 4245 32550 4265
rect 31635 4170 31675 4210
rect 31855 4170 31895 4210
rect 32075 4170 32115 4210
rect 32295 4170 32335 4210
rect 31150 4055 31875 4075
rect 31955 4055 32680 4075
rect 31150 3995 31170 4055
rect 31280 4025 31310 4035
rect 31280 4005 31285 4025
rect 31305 4005 31310 4025
rect 31280 3995 31310 4005
rect 31327 4025 31353 4035
rect 31327 4005 31330 4025
rect 31350 4005 31353 4025
rect 31327 3995 31353 4005
rect 31370 4025 31400 4035
rect 31370 4005 31375 4025
rect 31395 4005 31400 4025
rect 31370 3995 31400 4005
rect 31427 4025 31453 4035
rect 31427 4005 31430 4025
rect 31450 4005 31453 4025
rect 31427 3995 31453 4005
rect 31480 4025 31510 4035
rect 31480 4005 31485 4025
rect 31505 4005 31510 4025
rect 31480 3995 31510 4005
rect 31537 4025 31563 4035
rect 31537 4005 31540 4025
rect 31560 4005 31563 4025
rect 31537 3995 31563 4005
rect 31647 4025 31673 4035
rect 31647 4005 31650 4025
rect 31670 4005 31673 4025
rect 31647 3995 31673 4005
rect 31695 4025 31735 4035
rect 31695 4005 31705 4025
rect 31725 4005 31735 4025
rect 31695 3995 31735 4005
rect 31757 4025 31783 4035
rect 31757 4005 31760 4025
rect 31780 4005 31783 4025
rect 31757 3995 31783 4005
rect 32008 4025 32038 4035
rect 32008 4005 32013 4025
rect 32033 4005 32038 4025
rect 32008 3995 32038 4005
rect 32057 4025 32083 4035
rect 32057 4005 32060 4025
rect 32080 4005 32083 4025
rect 32057 3995 32083 4005
rect 32157 4025 32183 4035
rect 32157 4005 32160 4025
rect 32180 4005 32183 4025
rect 32157 3995 32183 4005
rect 32205 4025 32245 4035
rect 32205 4005 32215 4025
rect 32235 4005 32245 4025
rect 32205 3995 32245 4005
rect 32267 4025 32293 4035
rect 32267 4005 32270 4025
rect 32290 4005 32293 4025
rect 32267 3995 32293 4005
rect 32377 4025 32403 4035
rect 32377 4005 32380 4025
rect 32400 4005 32403 4025
rect 32377 3995 32403 4005
rect 32425 4025 32465 4035
rect 32425 4005 32435 4025
rect 32455 4005 32465 4025
rect 32425 3995 32465 4005
rect 32487 4025 32513 4035
rect 32487 4005 32490 4025
rect 32510 4005 32513 4025
rect 32487 3995 32513 4005
rect 32660 3995 32680 4055
rect 32875 4000 32905 4030
rect 31140 3935 31150 3975
rect 31327 3975 31345 3995
rect 31375 3975 31395 3995
rect 31430 3975 31450 3995
rect 31540 3975 31560 3995
rect 31650 3975 31670 3995
rect 31760 3975 31780 3995
rect 32057 3975 32075 3995
rect 32160 3975 32180 3995
rect 32270 3975 32290 3995
rect 32380 3975 32400 3995
rect 32490 3975 32510 3995
rect 31170 3935 31180 3975
rect 31205 3965 31235 3975
rect 31205 3945 31210 3965
rect 31230 3945 31235 3965
rect 31150 3855 31170 3915
rect 31205 3905 31235 3945
rect 31260 3965 31290 3975
rect 31260 3945 31265 3965
rect 31285 3945 31290 3965
rect 31260 3935 31290 3945
rect 31315 3965 31345 3975
rect 31315 3945 31320 3965
rect 31340 3945 31345 3965
rect 31315 3935 31345 3945
rect 31370 3965 31400 3975
rect 31370 3945 31375 3965
rect 31395 3945 31400 3965
rect 31370 3935 31400 3945
rect 31425 3965 31455 3975
rect 31425 3945 31430 3965
rect 31450 3945 31455 3965
rect 31425 3935 31455 3945
rect 31480 3965 31510 3975
rect 31480 3945 31485 3965
rect 31505 3945 31510 3965
rect 31480 3935 31510 3945
rect 31535 3965 31565 3975
rect 31535 3945 31540 3965
rect 31560 3945 31565 3965
rect 31535 3935 31565 3945
rect 31590 3965 31620 3975
rect 31590 3945 31595 3965
rect 31615 3945 31620 3965
rect 31590 3935 31620 3945
rect 31645 3965 31675 3975
rect 31645 3945 31650 3965
rect 31670 3945 31675 3965
rect 31645 3935 31675 3945
rect 31700 3965 31730 3975
rect 31700 3945 31705 3965
rect 31725 3945 31730 3965
rect 31700 3935 31730 3945
rect 31755 3965 31785 3975
rect 31755 3945 31760 3965
rect 31780 3945 31785 3965
rect 31755 3935 31785 3945
rect 31810 3965 31840 3975
rect 31810 3945 31815 3965
rect 31835 3945 31840 3965
rect 31810 3935 31840 3945
rect 31265 3915 31285 3935
rect 31370 3915 31390 3935
rect 31485 3915 31505 3935
rect 31590 3915 31610 3935
rect 31705 3915 31725 3935
rect 31820 3915 31840 3935
rect 31865 3965 31895 3975
rect 31865 3945 31870 3965
rect 31890 3945 31895 3965
rect 31205 3885 31210 3905
rect 31230 3885 31235 3905
rect 31205 3875 31235 3885
rect 31255 3905 31295 3915
rect 31255 3885 31265 3905
rect 31285 3885 31295 3905
rect 31255 3875 31295 3885
rect 31350 3905 31390 3915
rect 31350 3885 31360 3905
rect 31380 3885 31390 3905
rect 31350 3875 31390 3885
rect 31407 3905 31439 3915
rect 31407 3885 31413 3905
rect 31430 3885 31439 3905
rect 31407 3875 31439 3885
rect 31475 3905 31515 3915
rect 31475 3885 31485 3905
rect 31505 3885 31515 3905
rect 31475 3875 31515 3885
rect 31570 3905 31610 3915
rect 31570 3885 31580 3905
rect 31600 3885 31610 3905
rect 31570 3875 31610 3885
rect 31627 3905 31659 3915
rect 31627 3885 31633 3905
rect 31650 3885 31659 3905
rect 31627 3875 31659 3885
rect 31695 3905 31735 3915
rect 31695 3885 31705 3905
rect 31725 3885 31735 3905
rect 31695 3875 31735 3885
rect 31771 3905 31803 3915
rect 31771 3885 31780 3905
rect 31797 3885 31803 3905
rect 31771 3875 31803 3885
rect 31820 3905 31846 3915
rect 31820 3885 31823 3905
rect 31843 3885 31846 3905
rect 31820 3875 31846 3885
rect 31865 3905 31895 3945
rect 31865 3885 31870 3905
rect 31890 3885 31895 3905
rect 31865 3875 31895 3885
rect 31935 3965 31965 3975
rect 31935 3945 31940 3965
rect 31960 3945 31965 3965
rect 31935 3905 31965 3945
rect 31990 3965 32020 3975
rect 31990 3945 31995 3965
rect 32015 3945 32020 3965
rect 31990 3935 32020 3945
rect 32045 3965 32075 3975
rect 32045 3945 32050 3965
rect 32070 3945 32075 3965
rect 32045 3935 32075 3945
rect 32100 3965 32130 3975
rect 32100 3945 32105 3965
rect 32125 3945 32130 3965
rect 32100 3935 32130 3945
rect 32155 3965 32185 3975
rect 32155 3945 32160 3965
rect 32180 3945 32185 3965
rect 32155 3935 32185 3945
rect 32210 3965 32240 3975
rect 32210 3945 32215 3965
rect 32235 3945 32240 3965
rect 32210 3935 32240 3945
rect 32265 3965 32295 3975
rect 32265 3945 32270 3965
rect 32290 3945 32295 3965
rect 32265 3935 32295 3945
rect 32320 3965 32350 3975
rect 32320 3945 32325 3965
rect 32345 3945 32350 3965
rect 32320 3935 32350 3945
rect 32375 3965 32405 3975
rect 32375 3945 32380 3965
rect 32400 3945 32405 3965
rect 32375 3935 32405 3945
rect 32430 3965 32460 3975
rect 32430 3945 32435 3965
rect 32455 3945 32460 3965
rect 32430 3935 32460 3945
rect 32485 3965 32515 3975
rect 32485 3945 32490 3965
rect 32510 3945 32515 3965
rect 32485 3935 32515 3945
rect 32540 3965 32570 3975
rect 32540 3945 32545 3965
rect 32565 3945 32570 3965
rect 32540 3935 32570 3945
rect 31995 3915 32015 3935
rect 32100 3915 32120 3935
rect 32215 3915 32235 3935
rect 32320 3915 32340 3935
rect 32435 3915 32455 3935
rect 32550 3915 32570 3935
rect 32595 3965 32625 3975
rect 32595 3945 32600 3965
rect 32620 3945 32625 3965
rect 31935 3885 31940 3905
rect 31960 3885 31965 3905
rect 31935 3875 31965 3885
rect 31985 3905 32025 3915
rect 31985 3885 31995 3905
rect 32015 3885 32025 3905
rect 31985 3875 32025 3885
rect 32080 3905 32120 3915
rect 32080 3885 32090 3905
rect 32110 3885 32120 3905
rect 32080 3875 32120 3885
rect 32137 3905 32169 3915
rect 32137 3885 32143 3905
rect 32160 3885 32169 3905
rect 32137 3875 32169 3885
rect 32205 3905 32245 3915
rect 32205 3885 32215 3905
rect 32235 3885 32245 3905
rect 32205 3875 32245 3885
rect 32300 3905 32340 3915
rect 32300 3885 32310 3905
rect 32330 3885 32340 3905
rect 32300 3875 32340 3885
rect 32357 3905 32389 3915
rect 32357 3885 32363 3905
rect 32380 3885 32389 3905
rect 32357 3875 32389 3885
rect 32425 3905 32465 3915
rect 32425 3885 32435 3905
rect 32455 3885 32465 3905
rect 32425 3875 32465 3885
rect 32501 3905 32533 3915
rect 32501 3885 32510 3905
rect 32527 3885 32533 3905
rect 32501 3875 32533 3885
rect 32550 3905 32576 3915
rect 32550 3885 32553 3905
rect 32573 3885 32576 3905
rect 32550 3875 32576 3885
rect 32595 3905 32625 3945
rect 32595 3885 32600 3905
rect 32620 3885 32625 3905
rect 32595 3875 32625 3885
rect 31210 3855 31230 3875
rect 31870 3855 31890 3875
rect 31940 3855 31960 3875
rect 32600 3855 32620 3875
rect 32660 3855 32680 3915
rect 31150 3835 31875 3855
rect 31955 3835 32680 3855
rect 31815 3820 31845 3835
rect 32965 3820 32995 3850
rect 29905 3740 30265 3760
rect 30345 3740 30705 3760
rect 29485 3680 29765 3700
rect 29485 3375 29505 3680
rect 29554 3655 29695 3660
rect 29554 3625 29560 3655
rect 29590 3625 29610 3655
rect 29640 3625 29659 3655
rect 29689 3625 29695 3655
rect 29554 3620 29695 3625
rect 29485 2995 29505 3280
rect 29745 3375 29765 3680
rect 29554 3050 29695 3055
rect 29554 3020 29560 3050
rect 29590 3020 29610 3050
rect 29640 3020 29659 3050
rect 29689 3020 29695 3050
rect 29554 3015 29695 3020
rect 29745 2995 29765 3280
rect 29485 2985 29585 2995
rect 29485 2975 29535 2985
rect 29525 2965 29535 2975
rect 29555 2975 29585 2985
rect 29665 2975 29765 2995
rect 29905 3410 29925 3740
rect 29955 3710 29995 3720
rect 29955 3690 29965 3710
rect 29985 3690 29995 3710
rect 29955 3680 29995 3690
rect 30065 3710 30105 3720
rect 30065 3690 30075 3710
rect 30095 3690 30105 3710
rect 30065 3680 30105 3690
rect 30175 3710 30215 3720
rect 30175 3690 30185 3710
rect 30205 3690 30215 3710
rect 30175 3680 30215 3690
rect 30285 3710 30325 3720
rect 30285 3690 30295 3710
rect 30315 3690 30325 3710
rect 30285 3680 30325 3690
rect 30395 3710 30435 3720
rect 30395 3690 30405 3710
rect 30425 3690 30435 3710
rect 30395 3680 30435 3690
rect 30505 3710 30545 3720
rect 30505 3690 30515 3710
rect 30535 3690 30545 3710
rect 30505 3680 30545 3690
rect 30615 3710 30655 3720
rect 30615 3690 30625 3710
rect 30645 3690 30655 3710
rect 30615 3680 30655 3690
rect 29965 3660 29985 3680
rect 30075 3660 30095 3680
rect 30185 3660 30205 3680
rect 30295 3660 30315 3680
rect 30405 3660 30425 3680
rect 30515 3660 30535 3680
rect 30625 3660 30645 3680
rect 29905 2990 29925 3315
rect 29960 3650 29990 3660
rect 29960 3630 29965 3650
rect 29985 3630 29990 3650
rect 29960 3600 29990 3630
rect 29960 3580 29965 3600
rect 29985 3580 29990 3600
rect 29960 3550 29990 3580
rect 29960 3530 29965 3550
rect 29985 3530 29990 3550
rect 29960 3500 29990 3530
rect 29960 3480 29965 3500
rect 29985 3480 29990 3500
rect 29960 3450 29990 3480
rect 29960 3430 29965 3450
rect 29985 3430 29990 3450
rect 29960 3400 29990 3430
rect 29960 3380 29965 3400
rect 29985 3380 29990 3400
rect 29960 3350 29990 3380
rect 29960 3330 29965 3350
rect 29985 3330 29990 3350
rect 29960 3300 29990 3330
rect 29960 3280 29965 3300
rect 29985 3280 29990 3300
rect 29960 3250 29990 3280
rect 29960 3230 29965 3250
rect 29985 3230 29990 3250
rect 29960 3200 29990 3230
rect 29960 3180 29965 3200
rect 29985 3180 29990 3200
rect 29960 3150 29990 3180
rect 29960 3130 29965 3150
rect 29985 3130 29990 3150
rect 29960 3100 29990 3130
rect 29960 3080 29965 3100
rect 29985 3080 29990 3100
rect 29960 3040 29990 3080
rect 30015 3650 30045 3660
rect 30015 3630 30020 3650
rect 30040 3630 30045 3650
rect 30015 3600 30045 3630
rect 30015 3580 30020 3600
rect 30040 3580 30045 3600
rect 30015 3550 30045 3580
rect 30015 3530 30020 3550
rect 30040 3530 30045 3550
rect 30015 3500 30045 3530
rect 30015 3480 30020 3500
rect 30040 3480 30045 3500
rect 30015 3450 30045 3480
rect 30015 3430 30020 3450
rect 30040 3430 30045 3450
rect 30015 3400 30045 3430
rect 30015 3380 30020 3400
rect 30040 3380 30045 3400
rect 30015 3350 30045 3380
rect 30015 3330 30020 3350
rect 30040 3330 30045 3350
rect 30015 3300 30045 3330
rect 30015 3280 30020 3300
rect 30040 3280 30045 3300
rect 30015 3250 30045 3280
rect 30015 3230 30020 3250
rect 30040 3230 30045 3250
rect 30015 3200 30045 3230
rect 30015 3180 30020 3200
rect 30040 3180 30045 3200
rect 30015 3150 30045 3180
rect 30015 3130 30020 3150
rect 30040 3130 30045 3150
rect 30015 3100 30045 3130
rect 30015 3080 30020 3100
rect 30040 3080 30045 3100
rect 30015 3070 30045 3080
rect 30070 3650 30100 3660
rect 30070 3630 30075 3650
rect 30095 3630 30100 3650
rect 30070 3600 30100 3630
rect 30070 3580 30075 3600
rect 30095 3580 30100 3600
rect 30070 3550 30100 3580
rect 30070 3530 30075 3550
rect 30095 3530 30100 3550
rect 30070 3500 30100 3530
rect 30070 3480 30075 3500
rect 30095 3480 30100 3500
rect 30070 3450 30100 3480
rect 30070 3430 30075 3450
rect 30095 3430 30100 3450
rect 30070 3400 30100 3430
rect 30070 3380 30075 3400
rect 30095 3380 30100 3400
rect 30070 3350 30100 3380
rect 30070 3330 30075 3350
rect 30095 3330 30100 3350
rect 30070 3300 30100 3330
rect 30070 3280 30075 3300
rect 30095 3280 30100 3300
rect 30070 3250 30100 3280
rect 30070 3230 30075 3250
rect 30095 3230 30100 3250
rect 30070 3200 30100 3230
rect 30070 3180 30075 3200
rect 30095 3180 30100 3200
rect 30070 3150 30100 3180
rect 30070 3130 30075 3150
rect 30095 3130 30100 3150
rect 30070 3100 30100 3130
rect 30070 3080 30075 3100
rect 30095 3080 30100 3100
rect 30070 3070 30100 3080
rect 30125 3650 30155 3660
rect 30125 3630 30130 3650
rect 30150 3630 30155 3650
rect 30125 3600 30155 3630
rect 30125 3580 30130 3600
rect 30150 3580 30155 3600
rect 30125 3550 30155 3580
rect 30125 3530 30130 3550
rect 30150 3530 30155 3550
rect 30125 3500 30155 3530
rect 30125 3480 30130 3500
rect 30150 3480 30155 3500
rect 30125 3450 30155 3480
rect 30125 3430 30130 3450
rect 30150 3430 30155 3450
rect 30125 3400 30155 3430
rect 30125 3380 30130 3400
rect 30150 3380 30155 3400
rect 30125 3350 30155 3380
rect 30125 3330 30130 3350
rect 30150 3330 30155 3350
rect 30125 3300 30155 3330
rect 30125 3280 30130 3300
rect 30150 3280 30155 3300
rect 30125 3250 30155 3280
rect 30125 3230 30130 3250
rect 30150 3230 30155 3250
rect 30125 3200 30155 3230
rect 30125 3180 30130 3200
rect 30150 3180 30155 3200
rect 30125 3150 30155 3180
rect 30125 3130 30130 3150
rect 30150 3130 30155 3150
rect 30125 3100 30155 3130
rect 30125 3080 30130 3100
rect 30150 3080 30155 3100
rect 30125 3070 30155 3080
rect 30180 3650 30210 3660
rect 30180 3630 30185 3650
rect 30205 3630 30210 3650
rect 30180 3600 30210 3630
rect 30180 3580 30185 3600
rect 30205 3580 30210 3600
rect 30180 3550 30210 3580
rect 30180 3530 30185 3550
rect 30205 3530 30210 3550
rect 30180 3500 30210 3530
rect 30180 3480 30185 3500
rect 30205 3480 30210 3500
rect 30180 3450 30210 3480
rect 30180 3430 30185 3450
rect 30205 3430 30210 3450
rect 30180 3400 30210 3430
rect 30180 3380 30185 3400
rect 30205 3380 30210 3400
rect 30180 3350 30210 3380
rect 30180 3330 30185 3350
rect 30205 3330 30210 3350
rect 30180 3300 30210 3330
rect 30180 3280 30185 3300
rect 30205 3280 30210 3300
rect 30180 3250 30210 3280
rect 30180 3230 30185 3250
rect 30205 3230 30210 3250
rect 30180 3200 30210 3230
rect 30180 3180 30185 3200
rect 30205 3180 30210 3200
rect 30180 3150 30210 3180
rect 30180 3130 30185 3150
rect 30205 3130 30210 3150
rect 30180 3100 30210 3130
rect 30180 3080 30185 3100
rect 30205 3080 30210 3100
rect 30180 3070 30210 3080
rect 30235 3650 30265 3660
rect 30235 3630 30240 3650
rect 30260 3630 30265 3650
rect 30235 3600 30265 3630
rect 30235 3580 30240 3600
rect 30260 3580 30265 3600
rect 30235 3550 30265 3580
rect 30235 3530 30240 3550
rect 30260 3530 30265 3550
rect 30235 3500 30265 3530
rect 30235 3480 30240 3500
rect 30260 3480 30265 3500
rect 30235 3450 30265 3480
rect 30235 3430 30240 3450
rect 30260 3430 30265 3450
rect 30235 3400 30265 3430
rect 30235 3380 30240 3400
rect 30260 3380 30265 3400
rect 30235 3350 30265 3380
rect 30235 3330 30240 3350
rect 30260 3330 30265 3350
rect 30235 3300 30265 3330
rect 30235 3280 30240 3300
rect 30260 3280 30265 3300
rect 30235 3250 30265 3280
rect 30235 3230 30240 3250
rect 30260 3230 30265 3250
rect 30235 3200 30265 3230
rect 30235 3180 30240 3200
rect 30260 3180 30265 3200
rect 30235 3150 30265 3180
rect 30235 3130 30240 3150
rect 30260 3130 30265 3150
rect 30235 3100 30265 3130
rect 30235 3080 30240 3100
rect 30260 3080 30265 3100
rect 30235 3070 30265 3080
rect 30290 3650 30320 3660
rect 30290 3630 30295 3650
rect 30315 3630 30320 3650
rect 30290 3600 30320 3630
rect 30290 3580 30295 3600
rect 30315 3580 30320 3600
rect 30290 3550 30320 3580
rect 30290 3530 30295 3550
rect 30315 3530 30320 3550
rect 30290 3500 30320 3530
rect 30290 3480 30295 3500
rect 30315 3480 30320 3500
rect 30290 3450 30320 3480
rect 30290 3430 30295 3450
rect 30315 3430 30320 3450
rect 30290 3400 30320 3430
rect 30290 3380 30295 3400
rect 30315 3380 30320 3400
rect 30290 3350 30320 3380
rect 30290 3330 30295 3350
rect 30315 3330 30320 3350
rect 30290 3300 30320 3330
rect 30290 3280 30295 3300
rect 30315 3280 30320 3300
rect 30290 3250 30320 3280
rect 30290 3230 30295 3250
rect 30315 3230 30320 3250
rect 30290 3200 30320 3230
rect 30290 3180 30295 3200
rect 30315 3180 30320 3200
rect 30290 3150 30320 3180
rect 30290 3130 30295 3150
rect 30315 3130 30320 3150
rect 30290 3100 30320 3130
rect 30290 3080 30295 3100
rect 30315 3080 30320 3100
rect 30290 3070 30320 3080
rect 30345 3650 30375 3660
rect 30345 3630 30350 3650
rect 30370 3630 30375 3650
rect 30345 3600 30375 3630
rect 30345 3580 30350 3600
rect 30370 3580 30375 3600
rect 30345 3550 30375 3580
rect 30345 3530 30350 3550
rect 30370 3530 30375 3550
rect 30345 3500 30375 3530
rect 30345 3480 30350 3500
rect 30370 3480 30375 3500
rect 30345 3450 30375 3480
rect 30345 3430 30350 3450
rect 30370 3430 30375 3450
rect 30345 3400 30375 3430
rect 30345 3380 30350 3400
rect 30370 3380 30375 3400
rect 30345 3350 30375 3380
rect 30345 3330 30350 3350
rect 30370 3330 30375 3350
rect 30345 3300 30375 3330
rect 30345 3280 30350 3300
rect 30370 3280 30375 3300
rect 30345 3250 30375 3280
rect 30345 3230 30350 3250
rect 30370 3230 30375 3250
rect 30345 3200 30375 3230
rect 30345 3180 30350 3200
rect 30370 3180 30375 3200
rect 30345 3150 30375 3180
rect 30345 3130 30350 3150
rect 30370 3130 30375 3150
rect 30345 3100 30375 3130
rect 30345 3080 30350 3100
rect 30370 3080 30375 3100
rect 30345 3070 30375 3080
rect 30400 3650 30430 3660
rect 30400 3630 30405 3650
rect 30425 3630 30430 3650
rect 30400 3600 30430 3630
rect 30400 3580 30405 3600
rect 30425 3580 30430 3600
rect 30400 3550 30430 3580
rect 30400 3530 30405 3550
rect 30425 3530 30430 3550
rect 30400 3500 30430 3530
rect 30400 3480 30405 3500
rect 30425 3480 30430 3500
rect 30400 3450 30430 3480
rect 30400 3430 30405 3450
rect 30425 3430 30430 3450
rect 30400 3400 30430 3430
rect 30400 3380 30405 3400
rect 30425 3380 30430 3400
rect 30400 3350 30430 3380
rect 30400 3330 30405 3350
rect 30425 3330 30430 3350
rect 30400 3300 30430 3330
rect 30400 3280 30405 3300
rect 30425 3280 30430 3300
rect 30400 3250 30430 3280
rect 30400 3230 30405 3250
rect 30425 3230 30430 3250
rect 30400 3200 30430 3230
rect 30400 3180 30405 3200
rect 30425 3180 30430 3200
rect 30400 3150 30430 3180
rect 30400 3130 30405 3150
rect 30425 3130 30430 3150
rect 30400 3100 30430 3130
rect 30400 3080 30405 3100
rect 30425 3080 30430 3100
rect 30400 3070 30430 3080
rect 30455 3650 30485 3660
rect 30455 3630 30460 3650
rect 30480 3630 30485 3650
rect 30455 3600 30485 3630
rect 30455 3580 30460 3600
rect 30480 3580 30485 3600
rect 30455 3550 30485 3580
rect 30455 3530 30460 3550
rect 30480 3530 30485 3550
rect 30455 3500 30485 3530
rect 30455 3480 30460 3500
rect 30480 3480 30485 3500
rect 30455 3450 30485 3480
rect 30455 3430 30460 3450
rect 30480 3430 30485 3450
rect 30455 3400 30485 3430
rect 30455 3380 30460 3400
rect 30480 3380 30485 3400
rect 30455 3350 30485 3380
rect 30455 3330 30460 3350
rect 30480 3330 30485 3350
rect 30455 3300 30485 3330
rect 30455 3280 30460 3300
rect 30480 3280 30485 3300
rect 30455 3250 30485 3280
rect 30455 3230 30460 3250
rect 30480 3230 30485 3250
rect 30455 3200 30485 3230
rect 30455 3180 30460 3200
rect 30480 3180 30485 3200
rect 30455 3150 30485 3180
rect 30455 3130 30460 3150
rect 30480 3130 30485 3150
rect 30455 3100 30485 3130
rect 30455 3080 30460 3100
rect 30480 3080 30485 3100
rect 30455 3070 30485 3080
rect 30510 3650 30540 3660
rect 30510 3630 30515 3650
rect 30535 3630 30540 3650
rect 30510 3600 30540 3630
rect 30510 3580 30515 3600
rect 30535 3580 30540 3600
rect 30510 3550 30540 3580
rect 30510 3530 30515 3550
rect 30535 3530 30540 3550
rect 30510 3500 30540 3530
rect 30510 3480 30515 3500
rect 30535 3480 30540 3500
rect 30510 3450 30540 3480
rect 30510 3430 30515 3450
rect 30535 3430 30540 3450
rect 30510 3400 30540 3430
rect 30510 3380 30515 3400
rect 30535 3380 30540 3400
rect 30510 3350 30540 3380
rect 30510 3330 30515 3350
rect 30535 3330 30540 3350
rect 30510 3300 30540 3330
rect 30510 3280 30515 3300
rect 30535 3280 30540 3300
rect 30510 3250 30540 3280
rect 30510 3230 30515 3250
rect 30535 3230 30540 3250
rect 30510 3200 30540 3230
rect 30510 3180 30515 3200
rect 30535 3180 30540 3200
rect 30510 3150 30540 3180
rect 30510 3130 30515 3150
rect 30535 3130 30540 3150
rect 30510 3100 30540 3130
rect 30510 3080 30515 3100
rect 30535 3080 30540 3100
rect 30510 3070 30540 3080
rect 30565 3650 30595 3660
rect 30565 3630 30570 3650
rect 30590 3630 30595 3650
rect 30565 3600 30595 3630
rect 30565 3580 30570 3600
rect 30590 3580 30595 3600
rect 30565 3550 30595 3580
rect 30565 3530 30570 3550
rect 30590 3530 30595 3550
rect 30565 3500 30595 3530
rect 30565 3480 30570 3500
rect 30590 3480 30595 3500
rect 30565 3450 30595 3480
rect 30565 3430 30570 3450
rect 30590 3430 30595 3450
rect 30565 3400 30595 3430
rect 30565 3380 30570 3400
rect 30590 3380 30595 3400
rect 30565 3350 30595 3380
rect 30565 3330 30570 3350
rect 30590 3330 30595 3350
rect 30565 3300 30595 3330
rect 30565 3280 30570 3300
rect 30590 3280 30595 3300
rect 30565 3250 30595 3280
rect 30565 3230 30570 3250
rect 30590 3230 30595 3250
rect 30565 3200 30595 3230
rect 30565 3180 30570 3200
rect 30590 3180 30595 3200
rect 30565 3150 30595 3180
rect 30565 3130 30570 3150
rect 30590 3130 30595 3150
rect 30565 3100 30595 3130
rect 30565 3080 30570 3100
rect 30590 3080 30595 3100
rect 30565 3070 30595 3080
rect 30620 3650 30650 3660
rect 30620 3630 30625 3650
rect 30645 3630 30650 3650
rect 30620 3600 30650 3630
rect 30620 3580 30625 3600
rect 30645 3580 30650 3600
rect 30620 3550 30650 3580
rect 30620 3530 30625 3550
rect 30645 3530 30650 3550
rect 30620 3500 30650 3530
rect 30620 3480 30625 3500
rect 30645 3480 30650 3500
rect 30620 3450 30650 3480
rect 30620 3430 30625 3450
rect 30645 3430 30650 3450
rect 30620 3400 30650 3430
rect 30620 3380 30625 3400
rect 30645 3380 30650 3400
rect 30620 3350 30650 3380
rect 30620 3330 30625 3350
rect 30645 3330 30650 3350
rect 30620 3300 30650 3330
rect 30620 3280 30625 3300
rect 30645 3280 30650 3300
rect 30620 3250 30650 3280
rect 30620 3230 30625 3250
rect 30645 3230 30650 3250
rect 30620 3200 30650 3230
rect 30620 3180 30625 3200
rect 30645 3180 30650 3200
rect 30620 3150 30650 3180
rect 30620 3130 30625 3150
rect 30645 3130 30650 3150
rect 30620 3100 30650 3130
rect 30620 3080 30625 3100
rect 30645 3080 30650 3100
rect 30020 3050 30040 3070
rect 30130 3050 30150 3070
rect 30240 3050 30260 3070
rect 30350 3050 30370 3070
rect 30460 3050 30480 3070
rect 30570 3050 30590 3070
rect 29960 3020 29965 3040
rect 29985 3020 29990 3040
rect 29960 3010 29990 3020
rect 30010 3040 30050 3050
rect 30010 3020 30020 3040
rect 30040 3020 30050 3040
rect 30010 3010 30050 3020
rect 30120 3040 30160 3050
rect 30120 3020 30130 3040
rect 30150 3020 30160 3040
rect 30120 3010 30160 3020
rect 30178 3040 30212 3050
rect 30178 3020 30186 3040
rect 30204 3020 30212 3040
rect 30178 3010 30212 3020
rect 30230 3040 30270 3050
rect 30230 3020 30240 3040
rect 30260 3020 30270 3040
rect 30230 3010 30270 3020
rect 30340 3040 30380 3050
rect 30340 3020 30350 3040
rect 30370 3020 30380 3040
rect 30340 3010 30380 3020
rect 30450 3040 30490 3050
rect 30450 3020 30460 3040
rect 30480 3020 30490 3040
rect 30450 3010 30490 3020
rect 30560 3040 30600 3050
rect 30560 3020 30570 3040
rect 30590 3020 30600 3040
rect 30560 3010 30600 3020
rect 30620 3040 30650 3080
rect 30620 3020 30625 3040
rect 30645 3020 30650 3040
rect 30620 3010 30650 3020
rect 30685 3410 30705 3740
rect 32085 3730 32115 3760
rect 32305 3730 32335 3760
rect 32545 3730 32575 3760
rect 32920 3730 32950 3760
rect 33095 3740 33455 3760
rect 33535 3740 33895 3760
rect 31885 3695 31915 3725
rect 33010 3685 33040 3715
rect 31880 3660 31920 3670
rect 31880 3650 31890 3660
rect 31910 3650 31920 3660
rect 29965 2990 29985 3010
rect 30625 2990 30645 3010
rect 30685 2990 30705 3315
rect 31170 3630 31860 3650
rect 31940 3630 32630 3650
rect 31170 3445 31190 3630
rect 31340 3600 31380 3610
rect 31340 3580 31350 3600
rect 31370 3580 31380 3600
rect 31340 3570 31380 3580
rect 31460 3600 31500 3610
rect 31460 3580 31470 3600
rect 31490 3580 31500 3600
rect 31460 3570 31500 3580
rect 31580 3600 31620 3610
rect 31580 3580 31590 3600
rect 31610 3580 31620 3600
rect 31580 3570 31620 3580
rect 31700 3600 31740 3610
rect 31700 3580 31710 3600
rect 31730 3580 31740 3600
rect 31700 3570 31740 3580
rect 31820 3600 31860 3610
rect 31820 3580 31830 3600
rect 31850 3580 31860 3600
rect 31820 3570 31860 3580
rect 31885 3600 31915 3605
rect 31885 3580 31890 3600
rect 31910 3580 31915 3600
rect 31885 3575 31915 3580
rect 31940 3600 31980 3610
rect 31940 3580 31950 3600
rect 31970 3580 31980 3600
rect 31940 3570 31980 3580
rect 32060 3600 32100 3610
rect 32060 3580 32070 3600
rect 32090 3580 32100 3600
rect 32060 3570 32100 3580
rect 32180 3600 32220 3610
rect 32180 3580 32190 3600
rect 32210 3580 32220 3600
rect 32180 3570 32220 3580
rect 32300 3600 32340 3610
rect 32300 3580 32310 3600
rect 32330 3580 32340 3600
rect 32300 3570 32340 3580
rect 32420 3600 32460 3610
rect 32420 3580 32430 3600
rect 32450 3580 32460 3600
rect 32420 3570 32460 3580
rect 31350 3550 31370 3570
rect 31470 3550 31490 3570
rect 31590 3550 31610 3570
rect 31710 3550 31730 3570
rect 31830 3550 31850 3570
rect 31950 3550 31970 3570
rect 32070 3550 32090 3570
rect 32190 3550 32210 3570
rect 32310 3550 32330 3570
rect 32430 3550 32450 3570
rect 31170 3130 31190 3365
rect 31225 3540 31255 3550
rect 31225 3520 31230 3540
rect 31250 3520 31255 3540
rect 31225 3490 31255 3520
rect 31225 3470 31230 3490
rect 31250 3470 31255 3490
rect 31225 3440 31255 3470
rect 31225 3420 31230 3440
rect 31250 3420 31255 3440
rect 31225 3390 31255 3420
rect 31225 3370 31230 3390
rect 31250 3370 31255 3390
rect 31225 3340 31255 3370
rect 31225 3320 31230 3340
rect 31250 3320 31255 3340
rect 31225 3290 31255 3320
rect 31225 3270 31230 3290
rect 31250 3270 31255 3290
rect 31225 3240 31255 3270
rect 31225 3220 31230 3240
rect 31250 3220 31255 3240
rect 31225 3180 31255 3220
rect 31285 3540 31315 3550
rect 31285 3520 31290 3540
rect 31310 3520 31315 3540
rect 31285 3490 31315 3520
rect 31285 3470 31290 3490
rect 31310 3470 31315 3490
rect 31285 3440 31315 3470
rect 31285 3420 31290 3440
rect 31310 3420 31315 3440
rect 31285 3390 31315 3420
rect 31285 3370 31290 3390
rect 31310 3370 31315 3390
rect 31285 3340 31315 3370
rect 31285 3320 31290 3340
rect 31310 3320 31315 3340
rect 31285 3290 31315 3320
rect 31285 3270 31290 3290
rect 31310 3270 31315 3290
rect 31285 3240 31315 3270
rect 31285 3220 31290 3240
rect 31310 3220 31315 3240
rect 31285 3210 31315 3220
rect 31345 3540 31375 3550
rect 31345 3520 31350 3540
rect 31370 3520 31375 3540
rect 31345 3490 31375 3520
rect 31345 3470 31350 3490
rect 31370 3470 31375 3490
rect 31345 3440 31375 3470
rect 31345 3420 31350 3440
rect 31370 3420 31375 3440
rect 31345 3390 31375 3420
rect 31345 3370 31350 3390
rect 31370 3370 31375 3390
rect 31345 3340 31375 3370
rect 31345 3320 31350 3340
rect 31370 3320 31375 3340
rect 31345 3290 31375 3320
rect 31345 3270 31350 3290
rect 31370 3270 31375 3290
rect 31345 3240 31375 3270
rect 31345 3220 31350 3240
rect 31370 3220 31375 3240
rect 31345 3210 31375 3220
rect 31405 3540 31435 3550
rect 31405 3520 31410 3540
rect 31430 3520 31435 3540
rect 31405 3490 31435 3520
rect 31405 3470 31410 3490
rect 31430 3470 31435 3490
rect 31405 3440 31435 3470
rect 31405 3420 31410 3440
rect 31430 3420 31435 3440
rect 31405 3390 31435 3420
rect 31405 3370 31410 3390
rect 31430 3370 31435 3390
rect 31405 3340 31435 3370
rect 31405 3320 31410 3340
rect 31430 3320 31435 3340
rect 31405 3290 31435 3320
rect 31405 3270 31410 3290
rect 31430 3270 31435 3290
rect 31405 3240 31435 3270
rect 31405 3220 31410 3240
rect 31430 3220 31435 3240
rect 31405 3210 31435 3220
rect 31465 3540 31495 3550
rect 31465 3520 31470 3540
rect 31490 3520 31495 3540
rect 31465 3490 31495 3520
rect 31465 3470 31470 3490
rect 31490 3470 31495 3490
rect 31465 3440 31495 3470
rect 31465 3420 31470 3440
rect 31490 3420 31495 3440
rect 31465 3390 31495 3420
rect 31465 3370 31470 3390
rect 31490 3370 31495 3390
rect 31465 3340 31495 3370
rect 31465 3320 31470 3340
rect 31490 3320 31495 3340
rect 31465 3290 31495 3320
rect 31465 3270 31470 3290
rect 31490 3270 31495 3290
rect 31465 3240 31495 3270
rect 31465 3220 31470 3240
rect 31490 3220 31495 3240
rect 31465 3210 31495 3220
rect 31525 3540 31555 3550
rect 31525 3520 31530 3540
rect 31550 3520 31555 3540
rect 31525 3490 31555 3520
rect 31525 3470 31530 3490
rect 31550 3470 31555 3490
rect 31525 3440 31555 3470
rect 31525 3420 31530 3440
rect 31550 3420 31555 3440
rect 31525 3390 31555 3420
rect 31525 3370 31530 3390
rect 31550 3370 31555 3390
rect 31525 3340 31555 3370
rect 31525 3320 31530 3340
rect 31550 3320 31555 3340
rect 31525 3290 31555 3320
rect 31525 3270 31530 3290
rect 31550 3270 31555 3290
rect 31525 3240 31555 3270
rect 31525 3220 31530 3240
rect 31550 3220 31555 3240
rect 31525 3210 31555 3220
rect 31585 3540 31615 3550
rect 31585 3520 31590 3540
rect 31610 3520 31615 3540
rect 31585 3490 31615 3520
rect 31585 3470 31590 3490
rect 31610 3470 31615 3490
rect 31585 3440 31615 3470
rect 31585 3420 31590 3440
rect 31610 3420 31615 3440
rect 31585 3390 31615 3420
rect 31585 3370 31590 3390
rect 31610 3370 31615 3390
rect 31585 3340 31615 3370
rect 31585 3320 31590 3340
rect 31610 3320 31615 3340
rect 31585 3290 31615 3320
rect 31585 3270 31590 3290
rect 31610 3270 31615 3290
rect 31585 3240 31615 3270
rect 31585 3220 31590 3240
rect 31610 3220 31615 3240
rect 31585 3210 31615 3220
rect 31645 3540 31675 3550
rect 31645 3520 31650 3540
rect 31670 3520 31675 3540
rect 31645 3490 31675 3520
rect 31645 3470 31650 3490
rect 31670 3470 31675 3490
rect 31645 3440 31675 3470
rect 31645 3420 31650 3440
rect 31670 3420 31675 3440
rect 31645 3390 31675 3420
rect 31645 3370 31650 3390
rect 31670 3370 31675 3390
rect 31645 3340 31675 3370
rect 31645 3320 31650 3340
rect 31670 3320 31675 3340
rect 31645 3290 31675 3320
rect 31645 3270 31650 3290
rect 31670 3270 31675 3290
rect 31645 3240 31675 3270
rect 31645 3220 31650 3240
rect 31670 3220 31675 3240
rect 31645 3210 31675 3220
rect 31705 3540 31735 3550
rect 31705 3520 31710 3540
rect 31730 3520 31735 3540
rect 31705 3490 31735 3520
rect 31705 3470 31710 3490
rect 31730 3470 31735 3490
rect 31705 3440 31735 3470
rect 31705 3420 31710 3440
rect 31730 3420 31735 3440
rect 31705 3390 31735 3420
rect 31705 3370 31710 3390
rect 31730 3370 31735 3390
rect 31705 3340 31735 3370
rect 31705 3320 31710 3340
rect 31730 3320 31735 3340
rect 31705 3290 31735 3320
rect 31705 3270 31710 3290
rect 31730 3270 31735 3290
rect 31705 3240 31735 3270
rect 31705 3220 31710 3240
rect 31730 3220 31735 3240
rect 31705 3210 31735 3220
rect 31765 3540 31795 3550
rect 31765 3520 31770 3540
rect 31790 3520 31795 3540
rect 31765 3490 31795 3520
rect 31765 3470 31770 3490
rect 31790 3470 31795 3490
rect 31765 3440 31795 3470
rect 31765 3420 31770 3440
rect 31790 3420 31795 3440
rect 31765 3390 31795 3420
rect 31765 3370 31770 3390
rect 31790 3370 31795 3390
rect 31765 3340 31795 3370
rect 31765 3320 31770 3340
rect 31790 3320 31795 3340
rect 31765 3290 31795 3320
rect 31765 3270 31770 3290
rect 31790 3270 31795 3290
rect 31765 3240 31795 3270
rect 31765 3220 31770 3240
rect 31790 3220 31795 3240
rect 31765 3210 31795 3220
rect 31825 3540 31855 3550
rect 31825 3520 31830 3540
rect 31850 3520 31855 3540
rect 31825 3490 31855 3520
rect 31825 3470 31830 3490
rect 31850 3470 31855 3490
rect 31825 3440 31855 3470
rect 31825 3420 31830 3440
rect 31850 3420 31855 3440
rect 31825 3390 31855 3420
rect 31825 3370 31830 3390
rect 31850 3370 31855 3390
rect 31825 3340 31855 3370
rect 31825 3320 31830 3340
rect 31850 3320 31855 3340
rect 31825 3290 31855 3320
rect 31825 3270 31830 3290
rect 31850 3270 31855 3290
rect 31825 3240 31855 3270
rect 31825 3220 31830 3240
rect 31850 3220 31855 3240
rect 31825 3210 31855 3220
rect 31885 3540 31915 3550
rect 31885 3520 31890 3540
rect 31910 3520 31915 3540
rect 31885 3490 31915 3520
rect 31885 3470 31890 3490
rect 31910 3470 31915 3490
rect 31885 3440 31915 3470
rect 31885 3420 31890 3440
rect 31910 3420 31915 3440
rect 31885 3390 31915 3420
rect 31885 3370 31890 3390
rect 31910 3370 31915 3390
rect 31885 3340 31915 3370
rect 31885 3320 31890 3340
rect 31910 3320 31915 3340
rect 31885 3290 31915 3320
rect 31885 3270 31890 3290
rect 31910 3270 31915 3290
rect 31885 3240 31915 3270
rect 31885 3220 31890 3240
rect 31910 3220 31915 3240
rect 31885 3210 31915 3220
rect 31945 3540 31975 3550
rect 31945 3520 31950 3540
rect 31970 3520 31975 3540
rect 31945 3490 31975 3520
rect 31945 3470 31950 3490
rect 31970 3470 31975 3490
rect 31945 3440 31975 3470
rect 31945 3420 31950 3440
rect 31970 3420 31975 3440
rect 31945 3390 31975 3420
rect 31945 3370 31950 3390
rect 31970 3370 31975 3390
rect 31945 3340 31975 3370
rect 31945 3320 31950 3340
rect 31970 3320 31975 3340
rect 31945 3290 31975 3320
rect 31945 3270 31950 3290
rect 31970 3270 31975 3290
rect 31945 3240 31975 3270
rect 31945 3220 31950 3240
rect 31970 3220 31975 3240
rect 31945 3210 31975 3220
rect 32005 3540 32035 3550
rect 32005 3520 32010 3540
rect 32030 3520 32035 3540
rect 32005 3490 32035 3520
rect 32005 3470 32010 3490
rect 32030 3470 32035 3490
rect 32005 3440 32035 3470
rect 32005 3420 32010 3440
rect 32030 3420 32035 3440
rect 32005 3390 32035 3420
rect 32005 3370 32010 3390
rect 32030 3370 32035 3390
rect 32005 3340 32035 3370
rect 32005 3320 32010 3340
rect 32030 3320 32035 3340
rect 32005 3290 32035 3320
rect 32005 3270 32010 3290
rect 32030 3270 32035 3290
rect 32005 3240 32035 3270
rect 32005 3220 32010 3240
rect 32030 3220 32035 3240
rect 32005 3210 32035 3220
rect 32065 3540 32095 3550
rect 32065 3520 32070 3540
rect 32090 3520 32095 3540
rect 32065 3490 32095 3520
rect 32065 3470 32070 3490
rect 32090 3470 32095 3490
rect 32065 3440 32095 3470
rect 32065 3420 32070 3440
rect 32090 3420 32095 3440
rect 32065 3390 32095 3420
rect 32065 3370 32070 3390
rect 32090 3370 32095 3390
rect 32065 3340 32095 3370
rect 32065 3320 32070 3340
rect 32090 3320 32095 3340
rect 32065 3290 32095 3320
rect 32065 3270 32070 3290
rect 32090 3270 32095 3290
rect 32065 3240 32095 3270
rect 32065 3220 32070 3240
rect 32090 3220 32095 3240
rect 32065 3210 32095 3220
rect 32125 3540 32155 3550
rect 32125 3520 32130 3540
rect 32150 3520 32155 3540
rect 32125 3490 32155 3520
rect 32125 3470 32130 3490
rect 32150 3470 32155 3490
rect 32125 3440 32155 3470
rect 32125 3420 32130 3440
rect 32150 3420 32155 3440
rect 32125 3390 32155 3420
rect 32125 3370 32130 3390
rect 32150 3370 32155 3390
rect 32125 3340 32155 3370
rect 32125 3320 32130 3340
rect 32150 3320 32155 3340
rect 32125 3290 32155 3320
rect 32125 3270 32130 3290
rect 32150 3270 32155 3290
rect 32125 3240 32155 3270
rect 32125 3220 32130 3240
rect 32150 3220 32155 3240
rect 32125 3210 32155 3220
rect 32185 3540 32215 3550
rect 32185 3520 32190 3540
rect 32210 3520 32215 3540
rect 32185 3490 32215 3520
rect 32185 3470 32190 3490
rect 32210 3470 32215 3490
rect 32185 3440 32215 3470
rect 32185 3420 32190 3440
rect 32210 3420 32215 3440
rect 32185 3390 32215 3420
rect 32185 3370 32190 3390
rect 32210 3370 32215 3390
rect 32185 3340 32215 3370
rect 32185 3320 32190 3340
rect 32210 3320 32215 3340
rect 32185 3290 32215 3320
rect 32185 3270 32190 3290
rect 32210 3270 32215 3290
rect 32185 3240 32215 3270
rect 32185 3220 32190 3240
rect 32210 3220 32215 3240
rect 32185 3210 32215 3220
rect 32245 3540 32275 3550
rect 32245 3520 32250 3540
rect 32270 3520 32275 3540
rect 32245 3490 32275 3520
rect 32245 3470 32250 3490
rect 32270 3470 32275 3490
rect 32245 3440 32275 3470
rect 32245 3420 32250 3440
rect 32270 3420 32275 3440
rect 32245 3390 32275 3420
rect 32245 3370 32250 3390
rect 32270 3370 32275 3390
rect 32245 3340 32275 3370
rect 32245 3320 32250 3340
rect 32270 3320 32275 3340
rect 32245 3290 32275 3320
rect 32245 3270 32250 3290
rect 32270 3270 32275 3290
rect 32245 3240 32275 3270
rect 32245 3220 32250 3240
rect 32270 3220 32275 3240
rect 32245 3210 32275 3220
rect 32305 3540 32335 3550
rect 32305 3520 32310 3540
rect 32330 3520 32335 3540
rect 32305 3490 32335 3520
rect 32305 3470 32310 3490
rect 32330 3470 32335 3490
rect 32305 3440 32335 3470
rect 32305 3420 32310 3440
rect 32330 3420 32335 3440
rect 32305 3390 32335 3420
rect 32305 3370 32310 3390
rect 32330 3370 32335 3390
rect 32305 3340 32335 3370
rect 32305 3320 32310 3340
rect 32330 3320 32335 3340
rect 32305 3290 32335 3320
rect 32305 3270 32310 3290
rect 32330 3270 32335 3290
rect 32305 3240 32335 3270
rect 32305 3220 32310 3240
rect 32330 3220 32335 3240
rect 32305 3210 32335 3220
rect 32365 3540 32395 3550
rect 32365 3520 32370 3540
rect 32390 3520 32395 3540
rect 32365 3490 32395 3520
rect 32365 3470 32370 3490
rect 32390 3470 32395 3490
rect 32365 3440 32395 3470
rect 32365 3420 32370 3440
rect 32390 3420 32395 3440
rect 32365 3390 32395 3420
rect 32365 3370 32370 3390
rect 32390 3370 32395 3390
rect 32365 3340 32395 3370
rect 32365 3320 32370 3340
rect 32390 3320 32395 3340
rect 32365 3290 32395 3320
rect 32365 3270 32370 3290
rect 32390 3270 32395 3290
rect 32365 3240 32395 3270
rect 32365 3220 32370 3240
rect 32390 3220 32395 3240
rect 32365 3210 32395 3220
rect 32425 3540 32455 3550
rect 32425 3520 32430 3540
rect 32450 3520 32455 3540
rect 32425 3490 32455 3520
rect 32425 3470 32430 3490
rect 32450 3470 32455 3490
rect 32425 3440 32455 3470
rect 32425 3420 32430 3440
rect 32450 3420 32455 3440
rect 32425 3390 32455 3420
rect 32425 3370 32430 3390
rect 32450 3370 32455 3390
rect 32425 3340 32455 3370
rect 32425 3320 32430 3340
rect 32450 3320 32455 3340
rect 32425 3290 32455 3320
rect 32425 3270 32430 3290
rect 32450 3270 32455 3290
rect 32425 3240 32455 3270
rect 32425 3220 32430 3240
rect 32450 3220 32455 3240
rect 32425 3210 32455 3220
rect 32485 3540 32515 3550
rect 32485 3520 32490 3540
rect 32510 3520 32515 3540
rect 32485 3490 32515 3520
rect 32485 3470 32490 3490
rect 32510 3470 32515 3490
rect 32485 3440 32515 3470
rect 32485 3420 32490 3440
rect 32510 3420 32515 3440
rect 32485 3390 32515 3420
rect 32485 3370 32490 3390
rect 32510 3370 32515 3390
rect 32485 3340 32515 3370
rect 32485 3320 32490 3340
rect 32510 3320 32515 3340
rect 32485 3290 32515 3320
rect 32485 3270 32490 3290
rect 32510 3270 32515 3290
rect 32485 3240 32515 3270
rect 32485 3220 32490 3240
rect 32510 3220 32515 3240
rect 32485 3210 32515 3220
rect 32545 3540 32575 3550
rect 32545 3520 32550 3540
rect 32570 3520 32575 3540
rect 32545 3490 32575 3520
rect 32545 3470 32550 3490
rect 32570 3470 32575 3490
rect 32545 3440 32575 3470
rect 32545 3420 32550 3440
rect 32570 3420 32575 3440
rect 32545 3390 32575 3420
rect 32545 3370 32550 3390
rect 32570 3370 32575 3390
rect 32545 3340 32575 3370
rect 32545 3320 32550 3340
rect 32570 3320 32575 3340
rect 32545 3290 32575 3320
rect 32545 3270 32550 3290
rect 32570 3270 32575 3290
rect 32545 3240 32575 3270
rect 32545 3220 32550 3240
rect 32570 3220 32575 3240
rect 31290 3190 31310 3210
rect 31410 3190 31430 3210
rect 31530 3190 31550 3210
rect 31650 3190 31670 3210
rect 31770 3190 31790 3210
rect 31890 3190 31910 3210
rect 32010 3190 32030 3210
rect 32130 3190 32150 3210
rect 32250 3190 32270 3210
rect 32370 3190 32390 3210
rect 32490 3190 32510 3210
rect 31225 3160 31230 3180
rect 31250 3160 31255 3180
rect 31225 3150 31255 3160
rect 31280 3180 31320 3190
rect 31280 3160 31290 3180
rect 31310 3160 31320 3180
rect 31280 3150 31320 3160
rect 31400 3180 31440 3190
rect 31400 3160 31410 3180
rect 31430 3160 31440 3180
rect 31400 3150 31440 3160
rect 31520 3180 31560 3190
rect 31520 3160 31530 3180
rect 31550 3160 31560 3180
rect 31520 3150 31560 3160
rect 31640 3180 31680 3190
rect 31640 3160 31650 3180
rect 31670 3160 31680 3180
rect 31640 3150 31680 3160
rect 31760 3180 31800 3190
rect 31760 3160 31770 3180
rect 31790 3160 31800 3180
rect 31760 3150 31800 3160
rect 31823 3180 31857 3190
rect 31823 3160 31831 3180
rect 31849 3160 31857 3180
rect 31823 3150 31857 3160
rect 31880 3180 31920 3190
rect 31880 3160 31890 3180
rect 31910 3160 31920 3180
rect 31880 3150 31920 3160
rect 32000 3180 32040 3190
rect 32000 3160 32010 3180
rect 32030 3160 32040 3180
rect 32000 3150 32040 3160
rect 32120 3180 32160 3190
rect 32120 3160 32130 3180
rect 32150 3160 32160 3180
rect 32120 3150 32160 3160
rect 32240 3180 32280 3190
rect 32240 3160 32250 3180
rect 32270 3160 32280 3180
rect 32240 3150 32280 3160
rect 32360 3180 32400 3190
rect 32360 3160 32370 3180
rect 32390 3160 32400 3180
rect 32360 3150 32400 3160
rect 32480 3180 32520 3190
rect 32480 3160 32490 3180
rect 32510 3160 32520 3180
rect 32480 3150 32520 3160
rect 32545 3180 32575 3220
rect 32545 3160 32550 3180
rect 32570 3160 32575 3180
rect 32545 3150 32575 3160
rect 32610 3445 32630 3630
rect 31230 3130 31250 3150
rect 32550 3130 32570 3150
rect 32610 3130 32630 3365
rect 31170 3110 31860 3130
rect 31940 3110 32630 3130
rect 33095 3410 33115 3740
rect 33145 3710 33185 3720
rect 33145 3690 33155 3710
rect 33175 3690 33185 3710
rect 33145 3680 33185 3690
rect 33255 3710 33295 3720
rect 33255 3690 33265 3710
rect 33285 3690 33295 3710
rect 33255 3680 33295 3690
rect 33365 3710 33405 3720
rect 33365 3690 33375 3710
rect 33395 3690 33405 3710
rect 33365 3680 33405 3690
rect 33475 3710 33515 3720
rect 33475 3690 33485 3710
rect 33505 3690 33515 3710
rect 33475 3680 33515 3690
rect 33585 3710 33625 3720
rect 33585 3690 33595 3710
rect 33615 3690 33625 3710
rect 33585 3680 33625 3690
rect 33695 3710 33735 3720
rect 33695 3690 33705 3710
rect 33725 3690 33735 3710
rect 33695 3680 33735 3690
rect 33805 3710 33845 3720
rect 33805 3690 33815 3710
rect 33835 3690 33845 3710
rect 33805 3680 33845 3690
rect 33155 3660 33175 3680
rect 33265 3660 33285 3680
rect 33375 3660 33395 3680
rect 33485 3660 33505 3680
rect 33595 3660 33615 3680
rect 33705 3660 33725 3680
rect 33815 3660 33835 3680
rect 29555 2965 29565 2975
rect 29905 2970 30265 2990
rect 30345 2970 30705 2990
rect 33095 2990 33115 3315
rect 33150 3650 33180 3660
rect 33150 3630 33155 3650
rect 33175 3630 33180 3650
rect 33150 3600 33180 3630
rect 33150 3580 33155 3600
rect 33175 3580 33180 3600
rect 33150 3550 33180 3580
rect 33150 3530 33155 3550
rect 33175 3530 33180 3550
rect 33150 3500 33180 3530
rect 33150 3480 33155 3500
rect 33175 3480 33180 3500
rect 33150 3450 33180 3480
rect 33150 3430 33155 3450
rect 33175 3430 33180 3450
rect 33150 3400 33180 3430
rect 33150 3380 33155 3400
rect 33175 3380 33180 3400
rect 33150 3350 33180 3380
rect 33150 3330 33155 3350
rect 33175 3330 33180 3350
rect 33150 3300 33180 3330
rect 33150 3280 33155 3300
rect 33175 3280 33180 3300
rect 33150 3250 33180 3280
rect 33150 3230 33155 3250
rect 33175 3230 33180 3250
rect 33150 3200 33180 3230
rect 33150 3180 33155 3200
rect 33175 3180 33180 3200
rect 33150 3150 33180 3180
rect 33150 3130 33155 3150
rect 33175 3130 33180 3150
rect 33150 3100 33180 3130
rect 33150 3080 33155 3100
rect 33175 3080 33180 3100
rect 33150 3040 33180 3080
rect 33205 3650 33235 3660
rect 33205 3630 33210 3650
rect 33230 3630 33235 3650
rect 33205 3600 33235 3630
rect 33205 3580 33210 3600
rect 33230 3580 33235 3600
rect 33205 3550 33235 3580
rect 33205 3530 33210 3550
rect 33230 3530 33235 3550
rect 33205 3500 33235 3530
rect 33205 3480 33210 3500
rect 33230 3480 33235 3500
rect 33205 3450 33235 3480
rect 33205 3430 33210 3450
rect 33230 3430 33235 3450
rect 33205 3400 33235 3430
rect 33205 3380 33210 3400
rect 33230 3380 33235 3400
rect 33205 3350 33235 3380
rect 33205 3330 33210 3350
rect 33230 3330 33235 3350
rect 33205 3300 33235 3330
rect 33205 3280 33210 3300
rect 33230 3280 33235 3300
rect 33205 3250 33235 3280
rect 33205 3230 33210 3250
rect 33230 3230 33235 3250
rect 33205 3200 33235 3230
rect 33205 3180 33210 3200
rect 33230 3180 33235 3200
rect 33205 3150 33235 3180
rect 33205 3130 33210 3150
rect 33230 3130 33235 3150
rect 33205 3100 33235 3130
rect 33205 3080 33210 3100
rect 33230 3080 33235 3100
rect 33205 3070 33235 3080
rect 33260 3650 33290 3660
rect 33260 3630 33265 3650
rect 33285 3630 33290 3650
rect 33260 3600 33290 3630
rect 33260 3580 33265 3600
rect 33285 3580 33290 3600
rect 33260 3550 33290 3580
rect 33260 3530 33265 3550
rect 33285 3530 33290 3550
rect 33260 3500 33290 3530
rect 33260 3480 33265 3500
rect 33285 3480 33290 3500
rect 33260 3450 33290 3480
rect 33260 3430 33265 3450
rect 33285 3430 33290 3450
rect 33260 3400 33290 3430
rect 33260 3380 33265 3400
rect 33285 3380 33290 3400
rect 33260 3350 33290 3380
rect 33260 3330 33265 3350
rect 33285 3330 33290 3350
rect 33260 3300 33290 3330
rect 33260 3280 33265 3300
rect 33285 3280 33290 3300
rect 33260 3250 33290 3280
rect 33260 3230 33265 3250
rect 33285 3230 33290 3250
rect 33260 3200 33290 3230
rect 33260 3180 33265 3200
rect 33285 3180 33290 3200
rect 33260 3150 33290 3180
rect 33260 3130 33265 3150
rect 33285 3130 33290 3150
rect 33260 3100 33290 3130
rect 33260 3080 33265 3100
rect 33285 3080 33290 3100
rect 33260 3070 33290 3080
rect 33315 3650 33345 3660
rect 33315 3630 33320 3650
rect 33340 3630 33345 3650
rect 33315 3600 33345 3630
rect 33315 3580 33320 3600
rect 33340 3580 33345 3600
rect 33315 3550 33345 3580
rect 33315 3530 33320 3550
rect 33340 3530 33345 3550
rect 33315 3500 33345 3530
rect 33315 3480 33320 3500
rect 33340 3480 33345 3500
rect 33315 3450 33345 3480
rect 33315 3430 33320 3450
rect 33340 3430 33345 3450
rect 33315 3400 33345 3430
rect 33315 3380 33320 3400
rect 33340 3380 33345 3400
rect 33315 3350 33345 3380
rect 33315 3330 33320 3350
rect 33340 3330 33345 3350
rect 33315 3300 33345 3330
rect 33315 3280 33320 3300
rect 33340 3280 33345 3300
rect 33315 3250 33345 3280
rect 33315 3230 33320 3250
rect 33340 3230 33345 3250
rect 33315 3200 33345 3230
rect 33315 3180 33320 3200
rect 33340 3180 33345 3200
rect 33315 3150 33345 3180
rect 33315 3130 33320 3150
rect 33340 3130 33345 3150
rect 33315 3100 33345 3130
rect 33315 3080 33320 3100
rect 33340 3080 33345 3100
rect 33315 3070 33345 3080
rect 33370 3650 33400 3660
rect 33370 3630 33375 3650
rect 33395 3630 33400 3650
rect 33370 3600 33400 3630
rect 33370 3580 33375 3600
rect 33395 3580 33400 3600
rect 33370 3550 33400 3580
rect 33370 3530 33375 3550
rect 33395 3530 33400 3550
rect 33370 3500 33400 3530
rect 33370 3480 33375 3500
rect 33395 3480 33400 3500
rect 33370 3450 33400 3480
rect 33370 3430 33375 3450
rect 33395 3430 33400 3450
rect 33370 3400 33400 3430
rect 33370 3380 33375 3400
rect 33395 3380 33400 3400
rect 33370 3350 33400 3380
rect 33370 3330 33375 3350
rect 33395 3330 33400 3350
rect 33370 3300 33400 3330
rect 33370 3280 33375 3300
rect 33395 3280 33400 3300
rect 33370 3250 33400 3280
rect 33370 3230 33375 3250
rect 33395 3230 33400 3250
rect 33370 3200 33400 3230
rect 33370 3180 33375 3200
rect 33395 3180 33400 3200
rect 33370 3150 33400 3180
rect 33370 3130 33375 3150
rect 33395 3130 33400 3150
rect 33370 3100 33400 3130
rect 33370 3080 33375 3100
rect 33395 3080 33400 3100
rect 33370 3070 33400 3080
rect 33425 3650 33455 3660
rect 33425 3630 33430 3650
rect 33450 3630 33455 3650
rect 33425 3600 33455 3630
rect 33425 3580 33430 3600
rect 33450 3580 33455 3600
rect 33425 3550 33455 3580
rect 33425 3530 33430 3550
rect 33450 3530 33455 3550
rect 33425 3500 33455 3530
rect 33425 3480 33430 3500
rect 33450 3480 33455 3500
rect 33425 3450 33455 3480
rect 33425 3430 33430 3450
rect 33450 3430 33455 3450
rect 33425 3400 33455 3430
rect 33425 3380 33430 3400
rect 33450 3380 33455 3400
rect 33425 3350 33455 3380
rect 33425 3330 33430 3350
rect 33450 3330 33455 3350
rect 33425 3300 33455 3330
rect 33425 3280 33430 3300
rect 33450 3280 33455 3300
rect 33425 3250 33455 3280
rect 33425 3230 33430 3250
rect 33450 3230 33455 3250
rect 33425 3200 33455 3230
rect 33425 3180 33430 3200
rect 33450 3180 33455 3200
rect 33425 3150 33455 3180
rect 33425 3130 33430 3150
rect 33450 3130 33455 3150
rect 33425 3100 33455 3130
rect 33425 3080 33430 3100
rect 33450 3080 33455 3100
rect 33425 3070 33455 3080
rect 33480 3650 33510 3660
rect 33480 3630 33485 3650
rect 33505 3630 33510 3650
rect 33480 3600 33510 3630
rect 33480 3580 33485 3600
rect 33505 3580 33510 3600
rect 33480 3550 33510 3580
rect 33480 3530 33485 3550
rect 33505 3530 33510 3550
rect 33480 3500 33510 3530
rect 33480 3480 33485 3500
rect 33505 3480 33510 3500
rect 33480 3450 33510 3480
rect 33480 3430 33485 3450
rect 33505 3430 33510 3450
rect 33480 3400 33510 3430
rect 33480 3380 33485 3400
rect 33505 3380 33510 3400
rect 33480 3350 33510 3380
rect 33480 3330 33485 3350
rect 33505 3330 33510 3350
rect 33480 3300 33510 3330
rect 33480 3280 33485 3300
rect 33505 3280 33510 3300
rect 33480 3250 33510 3280
rect 33480 3230 33485 3250
rect 33505 3230 33510 3250
rect 33480 3200 33510 3230
rect 33480 3180 33485 3200
rect 33505 3180 33510 3200
rect 33480 3150 33510 3180
rect 33480 3130 33485 3150
rect 33505 3130 33510 3150
rect 33480 3100 33510 3130
rect 33480 3080 33485 3100
rect 33505 3080 33510 3100
rect 33480 3070 33510 3080
rect 33535 3650 33565 3660
rect 33535 3630 33540 3650
rect 33560 3630 33565 3650
rect 33535 3600 33565 3630
rect 33535 3580 33540 3600
rect 33560 3580 33565 3600
rect 33535 3550 33565 3580
rect 33535 3530 33540 3550
rect 33560 3530 33565 3550
rect 33535 3500 33565 3530
rect 33535 3480 33540 3500
rect 33560 3480 33565 3500
rect 33535 3450 33565 3480
rect 33535 3430 33540 3450
rect 33560 3430 33565 3450
rect 33535 3400 33565 3430
rect 33535 3380 33540 3400
rect 33560 3380 33565 3400
rect 33535 3350 33565 3380
rect 33535 3330 33540 3350
rect 33560 3330 33565 3350
rect 33535 3300 33565 3330
rect 33535 3280 33540 3300
rect 33560 3280 33565 3300
rect 33535 3250 33565 3280
rect 33535 3230 33540 3250
rect 33560 3230 33565 3250
rect 33535 3200 33565 3230
rect 33535 3180 33540 3200
rect 33560 3180 33565 3200
rect 33535 3150 33565 3180
rect 33535 3130 33540 3150
rect 33560 3130 33565 3150
rect 33535 3100 33565 3130
rect 33535 3080 33540 3100
rect 33560 3080 33565 3100
rect 33535 3070 33565 3080
rect 33590 3650 33620 3660
rect 33590 3630 33595 3650
rect 33615 3630 33620 3650
rect 33590 3600 33620 3630
rect 33590 3580 33595 3600
rect 33615 3580 33620 3600
rect 33590 3550 33620 3580
rect 33590 3530 33595 3550
rect 33615 3530 33620 3550
rect 33590 3500 33620 3530
rect 33590 3480 33595 3500
rect 33615 3480 33620 3500
rect 33590 3450 33620 3480
rect 33590 3430 33595 3450
rect 33615 3430 33620 3450
rect 33590 3400 33620 3430
rect 33590 3380 33595 3400
rect 33615 3380 33620 3400
rect 33590 3350 33620 3380
rect 33590 3330 33595 3350
rect 33615 3330 33620 3350
rect 33590 3300 33620 3330
rect 33590 3280 33595 3300
rect 33615 3280 33620 3300
rect 33590 3250 33620 3280
rect 33590 3230 33595 3250
rect 33615 3230 33620 3250
rect 33590 3200 33620 3230
rect 33590 3180 33595 3200
rect 33615 3180 33620 3200
rect 33590 3150 33620 3180
rect 33590 3130 33595 3150
rect 33615 3130 33620 3150
rect 33590 3100 33620 3130
rect 33590 3080 33595 3100
rect 33615 3080 33620 3100
rect 33590 3070 33620 3080
rect 33645 3650 33675 3660
rect 33645 3630 33650 3650
rect 33670 3630 33675 3650
rect 33645 3600 33675 3630
rect 33645 3580 33650 3600
rect 33670 3580 33675 3600
rect 33645 3550 33675 3580
rect 33645 3530 33650 3550
rect 33670 3530 33675 3550
rect 33645 3500 33675 3530
rect 33645 3480 33650 3500
rect 33670 3480 33675 3500
rect 33645 3450 33675 3480
rect 33645 3430 33650 3450
rect 33670 3430 33675 3450
rect 33645 3400 33675 3430
rect 33645 3380 33650 3400
rect 33670 3380 33675 3400
rect 33645 3350 33675 3380
rect 33645 3330 33650 3350
rect 33670 3330 33675 3350
rect 33645 3300 33675 3330
rect 33645 3280 33650 3300
rect 33670 3280 33675 3300
rect 33645 3250 33675 3280
rect 33645 3230 33650 3250
rect 33670 3230 33675 3250
rect 33645 3200 33675 3230
rect 33645 3180 33650 3200
rect 33670 3180 33675 3200
rect 33645 3150 33675 3180
rect 33645 3130 33650 3150
rect 33670 3130 33675 3150
rect 33645 3100 33675 3130
rect 33645 3080 33650 3100
rect 33670 3080 33675 3100
rect 33645 3070 33675 3080
rect 33700 3650 33730 3660
rect 33700 3630 33705 3650
rect 33725 3630 33730 3650
rect 33700 3600 33730 3630
rect 33700 3580 33705 3600
rect 33725 3580 33730 3600
rect 33700 3550 33730 3580
rect 33700 3530 33705 3550
rect 33725 3530 33730 3550
rect 33700 3500 33730 3530
rect 33700 3480 33705 3500
rect 33725 3480 33730 3500
rect 33700 3450 33730 3480
rect 33700 3430 33705 3450
rect 33725 3430 33730 3450
rect 33700 3400 33730 3430
rect 33700 3380 33705 3400
rect 33725 3380 33730 3400
rect 33700 3350 33730 3380
rect 33700 3330 33705 3350
rect 33725 3330 33730 3350
rect 33700 3300 33730 3330
rect 33700 3280 33705 3300
rect 33725 3280 33730 3300
rect 33700 3250 33730 3280
rect 33700 3230 33705 3250
rect 33725 3230 33730 3250
rect 33700 3200 33730 3230
rect 33700 3180 33705 3200
rect 33725 3180 33730 3200
rect 33700 3150 33730 3180
rect 33700 3130 33705 3150
rect 33725 3130 33730 3150
rect 33700 3100 33730 3130
rect 33700 3080 33705 3100
rect 33725 3080 33730 3100
rect 33700 3070 33730 3080
rect 33755 3650 33785 3660
rect 33755 3630 33760 3650
rect 33780 3630 33785 3650
rect 33755 3600 33785 3630
rect 33755 3580 33760 3600
rect 33780 3580 33785 3600
rect 33755 3550 33785 3580
rect 33755 3530 33760 3550
rect 33780 3530 33785 3550
rect 33755 3500 33785 3530
rect 33755 3480 33760 3500
rect 33780 3480 33785 3500
rect 33755 3450 33785 3480
rect 33755 3430 33760 3450
rect 33780 3430 33785 3450
rect 33755 3400 33785 3430
rect 33755 3380 33760 3400
rect 33780 3380 33785 3400
rect 33755 3350 33785 3380
rect 33755 3330 33760 3350
rect 33780 3330 33785 3350
rect 33755 3300 33785 3330
rect 33755 3280 33760 3300
rect 33780 3280 33785 3300
rect 33755 3250 33785 3280
rect 33755 3230 33760 3250
rect 33780 3230 33785 3250
rect 33755 3200 33785 3230
rect 33755 3180 33760 3200
rect 33780 3180 33785 3200
rect 33755 3150 33785 3180
rect 33755 3130 33760 3150
rect 33780 3130 33785 3150
rect 33755 3100 33785 3130
rect 33755 3080 33760 3100
rect 33780 3080 33785 3100
rect 33755 3070 33785 3080
rect 33810 3650 33840 3660
rect 33810 3630 33815 3650
rect 33835 3630 33840 3650
rect 33810 3600 33840 3630
rect 33810 3580 33815 3600
rect 33835 3580 33840 3600
rect 33810 3550 33840 3580
rect 33810 3530 33815 3550
rect 33835 3530 33840 3550
rect 33810 3500 33840 3530
rect 33810 3480 33815 3500
rect 33835 3480 33840 3500
rect 33810 3450 33840 3480
rect 33810 3430 33815 3450
rect 33835 3430 33840 3450
rect 33810 3400 33840 3430
rect 33810 3380 33815 3400
rect 33835 3380 33840 3400
rect 33810 3350 33840 3380
rect 33810 3330 33815 3350
rect 33835 3330 33840 3350
rect 33810 3300 33840 3330
rect 33810 3280 33815 3300
rect 33835 3280 33840 3300
rect 33810 3250 33840 3280
rect 33810 3230 33815 3250
rect 33835 3230 33840 3250
rect 33810 3200 33840 3230
rect 33810 3180 33815 3200
rect 33835 3180 33840 3200
rect 33810 3150 33840 3180
rect 33810 3130 33815 3150
rect 33835 3130 33840 3150
rect 33810 3100 33840 3130
rect 33810 3080 33815 3100
rect 33835 3080 33840 3100
rect 33210 3050 33230 3070
rect 33320 3050 33340 3070
rect 33430 3050 33450 3070
rect 33540 3050 33560 3070
rect 33650 3050 33670 3070
rect 33760 3050 33780 3070
rect 33150 3020 33155 3040
rect 33175 3020 33180 3040
rect 33150 3010 33180 3020
rect 33200 3040 33240 3050
rect 33200 3020 33210 3040
rect 33230 3020 33240 3040
rect 33200 3010 33240 3020
rect 33310 3040 33350 3050
rect 33310 3020 33320 3040
rect 33340 3020 33350 3040
rect 33310 3010 33350 3020
rect 33420 3040 33460 3050
rect 33420 3020 33430 3040
rect 33450 3020 33460 3040
rect 33420 3010 33460 3020
rect 33530 3040 33570 3050
rect 33530 3020 33540 3040
rect 33560 3020 33570 3040
rect 33530 3010 33570 3020
rect 33588 3040 33622 3050
rect 33588 3020 33596 3040
rect 33614 3020 33622 3040
rect 33588 3010 33622 3020
rect 33640 3040 33680 3050
rect 33640 3020 33650 3040
rect 33670 3020 33680 3040
rect 33640 3010 33680 3020
rect 33750 3040 33790 3050
rect 33750 3020 33760 3040
rect 33780 3020 33790 3040
rect 33750 3010 33790 3020
rect 33810 3040 33840 3080
rect 33810 3020 33815 3040
rect 33835 3020 33840 3040
rect 33810 3010 33840 3020
rect 33875 3410 33895 3740
rect 33155 2990 33175 3010
rect 33815 2990 33835 3010
rect 33875 2990 33895 3315
rect 33095 2970 33455 2990
rect 33535 2970 33895 2990
rect 34035 3680 34315 3700
rect 34035 3375 34055 3680
rect 34105 3655 34246 3660
rect 34105 3625 34111 3655
rect 34141 3625 34160 3655
rect 34190 3625 34210 3655
rect 34240 3625 34246 3655
rect 34105 3620 34246 3625
rect 34035 2995 34055 3280
rect 34295 3375 34315 3680
rect 34105 3050 34246 3055
rect 34105 3020 34111 3050
rect 34141 3020 34160 3050
rect 34190 3020 34210 3050
rect 34240 3020 34246 3050
rect 34105 3015 34246 3020
rect 34295 2995 34315 3280
rect 34035 2975 34135 2995
rect 34215 2985 34315 2995
rect 34215 2975 34245 2985
rect 29525 2955 29565 2965
rect 30285 2960 30295 2970
rect 30315 2960 30325 2970
rect 30285 2950 30325 2960
rect 33475 2960 33485 2970
rect 33505 2960 33515 2970
rect 33475 2950 33515 2960
rect 34235 2965 34245 2975
rect 34265 2975 34315 2985
rect 34265 2965 34275 2975
rect 34235 2955 34275 2965
rect 30955 2920 31345 2940
rect 31425 2920 31815 2940
rect 30285 2810 30325 2820
rect 30285 2800 30295 2810
rect 30315 2800 30325 2810
rect 29905 2780 30265 2800
rect 30345 2780 30705 2800
rect 29525 2679 29565 2689
rect 29525 2669 29535 2679
rect 29555 2669 29565 2679
rect 29400 2649 29535 2669
rect 29615 2649 29755 2669
rect 29400 2335 29420 2649
rect 29470 2609 29685 2629
rect 29470 2589 29505 2609
rect 29650 2589 29685 2609
rect 29565 2539 29590 2589
rect 29400 1925 29420 2255
rect 29735 2335 29755 2649
rect 29905 2645 29925 2780
rect 30010 2750 30050 2760
rect 30010 2730 30020 2750
rect 30040 2730 30050 2750
rect 30010 2720 30050 2730
rect 30120 2750 30160 2760
rect 30120 2730 30130 2750
rect 30150 2730 30160 2750
rect 30120 2720 30160 2730
rect 30230 2750 30270 2760
rect 30230 2730 30240 2750
rect 30260 2730 30270 2750
rect 30230 2720 30270 2730
rect 30340 2750 30380 2760
rect 30340 2730 30350 2750
rect 30370 2730 30380 2750
rect 30340 2720 30380 2730
rect 30450 2750 30490 2760
rect 30450 2730 30460 2750
rect 30480 2730 30490 2750
rect 30450 2720 30490 2730
rect 30560 2750 30600 2760
rect 30560 2730 30570 2750
rect 30590 2730 30600 2750
rect 30560 2720 30600 2730
rect 30020 2700 30040 2720
rect 30130 2700 30150 2720
rect 30240 2700 30260 2720
rect 30350 2700 30370 2720
rect 30460 2700 30480 2720
rect 30570 2700 30590 2720
rect 29905 2430 29925 2565
rect 29960 2690 29990 2700
rect 29960 2670 29965 2690
rect 29985 2670 29990 2690
rect 29960 2640 29990 2670
rect 29960 2620 29965 2640
rect 29985 2620 29990 2640
rect 29960 2590 29990 2620
rect 29960 2570 29965 2590
rect 29985 2570 29990 2590
rect 29960 2540 29990 2570
rect 29960 2520 29965 2540
rect 29985 2520 29990 2540
rect 29960 2480 29990 2520
rect 30015 2690 30045 2700
rect 30015 2670 30020 2690
rect 30040 2670 30045 2690
rect 30015 2640 30045 2670
rect 30015 2620 30020 2640
rect 30040 2620 30045 2640
rect 30015 2590 30045 2620
rect 30015 2570 30020 2590
rect 30040 2570 30045 2590
rect 30015 2540 30045 2570
rect 30015 2520 30020 2540
rect 30040 2520 30045 2540
rect 30015 2510 30045 2520
rect 30070 2690 30100 2700
rect 30070 2670 30075 2690
rect 30095 2670 30100 2690
rect 30070 2640 30100 2670
rect 30070 2620 30075 2640
rect 30095 2620 30100 2640
rect 30070 2590 30100 2620
rect 30070 2570 30075 2590
rect 30095 2570 30100 2590
rect 30070 2540 30100 2570
rect 30070 2520 30075 2540
rect 30095 2520 30100 2540
rect 30070 2510 30100 2520
rect 30125 2690 30155 2700
rect 30125 2670 30130 2690
rect 30150 2670 30155 2690
rect 30125 2640 30155 2670
rect 30125 2620 30130 2640
rect 30150 2620 30155 2640
rect 30125 2590 30155 2620
rect 30125 2570 30130 2590
rect 30150 2570 30155 2590
rect 30125 2540 30155 2570
rect 30125 2520 30130 2540
rect 30150 2520 30155 2540
rect 30125 2510 30155 2520
rect 30180 2690 30210 2700
rect 30180 2670 30185 2690
rect 30205 2670 30210 2690
rect 30180 2640 30210 2670
rect 30180 2620 30185 2640
rect 30205 2620 30210 2640
rect 30180 2590 30210 2620
rect 30180 2570 30185 2590
rect 30205 2570 30210 2590
rect 30180 2540 30210 2570
rect 30180 2520 30185 2540
rect 30205 2520 30210 2540
rect 30180 2510 30210 2520
rect 30235 2690 30265 2700
rect 30235 2670 30240 2690
rect 30260 2670 30265 2690
rect 30235 2640 30265 2670
rect 30235 2620 30240 2640
rect 30260 2620 30265 2640
rect 30235 2590 30265 2620
rect 30235 2570 30240 2590
rect 30260 2570 30265 2590
rect 30235 2540 30265 2570
rect 30235 2520 30240 2540
rect 30260 2520 30265 2540
rect 30235 2510 30265 2520
rect 30290 2690 30320 2700
rect 30290 2670 30295 2690
rect 30315 2670 30320 2690
rect 30290 2640 30320 2670
rect 30290 2620 30295 2640
rect 30315 2620 30320 2640
rect 30290 2590 30320 2620
rect 30290 2570 30295 2590
rect 30315 2570 30320 2590
rect 30290 2540 30320 2570
rect 30290 2520 30295 2540
rect 30315 2520 30320 2540
rect 30290 2510 30320 2520
rect 30345 2690 30375 2700
rect 30345 2670 30350 2690
rect 30370 2670 30375 2690
rect 30345 2640 30375 2670
rect 30345 2620 30350 2640
rect 30370 2620 30375 2640
rect 30345 2590 30375 2620
rect 30345 2570 30350 2590
rect 30370 2570 30375 2590
rect 30345 2540 30375 2570
rect 30345 2520 30350 2540
rect 30370 2520 30375 2540
rect 30345 2510 30375 2520
rect 30400 2690 30430 2700
rect 30400 2670 30405 2690
rect 30425 2670 30430 2690
rect 30400 2640 30430 2670
rect 30400 2620 30405 2640
rect 30425 2620 30430 2640
rect 30400 2590 30430 2620
rect 30400 2570 30405 2590
rect 30425 2570 30430 2590
rect 30400 2540 30430 2570
rect 30400 2520 30405 2540
rect 30425 2520 30430 2540
rect 30400 2510 30430 2520
rect 30455 2690 30485 2700
rect 30455 2670 30460 2690
rect 30480 2670 30485 2690
rect 30455 2640 30485 2670
rect 30455 2620 30460 2640
rect 30480 2620 30485 2640
rect 30455 2590 30485 2620
rect 30455 2570 30460 2590
rect 30480 2570 30485 2590
rect 30455 2540 30485 2570
rect 30455 2520 30460 2540
rect 30480 2520 30485 2540
rect 30455 2510 30485 2520
rect 30510 2690 30540 2700
rect 30510 2670 30515 2690
rect 30535 2670 30540 2690
rect 30510 2640 30540 2670
rect 30510 2620 30515 2640
rect 30535 2620 30540 2640
rect 30510 2590 30540 2620
rect 30510 2570 30515 2590
rect 30535 2570 30540 2590
rect 30510 2540 30540 2570
rect 30510 2520 30515 2540
rect 30535 2520 30540 2540
rect 30510 2510 30540 2520
rect 30565 2690 30595 2700
rect 30565 2670 30570 2690
rect 30590 2670 30595 2690
rect 30565 2640 30595 2670
rect 30565 2620 30570 2640
rect 30590 2620 30595 2640
rect 30565 2590 30595 2620
rect 30565 2570 30570 2590
rect 30590 2570 30595 2590
rect 30565 2540 30595 2570
rect 30565 2520 30570 2540
rect 30590 2520 30595 2540
rect 30565 2510 30595 2520
rect 30620 2690 30650 2700
rect 30620 2670 30625 2690
rect 30645 2670 30650 2690
rect 30620 2640 30650 2670
rect 30620 2620 30625 2640
rect 30645 2620 30650 2640
rect 30620 2590 30650 2620
rect 30620 2570 30625 2590
rect 30645 2570 30650 2590
rect 30620 2540 30650 2570
rect 30620 2520 30625 2540
rect 30645 2520 30650 2540
rect 30075 2490 30095 2510
rect 30185 2490 30205 2510
rect 30295 2490 30315 2510
rect 30405 2490 30425 2510
rect 30515 2490 30535 2510
rect 29960 2460 29965 2480
rect 29985 2460 29990 2480
rect 29960 2450 29990 2460
rect 30065 2480 30105 2490
rect 30065 2460 30075 2480
rect 30095 2460 30105 2480
rect 30065 2450 30105 2460
rect 30175 2480 30215 2490
rect 30175 2460 30185 2480
rect 30205 2460 30215 2480
rect 30175 2450 30215 2460
rect 30285 2480 30325 2490
rect 30285 2460 30295 2480
rect 30315 2460 30325 2480
rect 30285 2450 30325 2460
rect 30395 2480 30435 2490
rect 30395 2460 30405 2480
rect 30425 2460 30435 2480
rect 30395 2450 30435 2460
rect 30453 2480 30487 2490
rect 30453 2460 30461 2480
rect 30479 2460 30487 2480
rect 30453 2450 30487 2460
rect 30505 2480 30545 2490
rect 30505 2460 30515 2480
rect 30535 2460 30545 2480
rect 30505 2450 30545 2460
rect 30620 2480 30650 2520
rect 30620 2460 30625 2480
rect 30645 2460 30650 2480
rect 30620 2450 30650 2460
rect 30685 2645 30705 2780
rect 29965 2430 29985 2450
rect 30625 2430 30645 2450
rect 30685 2430 30705 2565
rect 29905 2410 30265 2430
rect 30345 2410 30705 2430
rect 30955 2710 30975 2920
rect 31375 2900 31395 2920
rect 31125 2890 31165 2900
rect 31125 2870 31135 2890
rect 31155 2870 31165 2890
rect 31125 2860 31165 2870
rect 31245 2890 31285 2900
rect 31245 2870 31255 2890
rect 31275 2870 31285 2890
rect 31245 2860 31285 2870
rect 31365 2890 31405 2900
rect 31365 2870 31375 2890
rect 31395 2870 31405 2890
rect 31365 2860 31405 2870
rect 31485 2890 31525 2900
rect 31485 2870 31495 2890
rect 31515 2870 31525 2890
rect 31485 2860 31525 2870
rect 31605 2890 31645 2900
rect 31605 2870 31615 2890
rect 31635 2870 31645 2890
rect 31605 2860 31645 2870
rect 31135 2840 31155 2860
rect 31255 2840 31275 2860
rect 31375 2840 31395 2860
rect 31495 2840 31515 2860
rect 31615 2840 31635 2860
rect 30955 2420 30975 2630
rect 31010 2830 31040 2840
rect 31010 2810 31015 2830
rect 31035 2810 31040 2830
rect 31010 2780 31040 2810
rect 31010 2760 31015 2780
rect 31035 2760 31040 2780
rect 31010 2730 31040 2760
rect 31010 2710 31015 2730
rect 31035 2710 31040 2730
rect 31010 2680 31040 2710
rect 31010 2660 31015 2680
rect 31035 2660 31040 2680
rect 31010 2630 31040 2660
rect 31010 2610 31015 2630
rect 31035 2610 31040 2630
rect 31010 2580 31040 2610
rect 31010 2560 31015 2580
rect 31035 2560 31040 2580
rect 31010 2530 31040 2560
rect 31010 2510 31015 2530
rect 31035 2510 31040 2530
rect 31010 2470 31040 2510
rect 31070 2830 31100 2840
rect 31070 2810 31075 2830
rect 31095 2810 31100 2830
rect 31070 2780 31100 2810
rect 31070 2760 31075 2780
rect 31095 2760 31100 2780
rect 31070 2730 31100 2760
rect 31070 2710 31075 2730
rect 31095 2710 31100 2730
rect 31070 2680 31100 2710
rect 31070 2660 31075 2680
rect 31095 2660 31100 2680
rect 31070 2630 31100 2660
rect 31070 2610 31075 2630
rect 31095 2610 31100 2630
rect 31070 2580 31100 2610
rect 31070 2560 31075 2580
rect 31095 2560 31100 2580
rect 31070 2530 31100 2560
rect 31070 2510 31075 2530
rect 31095 2510 31100 2530
rect 31070 2500 31100 2510
rect 31130 2830 31160 2840
rect 31130 2810 31135 2830
rect 31155 2810 31160 2830
rect 31130 2780 31160 2810
rect 31130 2760 31135 2780
rect 31155 2760 31160 2780
rect 31130 2730 31160 2760
rect 31130 2710 31135 2730
rect 31155 2710 31160 2730
rect 31130 2680 31160 2710
rect 31130 2660 31135 2680
rect 31155 2660 31160 2680
rect 31130 2630 31160 2660
rect 31130 2610 31135 2630
rect 31155 2610 31160 2630
rect 31130 2580 31160 2610
rect 31130 2560 31135 2580
rect 31155 2560 31160 2580
rect 31130 2530 31160 2560
rect 31130 2510 31135 2530
rect 31155 2510 31160 2530
rect 31130 2500 31160 2510
rect 31190 2830 31220 2840
rect 31190 2810 31195 2830
rect 31215 2810 31220 2830
rect 31190 2780 31220 2810
rect 31190 2760 31195 2780
rect 31215 2760 31220 2780
rect 31190 2730 31220 2760
rect 31190 2710 31195 2730
rect 31215 2710 31220 2730
rect 31190 2680 31220 2710
rect 31190 2660 31195 2680
rect 31215 2660 31220 2680
rect 31190 2630 31220 2660
rect 31190 2610 31195 2630
rect 31215 2610 31220 2630
rect 31190 2580 31220 2610
rect 31190 2560 31195 2580
rect 31215 2560 31220 2580
rect 31190 2530 31220 2560
rect 31190 2510 31195 2530
rect 31215 2510 31220 2530
rect 31190 2500 31220 2510
rect 31250 2830 31280 2840
rect 31250 2810 31255 2830
rect 31275 2810 31280 2830
rect 31250 2780 31280 2810
rect 31250 2760 31255 2780
rect 31275 2760 31280 2780
rect 31250 2730 31280 2760
rect 31250 2710 31255 2730
rect 31275 2710 31280 2730
rect 31250 2680 31280 2710
rect 31250 2660 31255 2680
rect 31275 2660 31280 2680
rect 31250 2630 31280 2660
rect 31250 2610 31255 2630
rect 31275 2610 31280 2630
rect 31250 2580 31280 2610
rect 31250 2560 31255 2580
rect 31275 2560 31280 2580
rect 31250 2530 31280 2560
rect 31250 2510 31255 2530
rect 31275 2510 31280 2530
rect 31250 2500 31280 2510
rect 31310 2830 31340 2840
rect 31310 2810 31315 2830
rect 31335 2810 31340 2830
rect 31310 2780 31340 2810
rect 31310 2760 31315 2780
rect 31335 2760 31340 2780
rect 31310 2730 31340 2760
rect 31310 2710 31315 2730
rect 31335 2710 31340 2730
rect 31310 2680 31340 2710
rect 31310 2660 31315 2680
rect 31335 2660 31340 2680
rect 31310 2630 31340 2660
rect 31310 2610 31315 2630
rect 31335 2610 31340 2630
rect 31310 2580 31340 2610
rect 31310 2560 31315 2580
rect 31335 2560 31340 2580
rect 31310 2530 31340 2560
rect 31310 2510 31315 2530
rect 31335 2510 31340 2530
rect 31310 2500 31340 2510
rect 31370 2830 31400 2840
rect 31370 2810 31375 2830
rect 31395 2810 31400 2830
rect 31370 2780 31400 2810
rect 31370 2760 31375 2780
rect 31395 2760 31400 2780
rect 31370 2730 31400 2760
rect 31370 2710 31375 2730
rect 31395 2710 31400 2730
rect 31370 2680 31400 2710
rect 31370 2660 31375 2680
rect 31395 2660 31400 2680
rect 31370 2630 31400 2660
rect 31370 2610 31375 2630
rect 31395 2610 31400 2630
rect 31370 2580 31400 2610
rect 31370 2560 31375 2580
rect 31395 2560 31400 2580
rect 31370 2530 31400 2560
rect 31370 2510 31375 2530
rect 31395 2510 31400 2530
rect 31370 2500 31400 2510
rect 31430 2830 31460 2840
rect 31430 2810 31435 2830
rect 31455 2810 31460 2830
rect 31430 2780 31460 2810
rect 31430 2760 31435 2780
rect 31455 2760 31460 2780
rect 31430 2730 31460 2760
rect 31430 2710 31435 2730
rect 31455 2710 31460 2730
rect 31430 2680 31460 2710
rect 31430 2660 31435 2680
rect 31455 2660 31460 2680
rect 31430 2630 31460 2660
rect 31430 2610 31435 2630
rect 31455 2610 31460 2630
rect 31430 2580 31460 2610
rect 31430 2560 31435 2580
rect 31455 2560 31460 2580
rect 31430 2530 31460 2560
rect 31430 2510 31435 2530
rect 31455 2510 31460 2530
rect 31430 2500 31460 2510
rect 31490 2830 31520 2840
rect 31490 2810 31495 2830
rect 31515 2810 31520 2830
rect 31490 2780 31520 2810
rect 31490 2760 31495 2780
rect 31515 2760 31520 2780
rect 31490 2730 31520 2760
rect 31490 2710 31495 2730
rect 31515 2710 31520 2730
rect 31490 2680 31520 2710
rect 31490 2660 31495 2680
rect 31515 2660 31520 2680
rect 31490 2630 31520 2660
rect 31490 2610 31495 2630
rect 31515 2610 31520 2630
rect 31490 2580 31520 2610
rect 31490 2560 31495 2580
rect 31515 2560 31520 2580
rect 31490 2530 31520 2560
rect 31490 2510 31495 2530
rect 31515 2510 31520 2530
rect 31490 2500 31520 2510
rect 31550 2830 31580 2840
rect 31550 2810 31555 2830
rect 31575 2810 31580 2830
rect 31550 2780 31580 2810
rect 31550 2760 31555 2780
rect 31575 2760 31580 2780
rect 31550 2730 31580 2760
rect 31550 2710 31555 2730
rect 31575 2710 31580 2730
rect 31550 2680 31580 2710
rect 31550 2660 31555 2680
rect 31575 2660 31580 2680
rect 31550 2630 31580 2660
rect 31550 2610 31555 2630
rect 31575 2610 31580 2630
rect 31550 2580 31580 2610
rect 31550 2560 31555 2580
rect 31575 2560 31580 2580
rect 31550 2530 31580 2560
rect 31550 2510 31555 2530
rect 31575 2510 31580 2530
rect 31550 2500 31580 2510
rect 31610 2830 31640 2840
rect 31610 2810 31615 2830
rect 31635 2810 31640 2830
rect 31610 2780 31640 2810
rect 31610 2760 31615 2780
rect 31635 2760 31640 2780
rect 31610 2730 31640 2760
rect 31610 2710 31615 2730
rect 31635 2710 31640 2730
rect 31610 2680 31640 2710
rect 31610 2660 31615 2680
rect 31635 2660 31640 2680
rect 31610 2630 31640 2660
rect 31610 2610 31615 2630
rect 31635 2610 31640 2630
rect 31610 2580 31640 2610
rect 31610 2560 31615 2580
rect 31635 2560 31640 2580
rect 31610 2530 31640 2560
rect 31610 2510 31615 2530
rect 31635 2510 31640 2530
rect 31610 2500 31640 2510
rect 31670 2830 31700 2840
rect 31670 2810 31675 2830
rect 31695 2810 31700 2830
rect 31670 2780 31700 2810
rect 31670 2760 31675 2780
rect 31695 2760 31700 2780
rect 31670 2730 31700 2760
rect 31670 2710 31675 2730
rect 31695 2710 31700 2730
rect 31670 2680 31700 2710
rect 31670 2660 31675 2680
rect 31695 2660 31700 2680
rect 31670 2630 31700 2660
rect 31670 2610 31675 2630
rect 31695 2610 31700 2630
rect 31670 2580 31700 2610
rect 31670 2560 31675 2580
rect 31695 2560 31700 2580
rect 31670 2530 31700 2560
rect 31670 2510 31675 2530
rect 31695 2510 31700 2530
rect 31670 2500 31700 2510
rect 31730 2830 31760 2840
rect 31730 2810 31735 2830
rect 31755 2810 31760 2830
rect 31730 2780 31760 2810
rect 31730 2760 31735 2780
rect 31755 2760 31760 2780
rect 31730 2730 31760 2760
rect 31730 2710 31735 2730
rect 31755 2710 31760 2730
rect 31730 2680 31760 2710
rect 31730 2660 31735 2680
rect 31755 2660 31760 2680
rect 31730 2630 31760 2660
rect 31730 2610 31735 2630
rect 31755 2610 31760 2630
rect 31730 2580 31760 2610
rect 31730 2560 31735 2580
rect 31755 2560 31760 2580
rect 31730 2530 31760 2560
rect 31730 2510 31735 2530
rect 31755 2510 31760 2530
rect 31075 2480 31095 2500
rect 31195 2480 31215 2500
rect 31315 2480 31335 2500
rect 31435 2480 31455 2500
rect 31555 2480 31575 2500
rect 31675 2480 31695 2500
rect 31010 2450 31015 2470
rect 31035 2450 31040 2470
rect 31010 2440 31040 2450
rect 31065 2470 31105 2480
rect 31065 2450 31075 2470
rect 31095 2450 31105 2470
rect 31065 2440 31105 2450
rect 31185 2470 31225 2480
rect 31185 2450 31195 2470
rect 31215 2450 31225 2470
rect 31185 2440 31225 2450
rect 31305 2470 31345 2480
rect 31305 2450 31315 2470
rect 31335 2450 31345 2470
rect 31305 2440 31345 2450
rect 31368 2470 31402 2480
rect 31368 2450 31376 2470
rect 31394 2450 31402 2470
rect 31368 2440 31402 2450
rect 31425 2470 31465 2480
rect 31425 2450 31435 2470
rect 31455 2450 31465 2470
rect 31425 2440 31465 2450
rect 31545 2470 31585 2480
rect 31545 2450 31555 2470
rect 31575 2450 31585 2470
rect 31545 2440 31585 2450
rect 31665 2470 31705 2480
rect 31665 2450 31675 2470
rect 31695 2450 31705 2470
rect 31665 2440 31705 2450
rect 31730 2470 31760 2510
rect 31730 2450 31735 2470
rect 31755 2450 31760 2470
rect 31730 2440 31760 2450
rect 31795 2710 31815 2920
rect 31015 2420 31035 2440
rect 31735 2420 31755 2440
rect 31795 2420 31815 2630
rect 30955 2400 31345 2420
rect 31425 2400 31815 2420
rect 31985 2920 32375 2940
rect 32455 2920 32845 2940
rect 31985 2710 32005 2920
rect 32405 2900 32425 2920
rect 32155 2890 32195 2900
rect 32155 2870 32165 2890
rect 32185 2870 32195 2890
rect 32155 2860 32195 2870
rect 32275 2890 32315 2900
rect 32275 2870 32285 2890
rect 32305 2870 32315 2890
rect 32275 2860 32315 2870
rect 32395 2890 32435 2900
rect 32395 2870 32405 2890
rect 32425 2870 32435 2890
rect 32395 2860 32435 2870
rect 32515 2890 32555 2900
rect 32515 2870 32525 2890
rect 32545 2870 32555 2890
rect 32515 2860 32555 2870
rect 32635 2890 32675 2900
rect 32635 2870 32645 2890
rect 32665 2870 32675 2890
rect 32635 2860 32675 2870
rect 32165 2840 32185 2860
rect 32285 2840 32305 2860
rect 32405 2840 32425 2860
rect 32525 2840 32545 2860
rect 32645 2840 32665 2860
rect 31985 2420 32005 2630
rect 32040 2830 32070 2840
rect 32040 2810 32045 2830
rect 32065 2810 32070 2830
rect 32040 2780 32070 2810
rect 32040 2760 32045 2780
rect 32065 2760 32070 2780
rect 32040 2730 32070 2760
rect 32040 2710 32045 2730
rect 32065 2710 32070 2730
rect 32040 2680 32070 2710
rect 32040 2660 32045 2680
rect 32065 2660 32070 2680
rect 32040 2630 32070 2660
rect 32040 2610 32045 2630
rect 32065 2610 32070 2630
rect 32040 2580 32070 2610
rect 32040 2560 32045 2580
rect 32065 2560 32070 2580
rect 32040 2530 32070 2560
rect 32040 2510 32045 2530
rect 32065 2510 32070 2530
rect 32040 2470 32070 2510
rect 32100 2830 32130 2840
rect 32100 2810 32105 2830
rect 32125 2810 32130 2830
rect 32100 2780 32130 2810
rect 32100 2760 32105 2780
rect 32125 2760 32130 2780
rect 32100 2730 32130 2760
rect 32100 2710 32105 2730
rect 32125 2710 32130 2730
rect 32100 2680 32130 2710
rect 32100 2660 32105 2680
rect 32125 2660 32130 2680
rect 32100 2630 32130 2660
rect 32100 2610 32105 2630
rect 32125 2610 32130 2630
rect 32100 2580 32130 2610
rect 32100 2560 32105 2580
rect 32125 2560 32130 2580
rect 32100 2530 32130 2560
rect 32100 2510 32105 2530
rect 32125 2510 32130 2530
rect 32100 2500 32130 2510
rect 32160 2830 32190 2840
rect 32160 2810 32165 2830
rect 32185 2810 32190 2830
rect 32160 2780 32190 2810
rect 32160 2760 32165 2780
rect 32185 2760 32190 2780
rect 32160 2730 32190 2760
rect 32160 2710 32165 2730
rect 32185 2710 32190 2730
rect 32160 2680 32190 2710
rect 32160 2660 32165 2680
rect 32185 2660 32190 2680
rect 32160 2630 32190 2660
rect 32160 2610 32165 2630
rect 32185 2610 32190 2630
rect 32160 2580 32190 2610
rect 32160 2560 32165 2580
rect 32185 2560 32190 2580
rect 32160 2530 32190 2560
rect 32160 2510 32165 2530
rect 32185 2510 32190 2530
rect 32160 2500 32190 2510
rect 32220 2830 32250 2840
rect 32220 2810 32225 2830
rect 32245 2810 32250 2830
rect 32220 2780 32250 2810
rect 32220 2760 32225 2780
rect 32245 2760 32250 2780
rect 32220 2730 32250 2760
rect 32220 2710 32225 2730
rect 32245 2710 32250 2730
rect 32220 2680 32250 2710
rect 32220 2660 32225 2680
rect 32245 2660 32250 2680
rect 32220 2630 32250 2660
rect 32220 2610 32225 2630
rect 32245 2610 32250 2630
rect 32220 2580 32250 2610
rect 32220 2560 32225 2580
rect 32245 2560 32250 2580
rect 32220 2530 32250 2560
rect 32220 2510 32225 2530
rect 32245 2510 32250 2530
rect 32220 2500 32250 2510
rect 32280 2830 32310 2840
rect 32280 2810 32285 2830
rect 32305 2810 32310 2830
rect 32280 2780 32310 2810
rect 32280 2760 32285 2780
rect 32305 2760 32310 2780
rect 32280 2730 32310 2760
rect 32280 2710 32285 2730
rect 32305 2710 32310 2730
rect 32280 2680 32310 2710
rect 32280 2660 32285 2680
rect 32305 2660 32310 2680
rect 32280 2630 32310 2660
rect 32280 2610 32285 2630
rect 32305 2610 32310 2630
rect 32280 2580 32310 2610
rect 32280 2560 32285 2580
rect 32305 2560 32310 2580
rect 32280 2530 32310 2560
rect 32280 2510 32285 2530
rect 32305 2510 32310 2530
rect 32280 2500 32310 2510
rect 32340 2830 32370 2840
rect 32340 2810 32345 2830
rect 32365 2810 32370 2830
rect 32340 2780 32370 2810
rect 32340 2760 32345 2780
rect 32365 2760 32370 2780
rect 32340 2730 32370 2760
rect 32340 2710 32345 2730
rect 32365 2710 32370 2730
rect 32340 2680 32370 2710
rect 32340 2660 32345 2680
rect 32365 2660 32370 2680
rect 32340 2630 32370 2660
rect 32340 2610 32345 2630
rect 32365 2610 32370 2630
rect 32340 2580 32370 2610
rect 32340 2560 32345 2580
rect 32365 2560 32370 2580
rect 32340 2530 32370 2560
rect 32340 2510 32345 2530
rect 32365 2510 32370 2530
rect 32340 2500 32370 2510
rect 32400 2830 32430 2840
rect 32400 2810 32405 2830
rect 32425 2810 32430 2830
rect 32400 2780 32430 2810
rect 32400 2760 32405 2780
rect 32425 2760 32430 2780
rect 32400 2730 32430 2760
rect 32400 2710 32405 2730
rect 32425 2710 32430 2730
rect 32400 2680 32430 2710
rect 32400 2660 32405 2680
rect 32425 2660 32430 2680
rect 32400 2630 32430 2660
rect 32400 2610 32405 2630
rect 32425 2610 32430 2630
rect 32400 2580 32430 2610
rect 32400 2560 32405 2580
rect 32425 2560 32430 2580
rect 32400 2530 32430 2560
rect 32400 2510 32405 2530
rect 32425 2510 32430 2530
rect 32400 2500 32430 2510
rect 32460 2830 32490 2840
rect 32460 2810 32465 2830
rect 32485 2810 32490 2830
rect 32460 2780 32490 2810
rect 32460 2760 32465 2780
rect 32485 2760 32490 2780
rect 32460 2730 32490 2760
rect 32460 2710 32465 2730
rect 32485 2710 32490 2730
rect 32460 2680 32490 2710
rect 32460 2660 32465 2680
rect 32485 2660 32490 2680
rect 32460 2630 32490 2660
rect 32460 2610 32465 2630
rect 32485 2610 32490 2630
rect 32460 2580 32490 2610
rect 32460 2560 32465 2580
rect 32485 2560 32490 2580
rect 32460 2530 32490 2560
rect 32460 2510 32465 2530
rect 32485 2510 32490 2530
rect 32460 2500 32490 2510
rect 32520 2830 32550 2840
rect 32520 2810 32525 2830
rect 32545 2810 32550 2830
rect 32520 2780 32550 2810
rect 32520 2760 32525 2780
rect 32545 2760 32550 2780
rect 32520 2730 32550 2760
rect 32520 2710 32525 2730
rect 32545 2710 32550 2730
rect 32520 2680 32550 2710
rect 32520 2660 32525 2680
rect 32545 2660 32550 2680
rect 32520 2630 32550 2660
rect 32520 2610 32525 2630
rect 32545 2610 32550 2630
rect 32520 2580 32550 2610
rect 32520 2560 32525 2580
rect 32545 2560 32550 2580
rect 32520 2530 32550 2560
rect 32520 2510 32525 2530
rect 32545 2510 32550 2530
rect 32520 2500 32550 2510
rect 32580 2830 32610 2840
rect 32580 2810 32585 2830
rect 32605 2810 32610 2830
rect 32580 2780 32610 2810
rect 32580 2760 32585 2780
rect 32605 2760 32610 2780
rect 32580 2730 32610 2760
rect 32580 2710 32585 2730
rect 32605 2710 32610 2730
rect 32580 2680 32610 2710
rect 32580 2660 32585 2680
rect 32605 2660 32610 2680
rect 32580 2630 32610 2660
rect 32580 2610 32585 2630
rect 32605 2610 32610 2630
rect 32580 2580 32610 2610
rect 32580 2560 32585 2580
rect 32605 2560 32610 2580
rect 32580 2530 32610 2560
rect 32580 2510 32585 2530
rect 32605 2510 32610 2530
rect 32580 2500 32610 2510
rect 32640 2830 32670 2840
rect 32640 2810 32645 2830
rect 32665 2810 32670 2830
rect 32640 2780 32670 2810
rect 32640 2760 32645 2780
rect 32665 2760 32670 2780
rect 32640 2730 32670 2760
rect 32640 2710 32645 2730
rect 32665 2710 32670 2730
rect 32640 2680 32670 2710
rect 32640 2660 32645 2680
rect 32665 2660 32670 2680
rect 32640 2630 32670 2660
rect 32640 2610 32645 2630
rect 32665 2610 32670 2630
rect 32640 2580 32670 2610
rect 32640 2560 32645 2580
rect 32665 2560 32670 2580
rect 32640 2530 32670 2560
rect 32640 2510 32645 2530
rect 32665 2510 32670 2530
rect 32640 2500 32670 2510
rect 32700 2830 32730 2840
rect 32700 2810 32705 2830
rect 32725 2810 32730 2830
rect 32700 2780 32730 2810
rect 32700 2760 32705 2780
rect 32725 2760 32730 2780
rect 32700 2730 32730 2760
rect 32700 2710 32705 2730
rect 32725 2710 32730 2730
rect 32700 2680 32730 2710
rect 32700 2660 32705 2680
rect 32725 2660 32730 2680
rect 32700 2630 32730 2660
rect 32700 2610 32705 2630
rect 32725 2610 32730 2630
rect 32700 2580 32730 2610
rect 32700 2560 32705 2580
rect 32725 2560 32730 2580
rect 32700 2530 32730 2560
rect 32700 2510 32705 2530
rect 32725 2510 32730 2530
rect 32700 2500 32730 2510
rect 32760 2830 32790 2840
rect 32760 2810 32765 2830
rect 32785 2810 32790 2830
rect 32760 2780 32790 2810
rect 32760 2760 32765 2780
rect 32785 2760 32790 2780
rect 32760 2730 32790 2760
rect 32760 2710 32765 2730
rect 32785 2710 32790 2730
rect 32760 2680 32790 2710
rect 32760 2660 32765 2680
rect 32785 2660 32790 2680
rect 32760 2630 32790 2660
rect 32760 2610 32765 2630
rect 32785 2610 32790 2630
rect 32760 2580 32790 2610
rect 32760 2560 32765 2580
rect 32785 2560 32790 2580
rect 32760 2530 32790 2560
rect 32760 2510 32765 2530
rect 32785 2510 32790 2530
rect 32105 2480 32125 2500
rect 32225 2480 32245 2500
rect 32345 2480 32365 2500
rect 32465 2480 32485 2500
rect 32585 2480 32605 2500
rect 32705 2480 32725 2500
rect 32040 2450 32045 2470
rect 32065 2450 32070 2470
rect 32040 2440 32070 2450
rect 32095 2470 32135 2480
rect 32095 2450 32105 2470
rect 32125 2450 32135 2470
rect 32095 2440 32135 2450
rect 32215 2470 32255 2480
rect 32215 2450 32225 2470
rect 32245 2450 32255 2470
rect 32215 2440 32255 2450
rect 32335 2470 32375 2480
rect 32335 2450 32345 2470
rect 32365 2450 32375 2470
rect 32335 2440 32375 2450
rect 32398 2470 32432 2480
rect 32398 2450 32406 2470
rect 32424 2450 32432 2470
rect 32398 2440 32432 2450
rect 32455 2470 32495 2480
rect 32455 2450 32465 2470
rect 32485 2450 32495 2470
rect 32455 2440 32495 2450
rect 32575 2470 32615 2480
rect 32575 2450 32585 2470
rect 32605 2450 32615 2470
rect 32575 2440 32615 2450
rect 32695 2470 32735 2480
rect 32695 2450 32705 2470
rect 32725 2450 32735 2470
rect 32695 2440 32735 2450
rect 32760 2470 32790 2510
rect 32760 2450 32765 2470
rect 32785 2450 32790 2470
rect 32760 2440 32790 2450
rect 32825 2710 32845 2920
rect 33475 2810 33515 2820
rect 33475 2800 33485 2810
rect 33505 2800 33515 2810
rect 32045 2420 32065 2440
rect 32765 2420 32785 2440
rect 32825 2420 32845 2630
rect 31985 2400 32375 2420
rect 32455 2400 32845 2420
rect 33095 2780 33455 2800
rect 33535 2780 33895 2800
rect 33095 2645 33115 2780
rect 33200 2750 33240 2760
rect 33200 2730 33210 2750
rect 33230 2730 33240 2750
rect 33200 2720 33240 2730
rect 33310 2750 33350 2760
rect 33310 2730 33320 2750
rect 33340 2730 33350 2750
rect 33310 2720 33350 2730
rect 33420 2750 33460 2760
rect 33420 2730 33430 2750
rect 33450 2730 33460 2750
rect 33420 2720 33460 2730
rect 33530 2750 33570 2760
rect 33530 2730 33540 2750
rect 33560 2730 33570 2750
rect 33530 2720 33570 2730
rect 33640 2750 33680 2760
rect 33640 2730 33650 2750
rect 33670 2730 33680 2750
rect 33640 2720 33680 2730
rect 33750 2750 33790 2760
rect 33750 2730 33760 2750
rect 33780 2730 33790 2750
rect 33750 2720 33790 2730
rect 33210 2700 33230 2720
rect 33320 2700 33340 2720
rect 33430 2700 33450 2720
rect 33540 2700 33560 2720
rect 33650 2700 33670 2720
rect 33760 2700 33780 2720
rect 33095 2430 33115 2565
rect 33150 2690 33180 2700
rect 33150 2670 33155 2690
rect 33175 2670 33180 2690
rect 33150 2640 33180 2670
rect 33150 2620 33155 2640
rect 33175 2620 33180 2640
rect 33150 2590 33180 2620
rect 33150 2570 33155 2590
rect 33175 2570 33180 2590
rect 33150 2540 33180 2570
rect 33150 2520 33155 2540
rect 33175 2520 33180 2540
rect 33150 2480 33180 2520
rect 33205 2690 33235 2700
rect 33205 2670 33210 2690
rect 33230 2670 33235 2690
rect 33205 2640 33235 2670
rect 33205 2620 33210 2640
rect 33230 2620 33235 2640
rect 33205 2590 33235 2620
rect 33205 2570 33210 2590
rect 33230 2570 33235 2590
rect 33205 2540 33235 2570
rect 33205 2520 33210 2540
rect 33230 2520 33235 2540
rect 33205 2510 33235 2520
rect 33260 2690 33290 2700
rect 33260 2670 33265 2690
rect 33285 2670 33290 2690
rect 33260 2640 33290 2670
rect 33260 2620 33265 2640
rect 33285 2620 33290 2640
rect 33260 2590 33290 2620
rect 33260 2570 33265 2590
rect 33285 2570 33290 2590
rect 33260 2540 33290 2570
rect 33260 2520 33265 2540
rect 33285 2520 33290 2540
rect 33260 2510 33290 2520
rect 33315 2690 33345 2700
rect 33315 2670 33320 2690
rect 33340 2670 33345 2690
rect 33315 2640 33345 2670
rect 33315 2620 33320 2640
rect 33340 2620 33345 2640
rect 33315 2590 33345 2620
rect 33315 2570 33320 2590
rect 33340 2570 33345 2590
rect 33315 2540 33345 2570
rect 33315 2520 33320 2540
rect 33340 2520 33345 2540
rect 33315 2510 33345 2520
rect 33370 2690 33400 2700
rect 33370 2670 33375 2690
rect 33395 2670 33400 2690
rect 33370 2640 33400 2670
rect 33370 2620 33375 2640
rect 33395 2620 33400 2640
rect 33370 2590 33400 2620
rect 33370 2570 33375 2590
rect 33395 2570 33400 2590
rect 33370 2540 33400 2570
rect 33370 2520 33375 2540
rect 33395 2520 33400 2540
rect 33370 2510 33400 2520
rect 33425 2690 33455 2700
rect 33425 2670 33430 2690
rect 33450 2670 33455 2690
rect 33425 2640 33455 2670
rect 33425 2620 33430 2640
rect 33450 2620 33455 2640
rect 33425 2590 33455 2620
rect 33425 2570 33430 2590
rect 33450 2570 33455 2590
rect 33425 2540 33455 2570
rect 33425 2520 33430 2540
rect 33450 2520 33455 2540
rect 33425 2510 33455 2520
rect 33480 2690 33510 2700
rect 33480 2670 33485 2690
rect 33505 2670 33510 2690
rect 33480 2640 33510 2670
rect 33480 2620 33485 2640
rect 33505 2620 33510 2640
rect 33480 2590 33510 2620
rect 33480 2570 33485 2590
rect 33505 2570 33510 2590
rect 33480 2540 33510 2570
rect 33480 2520 33485 2540
rect 33505 2520 33510 2540
rect 33480 2510 33510 2520
rect 33535 2690 33565 2700
rect 33535 2670 33540 2690
rect 33560 2670 33565 2690
rect 33535 2640 33565 2670
rect 33535 2620 33540 2640
rect 33560 2620 33565 2640
rect 33535 2590 33565 2620
rect 33535 2570 33540 2590
rect 33560 2570 33565 2590
rect 33535 2540 33565 2570
rect 33535 2520 33540 2540
rect 33560 2520 33565 2540
rect 33535 2510 33565 2520
rect 33590 2690 33620 2700
rect 33590 2670 33595 2690
rect 33615 2670 33620 2690
rect 33590 2640 33620 2670
rect 33590 2620 33595 2640
rect 33615 2620 33620 2640
rect 33590 2590 33620 2620
rect 33590 2570 33595 2590
rect 33615 2570 33620 2590
rect 33590 2540 33620 2570
rect 33590 2520 33595 2540
rect 33615 2520 33620 2540
rect 33590 2510 33620 2520
rect 33645 2690 33675 2700
rect 33645 2670 33650 2690
rect 33670 2670 33675 2690
rect 33645 2640 33675 2670
rect 33645 2620 33650 2640
rect 33670 2620 33675 2640
rect 33645 2590 33675 2620
rect 33645 2570 33650 2590
rect 33670 2570 33675 2590
rect 33645 2540 33675 2570
rect 33645 2520 33650 2540
rect 33670 2520 33675 2540
rect 33645 2510 33675 2520
rect 33700 2690 33730 2700
rect 33700 2670 33705 2690
rect 33725 2670 33730 2690
rect 33700 2640 33730 2670
rect 33700 2620 33705 2640
rect 33725 2620 33730 2640
rect 33700 2590 33730 2620
rect 33700 2570 33705 2590
rect 33725 2570 33730 2590
rect 33700 2540 33730 2570
rect 33700 2520 33705 2540
rect 33725 2520 33730 2540
rect 33700 2510 33730 2520
rect 33755 2690 33785 2700
rect 33755 2670 33760 2690
rect 33780 2670 33785 2690
rect 33755 2640 33785 2670
rect 33755 2620 33760 2640
rect 33780 2620 33785 2640
rect 33755 2590 33785 2620
rect 33755 2570 33760 2590
rect 33780 2570 33785 2590
rect 33755 2540 33785 2570
rect 33755 2520 33760 2540
rect 33780 2520 33785 2540
rect 33755 2510 33785 2520
rect 33810 2690 33840 2700
rect 33810 2670 33815 2690
rect 33835 2670 33840 2690
rect 33810 2640 33840 2670
rect 33810 2620 33815 2640
rect 33835 2620 33840 2640
rect 33810 2590 33840 2620
rect 33810 2570 33815 2590
rect 33835 2570 33840 2590
rect 33810 2540 33840 2570
rect 33810 2520 33815 2540
rect 33835 2520 33840 2540
rect 33265 2490 33285 2510
rect 33375 2490 33395 2510
rect 33485 2490 33505 2510
rect 33595 2490 33615 2510
rect 33705 2490 33725 2510
rect 33150 2460 33155 2480
rect 33175 2460 33180 2480
rect 33150 2450 33180 2460
rect 33255 2480 33295 2490
rect 33255 2460 33265 2480
rect 33285 2460 33295 2480
rect 33255 2450 33295 2460
rect 33313 2480 33347 2490
rect 33313 2460 33321 2480
rect 33339 2460 33347 2480
rect 33313 2450 33347 2460
rect 33365 2480 33405 2490
rect 33365 2460 33375 2480
rect 33395 2460 33405 2480
rect 33365 2450 33405 2460
rect 33475 2480 33515 2490
rect 33475 2460 33485 2480
rect 33505 2460 33515 2480
rect 33475 2450 33515 2460
rect 33585 2480 33625 2490
rect 33585 2460 33595 2480
rect 33615 2460 33625 2480
rect 33585 2450 33625 2460
rect 33695 2480 33735 2490
rect 33695 2460 33705 2480
rect 33725 2460 33735 2480
rect 33695 2450 33735 2460
rect 33810 2480 33840 2520
rect 33810 2460 33815 2480
rect 33835 2460 33840 2480
rect 33810 2450 33840 2460
rect 33875 2645 33895 2780
rect 34235 2679 34275 2689
rect 34235 2669 34245 2679
rect 34265 2669 34275 2679
rect 33155 2430 33175 2450
rect 33815 2430 33835 2450
rect 33875 2430 33895 2565
rect 33095 2410 33455 2430
rect 33535 2410 33895 2430
rect 34045 2649 34185 2669
rect 34265 2649 34400 2669
rect 29470 1980 29505 1990
rect 29470 1955 29475 1980
rect 29500 1955 29505 1980
rect 29470 1945 29505 1955
rect 29530 1980 29565 1990
rect 29530 1955 29535 1980
rect 29560 1955 29565 1980
rect 29530 1945 29565 1955
rect 29590 1980 29625 1990
rect 29590 1955 29595 1980
rect 29620 1955 29625 1980
rect 29590 1945 29625 1955
rect 29650 1980 29685 1990
rect 29650 1955 29655 1980
rect 29680 1955 29685 1980
rect 29650 1945 29685 1955
rect 29735 2115 29755 2255
rect 29905 2320 30265 2340
rect 30345 2320 30705 2340
rect 29905 2135 29925 2320
rect 29965 2300 29985 2320
rect 30625 2300 30645 2320
rect 29735 2105 29775 2115
rect 29735 2085 29745 2105
rect 29765 2085 29775 2105
rect 29735 2075 29775 2085
rect 29885 2105 29905 2115
rect 29885 2085 29895 2105
rect 29885 2075 29905 2085
rect 29735 1925 29755 2075
rect 29400 1905 29535 1925
rect 29615 1905 29755 1925
rect 29905 1870 29925 2055
rect 29960 2290 29990 2300
rect 29960 2270 29965 2290
rect 29985 2270 29990 2290
rect 29960 2230 29990 2270
rect 30065 2290 30105 2300
rect 30065 2270 30075 2290
rect 30095 2270 30105 2290
rect 30065 2260 30105 2270
rect 30175 2290 30215 2300
rect 30175 2270 30185 2290
rect 30205 2270 30215 2290
rect 30175 2260 30215 2270
rect 30285 2290 30325 2300
rect 30285 2270 30295 2290
rect 30315 2270 30325 2290
rect 30285 2260 30325 2270
rect 30395 2290 30435 2300
rect 30395 2270 30405 2290
rect 30425 2270 30435 2290
rect 30395 2260 30435 2270
rect 30453 2290 30487 2300
rect 30453 2270 30461 2290
rect 30479 2270 30487 2290
rect 30453 2260 30487 2270
rect 30505 2290 30545 2300
rect 30505 2270 30515 2290
rect 30535 2270 30545 2290
rect 30505 2260 30545 2270
rect 30620 2290 30650 2300
rect 30620 2270 30625 2290
rect 30645 2270 30650 2290
rect 30075 2240 30095 2260
rect 30185 2240 30205 2260
rect 30295 2240 30315 2260
rect 30405 2240 30425 2260
rect 30515 2240 30535 2260
rect 29960 2210 29965 2230
rect 29985 2210 29990 2230
rect 29960 2180 29990 2210
rect 29960 2160 29965 2180
rect 29985 2160 29990 2180
rect 29960 2130 29990 2160
rect 29960 2110 29965 2130
rect 29985 2110 29990 2130
rect 29960 2080 29990 2110
rect 29960 2060 29965 2080
rect 29985 2060 29990 2080
rect 29960 2030 29990 2060
rect 29960 2010 29965 2030
rect 29985 2010 29990 2030
rect 29960 1980 29990 2010
rect 29960 1960 29965 1980
rect 29985 1960 29990 1980
rect 29960 1950 29990 1960
rect 30015 2230 30045 2240
rect 30015 2210 30020 2230
rect 30040 2210 30045 2230
rect 30015 2180 30045 2210
rect 30015 2160 30020 2180
rect 30040 2160 30045 2180
rect 30015 2130 30045 2160
rect 30015 2110 30020 2130
rect 30040 2110 30045 2130
rect 30015 2080 30045 2110
rect 30015 2060 30020 2080
rect 30040 2060 30045 2080
rect 30015 2030 30045 2060
rect 30015 2010 30020 2030
rect 30040 2010 30045 2030
rect 30015 1980 30045 2010
rect 30015 1960 30020 1980
rect 30040 1960 30045 1980
rect 30015 1950 30045 1960
rect 30070 2230 30100 2240
rect 30070 2210 30075 2230
rect 30095 2210 30100 2230
rect 30070 2180 30100 2210
rect 30070 2160 30075 2180
rect 30095 2160 30100 2180
rect 30070 2130 30100 2160
rect 30070 2110 30075 2130
rect 30095 2110 30100 2130
rect 30070 2080 30100 2110
rect 30070 2060 30075 2080
rect 30095 2060 30100 2080
rect 30070 2030 30100 2060
rect 30070 2010 30075 2030
rect 30095 2010 30100 2030
rect 30070 1980 30100 2010
rect 30070 1960 30075 1980
rect 30095 1960 30100 1980
rect 30070 1950 30100 1960
rect 30125 2230 30155 2240
rect 30125 2210 30130 2230
rect 30150 2210 30155 2230
rect 30125 2180 30155 2210
rect 30125 2160 30130 2180
rect 30150 2160 30155 2180
rect 30125 2130 30155 2160
rect 30125 2110 30130 2130
rect 30150 2110 30155 2130
rect 30125 2080 30155 2110
rect 30125 2060 30130 2080
rect 30150 2060 30155 2080
rect 30125 2030 30155 2060
rect 30125 2010 30130 2030
rect 30150 2010 30155 2030
rect 30125 1980 30155 2010
rect 30125 1960 30130 1980
rect 30150 1960 30155 1980
rect 30125 1950 30155 1960
rect 30180 2230 30210 2240
rect 30180 2210 30185 2230
rect 30205 2210 30210 2230
rect 30180 2180 30210 2210
rect 30180 2160 30185 2180
rect 30205 2160 30210 2180
rect 30180 2130 30210 2160
rect 30180 2110 30185 2130
rect 30205 2110 30210 2130
rect 30180 2080 30210 2110
rect 30180 2060 30185 2080
rect 30205 2060 30210 2080
rect 30180 2030 30210 2060
rect 30180 2010 30185 2030
rect 30205 2010 30210 2030
rect 30180 1980 30210 2010
rect 30180 1960 30185 1980
rect 30205 1960 30210 1980
rect 30180 1950 30210 1960
rect 30235 2230 30265 2240
rect 30235 2210 30240 2230
rect 30260 2210 30265 2230
rect 30235 2180 30265 2210
rect 30235 2160 30240 2180
rect 30260 2160 30265 2180
rect 30235 2130 30265 2160
rect 30235 2110 30240 2130
rect 30260 2110 30265 2130
rect 30235 2080 30265 2110
rect 30235 2060 30240 2080
rect 30260 2060 30265 2080
rect 30235 2030 30265 2060
rect 30235 2010 30240 2030
rect 30260 2010 30265 2030
rect 30235 1980 30265 2010
rect 30235 1960 30240 1980
rect 30260 1960 30265 1980
rect 30235 1950 30265 1960
rect 30290 2230 30320 2240
rect 30290 2210 30295 2230
rect 30315 2210 30320 2230
rect 30290 2180 30320 2210
rect 30290 2160 30295 2180
rect 30315 2160 30320 2180
rect 30290 2130 30320 2160
rect 30290 2110 30295 2130
rect 30315 2110 30320 2130
rect 30290 2080 30320 2110
rect 30290 2060 30295 2080
rect 30315 2060 30320 2080
rect 30290 2030 30320 2060
rect 30290 2010 30295 2030
rect 30315 2010 30320 2030
rect 30290 1980 30320 2010
rect 30290 1960 30295 1980
rect 30315 1960 30320 1980
rect 30290 1950 30320 1960
rect 30345 2230 30375 2240
rect 30345 2210 30350 2230
rect 30370 2210 30375 2230
rect 30345 2180 30375 2210
rect 30345 2160 30350 2180
rect 30370 2160 30375 2180
rect 30345 2130 30375 2160
rect 30345 2110 30350 2130
rect 30370 2110 30375 2130
rect 30345 2080 30375 2110
rect 30345 2060 30350 2080
rect 30370 2060 30375 2080
rect 30345 2030 30375 2060
rect 30345 2010 30350 2030
rect 30370 2010 30375 2030
rect 30345 1980 30375 2010
rect 30345 1960 30350 1980
rect 30370 1960 30375 1980
rect 30345 1950 30375 1960
rect 30400 2230 30430 2240
rect 30400 2210 30405 2230
rect 30425 2210 30430 2230
rect 30400 2180 30430 2210
rect 30400 2160 30405 2180
rect 30425 2160 30430 2180
rect 30400 2130 30430 2160
rect 30400 2110 30405 2130
rect 30425 2110 30430 2130
rect 30400 2080 30430 2110
rect 30400 2060 30405 2080
rect 30425 2060 30430 2080
rect 30400 2030 30430 2060
rect 30400 2010 30405 2030
rect 30425 2010 30430 2030
rect 30400 1980 30430 2010
rect 30400 1960 30405 1980
rect 30425 1960 30430 1980
rect 30400 1950 30430 1960
rect 30455 2230 30485 2240
rect 30455 2210 30460 2230
rect 30480 2210 30485 2230
rect 30455 2180 30485 2210
rect 30455 2160 30460 2180
rect 30480 2160 30485 2180
rect 30455 2130 30485 2160
rect 30455 2110 30460 2130
rect 30480 2110 30485 2130
rect 30455 2080 30485 2110
rect 30455 2060 30460 2080
rect 30480 2060 30485 2080
rect 30455 2030 30485 2060
rect 30455 2010 30460 2030
rect 30480 2010 30485 2030
rect 30455 1980 30485 2010
rect 30455 1960 30460 1980
rect 30480 1960 30485 1980
rect 30455 1950 30485 1960
rect 30510 2230 30540 2240
rect 30510 2210 30515 2230
rect 30535 2210 30540 2230
rect 30510 2180 30540 2210
rect 30510 2160 30515 2180
rect 30535 2160 30540 2180
rect 30510 2130 30540 2160
rect 30510 2110 30515 2130
rect 30535 2110 30540 2130
rect 30510 2080 30540 2110
rect 30510 2060 30515 2080
rect 30535 2060 30540 2080
rect 30510 2030 30540 2060
rect 30510 2010 30515 2030
rect 30535 2010 30540 2030
rect 30510 1980 30540 2010
rect 30510 1960 30515 1980
rect 30535 1960 30540 1980
rect 30510 1950 30540 1960
rect 30565 2230 30595 2240
rect 30565 2210 30570 2230
rect 30590 2210 30595 2230
rect 30565 2180 30595 2210
rect 30565 2160 30570 2180
rect 30590 2160 30595 2180
rect 30565 2130 30595 2160
rect 30565 2110 30570 2130
rect 30590 2110 30595 2130
rect 30565 2080 30595 2110
rect 30565 2060 30570 2080
rect 30590 2060 30595 2080
rect 30565 2030 30595 2060
rect 30565 2010 30570 2030
rect 30590 2010 30595 2030
rect 30565 1980 30595 2010
rect 30565 1960 30570 1980
rect 30590 1960 30595 1980
rect 30565 1950 30595 1960
rect 30620 2230 30650 2270
rect 30620 2210 30625 2230
rect 30645 2210 30650 2230
rect 30620 2180 30650 2210
rect 30620 2160 30625 2180
rect 30645 2160 30650 2180
rect 30620 2130 30650 2160
rect 30620 2110 30625 2130
rect 30645 2110 30650 2130
rect 30620 2080 30650 2110
rect 30620 2060 30625 2080
rect 30645 2060 30650 2080
rect 30620 2030 30650 2060
rect 30620 2010 30625 2030
rect 30645 2010 30650 2030
rect 30620 1980 30650 2010
rect 30620 1960 30625 1980
rect 30645 1960 30650 1980
rect 30620 1950 30650 1960
rect 30685 2135 30705 2320
rect 33095 2320 33455 2340
rect 33535 2320 33895 2340
rect 30020 1930 30040 1950
rect 30130 1930 30150 1950
rect 30240 1930 30260 1950
rect 30350 1930 30370 1950
rect 30460 1930 30480 1950
rect 30570 1930 30590 1950
rect 30010 1920 30050 1930
rect 30010 1900 30020 1920
rect 30038 1900 30050 1920
rect 30010 1890 30050 1900
rect 30120 1920 30160 1930
rect 30120 1900 30130 1920
rect 30148 1900 30160 1920
rect 30120 1890 30160 1900
rect 30230 1920 30270 1930
rect 30230 1900 30240 1920
rect 30258 1900 30270 1920
rect 30230 1890 30270 1900
rect 30340 1920 30380 1930
rect 30340 1900 30350 1920
rect 30368 1900 30380 1920
rect 30340 1890 30380 1900
rect 30450 1920 30490 1930
rect 30450 1900 30460 1920
rect 30478 1900 30490 1920
rect 30450 1890 30490 1900
rect 30560 1920 30600 1930
rect 30560 1900 30570 1920
rect 30588 1900 30600 1920
rect 30560 1890 30600 1900
rect 30685 1870 30705 2055
rect 31095 2255 31860 2275
rect 31940 2255 32705 2275
rect 31095 2145 31115 2255
rect 31195 2235 31215 2255
rect 31855 2235 31875 2255
rect 31925 2235 31945 2255
rect 32585 2235 32605 2255
rect 31095 1955 31115 2065
rect 31190 2225 31220 2235
rect 31190 2205 31195 2225
rect 31215 2205 31220 2225
rect 31190 2165 31220 2205
rect 31240 2225 31280 2235
rect 31240 2205 31250 2225
rect 31270 2205 31280 2225
rect 31240 2195 31280 2205
rect 31350 2225 31390 2235
rect 31350 2205 31360 2225
rect 31380 2205 31390 2225
rect 31350 2195 31390 2205
rect 31460 2225 31500 2235
rect 31460 2205 31470 2225
rect 31490 2205 31500 2225
rect 31460 2195 31500 2205
rect 31520 2225 31550 2235
rect 31520 2205 31525 2225
rect 31545 2205 31550 2225
rect 31520 2195 31550 2205
rect 31570 2225 31610 2235
rect 31570 2205 31580 2225
rect 31600 2205 31610 2225
rect 31570 2195 31610 2205
rect 31680 2225 31720 2235
rect 31680 2205 31690 2225
rect 31710 2205 31720 2225
rect 31680 2195 31720 2205
rect 31790 2225 31830 2235
rect 31790 2205 31800 2225
rect 31820 2205 31830 2225
rect 31790 2195 31830 2205
rect 31850 2225 31880 2235
rect 31850 2205 31855 2225
rect 31875 2205 31880 2225
rect 31250 2175 31270 2195
rect 31360 2175 31380 2195
rect 31470 2175 31490 2195
rect 31580 2175 31600 2195
rect 31690 2175 31710 2195
rect 31800 2175 31820 2195
rect 31190 2145 31195 2165
rect 31215 2145 31220 2165
rect 31190 2115 31220 2145
rect 31190 2095 31195 2115
rect 31215 2095 31220 2115
rect 31190 2065 31220 2095
rect 31190 2045 31195 2065
rect 31215 2045 31220 2065
rect 31190 2035 31220 2045
rect 31245 2165 31275 2175
rect 31245 2145 31250 2165
rect 31270 2145 31275 2165
rect 31245 2115 31275 2145
rect 31245 2095 31250 2115
rect 31270 2095 31275 2115
rect 31245 2065 31275 2095
rect 31245 2045 31250 2065
rect 31270 2045 31275 2065
rect 31245 2035 31275 2045
rect 31300 2165 31330 2175
rect 31300 2145 31305 2165
rect 31325 2145 31330 2165
rect 31300 2115 31330 2145
rect 31300 2095 31305 2115
rect 31325 2095 31330 2115
rect 31300 2065 31330 2095
rect 31300 2045 31305 2065
rect 31325 2045 31330 2065
rect 31300 2035 31330 2045
rect 31355 2165 31385 2175
rect 31355 2145 31360 2165
rect 31380 2145 31385 2165
rect 31355 2115 31385 2145
rect 31355 2095 31360 2115
rect 31380 2095 31385 2115
rect 31355 2065 31385 2095
rect 31355 2045 31360 2065
rect 31380 2045 31385 2065
rect 31355 2035 31385 2045
rect 31410 2165 31440 2175
rect 31410 2145 31415 2165
rect 31435 2145 31440 2165
rect 31410 2115 31440 2145
rect 31410 2095 31415 2115
rect 31435 2095 31440 2115
rect 31410 2065 31440 2095
rect 31410 2045 31415 2065
rect 31435 2045 31440 2065
rect 31410 2035 31440 2045
rect 31465 2165 31495 2175
rect 31465 2145 31470 2165
rect 31490 2145 31495 2165
rect 31465 2115 31495 2145
rect 31465 2095 31470 2115
rect 31490 2095 31495 2115
rect 31465 2065 31495 2095
rect 31465 2045 31470 2065
rect 31490 2045 31495 2065
rect 31465 2035 31495 2045
rect 31520 2165 31550 2175
rect 31520 2145 31525 2165
rect 31545 2145 31550 2165
rect 31520 2115 31550 2145
rect 31520 2095 31525 2115
rect 31545 2095 31550 2115
rect 31520 2065 31550 2095
rect 31520 2045 31525 2065
rect 31545 2045 31550 2065
rect 31520 2035 31550 2045
rect 31575 2165 31605 2175
rect 31575 2145 31580 2165
rect 31600 2145 31605 2165
rect 31575 2115 31605 2145
rect 31575 2095 31580 2115
rect 31600 2095 31605 2115
rect 31575 2065 31605 2095
rect 31575 2045 31580 2065
rect 31600 2045 31605 2065
rect 31575 2035 31605 2045
rect 31630 2165 31660 2175
rect 31630 2145 31635 2165
rect 31655 2145 31660 2165
rect 31630 2115 31660 2145
rect 31630 2095 31635 2115
rect 31655 2095 31660 2115
rect 31630 2065 31660 2095
rect 31630 2045 31635 2065
rect 31655 2045 31660 2065
rect 31630 2035 31660 2045
rect 31685 2165 31715 2175
rect 31685 2145 31690 2165
rect 31710 2145 31715 2165
rect 31685 2115 31715 2145
rect 31685 2095 31690 2115
rect 31710 2095 31715 2115
rect 31685 2065 31715 2095
rect 31685 2045 31690 2065
rect 31710 2045 31715 2065
rect 31685 2035 31715 2045
rect 31740 2165 31770 2175
rect 31740 2145 31745 2165
rect 31765 2145 31770 2165
rect 31740 2115 31770 2145
rect 31740 2095 31745 2115
rect 31765 2095 31770 2115
rect 31740 2065 31770 2095
rect 31740 2045 31745 2065
rect 31765 2045 31770 2065
rect 31740 2035 31770 2045
rect 31795 2165 31825 2175
rect 31795 2145 31800 2165
rect 31820 2145 31825 2165
rect 31795 2115 31825 2145
rect 31795 2095 31800 2115
rect 31820 2095 31825 2115
rect 31795 2065 31825 2095
rect 31795 2045 31800 2065
rect 31820 2045 31825 2065
rect 31795 2035 31825 2045
rect 31850 2165 31880 2205
rect 31850 2145 31855 2165
rect 31875 2145 31880 2165
rect 31850 2115 31880 2145
rect 31850 2095 31855 2115
rect 31875 2095 31880 2115
rect 31850 2065 31880 2095
rect 31850 2045 31855 2065
rect 31875 2045 31880 2065
rect 31850 2035 31880 2045
rect 31920 2225 31950 2235
rect 31920 2205 31925 2225
rect 31945 2205 31950 2225
rect 31920 2165 31950 2205
rect 31970 2225 32010 2235
rect 31970 2205 31980 2225
rect 32000 2205 32010 2225
rect 31970 2195 32010 2205
rect 32080 2225 32120 2235
rect 32080 2205 32090 2225
rect 32110 2205 32120 2225
rect 32080 2195 32120 2205
rect 32190 2225 32230 2235
rect 32190 2205 32200 2225
rect 32220 2205 32230 2225
rect 32190 2195 32230 2205
rect 32250 2225 32280 2235
rect 32250 2205 32255 2225
rect 32275 2205 32280 2225
rect 32250 2195 32280 2205
rect 32300 2225 32340 2235
rect 32300 2205 32310 2225
rect 32330 2205 32340 2225
rect 32300 2195 32340 2205
rect 32410 2225 32450 2235
rect 32410 2205 32420 2225
rect 32440 2205 32450 2225
rect 32410 2195 32450 2205
rect 32520 2225 32560 2235
rect 32520 2205 32530 2225
rect 32550 2205 32560 2225
rect 32520 2195 32560 2205
rect 32580 2225 32610 2235
rect 32580 2205 32585 2225
rect 32605 2205 32610 2225
rect 31980 2175 32000 2195
rect 32090 2175 32110 2195
rect 32200 2175 32220 2195
rect 32310 2175 32330 2195
rect 32420 2175 32440 2195
rect 32530 2175 32550 2195
rect 31920 2145 31925 2165
rect 31945 2145 31950 2165
rect 31920 2115 31950 2145
rect 31920 2095 31925 2115
rect 31945 2095 31950 2115
rect 31920 2065 31950 2095
rect 31920 2045 31925 2065
rect 31945 2045 31950 2065
rect 31920 2035 31950 2045
rect 31975 2165 32005 2175
rect 31975 2145 31980 2165
rect 32000 2145 32005 2165
rect 31975 2115 32005 2145
rect 31975 2095 31980 2115
rect 32000 2095 32005 2115
rect 31975 2065 32005 2095
rect 31975 2045 31980 2065
rect 32000 2045 32005 2065
rect 31975 2035 32005 2045
rect 32030 2165 32060 2175
rect 32030 2145 32035 2165
rect 32055 2145 32060 2165
rect 32030 2115 32060 2145
rect 32030 2095 32035 2115
rect 32055 2095 32060 2115
rect 32030 2065 32060 2095
rect 32030 2045 32035 2065
rect 32055 2045 32060 2065
rect 32030 2035 32060 2045
rect 32085 2165 32115 2175
rect 32085 2145 32090 2165
rect 32110 2145 32115 2165
rect 32085 2115 32115 2145
rect 32085 2095 32090 2115
rect 32110 2095 32115 2115
rect 32085 2065 32115 2095
rect 32085 2045 32090 2065
rect 32110 2045 32115 2065
rect 32085 2035 32115 2045
rect 32140 2165 32170 2175
rect 32140 2145 32145 2165
rect 32165 2145 32170 2165
rect 32140 2115 32170 2145
rect 32140 2095 32145 2115
rect 32165 2095 32170 2115
rect 32140 2065 32170 2095
rect 32140 2045 32145 2065
rect 32165 2045 32170 2065
rect 32140 2035 32170 2045
rect 32195 2165 32225 2175
rect 32195 2145 32200 2165
rect 32220 2145 32225 2165
rect 32195 2115 32225 2145
rect 32195 2095 32200 2115
rect 32220 2095 32225 2115
rect 32195 2065 32225 2095
rect 32195 2045 32200 2065
rect 32220 2045 32225 2065
rect 32195 2035 32225 2045
rect 32250 2165 32280 2175
rect 32250 2145 32255 2165
rect 32275 2145 32280 2165
rect 32250 2115 32280 2145
rect 32250 2095 32255 2115
rect 32275 2095 32280 2115
rect 32250 2065 32280 2095
rect 32250 2045 32255 2065
rect 32275 2045 32280 2065
rect 32250 2035 32280 2045
rect 32305 2165 32335 2175
rect 32305 2145 32310 2165
rect 32330 2145 32335 2165
rect 32305 2115 32335 2145
rect 32305 2095 32310 2115
rect 32330 2095 32335 2115
rect 32305 2065 32335 2095
rect 32305 2045 32310 2065
rect 32330 2045 32335 2065
rect 32305 2035 32335 2045
rect 32360 2165 32390 2175
rect 32360 2145 32365 2165
rect 32385 2145 32390 2165
rect 32360 2115 32390 2145
rect 32360 2095 32365 2115
rect 32385 2095 32390 2115
rect 32360 2065 32390 2095
rect 32360 2045 32365 2065
rect 32385 2045 32390 2065
rect 32360 2035 32390 2045
rect 32415 2165 32445 2175
rect 32415 2145 32420 2165
rect 32440 2145 32445 2165
rect 32415 2115 32445 2145
rect 32415 2095 32420 2115
rect 32440 2095 32445 2115
rect 32415 2065 32445 2095
rect 32415 2045 32420 2065
rect 32440 2045 32445 2065
rect 32415 2035 32445 2045
rect 32470 2165 32500 2175
rect 32470 2145 32475 2165
rect 32495 2145 32500 2165
rect 32470 2115 32500 2145
rect 32470 2095 32475 2115
rect 32495 2095 32500 2115
rect 32470 2065 32500 2095
rect 32470 2045 32475 2065
rect 32495 2045 32500 2065
rect 32470 2035 32500 2045
rect 32525 2165 32555 2175
rect 32525 2145 32530 2165
rect 32550 2145 32555 2165
rect 32525 2115 32555 2145
rect 32525 2095 32530 2115
rect 32550 2095 32555 2115
rect 32525 2065 32555 2095
rect 32525 2045 32530 2065
rect 32550 2045 32555 2065
rect 32525 2035 32555 2045
rect 32580 2165 32610 2205
rect 32580 2145 32585 2165
rect 32605 2145 32610 2165
rect 32580 2115 32610 2145
rect 32580 2095 32585 2115
rect 32605 2095 32610 2115
rect 32580 2065 32610 2095
rect 32580 2045 32585 2065
rect 32605 2045 32610 2065
rect 32580 2035 32610 2045
rect 32685 2145 32705 2255
rect 31305 2015 31325 2035
rect 31415 2015 31435 2035
rect 31525 2015 31545 2035
rect 31635 2015 31655 2035
rect 31745 2015 31765 2035
rect 32035 2015 32055 2035
rect 32145 2015 32165 2035
rect 32255 2015 32275 2035
rect 32365 2015 32385 2035
rect 32475 2015 32495 2035
rect 31295 2005 31335 2015
rect 31295 1985 31305 2005
rect 31325 1985 31335 2005
rect 31295 1975 31335 1985
rect 31405 2005 31445 2015
rect 31405 1985 31415 2005
rect 31435 1985 31445 2005
rect 31405 1975 31445 1985
rect 31515 2005 31555 2015
rect 31515 1985 31525 2005
rect 31545 1985 31555 2005
rect 31515 1975 31555 1985
rect 31625 2005 31665 2015
rect 31625 1985 31635 2005
rect 31655 1985 31665 2005
rect 31625 1975 31665 1985
rect 31735 2005 31775 2015
rect 31735 1985 31745 2005
rect 31765 1985 31775 2005
rect 31735 1975 31775 1985
rect 32025 2005 32065 2015
rect 32025 1985 32035 2005
rect 32055 1985 32065 2005
rect 32025 1975 32065 1985
rect 32135 2005 32175 2015
rect 32135 1985 32145 2005
rect 32165 1985 32175 2005
rect 32135 1975 32175 1985
rect 32245 2005 32285 2015
rect 32245 1985 32255 2005
rect 32275 1985 32285 2005
rect 32245 1975 32285 1985
rect 32355 2005 32395 2015
rect 32355 1985 32365 2005
rect 32385 1985 32395 2005
rect 32355 1975 32395 1985
rect 32465 2005 32505 2015
rect 32465 1985 32475 2005
rect 32495 1985 32505 2005
rect 32465 1975 32505 1985
rect 32685 1955 32705 2065
rect 31095 1935 31860 1955
rect 31940 1935 32705 1955
rect 33095 2135 33115 2320
rect 33155 2300 33175 2320
rect 33815 2300 33835 2320
rect 31880 1925 31890 1935
rect 31910 1925 31920 1935
rect 31880 1915 31920 1925
rect 29905 1850 30265 1870
rect 30345 1850 30705 1870
rect 33095 1870 33115 2055
rect 33150 2290 33180 2300
rect 33150 2270 33155 2290
rect 33175 2270 33180 2290
rect 33150 2230 33180 2270
rect 33255 2290 33295 2300
rect 33255 2270 33265 2290
rect 33285 2270 33295 2290
rect 33255 2260 33295 2270
rect 33313 2290 33347 2300
rect 33313 2270 33321 2290
rect 33339 2270 33347 2290
rect 33313 2260 33347 2270
rect 33365 2290 33405 2300
rect 33365 2270 33375 2290
rect 33395 2270 33405 2290
rect 33365 2260 33405 2270
rect 33475 2290 33515 2300
rect 33475 2270 33485 2290
rect 33505 2270 33515 2290
rect 33475 2260 33515 2270
rect 33585 2290 33625 2300
rect 33585 2270 33595 2290
rect 33615 2270 33625 2290
rect 33585 2260 33625 2270
rect 33695 2290 33735 2300
rect 33695 2270 33705 2290
rect 33725 2270 33735 2290
rect 33695 2260 33735 2270
rect 33810 2290 33840 2300
rect 33810 2270 33815 2290
rect 33835 2270 33840 2290
rect 33265 2240 33285 2260
rect 33375 2240 33395 2260
rect 33485 2240 33505 2260
rect 33595 2240 33615 2260
rect 33705 2240 33725 2260
rect 33150 2210 33155 2230
rect 33175 2210 33180 2230
rect 33150 2180 33180 2210
rect 33150 2160 33155 2180
rect 33175 2160 33180 2180
rect 33150 2130 33180 2160
rect 33150 2110 33155 2130
rect 33175 2110 33180 2130
rect 33150 2080 33180 2110
rect 33150 2060 33155 2080
rect 33175 2060 33180 2080
rect 33150 2030 33180 2060
rect 33150 2010 33155 2030
rect 33175 2010 33180 2030
rect 33150 1980 33180 2010
rect 33150 1960 33155 1980
rect 33175 1960 33180 1980
rect 33150 1950 33180 1960
rect 33205 2230 33235 2240
rect 33205 2210 33210 2230
rect 33230 2210 33235 2230
rect 33205 2180 33235 2210
rect 33205 2160 33210 2180
rect 33230 2160 33235 2180
rect 33205 2130 33235 2160
rect 33205 2110 33210 2130
rect 33230 2110 33235 2130
rect 33205 2080 33235 2110
rect 33205 2060 33210 2080
rect 33230 2060 33235 2080
rect 33205 2030 33235 2060
rect 33205 2010 33210 2030
rect 33230 2010 33235 2030
rect 33205 1980 33235 2010
rect 33205 1960 33210 1980
rect 33230 1960 33235 1980
rect 33205 1950 33235 1960
rect 33260 2230 33290 2240
rect 33260 2210 33265 2230
rect 33285 2210 33290 2230
rect 33260 2180 33290 2210
rect 33260 2160 33265 2180
rect 33285 2160 33290 2180
rect 33260 2130 33290 2160
rect 33260 2110 33265 2130
rect 33285 2110 33290 2130
rect 33260 2080 33290 2110
rect 33260 2060 33265 2080
rect 33285 2060 33290 2080
rect 33260 2030 33290 2060
rect 33260 2010 33265 2030
rect 33285 2010 33290 2030
rect 33260 1980 33290 2010
rect 33260 1960 33265 1980
rect 33285 1960 33290 1980
rect 33260 1950 33290 1960
rect 33315 2230 33345 2240
rect 33315 2210 33320 2230
rect 33340 2210 33345 2230
rect 33315 2180 33345 2210
rect 33315 2160 33320 2180
rect 33340 2160 33345 2180
rect 33315 2130 33345 2160
rect 33315 2110 33320 2130
rect 33340 2110 33345 2130
rect 33315 2080 33345 2110
rect 33315 2060 33320 2080
rect 33340 2060 33345 2080
rect 33315 2030 33345 2060
rect 33315 2010 33320 2030
rect 33340 2010 33345 2030
rect 33315 1980 33345 2010
rect 33315 1960 33320 1980
rect 33340 1960 33345 1980
rect 33315 1950 33345 1960
rect 33370 2230 33400 2240
rect 33370 2210 33375 2230
rect 33395 2210 33400 2230
rect 33370 2180 33400 2210
rect 33370 2160 33375 2180
rect 33395 2160 33400 2180
rect 33370 2130 33400 2160
rect 33370 2110 33375 2130
rect 33395 2110 33400 2130
rect 33370 2080 33400 2110
rect 33370 2060 33375 2080
rect 33395 2060 33400 2080
rect 33370 2030 33400 2060
rect 33370 2010 33375 2030
rect 33395 2010 33400 2030
rect 33370 1980 33400 2010
rect 33370 1960 33375 1980
rect 33395 1960 33400 1980
rect 33370 1950 33400 1960
rect 33425 2230 33455 2240
rect 33425 2210 33430 2230
rect 33450 2210 33455 2230
rect 33425 2180 33455 2210
rect 33425 2160 33430 2180
rect 33450 2160 33455 2180
rect 33425 2130 33455 2160
rect 33425 2110 33430 2130
rect 33450 2110 33455 2130
rect 33425 2080 33455 2110
rect 33425 2060 33430 2080
rect 33450 2060 33455 2080
rect 33425 2030 33455 2060
rect 33425 2010 33430 2030
rect 33450 2010 33455 2030
rect 33425 1980 33455 2010
rect 33425 1960 33430 1980
rect 33450 1960 33455 1980
rect 33425 1950 33455 1960
rect 33480 2230 33510 2240
rect 33480 2210 33485 2230
rect 33505 2210 33510 2230
rect 33480 2180 33510 2210
rect 33480 2160 33485 2180
rect 33505 2160 33510 2180
rect 33480 2130 33510 2160
rect 33480 2110 33485 2130
rect 33505 2110 33510 2130
rect 33480 2080 33510 2110
rect 33480 2060 33485 2080
rect 33505 2060 33510 2080
rect 33480 2030 33510 2060
rect 33480 2010 33485 2030
rect 33505 2010 33510 2030
rect 33480 1980 33510 2010
rect 33480 1960 33485 1980
rect 33505 1960 33510 1980
rect 33480 1950 33510 1960
rect 33535 2230 33565 2240
rect 33535 2210 33540 2230
rect 33560 2210 33565 2230
rect 33535 2180 33565 2210
rect 33535 2160 33540 2180
rect 33560 2160 33565 2180
rect 33535 2130 33565 2160
rect 33535 2110 33540 2130
rect 33560 2110 33565 2130
rect 33535 2080 33565 2110
rect 33535 2060 33540 2080
rect 33560 2060 33565 2080
rect 33535 2030 33565 2060
rect 33535 2010 33540 2030
rect 33560 2010 33565 2030
rect 33535 1980 33565 2010
rect 33535 1960 33540 1980
rect 33560 1960 33565 1980
rect 33535 1950 33565 1960
rect 33590 2230 33620 2240
rect 33590 2210 33595 2230
rect 33615 2210 33620 2230
rect 33590 2180 33620 2210
rect 33590 2160 33595 2180
rect 33615 2160 33620 2180
rect 33590 2130 33620 2160
rect 33590 2110 33595 2130
rect 33615 2110 33620 2130
rect 33590 2080 33620 2110
rect 33590 2060 33595 2080
rect 33615 2060 33620 2080
rect 33590 2030 33620 2060
rect 33590 2010 33595 2030
rect 33615 2010 33620 2030
rect 33590 1980 33620 2010
rect 33590 1960 33595 1980
rect 33615 1960 33620 1980
rect 33590 1950 33620 1960
rect 33645 2230 33675 2240
rect 33645 2210 33650 2230
rect 33670 2210 33675 2230
rect 33645 2180 33675 2210
rect 33645 2160 33650 2180
rect 33670 2160 33675 2180
rect 33645 2130 33675 2160
rect 33645 2110 33650 2130
rect 33670 2110 33675 2130
rect 33645 2080 33675 2110
rect 33645 2060 33650 2080
rect 33670 2060 33675 2080
rect 33645 2030 33675 2060
rect 33645 2010 33650 2030
rect 33670 2010 33675 2030
rect 33645 1980 33675 2010
rect 33645 1960 33650 1980
rect 33670 1960 33675 1980
rect 33645 1950 33675 1960
rect 33700 2230 33730 2240
rect 33700 2210 33705 2230
rect 33725 2210 33730 2230
rect 33700 2180 33730 2210
rect 33700 2160 33705 2180
rect 33725 2160 33730 2180
rect 33700 2130 33730 2160
rect 33700 2110 33705 2130
rect 33725 2110 33730 2130
rect 33700 2080 33730 2110
rect 33700 2060 33705 2080
rect 33725 2060 33730 2080
rect 33700 2030 33730 2060
rect 33700 2010 33705 2030
rect 33725 2010 33730 2030
rect 33700 1980 33730 2010
rect 33700 1960 33705 1980
rect 33725 1960 33730 1980
rect 33700 1950 33730 1960
rect 33755 2230 33785 2240
rect 33755 2210 33760 2230
rect 33780 2210 33785 2230
rect 33755 2180 33785 2210
rect 33755 2160 33760 2180
rect 33780 2160 33785 2180
rect 33755 2130 33785 2160
rect 33755 2110 33760 2130
rect 33780 2110 33785 2130
rect 33755 2080 33785 2110
rect 33755 2060 33760 2080
rect 33780 2060 33785 2080
rect 33755 2030 33785 2060
rect 33755 2010 33760 2030
rect 33780 2010 33785 2030
rect 33755 1980 33785 2010
rect 33755 1960 33760 1980
rect 33780 1960 33785 1980
rect 33755 1950 33785 1960
rect 33810 2230 33840 2270
rect 33810 2210 33815 2230
rect 33835 2210 33840 2230
rect 33810 2180 33840 2210
rect 33810 2160 33815 2180
rect 33835 2160 33840 2180
rect 33810 2130 33840 2160
rect 33810 2110 33815 2130
rect 33835 2110 33840 2130
rect 33810 2080 33840 2110
rect 33810 2060 33815 2080
rect 33835 2060 33840 2080
rect 33810 2030 33840 2060
rect 33810 2010 33815 2030
rect 33835 2010 33840 2030
rect 33810 1980 33840 2010
rect 33810 1960 33815 1980
rect 33835 1960 33840 1980
rect 33810 1950 33840 1960
rect 33875 2135 33895 2320
rect 34045 2335 34065 2649
rect 34115 2609 34330 2629
rect 34115 2589 34150 2609
rect 34295 2589 34330 2609
rect 34210 2539 34235 2589
rect 34045 2115 34065 2255
rect 34380 2335 34400 2649
rect 33895 2105 33915 2115
rect 33905 2085 33915 2105
rect 33895 2075 33915 2085
rect 34025 2105 34065 2115
rect 34025 2085 34035 2105
rect 34055 2085 34065 2105
rect 34025 2075 34065 2085
rect 33210 1930 33230 1950
rect 33320 1930 33340 1950
rect 33430 1930 33450 1950
rect 33540 1930 33560 1950
rect 33650 1930 33670 1950
rect 33760 1930 33780 1950
rect 33200 1920 33240 1930
rect 33200 1900 33212 1920
rect 33230 1900 33240 1920
rect 33200 1890 33240 1900
rect 33310 1920 33350 1930
rect 33310 1900 33322 1920
rect 33340 1900 33350 1920
rect 33310 1890 33350 1900
rect 33420 1920 33460 1930
rect 33420 1900 33432 1920
rect 33450 1900 33460 1920
rect 33420 1890 33460 1900
rect 33530 1920 33570 1930
rect 33530 1900 33542 1920
rect 33560 1900 33570 1920
rect 33530 1890 33570 1900
rect 33640 1920 33680 1930
rect 33640 1900 33652 1920
rect 33670 1900 33680 1920
rect 33640 1890 33680 1900
rect 33750 1920 33790 1930
rect 33750 1900 33762 1920
rect 33780 1900 33790 1920
rect 33750 1890 33790 1900
rect 33875 1870 33895 2055
rect 34045 1925 34065 2075
rect 34115 1980 34150 1990
rect 34115 1955 34120 1980
rect 34145 1955 34150 1980
rect 34115 1945 34150 1955
rect 34175 1980 34210 1990
rect 34175 1955 34180 1980
rect 34205 1955 34210 1980
rect 34175 1945 34210 1955
rect 34235 1980 34270 1990
rect 34235 1955 34240 1980
rect 34265 1955 34270 1980
rect 34235 1945 34270 1955
rect 34295 1980 34330 1990
rect 34295 1955 34300 1980
rect 34325 1955 34330 1980
rect 34295 1945 34330 1955
rect 34380 1925 34400 2255
rect 34045 1905 34185 1925
rect 34265 1905 34400 1925
rect 33095 1850 33455 1870
rect 33535 1850 33895 1870
rect 30285 1840 30295 1850
rect 30315 1840 30325 1850
rect 30285 1830 30325 1840
rect 33475 1840 33485 1850
rect 33505 1840 33515 1850
rect 33475 1830 33515 1840
rect 31880 1815 31920 1825
rect 31880 1805 31890 1815
rect 31910 1805 31920 1815
rect 30940 1785 31860 1805
rect 31940 1785 32860 1805
rect 30285 1760 30325 1770
rect 30285 1750 30295 1760
rect 29985 1740 30295 1750
rect 30315 1750 30325 1760
rect 29985 1730 30315 1740
rect 30395 1730 30725 1750
rect 29660 1675 29735 1695
rect 29815 1675 29895 1695
rect 29660 1300 29680 1675
rect 29730 1640 29765 1650
rect 29730 1615 29735 1640
rect 29760 1615 29765 1640
rect 29730 1605 29765 1615
rect 29790 1640 29825 1650
rect 29790 1615 29795 1640
rect 29820 1615 29825 1640
rect 29790 1605 29825 1615
rect 29660 868 29680 1220
rect 29875 1325 29895 1675
rect 29985 1345 30005 1730
rect 30045 1710 30065 1730
rect 30645 1710 30665 1730
rect 29875 1315 29915 1325
rect 29875 1300 29885 1315
rect 29905 1295 29915 1315
rect 29895 1285 29915 1295
rect 29965 1315 29985 1325
rect 29965 1295 29975 1315
rect 29965 1285 29985 1295
rect 29765 918 29790 968
rect 29875 868 29895 1220
rect 29660 848 29735 868
rect 29815 848 29895 868
rect 29985 880 30005 1265
rect 30040 1700 30070 1710
rect 30040 1680 30045 1700
rect 30065 1680 30070 1700
rect 30040 1640 30070 1680
rect 30135 1700 30175 1710
rect 30135 1680 30145 1700
rect 30165 1680 30175 1700
rect 30135 1670 30175 1680
rect 30335 1700 30375 1710
rect 30335 1680 30345 1700
rect 30365 1680 30375 1700
rect 30335 1670 30375 1680
rect 30438 1700 30472 1710
rect 30438 1680 30446 1700
rect 30464 1680 30472 1700
rect 30438 1670 30472 1680
rect 30535 1700 30575 1710
rect 30535 1680 30545 1700
rect 30565 1680 30575 1700
rect 30535 1670 30575 1680
rect 30640 1700 30670 1710
rect 30640 1680 30645 1700
rect 30665 1680 30670 1700
rect 30145 1650 30165 1670
rect 30345 1650 30365 1670
rect 30545 1650 30565 1670
rect 30040 1620 30045 1640
rect 30065 1620 30070 1640
rect 30040 1590 30070 1620
rect 30040 1570 30045 1590
rect 30065 1570 30070 1590
rect 30040 1540 30070 1570
rect 30040 1520 30045 1540
rect 30065 1520 30070 1540
rect 30040 1490 30070 1520
rect 30040 1470 30045 1490
rect 30065 1470 30070 1490
rect 30040 1440 30070 1470
rect 30040 1420 30045 1440
rect 30065 1420 30070 1440
rect 30040 1390 30070 1420
rect 30040 1370 30045 1390
rect 30065 1370 30070 1390
rect 30040 1340 30070 1370
rect 30040 1320 30045 1340
rect 30065 1320 30070 1340
rect 30040 1290 30070 1320
rect 30040 1270 30045 1290
rect 30065 1270 30070 1290
rect 30040 1240 30070 1270
rect 30040 1220 30045 1240
rect 30065 1220 30070 1240
rect 30040 1190 30070 1220
rect 30040 1170 30045 1190
rect 30065 1170 30070 1190
rect 30040 1140 30070 1170
rect 30040 1120 30045 1140
rect 30065 1120 30070 1140
rect 30040 1090 30070 1120
rect 30040 1070 30045 1090
rect 30065 1070 30070 1090
rect 30040 1040 30070 1070
rect 30040 1020 30045 1040
rect 30065 1020 30070 1040
rect 30040 990 30070 1020
rect 30040 970 30045 990
rect 30065 970 30070 990
rect 30040 960 30070 970
rect 30140 1640 30170 1650
rect 30140 1620 30145 1640
rect 30165 1620 30170 1640
rect 30140 1590 30170 1620
rect 30140 1570 30145 1590
rect 30165 1570 30170 1590
rect 30140 1540 30170 1570
rect 30140 1520 30145 1540
rect 30165 1520 30170 1540
rect 30140 1490 30170 1520
rect 30140 1470 30145 1490
rect 30165 1470 30170 1490
rect 30140 1440 30170 1470
rect 30140 1420 30145 1440
rect 30165 1420 30170 1440
rect 30140 1390 30170 1420
rect 30140 1370 30145 1390
rect 30165 1370 30170 1390
rect 30140 1340 30170 1370
rect 30140 1320 30145 1340
rect 30165 1320 30170 1340
rect 30140 1290 30170 1320
rect 30140 1270 30145 1290
rect 30165 1270 30170 1290
rect 30140 1240 30170 1270
rect 30140 1220 30145 1240
rect 30165 1220 30170 1240
rect 30140 1190 30170 1220
rect 30140 1170 30145 1190
rect 30165 1170 30170 1190
rect 30140 1140 30170 1170
rect 30140 1120 30145 1140
rect 30165 1120 30170 1140
rect 30140 1090 30170 1120
rect 30140 1070 30145 1090
rect 30165 1070 30170 1090
rect 30140 1040 30170 1070
rect 30140 1020 30145 1040
rect 30165 1020 30170 1040
rect 30140 990 30170 1020
rect 30140 970 30145 990
rect 30165 970 30170 990
rect 30140 960 30170 970
rect 30240 1640 30270 1650
rect 30240 1620 30245 1640
rect 30265 1620 30270 1640
rect 30240 1590 30270 1620
rect 30240 1570 30245 1590
rect 30265 1570 30270 1590
rect 30240 1540 30270 1570
rect 30240 1520 30245 1540
rect 30265 1520 30270 1540
rect 30240 1490 30270 1520
rect 30240 1470 30245 1490
rect 30265 1470 30270 1490
rect 30240 1440 30270 1470
rect 30240 1420 30245 1440
rect 30265 1420 30270 1440
rect 30240 1390 30270 1420
rect 30240 1370 30245 1390
rect 30265 1370 30270 1390
rect 30240 1340 30270 1370
rect 30240 1320 30245 1340
rect 30265 1320 30270 1340
rect 30240 1290 30270 1320
rect 30240 1270 30245 1290
rect 30265 1270 30270 1290
rect 30240 1240 30270 1270
rect 30240 1220 30245 1240
rect 30265 1220 30270 1240
rect 30240 1190 30270 1220
rect 30240 1170 30245 1190
rect 30265 1170 30270 1190
rect 30240 1140 30270 1170
rect 30240 1120 30245 1140
rect 30265 1120 30270 1140
rect 30240 1090 30270 1120
rect 30240 1070 30245 1090
rect 30265 1070 30270 1090
rect 30240 1040 30270 1070
rect 30240 1020 30245 1040
rect 30265 1020 30270 1040
rect 30240 990 30270 1020
rect 30240 970 30245 990
rect 30265 970 30270 990
rect 30240 960 30270 970
rect 30340 1640 30370 1650
rect 30340 1620 30345 1640
rect 30365 1620 30370 1640
rect 30340 1590 30370 1620
rect 30340 1570 30345 1590
rect 30365 1570 30370 1590
rect 30340 1540 30370 1570
rect 30340 1520 30345 1540
rect 30365 1520 30370 1540
rect 30340 1490 30370 1520
rect 30340 1470 30345 1490
rect 30365 1470 30370 1490
rect 30340 1440 30370 1470
rect 30340 1420 30345 1440
rect 30365 1420 30370 1440
rect 30340 1390 30370 1420
rect 30340 1370 30345 1390
rect 30365 1370 30370 1390
rect 30340 1340 30370 1370
rect 30340 1320 30345 1340
rect 30365 1320 30370 1340
rect 30340 1290 30370 1320
rect 30340 1270 30345 1290
rect 30365 1270 30370 1290
rect 30340 1240 30370 1270
rect 30340 1220 30345 1240
rect 30365 1220 30370 1240
rect 30340 1190 30370 1220
rect 30340 1170 30345 1190
rect 30365 1170 30370 1190
rect 30340 1140 30370 1170
rect 30340 1120 30345 1140
rect 30365 1120 30370 1140
rect 30340 1090 30370 1120
rect 30340 1070 30345 1090
rect 30365 1070 30370 1090
rect 30340 1040 30370 1070
rect 30340 1020 30345 1040
rect 30365 1020 30370 1040
rect 30340 990 30370 1020
rect 30340 970 30345 990
rect 30365 970 30370 990
rect 30340 960 30370 970
rect 30440 1640 30470 1650
rect 30440 1620 30445 1640
rect 30465 1620 30470 1640
rect 30440 1590 30470 1620
rect 30440 1570 30445 1590
rect 30465 1570 30470 1590
rect 30440 1540 30470 1570
rect 30440 1520 30445 1540
rect 30465 1520 30470 1540
rect 30440 1490 30470 1520
rect 30440 1470 30445 1490
rect 30465 1470 30470 1490
rect 30440 1440 30470 1470
rect 30440 1420 30445 1440
rect 30465 1420 30470 1440
rect 30440 1390 30470 1420
rect 30440 1370 30445 1390
rect 30465 1370 30470 1390
rect 30440 1340 30470 1370
rect 30440 1320 30445 1340
rect 30465 1320 30470 1340
rect 30440 1290 30470 1320
rect 30440 1270 30445 1290
rect 30465 1270 30470 1290
rect 30440 1240 30470 1270
rect 30440 1220 30445 1240
rect 30465 1220 30470 1240
rect 30440 1190 30470 1220
rect 30440 1170 30445 1190
rect 30465 1170 30470 1190
rect 30440 1140 30470 1170
rect 30440 1120 30445 1140
rect 30465 1120 30470 1140
rect 30440 1090 30470 1120
rect 30440 1070 30445 1090
rect 30465 1070 30470 1090
rect 30440 1040 30470 1070
rect 30440 1020 30445 1040
rect 30465 1020 30470 1040
rect 30440 990 30470 1020
rect 30440 970 30445 990
rect 30465 970 30470 990
rect 30440 960 30470 970
rect 30540 1640 30570 1650
rect 30540 1620 30545 1640
rect 30565 1620 30570 1640
rect 30540 1590 30570 1620
rect 30540 1570 30545 1590
rect 30565 1570 30570 1590
rect 30540 1540 30570 1570
rect 30540 1520 30545 1540
rect 30565 1520 30570 1540
rect 30540 1490 30570 1520
rect 30540 1470 30545 1490
rect 30565 1470 30570 1490
rect 30540 1440 30570 1470
rect 30540 1420 30545 1440
rect 30565 1420 30570 1440
rect 30540 1390 30570 1420
rect 30540 1370 30545 1390
rect 30565 1370 30570 1390
rect 30540 1340 30570 1370
rect 30540 1320 30545 1340
rect 30565 1320 30570 1340
rect 30540 1290 30570 1320
rect 30540 1270 30545 1290
rect 30565 1270 30570 1290
rect 30540 1240 30570 1270
rect 30540 1220 30545 1240
rect 30565 1220 30570 1240
rect 30540 1190 30570 1220
rect 30540 1170 30545 1190
rect 30565 1170 30570 1190
rect 30540 1140 30570 1170
rect 30540 1120 30545 1140
rect 30565 1120 30570 1140
rect 30540 1090 30570 1120
rect 30540 1070 30545 1090
rect 30565 1070 30570 1090
rect 30540 1040 30570 1070
rect 30540 1020 30545 1040
rect 30565 1020 30570 1040
rect 30540 990 30570 1020
rect 30540 970 30545 990
rect 30565 970 30570 990
rect 30540 960 30570 970
rect 30640 1640 30670 1680
rect 30640 1620 30645 1640
rect 30665 1620 30670 1640
rect 30640 1590 30670 1620
rect 30640 1570 30645 1590
rect 30665 1570 30670 1590
rect 30640 1540 30670 1570
rect 30640 1520 30645 1540
rect 30665 1520 30670 1540
rect 30640 1490 30670 1520
rect 30640 1470 30645 1490
rect 30665 1470 30670 1490
rect 30640 1440 30670 1470
rect 30640 1420 30645 1440
rect 30665 1420 30670 1440
rect 30640 1390 30670 1420
rect 30640 1370 30645 1390
rect 30665 1370 30670 1390
rect 30640 1340 30670 1370
rect 30640 1320 30645 1340
rect 30665 1320 30670 1340
rect 30640 1290 30670 1320
rect 30640 1270 30645 1290
rect 30665 1270 30670 1290
rect 30640 1240 30670 1270
rect 30640 1220 30645 1240
rect 30665 1220 30670 1240
rect 30640 1190 30670 1220
rect 30640 1170 30645 1190
rect 30665 1170 30670 1190
rect 30640 1140 30670 1170
rect 30640 1120 30645 1140
rect 30665 1120 30670 1140
rect 30640 1090 30670 1120
rect 30640 1070 30645 1090
rect 30665 1070 30670 1090
rect 30640 1040 30670 1070
rect 30640 1020 30645 1040
rect 30665 1020 30670 1040
rect 30640 990 30670 1020
rect 30640 970 30645 990
rect 30665 970 30670 990
rect 30640 960 30670 970
rect 30705 1345 30725 1730
rect 30940 1675 30960 1785
rect 31040 1765 31060 1785
rect 31700 1765 31720 1785
rect 31780 1765 31800 1785
rect 32000 1765 32020 1785
rect 32080 1765 32100 1785
rect 32740 1765 32760 1785
rect 31035 1755 31065 1765
rect 31237 1755 31269 1765
rect 31457 1755 31489 1765
rect 31601 1755 31633 1765
rect 31695 1755 31725 1765
rect 31035 1735 31040 1755
rect 31060 1735 31065 1755
rect 31035 1695 31065 1735
rect 31100 1745 31126 1755
rect 31100 1725 31103 1745
rect 31123 1725 31126 1745
rect 31100 1715 31126 1725
rect 31194 1745 31220 1755
rect 31194 1725 31197 1745
rect 31217 1725 31220 1745
rect 31237 1735 31243 1755
rect 31260 1735 31269 1755
rect 31237 1725 31269 1735
rect 31320 1745 31346 1755
rect 31320 1725 31323 1745
rect 31343 1725 31346 1745
rect 31194 1715 31220 1725
rect 31100 1705 31120 1715
rect 31200 1705 31220 1715
rect 31320 1715 31346 1725
rect 31414 1745 31440 1755
rect 31414 1725 31417 1745
rect 31437 1725 31440 1745
rect 31457 1735 31463 1755
rect 31480 1735 31489 1755
rect 31457 1725 31489 1735
rect 31540 1745 31566 1755
rect 31540 1725 31543 1745
rect 31563 1725 31566 1745
rect 31601 1735 31610 1755
rect 31627 1735 31633 1755
rect 31601 1725 31633 1735
rect 31650 1745 31676 1755
rect 31650 1725 31653 1745
rect 31673 1725 31676 1745
rect 31414 1715 31440 1725
rect 31320 1705 31340 1715
rect 31420 1705 31440 1715
rect 31540 1715 31566 1725
rect 31650 1715 31676 1725
rect 31695 1735 31700 1755
rect 31720 1735 31725 1755
rect 31540 1705 31560 1715
rect 31650 1705 31670 1715
rect 31035 1675 31040 1695
rect 31060 1675 31065 1695
rect 30960 1645 30980 1655
rect 30970 1625 30980 1645
rect 30960 1615 30980 1625
rect 31035 1645 31065 1675
rect 31035 1625 31040 1645
rect 31060 1625 31065 1645
rect 30940 1485 30960 1595
rect 31035 1595 31065 1625
rect 31035 1575 31040 1595
rect 31060 1575 31065 1595
rect 31035 1565 31065 1575
rect 31090 1695 31120 1705
rect 31090 1675 31095 1695
rect 31115 1675 31120 1695
rect 31090 1645 31120 1675
rect 31090 1625 31095 1645
rect 31115 1625 31120 1645
rect 31090 1595 31120 1625
rect 31090 1575 31095 1595
rect 31115 1575 31120 1595
rect 31090 1565 31120 1575
rect 31145 1695 31175 1705
rect 31145 1675 31150 1695
rect 31170 1675 31175 1695
rect 31145 1645 31175 1675
rect 31145 1625 31150 1645
rect 31170 1625 31175 1645
rect 31145 1595 31175 1625
rect 31145 1575 31150 1595
rect 31170 1575 31175 1595
rect 31145 1565 31175 1575
rect 31200 1695 31230 1705
rect 31200 1675 31205 1695
rect 31225 1675 31230 1695
rect 31200 1645 31230 1675
rect 31200 1625 31205 1645
rect 31225 1625 31230 1645
rect 31200 1595 31230 1625
rect 31200 1575 31205 1595
rect 31225 1575 31230 1595
rect 31200 1565 31230 1575
rect 31255 1695 31285 1705
rect 31255 1675 31260 1695
rect 31280 1675 31285 1695
rect 31255 1645 31285 1675
rect 31255 1625 31260 1645
rect 31280 1625 31285 1645
rect 31255 1595 31285 1625
rect 31255 1575 31260 1595
rect 31280 1575 31285 1595
rect 31255 1565 31285 1575
rect 31310 1695 31340 1705
rect 31310 1675 31315 1695
rect 31335 1675 31340 1695
rect 31310 1645 31340 1675
rect 31310 1625 31315 1645
rect 31335 1625 31340 1645
rect 31310 1595 31340 1625
rect 31310 1575 31315 1595
rect 31335 1575 31340 1595
rect 31310 1565 31340 1575
rect 31365 1695 31395 1705
rect 31365 1675 31370 1695
rect 31390 1675 31395 1695
rect 31365 1645 31395 1675
rect 31365 1625 31370 1645
rect 31390 1625 31395 1645
rect 31365 1595 31395 1625
rect 31365 1575 31370 1595
rect 31390 1575 31395 1595
rect 31365 1565 31395 1575
rect 31420 1695 31450 1705
rect 31420 1675 31425 1695
rect 31445 1675 31450 1695
rect 31420 1645 31450 1675
rect 31420 1625 31425 1645
rect 31445 1625 31450 1645
rect 31420 1595 31450 1625
rect 31420 1575 31425 1595
rect 31445 1575 31450 1595
rect 31420 1565 31450 1575
rect 31475 1695 31505 1705
rect 31475 1675 31480 1695
rect 31500 1675 31505 1695
rect 31475 1645 31505 1675
rect 31475 1625 31480 1645
rect 31500 1625 31505 1645
rect 31475 1595 31505 1625
rect 31475 1575 31480 1595
rect 31500 1575 31505 1595
rect 31475 1565 31505 1575
rect 31530 1695 31560 1705
rect 31530 1675 31535 1695
rect 31555 1675 31560 1695
rect 31530 1645 31560 1675
rect 31530 1625 31535 1645
rect 31555 1625 31560 1645
rect 31530 1595 31560 1625
rect 31530 1575 31535 1595
rect 31555 1575 31560 1595
rect 31530 1565 31560 1575
rect 31585 1695 31615 1705
rect 31585 1675 31590 1695
rect 31610 1675 31615 1695
rect 31585 1645 31615 1675
rect 31585 1625 31590 1645
rect 31610 1625 31615 1645
rect 31585 1595 31615 1625
rect 31585 1575 31590 1595
rect 31610 1575 31615 1595
rect 31585 1565 31615 1575
rect 31640 1695 31670 1705
rect 31640 1675 31645 1695
rect 31665 1675 31670 1695
rect 31640 1645 31670 1675
rect 31640 1625 31645 1645
rect 31665 1625 31670 1645
rect 31640 1595 31670 1625
rect 31640 1575 31645 1595
rect 31665 1575 31670 1595
rect 31640 1565 31670 1575
rect 31695 1695 31725 1735
rect 31695 1675 31700 1695
rect 31720 1675 31725 1695
rect 31695 1645 31725 1675
rect 31695 1625 31700 1645
rect 31720 1625 31725 1645
rect 31695 1595 31725 1625
rect 31695 1575 31700 1595
rect 31720 1575 31725 1595
rect 31695 1565 31725 1575
rect 31775 1755 31805 1765
rect 31775 1735 31780 1755
rect 31800 1735 31805 1755
rect 31775 1695 31805 1735
rect 31824 1755 31850 1765
rect 31824 1735 31827 1755
rect 31847 1735 31850 1755
rect 31824 1725 31850 1735
rect 31867 1755 31899 1765
rect 31867 1735 31873 1755
rect 31890 1735 31899 1755
rect 31867 1725 31899 1735
rect 31947 1755 31973 1765
rect 31947 1735 31950 1755
rect 31970 1735 31973 1755
rect 31947 1725 31973 1735
rect 31995 1755 32025 1765
rect 31995 1735 32000 1755
rect 32020 1735 32025 1755
rect 31775 1675 31780 1695
rect 31800 1675 31805 1695
rect 31775 1645 31805 1675
rect 31775 1625 31780 1645
rect 31800 1625 31805 1645
rect 31775 1595 31805 1625
rect 31775 1575 31780 1595
rect 31800 1575 31805 1595
rect 31775 1565 31805 1575
rect 31830 1705 31850 1725
rect 31950 1705 31970 1725
rect 31830 1695 31860 1705
rect 31830 1675 31835 1695
rect 31855 1675 31860 1695
rect 31830 1645 31860 1675
rect 31830 1625 31835 1645
rect 31855 1625 31860 1645
rect 31830 1595 31860 1625
rect 31830 1575 31835 1595
rect 31855 1575 31860 1595
rect 31830 1565 31860 1575
rect 31885 1695 31915 1705
rect 31885 1675 31890 1695
rect 31910 1675 31915 1695
rect 31885 1645 31915 1675
rect 31885 1625 31890 1645
rect 31910 1625 31915 1645
rect 31885 1595 31915 1625
rect 31885 1575 31890 1595
rect 31910 1575 31915 1595
rect 31885 1565 31915 1575
rect 31940 1695 31970 1705
rect 31940 1675 31945 1695
rect 31965 1675 31970 1695
rect 31940 1645 31970 1675
rect 31940 1625 31945 1645
rect 31965 1625 31970 1645
rect 31940 1595 31970 1625
rect 31940 1575 31945 1595
rect 31965 1575 31970 1595
rect 31940 1565 31970 1575
rect 31995 1695 32025 1735
rect 31995 1675 32000 1695
rect 32020 1675 32025 1695
rect 31995 1645 32025 1675
rect 31995 1625 32000 1645
rect 32020 1625 32025 1645
rect 31995 1595 32025 1625
rect 31995 1575 32000 1595
rect 32020 1575 32025 1595
rect 31995 1565 32025 1575
rect 32075 1755 32105 1765
rect 32277 1755 32309 1765
rect 32497 1755 32529 1765
rect 32641 1755 32673 1765
rect 32735 1755 32765 1765
rect 32075 1735 32080 1755
rect 32100 1735 32105 1755
rect 32075 1695 32105 1735
rect 32140 1745 32166 1755
rect 32140 1725 32143 1745
rect 32163 1725 32166 1745
rect 32140 1715 32166 1725
rect 32234 1745 32260 1755
rect 32234 1725 32237 1745
rect 32257 1725 32260 1745
rect 32277 1735 32283 1755
rect 32300 1735 32309 1755
rect 32277 1725 32309 1735
rect 32360 1745 32386 1755
rect 32360 1725 32363 1745
rect 32383 1725 32386 1745
rect 32234 1715 32260 1725
rect 32140 1705 32160 1715
rect 32240 1705 32260 1715
rect 32360 1715 32386 1725
rect 32454 1745 32480 1755
rect 32454 1725 32457 1745
rect 32477 1725 32480 1745
rect 32497 1735 32503 1755
rect 32520 1735 32529 1755
rect 32497 1725 32529 1735
rect 32580 1745 32606 1755
rect 32580 1725 32583 1745
rect 32603 1725 32606 1745
rect 32641 1735 32650 1755
rect 32667 1735 32673 1755
rect 32641 1725 32673 1735
rect 32690 1745 32716 1755
rect 32690 1725 32693 1745
rect 32713 1725 32716 1745
rect 32454 1715 32480 1725
rect 32360 1705 32380 1715
rect 32460 1705 32480 1715
rect 32580 1715 32606 1725
rect 32690 1715 32716 1725
rect 32735 1735 32740 1755
rect 32760 1735 32765 1755
rect 32580 1705 32600 1715
rect 32690 1705 32710 1715
rect 32075 1675 32080 1695
rect 32100 1675 32105 1695
rect 32075 1645 32105 1675
rect 32075 1625 32080 1645
rect 32100 1625 32105 1645
rect 32075 1595 32105 1625
rect 32075 1575 32080 1595
rect 32100 1575 32105 1595
rect 32075 1565 32105 1575
rect 32130 1695 32160 1705
rect 32130 1675 32135 1695
rect 32155 1675 32160 1695
rect 32130 1645 32160 1675
rect 32130 1625 32135 1645
rect 32155 1625 32160 1645
rect 32130 1595 32160 1625
rect 32130 1575 32135 1595
rect 32155 1575 32160 1595
rect 32130 1565 32160 1575
rect 32185 1695 32215 1705
rect 32185 1675 32190 1695
rect 32210 1675 32215 1695
rect 32185 1645 32215 1675
rect 32185 1625 32190 1645
rect 32210 1625 32215 1645
rect 32185 1595 32215 1625
rect 32185 1575 32190 1595
rect 32210 1575 32215 1595
rect 32185 1565 32215 1575
rect 32240 1695 32270 1705
rect 32240 1675 32245 1695
rect 32265 1675 32270 1695
rect 32240 1645 32270 1675
rect 32240 1625 32245 1645
rect 32265 1625 32270 1645
rect 32240 1595 32270 1625
rect 32240 1575 32245 1595
rect 32265 1575 32270 1595
rect 32240 1565 32270 1575
rect 32295 1695 32325 1705
rect 32295 1675 32300 1695
rect 32320 1675 32325 1695
rect 32295 1645 32325 1675
rect 32295 1625 32300 1645
rect 32320 1625 32325 1645
rect 32295 1595 32325 1625
rect 32295 1575 32300 1595
rect 32320 1575 32325 1595
rect 32295 1565 32325 1575
rect 32350 1695 32380 1705
rect 32350 1675 32355 1695
rect 32375 1675 32380 1695
rect 32350 1645 32380 1675
rect 32350 1625 32355 1645
rect 32375 1625 32380 1645
rect 32350 1595 32380 1625
rect 32350 1575 32355 1595
rect 32375 1575 32380 1595
rect 32350 1565 32380 1575
rect 32405 1695 32435 1705
rect 32405 1675 32410 1695
rect 32430 1675 32435 1695
rect 32405 1645 32435 1675
rect 32405 1625 32410 1645
rect 32430 1625 32435 1645
rect 32405 1595 32435 1625
rect 32405 1575 32410 1595
rect 32430 1575 32435 1595
rect 32405 1565 32435 1575
rect 32460 1695 32490 1705
rect 32460 1675 32465 1695
rect 32485 1675 32490 1695
rect 32460 1645 32490 1675
rect 32460 1625 32465 1645
rect 32485 1625 32490 1645
rect 32460 1595 32490 1625
rect 32460 1575 32465 1595
rect 32485 1575 32490 1595
rect 32460 1565 32490 1575
rect 32515 1695 32545 1705
rect 32515 1675 32520 1695
rect 32540 1675 32545 1695
rect 32515 1645 32545 1675
rect 32515 1625 32520 1645
rect 32540 1625 32545 1645
rect 32515 1595 32545 1625
rect 32515 1575 32520 1595
rect 32540 1575 32545 1595
rect 32515 1565 32545 1575
rect 32570 1695 32600 1705
rect 32570 1675 32575 1695
rect 32595 1675 32600 1695
rect 32570 1645 32600 1675
rect 32570 1625 32575 1645
rect 32595 1625 32600 1645
rect 32570 1595 32600 1625
rect 32570 1575 32575 1595
rect 32595 1575 32600 1595
rect 32570 1565 32600 1575
rect 32625 1695 32655 1705
rect 32625 1675 32630 1695
rect 32650 1675 32655 1695
rect 32625 1645 32655 1675
rect 32625 1625 32630 1645
rect 32650 1625 32655 1645
rect 32625 1595 32655 1625
rect 32625 1575 32630 1595
rect 32650 1575 32655 1595
rect 32625 1565 32655 1575
rect 32680 1695 32710 1705
rect 32680 1675 32685 1695
rect 32705 1675 32710 1695
rect 32680 1645 32710 1675
rect 32680 1625 32685 1645
rect 32705 1625 32710 1645
rect 32680 1595 32710 1625
rect 32680 1575 32685 1595
rect 32705 1575 32710 1595
rect 32680 1565 32710 1575
rect 32735 1695 32765 1735
rect 32735 1675 32740 1695
rect 32760 1675 32765 1695
rect 32735 1645 32765 1675
rect 32735 1625 32740 1645
rect 32760 1625 32765 1645
rect 32735 1595 32765 1625
rect 32735 1575 32740 1595
rect 32760 1575 32765 1595
rect 32735 1565 32765 1575
rect 32840 1675 32860 1785
rect 33475 1760 33515 1770
rect 33475 1750 33485 1760
rect 31155 1545 31175 1565
rect 31260 1545 31280 1565
rect 31370 1545 31390 1565
rect 31480 1545 31500 1565
rect 31590 1545 31610 1565
rect 31830 1545 31850 1565
rect 31885 1545 31905 1565
rect 32195 1545 32215 1565
rect 32300 1545 32320 1565
rect 32410 1545 32430 1565
rect 32520 1545 32540 1565
rect 32630 1545 32650 1565
rect 31106 1535 31138 1545
rect 31106 1515 31112 1535
rect 31129 1515 31138 1535
rect 31106 1505 31138 1515
rect 31155 1535 31181 1545
rect 31155 1515 31158 1535
rect 31178 1515 31181 1535
rect 31155 1505 31181 1515
rect 31256 1535 31283 1545
rect 31256 1515 31260 1535
rect 31280 1515 31283 1535
rect 31256 1505 31283 1515
rect 31305 1535 31345 1545
rect 31305 1515 31315 1535
rect 31335 1515 31345 1535
rect 31305 1505 31345 1515
rect 31366 1535 31393 1545
rect 31366 1515 31370 1535
rect 31390 1515 31393 1535
rect 31366 1505 31393 1515
rect 31476 1535 31503 1545
rect 31476 1515 31480 1535
rect 31500 1515 31503 1535
rect 31476 1505 31503 1515
rect 31525 1535 31565 1545
rect 31525 1515 31535 1535
rect 31555 1515 31565 1535
rect 31525 1505 31565 1515
rect 31586 1535 31613 1545
rect 31586 1515 31590 1535
rect 31610 1515 31613 1535
rect 31586 1505 31613 1515
rect 31825 1535 31855 1545
rect 31825 1515 31830 1535
rect 31850 1515 31855 1535
rect 31825 1505 31855 1515
rect 31875 1535 31905 1545
rect 31875 1515 31880 1535
rect 31900 1515 31905 1535
rect 31875 1505 31905 1515
rect 31922 1535 31954 1545
rect 31922 1515 31928 1535
rect 31945 1515 31954 1535
rect 31922 1505 31954 1515
rect 32146 1535 32178 1545
rect 32146 1515 32152 1535
rect 32169 1515 32178 1535
rect 32146 1505 32178 1515
rect 32195 1535 32221 1545
rect 32195 1515 32198 1535
rect 32218 1515 32221 1535
rect 32195 1505 32221 1515
rect 32296 1535 32323 1545
rect 32296 1515 32300 1535
rect 32320 1515 32323 1535
rect 32296 1505 32323 1515
rect 32345 1535 32385 1545
rect 32345 1515 32355 1535
rect 32375 1515 32385 1535
rect 32345 1505 32385 1515
rect 32406 1535 32433 1545
rect 32406 1515 32410 1535
rect 32430 1515 32433 1535
rect 32406 1505 32433 1515
rect 32516 1535 32543 1545
rect 32516 1515 32520 1535
rect 32540 1515 32543 1535
rect 32516 1505 32543 1515
rect 32565 1535 32605 1545
rect 32565 1515 32575 1535
rect 32595 1515 32605 1535
rect 32565 1505 32605 1515
rect 32626 1535 32653 1545
rect 32626 1515 32630 1535
rect 32650 1515 32653 1535
rect 32626 1505 32653 1515
rect 32840 1485 32860 1595
rect 30940 1465 31860 1485
rect 31940 1465 32860 1485
rect 33075 1730 33405 1750
rect 33505 1750 33515 1760
rect 33505 1740 33815 1750
rect 33485 1730 33815 1740
rect 33075 1345 33095 1730
rect 33135 1710 33155 1730
rect 33735 1710 33755 1730
rect 30245 940 30265 960
rect 30445 940 30465 960
rect 30235 930 30275 940
rect 30235 910 30245 930
rect 30265 910 30275 930
rect 30235 900 30275 910
rect 30435 930 30475 940
rect 30435 910 30445 930
rect 30465 910 30475 930
rect 30435 900 30475 910
rect 30705 880 30725 1265
rect 29985 860 30315 880
rect 30395 860 30725 880
rect 31155 1280 31845 1300
rect 31925 1280 32565 1300
rect 31155 1100 31175 1280
rect 31315 1250 31355 1260
rect 31315 1230 31325 1250
rect 31345 1230 31355 1250
rect 31315 1220 31355 1230
rect 31425 1250 31465 1260
rect 31425 1230 31435 1250
rect 31455 1230 31465 1250
rect 31425 1220 31465 1230
rect 31535 1250 31575 1260
rect 31535 1230 31545 1250
rect 31565 1230 31575 1250
rect 31535 1220 31575 1230
rect 31645 1250 31685 1260
rect 31645 1230 31655 1250
rect 31675 1230 31685 1250
rect 31645 1220 31685 1230
rect 31755 1250 31795 1260
rect 31755 1230 31765 1250
rect 31785 1230 31795 1250
rect 31755 1220 31795 1230
rect 31815 1250 31845 1260
rect 31815 1230 31820 1250
rect 31840 1230 31845 1250
rect 31815 1220 31845 1230
rect 31865 1250 31905 1260
rect 31865 1230 31875 1250
rect 31895 1230 31905 1250
rect 31865 1220 31905 1230
rect 31975 1250 32015 1260
rect 31975 1230 31985 1250
rect 32005 1230 32015 1250
rect 31975 1220 32015 1230
rect 32085 1250 32125 1260
rect 32085 1230 32095 1250
rect 32115 1230 32125 1250
rect 32085 1220 32125 1230
rect 32195 1250 32235 1260
rect 32195 1230 32205 1250
rect 32225 1230 32235 1250
rect 32195 1220 32235 1230
rect 32305 1250 32345 1260
rect 32305 1230 32315 1250
rect 32335 1230 32345 1250
rect 32305 1220 32345 1230
rect 32381 1250 32411 1260
rect 32381 1230 32386 1250
rect 32406 1230 32411 1250
rect 32381 1220 32411 1230
rect 32430 1250 32470 1260
rect 32430 1230 32440 1250
rect 32460 1230 32470 1250
rect 32430 1220 32470 1230
rect 31325 1200 31345 1220
rect 31435 1200 31455 1220
rect 31545 1200 31565 1220
rect 31655 1200 31675 1220
rect 31765 1200 31785 1220
rect 31875 1200 31895 1220
rect 31985 1200 32005 1220
rect 32095 1200 32115 1220
rect 32205 1200 32225 1220
rect 32315 1200 32335 1220
rect 32430 1200 32450 1220
rect 31155 875 31175 1020
rect 31210 1190 31240 1200
rect 31210 1170 31215 1190
rect 31235 1170 31240 1190
rect 31210 1140 31240 1170
rect 31210 1120 31215 1140
rect 31235 1120 31240 1140
rect 31210 1090 31240 1120
rect 31210 1070 31215 1090
rect 31235 1070 31240 1090
rect 31210 1040 31240 1070
rect 31210 1020 31215 1040
rect 31235 1020 31240 1040
rect 31210 990 31240 1020
rect 31210 970 31215 990
rect 31235 970 31240 990
rect 31210 960 31240 970
rect 31265 1190 31295 1200
rect 31265 1170 31270 1190
rect 31290 1170 31295 1190
rect 31265 1140 31295 1170
rect 31265 1120 31270 1140
rect 31290 1120 31295 1140
rect 31265 1090 31295 1120
rect 31265 1070 31270 1090
rect 31290 1070 31295 1090
rect 31265 1040 31295 1070
rect 31265 1020 31270 1040
rect 31290 1020 31295 1040
rect 31265 990 31295 1020
rect 31265 970 31270 990
rect 31290 970 31295 990
rect 31265 960 31295 970
rect 31320 1190 31350 1200
rect 31320 1170 31325 1190
rect 31345 1170 31350 1190
rect 31320 1140 31350 1170
rect 31320 1120 31325 1140
rect 31345 1120 31350 1140
rect 31320 1090 31350 1120
rect 31320 1070 31325 1090
rect 31345 1070 31350 1090
rect 31320 1040 31350 1070
rect 31320 1020 31325 1040
rect 31345 1020 31350 1040
rect 31320 990 31350 1020
rect 31320 970 31325 990
rect 31345 970 31350 990
rect 31320 960 31350 970
rect 31375 1190 31405 1200
rect 31375 1170 31380 1190
rect 31400 1170 31405 1190
rect 31375 1140 31405 1170
rect 31375 1120 31380 1140
rect 31400 1120 31405 1140
rect 31375 1090 31405 1120
rect 31375 1070 31380 1090
rect 31400 1070 31405 1090
rect 31375 1040 31405 1070
rect 31375 1020 31380 1040
rect 31400 1020 31405 1040
rect 31375 990 31405 1020
rect 31375 970 31380 990
rect 31400 970 31405 990
rect 31375 960 31405 970
rect 31430 1190 31460 1200
rect 31430 1170 31435 1190
rect 31455 1170 31460 1190
rect 31430 1140 31460 1170
rect 31430 1120 31435 1140
rect 31455 1120 31460 1140
rect 31430 1090 31460 1120
rect 31430 1070 31435 1090
rect 31455 1070 31460 1090
rect 31430 1040 31460 1070
rect 31430 1020 31435 1040
rect 31455 1020 31460 1040
rect 31430 990 31460 1020
rect 31430 970 31435 990
rect 31455 970 31460 990
rect 31430 960 31460 970
rect 31485 1190 31515 1200
rect 31485 1170 31490 1190
rect 31510 1170 31515 1190
rect 31485 1140 31515 1170
rect 31485 1120 31490 1140
rect 31510 1120 31515 1140
rect 31485 1090 31515 1120
rect 31485 1070 31490 1090
rect 31510 1070 31515 1090
rect 31485 1040 31515 1070
rect 31485 1020 31490 1040
rect 31510 1020 31515 1040
rect 31485 990 31515 1020
rect 31485 970 31490 990
rect 31510 970 31515 990
rect 31485 960 31515 970
rect 31540 1190 31570 1200
rect 31540 1170 31545 1190
rect 31565 1170 31570 1190
rect 31540 1140 31570 1170
rect 31540 1120 31545 1140
rect 31565 1120 31570 1140
rect 31540 1090 31570 1120
rect 31540 1070 31545 1090
rect 31565 1070 31570 1090
rect 31540 1040 31570 1070
rect 31540 1020 31545 1040
rect 31565 1020 31570 1040
rect 31540 990 31570 1020
rect 31540 970 31545 990
rect 31565 970 31570 990
rect 31540 960 31570 970
rect 31595 1190 31625 1200
rect 31595 1170 31600 1190
rect 31620 1170 31625 1190
rect 31595 1140 31625 1170
rect 31595 1120 31600 1140
rect 31620 1120 31625 1140
rect 31595 1090 31625 1120
rect 31595 1070 31600 1090
rect 31620 1070 31625 1090
rect 31595 1040 31625 1070
rect 31595 1020 31600 1040
rect 31620 1020 31625 1040
rect 31595 990 31625 1020
rect 31595 970 31600 990
rect 31620 970 31625 990
rect 31595 960 31625 970
rect 31650 1190 31680 1200
rect 31650 1170 31655 1190
rect 31675 1170 31680 1190
rect 31650 1140 31680 1170
rect 31650 1120 31655 1140
rect 31675 1120 31680 1140
rect 31650 1090 31680 1120
rect 31650 1070 31655 1090
rect 31675 1070 31680 1090
rect 31650 1040 31680 1070
rect 31650 1020 31655 1040
rect 31675 1020 31680 1040
rect 31650 990 31680 1020
rect 31650 970 31655 990
rect 31675 970 31680 990
rect 31650 960 31680 970
rect 31705 1190 31735 1200
rect 31705 1170 31710 1190
rect 31730 1170 31735 1190
rect 31705 1140 31735 1170
rect 31705 1120 31710 1140
rect 31730 1120 31735 1140
rect 31705 1090 31735 1120
rect 31705 1070 31710 1090
rect 31730 1070 31735 1090
rect 31705 1040 31735 1070
rect 31705 1020 31710 1040
rect 31730 1020 31735 1040
rect 31705 990 31735 1020
rect 31705 970 31710 990
rect 31730 970 31735 990
rect 31705 960 31735 970
rect 31760 1190 31790 1200
rect 31760 1170 31765 1190
rect 31785 1170 31790 1190
rect 31760 1140 31790 1170
rect 31760 1120 31765 1140
rect 31785 1120 31790 1140
rect 31760 1090 31790 1120
rect 31760 1070 31765 1090
rect 31785 1070 31790 1090
rect 31760 1040 31790 1070
rect 31760 1020 31765 1040
rect 31785 1020 31790 1040
rect 31760 990 31790 1020
rect 31760 970 31765 990
rect 31785 970 31790 990
rect 31760 960 31790 970
rect 31815 1190 31845 1200
rect 31815 1170 31820 1190
rect 31840 1170 31845 1190
rect 31815 1140 31845 1170
rect 31815 1120 31820 1140
rect 31840 1120 31845 1140
rect 31815 1090 31845 1120
rect 31815 1070 31820 1090
rect 31840 1070 31845 1090
rect 31815 1040 31845 1070
rect 31815 1020 31820 1040
rect 31840 1020 31845 1040
rect 31815 990 31845 1020
rect 31815 970 31820 990
rect 31840 970 31845 990
rect 31815 960 31845 970
rect 31870 1190 31900 1200
rect 31870 1170 31875 1190
rect 31895 1170 31900 1190
rect 31870 1140 31900 1170
rect 31870 1120 31875 1140
rect 31895 1120 31900 1140
rect 31870 1090 31900 1120
rect 31870 1070 31875 1090
rect 31895 1070 31900 1090
rect 31870 1040 31900 1070
rect 31870 1020 31875 1040
rect 31895 1020 31900 1040
rect 31870 990 31900 1020
rect 31870 970 31875 990
rect 31895 970 31900 990
rect 31870 960 31900 970
rect 31925 1190 31955 1200
rect 31925 1170 31930 1190
rect 31950 1170 31955 1190
rect 31925 1140 31955 1170
rect 31925 1120 31930 1140
rect 31950 1120 31955 1140
rect 31925 1090 31955 1120
rect 31925 1070 31930 1090
rect 31950 1070 31955 1090
rect 31925 1040 31955 1070
rect 31925 1020 31930 1040
rect 31950 1020 31955 1040
rect 31925 990 31955 1020
rect 31925 970 31930 990
rect 31950 970 31955 990
rect 31925 960 31955 970
rect 31980 1190 32010 1200
rect 31980 1170 31985 1190
rect 32005 1170 32010 1190
rect 31980 1140 32010 1170
rect 31980 1120 31985 1140
rect 32005 1120 32010 1140
rect 31980 1090 32010 1120
rect 31980 1070 31985 1090
rect 32005 1070 32010 1090
rect 31980 1040 32010 1070
rect 31980 1020 31985 1040
rect 32005 1020 32010 1040
rect 31980 990 32010 1020
rect 31980 970 31985 990
rect 32005 970 32010 990
rect 31980 960 32010 970
rect 32035 1190 32065 1200
rect 32035 1170 32040 1190
rect 32060 1170 32065 1190
rect 32035 1140 32065 1170
rect 32035 1120 32040 1140
rect 32060 1120 32065 1140
rect 32035 1090 32065 1120
rect 32035 1070 32040 1090
rect 32060 1070 32065 1090
rect 32035 1040 32065 1070
rect 32035 1020 32040 1040
rect 32060 1020 32065 1040
rect 32035 990 32065 1020
rect 32035 970 32040 990
rect 32060 970 32065 990
rect 32035 960 32065 970
rect 32090 1190 32120 1200
rect 32090 1170 32095 1190
rect 32115 1170 32120 1190
rect 32090 1140 32120 1170
rect 32090 1120 32095 1140
rect 32115 1120 32120 1140
rect 32090 1090 32120 1120
rect 32090 1070 32095 1090
rect 32115 1070 32120 1090
rect 32090 1040 32120 1070
rect 32090 1020 32095 1040
rect 32115 1020 32120 1040
rect 32090 990 32120 1020
rect 32090 970 32095 990
rect 32115 970 32120 990
rect 32090 960 32120 970
rect 32145 1190 32175 1200
rect 32145 1170 32150 1190
rect 32170 1170 32175 1190
rect 32145 1140 32175 1170
rect 32145 1120 32150 1140
rect 32170 1120 32175 1140
rect 32145 1090 32175 1120
rect 32145 1070 32150 1090
rect 32170 1070 32175 1090
rect 32145 1040 32175 1070
rect 32145 1020 32150 1040
rect 32170 1020 32175 1040
rect 32145 990 32175 1020
rect 32145 970 32150 990
rect 32170 970 32175 990
rect 32145 960 32175 970
rect 32200 1190 32230 1200
rect 32200 1170 32205 1190
rect 32225 1170 32230 1190
rect 32200 1140 32230 1170
rect 32200 1120 32205 1140
rect 32225 1120 32230 1140
rect 32200 1090 32230 1120
rect 32200 1070 32205 1090
rect 32225 1070 32230 1090
rect 32200 1040 32230 1070
rect 32200 1020 32205 1040
rect 32225 1020 32230 1040
rect 32200 990 32230 1020
rect 32200 970 32205 990
rect 32225 970 32230 990
rect 32200 960 32230 970
rect 32255 1190 32285 1200
rect 32255 1170 32260 1190
rect 32280 1170 32285 1190
rect 32255 1140 32285 1170
rect 32255 1120 32260 1140
rect 32280 1120 32285 1140
rect 32255 1090 32285 1120
rect 32255 1070 32260 1090
rect 32280 1070 32285 1090
rect 32255 1040 32285 1070
rect 32255 1020 32260 1040
rect 32280 1020 32285 1040
rect 32255 990 32285 1020
rect 32255 970 32260 990
rect 32280 970 32285 990
rect 32255 960 32285 970
rect 32310 1190 32340 1200
rect 32310 1170 32315 1190
rect 32335 1170 32340 1190
rect 32310 1140 32340 1170
rect 32310 1120 32315 1140
rect 32335 1120 32340 1140
rect 32310 1090 32340 1120
rect 32310 1070 32315 1090
rect 32335 1070 32340 1090
rect 32310 1040 32340 1070
rect 32310 1020 32315 1040
rect 32335 1020 32340 1040
rect 32310 990 32340 1020
rect 32310 970 32315 990
rect 32335 970 32340 990
rect 32310 960 32340 970
rect 32365 1190 32395 1200
rect 32365 1170 32370 1190
rect 32390 1170 32395 1190
rect 32365 1140 32395 1170
rect 32365 1120 32370 1140
rect 32390 1120 32395 1140
rect 32365 1090 32395 1120
rect 32365 1070 32370 1090
rect 32390 1070 32395 1090
rect 32365 1040 32395 1070
rect 32365 1020 32370 1040
rect 32390 1020 32395 1040
rect 32365 990 32395 1020
rect 32365 970 32370 990
rect 32390 970 32395 990
rect 32365 960 32395 970
rect 32420 1190 32450 1200
rect 32420 1170 32425 1190
rect 32445 1170 32450 1190
rect 32420 1140 32450 1170
rect 32420 1120 32425 1140
rect 32445 1120 32450 1140
rect 32420 1090 32450 1120
rect 32420 1070 32425 1090
rect 32445 1070 32450 1090
rect 32420 1040 32450 1070
rect 32420 1020 32425 1040
rect 32445 1020 32450 1040
rect 32420 990 32450 1020
rect 32420 970 32425 990
rect 32445 970 32450 990
rect 32420 960 32450 970
rect 32475 1190 32505 1200
rect 32475 1170 32480 1190
rect 32500 1170 32505 1190
rect 32475 1140 32505 1170
rect 32475 1120 32480 1140
rect 32500 1120 32505 1140
rect 32475 1090 32505 1120
rect 32475 1070 32480 1090
rect 32500 1070 32505 1090
rect 32475 1040 32505 1070
rect 32475 1020 32480 1040
rect 32500 1020 32505 1040
rect 32475 990 32505 1020
rect 32475 970 32480 990
rect 32500 970 32505 990
rect 32475 960 32505 970
rect 32545 1100 32565 1280
rect 31215 940 31235 960
rect 31270 940 31290 960
rect 31380 940 31400 960
rect 31490 940 31510 960
rect 31600 940 31620 960
rect 31710 940 31730 960
rect 31820 940 31840 960
rect 31930 940 31950 960
rect 32040 940 32060 960
rect 32150 940 32170 960
rect 32260 940 32280 960
rect 32370 940 32390 960
rect 32480 940 32500 960
rect 31195 930 31235 940
rect 31195 910 31205 930
rect 31225 910 31235 930
rect 31195 900 31235 910
rect 31260 930 31300 940
rect 31260 910 31270 930
rect 31290 910 31300 930
rect 31260 900 31300 910
rect 31370 930 31410 940
rect 31370 910 31380 930
rect 31400 910 31410 930
rect 31370 900 31410 910
rect 31480 930 31520 940
rect 31480 910 31490 930
rect 31510 910 31520 930
rect 31480 900 31520 910
rect 31590 930 31630 940
rect 31590 910 31600 930
rect 31620 910 31630 930
rect 31590 900 31630 910
rect 31700 930 31740 940
rect 31700 910 31710 930
rect 31730 910 31740 930
rect 31700 900 31740 910
rect 31810 930 31850 940
rect 31810 910 31820 930
rect 31840 910 31850 930
rect 31810 900 31850 910
rect 31920 930 31960 940
rect 31920 910 31930 930
rect 31950 910 31960 930
rect 31920 900 31960 910
rect 32030 930 32070 940
rect 32030 910 32040 930
rect 32060 910 32070 930
rect 32030 900 32070 910
rect 32140 930 32180 940
rect 32140 910 32150 930
rect 32170 910 32180 930
rect 32140 900 32180 910
rect 32250 930 32290 940
rect 32250 910 32260 930
rect 32280 910 32290 930
rect 32250 900 32290 910
rect 32360 930 32400 940
rect 32360 910 32370 930
rect 32390 910 32400 930
rect 32360 900 32400 910
rect 32475 930 32515 940
rect 32475 910 32485 930
rect 32505 910 32515 930
rect 32475 900 32515 910
rect 31205 875 31225 900
rect 32485 875 32505 900
rect 32545 875 32565 1020
rect 30335 850 30345 860
rect 30365 850 30375 860
rect 31155 855 31845 875
rect 31925 855 32565 875
rect 33075 880 33095 1265
rect 33130 1700 33160 1710
rect 33130 1680 33135 1700
rect 33155 1680 33160 1700
rect 33130 1640 33160 1680
rect 33225 1700 33265 1710
rect 33225 1680 33235 1700
rect 33255 1680 33265 1700
rect 33225 1670 33265 1680
rect 33328 1700 33362 1710
rect 33328 1680 33336 1700
rect 33354 1680 33362 1700
rect 33328 1670 33362 1680
rect 33425 1700 33465 1710
rect 33425 1680 33435 1700
rect 33455 1680 33465 1700
rect 33425 1670 33465 1680
rect 33625 1700 33665 1710
rect 33625 1680 33635 1700
rect 33655 1680 33665 1700
rect 33625 1670 33665 1680
rect 33730 1700 33760 1710
rect 33730 1680 33735 1700
rect 33755 1680 33760 1700
rect 33235 1650 33255 1670
rect 33435 1650 33455 1670
rect 33635 1650 33655 1670
rect 33130 1620 33135 1640
rect 33155 1620 33160 1640
rect 33130 1590 33160 1620
rect 33130 1570 33135 1590
rect 33155 1570 33160 1590
rect 33130 1540 33160 1570
rect 33130 1520 33135 1540
rect 33155 1520 33160 1540
rect 33130 1490 33160 1520
rect 33130 1470 33135 1490
rect 33155 1470 33160 1490
rect 33130 1440 33160 1470
rect 33130 1420 33135 1440
rect 33155 1420 33160 1440
rect 33130 1390 33160 1420
rect 33130 1370 33135 1390
rect 33155 1370 33160 1390
rect 33130 1340 33160 1370
rect 33130 1320 33135 1340
rect 33155 1320 33160 1340
rect 33130 1290 33160 1320
rect 33130 1270 33135 1290
rect 33155 1270 33160 1290
rect 33130 1240 33160 1270
rect 33130 1220 33135 1240
rect 33155 1220 33160 1240
rect 33130 1190 33160 1220
rect 33130 1170 33135 1190
rect 33155 1170 33160 1190
rect 33130 1140 33160 1170
rect 33130 1120 33135 1140
rect 33155 1120 33160 1140
rect 33130 1090 33160 1120
rect 33130 1070 33135 1090
rect 33155 1070 33160 1090
rect 33130 1040 33160 1070
rect 33130 1020 33135 1040
rect 33155 1020 33160 1040
rect 33130 990 33160 1020
rect 33130 970 33135 990
rect 33155 970 33160 990
rect 33130 960 33160 970
rect 33230 1640 33260 1650
rect 33230 1620 33235 1640
rect 33255 1620 33260 1640
rect 33230 1590 33260 1620
rect 33230 1570 33235 1590
rect 33255 1570 33260 1590
rect 33230 1540 33260 1570
rect 33230 1520 33235 1540
rect 33255 1520 33260 1540
rect 33230 1490 33260 1520
rect 33230 1470 33235 1490
rect 33255 1470 33260 1490
rect 33230 1440 33260 1470
rect 33230 1420 33235 1440
rect 33255 1420 33260 1440
rect 33230 1390 33260 1420
rect 33230 1370 33235 1390
rect 33255 1370 33260 1390
rect 33230 1340 33260 1370
rect 33230 1320 33235 1340
rect 33255 1320 33260 1340
rect 33230 1290 33260 1320
rect 33230 1270 33235 1290
rect 33255 1270 33260 1290
rect 33230 1240 33260 1270
rect 33230 1220 33235 1240
rect 33255 1220 33260 1240
rect 33230 1190 33260 1220
rect 33230 1170 33235 1190
rect 33255 1170 33260 1190
rect 33230 1140 33260 1170
rect 33230 1120 33235 1140
rect 33255 1120 33260 1140
rect 33230 1090 33260 1120
rect 33230 1070 33235 1090
rect 33255 1070 33260 1090
rect 33230 1040 33260 1070
rect 33230 1020 33235 1040
rect 33255 1020 33260 1040
rect 33230 990 33260 1020
rect 33230 970 33235 990
rect 33255 970 33260 990
rect 33230 960 33260 970
rect 33330 1640 33360 1650
rect 33330 1620 33335 1640
rect 33355 1620 33360 1640
rect 33330 1590 33360 1620
rect 33330 1570 33335 1590
rect 33355 1570 33360 1590
rect 33330 1540 33360 1570
rect 33330 1520 33335 1540
rect 33355 1520 33360 1540
rect 33330 1490 33360 1520
rect 33330 1470 33335 1490
rect 33355 1470 33360 1490
rect 33330 1440 33360 1470
rect 33330 1420 33335 1440
rect 33355 1420 33360 1440
rect 33330 1390 33360 1420
rect 33330 1370 33335 1390
rect 33355 1370 33360 1390
rect 33330 1340 33360 1370
rect 33330 1320 33335 1340
rect 33355 1320 33360 1340
rect 33330 1290 33360 1320
rect 33330 1270 33335 1290
rect 33355 1270 33360 1290
rect 33330 1240 33360 1270
rect 33330 1220 33335 1240
rect 33355 1220 33360 1240
rect 33330 1190 33360 1220
rect 33330 1170 33335 1190
rect 33355 1170 33360 1190
rect 33330 1140 33360 1170
rect 33330 1120 33335 1140
rect 33355 1120 33360 1140
rect 33330 1090 33360 1120
rect 33330 1070 33335 1090
rect 33355 1070 33360 1090
rect 33330 1040 33360 1070
rect 33330 1020 33335 1040
rect 33355 1020 33360 1040
rect 33330 990 33360 1020
rect 33330 970 33335 990
rect 33355 970 33360 990
rect 33330 960 33360 970
rect 33430 1640 33460 1650
rect 33430 1620 33435 1640
rect 33455 1620 33460 1640
rect 33430 1590 33460 1620
rect 33430 1570 33435 1590
rect 33455 1570 33460 1590
rect 33430 1540 33460 1570
rect 33430 1520 33435 1540
rect 33455 1520 33460 1540
rect 33430 1490 33460 1520
rect 33430 1470 33435 1490
rect 33455 1470 33460 1490
rect 33430 1440 33460 1470
rect 33430 1420 33435 1440
rect 33455 1420 33460 1440
rect 33430 1390 33460 1420
rect 33430 1370 33435 1390
rect 33455 1370 33460 1390
rect 33430 1340 33460 1370
rect 33430 1320 33435 1340
rect 33455 1320 33460 1340
rect 33430 1290 33460 1320
rect 33430 1270 33435 1290
rect 33455 1270 33460 1290
rect 33430 1240 33460 1270
rect 33430 1220 33435 1240
rect 33455 1220 33460 1240
rect 33430 1190 33460 1220
rect 33430 1170 33435 1190
rect 33455 1170 33460 1190
rect 33430 1140 33460 1170
rect 33430 1120 33435 1140
rect 33455 1120 33460 1140
rect 33430 1090 33460 1120
rect 33430 1070 33435 1090
rect 33455 1070 33460 1090
rect 33430 1040 33460 1070
rect 33430 1020 33435 1040
rect 33455 1020 33460 1040
rect 33430 990 33460 1020
rect 33430 970 33435 990
rect 33455 970 33460 990
rect 33430 960 33460 970
rect 33530 1640 33560 1650
rect 33530 1620 33535 1640
rect 33555 1620 33560 1640
rect 33530 1590 33560 1620
rect 33530 1570 33535 1590
rect 33555 1570 33560 1590
rect 33530 1540 33560 1570
rect 33530 1520 33535 1540
rect 33555 1520 33560 1540
rect 33530 1490 33560 1520
rect 33530 1470 33535 1490
rect 33555 1470 33560 1490
rect 33530 1440 33560 1470
rect 33530 1420 33535 1440
rect 33555 1420 33560 1440
rect 33530 1390 33560 1420
rect 33530 1370 33535 1390
rect 33555 1370 33560 1390
rect 33530 1340 33560 1370
rect 33530 1320 33535 1340
rect 33555 1320 33560 1340
rect 33530 1290 33560 1320
rect 33530 1270 33535 1290
rect 33555 1270 33560 1290
rect 33530 1240 33560 1270
rect 33530 1220 33535 1240
rect 33555 1220 33560 1240
rect 33530 1190 33560 1220
rect 33530 1170 33535 1190
rect 33555 1170 33560 1190
rect 33530 1140 33560 1170
rect 33530 1120 33535 1140
rect 33555 1120 33560 1140
rect 33530 1090 33560 1120
rect 33530 1070 33535 1090
rect 33555 1070 33560 1090
rect 33530 1040 33560 1070
rect 33530 1020 33535 1040
rect 33555 1020 33560 1040
rect 33530 990 33560 1020
rect 33530 970 33535 990
rect 33555 970 33560 990
rect 33530 960 33560 970
rect 33630 1640 33660 1650
rect 33630 1620 33635 1640
rect 33655 1620 33660 1640
rect 33630 1590 33660 1620
rect 33630 1570 33635 1590
rect 33655 1570 33660 1590
rect 33630 1540 33660 1570
rect 33630 1520 33635 1540
rect 33655 1520 33660 1540
rect 33630 1490 33660 1520
rect 33630 1470 33635 1490
rect 33655 1470 33660 1490
rect 33630 1440 33660 1470
rect 33630 1420 33635 1440
rect 33655 1420 33660 1440
rect 33630 1390 33660 1420
rect 33630 1370 33635 1390
rect 33655 1370 33660 1390
rect 33630 1340 33660 1370
rect 33630 1320 33635 1340
rect 33655 1320 33660 1340
rect 33630 1290 33660 1320
rect 33630 1270 33635 1290
rect 33655 1270 33660 1290
rect 33630 1240 33660 1270
rect 33630 1220 33635 1240
rect 33655 1220 33660 1240
rect 33630 1190 33660 1220
rect 33630 1170 33635 1190
rect 33655 1170 33660 1190
rect 33630 1140 33660 1170
rect 33630 1120 33635 1140
rect 33655 1120 33660 1140
rect 33630 1090 33660 1120
rect 33630 1070 33635 1090
rect 33655 1070 33660 1090
rect 33630 1040 33660 1070
rect 33630 1020 33635 1040
rect 33655 1020 33660 1040
rect 33630 990 33660 1020
rect 33630 970 33635 990
rect 33655 970 33660 990
rect 33630 960 33660 970
rect 33730 1640 33760 1680
rect 33730 1620 33735 1640
rect 33755 1620 33760 1640
rect 33730 1590 33760 1620
rect 33730 1570 33735 1590
rect 33755 1570 33760 1590
rect 33730 1540 33760 1570
rect 33730 1520 33735 1540
rect 33755 1520 33760 1540
rect 33730 1490 33760 1520
rect 33730 1470 33735 1490
rect 33755 1470 33760 1490
rect 33730 1440 33760 1470
rect 33730 1420 33735 1440
rect 33755 1420 33760 1440
rect 33730 1390 33760 1420
rect 33730 1370 33735 1390
rect 33755 1370 33760 1390
rect 33730 1340 33760 1370
rect 33730 1320 33735 1340
rect 33755 1320 33760 1340
rect 33730 1290 33760 1320
rect 33730 1270 33735 1290
rect 33755 1270 33760 1290
rect 33730 1240 33760 1270
rect 33730 1220 33735 1240
rect 33755 1220 33760 1240
rect 33730 1190 33760 1220
rect 33730 1170 33735 1190
rect 33755 1170 33760 1190
rect 33730 1140 33760 1170
rect 33730 1120 33735 1140
rect 33755 1120 33760 1140
rect 33730 1090 33760 1120
rect 33730 1070 33735 1090
rect 33755 1070 33760 1090
rect 33730 1040 33760 1070
rect 33730 1020 33735 1040
rect 33755 1020 33760 1040
rect 33730 990 33760 1020
rect 33730 970 33735 990
rect 33755 970 33760 990
rect 33730 960 33760 970
rect 33795 1345 33815 1730
rect 33905 1675 33985 1695
rect 34065 1675 34140 1695
rect 33905 1325 33925 1675
rect 33975 1640 34010 1650
rect 33975 1615 33980 1640
rect 34005 1615 34010 1640
rect 33975 1605 34010 1615
rect 34035 1640 34070 1650
rect 34035 1615 34040 1640
rect 34065 1615 34070 1640
rect 34035 1605 34070 1615
rect 33815 1315 33835 1325
rect 33825 1295 33835 1315
rect 33815 1285 33835 1295
rect 33885 1315 33925 1325
rect 33885 1295 33895 1315
rect 33915 1300 33925 1315
rect 33885 1285 33905 1295
rect 33335 940 33355 960
rect 33535 940 33555 960
rect 33325 930 33365 940
rect 33325 910 33335 930
rect 33355 910 33365 930
rect 33325 900 33365 910
rect 33525 930 33565 940
rect 33525 910 33535 930
rect 33555 910 33565 930
rect 33525 900 33565 910
rect 33795 880 33815 1265
rect 33075 860 33405 880
rect 33485 860 33815 880
rect 33905 868 33925 1220
rect 34120 1300 34140 1675
rect 34010 918 34035 968
rect 34120 868 34140 1220
rect 30335 840 30375 850
rect 33425 850 33435 860
rect 33455 850 33465 860
rect 33425 840 33465 850
rect 33905 848 33985 868
rect 34065 848 34140 868
rect 31210 765 31355 785
rect 31435 765 31585 785
rect 31210 695 31230 765
rect 31305 735 31345 745
rect 31305 725 31315 735
rect 31275 715 31315 725
rect 31335 715 31345 735
rect 31275 705 31345 715
rect 31375 735 31415 745
rect 31375 715 31385 735
rect 31405 715 31415 735
rect 31375 705 31415 715
rect 31445 735 31485 745
rect 31445 715 31455 735
rect 31475 715 31485 735
rect 31445 705 31485 715
rect 31505 735 31545 745
rect 31505 715 31515 735
rect 31535 715 31545 735
rect 31505 705 31545 715
rect 31275 685 31295 705
rect 31505 685 31525 705
rect 31210 555 31230 615
rect 31265 675 31295 685
rect 31265 655 31270 675
rect 31290 655 31295 675
rect 31265 625 31295 655
rect 31265 605 31270 625
rect 31290 605 31295 625
rect 31265 595 31295 605
rect 31495 675 31525 685
rect 31495 655 31500 675
rect 31520 655 31525 675
rect 31495 625 31525 655
rect 31495 605 31500 625
rect 31520 605 31525 625
rect 31495 595 31525 605
rect 31565 695 31585 765
rect 31565 555 31585 615
rect 31210 535 31355 555
rect 31435 535 31585 555
rect 31830 760 32190 780
rect 32270 760 32630 780
rect 31830 690 31850 760
rect 31890 740 31910 760
rect 32550 740 32570 760
rect 31885 730 31915 740
rect 31885 710 31890 730
rect 31910 710 31915 730
rect 31885 670 31915 710
rect 31935 730 31975 740
rect 31935 710 31945 730
rect 31965 710 31975 730
rect 31935 700 31975 710
rect 32045 730 32085 740
rect 32045 710 32055 730
rect 32075 710 32085 730
rect 32045 700 32085 710
rect 32155 730 32195 740
rect 32155 710 32165 730
rect 32185 710 32195 730
rect 32155 700 32195 710
rect 32265 730 32305 740
rect 32265 710 32275 730
rect 32295 710 32305 730
rect 32265 700 32305 710
rect 32375 730 32415 740
rect 32375 710 32385 730
rect 32405 710 32415 730
rect 32375 700 32415 710
rect 32485 730 32525 740
rect 32485 710 32495 730
rect 32515 710 32525 730
rect 32485 700 32525 710
rect 32545 730 32575 740
rect 32545 710 32550 730
rect 32570 710 32575 730
rect 31945 680 31965 700
rect 32055 680 32075 700
rect 32165 680 32185 700
rect 32275 680 32295 700
rect 32385 680 32405 700
rect 32495 680 32515 700
rect 31885 650 31890 670
rect 31910 650 31915 670
rect 31885 640 31915 650
rect 31940 670 31970 680
rect 31940 650 31945 670
rect 31965 650 31970 670
rect 31940 640 31970 650
rect 31995 670 32025 680
rect 31995 650 32000 670
rect 32020 650 32025 670
rect 31995 640 32025 650
rect 32050 670 32080 680
rect 32050 650 32055 670
rect 32075 650 32080 670
rect 32050 640 32080 650
rect 32105 670 32135 680
rect 32105 650 32110 670
rect 32130 650 32135 670
rect 32105 640 32135 650
rect 32160 670 32190 680
rect 32160 650 32165 670
rect 32185 650 32190 670
rect 32160 640 32190 650
rect 32215 670 32245 680
rect 32215 650 32220 670
rect 32240 650 32245 670
rect 32215 640 32245 650
rect 32270 670 32300 680
rect 32270 650 32275 670
rect 32295 650 32300 670
rect 32270 640 32300 650
rect 32325 670 32355 680
rect 32325 650 32330 670
rect 32350 650 32355 670
rect 32325 640 32355 650
rect 32380 670 32410 680
rect 32380 650 32385 670
rect 32405 650 32410 670
rect 32380 640 32410 650
rect 32435 670 32465 680
rect 32435 650 32440 670
rect 32460 650 32465 670
rect 32435 640 32465 650
rect 32490 670 32520 680
rect 32490 650 32495 670
rect 32515 650 32520 670
rect 32490 640 32520 650
rect 32545 670 32575 710
rect 32545 650 32550 670
rect 32570 650 32575 670
rect 32545 640 32575 650
rect 32610 690 32630 760
rect 32000 620 32020 640
rect 32110 620 32130 640
rect 32220 620 32240 640
rect 32330 620 32350 640
rect 32440 620 32460 640
rect 31830 560 31850 610
rect 31990 610 32030 620
rect 31990 590 32000 610
rect 32020 590 32030 610
rect 31990 580 32030 590
rect 32100 610 32140 620
rect 32100 590 32110 610
rect 32130 590 32140 610
rect 32100 580 32140 590
rect 32210 610 32250 620
rect 32210 590 32220 610
rect 32240 590 32250 610
rect 32210 580 32250 590
rect 32320 610 32360 620
rect 32320 590 32330 610
rect 32350 590 32360 610
rect 32320 580 32360 590
rect 32430 610 32470 620
rect 32430 590 32440 610
rect 32460 590 32470 610
rect 32430 580 32470 590
rect 32610 560 32630 610
rect 31830 540 32190 560
rect 32270 540 32630 560
rect 31375 525 31385 535
rect 31405 525 31415 535
rect 31375 515 31415 525
rect 32210 530 32220 540
rect 32240 530 32250 540
rect 32210 520 32250 530
<< viali >>
rect 31290 4845 31310 4865
rect 31480 4860 31500 4880
rect 31540 4860 31560 4880
rect 31600 4860 31620 4880
rect 31660 4860 31680 4880
rect 31720 4860 31740 4880
rect 31780 4860 31800 4880
rect 31840 4860 31860 4880
rect 31320 4710 31340 4730
rect 31660 4705 31680 4725
rect 32210 4835 32230 4855
rect 32330 4835 32350 4855
rect 32450 4835 32470 4855
rect 32570 4835 32590 4855
rect 32690 4835 32710 4855
rect 32270 4705 32290 4725
rect 32331 4705 32349 4725
rect 32390 4705 32410 4725
rect 32510 4705 32530 4725
rect 32630 4705 32650 4725
rect 31260 4415 31280 4435
rect 31370 4415 31390 4435
rect 31480 4415 31500 4435
rect 31590 4415 31610 4435
rect 31700 4415 31720 4435
rect 31810 4415 31830 4435
rect 31920 4415 31940 4435
rect 32030 4415 32050 4435
rect 32140 4415 32160 4435
rect 32250 4415 32270 4435
rect 32360 4415 32380 4435
rect 32470 4415 32490 4435
rect 31315 4295 31335 4315
rect 31370 4295 31390 4315
rect 31425 4295 31445 4315
rect 31535 4295 31555 4315
rect 31645 4295 31665 4315
rect 31755 4295 31775 4315
rect 31865 4295 31885 4315
rect 31975 4295 31995 4315
rect 32085 4295 32105 4315
rect 32195 4295 32215 4315
rect 32305 4295 32325 4315
rect 32415 4295 32435 4315
rect 31285 4005 31305 4025
rect 31330 4005 31350 4025
rect 31375 4005 31395 4025
rect 31430 4005 31450 4025
rect 31485 4005 31505 4025
rect 31540 4005 31560 4025
rect 31650 4005 31670 4025
rect 31705 4005 31725 4025
rect 31760 4005 31780 4025
rect 32013 4005 32033 4025
rect 32060 4005 32080 4025
rect 32160 4005 32180 4025
rect 32215 4005 32235 4025
rect 32270 4005 32290 4025
rect 32380 4005 32400 4025
rect 32435 4005 32455 4025
rect 32490 4005 32510 4025
rect 31150 3945 31170 3965
rect 31265 3885 31285 3905
rect 31360 3885 31380 3905
rect 31413 3885 31430 3905
rect 31485 3885 31505 3905
rect 31580 3885 31600 3905
rect 31633 3885 31650 3905
rect 31705 3885 31725 3905
rect 31780 3885 31797 3905
rect 31823 3885 31843 3905
rect 31995 3885 32015 3905
rect 32090 3885 32110 3905
rect 32143 3885 32160 3905
rect 32215 3885 32235 3905
rect 32310 3885 32330 3905
rect 32363 3885 32380 3905
rect 32435 3885 32455 3905
rect 32510 3885 32527 3905
rect 32553 3885 32573 3905
rect 29560 3625 29590 3655
rect 29610 3625 29640 3655
rect 29659 3625 29689 3655
rect 29560 3020 29590 3050
rect 29610 3020 29640 3050
rect 29659 3020 29689 3050
rect 29535 2965 29555 2985
rect 29965 3690 29985 3710
rect 30075 3690 30095 3710
rect 30185 3690 30205 3710
rect 30295 3690 30315 3710
rect 30405 3690 30425 3710
rect 30515 3690 30535 3710
rect 30625 3690 30645 3710
rect 30020 3020 30040 3040
rect 30130 3020 30150 3040
rect 30186 3020 30204 3040
rect 30240 3020 30260 3040
rect 30350 3020 30370 3040
rect 30460 3020 30480 3040
rect 30570 3020 30590 3040
rect 31890 3650 31910 3660
rect 31890 3640 31910 3650
rect 31350 3580 31370 3600
rect 31470 3580 31490 3600
rect 31590 3580 31610 3600
rect 31710 3580 31730 3600
rect 31830 3580 31850 3600
rect 31890 3580 31910 3600
rect 31950 3580 31970 3600
rect 32070 3580 32090 3600
rect 32190 3580 32210 3600
rect 32310 3580 32330 3600
rect 32430 3580 32450 3600
rect 31290 3160 31310 3180
rect 31410 3160 31430 3180
rect 31530 3160 31550 3180
rect 31650 3160 31670 3180
rect 31770 3160 31790 3180
rect 31831 3160 31849 3180
rect 31890 3160 31910 3180
rect 32010 3160 32030 3180
rect 32130 3160 32150 3180
rect 32250 3160 32270 3180
rect 32370 3160 32390 3180
rect 32490 3160 32510 3180
rect 33155 3690 33175 3710
rect 33265 3690 33285 3710
rect 33375 3690 33395 3710
rect 33485 3690 33505 3710
rect 33595 3690 33615 3710
rect 33705 3690 33725 3710
rect 33815 3690 33835 3710
rect 30295 2970 30315 2980
rect 33210 3020 33230 3040
rect 33320 3020 33340 3040
rect 33430 3020 33450 3040
rect 33540 3020 33560 3040
rect 33596 3020 33614 3040
rect 33650 3020 33670 3040
rect 33760 3020 33780 3040
rect 33485 2970 33505 2980
rect 34111 3625 34141 3655
rect 34160 3625 34190 3655
rect 34210 3625 34240 3655
rect 34111 3020 34141 3050
rect 34160 3020 34190 3050
rect 34210 3020 34240 3050
rect 30295 2960 30315 2970
rect 33485 2960 33505 2970
rect 34245 2965 34265 2985
rect 30295 2800 30315 2810
rect 30295 2790 30315 2800
rect 29535 2669 29555 2679
rect 29535 2659 29555 2669
rect 30020 2730 30040 2750
rect 30130 2730 30150 2750
rect 30240 2730 30260 2750
rect 30350 2730 30370 2750
rect 30460 2730 30480 2750
rect 30570 2730 30590 2750
rect 30075 2460 30095 2480
rect 30185 2460 30205 2480
rect 30295 2460 30315 2480
rect 30405 2460 30425 2480
rect 30461 2460 30479 2480
rect 30515 2460 30535 2480
rect 31135 2870 31155 2890
rect 31255 2870 31275 2890
rect 31375 2870 31395 2890
rect 31495 2870 31515 2890
rect 31615 2870 31635 2890
rect 31075 2450 31095 2470
rect 31195 2450 31215 2470
rect 31315 2450 31335 2470
rect 31376 2450 31394 2470
rect 31435 2450 31455 2470
rect 31555 2450 31575 2470
rect 31675 2450 31695 2470
rect 32165 2870 32185 2890
rect 32285 2870 32305 2890
rect 32405 2870 32425 2890
rect 32525 2870 32545 2890
rect 32645 2870 32665 2890
rect 32105 2450 32125 2470
rect 32225 2450 32245 2470
rect 32345 2450 32365 2470
rect 32406 2450 32424 2470
rect 32465 2450 32485 2470
rect 32585 2450 32605 2470
rect 32705 2450 32725 2470
rect 33485 2800 33505 2810
rect 33485 2790 33505 2800
rect 33210 2730 33230 2750
rect 33320 2730 33340 2750
rect 33430 2730 33450 2750
rect 33540 2730 33560 2750
rect 33650 2730 33670 2750
rect 33760 2730 33780 2750
rect 33265 2460 33285 2480
rect 33321 2460 33339 2480
rect 33375 2460 33395 2480
rect 33485 2460 33505 2480
rect 33595 2460 33615 2480
rect 33705 2460 33725 2480
rect 34245 2669 34265 2679
rect 34245 2659 34265 2669
rect 29475 1955 29500 1980
rect 29535 1955 29560 1980
rect 29595 1955 29620 1980
rect 29655 1955 29680 1980
rect 29745 2085 29765 2105
rect 29895 2085 29905 2105
rect 29905 2085 29915 2105
rect 30075 2270 30095 2290
rect 30185 2270 30205 2290
rect 30295 2270 30315 2290
rect 30405 2270 30425 2290
rect 30461 2270 30479 2290
rect 30515 2270 30535 2290
rect 30020 1900 30038 1920
rect 30130 1900 30148 1920
rect 30240 1900 30258 1920
rect 30350 1900 30368 1920
rect 30460 1900 30478 1920
rect 30570 1900 30588 1920
rect 31250 2205 31270 2225
rect 31360 2205 31380 2225
rect 31470 2205 31490 2225
rect 31525 2205 31545 2225
rect 31580 2205 31600 2225
rect 31690 2205 31710 2225
rect 31800 2205 31820 2225
rect 31980 2205 32000 2225
rect 32090 2205 32110 2225
rect 32200 2205 32220 2225
rect 32255 2205 32275 2225
rect 32310 2205 32330 2225
rect 32420 2205 32440 2225
rect 32530 2205 32550 2225
rect 31305 1985 31325 2005
rect 31415 1985 31435 2005
rect 31525 1985 31545 2005
rect 31635 1985 31655 2005
rect 31745 1985 31765 2005
rect 32035 1985 32055 2005
rect 32145 1985 32165 2005
rect 32255 1985 32275 2005
rect 32365 1985 32385 2005
rect 32475 1985 32495 2005
rect 31890 1935 31910 1945
rect 31890 1925 31910 1935
rect 30295 1850 30315 1860
rect 33265 2270 33285 2290
rect 33321 2270 33339 2290
rect 33375 2270 33395 2290
rect 33485 2270 33505 2290
rect 33595 2270 33615 2290
rect 33705 2270 33725 2290
rect 33885 2085 33895 2105
rect 33895 2085 33905 2105
rect 34035 2085 34055 2105
rect 33212 1900 33230 1920
rect 33322 1900 33340 1920
rect 33432 1900 33450 1920
rect 33542 1900 33560 1920
rect 33652 1900 33670 1920
rect 33762 1900 33780 1920
rect 34120 1955 34145 1980
rect 34180 1955 34205 1980
rect 34240 1955 34265 1980
rect 34300 1955 34325 1980
rect 33485 1850 33505 1860
rect 30295 1840 30315 1850
rect 33485 1840 33505 1850
rect 31890 1805 31910 1815
rect 31890 1795 31910 1805
rect 30295 1740 30315 1760
rect 29735 1615 29760 1640
rect 29795 1615 29820 1640
rect 29885 1300 29905 1315
rect 29885 1295 29895 1300
rect 29895 1295 29905 1300
rect 29975 1295 29985 1315
rect 29985 1295 29995 1315
rect 30145 1680 30165 1700
rect 30345 1680 30365 1700
rect 30446 1680 30464 1700
rect 30545 1680 30565 1700
rect 31103 1725 31123 1745
rect 31197 1725 31217 1745
rect 31243 1735 31260 1755
rect 31323 1725 31343 1745
rect 31417 1725 31437 1745
rect 31463 1735 31480 1755
rect 31543 1725 31563 1745
rect 31610 1735 31627 1755
rect 31653 1725 31673 1745
rect 30950 1625 30960 1645
rect 30960 1625 30970 1645
rect 31827 1735 31847 1755
rect 31873 1735 31890 1755
rect 31950 1735 31970 1755
rect 32143 1725 32163 1745
rect 32237 1725 32257 1745
rect 32283 1735 32300 1755
rect 32363 1725 32383 1745
rect 32457 1725 32477 1745
rect 32503 1735 32520 1755
rect 32583 1725 32603 1745
rect 32650 1735 32667 1755
rect 32693 1725 32713 1745
rect 31112 1515 31129 1535
rect 31158 1515 31178 1535
rect 31260 1515 31280 1535
rect 31315 1515 31335 1535
rect 31370 1515 31390 1535
rect 31480 1515 31500 1535
rect 31535 1515 31555 1535
rect 31590 1515 31610 1535
rect 31830 1515 31850 1535
rect 31880 1515 31900 1535
rect 31928 1515 31945 1535
rect 32152 1515 32169 1535
rect 32198 1515 32218 1535
rect 32300 1515 32320 1535
rect 32355 1515 32375 1535
rect 32410 1515 32430 1535
rect 32520 1515 32540 1535
rect 32575 1515 32595 1535
rect 32630 1515 32650 1535
rect 33485 1740 33505 1760
rect 30245 910 30265 930
rect 30445 910 30465 930
rect 30345 860 30365 870
rect 31325 1230 31345 1250
rect 31435 1230 31455 1250
rect 31545 1230 31565 1250
rect 31655 1230 31675 1250
rect 31765 1230 31785 1250
rect 31820 1230 31840 1250
rect 31875 1230 31895 1250
rect 31985 1230 32005 1250
rect 32095 1230 32115 1250
rect 32205 1230 32225 1250
rect 32315 1230 32335 1250
rect 32386 1230 32406 1250
rect 32440 1230 32460 1250
rect 31205 910 31225 930
rect 31270 910 31290 930
rect 31380 910 31400 930
rect 31490 910 31510 930
rect 31600 910 31620 930
rect 31710 910 31730 930
rect 31820 910 31840 930
rect 31930 910 31950 930
rect 32040 910 32060 930
rect 32150 910 32170 930
rect 32260 910 32280 930
rect 32370 910 32390 930
rect 32485 910 32505 930
rect 30345 850 30365 860
rect 33235 1680 33255 1700
rect 33336 1680 33354 1700
rect 33435 1680 33455 1700
rect 33635 1680 33655 1700
rect 33980 1615 34005 1640
rect 34040 1615 34065 1640
rect 33805 1295 33815 1315
rect 33815 1295 33825 1315
rect 33895 1300 33915 1315
rect 33895 1295 33905 1300
rect 33905 1295 33915 1300
rect 33335 910 33355 930
rect 33535 910 33555 930
rect 33435 860 33455 870
rect 33435 850 33455 860
rect 31315 715 31335 735
rect 31385 715 31405 735
rect 31455 715 31475 735
rect 31515 715 31535 735
rect 31385 535 31405 545
rect 31945 710 31965 730
rect 32055 710 32075 730
rect 32165 710 32185 730
rect 32275 710 32295 730
rect 32385 710 32405 730
rect 32495 710 32515 730
rect 32000 590 32020 610
rect 32110 590 32130 610
rect 32220 590 32240 610
rect 32330 590 32350 610
rect 32440 590 32460 610
rect 32220 540 32240 550
rect 31385 525 31405 535
rect 32220 530 32240 540
<< metal1 >>
rect 30785 6185 30825 6190
rect 30785 6155 30790 6185
rect 30820 6155 30825 6185
rect 30785 6150 30825 6155
rect 30795 4875 30815 6150
rect 31530 4945 31570 4950
rect 31530 4915 31535 4945
rect 31565 4915 31570 4945
rect 31530 4910 31570 4915
rect 31650 4945 31690 4950
rect 31650 4915 31655 4945
rect 31685 4915 31690 4945
rect 31650 4910 31690 4915
rect 31770 4945 31810 4950
rect 31770 4915 31775 4945
rect 31805 4915 31810 4945
rect 31770 4910 31810 4915
rect 32440 4930 32480 4935
rect 31540 4890 31560 4910
rect 31660 4890 31680 4910
rect 31780 4890 31800 4910
rect 32440 4900 32445 4930
rect 32475 4900 32480 4930
rect 32440 4895 32480 4900
rect 31470 4885 31510 4890
rect 30785 4870 30825 4875
rect 30785 4840 30790 4870
rect 30820 4840 30825 4870
rect 30785 4835 30825 4840
rect 31280 4870 31320 4875
rect 31280 4840 31285 4870
rect 31315 4840 31320 4870
rect 31470 4855 31475 4885
rect 31505 4855 31510 4885
rect 31470 4850 31510 4855
rect 31537 4880 31563 4890
rect 31537 4860 31540 4880
rect 31560 4860 31563 4880
rect 31537 4850 31563 4860
rect 31590 4885 31630 4890
rect 31590 4855 31595 4885
rect 31625 4855 31630 4885
rect 31590 4850 31630 4855
rect 31657 4880 31683 4890
rect 31657 4860 31660 4880
rect 31680 4860 31683 4880
rect 31657 4850 31683 4860
rect 31710 4885 31750 4890
rect 31710 4855 31715 4885
rect 31745 4855 31750 4885
rect 31710 4850 31750 4855
rect 31777 4880 31803 4890
rect 31777 4860 31780 4880
rect 31800 4860 31803 4880
rect 31777 4850 31803 4860
rect 31830 4885 31870 4890
rect 31830 4855 31835 4885
rect 31865 4855 31870 4885
rect 32450 4865 32470 4895
rect 31830 4850 31870 4855
rect 32200 4860 32240 4865
rect 31280 4835 31320 4840
rect 30795 4445 30815 4835
rect 32200 4830 32205 4860
rect 32235 4830 32240 4860
rect 32200 4825 32240 4830
rect 32320 4860 32360 4865
rect 32320 4830 32325 4860
rect 32355 4830 32360 4860
rect 32320 4825 32360 4830
rect 32440 4860 32480 4865
rect 32440 4830 32445 4860
rect 32475 4830 32480 4860
rect 32440 4825 32480 4830
rect 32560 4860 32600 4865
rect 32560 4830 32565 4860
rect 32595 4830 32600 4860
rect 32560 4825 32600 4830
rect 32680 4860 32720 4865
rect 32680 4830 32685 4860
rect 32715 4830 32720 4860
rect 32680 4825 32720 4830
rect 31000 4730 31040 4735
rect 31000 4700 31005 4730
rect 31035 4700 31040 4730
rect 31310 4730 31350 4740
rect 31310 4710 31320 4730
rect 31340 4710 31350 4730
rect 31310 4700 31350 4710
rect 31650 4730 31690 4735
rect 31650 4700 31655 4730
rect 31685 4700 31690 4730
rect 31000 4695 31040 4700
rect 30785 4440 30825 4445
rect 30785 4410 30790 4440
rect 30820 4410 30825 4440
rect 30785 4405 30825 4410
rect 30795 3975 30815 4405
rect 30785 3970 30825 3975
rect 30785 3940 30790 3970
rect 30820 3940 30825 3970
rect 30785 3935 30825 3940
rect 29605 3735 29645 3740
rect 29605 3705 29610 3735
rect 29640 3705 29645 3735
rect 30795 3720 30815 3935
rect 29605 3700 29645 3705
rect 29955 3715 29995 3720
rect 29615 3660 29635 3700
rect 29955 3685 29960 3715
rect 29990 3685 29995 3715
rect 29955 3680 29995 3685
rect 30065 3715 30105 3720
rect 30065 3685 30070 3715
rect 30100 3685 30105 3715
rect 30065 3680 30105 3685
rect 30175 3715 30215 3720
rect 30175 3685 30180 3715
rect 30210 3685 30215 3715
rect 30175 3680 30215 3685
rect 30285 3715 30325 3720
rect 30285 3685 30290 3715
rect 30320 3685 30325 3715
rect 30285 3680 30325 3685
rect 30395 3715 30435 3720
rect 30395 3685 30400 3715
rect 30430 3685 30435 3715
rect 30395 3680 30435 3685
rect 30505 3715 30545 3720
rect 30505 3685 30510 3715
rect 30540 3685 30545 3715
rect 30505 3680 30545 3685
rect 30615 3715 30655 3720
rect 30615 3685 30620 3715
rect 30650 3685 30655 3715
rect 30615 3680 30655 3685
rect 30785 3715 30825 3720
rect 30785 3685 30790 3715
rect 30820 3685 30825 3715
rect 30785 3680 30825 3685
rect 29554 3655 29695 3660
rect 29554 3625 29560 3655
rect 29590 3625 29610 3655
rect 29640 3625 29659 3655
rect 29689 3625 29695 3655
rect 29554 3620 29695 3625
rect 29554 3050 29695 3055
rect 29554 3020 29560 3050
rect 29590 3020 29610 3050
rect 29640 3020 29659 3050
rect 29689 3020 29695 3050
rect 29554 3015 29695 3020
rect 30010 3045 30050 3050
rect 30010 3015 30015 3045
rect 30045 3015 30050 3045
rect 29525 2985 29565 2995
rect 29525 2965 29535 2985
rect 29555 2965 29565 2985
rect 29525 2955 29565 2965
rect 29315 2870 29355 2875
rect 29315 2840 29320 2870
rect 29350 2840 29355 2870
rect 29315 2835 29355 2840
rect 29265 2755 29305 2760
rect 29265 2725 29270 2755
rect 29300 2725 29305 2755
rect 29265 2720 29305 2725
rect 29275 500 29295 2720
rect 29325 2270 29345 2835
rect 29535 2689 29555 2955
rect 29615 2930 29635 3015
rect 30010 3010 30050 3015
rect 30120 3045 30160 3050
rect 30120 3015 30125 3045
rect 30155 3015 30160 3045
rect 30120 3010 30160 3015
rect 30178 3040 30212 3050
rect 30178 3020 30186 3040
rect 30204 3020 30212 3040
rect 30178 3010 30212 3020
rect 30230 3045 30270 3050
rect 30230 3015 30235 3045
rect 30265 3015 30270 3045
rect 30230 3010 30270 3015
rect 30340 3045 30380 3050
rect 30340 3015 30345 3045
rect 30375 3015 30380 3045
rect 30340 3010 30380 3015
rect 30450 3045 30490 3050
rect 30450 3015 30455 3045
rect 30485 3015 30490 3045
rect 30450 3010 30490 3015
rect 30560 3045 30600 3050
rect 30560 3015 30565 3045
rect 30595 3015 30600 3045
rect 30560 3010 30600 3015
rect 30185 2930 30205 3010
rect 30285 2980 30325 2990
rect 30285 2960 30295 2980
rect 30315 2960 30325 2980
rect 30285 2950 30325 2960
rect 29605 2925 29645 2930
rect 29605 2895 29610 2925
rect 29640 2895 29645 2925
rect 29605 2890 29645 2895
rect 30175 2925 30215 2930
rect 30175 2895 30180 2925
rect 30210 2895 30215 2925
rect 30175 2890 30215 2895
rect 30295 2820 30315 2950
rect 30460 2875 30480 3010
rect 30740 2925 30780 2930
rect 30740 2895 30745 2925
rect 30775 2895 30780 2925
rect 30740 2890 30780 2895
rect 30450 2870 30490 2875
rect 30450 2840 30455 2870
rect 30485 2840 30490 2870
rect 30450 2835 30490 2840
rect 30285 2810 30325 2820
rect 30285 2790 30295 2810
rect 30315 2790 30325 2810
rect 30285 2780 30325 2790
rect 30010 2755 30050 2760
rect 30010 2725 30015 2755
rect 30045 2725 30050 2755
rect 30010 2720 30050 2725
rect 30120 2755 30160 2760
rect 30120 2725 30125 2755
rect 30155 2725 30160 2755
rect 30120 2720 30160 2725
rect 30230 2755 30270 2760
rect 30230 2725 30235 2755
rect 30265 2725 30270 2755
rect 30230 2720 30270 2725
rect 30340 2755 30380 2760
rect 30340 2725 30345 2755
rect 30375 2725 30380 2755
rect 30340 2720 30380 2725
rect 30450 2755 30490 2760
rect 30450 2725 30455 2755
rect 30485 2725 30490 2755
rect 30450 2720 30490 2725
rect 30560 2755 30600 2760
rect 30560 2725 30565 2755
rect 30595 2725 30600 2755
rect 30560 2720 30600 2725
rect 29525 2679 29565 2689
rect 29525 2659 29535 2679
rect 29555 2659 29565 2679
rect 29525 2649 29565 2659
rect 29790 2485 29830 2490
rect 29790 2455 29795 2485
rect 29825 2455 29830 2485
rect 29790 2450 29830 2455
rect 30065 2485 30105 2490
rect 30065 2455 30070 2485
rect 30100 2455 30105 2485
rect 30065 2450 30105 2455
rect 30175 2485 30215 2490
rect 30175 2455 30180 2485
rect 30210 2455 30215 2485
rect 30175 2450 30215 2455
rect 30285 2485 30325 2490
rect 30285 2455 30290 2485
rect 30320 2455 30325 2485
rect 30285 2450 30325 2455
rect 30395 2485 30435 2490
rect 30395 2455 30400 2485
rect 30430 2455 30435 2485
rect 30395 2450 30435 2455
rect 30453 2480 30487 2490
rect 30453 2460 30461 2480
rect 30479 2460 30487 2480
rect 30453 2450 30487 2460
rect 30505 2485 30545 2490
rect 30505 2455 30510 2485
rect 30540 2455 30545 2485
rect 30505 2450 30545 2455
rect 29310 2260 29360 2270
rect 29310 2230 29320 2260
rect 29350 2230 29360 2260
rect 29310 2220 29360 2230
rect 29325 1710 29345 2220
rect 29735 2110 29775 2115
rect 29735 2080 29740 2110
rect 29770 2080 29775 2110
rect 29735 2075 29775 2080
rect 29470 1985 29505 1990
rect 29470 1945 29505 1950
rect 29530 1985 29565 1990
rect 29530 1945 29565 1950
rect 29590 1985 29625 1991
rect 29590 1945 29625 1950
rect 29650 1985 29685 1990
rect 29800 1985 29820 2450
rect 30460 2380 30480 2450
rect 30750 2380 30770 2890
rect 30450 2375 30490 2380
rect 30450 2345 30455 2375
rect 30485 2345 30490 2375
rect 30450 2340 30490 2345
rect 30740 2375 30780 2380
rect 30740 2345 30745 2375
rect 30775 2345 30780 2375
rect 30740 2340 30780 2345
rect 30460 2300 30480 2340
rect 29835 2295 29875 2300
rect 29835 2265 29840 2295
rect 29870 2265 29875 2295
rect 29835 2260 29875 2265
rect 30065 2295 30105 2300
rect 30065 2265 30070 2295
rect 30100 2265 30105 2295
rect 30065 2260 30105 2265
rect 30175 2295 30215 2300
rect 30175 2265 30180 2295
rect 30210 2265 30215 2295
rect 30175 2260 30215 2265
rect 30285 2295 30325 2300
rect 30285 2265 30290 2295
rect 30320 2265 30325 2295
rect 30285 2260 30325 2265
rect 30395 2295 30435 2300
rect 30395 2265 30400 2295
rect 30430 2265 30435 2295
rect 30395 2260 30435 2265
rect 30453 2290 30487 2300
rect 30453 2270 30461 2290
rect 30479 2270 30487 2290
rect 30453 2260 30487 2270
rect 30505 2295 30545 2300
rect 30505 2265 30510 2295
rect 30540 2265 30545 2295
rect 30505 2260 30545 2265
rect 29650 1945 29685 1950
rect 29790 1980 29830 1985
rect 29790 1950 29795 1980
rect 29825 1950 29830 1980
rect 29790 1945 29830 1950
rect 29480 1825 29500 1945
rect 29600 1930 29620 1945
rect 29845 1930 29865 2260
rect 29885 2110 29925 2115
rect 29885 2080 29890 2110
rect 29920 2080 29925 2110
rect 29885 2075 29925 2080
rect 30795 1930 30815 3680
rect 31010 3190 31030 4695
rect 31320 4550 31340 4700
rect 31650 4695 31690 4700
rect 32260 4730 32300 4735
rect 32260 4700 32265 4730
rect 32295 4700 32300 4730
rect 32260 4695 32300 4700
rect 32323 4725 32357 4735
rect 32323 4705 32331 4725
rect 32349 4705 32357 4725
rect 32323 4695 32357 4705
rect 32380 4730 32420 4735
rect 32380 4700 32385 4730
rect 32415 4700 32420 4730
rect 32380 4695 32420 4700
rect 32500 4730 32540 4735
rect 32500 4700 32505 4730
rect 32535 4700 32540 4730
rect 32500 4695 32540 4700
rect 32620 4730 32660 4735
rect 32620 4700 32625 4730
rect 32655 4700 32660 4730
rect 32620 4695 32660 4700
rect 32330 4550 32350 4695
rect 31055 4545 31095 4550
rect 31055 4515 31060 4545
rect 31090 4515 31095 4545
rect 31055 4510 31095 4515
rect 31310 4545 31350 4550
rect 31310 4515 31315 4545
rect 31345 4515 31350 4545
rect 31310 4510 31350 4515
rect 32320 4545 32360 4550
rect 32320 4515 32325 4545
rect 32355 4515 32360 4545
rect 32320 4510 32360 4515
rect 31000 3185 31040 3190
rect 31000 3155 31005 3185
rect 31035 3155 31040 3185
rect 31000 3150 31040 3155
rect 31065 2995 31085 4510
rect 31250 4440 31290 4445
rect 31250 4410 31255 4440
rect 31285 4410 31290 4440
rect 31250 4405 31290 4410
rect 31360 4440 31400 4445
rect 31360 4410 31365 4440
rect 31395 4410 31400 4440
rect 31360 4405 31400 4410
rect 31470 4440 31510 4445
rect 31470 4410 31475 4440
rect 31505 4410 31510 4440
rect 31470 4405 31510 4410
rect 31580 4440 31620 4445
rect 31580 4410 31585 4440
rect 31615 4410 31620 4440
rect 31580 4405 31620 4410
rect 31690 4440 31730 4445
rect 31690 4410 31695 4440
rect 31725 4410 31730 4440
rect 31690 4405 31730 4410
rect 31800 4440 31840 4445
rect 31800 4410 31805 4440
rect 31835 4410 31840 4440
rect 31800 4405 31840 4410
rect 31910 4440 31950 4445
rect 31910 4410 31915 4440
rect 31945 4410 31950 4440
rect 31910 4405 31950 4410
rect 32020 4440 32060 4445
rect 32020 4410 32025 4440
rect 32055 4410 32060 4440
rect 32020 4405 32060 4410
rect 32130 4440 32170 4445
rect 32130 4410 32135 4440
rect 32165 4410 32170 4440
rect 32130 4405 32170 4410
rect 32240 4440 32280 4445
rect 32240 4410 32245 4440
rect 32275 4410 32280 4440
rect 32240 4405 32280 4410
rect 32350 4440 32390 4445
rect 32350 4410 32355 4440
rect 32385 4410 32390 4440
rect 32350 4405 32390 4410
rect 32460 4440 32500 4445
rect 32460 4410 32465 4440
rect 32495 4410 32500 4440
rect 32460 4405 32500 4410
rect 31305 4320 31345 4325
rect 31305 4290 31310 4320
rect 31340 4290 31345 4320
rect 31305 4285 31345 4290
rect 31362 4315 31398 4325
rect 31362 4295 31370 4315
rect 31390 4295 31398 4315
rect 31362 4285 31398 4295
rect 31415 4315 31455 4325
rect 31415 4295 31425 4315
rect 31445 4295 31455 4315
rect 31415 4285 31455 4295
rect 31525 4320 31565 4325
rect 31525 4290 31530 4320
rect 31560 4290 31565 4320
rect 31525 4285 31565 4290
rect 31635 4315 31675 4325
rect 31635 4295 31645 4315
rect 31665 4295 31675 4315
rect 31635 4285 31675 4295
rect 31745 4320 31785 4325
rect 31745 4290 31750 4320
rect 31780 4290 31785 4320
rect 31745 4285 31785 4290
rect 31855 4315 31895 4325
rect 31855 4295 31865 4315
rect 31885 4295 31895 4315
rect 31855 4285 31895 4295
rect 31965 4320 32005 4325
rect 31965 4290 31970 4320
rect 32000 4290 32005 4320
rect 31965 4285 32005 4290
rect 32075 4315 32115 4325
rect 32075 4295 32085 4315
rect 32105 4295 32115 4315
rect 32075 4285 32115 4295
rect 32185 4320 32225 4325
rect 32185 4290 32190 4320
rect 32220 4290 32225 4320
rect 32185 4285 32225 4290
rect 32295 4315 32335 4325
rect 32295 4295 32305 4315
rect 32325 4295 32335 4315
rect 32295 4285 32335 4295
rect 32390 4320 32445 4325
rect 32390 4290 32410 4320
rect 32440 4290 32445 4320
rect 32390 4285 32445 4290
rect 31320 4090 31360 4095
rect 31320 4060 31325 4090
rect 31355 4060 31360 4090
rect 31320 4055 31360 4060
rect 31330 4035 31350 4055
rect 31375 4035 31395 4285
rect 31430 4210 31450 4285
rect 31645 4210 31665 4285
rect 31865 4210 31885 4285
rect 32085 4210 32105 4285
rect 32305 4210 32325 4285
rect 31420 4205 31460 4210
rect 31420 4175 31425 4205
rect 31455 4175 31460 4205
rect 31420 4170 31460 4175
rect 31635 4205 31675 4210
rect 31635 4175 31640 4205
rect 31670 4175 31675 4205
rect 31635 4170 31675 4175
rect 31855 4205 31895 4210
rect 31855 4175 31860 4205
rect 31890 4175 31895 4205
rect 31855 4170 31895 4175
rect 32075 4205 32115 4210
rect 32075 4175 32080 4205
rect 32110 4175 32115 4205
rect 32075 4170 32115 4175
rect 32295 4205 32335 4210
rect 32295 4175 32300 4205
rect 32330 4175 32335 4205
rect 32295 4170 32335 4175
rect 31430 4095 31450 4170
rect 32390 4095 32410 4285
rect 31420 4090 31460 4095
rect 31420 4060 31425 4090
rect 31455 4060 31460 4090
rect 31420 4055 31460 4060
rect 31530 4090 31570 4095
rect 31530 4060 31535 4090
rect 31565 4060 31570 4090
rect 31530 4055 31570 4060
rect 31640 4090 31680 4095
rect 31640 4060 31645 4090
rect 31675 4060 31680 4090
rect 31640 4055 31680 4060
rect 31750 4090 31790 4095
rect 31750 4060 31755 4090
rect 31785 4060 31790 4090
rect 31750 4055 31790 4060
rect 32050 4090 32090 4095
rect 32050 4060 32055 4090
rect 32085 4060 32090 4090
rect 32050 4055 32090 4060
rect 32150 4090 32190 4095
rect 32150 4060 32155 4090
rect 32185 4060 32190 4090
rect 32150 4055 32190 4060
rect 32260 4090 32300 4095
rect 32260 4060 32265 4090
rect 32295 4060 32300 4090
rect 32260 4055 32300 4060
rect 32370 4090 32410 4095
rect 32370 4060 32375 4090
rect 32405 4060 32410 4090
rect 32370 4055 32410 4060
rect 32480 4090 32520 4095
rect 32480 4060 32485 4090
rect 32515 4060 32520 4090
rect 32480 4055 32520 4060
rect 31430 4035 31450 4055
rect 31540 4035 31560 4055
rect 31650 4035 31670 4055
rect 31760 4035 31780 4055
rect 32060 4035 32080 4055
rect 32160 4035 32180 4055
rect 32270 4035 32290 4055
rect 32380 4035 32400 4055
rect 32490 4035 32510 4055
rect 31280 4029 31310 4035
rect 31280 4001 31282 4029
rect 31308 4001 31310 4029
rect 31280 3995 31310 4001
rect 31327 4025 31353 4035
rect 31327 4005 31330 4025
rect 31350 4005 31353 4025
rect 31327 3995 31353 4005
rect 31370 4025 31400 4035
rect 31370 4005 31375 4025
rect 31395 4005 31400 4025
rect 31370 3995 31400 4005
rect 31427 4025 31453 4035
rect 31427 4005 31430 4025
rect 31450 4005 31453 4025
rect 31427 3995 31453 4005
rect 31480 4029 31510 4035
rect 31480 4001 31482 4029
rect 31508 4001 31510 4029
rect 31480 3995 31510 4001
rect 31537 4025 31563 4035
rect 31537 4005 31540 4025
rect 31560 4005 31563 4025
rect 31537 3995 31563 4005
rect 31647 4025 31673 4035
rect 31647 4005 31650 4025
rect 31670 4005 31673 4025
rect 31647 3995 31673 4005
rect 31695 4030 31735 4035
rect 31695 4000 31700 4030
rect 31730 4000 31735 4030
rect 31695 3995 31735 4000
rect 31757 4025 31783 4035
rect 31757 4005 31760 4025
rect 31780 4005 31783 4025
rect 31757 3995 31783 4005
rect 32008 4029 32038 4035
rect 32008 4001 32010 4029
rect 32036 4001 32038 4029
rect 32008 3995 32038 4001
rect 32057 4025 32083 4035
rect 32057 4005 32060 4025
rect 32080 4005 32083 4025
rect 32057 3995 32083 4005
rect 32157 4025 32183 4035
rect 32157 4005 32160 4025
rect 32180 4005 32183 4025
rect 32157 3995 32183 4005
rect 32205 4030 32245 4035
rect 32205 4000 32210 4030
rect 32240 4000 32245 4030
rect 32205 3995 32245 4000
rect 32267 4025 32293 4035
rect 32267 4005 32270 4025
rect 32290 4005 32293 4025
rect 32267 3995 32293 4005
rect 32377 4025 32403 4035
rect 32377 4005 32380 4025
rect 32400 4005 32403 4025
rect 32377 3995 32403 4005
rect 32425 4030 32465 4035
rect 32425 4000 32430 4030
rect 32460 4000 32465 4030
rect 32425 3995 32465 4000
rect 32487 4025 32513 4035
rect 32487 4005 32490 4025
rect 32510 4005 32513 4025
rect 32487 3995 32513 4005
rect 32870 4030 32910 4035
rect 32870 4000 32875 4030
rect 32905 4000 32910 4030
rect 32870 3995 32910 4000
rect 31140 3970 31180 3975
rect 31140 3940 31145 3970
rect 31175 3940 31180 3970
rect 31140 3935 31180 3940
rect 31255 3905 31295 3915
rect 31255 3885 31265 3905
rect 31285 3885 31295 3905
rect 31255 3875 31295 3885
rect 31350 3905 31390 3915
rect 31350 3885 31360 3905
rect 31380 3885 31390 3905
rect 31350 3875 31390 3885
rect 31407 3910 31439 3915
rect 31407 3880 31410 3910
rect 31436 3880 31439 3910
rect 31407 3875 31439 3880
rect 31475 3905 31515 3915
rect 31475 3885 31485 3905
rect 31505 3885 31515 3905
rect 31475 3875 31515 3885
rect 31570 3905 31610 3915
rect 31570 3885 31580 3905
rect 31600 3885 31610 3905
rect 31570 3875 31610 3885
rect 31627 3910 31659 3915
rect 31627 3880 31630 3910
rect 31656 3880 31659 3910
rect 31627 3875 31659 3880
rect 31695 3905 31735 3915
rect 31695 3885 31705 3905
rect 31725 3885 31735 3905
rect 31695 3875 31735 3885
rect 31771 3910 31803 3915
rect 31771 3880 31774 3910
rect 31800 3880 31803 3910
rect 31771 3875 31803 3880
rect 31820 3905 31846 3915
rect 31820 3885 31823 3905
rect 31843 3885 31846 3905
rect 31820 3875 31846 3885
rect 31985 3905 32025 3915
rect 31985 3885 31995 3905
rect 32015 3885 32025 3905
rect 31985 3875 32025 3885
rect 32080 3905 32120 3915
rect 32080 3885 32090 3905
rect 32110 3885 32120 3905
rect 32080 3875 32120 3885
rect 32137 3910 32169 3915
rect 32137 3880 32140 3910
rect 32166 3880 32169 3910
rect 32137 3875 32169 3880
rect 32205 3905 32245 3915
rect 32205 3885 32215 3905
rect 32235 3885 32245 3905
rect 32205 3875 32245 3885
rect 32300 3905 32340 3915
rect 32300 3885 32310 3905
rect 32330 3885 32340 3905
rect 32300 3875 32340 3885
rect 32357 3910 32389 3915
rect 32357 3880 32360 3910
rect 32386 3880 32389 3910
rect 32357 3875 32389 3880
rect 32425 3905 32465 3915
rect 32425 3885 32435 3905
rect 32455 3885 32465 3905
rect 32425 3875 32465 3885
rect 32501 3910 32533 3915
rect 32501 3880 32504 3910
rect 32530 3880 32533 3910
rect 32501 3875 32533 3880
rect 32550 3905 32576 3915
rect 32550 3885 32553 3905
rect 32573 3885 32576 3905
rect 32550 3875 32576 3885
rect 31265 3855 31285 3875
rect 31370 3855 31390 3875
rect 31485 3855 31505 3875
rect 31590 3855 31610 3875
rect 31705 3855 31725 3875
rect 31820 3855 31840 3875
rect 31995 3855 32015 3875
rect 31255 3850 31295 3855
rect 31255 3820 31260 3850
rect 31290 3820 31295 3850
rect 31255 3815 31295 3820
rect 31360 3850 31400 3855
rect 31360 3820 31365 3850
rect 31395 3820 31400 3850
rect 31360 3815 31400 3820
rect 31475 3850 31515 3855
rect 31475 3820 31480 3850
rect 31510 3820 31515 3850
rect 31475 3815 31515 3820
rect 31580 3850 31620 3855
rect 31580 3820 31585 3850
rect 31615 3820 31620 3850
rect 31580 3815 31620 3820
rect 31695 3850 31735 3855
rect 31695 3820 31700 3850
rect 31730 3820 31735 3850
rect 31695 3815 31735 3820
rect 31810 3850 31850 3855
rect 31810 3820 31815 3850
rect 31845 3820 31850 3850
rect 31810 3815 31850 3820
rect 31985 3850 32025 3855
rect 31985 3820 31990 3850
rect 32020 3820 32025 3850
rect 31985 3815 32025 3820
rect 32090 3765 32110 3875
rect 32215 3855 32235 3875
rect 32205 3850 32245 3855
rect 32205 3820 32210 3850
rect 32240 3820 32245 3850
rect 32205 3815 32245 3820
rect 32310 3765 32330 3875
rect 32435 3855 32455 3875
rect 32425 3850 32465 3855
rect 32425 3820 32430 3850
rect 32460 3820 32465 3850
rect 32425 3815 32465 3820
rect 32550 3765 32570 3875
rect 32080 3760 32120 3765
rect 32080 3730 32085 3760
rect 32115 3730 32120 3760
rect 31880 3725 31920 3730
rect 32080 3725 32120 3730
rect 32300 3760 32340 3765
rect 32300 3730 32305 3760
rect 32335 3730 32340 3760
rect 32300 3725 32340 3730
rect 32540 3760 32580 3765
rect 32540 3730 32545 3760
rect 32575 3730 32580 3760
rect 32540 3725 32580 3730
rect 31880 3695 31885 3725
rect 31915 3695 31920 3725
rect 31880 3690 31920 3695
rect 31890 3670 31910 3690
rect 31880 3665 31920 3670
rect 31880 3635 31885 3665
rect 31915 3635 31920 3665
rect 31880 3630 31920 3635
rect 31890 3610 31910 3630
rect 31340 3605 31380 3610
rect 31340 3575 31345 3605
rect 31375 3575 31380 3605
rect 31340 3570 31380 3575
rect 31460 3605 31500 3610
rect 31460 3575 31465 3605
rect 31495 3575 31500 3605
rect 31460 3570 31500 3575
rect 31580 3605 31620 3610
rect 31580 3575 31585 3605
rect 31615 3575 31620 3605
rect 31580 3570 31620 3575
rect 31700 3605 31740 3610
rect 31700 3575 31705 3605
rect 31735 3575 31740 3605
rect 31700 3570 31740 3575
rect 31820 3605 31860 3610
rect 31820 3575 31825 3605
rect 31855 3575 31860 3605
rect 31820 3570 31860 3575
rect 31880 3605 31920 3610
rect 31880 3575 31885 3605
rect 31915 3575 31920 3605
rect 31880 3570 31920 3575
rect 31940 3605 31980 3610
rect 31940 3575 31945 3605
rect 31975 3575 31980 3605
rect 31940 3570 31980 3575
rect 32060 3605 32100 3610
rect 32060 3575 32065 3605
rect 32095 3575 32100 3605
rect 32060 3570 32100 3575
rect 32180 3605 32220 3610
rect 32180 3575 32185 3605
rect 32215 3575 32220 3605
rect 32180 3570 32220 3575
rect 32300 3605 32340 3610
rect 32300 3575 32305 3605
rect 32335 3575 32340 3605
rect 32300 3570 32340 3575
rect 32420 3605 32460 3610
rect 32420 3575 32425 3605
rect 32455 3575 32460 3605
rect 32420 3570 32460 3575
rect 31280 3180 31320 3190
rect 31280 3160 31290 3180
rect 31310 3160 31320 3180
rect 31280 3150 31320 3160
rect 31400 3180 31440 3190
rect 31400 3160 31410 3180
rect 31430 3160 31440 3180
rect 31400 3150 31440 3160
rect 31520 3180 31560 3190
rect 31520 3160 31530 3180
rect 31550 3160 31560 3180
rect 31520 3150 31560 3160
rect 31640 3180 31680 3190
rect 31640 3160 31650 3180
rect 31670 3160 31680 3180
rect 31640 3150 31680 3160
rect 31760 3180 31800 3190
rect 31760 3160 31770 3180
rect 31790 3160 31800 3180
rect 31760 3150 31800 3160
rect 31823 3185 31857 3190
rect 31823 3155 31826 3185
rect 31854 3155 31857 3185
rect 31823 3150 31857 3155
rect 31880 3180 31920 3190
rect 31880 3160 31890 3180
rect 31910 3160 31920 3180
rect 31880 3150 31920 3160
rect 32000 3180 32040 3190
rect 32000 3160 32010 3180
rect 32030 3160 32040 3180
rect 32000 3150 32040 3160
rect 32120 3180 32160 3190
rect 32120 3160 32130 3180
rect 32150 3160 32160 3180
rect 32120 3150 32160 3160
rect 32240 3180 32280 3190
rect 32240 3160 32250 3180
rect 32270 3160 32280 3180
rect 32240 3150 32280 3160
rect 32360 3180 32400 3190
rect 32360 3160 32370 3180
rect 32390 3160 32400 3180
rect 32360 3150 32400 3160
rect 32480 3180 32520 3190
rect 32480 3160 32490 3180
rect 32510 3160 32520 3180
rect 32480 3150 32520 3160
rect 31290 3135 31310 3150
rect 31260 3130 31320 3135
rect 31260 3100 31285 3130
rect 31315 3100 31320 3130
rect 31260 3095 31320 3100
rect 31055 2990 31095 2995
rect 31055 2960 31060 2990
rect 31090 2960 31095 2990
rect 31055 2955 31095 2960
rect 31260 2900 31280 3095
rect 31410 3050 31430 3150
rect 31530 3135 31550 3150
rect 31520 3130 31560 3135
rect 31520 3100 31525 3130
rect 31555 3100 31560 3130
rect 31520 3095 31560 3100
rect 31650 3050 31670 3150
rect 31770 3135 31790 3150
rect 31760 3130 31800 3135
rect 31760 3100 31765 3130
rect 31795 3100 31800 3130
rect 31760 3095 31800 3100
rect 31890 3050 31910 3150
rect 32010 3135 32030 3150
rect 32000 3130 32040 3135
rect 32000 3100 32005 3130
rect 32035 3100 32040 3130
rect 32000 3095 32040 3100
rect 32130 3050 32150 3150
rect 32250 3135 32270 3150
rect 32240 3130 32280 3135
rect 32240 3100 32245 3130
rect 32275 3100 32280 3130
rect 32240 3095 32280 3100
rect 32370 3050 32390 3150
rect 32490 3135 32510 3150
rect 32480 3130 32520 3135
rect 32480 3100 32485 3130
rect 32515 3100 32520 3130
rect 32480 3095 32520 3100
rect 31400 3045 31440 3050
rect 31400 3015 31405 3045
rect 31435 3015 31440 3045
rect 31400 3010 31440 3015
rect 31640 3045 31680 3050
rect 31640 3015 31645 3045
rect 31675 3015 31680 3045
rect 31640 3010 31680 3015
rect 31880 3045 31920 3050
rect 31880 3015 31885 3045
rect 31915 3015 31920 3045
rect 31880 3010 31920 3015
rect 32120 3045 32160 3050
rect 32120 3015 32125 3045
rect 32155 3015 32160 3045
rect 32120 3010 32160 3015
rect 32360 3045 32415 3050
rect 32360 3015 32365 3045
rect 32395 3015 32415 3045
rect 32360 3010 32415 3015
rect 31880 2990 31920 2995
rect 31880 2960 31885 2990
rect 31915 2960 31920 2990
rect 31880 2955 31920 2960
rect 31125 2895 31165 2900
rect 31125 2865 31130 2895
rect 31160 2865 31165 2895
rect 31125 2860 31165 2865
rect 31245 2895 31285 2900
rect 31245 2865 31250 2895
rect 31280 2865 31285 2895
rect 31245 2860 31285 2865
rect 31365 2895 31405 2900
rect 31365 2865 31370 2895
rect 31400 2865 31405 2895
rect 31365 2860 31405 2865
rect 31485 2895 31525 2900
rect 31485 2865 31490 2895
rect 31520 2865 31525 2895
rect 31485 2860 31525 2865
rect 31605 2895 31645 2900
rect 31605 2865 31610 2895
rect 31640 2865 31645 2895
rect 31605 2860 31645 2865
rect 31065 2475 31105 2480
rect 31065 2445 31070 2475
rect 31100 2445 31105 2475
rect 31065 2440 31105 2445
rect 31185 2475 31225 2480
rect 31185 2445 31190 2475
rect 31220 2445 31225 2475
rect 31185 2440 31225 2445
rect 31305 2475 31345 2480
rect 31305 2445 31310 2475
rect 31340 2445 31345 2475
rect 31305 2440 31345 2445
rect 31368 2470 31402 2480
rect 31368 2450 31376 2470
rect 31394 2450 31402 2470
rect 31368 2440 31402 2450
rect 31425 2475 31465 2480
rect 31425 2445 31430 2475
rect 31460 2445 31465 2475
rect 31425 2440 31465 2445
rect 31545 2475 31585 2480
rect 31545 2445 31550 2475
rect 31580 2445 31585 2475
rect 31545 2440 31585 2445
rect 31665 2475 31705 2480
rect 31665 2445 31670 2475
rect 31700 2445 31705 2475
rect 31665 2440 31705 2445
rect 31375 2425 31395 2440
rect 31365 2420 31405 2425
rect 31365 2390 31370 2420
rect 31400 2390 31405 2420
rect 31365 2385 31405 2390
rect 31680 2380 31700 2440
rect 31890 2425 31910 2955
rect 32395 2900 32415 3010
rect 32155 2895 32195 2900
rect 32155 2865 32160 2895
rect 32190 2865 32195 2895
rect 32155 2860 32195 2865
rect 32275 2895 32315 2900
rect 32275 2865 32280 2895
rect 32310 2865 32315 2895
rect 32275 2860 32315 2865
rect 32395 2895 32435 2900
rect 32395 2865 32400 2895
rect 32430 2865 32435 2895
rect 32395 2860 32435 2865
rect 32515 2895 32555 2900
rect 32515 2865 32520 2895
rect 32550 2865 32555 2895
rect 32515 2860 32555 2865
rect 32635 2895 32675 2900
rect 32635 2865 32640 2895
rect 32670 2865 32675 2895
rect 32635 2860 32675 2865
rect 32095 2475 32135 2480
rect 32095 2445 32100 2475
rect 32130 2445 32135 2475
rect 32095 2440 32135 2445
rect 32215 2475 32255 2480
rect 32215 2445 32220 2475
rect 32250 2445 32255 2475
rect 32215 2440 32255 2445
rect 32335 2475 32375 2480
rect 32335 2445 32340 2475
rect 32370 2445 32375 2475
rect 32335 2440 32375 2445
rect 32398 2470 32432 2480
rect 32398 2450 32406 2470
rect 32424 2450 32432 2470
rect 32398 2440 32432 2450
rect 32455 2475 32495 2480
rect 32455 2445 32460 2475
rect 32490 2445 32495 2475
rect 32455 2440 32495 2445
rect 32575 2475 32615 2480
rect 32575 2445 32580 2475
rect 32610 2445 32615 2475
rect 32575 2440 32615 2445
rect 32695 2475 32735 2480
rect 32695 2445 32700 2475
rect 32730 2445 32735 2475
rect 32695 2440 32735 2445
rect 31880 2420 31920 2425
rect 31880 2390 31885 2420
rect 31915 2390 31920 2420
rect 31880 2385 31920 2390
rect 32100 2380 32120 2440
rect 32405 2425 32425 2440
rect 32395 2420 32435 2425
rect 32395 2390 32400 2420
rect 32430 2390 32435 2420
rect 32395 2385 32435 2390
rect 31670 2375 31710 2380
rect 31670 2345 31675 2375
rect 31705 2345 31710 2375
rect 31670 2340 31710 2345
rect 32090 2375 32130 2380
rect 32090 2345 32095 2375
rect 32125 2345 32130 2375
rect 32090 2340 32130 2345
rect 30875 2330 30915 2335
rect 30875 2300 30880 2330
rect 30910 2300 30915 2330
rect 30875 2295 30915 2300
rect 30830 2230 30870 2235
rect 30830 2200 30835 2230
rect 30865 2200 30870 2230
rect 30830 2195 30870 2200
rect 29590 1925 29630 1930
rect 29590 1895 29595 1925
rect 29625 1895 29630 1925
rect 29590 1890 29630 1895
rect 29835 1925 29875 1930
rect 29835 1895 29840 1925
rect 29870 1895 29875 1925
rect 29835 1890 29875 1895
rect 30010 1925 30050 1930
rect 30010 1895 30015 1925
rect 30045 1895 30050 1925
rect 30010 1890 30050 1895
rect 30120 1925 30160 1930
rect 30120 1895 30125 1925
rect 30155 1895 30160 1925
rect 30120 1890 30160 1895
rect 30230 1925 30270 1930
rect 30230 1895 30235 1925
rect 30265 1895 30270 1925
rect 30230 1890 30270 1895
rect 30340 1925 30380 1930
rect 30340 1895 30345 1925
rect 30375 1895 30380 1925
rect 30340 1890 30380 1895
rect 30450 1925 30490 1930
rect 30450 1895 30455 1925
rect 30485 1895 30490 1925
rect 30450 1890 30490 1895
rect 30560 1925 30600 1930
rect 30560 1895 30565 1925
rect 30595 1895 30600 1925
rect 30560 1890 30600 1895
rect 30785 1925 30825 1930
rect 30785 1895 30790 1925
rect 30820 1895 30825 1925
rect 30785 1890 30825 1895
rect 30285 1860 30325 1870
rect 30285 1840 30295 1860
rect 30315 1840 30325 1860
rect 30285 1830 30325 1840
rect 29470 1820 29510 1825
rect 29470 1790 29475 1820
rect 29505 1790 29510 1820
rect 29470 1785 29510 1790
rect 30295 1770 30315 1830
rect 29725 1760 29765 1765
rect 29725 1730 29730 1760
rect 29760 1730 29765 1760
rect 30285 1760 30325 1770
rect 30285 1740 30295 1760
rect 30315 1740 30325 1760
rect 30285 1730 30325 1740
rect 30435 1760 30475 1765
rect 30435 1730 30440 1760
rect 30470 1730 30475 1760
rect 29725 1725 29765 1730
rect 30435 1725 30475 1730
rect 30740 1760 30780 1765
rect 30740 1730 30745 1760
rect 30775 1730 30780 1760
rect 30740 1725 30780 1730
rect 29315 1705 29355 1710
rect 29315 1675 29320 1705
rect 29350 1675 29355 1705
rect 29315 1670 29355 1675
rect 29735 1650 29755 1725
rect 30445 1710 30465 1725
rect 29790 1705 29830 1710
rect 29790 1675 29795 1705
rect 29825 1675 29830 1705
rect 29790 1670 29830 1675
rect 30135 1705 30175 1710
rect 30135 1675 30140 1705
rect 30170 1675 30175 1705
rect 30135 1670 30175 1675
rect 30335 1705 30375 1710
rect 30335 1675 30340 1705
rect 30370 1675 30375 1705
rect 30335 1670 30375 1675
rect 30438 1700 30472 1710
rect 30438 1680 30446 1700
rect 30464 1680 30472 1700
rect 30438 1670 30472 1680
rect 30535 1705 30575 1710
rect 30535 1675 30540 1705
rect 30570 1675 30575 1705
rect 30535 1670 30575 1675
rect 29800 1650 29820 1670
rect 29730 1645 29765 1650
rect 29730 1605 29765 1610
rect 29790 1645 29825 1650
rect 29790 1605 29825 1610
rect 30750 1440 30770 1725
rect 30785 1650 30825 1655
rect 30785 1620 30790 1650
rect 30820 1620 30825 1650
rect 30785 1615 30825 1620
rect 30740 1435 30780 1440
rect 30740 1405 30745 1435
rect 30775 1405 30780 1435
rect 30740 1400 30780 1405
rect 29875 1320 29915 1325
rect 29875 1290 29880 1320
rect 29910 1290 29915 1320
rect 29875 1285 29915 1290
rect 29965 1320 30005 1325
rect 29965 1290 29970 1320
rect 30000 1290 30005 1320
rect 29965 1285 30005 1290
rect 30795 940 30815 1615
rect 30235 935 30275 940
rect 30235 905 30240 935
rect 30270 905 30275 935
rect 30235 900 30275 905
rect 30335 935 30375 940
rect 30335 905 30340 935
rect 30370 905 30375 935
rect 30335 900 30375 905
rect 30435 935 30475 940
rect 30435 905 30440 935
rect 30470 905 30475 935
rect 30435 900 30475 905
rect 30785 935 30825 940
rect 30785 905 30790 935
rect 30820 905 30825 935
rect 30785 900 30825 905
rect 30345 880 30365 900
rect 30335 875 30375 880
rect 30335 845 30340 875
rect 30370 845 30375 875
rect 30795 865 30815 900
rect 30335 840 30375 845
rect 30785 860 30825 865
rect 30785 830 30790 860
rect 30820 830 30825 860
rect 30785 825 30825 830
rect 30795 500 30815 825
rect 30840 745 30860 2195
rect 30885 1825 30905 2295
rect 31680 2290 31700 2340
rect 32100 2290 32120 2340
rect 32880 2335 32900 3995
rect 32960 3850 33000 3855
rect 32960 3820 32965 3850
rect 32995 3820 33000 3850
rect 32960 3815 33000 3820
rect 32915 3760 32955 3765
rect 32915 3730 32920 3760
rect 32950 3730 32955 3760
rect 32915 3725 32955 3730
rect 32870 2330 32910 2335
rect 32870 2300 32875 2330
rect 32905 2300 32910 2330
rect 32870 2295 32910 2300
rect 31240 2285 31280 2290
rect 31240 2255 31245 2285
rect 31275 2255 31280 2285
rect 31240 2250 31280 2255
rect 31350 2285 31390 2290
rect 31350 2255 31355 2285
rect 31385 2255 31390 2285
rect 31350 2250 31390 2255
rect 31460 2285 31500 2290
rect 31460 2255 31465 2285
rect 31495 2255 31500 2285
rect 31460 2250 31500 2255
rect 31570 2285 31610 2290
rect 31570 2255 31575 2285
rect 31605 2255 31610 2285
rect 31570 2250 31610 2255
rect 31680 2285 31720 2290
rect 31680 2255 31685 2285
rect 31715 2255 31720 2285
rect 31680 2250 31720 2255
rect 31790 2285 31830 2290
rect 31790 2255 31795 2285
rect 31825 2255 31830 2285
rect 31790 2250 31830 2255
rect 31970 2285 32010 2290
rect 31970 2255 31975 2285
rect 32005 2255 32010 2285
rect 31970 2250 32010 2255
rect 32080 2285 32120 2290
rect 32080 2255 32085 2285
rect 32115 2255 32120 2285
rect 32080 2250 32120 2255
rect 32190 2285 32230 2290
rect 32190 2255 32195 2285
rect 32225 2255 32230 2285
rect 32190 2250 32230 2255
rect 32300 2285 32340 2290
rect 32300 2255 32305 2285
rect 32335 2255 32340 2285
rect 32300 2250 32340 2255
rect 32410 2285 32450 2290
rect 32410 2255 32415 2285
rect 32445 2255 32450 2285
rect 32410 2250 32450 2255
rect 32520 2285 32560 2290
rect 32520 2255 32525 2285
rect 32555 2255 32560 2285
rect 32520 2250 32560 2255
rect 31250 2235 31270 2250
rect 31360 2235 31380 2250
rect 31470 2235 31490 2250
rect 31580 2235 31600 2250
rect 31690 2235 31710 2250
rect 31800 2235 31820 2250
rect 31980 2235 32000 2250
rect 32090 2235 32110 2250
rect 32200 2235 32220 2250
rect 32310 2235 32330 2250
rect 32420 2235 32440 2250
rect 32530 2235 32550 2250
rect 31240 2225 31280 2235
rect 31240 2205 31250 2225
rect 31270 2205 31280 2225
rect 31240 2195 31280 2205
rect 31350 2225 31390 2235
rect 31350 2205 31360 2225
rect 31380 2205 31390 2225
rect 31350 2195 31390 2205
rect 31460 2225 31500 2235
rect 31460 2205 31470 2225
rect 31490 2205 31500 2225
rect 31460 2195 31500 2205
rect 31520 2230 31550 2235
rect 31520 2195 31550 2200
rect 31570 2225 31610 2235
rect 31570 2205 31580 2225
rect 31600 2205 31610 2225
rect 31570 2195 31610 2205
rect 31680 2225 31720 2235
rect 31680 2205 31690 2225
rect 31710 2205 31720 2225
rect 31680 2195 31720 2205
rect 31790 2225 31830 2235
rect 31790 2205 31800 2225
rect 31820 2205 31830 2225
rect 31790 2195 31830 2205
rect 31970 2225 32010 2235
rect 31970 2205 31980 2225
rect 32000 2205 32010 2225
rect 31970 2195 32010 2205
rect 32080 2225 32120 2235
rect 32080 2205 32090 2225
rect 32110 2205 32120 2225
rect 32080 2195 32120 2205
rect 32190 2225 32230 2235
rect 32190 2205 32200 2225
rect 32220 2205 32230 2225
rect 32190 2195 32230 2205
rect 32250 2230 32280 2235
rect 32250 2195 32280 2200
rect 32300 2225 32340 2235
rect 32300 2205 32310 2225
rect 32330 2205 32340 2225
rect 32300 2195 32340 2205
rect 32410 2225 32450 2235
rect 32410 2205 32420 2225
rect 32440 2205 32450 2225
rect 32410 2195 32450 2205
rect 32520 2225 32560 2235
rect 32520 2205 32530 2225
rect 32550 2205 32560 2225
rect 32520 2195 32560 2205
rect 31295 2005 31335 2015
rect 31295 1985 31305 2005
rect 31325 1985 31335 2005
rect 31295 1975 31335 1985
rect 31405 2005 31445 2015
rect 31405 1985 31415 2005
rect 31435 1985 31445 2005
rect 31405 1975 31445 1985
rect 31515 2005 31555 2015
rect 31515 1985 31525 2005
rect 31545 1985 31555 2005
rect 31515 1975 31555 1985
rect 31625 2005 31665 2015
rect 31625 1985 31635 2005
rect 31655 1985 31665 2005
rect 31625 1975 31665 1985
rect 31735 2005 31775 2015
rect 31735 1985 31745 2005
rect 31765 1985 31775 2005
rect 31735 1975 31775 1985
rect 32025 2005 32065 2015
rect 32025 1985 32035 2005
rect 32055 1985 32065 2005
rect 32025 1975 32065 1985
rect 32135 2005 32175 2015
rect 32135 1985 32145 2005
rect 32165 1985 32175 2005
rect 32135 1975 32175 1985
rect 32245 2005 32285 2015
rect 32245 1985 32255 2005
rect 32275 1985 32285 2005
rect 32245 1975 32285 1985
rect 32355 2005 32395 2015
rect 32355 1985 32365 2005
rect 32385 1985 32395 2005
rect 32355 1975 32395 1985
rect 32465 2005 32505 2015
rect 32465 1985 32475 2005
rect 32495 1985 32505 2005
rect 32465 1975 32505 1985
rect 31305 1955 31325 1975
rect 31415 1955 31435 1975
rect 31525 1955 31545 1975
rect 31635 1955 31655 1975
rect 31745 1955 31765 1975
rect 32035 1955 32055 1975
rect 32145 1955 32165 1975
rect 32255 1955 32275 1975
rect 32365 1955 32385 1975
rect 32475 1955 32495 1975
rect 31295 1950 31335 1955
rect 31295 1920 31300 1950
rect 31330 1920 31335 1950
rect 31295 1915 31335 1920
rect 31405 1950 31445 1955
rect 31405 1920 31410 1950
rect 31440 1920 31445 1950
rect 31405 1915 31445 1920
rect 31515 1950 31555 1955
rect 31515 1920 31520 1950
rect 31550 1920 31555 1950
rect 31515 1915 31555 1920
rect 31625 1950 31665 1955
rect 31625 1920 31630 1950
rect 31660 1920 31665 1950
rect 31625 1915 31665 1920
rect 31735 1950 31775 1955
rect 31735 1920 31740 1950
rect 31770 1920 31775 1950
rect 31735 1915 31775 1920
rect 31880 1945 31920 1955
rect 31880 1925 31890 1945
rect 31910 1925 31920 1945
rect 31880 1915 31920 1925
rect 32025 1950 32065 1955
rect 32025 1920 32030 1950
rect 32060 1920 32065 1950
rect 32025 1915 32065 1920
rect 32135 1950 32175 1955
rect 32135 1920 32140 1950
rect 32170 1920 32175 1950
rect 32135 1915 32175 1920
rect 32245 1950 32285 1955
rect 32245 1920 32250 1950
rect 32280 1920 32285 1950
rect 32245 1915 32285 1920
rect 32355 1950 32395 1955
rect 32355 1920 32360 1950
rect 32390 1920 32395 1950
rect 32355 1915 32395 1920
rect 32465 1950 32505 1955
rect 32465 1920 32470 1950
rect 32500 1920 32505 1950
rect 32465 1915 32505 1920
rect 31190 1895 31230 1900
rect 31190 1865 31195 1895
rect 31225 1865 31230 1895
rect 31190 1860 31230 1865
rect 31410 1895 31450 1900
rect 31410 1865 31415 1895
rect 31445 1865 31450 1895
rect 31410 1860 31450 1865
rect 30875 1820 30915 1825
rect 30875 1790 30880 1820
rect 30910 1790 30915 1820
rect 30875 1785 30915 1790
rect 31085 1805 31125 1810
rect 31085 1775 31090 1805
rect 31120 1775 31125 1805
rect 31085 1770 31125 1775
rect 31100 1755 31120 1770
rect 31200 1755 31220 1860
rect 31305 1805 31345 1810
rect 31305 1775 31310 1805
rect 31340 1775 31345 1805
rect 31305 1770 31345 1775
rect 31100 1745 31126 1755
rect 31100 1725 31103 1745
rect 31123 1725 31126 1745
rect 31100 1715 31126 1725
rect 31194 1745 31220 1755
rect 31194 1725 31197 1745
rect 31217 1725 31220 1745
rect 31237 1760 31269 1765
rect 31237 1730 31240 1760
rect 31266 1730 31269 1760
rect 31237 1725 31269 1730
rect 31320 1755 31340 1770
rect 31420 1755 31440 1860
rect 31535 1810 31555 1915
rect 31640 1895 31680 1900
rect 31640 1865 31645 1895
rect 31675 1865 31680 1895
rect 31640 1860 31680 1865
rect 31525 1805 31565 1810
rect 31525 1775 31530 1805
rect 31560 1775 31565 1805
rect 31525 1770 31565 1775
rect 31320 1745 31346 1755
rect 31320 1725 31323 1745
rect 31343 1725 31346 1745
rect 31194 1715 31220 1725
rect 31320 1715 31346 1725
rect 31414 1745 31440 1755
rect 31414 1725 31417 1745
rect 31437 1725 31440 1745
rect 31457 1760 31489 1765
rect 31457 1730 31460 1760
rect 31486 1730 31489 1760
rect 31457 1725 31489 1730
rect 31540 1755 31560 1770
rect 31601 1760 31633 1765
rect 31540 1745 31566 1755
rect 31540 1725 31543 1745
rect 31563 1725 31566 1745
rect 31601 1730 31604 1760
rect 31630 1730 31633 1760
rect 31601 1725 31633 1730
rect 31650 1755 31670 1860
rect 31820 1850 31860 1855
rect 31820 1820 31825 1850
rect 31855 1820 31860 1850
rect 31890 1825 31910 1915
rect 32245 1900 32265 1915
rect 32230 1895 32270 1900
rect 32230 1865 32235 1895
rect 32265 1865 32270 1895
rect 32230 1860 32270 1865
rect 32450 1895 32490 1900
rect 32450 1865 32455 1895
rect 32485 1865 32490 1895
rect 32450 1860 32490 1865
rect 32680 1895 32720 1900
rect 32680 1865 32685 1895
rect 32715 1865 32720 1895
rect 32680 1860 32720 1865
rect 31940 1850 31980 1855
rect 31820 1815 31860 1820
rect 31880 1815 31920 1825
rect 31940 1820 31945 1850
rect 31975 1820 31980 1850
rect 31940 1815 31980 1820
rect 31830 1765 31850 1815
rect 31880 1795 31890 1815
rect 31910 1795 31920 1815
rect 31880 1785 31920 1795
rect 31950 1765 31970 1815
rect 32125 1805 32165 1810
rect 32125 1775 32130 1805
rect 32160 1775 32165 1805
rect 32125 1770 32165 1775
rect 31824 1755 31850 1765
rect 31650 1745 31676 1755
rect 31650 1725 31653 1745
rect 31673 1725 31676 1745
rect 31824 1735 31827 1755
rect 31847 1735 31850 1755
rect 31824 1725 31850 1735
rect 31867 1760 31899 1765
rect 31867 1730 31870 1760
rect 31896 1730 31899 1760
rect 31867 1725 31899 1730
rect 31947 1755 31973 1765
rect 31947 1735 31950 1755
rect 31970 1735 31973 1755
rect 31947 1725 31973 1735
rect 32140 1755 32160 1770
rect 32240 1755 32260 1860
rect 32345 1805 32385 1810
rect 32345 1775 32350 1805
rect 32380 1775 32385 1805
rect 32345 1770 32385 1775
rect 32140 1745 32166 1755
rect 32140 1725 32143 1745
rect 32163 1725 32166 1745
rect 31414 1715 31440 1725
rect 31540 1715 31566 1725
rect 31650 1715 31676 1725
rect 32140 1715 32166 1725
rect 32234 1745 32260 1755
rect 32234 1725 32237 1745
rect 32257 1725 32260 1745
rect 32277 1760 32309 1765
rect 32277 1730 32280 1760
rect 32306 1730 32309 1760
rect 32277 1725 32309 1730
rect 32360 1755 32380 1770
rect 32460 1755 32480 1860
rect 32565 1805 32605 1810
rect 32565 1775 32570 1805
rect 32600 1775 32605 1805
rect 32565 1770 32605 1775
rect 32360 1745 32386 1755
rect 32360 1725 32363 1745
rect 32383 1725 32386 1745
rect 32234 1715 32260 1725
rect 32360 1715 32386 1725
rect 32454 1745 32480 1755
rect 32454 1725 32457 1745
rect 32477 1725 32480 1745
rect 32497 1760 32529 1765
rect 32497 1730 32500 1760
rect 32526 1730 32529 1760
rect 32497 1725 32529 1730
rect 32580 1755 32600 1770
rect 32641 1760 32673 1765
rect 32580 1745 32606 1755
rect 32580 1725 32583 1745
rect 32603 1725 32606 1745
rect 32641 1730 32644 1760
rect 32670 1730 32673 1760
rect 32641 1725 32673 1730
rect 32690 1755 32710 1860
rect 32880 1830 32900 2295
rect 32870 1825 32910 1830
rect 32870 1795 32875 1825
rect 32905 1795 32910 1825
rect 32870 1790 32910 1795
rect 32690 1745 32716 1755
rect 32690 1725 32693 1745
rect 32713 1725 32716 1745
rect 32454 1715 32480 1725
rect 32580 1715 32606 1725
rect 32690 1715 32716 1725
rect 30940 1650 30980 1655
rect 30940 1620 30945 1650
rect 30975 1620 30980 1650
rect 30940 1615 30980 1620
rect 31106 1540 31138 1545
rect 31106 1510 31109 1540
rect 31135 1510 31138 1540
rect 31106 1505 31138 1510
rect 31155 1535 31181 1545
rect 31155 1515 31158 1535
rect 31178 1515 31181 1535
rect 31155 1505 31181 1515
rect 31256 1535 31283 1545
rect 31256 1515 31260 1535
rect 31280 1515 31283 1535
rect 31256 1505 31283 1515
rect 31305 1540 31345 1545
rect 31305 1510 31310 1540
rect 31340 1510 31345 1540
rect 31305 1505 31345 1510
rect 31366 1535 31393 1545
rect 31366 1515 31370 1535
rect 31390 1515 31393 1535
rect 31366 1505 31393 1515
rect 31476 1535 31503 1545
rect 31476 1515 31480 1535
rect 31500 1515 31503 1535
rect 31476 1505 31503 1515
rect 31525 1540 31565 1545
rect 31525 1510 31530 1540
rect 31560 1510 31565 1540
rect 31525 1505 31565 1510
rect 31586 1535 31613 1545
rect 31586 1515 31590 1535
rect 31610 1515 31613 1535
rect 31586 1505 31613 1515
rect 31825 1535 31855 1545
rect 31825 1515 31830 1535
rect 31850 1515 31855 1535
rect 31825 1505 31855 1515
rect 31875 1535 31905 1545
rect 31875 1515 31880 1535
rect 31900 1515 31905 1535
rect 31875 1505 31905 1515
rect 31922 1540 31954 1545
rect 31922 1510 31925 1540
rect 31951 1510 31954 1540
rect 31922 1505 31954 1510
rect 32146 1540 32178 1545
rect 32146 1510 32149 1540
rect 32175 1510 32178 1540
rect 32146 1505 32178 1510
rect 32195 1535 32221 1545
rect 32195 1515 32198 1535
rect 32218 1515 32221 1535
rect 32195 1505 32221 1515
rect 32296 1535 32323 1545
rect 32296 1515 32300 1535
rect 32320 1515 32323 1535
rect 32296 1505 32323 1515
rect 32345 1540 32385 1545
rect 32345 1510 32350 1540
rect 32380 1510 32385 1540
rect 32345 1505 32385 1510
rect 32406 1535 32433 1545
rect 32406 1515 32410 1535
rect 32430 1515 32433 1535
rect 32406 1505 32433 1515
rect 32516 1535 32543 1545
rect 32516 1515 32520 1535
rect 32540 1515 32543 1535
rect 32516 1505 32543 1515
rect 32565 1540 32605 1545
rect 32565 1510 32570 1540
rect 32600 1510 32605 1540
rect 32565 1505 32605 1510
rect 32626 1535 32653 1545
rect 32626 1515 32630 1535
rect 32650 1515 32653 1535
rect 32626 1505 32653 1515
rect 31155 1485 31175 1505
rect 31260 1485 31280 1505
rect 31370 1485 31390 1505
rect 31480 1485 31500 1505
rect 31590 1485 31610 1505
rect 31145 1480 31185 1485
rect 31145 1450 31150 1480
rect 31180 1450 31185 1480
rect 31145 1445 31185 1450
rect 31250 1480 31290 1485
rect 31250 1450 31255 1480
rect 31285 1450 31290 1480
rect 31250 1445 31290 1450
rect 31360 1480 31400 1485
rect 31360 1450 31365 1480
rect 31395 1450 31400 1480
rect 31360 1445 31400 1450
rect 31470 1480 31510 1485
rect 31470 1450 31475 1480
rect 31505 1450 31510 1480
rect 31470 1445 31510 1450
rect 31580 1480 31620 1485
rect 31580 1450 31585 1480
rect 31615 1450 31620 1480
rect 31580 1445 31620 1450
rect 31005 1390 31045 1395
rect 31005 1360 31010 1390
rect 31040 1360 31045 1390
rect 31005 1355 31045 1360
rect 31755 1390 31795 1395
rect 31755 1360 31760 1390
rect 31790 1360 31795 1390
rect 31755 1355 31795 1360
rect 31015 845 31035 1355
rect 31315 1345 31355 1350
rect 31315 1315 31320 1345
rect 31350 1315 31355 1345
rect 31315 1310 31355 1315
rect 31325 1260 31345 1310
rect 31765 1260 31785 1355
rect 31825 1260 31845 1505
rect 31880 1350 31900 1505
rect 32195 1485 32215 1505
rect 32300 1485 32320 1505
rect 32410 1485 32430 1505
rect 32520 1485 32540 1505
rect 32630 1485 32650 1505
rect 32185 1480 32225 1485
rect 32185 1450 32190 1480
rect 32220 1450 32225 1480
rect 32185 1445 32225 1450
rect 32290 1480 32330 1485
rect 32290 1450 32295 1480
rect 32325 1450 32330 1480
rect 32290 1445 32330 1450
rect 32400 1480 32440 1485
rect 32400 1450 32405 1480
rect 32435 1450 32440 1480
rect 32400 1445 32440 1450
rect 32510 1480 32550 1485
rect 32510 1450 32515 1480
rect 32545 1450 32550 1480
rect 32510 1445 32550 1450
rect 32620 1480 32660 1485
rect 32620 1450 32625 1480
rect 32655 1450 32660 1480
rect 32620 1445 32660 1450
rect 31870 1345 31910 1350
rect 31870 1315 31875 1345
rect 31905 1315 31910 1345
rect 31870 1310 31910 1315
rect 32195 1260 32215 1445
rect 32925 1370 32945 3725
rect 32375 1365 32415 1370
rect 32375 1335 32380 1365
rect 32410 1335 32415 1365
rect 32375 1330 32415 1335
rect 32915 1365 32955 1370
rect 32915 1335 32920 1365
rect 32950 1335 32955 1365
rect 32915 1330 32955 1335
rect 32385 1260 32405 1330
rect 31315 1250 31355 1260
rect 31315 1230 31325 1250
rect 31345 1230 31355 1250
rect 31315 1220 31355 1230
rect 31425 1255 31465 1260
rect 31425 1225 31430 1255
rect 31460 1225 31465 1255
rect 31425 1220 31465 1225
rect 31535 1255 31575 1260
rect 31535 1225 31540 1255
rect 31570 1225 31575 1255
rect 31535 1220 31575 1225
rect 31645 1255 31685 1260
rect 31645 1225 31650 1255
rect 31680 1225 31685 1255
rect 31645 1220 31685 1225
rect 31755 1255 31795 1260
rect 31755 1225 31760 1255
rect 31790 1225 31795 1255
rect 31755 1220 31795 1225
rect 31815 1250 31845 1260
rect 31815 1230 31820 1250
rect 31840 1230 31845 1250
rect 31815 1220 31845 1230
rect 31865 1255 31905 1260
rect 31865 1225 31870 1255
rect 31900 1225 31905 1255
rect 31865 1220 31905 1225
rect 31975 1255 32015 1260
rect 31975 1225 31980 1255
rect 32010 1225 32015 1255
rect 31975 1220 32015 1225
rect 32085 1255 32125 1260
rect 32085 1225 32090 1255
rect 32120 1225 32125 1255
rect 32085 1220 32125 1225
rect 32195 1255 32235 1260
rect 32195 1225 32200 1255
rect 32230 1225 32235 1255
rect 32195 1220 32235 1225
rect 32305 1255 32345 1260
rect 32305 1225 32310 1255
rect 32340 1225 32345 1255
rect 32305 1220 32345 1225
rect 32381 1250 32411 1260
rect 32381 1230 32386 1250
rect 32406 1230 32411 1250
rect 32381 1220 32411 1230
rect 32430 1255 32470 1260
rect 32430 1225 32435 1255
rect 32465 1225 32470 1255
rect 32430 1220 32470 1225
rect 31195 935 31235 940
rect 31195 905 31200 935
rect 31230 905 31235 935
rect 31195 900 31235 905
rect 31260 935 31300 940
rect 31260 905 31265 935
rect 31295 905 31300 935
rect 31260 900 31300 905
rect 31370 935 31410 940
rect 31370 905 31375 935
rect 31405 905 31410 935
rect 31370 900 31410 905
rect 31480 935 31520 940
rect 31480 905 31485 935
rect 31515 905 31520 935
rect 31480 900 31520 905
rect 31590 935 31630 940
rect 31590 905 31595 935
rect 31625 905 31630 935
rect 31590 900 31630 905
rect 31700 935 31740 940
rect 31700 905 31705 935
rect 31735 905 31740 935
rect 31700 900 31740 905
rect 31810 935 31850 940
rect 31810 905 31815 935
rect 31845 905 31850 935
rect 31810 900 31850 905
rect 31920 935 31960 940
rect 31920 905 31925 935
rect 31955 905 31960 935
rect 31920 900 31960 905
rect 32030 935 32070 940
rect 32030 905 32035 935
rect 32065 905 32070 935
rect 32030 900 32070 905
rect 32140 935 32180 940
rect 32140 905 32145 935
rect 32175 905 32180 935
rect 32140 900 32180 905
rect 32250 935 32290 940
rect 32250 905 32255 935
rect 32285 905 32290 935
rect 32250 900 32290 905
rect 32360 935 32400 940
rect 32360 905 32365 935
rect 32395 905 32400 935
rect 32360 900 32400 905
rect 32475 935 32515 940
rect 32475 905 32480 935
rect 32510 905 32515 935
rect 32475 900 32515 905
rect 31005 840 31045 845
rect 31005 810 31010 840
rect 31040 810 31045 840
rect 31005 805 31045 810
rect 31505 840 31545 845
rect 31505 810 31510 840
rect 31540 810 31545 840
rect 31505 805 31545 810
rect 31935 840 31975 845
rect 31935 810 31940 840
rect 31970 810 31975 840
rect 31935 805 31975 810
rect 32155 840 32195 845
rect 32155 810 32160 840
rect 32190 810 32195 840
rect 32155 805 32195 810
rect 32375 840 32415 845
rect 32375 810 32380 840
rect 32410 810 32415 840
rect 32375 805 32415 810
rect 31515 745 31535 805
rect 30830 740 30870 745
rect 30830 710 30835 740
rect 30865 710 30870 740
rect 30830 705 30870 710
rect 31305 740 31345 745
rect 31305 710 31310 740
rect 31340 710 31345 740
rect 31305 705 31345 710
rect 31375 740 31415 745
rect 31375 710 31380 740
rect 31410 710 31415 740
rect 31375 705 31415 710
rect 31445 740 31485 745
rect 31445 710 31450 740
rect 31480 710 31485 740
rect 31445 705 31485 710
rect 31505 735 31545 745
rect 31945 740 31965 805
rect 32165 740 32185 805
rect 32385 740 32405 805
rect 32925 740 32945 1330
rect 32970 845 32990 3815
rect 34155 3735 34195 3740
rect 33005 3715 33045 3720
rect 33005 3685 33010 3715
rect 33040 3685 33045 3715
rect 33005 3680 33045 3685
rect 33145 3715 33185 3720
rect 33145 3685 33150 3715
rect 33180 3685 33185 3715
rect 33145 3680 33185 3685
rect 33255 3715 33295 3720
rect 33255 3685 33260 3715
rect 33290 3685 33295 3715
rect 33255 3680 33295 3685
rect 33365 3715 33405 3720
rect 33365 3685 33370 3715
rect 33400 3685 33405 3715
rect 33365 3680 33405 3685
rect 33475 3715 33515 3720
rect 33475 3685 33480 3715
rect 33510 3685 33515 3715
rect 33475 3680 33515 3685
rect 33585 3715 33625 3720
rect 33585 3685 33590 3715
rect 33620 3685 33625 3715
rect 33585 3680 33625 3685
rect 33695 3715 33735 3720
rect 33695 3685 33700 3715
rect 33730 3685 33735 3715
rect 33695 3680 33735 3685
rect 33805 3715 33845 3720
rect 33805 3685 33810 3715
rect 33840 3685 33845 3715
rect 34155 3705 34160 3735
rect 34190 3705 34195 3735
rect 34155 3700 34195 3705
rect 33805 3680 33845 3685
rect 33005 1930 33025 3680
rect 34165 3660 34185 3700
rect 34105 3655 34246 3660
rect 34105 3625 34111 3655
rect 34141 3625 34160 3655
rect 34190 3625 34210 3655
rect 34240 3625 34246 3655
rect 34105 3620 34246 3625
rect 34105 3050 34246 3055
rect 33200 3045 33240 3050
rect 33200 3015 33205 3045
rect 33235 3015 33240 3045
rect 33200 3010 33240 3015
rect 33310 3045 33350 3050
rect 33310 3015 33315 3045
rect 33345 3015 33350 3045
rect 33310 3010 33350 3015
rect 33420 3045 33460 3050
rect 33420 3015 33425 3045
rect 33455 3015 33460 3045
rect 33420 3010 33460 3015
rect 33530 3045 33570 3050
rect 33530 3015 33535 3045
rect 33565 3015 33570 3045
rect 33530 3010 33570 3015
rect 33588 3040 33622 3050
rect 33588 3020 33596 3040
rect 33614 3020 33622 3040
rect 33588 3010 33622 3020
rect 33640 3045 33680 3050
rect 33640 3015 33645 3045
rect 33675 3015 33680 3045
rect 33640 3010 33680 3015
rect 33750 3045 33790 3050
rect 33750 3015 33755 3045
rect 33785 3015 33790 3045
rect 34105 3020 34111 3050
rect 34141 3020 34160 3050
rect 34190 3020 34210 3050
rect 34240 3020 34246 3050
rect 34105 3015 34246 3020
rect 33750 3010 33790 3015
rect 33040 2935 33080 2940
rect 33040 2905 33045 2935
rect 33075 2905 33080 2935
rect 33040 2900 33080 2905
rect 33050 2380 33070 2900
rect 33320 2895 33340 3010
rect 33475 2980 33515 2990
rect 33475 2960 33485 2980
rect 33505 2960 33515 2980
rect 33475 2950 33515 2960
rect 33310 2890 33350 2895
rect 33310 2860 33315 2890
rect 33345 2860 33350 2890
rect 33310 2855 33350 2860
rect 33485 2820 33505 2950
rect 33595 2940 33615 3010
rect 34165 2940 34185 3015
rect 34235 2985 34275 2995
rect 34235 2965 34245 2985
rect 34265 2965 34275 2985
rect 34235 2955 34275 2965
rect 33585 2935 33625 2940
rect 33585 2905 33590 2935
rect 33620 2905 33625 2935
rect 33585 2900 33625 2905
rect 34155 2935 34195 2940
rect 34155 2905 34160 2935
rect 34190 2905 34195 2935
rect 34155 2900 34195 2905
rect 33475 2810 33515 2820
rect 33475 2790 33485 2810
rect 33505 2790 33515 2810
rect 33475 2780 33515 2790
rect 33200 2755 33240 2760
rect 33200 2725 33205 2755
rect 33235 2725 33240 2755
rect 33200 2720 33240 2725
rect 33310 2755 33350 2760
rect 33310 2725 33315 2755
rect 33345 2725 33350 2755
rect 33310 2720 33350 2725
rect 33420 2755 33460 2760
rect 33420 2725 33425 2755
rect 33455 2725 33460 2755
rect 33420 2720 33460 2725
rect 33530 2755 33570 2760
rect 33530 2725 33535 2755
rect 33565 2725 33570 2755
rect 33530 2720 33570 2725
rect 33640 2755 33680 2760
rect 33640 2725 33645 2755
rect 33675 2725 33680 2755
rect 33640 2720 33680 2725
rect 33750 2755 33790 2760
rect 33750 2725 33755 2755
rect 33785 2725 33790 2755
rect 33750 2720 33790 2725
rect 34245 2689 34265 2955
rect 34445 2890 34485 2895
rect 34445 2860 34450 2890
rect 34480 2860 34485 2890
rect 34445 2855 34485 2860
rect 34235 2679 34275 2689
rect 34235 2659 34245 2679
rect 34265 2659 34275 2679
rect 34235 2649 34275 2659
rect 33255 2485 33295 2490
rect 33255 2455 33260 2485
rect 33290 2455 33295 2485
rect 33255 2450 33295 2455
rect 33313 2480 33347 2490
rect 33313 2460 33321 2480
rect 33339 2460 33347 2480
rect 33313 2450 33347 2460
rect 33365 2485 33405 2490
rect 33365 2455 33370 2485
rect 33400 2455 33405 2485
rect 33365 2450 33405 2455
rect 33475 2485 33515 2490
rect 33475 2455 33480 2485
rect 33510 2455 33515 2485
rect 33475 2450 33515 2455
rect 33585 2485 33625 2490
rect 33585 2455 33590 2485
rect 33620 2455 33625 2485
rect 33585 2450 33625 2455
rect 33695 2485 33735 2490
rect 33695 2455 33700 2485
rect 33730 2455 33735 2485
rect 33695 2450 33735 2455
rect 33975 2485 34015 2490
rect 33975 2455 33980 2485
rect 34010 2455 34015 2485
rect 33975 2450 34015 2455
rect 33320 2380 33340 2450
rect 33040 2375 33080 2380
rect 33040 2345 33045 2375
rect 33075 2345 33080 2375
rect 33040 2340 33080 2345
rect 33310 2375 33350 2380
rect 33310 2345 33315 2375
rect 33345 2345 33350 2375
rect 33310 2340 33350 2345
rect 33320 2300 33340 2340
rect 33255 2295 33295 2300
rect 33255 2265 33260 2295
rect 33290 2265 33295 2295
rect 33255 2260 33295 2265
rect 33313 2290 33347 2300
rect 33313 2270 33321 2290
rect 33339 2270 33347 2290
rect 33313 2260 33347 2270
rect 33365 2295 33405 2300
rect 33365 2265 33370 2295
rect 33400 2265 33405 2295
rect 33365 2260 33405 2265
rect 33475 2295 33515 2300
rect 33475 2265 33480 2295
rect 33510 2265 33515 2295
rect 33475 2260 33515 2265
rect 33585 2295 33625 2300
rect 33585 2265 33590 2295
rect 33620 2265 33625 2295
rect 33585 2260 33625 2265
rect 33695 2295 33735 2300
rect 33695 2265 33700 2295
rect 33730 2265 33735 2295
rect 33695 2260 33735 2265
rect 33930 2295 33970 2300
rect 33930 2265 33935 2295
rect 33965 2265 33970 2295
rect 33930 2260 33970 2265
rect 33875 2110 33915 2115
rect 33875 2080 33880 2110
rect 33910 2080 33915 2110
rect 33875 2075 33915 2080
rect 33940 1930 33960 2260
rect 33985 1985 34005 2450
rect 34455 2270 34475 2855
rect 34495 2755 34535 2760
rect 34495 2725 34500 2755
rect 34530 2725 34535 2755
rect 34495 2720 34535 2725
rect 34440 2260 34490 2270
rect 34440 2230 34450 2260
rect 34480 2230 34490 2260
rect 34440 2220 34490 2230
rect 34025 2110 34065 2115
rect 34025 2080 34030 2110
rect 34060 2080 34065 2110
rect 34025 2075 34065 2080
rect 34115 1985 34150 1990
rect 33975 1980 34015 1985
rect 33975 1950 33980 1980
rect 34010 1950 34015 1980
rect 33975 1945 34015 1950
rect 34115 1945 34150 1950
rect 34175 1985 34210 1991
rect 34175 1945 34210 1950
rect 34235 1985 34270 1990
rect 34235 1945 34270 1950
rect 34295 1985 34330 1991
rect 34295 1945 34330 1950
rect 34180 1930 34200 1945
rect 33005 1925 33045 1930
rect 33005 1895 33010 1925
rect 33040 1895 33045 1925
rect 33005 1890 33045 1895
rect 33200 1925 33240 1930
rect 33200 1895 33205 1925
rect 33235 1895 33240 1925
rect 33200 1890 33240 1895
rect 33310 1925 33350 1930
rect 33310 1895 33315 1925
rect 33345 1895 33350 1925
rect 33310 1890 33350 1895
rect 33420 1925 33460 1930
rect 33420 1895 33425 1925
rect 33455 1895 33460 1925
rect 33420 1890 33460 1895
rect 33530 1925 33570 1930
rect 33530 1895 33535 1925
rect 33565 1895 33570 1925
rect 33530 1890 33570 1895
rect 33640 1925 33680 1930
rect 33640 1895 33645 1925
rect 33675 1895 33680 1925
rect 33640 1890 33680 1895
rect 33750 1925 33790 1930
rect 33750 1895 33755 1925
rect 33785 1895 33790 1925
rect 33750 1890 33790 1895
rect 33930 1925 33970 1930
rect 33930 1895 33935 1925
rect 33965 1895 33970 1925
rect 33930 1890 33970 1895
rect 34170 1925 34210 1930
rect 34170 1895 34175 1925
rect 34205 1895 34210 1925
rect 34170 1890 34210 1895
rect 33475 1860 33515 1870
rect 33475 1840 33485 1860
rect 33505 1840 33515 1860
rect 33475 1830 33515 1840
rect 34300 1830 34320 1945
rect 33485 1770 33505 1830
rect 34290 1825 34330 1830
rect 34290 1795 34295 1825
rect 34325 1795 34330 1825
rect 34290 1790 34330 1795
rect 33015 1760 33055 1765
rect 33015 1730 33020 1760
rect 33050 1730 33055 1760
rect 33015 1725 33055 1730
rect 33325 1760 33365 1765
rect 33325 1730 33330 1760
rect 33360 1730 33365 1760
rect 33475 1760 33515 1770
rect 33475 1740 33485 1760
rect 33505 1740 33515 1760
rect 33475 1730 33515 1740
rect 34035 1760 34075 1765
rect 34035 1730 34040 1760
rect 34070 1730 34075 1760
rect 33325 1725 33365 1730
rect 34035 1725 34075 1730
rect 33025 1440 33045 1725
rect 33335 1710 33355 1725
rect 33225 1705 33265 1710
rect 33225 1675 33230 1705
rect 33260 1675 33265 1705
rect 33225 1670 33265 1675
rect 33328 1700 33362 1710
rect 33328 1680 33336 1700
rect 33354 1680 33362 1700
rect 33328 1670 33362 1680
rect 33425 1705 33465 1710
rect 33425 1675 33430 1705
rect 33460 1675 33465 1705
rect 33425 1670 33465 1675
rect 33625 1705 33665 1710
rect 33625 1675 33630 1705
rect 33660 1675 33665 1705
rect 33625 1670 33665 1675
rect 33970 1705 34010 1710
rect 33970 1675 33975 1705
rect 34005 1675 34010 1705
rect 33970 1670 34010 1675
rect 33980 1650 34000 1670
rect 34045 1650 34065 1725
rect 34455 1710 34475 2220
rect 34445 1705 34485 1710
rect 34445 1675 34450 1705
rect 34480 1675 34485 1705
rect 34445 1670 34485 1675
rect 33975 1645 34010 1650
rect 33975 1605 34010 1610
rect 34035 1645 34070 1650
rect 34035 1605 34070 1610
rect 33015 1435 33055 1440
rect 33015 1405 33020 1435
rect 33050 1405 33055 1435
rect 33015 1400 33055 1405
rect 33795 1320 33835 1325
rect 33795 1290 33800 1320
rect 33830 1290 33835 1320
rect 33795 1285 33835 1290
rect 33885 1320 33925 1325
rect 33885 1290 33890 1320
rect 33920 1290 33925 1320
rect 33885 1285 33925 1290
rect 33015 935 33055 940
rect 33015 905 33020 935
rect 33050 905 33055 935
rect 33015 900 33055 905
rect 33325 935 33365 940
rect 33325 905 33330 935
rect 33360 905 33365 935
rect 33325 900 33365 905
rect 33425 935 33465 940
rect 33425 905 33430 935
rect 33460 905 33465 935
rect 33425 900 33465 905
rect 33525 935 33565 940
rect 33525 905 33530 935
rect 33560 905 33565 935
rect 33525 900 33565 905
rect 32960 840 33000 845
rect 32960 810 32965 840
rect 32995 810 33000 840
rect 32960 805 33000 810
rect 31505 715 31515 735
rect 31535 715 31545 735
rect 31505 705 31545 715
rect 31935 730 31975 740
rect 31935 710 31945 730
rect 31965 710 31975 730
rect 31935 700 31975 710
rect 32045 735 32085 740
rect 32045 705 32050 735
rect 32080 705 32085 735
rect 32045 700 32085 705
rect 32155 730 32195 740
rect 32155 710 32165 730
rect 32185 710 32195 730
rect 32155 700 32195 710
rect 32265 735 32305 740
rect 32265 705 32270 735
rect 32300 705 32305 735
rect 32265 700 32305 705
rect 32375 730 32415 740
rect 32375 710 32385 730
rect 32405 710 32415 730
rect 32375 700 32415 710
rect 32485 735 32525 740
rect 32485 705 32490 735
rect 32520 705 32525 735
rect 32485 700 32525 705
rect 32915 735 32955 740
rect 32915 705 32920 735
rect 32950 705 32955 735
rect 32915 700 32955 705
rect 31990 615 32030 620
rect 31990 585 31995 615
rect 32025 585 32030 615
rect 31990 580 32030 585
rect 32100 615 32140 620
rect 32100 585 32105 615
rect 32135 585 32140 615
rect 32100 580 32140 585
rect 32210 615 32250 620
rect 32210 585 32215 615
rect 32245 585 32250 615
rect 32210 580 32250 585
rect 32320 615 32360 620
rect 32320 585 32325 615
rect 32355 585 32360 615
rect 32320 580 32360 585
rect 32430 615 32470 620
rect 32430 585 32435 615
rect 32465 585 32470 615
rect 32430 580 32470 585
rect 32220 560 32240 580
rect 31375 545 31415 555
rect 31375 525 31385 545
rect 31405 525 31415 545
rect 31375 515 31415 525
rect 32210 550 32250 560
rect 32210 530 32220 550
rect 32240 530 32250 550
rect 32210 520 32250 530
rect 31385 500 31405 515
rect 32220 500 32240 520
rect 33025 500 33045 900
rect 33435 880 33455 900
rect 33425 875 33465 880
rect 33425 845 33430 875
rect 33460 845 33465 875
rect 33425 840 33465 845
rect 34505 500 34525 2720
rect 29265 495 29305 500
rect 29265 465 29270 495
rect 29300 465 29305 495
rect 29265 460 29305 465
rect 30785 495 30825 500
rect 30785 465 30790 495
rect 30820 465 30825 495
rect 30785 460 30825 465
rect 31375 495 31415 500
rect 31375 465 31380 495
rect 31410 465 31415 495
rect 31375 460 31415 465
rect 32210 495 32250 500
rect 32210 465 32215 495
rect 32245 465 32250 495
rect 32210 460 32250 465
rect 33015 495 33055 500
rect 33015 465 33020 495
rect 33050 465 33055 495
rect 33015 460 33055 465
rect 34495 495 34535 500
rect 34495 465 34500 495
rect 34530 465 34535 495
rect 34495 460 34535 465
rect 30795 -510 30815 460
rect 30785 -515 30825 -510
rect 30785 -545 30790 -515
rect 30820 -545 30825 -515
rect 30785 -550 30825 -545
<< via1 >>
rect 30790 6155 30820 6185
rect 31535 4915 31565 4945
rect 31655 4915 31685 4945
rect 31775 4915 31805 4945
rect 32445 4900 32475 4930
rect 30790 4840 30820 4870
rect 31285 4865 31315 4870
rect 31285 4845 31290 4865
rect 31290 4845 31310 4865
rect 31310 4845 31315 4865
rect 31285 4840 31315 4845
rect 31475 4880 31505 4885
rect 31475 4860 31480 4880
rect 31480 4860 31500 4880
rect 31500 4860 31505 4880
rect 31475 4855 31505 4860
rect 31595 4880 31625 4885
rect 31595 4860 31600 4880
rect 31600 4860 31620 4880
rect 31620 4860 31625 4880
rect 31595 4855 31625 4860
rect 31715 4880 31745 4885
rect 31715 4860 31720 4880
rect 31720 4860 31740 4880
rect 31740 4860 31745 4880
rect 31715 4855 31745 4860
rect 31835 4880 31865 4885
rect 31835 4860 31840 4880
rect 31840 4860 31860 4880
rect 31860 4860 31865 4880
rect 31835 4855 31865 4860
rect 32205 4855 32235 4860
rect 32205 4835 32210 4855
rect 32210 4835 32230 4855
rect 32230 4835 32235 4855
rect 32205 4830 32235 4835
rect 32325 4855 32355 4860
rect 32325 4835 32330 4855
rect 32330 4835 32350 4855
rect 32350 4835 32355 4855
rect 32325 4830 32355 4835
rect 32445 4855 32475 4860
rect 32445 4835 32450 4855
rect 32450 4835 32470 4855
rect 32470 4835 32475 4855
rect 32445 4830 32475 4835
rect 32565 4855 32595 4860
rect 32565 4835 32570 4855
rect 32570 4835 32590 4855
rect 32590 4835 32595 4855
rect 32565 4830 32595 4835
rect 32685 4855 32715 4860
rect 32685 4835 32690 4855
rect 32690 4835 32710 4855
rect 32710 4835 32715 4855
rect 32685 4830 32715 4835
rect 31005 4700 31035 4730
rect 31655 4725 31685 4730
rect 31655 4705 31660 4725
rect 31660 4705 31680 4725
rect 31680 4705 31685 4725
rect 31655 4700 31685 4705
rect 30790 4410 30820 4440
rect 30790 3940 30820 3970
rect 29610 3705 29640 3735
rect 29960 3710 29990 3715
rect 29960 3690 29965 3710
rect 29965 3690 29985 3710
rect 29985 3690 29990 3710
rect 29960 3685 29990 3690
rect 30070 3710 30100 3715
rect 30070 3690 30075 3710
rect 30075 3690 30095 3710
rect 30095 3690 30100 3710
rect 30070 3685 30100 3690
rect 30180 3710 30210 3715
rect 30180 3690 30185 3710
rect 30185 3690 30205 3710
rect 30205 3690 30210 3710
rect 30180 3685 30210 3690
rect 30290 3710 30320 3715
rect 30290 3690 30295 3710
rect 30295 3690 30315 3710
rect 30315 3690 30320 3710
rect 30290 3685 30320 3690
rect 30400 3710 30430 3715
rect 30400 3690 30405 3710
rect 30405 3690 30425 3710
rect 30425 3690 30430 3710
rect 30400 3685 30430 3690
rect 30510 3710 30540 3715
rect 30510 3690 30515 3710
rect 30515 3690 30535 3710
rect 30535 3690 30540 3710
rect 30510 3685 30540 3690
rect 30620 3710 30650 3715
rect 30620 3690 30625 3710
rect 30625 3690 30645 3710
rect 30645 3690 30650 3710
rect 30620 3685 30650 3690
rect 30790 3685 30820 3715
rect 29560 3625 29590 3655
rect 29610 3625 29640 3655
rect 29659 3625 29689 3655
rect 29560 3020 29590 3050
rect 29610 3020 29640 3050
rect 29659 3020 29689 3050
rect 30015 3040 30045 3045
rect 30015 3020 30020 3040
rect 30020 3020 30040 3040
rect 30040 3020 30045 3040
rect 30015 3015 30045 3020
rect 29320 2840 29350 2870
rect 29270 2725 29300 2755
rect 30125 3040 30155 3045
rect 30125 3020 30130 3040
rect 30130 3020 30150 3040
rect 30150 3020 30155 3040
rect 30125 3015 30155 3020
rect 30235 3040 30265 3045
rect 30235 3020 30240 3040
rect 30240 3020 30260 3040
rect 30260 3020 30265 3040
rect 30235 3015 30265 3020
rect 30345 3040 30375 3045
rect 30345 3020 30350 3040
rect 30350 3020 30370 3040
rect 30370 3020 30375 3040
rect 30345 3015 30375 3020
rect 30455 3040 30485 3045
rect 30455 3020 30460 3040
rect 30460 3020 30480 3040
rect 30480 3020 30485 3040
rect 30455 3015 30485 3020
rect 30565 3040 30595 3045
rect 30565 3020 30570 3040
rect 30570 3020 30590 3040
rect 30590 3020 30595 3040
rect 30565 3015 30595 3020
rect 29610 2895 29640 2925
rect 30180 2895 30210 2925
rect 30745 2895 30775 2925
rect 30455 2840 30485 2870
rect 30015 2750 30045 2755
rect 30015 2730 30020 2750
rect 30020 2730 30040 2750
rect 30040 2730 30045 2750
rect 30015 2725 30045 2730
rect 30125 2750 30155 2755
rect 30125 2730 30130 2750
rect 30130 2730 30150 2750
rect 30150 2730 30155 2750
rect 30125 2725 30155 2730
rect 30235 2750 30265 2755
rect 30235 2730 30240 2750
rect 30240 2730 30260 2750
rect 30260 2730 30265 2750
rect 30235 2725 30265 2730
rect 30345 2750 30375 2755
rect 30345 2730 30350 2750
rect 30350 2730 30370 2750
rect 30370 2730 30375 2750
rect 30345 2725 30375 2730
rect 30455 2750 30485 2755
rect 30455 2730 30460 2750
rect 30460 2730 30480 2750
rect 30480 2730 30485 2750
rect 30455 2725 30485 2730
rect 30565 2750 30595 2755
rect 30565 2730 30570 2750
rect 30570 2730 30590 2750
rect 30590 2730 30595 2750
rect 30565 2725 30595 2730
rect 29795 2455 29825 2485
rect 30070 2480 30100 2485
rect 30070 2460 30075 2480
rect 30075 2460 30095 2480
rect 30095 2460 30100 2480
rect 30070 2455 30100 2460
rect 30180 2480 30210 2485
rect 30180 2460 30185 2480
rect 30185 2460 30205 2480
rect 30205 2460 30210 2480
rect 30180 2455 30210 2460
rect 30290 2480 30320 2485
rect 30290 2460 30295 2480
rect 30295 2460 30315 2480
rect 30315 2460 30320 2480
rect 30290 2455 30320 2460
rect 30400 2480 30430 2485
rect 30400 2460 30405 2480
rect 30405 2460 30425 2480
rect 30425 2460 30430 2480
rect 30400 2455 30430 2460
rect 30510 2480 30540 2485
rect 30510 2460 30515 2480
rect 30515 2460 30535 2480
rect 30535 2460 30540 2480
rect 30510 2455 30540 2460
rect 29320 2230 29350 2260
rect 29740 2105 29770 2110
rect 29740 2085 29745 2105
rect 29745 2085 29765 2105
rect 29765 2085 29770 2105
rect 29740 2080 29770 2085
rect 29470 1980 29505 1985
rect 29470 1955 29475 1980
rect 29475 1955 29500 1980
rect 29500 1955 29505 1980
rect 29470 1950 29505 1955
rect 29530 1980 29565 1985
rect 29530 1955 29535 1980
rect 29535 1955 29560 1980
rect 29560 1955 29565 1980
rect 29530 1950 29565 1955
rect 29590 1980 29625 1985
rect 29590 1955 29595 1980
rect 29595 1955 29620 1980
rect 29620 1955 29625 1980
rect 29590 1950 29625 1955
rect 30455 2345 30485 2375
rect 30745 2345 30775 2375
rect 29840 2265 29870 2295
rect 30070 2290 30100 2295
rect 30070 2270 30075 2290
rect 30075 2270 30095 2290
rect 30095 2270 30100 2290
rect 30070 2265 30100 2270
rect 30180 2290 30210 2295
rect 30180 2270 30185 2290
rect 30185 2270 30205 2290
rect 30205 2270 30210 2290
rect 30180 2265 30210 2270
rect 30290 2290 30320 2295
rect 30290 2270 30295 2290
rect 30295 2270 30315 2290
rect 30315 2270 30320 2290
rect 30290 2265 30320 2270
rect 30400 2290 30430 2295
rect 30400 2270 30405 2290
rect 30405 2270 30425 2290
rect 30425 2270 30430 2290
rect 30400 2265 30430 2270
rect 30510 2290 30540 2295
rect 30510 2270 30515 2290
rect 30515 2270 30535 2290
rect 30535 2270 30540 2290
rect 30510 2265 30540 2270
rect 29650 1980 29685 1985
rect 29650 1955 29655 1980
rect 29655 1955 29680 1980
rect 29680 1955 29685 1980
rect 29650 1950 29685 1955
rect 29795 1950 29825 1980
rect 29890 2105 29920 2110
rect 29890 2085 29895 2105
rect 29895 2085 29915 2105
rect 29915 2085 29920 2105
rect 29890 2080 29920 2085
rect 32265 4725 32295 4730
rect 32265 4705 32270 4725
rect 32270 4705 32290 4725
rect 32290 4705 32295 4725
rect 32265 4700 32295 4705
rect 32385 4725 32415 4730
rect 32385 4705 32390 4725
rect 32390 4705 32410 4725
rect 32410 4705 32415 4725
rect 32385 4700 32415 4705
rect 32505 4725 32535 4730
rect 32505 4705 32510 4725
rect 32510 4705 32530 4725
rect 32530 4705 32535 4725
rect 32505 4700 32535 4705
rect 32625 4725 32655 4730
rect 32625 4705 32630 4725
rect 32630 4705 32650 4725
rect 32650 4705 32655 4725
rect 32625 4700 32655 4705
rect 31060 4515 31090 4545
rect 31315 4515 31345 4545
rect 32325 4515 32355 4545
rect 31005 3155 31035 3185
rect 31255 4435 31285 4440
rect 31255 4415 31260 4435
rect 31260 4415 31280 4435
rect 31280 4415 31285 4435
rect 31255 4410 31285 4415
rect 31365 4435 31395 4440
rect 31365 4415 31370 4435
rect 31370 4415 31390 4435
rect 31390 4415 31395 4435
rect 31365 4410 31395 4415
rect 31475 4435 31505 4440
rect 31475 4415 31480 4435
rect 31480 4415 31500 4435
rect 31500 4415 31505 4435
rect 31475 4410 31505 4415
rect 31585 4435 31615 4440
rect 31585 4415 31590 4435
rect 31590 4415 31610 4435
rect 31610 4415 31615 4435
rect 31585 4410 31615 4415
rect 31695 4435 31725 4440
rect 31695 4415 31700 4435
rect 31700 4415 31720 4435
rect 31720 4415 31725 4435
rect 31695 4410 31725 4415
rect 31805 4435 31835 4440
rect 31805 4415 31810 4435
rect 31810 4415 31830 4435
rect 31830 4415 31835 4435
rect 31805 4410 31835 4415
rect 31915 4435 31945 4440
rect 31915 4415 31920 4435
rect 31920 4415 31940 4435
rect 31940 4415 31945 4435
rect 31915 4410 31945 4415
rect 32025 4435 32055 4440
rect 32025 4415 32030 4435
rect 32030 4415 32050 4435
rect 32050 4415 32055 4435
rect 32025 4410 32055 4415
rect 32135 4435 32165 4440
rect 32135 4415 32140 4435
rect 32140 4415 32160 4435
rect 32160 4415 32165 4435
rect 32135 4410 32165 4415
rect 32245 4435 32275 4440
rect 32245 4415 32250 4435
rect 32250 4415 32270 4435
rect 32270 4415 32275 4435
rect 32245 4410 32275 4415
rect 32355 4435 32385 4440
rect 32355 4415 32360 4435
rect 32360 4415 32380 4435
rect 32380 4415 32385 4435
rect 32355 4410 32385 4415
rect 32465 4435 32495 4440
rect 32465 4415 32470 4435
rect 32470 4415 32490 4435
rect 32490 4415 32495 4435
rect 32465 4410 32495 4415
rect 31310 4315 31340 4320
rect 31310 4295 31315 4315
rect 31315 4295 31335 4315
rect 31335 4295 31340 4315
rect 31310 4290 31340 4295
rect 31530 4315 31560 4320
rect 31530 4295 31535 4315
rect 31535 4295 31555 4315
rect 31555 4295 31560 4315
rect 31530 4290 31560 4295
rect 31750 4315 31780 4320
rect 31750 4295 31755 4315
rect 31755 4295 31775 4315
rect 31775 4295 31780 4315
rect 31750 4290 31780 4295
rect 31970 4315 32000 4320
rect 31970 4295 31975 4315
rect 31975 4295 31995 4315
rect 31995 4295 32000 4315
rect 31970 4290 32000 4295
rect 32190 4315 32220 4320
rect 32190 4295 32195 4315
rect 32195 4295 32215 4315
rect 32215 4295 32220 4315
rect 32190 4290 32220 4295
rect 32410 4315 32440 4320
rect 32410 4295 32415 4315
rect 32415 4295 32435 4315
rect 32435 4295 32440 4315
rect 32410 4290 32440 4295
rect 31325 4060 31355 4090
rect 31425 4175 31455 4205
rect 31640 4175 31670 4205
rect 31860 4175 31890 4205
rect 32080 4175 32110 4205
rect 32300 4175 32330 4205
rect 31425 4060 31455 4090
rect 31535 4060 31565 4090
rect 31645 4060 31675 4090
rect 31755 4060 31785 4090
rect 32055 4060 32085 4090
rect 32155 4060 32185 4090
rect 32265 4060 32295 4090
rect 32375 4060 32405 4090
rect 32485 4060 32515 4090
rect 31282 4025 31308 4029
rect 31282 4005 31285 4025
rect 31285 4005 31305 4025
rect 31305 4005 31308 4025
rect 31282 4001 31308 4005
rect 31482 4025 31508 4029
rect 31482 4005 31485 4025
rect 31485 4005 31505 4025
rect 31505 4005 31508 4025
rect 31482 4001 31508 4005
rect 31700 4025 31730 4030
rect 31700 4005 31705 4025
rect 31705 4005 31725 4025
rect 31725 4005 31730 4025
rect 31700 4000 31730 4005
rect 32010 4025 32036 4029
rect 32010 4005 32013 4025
rect 32013 4005 32033 4025
rect 32033 4005 32036 4025
rect 32010 4001 32036 4005
rect 32210 4025 32240 4030
rect 32210 4005 32215 4025
rect 32215 4005 32235 4025
rect 32235 4005 32240 4025
rect 32210 4000 32240 4005
rect 32430 4025 32460 4030
rect 32430 4005 32435 4025
rect 32435 4005 32455 4025
rect 32455 4005 32460 4025
rect 32430 4000 32460 4005
rect 32875 4000 32905 4030
rect 31145 3965 31175 3970
rect 31145 3945 31150 3965
rect 31150 3945 31170 3965
rect 31170 3945 31175 3965
rect 31145 3940 31175 3945
rect 31410 3905 31436 3910
rect 31410 3885 31413 3905
rect 31413 3885 31430 3905
rect 31430 3885 31436 3905
rect 31410 3880 31436 3885
rect 31630 3905 31656 3910
rect 31630 3885 31633 3905
rect 31633 3885 31650 3905
rect 31650 3885 31656 3905
rect 31630 3880 31656 3885
rect 31774 3905 31800 3910
rect 31774 3885 31780 3905
rect 31780 3885 31797 3905
rect 31797 3885 31800 3905
rect 31774 3880 31800 3885
rect 32140 3905 32166 3910
rect 32140 3885 32143 3905
rect 32143 3885 32160 3905
rect 32160 3885 32166 3905
rect 32140 3880 32166 3885
rect 32360 3905 32386 3910
rect 32360 3885 32363 3905
rect 32363 3885 32380 3905
rect 32380 3885 32386 3905
rect 32360 3880 32386 3885
rect 32504 3905 32530 3910
rect 32504 3885 32510 3905
rect 32510 3885 32527 3905
rect 32527 3885 32530 3905
rect 32504 3880 32530 3885
rect 31260 3820 31290 3850
rect 31365 3820 31395 3850
rect 31480 3820 31510 3850
rect 31585 3820 31615 3850
rect 31700 3820 31730 3850
rect 31815 3820 31845 3850
rect 31990 3820 32020 3850
rect 32210 3820 32240 3850
rect 32430 3820 32460 3850
rect 32085 3730 32115 3760
rect 32305 3730 32335 3760
rect 32545 3730 32575 3760
rect 31885 3695 31915 3725
rect 31885 3660 31915 3665
rect 31885 3640 31890 3660
rect 31890 3640 31910 3660
rect 31910 3640 31915 3660
rect 31885 3635 31915 3640
rect 31345 3600 31375 3605
rect 31345 3580 31350 3600
rect 31350 3580 31370 3600
rect 31370 3580 31375 3600
rect 31345 3575 31375 3580
rect 31465 3600 31495 3605
rect 31465 3580 31470 3600
rect 31470 3580 31490 3600
rect 31490 3580 31495 3600
rect 31465 3575 31495 3580
rect 31585 3600 31615 3605
rect 31585 3580 31590 3600
rect 31590 3580 31610 3600
rect 31610 3580 31615 3600
rect 31585 3575 31615 3580
rect 31705 3600 31735 3605
rect 31705 3580 31710 3600
rect 31710 3580 31730 3600
rect 31730 3580 31735 3600
rect 31705 3575 31735 3580
rect 31825 3600 31855 3605
rect 31825 3580 31830 3600
rect 31830 3580 31850 3600
rect 31850 3580 31855 3600
rect 31825 3575 31855 3580
rect 31885 3600 31915 3605
rect 31885 3580 31890 3600
rect 31890 3580 31910 3600
rect 31910 3580 31915 3600
rect 31885 3575 31915 3580
rect 31945 3600 31975 3605
rect 31945 3580 31950 3600
rect 31950 3580 31970 3600
rect 31970 3580 31975 3600
rect 31945 3575 31975 3580
rect 32065 3600 32095 3605
rect 32065 3580 32070 3600
rect 32070 3580 32090 3600
rect 32090 3580 32095 3600
rect 32065 3575 32095 3580
rect 32185 3600 32215 3605
rect 32185 3580 32190 3600
rect 32190 3580 32210 3600
rect 32210 3580 32215 3600
rect 32185 3575 32215 3580
rect 32305 3600 32335 3605
rect 32305 3580 32310 3600
rect 32310 3580 32330 3600
rect 32330 3580 32335 3600
rect 32305 3575 32335 3580
rect 32425 3600 32455 3605
rect 32425 3580 32430 3600
rect 32430 3580 32450 3600
rect 32450 3580 32455 3600
rect 32425 3575 32455 3580
rect 31826 3180 31854 3185
rect 31826 3160 31831 3180
rect 31831 3160 31849 3180
rect 31849 3160 31854 3180
rect 31826 3155 31854 3160
rect 31285 3100 31315 3130
rect 31060 2960 31090 2990
rect 31525 3100 31555 3130
rect 31765 3100 31795 3130
rect 32005 3100 32035 3130
rect 32245 3100 32275 3130
rect 32485 3100 32515 3130
rect 31405 3015 31435 3045
rect 31645 3015 31675 3045
rect 31885 3015 31915 3045
rect 32125 3015 32155 3045
rect 32365 3015 32395 3045
rect 31885 2960 31915 2990
rect 31130 2890 31160 2895
rect 31130 2870 31135 2890
rect 31135 2870 31155 2890
rect 31155 2870 31160 2890
rect 31130 2865 31160 2870
rect 31250 2890 31280 2895
rect 31250 2870 31255 2890
rect 31255 2870 31275 2890
rect 31275 2870 31280 2890
rect 31250 2865 31280 2870
rect 31370 2890 31400 2895
rect 31370 2870 31375 2890
rect 31375 2870 31395 2890
rect 31395 2870 31400 2890
rect 31370 2865 31400 2870
rect 31490 2890 31520 2895
rect 31490 2870 31495 2890
rect 31495 2870 31515 2890
rect 31515 2870 31520 2890
rect 31490 2865 31520 2870
rect 31610 2890 31640 2895
rect 31610 2870 31615 2890
rect 31615 2870 31635 2890
rect 31635 2870 31640 2890
rect 31610 2865 31640 2870
rect 31070 2470 31100 2475
rect 31070 2450 31075 2470
rect 31075 2450 31095 2470
rect 31095 2450 31100 2470
rect 31070 2445 31100 2450
rect 31190 2470 31220 2475
rect 31190 2450 31195 2470
rect 31195 2450 31215 2470
rect 31215 2450 31220 2470
rect 31190 2445 31220 2450
rect 31310 2470 31340 2475
rect 31310 2450 31315 2470
rect 31315 2450 31335 2470
rect 31335 2450 31340 2470
rect 31310 2445 31340 2450
rect 31430 2470 31460 2475
rect 31430 2450 31435 2470
rect 31435 2450 31455 2470
rect 31455 2450 31460 2470
rect 31430 2445 31460 2450
rect 31550 2470 31580 2475
rect 31550 2450 31555 2470
rect 31555 2450 31575 2470
rect 31575 2450 31580 2470
rect 31550 2445 31580 2450
rect 31670 2470 31700 2475
rect 31670 2450 31675 2470
rect 31675 2450 31695 2470
rect 31695 2450 31700 2470
rect 31670 2445 31700 2450
rect 31370 2390 31400 2420
rect 32160 2890 32190 2895
rect 32160 2870 32165 2890
rect 32165 2870 32185 2890
rect 32185 2870 32190 2890
rect 32160 2865 32190 2870
rect 32280 2890 32310 2895
rect 32280 2870 32285 2890
rect 32285 2870 32305 2890
rect 32305 2870 32310 2890
rect 32280 2865 32310 2870
rect 32400 2890 32430 2895
rect 32400 2870 32405 2890
rect 32405 2870 32425 2890
rect 32425 2870 32430 2890
rect 32400 2865 32430 2870
rect 32520 2890 32550 2895
rect 32520 2870 32525 2890
rect 32525 2870 32545 2890
rect 32545 2870 32550 2890
rect 32520 2865 32550 2870
rect 32640 2890 32670 2895
rect 32640 2870 32645 2890
rect 32645 2870 32665 2890
rect 32665 2870 32670 2890
rect 32640 2865 32670 2870
rect 32100 2470 32130 2475
rect 32100 2450 32105 2470
rect 32105 2450 32125 2470
rect 32125 2450 32130 2470
rect 32100 2445 32130 2450
rect 32220 2470 32250 2475
rect 32220 2450 32225 2470
rect 32225 2450 32245 2470
rect 32245 2450 32250 2470
rect 32220 2445 32250 2450
rect 32340 2470 32370 2475
rect 32340 2450 32345 2470
rect 32345 2450 32365 2470
rect 32365 2450 32370 2470
rect 32340 2445 32370 2450
rect 32460 2470 32490 2475
rect 32460 2450 32465 2470
rect 32465 2450 32485 2470
rect 32485 2450 32490 2470
rect 32460 2445 32490 2450
rect 32580 2470 32610 2475
rect 32580 2450 32585 2470
rect 32585 2450 32605 2470
rect 32605 2450 32610 2470
rect 32580 2445 32610 2450
rect 32700 2470 32730 2475
rect 32700 2450 32705 2470
rect 32705 2450 32725 2470
rect 32725 2450 32730 2470
rect 32700 2445 32730 2450
rect 31885 2390 31915 2420
rect 32400 2390 32430 2420
rect 31675 2345 31705 2375
rect 32095 2345 32125 2375
rect 30880 2300 30910 2330
rect 30835 2200 30865 2230
rect 29595 1895 29625 1925
rect 29840 1895 29870 1925
rect 30015 1920 30045 1925
rect 30015 1900 30020 1920
rect 30020 1900 30038 1920
rect 30038 1900 30045 1920
rect 30015 1895 30045 1900
rect 30125 1920 30155 1925
rect 30125 1900 30130 1920
rect 30130 1900 30148 1920
rect 30148 1900 30155 1920
rect 30125 1895 30155 1900
rect 30235 1920 30265 1925
rect 30235 1900 30240 1920
rect 30240 1900 30258 1920
rect 30258 1900 30265 1920
rect 30235 1895 30265 1900
rect 30345 1920 30375 1925
rect 30345 1900 30350 1920
rect 30350 1900 30368 1920
rect 30368 1900 30375 1920
rect 30345 1895 30375 1900
rect 30455 1920 30485 1925
rect 30455 1900 30460 1920
rect 30460 1900 30478 1920
rect 30478 1900 30485 1920
rect 30455 1895 30485 1900
rect 30565 1920 30595 1925
rect 30565 1900 30570 1920
rect 30570 1900 30588 1920
rect 30588 1900 30595 1920
rect 30565 1895 30595 1900
rect 30790 1895 30820 1925
rect 29475 1790 29505 1820
rect 29730 1730 29760 1760
rect 30440 1730 30470 1760
rect 30745 1730 30775 1760
rect 29320 1675 29350 1705
rect 29795 1675 29825 1705
rect 30140 1700 30170 1705
rect 30140 1680 30145 1700
rect 30145 1680 30165 1700
rect 30165 1680 30170 1700
rect 30140 1675 30170 1680
rect 30340 1700 30370 1705
rect 30340 1680 30345 1700
rect 30345 1680 30365 1700
rect 30365 1680 30370 1700
rect 30340 1675 30370 1680
rect 30540 1700 30570 1705
rect 30540 1680 30545 1700
rect 30545 1680 30565 1700
rect 30565 1680 30570 1700
rect 30540 1675 30570 1680
rect 29730 1640 29765 1645
rect 29730 1615 29735 1640
rect 29735 1615 29760 1640
rect 29760 1615 29765 1640
rect 29730 1610 29765 1615
rect 29790 1640 29825 1645
rect 29790 1615 29795 1640
rect 29795 1615 29820 1640
rect 29820 1615 29825 1640
rect 29790 1610 29825 1615
rect 30790 1620 30820 1650
rect 30745 1405 30775 1435
rect 29880 1315 29910 1320
rect 29880 1295 29885 1315
rect 29885 1295 29905 1315
rect 29905 1295 29910 1315
rect 29880 1290 29910 1295
rect 29970 1315 30000 1320
rect 29970 1295 29975 1315
rect 29975 1295 29995 1315
rect 29995 1295 30000 1315
rect 29970 1290 30000 1295
rect 30240 930 30270 935
rect 30240 910 30245 930
rect 30245 910 30265 930
rect 30265 910 30270 930
rect 30240 905 30270 910
rect 30340 905 30370 935
rect 30440 930 30470 935
rect 30440 910 30445 930
rect 30445 910 30465 930
rect 30465 910 30470 930
rect 30440 905 30470 910
rect 30790 905 30820 935
rect 30340 870 30370 875
rect 30340 850 30345 870
rect 30345 850 30365 870
rect 30365 850 30370 870
rect 30340 845 30370 850
rect 30790 830 30820 860
rect 32965 3820 32995 3850
rect 32920 3730 32950 3760
rect 32875 2300 32905 2330
rect 31245 2255 31275 2285
rect 31355 2255 31385 2285
rect 31465 2255 31495 2285
rect 31575 2255 31605 2285
rect 31685 2255 31715 2285
rect 31795 2255 31825 2285
rect 31975 2255 32005 2285
rect 32085 2255 32115 2285
rect 32195 2255 32225 2285
rect 32305 2255 32335 2285
rect 32415 2255 32445 2285
rect 32525 2255 32555 2285
rect 31520 2225 31550 2230
rect 31520 2205 31525 2225
rect 31525 2205 31545 2225
rect 31545 2205 31550 2225
rect 31520 2200 31550 2205
rect 32250 2225 32280 2230
rect 32250 2205 32255 2225
rect 32255 2205 32275 2225
rect 32275 2205 32280 2225
rect 32250 2200 32280 2205
rect 31300 1920 31330 1950
rect 31410 1920 31440 1950
rect 31520 1920 31550 1950
rect 31630 1920 31660 1950
rect 31740 1920 31770 1950
rect 32030 1920 32060 1950
rect 32140 1920 32170 1950
rect 32250 1920 32280 1950
rect 32360 1920 32390 1950
rect 32470 1920 32500 1950
rect 31195 1865 31225 1895
rect 31415 1865 31445 1895
rect 30880 1790 30910 1820
rect 31090 1775 31120 1805
rect 31310 1775 31340 1805
rect 31240 1755 31266 1760
rect 31240 1735 31243 1755
rect 31243 1735 31260 1755
rect 31260 1735 31266 1755
rect 31240 1730 31266 1735
rect 31645 1865 31675 1895
rect 31530 1775 31560 1805
rect 31460 1755 31486 1760
rect 31460 1735 31463 1755
rect 31463 1735 31480 1755
rect 31480 1735 31486 1755
rect 31460 1730 31486 1735
rect 31604 1755 31630 1760
rect 31604 1735 31610 1755
rect 31610 1735 31627 1755
rect 31627 1735 31630 1755
rect 31604 1730 31630 1735
rect 31825 1820 31855 1850
rect 32235 1865 32265 1895
rect 32455 1865 32485 1895
rect 32685 1865 32715 1895
rect 31945 1820 31975 1850
rect 32130 1775 32160 1805
rect 31870 1755 31896 1760
rect 31870 1735 31873 1755
rect 31873 1735 31890 1755
rect 31890 1735 31896 1755
rect 31870 1730 31896 1735
rect 32350 1775 32380 1805
rect 32280 1755 32306 1760
rect 32280 1735 32283 1755
rect 32283 1735 32300 1755
rect 32300 1735 32306 1755
rect 32280 1730 32306 1735
rect 32570 1775 32600 1805
rect 32500 1755 32526 1760
rect 32500 1735 32503 1755
rect 32503 1735 32520 1755
rect 32520 1735 32526 1755
rect 32500 1730 32526 1735
rect 32644 1755 32670 1760
rect 32644 1735 32650 1755
rect 32650 1735 32667 1755
rect 32667 1735 32670 1755
rect 32644 1730 32670 1735
rect 32875 1795 32905 1825
rect 30945 1645 30975 1650
rect 30945 1625 30950 1645
rect 30950 1625 30970 1645
rect 30970 1625 30975 1645
rect 30945 1620 30975 1625
rect 31109 1535 31135 1540
rect 31109 1515 31112 1535
rect 31112 1515 31129 1535
rect 31129 1515 31135 1535
rect 31109 1510 31135 1515
rect 31310 1535 31340 1540
rect 31310 1515 31315 1535
rect 31315 1515 31335 1535
rect 31335 1515 31340 1535
rect 31310 1510 31340 1515
rect 31530 1535 31560 1540
rect 31530 1515 31535 1535
rect 31535 1515 31555 1535
rect 31555 1515 31560 1535
rect 31530 1510 31560 1515
rect 31925 1535 31951 1540
rect 31925 1515 31928 1535
rect 31928 1515 31945 1535
rect 31945 1515 31951 1535
rect 31925 1510 31951 1515
rect 32149 1535 32175 1540
rect 32149 1515 32152 1535
rect 32152 1515 32169 1535
rect 32169 1515 32175 1535
rect 32149 1510 32175 1515
rect 32350 1535 32380 1540
rect 32350 1515 32355 1535
rect 32355 1515 32375 1535
rect 32375 1515 32380 1535
rect 32350 1510 32380 1515
rect 32570 1535 32600 1540
rect 32570 1515 32575 1535
rect 32575 1515 32595 1535
rect 32595 1515 32600 1535
rect 32570 1510 32600 1515
rect 31150 1450 31180 1480
rect 31255 1450 31285 1480
rect 31365 1450 31395 1480
rect 31475 1450 31505 1480
rect 31585 1450 31615 1480
rect 31010 1360 31040 1390
rect 31760 1360 31790 1390
rect 31320 1315 31350 1345
rect 32190 1450 32220 1480
rect 32295 1450 32325 1480
rect 32405 1450 32435 1480
rect 32515 1450 32545 1480
rect 32625 1450 32655 1480
rect 31875 1315 31905 1345
rect 32380 1335 32410 1365
rect 32920 1335 32950 1365
rect 31430 1250 31460 1255
rect 31430 1230 31435 1250
rect 31435 1230 31455 1250
rect 31455 1230 31460 1250
rect 31430 1225 31460 1230
rect 31540 1250 31570 1255
rect 31540 1230 31545 1250
rect 31545 1230 31565 1250
rect 31565 1230 31570 1250
rect 31540 1225 31570 1230
rect 31650 1250 31680 1255
rect 31650 1230 31655 1250
rect 31655 1230 31675 1250
rect 31675 1230 31680 1250
rect 31650 1225 31680 1230
rect 31760 1250 31790 1255
rect 31760 1230 31765 1250
rect 31765 1230 31785 1250
rect 31785 1230 31790 1250
rect 31760 1225 31790 1230
rect 31870 1250 31900 1255
rect 31870 1230 31875 1250
rect 31875 1230 31895 1250
rect 31895 1230 31900 1250
rect 31870 1225 31900 1230
rect 31980 1250 32010 1255
rect 31980 1230 31985 1250
rect 31985 1230 32005 1250
rect 32005 1230 32010 1250
rect 31980 1225 32010 1230
rect 32090 1250 32120 1255
rect 32090 1230 32095 1250
rect 32095 1230 32115 1250
rect 32115 1230 32120 1250
rect 32090 1225 32120 1230
rect 32200 1250 32230 1255
rect 32200 1230 32205 1250
rect 32205 1230 32225 1250
rect 32225 1230 32230 1250
rect 32200 1225 32230 1230
rect 32310 1250 32340 1255
rect 32310 1230 32315 1250
rect 32315 1230 32335 1250
rect 32335 1230 32340 1250
rect 32310 1225 32340 1230
rect 32435 1250 32465 1255
rect 32435 1230 32440 1250
rect 32440 1230 32460 1250
rect 32460 1230 32465 1250
rect 32435 1225 32465 1230
rect 31200 930 31230 935
rect 31200 910 31205 930
rect 31205 910 31225 930
rect 31225 910 31230 930
rect 31200 905 31230 910
rect 31265 930 31295 935
rect 31265 910 31270 930
rect 31270 910 31290 930
rect 31290 910 31295 930
rect 31265 905 31295 910
rect 31375 930 31405 935
rect 31375 910 31380 930
rect 31380 910 31400 930
rect 31400 910 31405 930
rect 31375 905 31405 910
rect 31485 930 31515 935
rect 31485 910 31490 930
rect 31490 910 31510 930
rect 31510 910 31515 930
rect 31485 905 31515 910
rect 31595 930 31625 935
rect 31595 910 31600 930
rect 31600 910 31620 930
rect 31620 910 31625 930
rect 31595 905 31625 910
rect 31705 930 31735 935
rect 31705 910 31710 930
rect 31710 910 31730 930
rect 31730 910 31735 930
rect 31705 905 31735 910
rect 31815 930 31845 935
rect 31815 910 31820 930
rect 31820 910 31840 930
rect 31840 910 31845 930
rect 31815 905 31845 910
rect 31925 930 31955 935
rect 31925 910 31930 930
rect 31930 910 31950 930
rect 31950 910 31955 930
rect 31925 905 31955 910
rect 32035 930 32065 935
rect 32035 910 32040 930
rect 32040 910 32060 930
rect 32060 910 32065 930
rect 32035 905 32065 910
rect 32145 930 32175 935
rect 32145 910 32150 930
rect 32150 910 32170 930
rect 32170 910 32175 930
rect 32145 905 32175 910
rect 32255 930 32285 935
rect 32255 910 32260 930
rect 32260 910 32280 930
rect 32280 910 32285 930
rect 32255 905 32285 910
rect 32365 930 32395 935
rect 32365 910 32370 930
rect 32370 910 32390 930
rect 32390 910 32395 930
rect 32365 905 32395 910
rect 32480 930 32510 935
rect 32480 910 32485 930
rect 32485 910 32505 930
rect 32505 910 32510 930
rect 32480 905 32510 910
rect 31010 810 31040 840
rect 31510 810 31540 840
rect 31940 810 31970 840
rect 32160 810 32190 840
rect 32380 810 32410 840
rect 30835 710 30865 740
rect 31310 735 31340 740
rect 31310 715 31315 735
rect 31315 715 31335 735
rect 31335 715 31340 735
rect 31310 710 31340 715
rect 31380 735 31410 740
rect 31380 715 31385 735
rect 31385 715 31405 735
rect 31405 715 31410 735
rect 31380 710 31410 715
rect 31450 735 31480 740
rect 31450 715 31455 735
rect 31455 715 31475 735
rect 31475 715 31480 735
rect 31450 710 31480 715
rect 33010 3685 33040 3715
rect 33150 3710 33180 3715
rect 33150 3690 33155 3710
rect 33155 3690 33175 3710
rect 33175 3690 33180 3710
rect 33150 3685 33180 3690
rect 33260 3710 33290 3715
rect 33260 3690 33265 3710
rect 33265 3690 33285 3710
rect 33285 3690 33290 3710
rect 33260 3685 33290 3690
rect 33370 3710 33400 3715
rect 33370 3690 33375 3710
rect 33375 3690 33395 3710
rect 33395 3690 33400 3710
rect 33370 3685 33400 3690
rect 33480 3710 33510 3715
rect 33480 3690 33485 3710
rect 33485 3690 33505 3710
rect 33505 3690 33510 3710
rect 33480 3685 33510 3690
rect 33590 3710 33620 3715
rect 33590 3690 33595 3710
rect 33595 3690 33615 3710
rect 33615 3690 33620 3710
rect 33590 3685 33620 3690
rect 33700 3710 33730 3715
rect 33700 3690 33705 3710
rect 33705 3690 33725 3710
rect 33725 3690 33730 3710
rect 33700 3685 33730 3690
rect 33810 3710 33840 3715
rect 33810 3690 33815 3710
rect 33815 3690 33835 3710
rect 33835 3690 33840 3710
rect 33810 3685 33840 3690
rect 34160 3705 34190 3735
rect 34111 3625 34141 3655
rect 34160 3625 34190 3655
rect 34210 3625 34240 3655
rect 33205 3040 33235 3045
rect 33205 3020 33210 3040
rect 33210 3020 33230 3040
rect 33230 3020 33235 3040
rect 33205 3015 33235 3020
rect 33315 3040 33345 3045
rect 33315 3020 33320 3040
rect 33320 3020 33340 3040
rect 33340 3020 33345 3040
rect 33315 3015 33345 3020
rect 33425 3040 33455 3045
rect 33425 3020 33430 3040
rect 33430 3020 33450 3040
rect 33450 3020 33455 3040
rect 33425 3015 33455 3020
rect 33535 3040 33565 3045
rect 33535 3020 33540 3040
rect 33540 3020 33560 3040
rect 33560 3020 33565 3040
rect 33535 3015 33565 3020
rect 33645 3040 33675 3045
rect 33645 3020 33650 3040
rect 33650 3020 33670 3040
rect 33670 3020 33675 3040
rect 33645 3015 33675 3020
rect 33755 3040 33785 3045
rect 33755 3020 33760 3040
rect 33760 3020 33780 3040
rect 33780 3020 33785 3040
rect 33755 3015 33785 3020
rect 34111 3020 34141 3050
rect 34160 3020 34190 3050
rect 34210 3020 34240 3050
rect 33045 2905 33075 2935
rect 33315 2860 33345 2890
rect 33590 2905 33620 2935
rect 34160 2905 34190 2935
rect 33205 2750 33235 2755
rect 33205 2730 33210 2750
rect 33210 2730 33230 2750
rect 33230 2730 33235 2750
rect 33205 2725 33235 2730
rect 33315 2750 33345 2755
rect 33315 2730 33320 2750
rect 33320 2730 33340 2750
rect 33340 2730 33345 2750
rect 33315 2725 33345 2730
rect 33425 2750 33455 2755
rect 33425 2730 33430 2750
rect 33430 2730 33450 2750
rect 33450 2730 33455 2750
rect 33425 2725 33455 2730
rect 33535 2750 33565 2755
rect 33535 2730 33540 2750
rect 33540 2730 33560 2750
rect 33560 2730 33565 2750
rect 33535 2725 33565 2730
rect 33645 2750 33675 2755
rect 33645 2730 33650 2750
rect 33650 2730 33670 2750
rect 33670 2730 33675 2750
rect 33645 2725 33675 2730
rect 33755 2750 33785 2755
rect 33755 2730 33760 2750
rect 33760 2730 33780 2750
rect 33780 2730 33785 2750
rect 33755 2725 33785 2730
rect 34450 2860 34480 2890
rect 33260 2480 33290 2485
rect 33260 2460 33265 2480
rect 33265 2460 33285 2480
rect 33285 2460 33290 2480
rect 33260 2455 33290 2460
rect 33370 2480 33400 2485
rect 33370 2460 33375 2480
rect 33375 2460 33395 2480
rect 33395 2460 33400 2480
rect 33370 2455 33400 2460
rect 33480 2480 33510 2485
rect 33480 2460 33485 2480
rect 33485 2460 33505 2480
rect 33505 2460 33510 2480
rect 33480 2455 33510 2460
rect 33590 2480 33620 2485
rect 33590 2460 33595 2480
rect 33595 2460 33615 2480
rect 33615 2460 33620 2480
rect 33590 2455 33620 2460
rect 33700 2480 33730 2485
rect 33700 2460 33705 2480
rect 33705 2460 33725 2480
rect 33725 2460 33730 2480
rect 33700 2455 33730 2460
rect 33980 2455 34010 2485
rect 33045 2345 33075 2375
rect 33315 2345 33345 2375
rect 33260 2290 33290 2295
rect 33260 2270 33265 2290
rect 33265 2270 33285 2290
rect 33285 2270 33290 2290
rect 33260 2265 33290 2270
rect 33370 2290 33400 2295
rect 33370 2270 33375 2290
rect 33375 2270 33395 2290
rect 33395 2270 33400 2290
rect 33370 2265 33400 2270
rect 33480 2290 33510 2295
rect 33480 2270 33485 2290
rect 33485 2270 33505 2290
rect 33505 2270 33510 2290
rect 33480 2265 33510 2270
rect 33590 2290 33620 2295
rect 33590 2270 33595 2290
rect 33595 2270 33615 2290
rect 33615 2270 33620 2290
rect 33590 2265 33620 2270
rect 33700 2290 33730 2295
rect 33700 2270 33705 2290
rect 33705 2270 33725 2290
rect 33725 2270 33730 2290
rect 33700 2265 33730 2270
rect 33935 2265 33965 2295
rect 33880 2105 33910 2110
rect 33880 2085 33885 2105
rect 33885 2085 33905 2105
rect 33905 2085 33910 2105
rect 33880 2080 33910 2085
rect 34500 2725 34530 2755
rect 34450 2230 34480 2260
rect 34030 2105 34060 2110
rect 34030 2085 34035 2105
rect 34035 2085 34055 2105
rect 34055 2085 34060 2105
rect 34030 2080 34060 2085
rect 33980 1950 34010 1980
rect 34115 1980 34150 1985
rect 34115 1955 34120 1980
rect 34120 1955 34145 1980
rect 34145 1955 34150 1980
rect 34115 1950 34150 1955
rect 34175 1980 34210 1985
rect 34175 1955 34180 1980
rect 34180 1955 34205 1980
rect 34205 1955 34210 1980
rect 34175 1950 34210 1955
rect 34235 1980 34270 1985
rect 34235 1955 34240 1980
rect 34240 1955 34265 1980
rect 34265 1955 34270 1980
rect 34235 1950 34270 1955
rect 34295 1980 34330 1985
rect 34295 1955 34300 1980
rect 34300 1955 34325 1980
rect 34325 1955 34330 1980
rect 34295 1950 34330 1955
rect 33010 1895 33040 1925
rect 33205 1920 33235 1925
rect 33205 1900 33212 1920
rect 33212 1900 33230 1920
rect 33230 1900 33235 1920
rect 33205 1895 33235 1900
rect 33315 1920 33345 1925
rect 33315 1900 33322 1920
rect 33322 1900 33340 1920
rect 33340 1900 33345 1920
rect 33315 1895 33345 1900
rect 33425 1920 33455 1925
rect 33425 1900 33432 1920
rect 33432 1900 33450 1920
rect 33450 1900 33455 1920
rect 33425 1895 33455 1900
rect 33535 1920 33565 1925
rect 33535 1900 33542 1920
rect 33542 1900 33560 1920
rect 33560 1900 33565 1920
rect 33535 1895 33565 1900
rect 33645 1920 33675 1925
rect 33645 1900 33652 1920
rect 33652 1900 33670 1920
rect 33670 1900 33675 1920
rect 33645 1895 33675 1900
rect 33755 1920 33785 1925
rect 33755 1900 33762 1920
rect 33762 1900 33780 1920
rect 33780 1900 33785 1920
rect 33755 1895 33785 1900
rect 33935 1895 33965 1925
rect 34175 1895 34205 1925
rect 34295 1795 34325 1825
rect 33020 1730 33050 1760
rect 33330 1730 33360 1760
rect 34040 1730 34070 1760
rect 33230 1700 33260 1705
rect 33230 1680 33235 1700
rect 33235 1680 33255 1700
rect 33255 1680 33260 1700
rect 33230 1675 33260 1680
rect 33430 1700 33460 1705
rect 33430 1680 33435 1700
rect 33435 1680 33455 1700
rect 33455 1680 33460 1700
rect 33430 1675 33460 1680
rect 33630 1700 33660 1705
rect 33630 1680 33635 1700
rect 33635 1680 33655 1700
rect 33655 1680 33660 1700
rect 33630 1675 33660 1680
rect 33975 1675 34005 1705
rect 34450 1675 34480 1705
rect 33975 1640 34010 1645
rect 33975 1615 33980 1640
rect 33980 1615 34005 1640
rect 34005 1615 34010 1640
rect 33975 1610 34010 1615
rect 34035 1640 34070 1645
rect 34035 1615 34040 1640
rect 34040 1615 34065 1640
rect 34065 1615 34070 1640
rect 34035 1610 34070 1615
rect 33020 1405 33050 1435
rect 33800 1315 33830 1320
rect 33800 1295 33805 1315
rect 33805 1295 33825 1315
rect 33825 1295 33830 1315
rect 33800 1290 33830 1295
rect 33890 1315 33920 1320
rect 33890 1295 33895 1315
rect 33895 1295 33915 1315
rect 33915 1295 33920 1315
rect 33890 1290 33920 1295
rect 33020 905 33050 935
rect 33330 930 33360 935
rect 33330 910 33335 930
rect 33335 910 33355 930
rect 33355 910 33360 930
rect 33330 905 33360 910
rect 33430 905 33460 935
rect 33530 930 33560 935
rect 33530 910 33535 930
rect 33535 910 33555 930
rect 33555 910 33560 930
rect 33530 905 33560 910
rect 32965 810 32995 840
rect 32050 730 32080 735
rect 32050 710 32055 730
rect 32055 710 32075 730
rect 32075 710 32080 730
rect 32050 705 32080 710
rect 32270 730 32300 735
rect 32270 710 32275 730
rect 32275 710 32295 730
rect 32295 710 32300 730
rect 32270 705 32300 710
rect 32490 730 32520 735
rect 32490 710 32495 730
rect 32495 710 32515 730
rect 32515 710 32520 730
rect 32490 705 32520 710
rect 32920 705 32950 735
rect 31995 610 32025 615
rect 31995 590 32000 610
rect 32000 590 32020 610
rect 32020 590 32025 610
rect 31995 585 32025 590
rect 32105 610 32135 615
rect 32105 590 32110 610
rect 32110 590 32130 610
rect 32130 590 32135 610
rect 32105 585 32135 590
rect 32215 610 32245 615
rect 32215 590 32220 610
rect 32220 590 32240 610
rect 32240 590 32245 610
rect 32215 585 32245 590
rect 32325 610 32355 615
rect 32325 590 32330 610
rect 32330 590 32350 610
rect 32350 590 32355 610
rect 32325 585 32355 590
rect 32435 610 32465 615
rect 32435 590 32440 610
rect 32440 590 32460 610
rect 32460 590 32465 610
rect 32435 585 32465 590
rect 33430 870 33460 875
rect 33430 850 33435 870
rect 33435 850 33455 870
rect 33455 850 33460 870
rect 33430 845 33460 850
rect 29270 465 29300 495
rect 30790 465 30820 495
rect 31380 465 31410 495
rect 32215 465 32245 495
rect 33020 465 33050 495
rect 34500 465 34530 495
rect 30790 -545 30820 -515
<< metal2 >>
rect 30785 6185 30825 6190
rect 30785 6155 30790 6185
rect 30820 6155 30825 6185
rect 30785 6150 30825 6155
rect 31530 4945 31570 4950
rect 31530 4915 31535 4945
rect 31565 4940 31570 4945
rect 31650 4945 31690 4950
rect 31650 4940 31655 4945
rect 31565 4920 31655 4940
rect 31565 4915 31570 4920
rect 31530 4910 31570 4915
rect 31650 4915 31655 4920
rect 31685 4940 31690 4945
rect 31770 4945 31810 4950
rect 31770 4940 31775 4945
rect 31685 4920 31775 4940
rect 31685 4915 31690 4920
rect 31650 4910 31690 4915
rect 31770 4915 31775 4920
rect 31805 4930 31810 4945
rect 32440 4930 32480 4935
rect 31805 4915 32445 4930
rect 31770 4910 32445 4915
rect 32440 4900 32445 4910
rect 32475 4900 32480 4930
rect 32440 4895 32480 4900
rect 31470 4885 31510 4890
rect 31470 4875 31475 4885
rect 30785 4870 30825 4875
rect 30785 4840 30790 4870
rect 30820 4865 30825 4870
rect 31280 4870 31475 4875
rect 31280 4865 31285 4870
rect 30820 4845 31285 4865
rect 30820 4840 30825 4845
rect 30785 4835 30825 4840
rect 31280 4840 31285 4845
rect 31315 4855 31475 4870
rect 31505 4880 31510 4885
rect 31590 4885 31630 4890
rect 31590 4880 31595 4885
rect 31505 4860 31595 4880
rect 31505 4855 31510 4860
rect 31315 4840 31320 4855
rect 31470 4850 31510 4855
rect 31590 4855 31595 4860
rect 31625 4880 31630 4885
rect 31710 4885 31750 4890
rect 31710 4880 31715 4885
rect 31625 4860 31715 4880
rect 31625 4855 31630 4860
rect 31590 4850 31630 4855
rect 31710 4855 31715 4860
rect 31745 4880 31750 4885
rect 31830 4885 31870 4890
rect 31830 4880 31835 4885
rect 31745 4860 31835 4880
rect 31745 4855 31750 4860
rect 31710 4850 31750 4855
rect 31830 4855 31835 4860
rect 31865 4855 31870 4885
rect 31830 4850 31870 4855
rect 32200 4860 32240 4865
rect 31280 4835 31320 4840
rect 32200 4830 32205 4860
rect 32235 4855 32240 4860
rect 32320 4860 32360 4865
rect 32320 4855 32325 4860
rect 32235 4835 32325 4855
rect 32235 4830 32240 4835
rect 32200 4825 32240 4830
rect 32320 4830 32325 4835
rect 32355 4855 32360 4860
rect 32440 4860 32480 4865
rect 32440 4855 32445 4860
rect 32355 4835 32445 4855
rect 32355 4830 32360 4835
rect 32320 4825 32360 4830
rect 32440 4830 32445 4835
rect 32475 4855 32480 4860
rect 32560 4860 32600 4865
rect 32560 4855 32565 4860
rect 32475 4835 32565 4855
rect 32475 4830 32480 4835
rect 32440 4825 32480 4830
rect 32560 4830 32565 4835
rect 32595 4855 32600 4860
rect 32680 4860 32720 4865
rect 32680 4855 32685 4860
rect 32595 4835 32685 4855
rect 32595 4830 32600 4835
rect 32560 4825 32600 4830
rect 32680 4830 32685 4835
rect 32715 4830 32720 4860
rect 32680 4825 32720 4830
rect 31000 4730 31040 4735
rect 31000 4700 31005 4730
rect 31035 4725 31040 4730
rect 31650 4730 31690 4735
rect 31650 4725 31655 4730
rect 31035 4705 31655 4725
rect 31035 4700 31040 4705
rect 31000 4695 31040 4700
rect 31650 4700 31655 4705
rect 31685 4725 31690 4730
rect 32260 4730 32300 4735
rect 32260 4725 32265 4730
rect 31685 4705 32265 4725
rect 31685 4700 31690 4705
rect 31650 4695 31690 4700
rect 32260 4700 32265 4705
rect 32295 4725 32300 4730
rect 32380 4730 32420 4735
rect 32380 4725 32385 4730
rect 32295 4705 32385 4725
rect 32295 4700 32300 4705
rect 32260 4695 32300 4700
rect 32380 4700 32385 4705
rect 32415 4725 32420 4730
rect 32500 4730 32540 4735
rect 32500 4725 32505 4730
rect 32415 4705 32505 4725
rect 32415 4700 32420 4705
rect 32380 4695 32420 4700
rect 32500 4700 32505 4705
rect 32535 4725 32540 4730
rect 32620 4730 32660 4735
rect 32620 4725 32625 4730
rect 32535 4705 32625 4725
rect 32535 4700 32540 4705
rect 32500 4695 32540 4700
rect 32620 4700 32625 4705
rect 32655 4700 32660 4730
rect 32620 4695 32660 4700
rect 31055 4545 31095 4550
rect 31055 4515 31060 4545
rect 31090 4540 31095 4545
rect 31310 4545 31350 4550
rect 31310 4540 31315 4545
rect 31090 4520 31315 4540
rect 31090 4515 31095 4520
rect 31055 4510 31095 4515
rect 31310 4515 31315 4520
rect 31345 4540 31350 4545
rect 32320 4545 32360 4550
rect 32320 4540 32325 4545
rect 31345 4520 32325 4540
rect 31345 4515 31350 4520
rect 31310 4510 31350 4515
rect 32320 4515 32325 4520
rect 32355 4515 32360 4545
rect 32320 4510 32360 4515
rect 30785 4440 30825 4445
rect 30785 4410 30790 4440
rect 30820 4435 30825 4440
rect 31250 4440 31290 4445
rect 31250 4435 31255 4440
rect 30820 4415 31255 4435
rect 30820 4410 30825 4415
rect 30785 4405 30825 4410
rect 31250 4410 31255 4415
rect 31285 4435 31290 4440
rect 31360 4440 31400 4445
rect 31360 4435 31365 4440
rect 31285 4415 31365 4435
rect 31285 4410 31290 4415
rect 31250 4405 31290 4410
rect 31360 4410 31365 4415
rect 31395 4435 31400 4440
rect 31470 4440 31510 4445
rect 31470 4435 31475 4440
rect 31395 4415 31475 4435
rect 31395 4410 31400 4415
rect 31360 4405 31400 4410
rect 31470 4410 31475 4415
rect 31505 4435 31510 4440
rect 31580 4440 31620 4445
rect 31580 4435 31585 4440
rect 31505 4415 31585 4435
rect 31505 4410 31510 4415
rect 31470 4405 31510 4410
rect 31580 4410 31585 4415
rect 31615 4435 31620 4440
rect 31690 4440 31730 4445
rect 31690 4435 31695 4440
rect 31615 4415 31695 4435
rect 31615 4410 31620 4415
rect 31580 4405 31620 4410
rect 31690 4410 31695 4415
rect 31725 4435 31730 4440
rect 31800 4440 31840 4445
rect 31800 4435 31805 4440
rect 31725 4415 31805 4435
rect 31725 4410 31730 4415
rect 31690 4405 31730 4410
rect 31800 4410 31805 4415
rect 31835 4435 31840 4440
rect 31910 4440 31950 4445
rect 31910 4435 31915 4440
rect 31835 4415 31915 4435
rect 31835 4410 31840 4415
rect 31800 4405 31840 4410
rect 31910 4410 31915 4415
rect 31945 4435 31950 4440
rect 32020 4440 32060 4445
rect 32020 4435 32025 4440
rect 31945 4415 32025 4435
rect 31945 4410 31950 4415
rect 31910 4405 31950 4410
rect 32020 4410 32025 4415
rect 32055 4435 32060 4440
rect 32130 4440 32170 4445
rect 32130 4435 32135 4440
rect 32055 4415 32135 4435
rect 32055 4410 32060 4415
rect 32020 4405 32060 4410
rect 32130 4410 32135 4415
rect 32165 4435 32170 4440
rect 32240 4440 32280 4445
rect 32240 4435 32245 4440
rect 32165 4415 32245 4435
rect 32165 4410 32170 4415
rect 32130 4405 32170 4410
rect 32240 4410 32245 4415
rect 32275 4435 32280 4440
rect 32350 4440 32390 4445
rect 32350 4435 32355 4440
rect 32275 4415 32355 4435
rect 32275 4410 32280 4415
rect 32240 4405 32280 4410
rect 32350 4410 32355 4415
rect 32385 4435 32390 4440
rect 32460 4440 32500 4445
rect 32460 4435 32465 4440
rect 32385 4415 32465 4435
rect 32385 4410 32390 4415
rect 32350 4405 32390 4410
rect 32460 4410 32465 4415
rect 32495 4410 32500 4440
rect 32460 4405 32500 4410
rect 31305 4320 31345 4325
rect 31305 4290 31310 4320
rect 31340 4315 31345 4320
rect 31525 4320 31565 4325
rect 31525 4315 31530 4320
rect 31340 4295 31530 4315
rect 31340 4290 31345 4295
rect 31305 4285 31345 4290
rect 31525 4290 31530 4295
rect 31560 4315 31565 4320
rect 31745 4320 31785 4325
rect 31745 4315 31750 4320
rect 31560 4295 31750 4315
rect 31560 4290 31565 4295
rect 31525 4285 31565 4290
rect 31745 4290 31750 4295
rect 31780 4315 31785 4320
rect 31965 4320 32005 4325
rect 31965 4315 31970 4320
rect 31780 4295 31970 4315
rect 31780 4290 31785 4295
rect 31745 4285 31785 4290
rect 31965 4290 31970 4295
rect 32000 4315 32005 4320
rect 32185 4320 32225 4325
rect 32185 4315 32190 4320
rect 32000 4295 32190 4315
rect 32000 4290 32005 4295
rect 31965 4285 32005 4290
rect 32185 4290 32190 4295
rect 32220 4315 32225 4320
rect 32405 4320 32445 4325
rect 32405 4315 32410 4320
rect 32220 4295 32410 4315
rect 32220 4290 32225 4295
rect 32185 4285 32225 4290
rect 32405 4290 32410 4295
rect 32440 4290 32445 4320
rect 32405 4285 32445 4290
rect 31420 4205 31460 4210
rect 31420 4175 31425 4205
rect 31455 4200 31460 4205
rect 31635 4205 31675 4210
rect 31635 4200 31640 4205
rect 31455 4180 31640 4200
rect 31455 4175 31460 4180
rect 31420 4170 31460 4175
rect 31635 4175 31640 4180
rect 31670 4200 31675 4205
rect 31855 4205 31895 4210
rect 31855 4200 31860 4205
rect 31670 4180 31860 4200
rect 31670 4175 31675 4180
rect 31635 4170 31675 4175
rect 31855 4175 31860 4180
rect 31890 4200 31895 4205
rect 32075 4205 32115 4210
rect 32075 4200 32080 4205
rect 31890 4180 32080 4200
rect 31890 4175 31895 4180
rect 31855 4170 31895 4175
rect 32075 4175 32080 4180
rect 32110 4200 32115 4205
rect 32295 4205 32335 4210
rect 32295 4200 32300 4205
rect 32110 4180 32300 4200
rect 32110 4175 32115 4180
rect 32075 4170 32115 4175
rect 32295 4175 32300 4180
rect 32330 4175 32335 4205
rect 32295 4170 32335 4175
rect 31320 4090 31360 4095
rect 31320 4060 31325 4090
rect 31355 4085 31360 4090
rect 31420 4090 31460 4095
rect 31420 4085 31425 4090
rect 31355 4065 31425 4085
rect 31355 4060 31360 4065
rect 31320 4055 31360 4060
rect 31420 4060 31425 4065
rect 31455 4085 31460 4090
rect 31530 4090 31570 4095
rect 31530 4085 31535 4090
rect 31455 4065 31535 4085
rect 31455 4060 31460 4065
rect 31420 4055 31460 4060
rect 31530 4060 31535 4065
rect 31565 4085 31570 4090
rect 31640 4090 31680 4095
rect 31640 4085 31645 4090
rect 31565 4065 31645 4085
rect 31565 4060 31570 4065
rect 31530 4055 31570 4060
rect 31640 4060 31645 4065
rect 31675 4085 31680 4090
rect 31750 4090 31790 4095
rect 31750 4085 31755 4090
rect 31675 4065 31755 4085
rect 31675 4060 31680 4065
rect 31640 4055 31680 4060
rect 31750 4060 31755 4065
rect 31785 4060 31790 4090
rect 31750 4055 31790 4060
rect 32050 4090 32090 4095
rect 32050 4060 32055 4090
rect 32085 4085 32090 4090
rect 32150 4090 32190 4095
rect 32150 4085 32155 4090
rect 32085 4065 32155 4085
rect 32085 4060 32090 4065
rect 32050 4055 32090 4060
rect 32150 4060 32155 4065
rect 32185 4085 32190 4090
rect 32260 4090 32300 4095
rect 32260 4085 32265 4090
rect 32185 4065 32265 4085
rect 32185 4060 32190 4065
rect 32150 4055 32190 4060
rect 32260 4060 32265 4065
rect 32295 4085 32300 4090
rect 32370 4090 32410 4095
rect 32370 4085 32375 4090
rect 32295 4065 32375 4085
rect 32295 4060 32300 4065
rect 32260 4055 32300 4060
rect 32370 4060 32375 4065
rect 32405 4085 32410 4090
rect 32480 4090 32520 4095
rect 32480 4085 32485 4090
rect 32405 4065 32485 4085
rect 32405 4060 32410 4065
rect 32370 4055 32410 4060
rect 32480 4060 32485 4065
rect 32515 4060 32520 4090
rect 32480 4055 32520 4060
rect 31280 4029 31310 4035
rect 31280 4001 31282 4029
rect 31308 4025 31310 4029
rect 31480 4029 31510 4035
rect 31480 4025 31482 4029
rect 31308 4005 31482 4025
rect 31308 4001 31310 4005
rect 31280 3995 31310 4001
rect 31480 4001 31482 4005
rect 31508 4025 31510 4029
rect 31695 4030 31735 4035
rect 31695 4025 31700 4030
rect 31508 4005 31700 4025
rect 31508 4001 31510 4005
rect 31480 3995 31510 4001
rect 31695 4000 31700 4005
rect 31730 4025 31735 4030
rect 32008 4029 32038 4035
rect 32008 4025 32010 4029
rect 31730 4005 32010 4025
rect 31730 4000 31735 4005
rect 31695 3995 31735 4000
rect 32008 4001 32010 4005
rect 32036 4025 32038 4029
rect 32205 4030 32245 4035
rect 32205 4025 32210 4030
rect 32036 4005 32210 4025
rect 32036 4001 32038 4005
rect 32008 3995 32038 4001
rect 32205 4000 32210 4005
rect 32240 4025 32245 4030
rect 32425 4030 32465 4035
rect 32425 4025 32430 4030
rect 32240 4005 32430 4025
rect 32240 4000 32245 4005
rect 32205 3995 32245 4000
rect 32425 4000 32430 4005
rect 32460 4025 32465 4030
rect 32870 4030 32910 4035
rect 32870 4025 32875 4030
rect 32460 4005 32875 4025
rect 32460 4000 32465 4005
rect 32425 3995 32465 4000
rect 32870 4000 32875 4005
rect 32905 4000 32910 4030
rect 32870 3995 32910 4000
rect 30785 3970 30825 3975
rect 30785 3940 30790 3970
rect 30820 3965 30825 3970
rect 31140 3970 31180 3975
rect 31140 3965 31145 3970
rect 30820 3945 31145 3965
rect 30820 3940 30825 3945
rect 30785 3935 30825 3940
rect 31140 3940 31145 3945
rect 31175 3940 31180 3970
rect 31140 3935 31180 3940
rect 31407 3910 31439 3915
rect 31407 3905 31410 3910
rect 30950 3885 31410 3905
rect 31407 3880 31410 3885
rect 31436 3905 31439 3910
rect 31627 3910 31659 3915
rect 31627 3905 31630 3910
rect 31436 3885 31630 3905
rect 31436 3880 31439 3885
rect 31407 3875 31439 3880
rect 31627 3880 31630 3885
rect 31656 3905 31659 3910
rect 31771 3910 31803 3915
rect 31771 3905 31774 3910
rect 31656 3885 31774 3905
rect 31656 3880 31659 3885
rect 31627 3875 31659 3880
rect 31771 3880 31774 3885
rect 31800 3905 31803 3910
rect 32137 3910 32169 3915
rect 32137 3905 32140 3910
rect 31800 3885 32140 3905
rect 31800 3880 31803 3885
rect 31771 3875 31803 3880
rect 32137 3880 32140 3885
rect 32166 3905 32169 3910
rect 32357 3910 32389 3915
rect 32357 3905 32360 3910
rect 32166 3885 32360 3905
rect 32166 3880 32169 3885
rect 32137 3875 32169 3880
rect 32357 3880 32360 3885
rect 32386 3905 32389 3910
rect 32501 3910 32533 3915
rect 32501 3905 32504 3910
rect 32386 3885 32504 3905
rect 32386 3880 32389 3885
rect 32357 3875 32389 3880
rect 32501 3880 32504 3885
rect 32530 3905 32533 3910
rect 32530 3885 32535 3905
rect 32530 3880 32533 3885
rect 32501 3875 32533 3880
rect 31255 3850 31295 3855
rect 31255 3820 31260 3850
rect 31290 3845 31295 3850
rect 31360 3850 31400 3855
rect 31360 3845 31365 3850
rect 31290 3825 31365 3845
rect 31290 3820 31295 3825
rect 31255 3815 31295 3820
rect 31360 3820 31365 3825
rect 31395 3845 31400 3850
rect 31475 3850 31515 3855
rect 31475 3845 31480 3850
rect 31395 3825 31480 3845
rect 31395 3820 31400 3825
rect 31360 3815 31400 3820
rect 31475 3820 31480 3825
rect 31510 3845 31515 3850
rect 31580 3850 31620 3855
rect 31580 3845 31585 3850
rect 31510 3825 31585 3845
rect 31510 3820 31515 3825
rect 31475 3815 31515 3820
rect 31580 3820 31585 3825
rect 31615 3845 31620 3850
rect 31695 3850 31735 3855
rect 31695 3845 31700 3850
rect 31615 3825 31700 3845
rect 31615 3820 31620 3825
rect 31580 3815 31620 3820
rect 31695 3820 31700 3825
rect 31730 3845 31735 3850
rect 31810 3850 31850 3855
rect 31810 3845 31815 3850
rect 31730 3825 31815 3845
rect 31730 3820 31735 3825
rect 31695 3815 31735 3820
rect 31810 3820 31815 3825
rect 31845 3820 31850 3850
rect 31810 3815 31850 3820
rect 31985 3850 32025 3855
rect 31985 3820 31990 3850
rect 32020 3845 32025 3850
rect 32205 3850 32245 3855
rect 32205 3845 32210 3850
rect 32020 3825 32210 3845
rect 32020 3820 32025 3825
rect 31985 3815 32025 3820
rect 32205 3820 32210 3825
rect 32240 3845 32245 3850
rect 32425 3850 32465 3855
rect 32425 3845 32430 3850
rect 32240 3825 32430 3845
rect 32240 3820 32245 3825
rect 32205 3815 32245 3820
rect 32425 3820 32430 3825
rect 32460 3845 32465 3850
rect 32960 3850 33000 3855
rect 32960 3845 32965 3850
rect 32460 3825 32965 3845
rect 32460 3820 32465 3825
rect 32425 3815 32465 3820
rect 32960 3820 32965 3825
rect 32995 3820 33000 3850
rect 32960 3815 33000 3820
rect 32080 3760 32120 3765
rect 29605 3735 29645 3740
rect 29605 3705 29610 3735
rect 29640 3705 29645 3735
rect 32080 3730 32085 3760
rect 32115 3755 32120 3760
rect 32300 3760 32340 3765
rect 32300 3755 32305 3760
rect 32115 3735 32305 3755
rect 32115 3730 32120 3735
rect 31880 3725 31920 3730
rect 32080 3725 32120 3730
rect 32300 3730 32305 3735
rect 32335 3755 32340 3760
rect 32540 3760 32580 3765
rect 32540 3755 32545 3760
rect 32335 3735 32545 3755
rect 32335 3730 32340 3735
rect 32300 3725 32340 3730
rect 32540 3730 32545 3735
rect 32575 3755 32580 3760
rect 32915 3760 32955 3765
rect 32915 3755 32920 3760
rect 32575 3735 32920 3755
rect 32575 3730 32580 3735
rect 32540 3725 32580 3730
rect 32915 3730 32920 3735
rect 32950 3730 32955 3760
rect 32915 3725 32955 3730
rect 34155 3735 34195 3740
rect 29605 3700 29645 3705
rect 29955 3715 29995 3720
rect 29955 3685 29960 3715
rect 29990 3710 29995 3715
rect 30065 3715 30105 3720
rect 30065 3710 30070 3715
rect 29990 3690 30070 3710
rect 29990 3685 29995 3690
rect 29955 3680 29995 3685
rect 30065 3685 30070 3690
rect 30100 3710 30105 3715
rect 30175 3715 30215 3720
rect 30175 3710 30180 3715
rect 30100 3690 30180 3710
rect 30100 3685 30105 3690
rect 30065 3680 30105 3685
rect 30175 3685 30180 3690
rect 30210 3710 30215 3715
rect 30285 3715 30325 3720
rect 30285 3710 30290 3715
rect 30210 3690 30290 3710
rect 30210 3685 30215 3690
rect 30175 3680 30215 3685
rect 30285 3685 30290 3690
rect 30320 3710 30325 3715
rect 30395 3715 30435 3720
rect 30395 3710 30400 3715
rect 30320 3690 30400 3710
rect 30320 3685 30325 3690
rect 30285 3680 30325 3685
rect 30395 3685 30400 3690
rect 30430 3710 30435 3715
rect 30505 3715 30545 3720
rect 30505 3710 30510 3715
rect 30430 3690 30510 3710
rect 30430 3685 30435 3690
rect 30395 3680 30435 3685
rect 30505 3685 30510 3690
rect 30540 3710 30545 3715
rect 30615 3715 30655 3720
rect 30615 3710 30620 3715
rect 30540 3690 30620 3710
rect 30540 3685 30545 3690
rect 30505 3680 30545 3685
rect 30615 3685 30620 3690
rect 30650 3710 30655 3715
rect 30785 3715 30825 3720
rect 30785 3710 30790 3715
rect 30650 3690 30790 3710
rect 30650 3685 30655 3690
rect 30615 3680 30655 3685
rect 30785 3685 30790 3690
rect 30820 3710 30825 3715
rect 31880 3710 31885 3725
rect 30820 3695 31885 3710
rect 31915 3710 31920 3725
rect 33005 3715 33045 3720
rect 33005 3710 33010 3715
rect 31915 3695 33010 3710
rect 30820 3690 33010 3695
rect 30820 3685 30825 3690
rect 30785 3680 30825 3685
rect 33005 3685 33010 3690
rect 33040 3710 33045 3715
rect 33145 3715 33185 3720
rect 33145 3710 33150 3715
rect 33040 3690 33150 3710
rect 33040 3685 33045 3690
rect 33005 3680 33045 3685
rect 33145 3685 33150 3690
rect 33180 3710 33185 3715
rect 33255 3715 33295 3720
rect 33255 3710 33260 3715
rect 33180 3690 33260 3710
rect 33180 3685 33185 3690
rect 33145 3680 33185 3685
rect 33255 3685 33260 3690
rect 33290 3710 33295 3715
rect 33365 3715 33405 3720
rect 33365 3710 33370 3715
rect 33290 3690 33370 3710
rect 33290 3685 33295 3690
rect 33255 3680 33295 3685
rect 33365 3685 33370 3690
rect 33400 3710 33405 3715
rect 33475 3715 33515 3720
rect 33475 3710 33480 3715
rect 33400 3690 33480 3710
rect 33400 3685 33405 3690
rect 33365 3680 33405 3685
rect 33475 3685 33480 3690
rect 33510 3710 33515 3715
rect 33585 3715 33625 3720
rect 33585 3710 33590 3715
rect 33510 3690 33590 3710
rect 33510 3685 33515 3690
rect 33475 3680 33515 3685
rect 33585 3685 33590 3690
rect 33620 3710 33625 3715
rect 33695 3715 33735 3720
rect 33695 3710 33700 3715
rect 33620 3690 33700 3710
rect 33620 3685 33625 3690
rect 33585 3680 33625 3685
rect 33695 3685 33700 3690
rect 33730 3710 33735 3715
rect 33805 3715 33845 3720
rect 33805 3710 33810 3715
rect 33730 3690 33810 3710
rect 33730 3685 33735 3690
rect 33695 3680 33735 3685
rect 33805 3685 33810 3690
rect 33840 3685 33845 3715
rect 34155 3705 34160 3735
rect 34190 3705 34195 3735
rect 34155 3700 34195 3705
rect 33805 3680 33845 3685
rect 31880 3665 31920 3670
rect 29554 3655 29695 3660
rect 29554 3625 29560 3655
rect 29590 3625 29610 3655
rect 29640 3625 29659 3655
rect 29689 3625 29695 3655
rect 31880 3635 31885 3665
rect 31915 3635 31920 3665
rect 31880 3630 31920 3635
rect 34105 3655 34246 3660
rect 29554 3620 29695 3625
rect 34105 3625 34111 3655
rect 34141 3625 34160 3655
rect 34190 3625 34210 3655
rect 34240 3625 34246 3655
rect 34105 3620 34246 3625
rect 31340 3605 31380 3610
rect 31340 3575 31345 3605
rect 31375 3600 31380 3605
rect 31460 3605 31500 3610
rect 31460 3600 31465 3605
rect 31375 3580 31465 3600
rect 31375 3575 31380 3580
rect 31340 3570 31380 3575
rect 31460 3575 31465 3580
rect 31495 3600 31500 3605
rect 31580 3605 31620 3610
rect 31580 3600 31585 3605
rect 31495 3580 31585 3600
rect 31495 3575 31500 3580
rect 31460 3570 31500 3575
rect 31580 3575 31585 3580
rect 31615 3600 31620 3605
rect 31700 3605 31740 3610
rect 31700 3600 31705 3605
rect 31615 3580 31705 3600
rect 31615 3575 31620 3580
rect 31580 3570 31620 3575
rect 31700 3575 31705 3580
rect 31735 3600 31740 3605
rect 31820 3605 31860 3610
rect 31820 3600 31825 3605
rect 31735 3580 31825 3600
rect 31735 3575 31740 3580
rect 31700 3570 31740 3575
rect 31820 3575 31825 3580
rect 31855 3600 31860 3605
rect 31880 3605 31920 3610
rect 31880 3600 31885 3605
rect 31855 3580 31885 3600
rect 31855 3575 31860 3580
rect 31820 3570 31860 3575
rect 31880 3575 31885 3580
rect 31915 3600 31920 3605
rect 31940 3605 31980 3610
rect 31940 3600 31945 3605
rect 31915 3580 31945 3600
rect 31915 3575 31920 3580
rect 31880 3570 31920 3575
rect 31940 3575 31945 3580
rect 31975 3600 31980 3605
rect 32060 3605 32100 3610
rect 32060 3600 32065 3605
rect 31975 3580 32065 3600
rect 31975 3575 31980 3580
rect 31940 3570 31980 3575
rect 32060 3575 32065 3580
rect 32095 3600 32100 3605
rect 32180 3605 32220 3610
rect 32180 3600 32185 3605
rect 32095 3580 32185 3600
rect 32095 3575 32100 3580
rect 32060 3570 32100 3575
rect 32180 3575 32185 3580
rect 32215 3600 32220 3605
rect 32300 3605 32340 3610
rect 32300 3600 32305 3605
rect 32215 3580 32305 3600
rect 32215 3575 32220 3580
rect 32180 3570 32220 3575
rect 32300 3575 32305 3580
rect 32335 3600 32340 3605
rect 32420 3605 32460 3610
rect 32420 3600 32425 3605
rect 32335 3580 32425 3600
rect 32335 3575 32340 3580
rect 32300 3570 32340 3575
rect 32420 3575 32425 3580
rect 32455 3575 32460 3605
rect 32420 3570 32460 3575
rect 31000 3185 31040 3190
rect 31000 3155 31005 3185
rect 31035 3180 31040 3185
rect 31823 3185 31857 3190
rect 31823 3180 31826 3185
rect 31035 3160 31826 3180
rect 31035 3155 31040 3160
rect 31000 3150 31040 3155
rect 31823 3155 31826 3160
rect 31854 3155 31857 3185
rect 31823 3150 31857 3155
rect 31280 3130 31320 3135
rect 31280 3100 31285 3130
rect 31315 3125 31320 3130
rect 31520 3130 31560 3135
rect 31520 3125 31525 3130
rect 31315 3105 31525 3125
rect 31315 3100 31320 3105
rect 31280 3095 31320 3100
rect 31520 3100 31525 3105
rect 31555 3125 31560 3130
rect 31760 3130 31800 3135
rect 31760 3125 31765 3130
rect 31555 3105 31765 3125
rect 31555 3100 31560 3105
rect 31520 3095 31560 3100
rect 31760 3100 31765 3105
rect 31795 3125 31800 3130
rect 32000 3130 32040 3135
rect 32000 3125 32005 3130
rect 31795 3105 32005 3125
rect 31795 3100 31800 3105
rect 31760 3095 31800 3100
rect 32000 3100 32005 3105
rect 32035 3125 32040 3130
rect 32240 3130 32280 3135
rect 32240 3125 32245 3130
rect 32035 3105 32245 3125
rect 32035 3100 32040 3105
rect 32000 3095 32040 3100
rect 32240 3100 32245 3105
rect 32275 3125 32280 3130
rect 32480 3130 32520 3135
rect 32480 3125 32485 3130
rect 32275 3105 32485 3125
rect 32275 3100 32280 3105
rect 32240 3095 32280 3100
rect 32480 3100 32485 3105
rect 32515 3100 32520 3130
rect 32480 3095 32520 3100
rect 29554 3050 29695 3055
rect 34105 3050 34246 3055
rect 29554 3020 29560 3050
rect 29590 3020 29610 3050
rect 29640 3020 29659 3050
rect 29689 3020 29695 3050
rect 29554 3015 29695 3020
rect 30010 3045 30050 3050
rect 30010 3015 30015 3045
rect 30045 3040 30050 3045
rect 30120 3045 30160 3050
rect 30120 3040 30125 3045
rect 30045 3020 30125 3040
rect 30045 3015 30050 3020
rect 30010 3010 30050 3015
rect 30120 3015 30125 3020
rect 30155 3040 30160 3045
rect 30230 3045 30270 3050
rect 30230 3040 30235 3045
rect 30155 3020 30235 3040
rect 30155 3015 30160 3020
rect 30120 3010 30160 3015
rect 30230 3015 30235 3020
rect 30265 3040 30270 3045
rect 30340 3045 30380 3050
rect 30340 3040 30345 3045
rect 30265 3020 30345 3040
rect 30265 3015 30270 3020
rect 30230 3010 30270 3015
rect 30340 3015 30345 3020
rect 30375 3040 30380 3045
rect 30450 3045 30490 3050
rect 30450 3040 30455 3045
rect 30375 3020 30455 3040
rect 30375 3015 30380 3020
rect 30340 3010 30380 3015
rect 30450 3015 30455 3020
rect 30485 3040 30490 3045
rect 30560 3045 30600 3050
rect 30560 3040 30565 3045
rect 30485 3020 30565 3040
rect 30485 3015 30490 3020
rect 30450 3010 30490 3015
rect 30560 3015 30565 3020
rect 30595 3015 30600 3045
rect 30560 3010 30600 3015
rect 31400 3045 31440 3050
rect 31400 3015 31405 3045
rect 31435 3040 31440 3045
rect 31640 3045 31680 3050
rect 31640 3040 31645 3045
rect 31435 3020 31645 3040
rect 31435 3015 31440 3020
rect 31400 3010 31440 3015
rect 31640 3015 31645 3020
rect 31675 3040 31680 3045
rect 31880 3045 31920 3050
rect 31880 3040 31885 3045
rect 31675 3020 31885 3040
rect 31675 3015 31680 3020
rect 31640 3010 31680 3015
rect 31880 3015 31885 3020
rect 31915 3040 31920 3045
rect 32120 3045 32160 3050
rect 32120 3040 32125 3045
rect 31915 3020 32125 3040
rect 31915 3015 31920 3020
rect 31880 3010 31920 3015
rect 32120 3015 32125 3020
rect 32155 3040 32160 3045
rect 32360 3045 32400 3050
rect 32360 3040 32365 3045
rect 32155 3020 32365 3040
rect 32155 3015 32160 3020
rect 32120 3010 32160 3015
rect 32360 3015 32365 3020
rect 32395 3015 32400 3045
rect 32360 3010 32400 3015
rect 33200 3045 33240 3050
rect 33200 3015 33205 3045
rect 33235 3040 33240 3045
rect 33310 3045 33350 3050
rect 33310 3040 33315 3045
rect 33235 3020 33315 3040
rect 33235 3015 33240 3020
rect 33200 3010 33240 3015
rect 33310 3015 33315 3020
rect 33345 3040 33350 3045
rect 33420 3045 33460 3050
rect 33420 3040 33425 3045
rect 33345 3020 33425 3040
rect 33345 3015 33350 3020
rect 33310 3010 33350 3015
rect 33420 3015 33425 3020
rect 33455 3040 33460 3045
rect 33530 3045 33570 3050
rect 33530 3040 33535 3045
rect 33455 3020 33535 3040
rect 33455 3015 33460 3020
rect 33420 3010 33460 3015
rect 33530 3015 33535 3020
rect 33565 3040 33570 3045
rect 33640 3045 33680 3050
rect 33640 3040 33645 3045
rect 33565 3020 33645 3040
rect 33565 3015 33570 3020
rect 33530 3010 33570 3015
rect 33640 3015 33645 3020
rect 33675 3040 33680 3045
rect 33750 3045 33790 3050
rect 33750 3040 33755 3045
rect 33675 3020 33755 3040
rect 33675 3015 33680 3020
rect 33640 3010 33680 3015
rect 33750 3015 33755 3020
rect 33785 3015 33790 3045
rect 34105 3020 34111 3050
rect 34141 3020 34160 3050
rect 34190 3020 34210 3050
rect 34240 3020 34246 3050
rect 34105 3015 34246 3020
rect 33750 3010 33790 3015
rect 31055 2990 31095 2995
rect 31055 2960 31060 2990
rect 31090 2985 31095 2990
rect 31880 2990 31920 2995
rect 31880 2985 31885 2990
rect 31090 2965 31885 2985
rect 31090 2960 31095 2965
rect 31055 2955 31095 2960
rect 31880 2960 31885 2965
rect 31915 2960 31920 2990
rect 31880 2955 31920 2960
rect 33040 2935 33080 2940
rect 29605 2925 29645 2930
rect 29605 2895 29610 2925
rect 29640 2920 29645 2925
rect 30175 2925 30215 2930
rect 30175 2920 30180 2925
rect 29640 2900 30180 2920
rect 29640 2895 29645 2900
rect 29605 2890 29645 2895
rect 30175 2895 30180 2900
rect 30210 2920 30215 2925
rect 30740 2925 30780 2930
rect 30740 2920 30745 2925
rect 30210 2900 30745 2920
rect 30210 2895 30215 2900
rect 30175 2890 30215 2895
rect 30740 2895 30745 2900
rect 30775 2895 30780 2925
rect 33040 2905 33045 2935
rect 33075 2930 33080 2935
rect 33585 2935 33625 2940
rect 33585 2930 33590 2935
rect 33075 2910 33590 2930
rect 33075 2905 33080 2910
rect 33040 2900 33080 2905
rect 33585 2905 33590 2910
rect 33620 2930 33625 2935
rect 34155 2935 34195 2940
rect 34155 2930 34160 2935
rect 33620 2910 34160 2930
rect 33620 2905 33625 2910
rect 33585 2900 33625 2905
rect 34155 2905 34160 2910
rect 34190 2905 34195 2935
rect 34155 2900 34195 2905
rect 30740 2890 30780 2895
rect 31125 2895 31165 2900
rect 29315 2870 29355 2875
rect 29315 2840 29320 2870
rect 29350 2865 29355 2870
rect 30450 2870 30490 2875
rect 30450 2865 30455 2870
rect 29350 2845 30455 2865
rect 29350 2840 29355 2845
rect 29315 2835 29355 2840
rect 30450 2840 30455 2845
rect 30485 2840 30490 2870
rect 31125 2865 31130 2895
rect 31160 2890 31165 2895
rect 31245 2895 31285 2900
rect 31245 2890 31250 2895
rect 31160 2870 31250 2890
rect 31160 2865 31165 2870
rect 31125 2860 31165 2865
rect 31245 2865 31250 2870
rect 31280 2890 31285 2895
rect 31365 2895 31405 2900
rect 31365 2890 31370 2895
rect 31280 2870 31370 2890
rect 31280 2865 31285 2870
rect 31245 2860 31285 2865
rect 31365 2865 31370 2870
rect 31400 2890 31405 2895
rect 31485 2895 31525 2900
rect 31485 2890 31490 2895
rect 31400 2870 31490 2890
rect 31400 2865 31405 2870
rect 31365 2860 31405 2865
rect 31485 2865 31490 2870
rect 31520 2890 31525 2895
rect 31605 2895 31645 2900
rect 31605 2890 31610 2895
rect 31520 2870 31610 2890
rect 31520 2865 31525 2870
rect 31485 2860 31525 2865
rect 31605 2865 31610 2870
rect 31640 2865 31645 2895
rect 31605 2860 31645 2865
rect 32155 2895 32195 2900
rect 32155 2865 32160 2895
rect 32190 2890 32195 2895
rect 32275 2895 32315 2900
rect 32275 2890 32280 2895
rect 32190 2870 32280 2890
rect 32190 2865 32195 2870
rect 32155 2860 32195 2865
rect 32275 2865 32280 2870
rect 32310 2890 32315 2895
rect 32395 2895 32435 2900
rect 32395 2890 32400 2895
rect 32310 2870 32400 2890
rect 32310 2865 32315 2870
rect 32275 2860 32315 2865
rect 32395 2865 32400 2870
rect 32430 2890 32435 2895
rect 32515 2895 32555 2900
rect 32515 2890 32520 2895
rect 32430 2870 32520 2890
rect 32430 2865 32435 2870
rect 32395 2860 32435 2865
rect 32515 2865 32520 2870
rect 32550 2890 32555 2895
rect 32635 2895 32675 2900
rect 32635 2890 32640 2895
rect 32550 2870 32640 2890
rect 32550 2865 32555 2870
rect 32515 2860 32555 2865
rect 32635 2865 32640 2870
rect 32670 2865 32675 2895
rect 32635 2860 32675 2865
rect 33310 2890 33350 2895
rect 33310 2860 33315 2890
rect 33345 2885 33350 2890
rect 34445 2890 34485 2895
rect 34445 2885 34450 2890
rect 33345 2865 34450 2885
rect 33345 2860 33350 2865
rect 33310 2855 33350 2860
rect 34445 2860 34450 2865
rect 34480 2860 34485 2890
rect 34445 2855 34485 2860
rect 30450 2835 30490 2840
rect 29265 2755 29305 2760
rect 29265 2725 29270 2755
rect 29300 2750 29305 2755
rect 30010 2755 30050 2760
rect 30010 2750 30015 2755
rect 29300 2730 30015 2750
rect 29300 2725 29305 2730
rect 29265 2720 29305 2725
rect 30010 2725 30015 2730
rect 30045 2750 30050 2755
rect 30120 2755 30160 2760
rect 30120 2750 30125 2755
rect 30045 2730 30125 2750
rect 30045 2725 30050 2730
rect 30010 2720 30050 2725
rect 30120 2725 30125 2730
rect 30155 2750 30160 2755
rect 30230 2755 30270 2760
rect 30230 2750 30235 2755
rect 30155 2730 30235 2750
rect 30155 2725 30160 2730
rect 30120 2720 30160 2725
rect 30230 2725 30235 2730
rect 30265 2750 30270 2755
rect 30340 2755 30380 2760
rect 30340 2750 30345 2755
rect 30265 2730 30345 2750
rect 30265 2725 30270 2730
rect 30230 2720 30270 2725
rect 30340 2725 30345 2730
rect 30375 2750 30380 2755
rect 30450 2755 30490 2760
rect 30450 2750 30455 2755
rect 30375 2730 30455 2750
rect 30375 2725 30380 2730
rect 30340 2720 30380 2725
rect 30450 2725 30455 2730
rect 30485 2750 30490 2755
rect 30560 2755 30600 2760
rect 30560 2750 30565 2755
rect 30485 2730 30565 2750
rect 30485 2725 30490 2730
rect 30450 2720 30490 2725
rect 30560 2725 30565 2730
rect 30595 2725 30600 2755
rect 30560 2720 30600 2725
rect 33200 2755 33240 2760
rect 33200 2725 33205 2755
rect 33235 2750 33240 2755
rect 33310 2755 33350 2760
rect 33310 2750 33315 2755
rect 33235 2730 33315 2750
rect 33235 2725 33240 2730
rect 33200 2720 33240 2725
rect 33310 2725 33315 2730
rect 33345 2750 33350 2755
rect 33420 2755 33460 2760
rect 33420 2750 33425 2755
rect 33345 2730 33425 2750
rect 33345 2725 33350 2730
rect 33310 2720 33350 2725
rect 33420 2725 33425 2730
rect 33455 2750 33460 2755
rect 33530 2755 33570 2760
rect 33530 2750 33535 2755
rect 33455 2730 33535 2750
rect 33455 2725 33460 2730
rect 33420 2720 33460 2725
rect 33530 2725 33535 2730
rect 33565 2750 33570 2755
rect 33640 2755 33680 2760
rect 33640 2750 33645 2755
rect 33565 2730 33645 2750
rect 33565 2725 33570 2730
rect 33530 2720 33570 2725
rect 33640 2725 33645 2730
rect 33675 2750 33680 2755
rect 33750 2755 33790 2760
rect 33750 2750 33755 2755
rect 33675 2730 33755 2750
rect 33675 2725 33680 2730
rect 33640 2720 33680 2725
rect 33750 2725 33755 2730
rect 33785 2750 33790 2755
rect 34495 2755 34535 2760
rect 34495 2750 34500 2755
rect 33785 2730 34500 2750
rect 33785 2725 33790 2730
rect 33750 2720 33790 2725
rect 34495 2725 34500 2730
rect 34530 2725 34535 2755
rect 34495 2720 34535 2725
rect 29790 2485 29830 2490
rect 29790 2455 29795 2485
rect 29825 2480 29830 2485
rect 30065 2485 30105 2490
rect 30065 2480 30070 2485
rect 29825 2460 30070 2480
rect 29825 2455 29830 2460
rect 29790 2450 29830 2455
rect 30065 2455 30070 2460
rect 30100 2480 30105 2485
rect 30175 2485 30215 2490
rect 30175 2480 30180 2485
rect 30100 2460 30180 2480
rect 30100 2455 30105 2460
rect 30065 2450 30105 2455
rect 30175 2455 30180 2460
rect 30210 2480 30215 2485
rect 30285 2485 30325 2490
rect 30285 2480 30290 2485
rect 30210 2460 30290 2480
rect 30210 2455 30215 2460
rect 30175 2450 30215 2455
rect 30285 2455 30290 2460
rect 30320 2480 30325 2485
rect 30395 2485 30435 2490
rect 30395 2480 30400 2485
rect 30320 2460 30400 2480
rect 30320 2455 30325 2460
rect 30285 2450 30325 2455
rect 30395 2455 30400 2460
rect 30430 2480 30435 2485
rect 30505 2485 30545 2490
rect 30505 2480 30510 2485
rect 30430 2460 30510 2480
rect 30430 2455 30435 2460
rect 30395 2450 30435 2455
rect 30505 2455 30510 2460
rect 30540 2455 30545 2485
rect 33255 2485 33295 2490
rect 30505 2450 30545 2455
rect 31065 2475 31105 2480
rect 31065 2445 31070 2475
rect 31100 2470 31105 2475
rect 31185 2475 31225 2480
rect 31185 2470 31190 2475
rect 31100 2450 31190 2470
rect 31100 2445 31105 2450
rect 31065 2440 31105 2445
rect 31185 2445 31190 2450
rect 31220 2470 31225 2475
rect 31305 2475 31345 2480
rect 31305 2470 31310 2475
rect 31220 2450 31310 2470
rect 31220 2445 31225 2450
rect 31185 2440 31225 2445
rect 31305 2445 31310 2450
rect 31340 2470 31345 2475
rect 31425 2475 31465 2480
rect 31425 2470 31430 2475
rect 31340 2450 31430 2470
rect 31340 2445 31345 2450
rect 31305 2440 31345 2445
rect 31425 2445 31430 2450
rect 31460 2470 31465 2475
rect 31545 2475 31585 2480
rect 31545 2470 31550 2475
rect 31460 2450 31550 2470
rect 31460 2445 31465 2450
rect 31425 2440 31465 2445
rect 31545 2445 31550 2450
rect 31580 2470 31585 2475
rect 31665 2475 31705 2480
rect 31665 2470 31670 2475
rect 31580 2450 31670 2470
rect 31580 2445 31585 2450
rect 31545 2440 31585 2445
rect 31665 2445 31670 2450
rect 31700 2445 31705 2475
rect 31665 2440 31705 2445
rect 32095 2475 32135 2480
rect 32095 2445 32100 2475
rect 32130 2470 32135 2475
rect 32215 2475 32255 2480
rect 32215 2470 32220 2475
rect 32130 2450 32220 2470
rect 32130 2445 32135 2450
rect 32095 2440 32135 2445
rect 32215 2445 32220 2450
rect 32250 2470 32255 2475
rect 32335 2475 32375 2480
rect 32335 2470 32340 2475
rect 32250 2450 32340 2470
rect 32250 2445 32255 2450
rect 32215 2440 32255 2445
rect 32335 2445 32340 2450
rect 32370 2470 32375 2475
rect 32455 2475 32495 2480
rect 32455 2470 32460 2475
rect 32370 2450 32460 2470
rect 32370 2445 32375 2450
rect 32335 2440 32375 2445
rect 32455 2445 32460 2450
rect 32490 2470 32495 2475
rect 32575 2475 32615 2480
rect 32575 2470 32580 2475
rect 32490 2450 32580 2470
rect 32490 2445 32495 2450
rect 32455 2440 32495 2445
rect 32575 2445 32580 2450
rect 32610 2470 32615 2475
rect 32695 2475 32735 2480
rect 32695 2470 32700 2475
rect 32610 2450 32700 2470
rect 32610 2445 32615 2450
rect 32575 2440 32615 2445
rect 32695 2445 32700 2450
rect 32730 2445 32735 2475
rect 33255 2455 33260 2485
rect 33290 2480 33295 2485
rect 33365 2485 33405 2490
rect 33365 2480 33370 2485
rect 33290 2460 33370 2480
rect 33290 2455 33295 2460
rect 33255 2450 33295 2455
rect 33365 2455 33370 2460
rect 33400 2480 33405 2485
rect 33475 2485 33515 2490
rect 33475 2480 33480 2485
rect 33400 2460 33480 2480
rect 33400 2455 33405 2460
rect 33365 2450 33405 2455
rect 33475 2455 33480 2460
rect 33510 2480 33515 2485
rect 33585 2485 33625 2490
rect 33585 2480 33590 2485
rect 33510 2460 33590 2480
rect 33510 2455 33515 2460
rect 33475 2450 33515 2455
rect 33585 2455 33590 2460
rect 33620 2480 33625 2485
rect 33695 2485 33735 2490
rect 33695 2480 33700 2485
rect 33620 2460 33700 2480
rect 33620 2455 33625 2460
rect 33585 2450 33625 2455
rect 33695 2455 33700 2460
rect 33730 2480 33735 2485
rect 33975 2485 34015 2490
rect 33975 2480 33980 2485
rect 33730 2460 33980 2480
rect 33730 2455 33735 2460
rect 33695 2450 33735 2455
rect 33975 2455 33980 2460
rect 34010 2455 34015 2485
rect 33975 2450 34015 2455
rect 32695 2440 32735 2445
rect 31365 2420 31405 2425
rect 31365 2390 31370 2420
rect 31400 2415 31405 2420
rect 31880 2420 31920 2425
rect 31880 2415 31885 2420
rect 31400 2395 31885 2415
rect 31400 2390 31405 2395
rect 31365 2385 31405 2390
rect 31880 2390 31885 2395
rect 31915 2415 31920 2420
rect 32395 2420 32435 2425
rect 32395 2415 32400 2420
rect 31915 2395 32400 2415
rect 31915 2390 31920 2395
rect 31880 2385 31920 2390
rect 32395 2390 32400 2395
rect 32430 2390 32435 2420
rect 32395 2385 32435 2390
rect 30450 2375 30490 2380
rect 30450 2345 30455 2375
rect 30485 2370 30490 2375
rect 30740 2375 30780 2380
rect 30740 2370 30745 2375
rect 30485 2350 30745 2370
rect 30485 2345 30490 2350
rect 30450 2340 30490 2345
rect 30740 2345 30745 2350
rect 30775 2370 30780 2375
rect 31670 2375 31710 2380
rect 31670 2370 31675 2375
rect 30775 2350 31675 2370
rect 30775 2345 30780 2350
rect 30740 2340 30780 2345
rect 31670 2345 31675 2350
rect 31705 2345 31710 2375
rect 31670 2340 31710 2345
rect 32090 2375 32130 2380
rect 32090 2345 32095 2375
rect 32125 2370 32130 2375
rect 33040 2375 33080 2380
rect 33040 2370 33045 2375
rect 32125 2350 33045 2370
rect 32125 2345 32130 2350
rect 32090 2340 32130 2345
rect 33040 2345 33045 2350
rect 33075 2370 33080 2375
rect 33310 2375 33350 2380
rect 33310 2370 33315 2375
rect 33075 2350 33315 2370
rect 33075 2345 33080 2350
rect 33040 2340 33080 2345
rect 33310 2345 33315 2350
rect 33345 2345 33350 2375
rect 33310 2340 33350 2345
rect 30875 2330 30915 2335
rect 30875 2300 30880 2330
rect 30910 2325 30915 2330
rect 32870 2330 32910 2335
rect 32870 2325 32875 2330
rect 30910 2305 32875 2325
rect 30910 2300 30915 2305
rect 29835 2295 29875 2300
rect 29310 2260 29360 2270
rect 29835 2265 29840 2295
rect 29870 2290 29875 2295
rect 30065 2295 30105 2300
rect 30065 2290 30070 2295
rect 29870 2270 30070 2290
rect 29870 2265 29875 2270
rect 29835 2260 29875 2265
rect 30065 2265 30070 2270
rect 30100 2290 30105 2295
rect 30175 2295 30215 2300
rect 30175 2290 30180 2295
rect 30100 2270 30180 2290
rect 30100 2265 30105 2270
rect 30065 2260 30105 2265
rect 30175 2265 30180 2270
rect 30210 2290 30215 2295
rect 30285 2295 30325 2300
rect 30285 2290 30290 2295
rect 30210 2270 30290 2290
rect 30210 2265 30215 2270
rect 30175 2260 30215 2265
rect 30285 2265 30290 2270
rect 30320 2290 30325 2295
rect 30395 2295 30435 2300
rect 30395 2290 30400 2295
rect 30320 2270 30400 2290
rect 30320 2265 30325 2270
rect 30285 2260 30325 2265
rect 30395 2265 30400 2270
rect 30430 2290 30435 2295
rect 30505 2295 30545 2300
rect 30875 2295 30915 2300
rect 32870 2300 32875 2305
rect 32905 2300 32910 2330
rect 32870 2295 32910 2300
rect 33255 2295 33295 2300
rect 30505 2290 30510 2295
rect 30430 2270 30510 2290
rect 30430 2265 30435 2270
rect 30395 2260 30435 2265
rect 30505 2265 30510 2270
rect 30540 2265 30545 2295
rect 30505 2260 30545 2265
rect 31240 2285 31280 2290
rect 29310 2230 29320 2260
rect 29350 2230 29360 2260
rect 31240 2255 31245 2285
rect 31275 2280 31280 2285
rect 31350 2285 31390 2290
rect 31350 2280 31355 2285
rect 31275 2260 31355 2280
rect 31275 2255 31280 2260
rect 31240 2250 31280 2255
rect 31350 2255 31355 2260
rect 31385 2280 31390 2285
rect 31460 2285 31500 2290
rect 31460 2280 31465 2285
rect 31385 2260 31465 2280
rect 31385 2255 31390 2260
rect 31350 2250 31390 2255
rect 31460 2255 31465 2260
rect 31495 2280 31500 2285
rect 31570 2285 31610 2290
rect 31570 2280 31575 2285
rect 31495 2260 31575 2280
rect 31495 2255 31500 2260
rect 31460 2250 31500 2255
rect 31570 2255 31575 2260
rect 31605 2280 31610 2285
rect 31680 2285 31720 2290
rect 31680 2280 31685 2285
rect 31605 2260 31685 2280
rect 31605 2255 31610 2260
rect 31570 2250 31610 2255
rect 31680 2255 31685 2260
rect 31715 2280 31720 2285
rect 31790 2285 31830 2290
rect 31790 2280 31795 2285
rect 31715 2260 31795 2280
rect 31715 2255 31720 2260
rect 31680 2250 31720 2255
rect 31790 2255 31795 2260
rect 31825 2255 31830 2285
rect 31790 2250 31830 2255
rect 31970 2285 32010 2290
rect 31970 2255 31975 2285
rect 32005 2280 32010 2285
rect 32080 2285 32120 2290
rect 32080 2280 32085 2285
rect 32005 2260 32085 2280
rect 32005 2255 32010 2260
rect 31970 2250 32010 2255
rect 32080 2255 32085 2260
rect 32115 2280 32120 2285
rect 32190 2285 32230 2290
rect 32190 2280 32195 2285
rect 32115 2260 32195 2280
rect 32115 2255 32120 2260
rect 32080 2250 32120 2255
rect 32190 2255 32195 2260
rect 32225 2280 32230 2285
rect 32300 2285 32340 2290
rect 32300 2280 32305 2285
rect 32225 2260 32305 2280
rect 32225 2255 32230 2260
rect 32190 2250 32230 2255
rect 32300 2255 32305 2260
rect 32335 2280 32340 2285
rect 32410 2285 32450 2290
rect 32410 2280 32415 2285
rect 32335 2260 32415 2280
rect 32335 2255 32340 2260
rect 32300 2250 32340 2255
rect 32410 2255 32415 2260
rect 32445 2280 32450 2285
rect 32520 2285 32560 2290
rect 32520 2280 32525 2285
rect 32445 2260 32525 2280
rect 32445 2255 32450 2260
rect 32410 2250 32450 2255
rect 32520 2255 32525 2260
rect 32555 2255 32560 2285
rect 33255 2265 33260 2295
rect 33290 2290 33295 2295
rect 33365 2295 33405 2300
rect 33365 2290 33370 2295
rect 33290 2270 33370 2290
rect 33290 2265 33295 2270
rect 33255 2260 33295 2265
rect 33365 2265 33370 2270
rect 33400 2290 33405 2295
rect 33475 2295 33515 2300
rect 33475 2290 33480 2295
rect 33400 2270 33480 2290
rect 33400 2265 33405 2270
rect 33365 2260 33405 2265
rect 33475 2265 33480 2270
rect 33510 2290 33515 2295
rect 33585 2295 33625 2300
rect 33585 2290 33590 2295
rect 33510 2270 33590 2290
rect 33510 2265 33515 2270
rect 33475 2260 33515 2265
rect 33585 2265 33590 2270
rect 33620 2290 33625 2295
rect 33695 2295 33735 2300
rect 33695 2290 33700 2295
rect 33620 2270 33700 2290
rect 33620 2265 33625 2270
rect 33585 2260 33625 2265
rect 33695 2265 33700 2270
rect 33730 2290 33735 2295
rect 33930 2295 33970 2300
rect 33930 2290 33935 2295
rect 33730 2270 33935 2290
rect 33730 2265 33735 2270
rect 33695 2260 33735 2265
rect 33930 2265 33935 2270
rect 33965 2265 33970 2295
rect 33930 2260 33970 2265
rect 34440 2260 34490 2270
rect 32520 2250 32560 2255
rect 29310 2220 29360 2230
rect 30830 2230 30870 2235
rect 30830 2200 30835 2230
rect 30865 2225 30870 2230
rect 31520 2230 31550 2235
rect 30865 2205 31520 2225
rect 30865 2200 30870 2205
rect 30830 2195 30870 2200
rect 32250 2230 32280 2235
rect 31550 2205 32250 2225
rect 31520 2195 31550 2200
rect 34440 2230 34450 2260
rect 34480 2230 34490 2260
rect 34440 2220 34490 2230
rect 32250 2195 32280 2200
rect 29735 2110 29775 2115
rect 29735 2080 29740 2110
rect 29770 2105 29775 2110
rect 29885 2110 29925 2115
rect 29885 2105 29890 2110
rect 29770 2085 29890 2105
rect 29770 2080 29775 2085
rect 29735 2075 29775 2080
rect 29885 2080 29890 2085
rect 29920 2080 29925 2110
rect 29885 2075 29925 2080
rect 33875 2110 33915 2115
rect 33875 2080 33880 2110
rect 33910 2105 33915 2110
rect 34025 2110 34065 2115
rect 34025 2105 34030 2110
rect 33910 2085 34030 2105
rect 33910 2080 33915 2085
rect 33875 2075 33915 2080
rect 34025 2080 34030 2085
rect 34060 2080 34065 2110
rect 34025 2075 34065 2080
rect 29470 1985 29565 1990
rect 29505 1950 29530 1985
rect 29470 1945 29565 1950
rect 29590 1985 29625 1991
rect 29590 1945 29625 1950
rect 29650 1985 29685 1990
rect 34115 1985 34150 1990
rect 29790 1980 29830 1985
rect 29790 1975 29795 1980
rect 29685 1955 29795 1975
rect 29650 1945 29685 1950
rect 29790 1950 29795 1955
rect 29825 1950 29830 1980
rect 33975 1980 34015 1985
rect 29790 1945 29830 1950
rect 31295 1950 31335 1955
rect 29590 1925 29630 1930
rect 29590 1895 29595 1925
rect 29625 1920 29630 1925
rect 29835 1925 29875 1930
rect 29835 1920 29840 1925
rect 29625 1900 29840 1920
rect 29625 1895 29630 1900
rect 29590 1890 29630 1895
rect 29835 1895 29840 1900
rect 29870 1895 29875 1925
rect 29835 1890 29875 1895
rect 30010 1925 30050 1930
rect 30010 1895 30015 1925
rect 30045 1920 30050 1925
rect 30120 1925 30160 1930
rect 30120 1920 30125 1925
rect 30045 1900 30125 1920
rect 30045 1895 30050 1900
rect 30010 1890 30050 1895
rect 30120 1895 30125 1900
rect 30155 1920 30160 1925
rect 30230 1925 30270 1930
rect 30230 1920 30235 1925
rect 30155 1900 30235 1920
rect 30155 1895 30160 1900
rect 30120 1890 30160 1895
rect 30230 1895 30235 1900
rect 30265 1920 30270 1925
rect 30340 1925 30380 1930
rect 30340 1920 30345 1925
rect 30265 1900 30345 1920
rect 30265 1895 30270 1900
rect 30230 1890 30270 1895
rect 30340 1895 30345 1900
rect 30375 1920 30380 1925
rect 30450 1925 30490 1930
rect 30450 1920 30455 1925
rect 30375 1900 30455 1920
rect 30375 1895 30380 1900
rect 30340 1890 30380 1895
rect 30450 1895 30455 1900
rect 30485 1920 30490 1925
rect 30560 1925 30600 1930
rect 30560 1920 30565 1925
rect 30485 1900 30565 1920
rect 30485 1895 30490 1900
rect 30450 1890 30490 1895
rect 30560 1895 30565 1900
rect 30595 1920 30600 1925
rect 30785 1925 30825 1930
rect 30785 1920 30790 1925
rect 30595 1900 30790 1920
rect 30595 1895 30600 1900
rect 30560 1890 30600 1895
rect 30785 1895 30790 1900
rect 30820 1895 30825 1925
rect 31295 1920 31300 1950
rect 31330 1945 31335 1950
rect 31405 1950 31445 1955
rect 31405 1945 31410 1950
rect 31330 1925 31410 1945
rect 31330 1920 31335 1925
rect 31295 1915 31335 1920
rect 31405 1920 31410 1925
rect 31440 1945 31445 1950
rect 31515 1950 31555 1955
rect 31515 1945 31520 1950
rect 31440 1925 31520 1945
rect 31440 1920 31445 1925
rect 31405 1915 31445 1920
rect 31515 1920 31520 1925
rect 31550 1945 31555 1950
rect 31625 1950 31665 1955
rect 31625 1945 31630 1950
rect 31550 1925 31630 1945
rect 31550 1920 31555 1925
rect 31515 1915 31555 1920
rect 31625 1920 31630 1925
rect 31660 1945 31665 1950
rect 31735 1950 31775 1955
rect 31735 1945 31740 1950
rect 31660 1925 31740 1945
rect 31660 1920 31665 1925
rect 31625 1915 31665 1920
rect 31735 1920 31740 1925
rect 31770 1920 31775 1950
rect 31735 1915 31775 1920
rect 32025 1950 32065 1955
rect 32025 1920 32030 1950
rect 32060 1945 32065 1950
rect 32135 1950 32175 1955
rect 32135 1945 32140 1950
rect 32060 1925 32140 1945
rect 32060 1920 32065 1925
rect 32025 1915 32065 1920
rect 32135 1920 32140 1925
rect 32170 1945 32175 1950
rect 32245 1950 32285 1955
rect 32245 1945 32250 1950
rect 32170 1925 32250 1945
rect 32170 1920 32175 1925
rect 32135 1915 32175 1920
rect 32245 1920 32250 1925
rect 32280 1945 32285 1950
rect 32355 1950 32395 1955
rect 32355 1945 32360 1950
rect 32280 1925 32360 1945
rect 32280 1920 32285 1925
rect 32245 1915 32285 1920
rect 32355 1920 32360 1925
rect 32390 1945 32395 1950
rect 32465 1950 32505 1955
rect 32465 1945 32470 1950
rect 32390 1925 32470 1945
rect 32390 1920 32395 1925
rect 32355 1915 32395 1920
rect 32465 1920 32470 1925
rect 32500 1920 32505 1950
rect 33975 1950 33980 1980
rect 34010 1975 34015 1980
rect 34010 1955 34115 1975
rect 34010 1950 34015 1955
rect 33975 1945 34015 1950
rect 34115 1945 34150 1950
rect 34175 1985 34210 1991
rect 34295 1990 34330 1991
rect 34175 1945 34210 1950
rect 34235 1985 34330 1990
rect 34270 1950 34295 1985
rect 34235 1945 34330 1950
rect 32465 1915 32505 1920
rect 33005 1925 33045 1930
rect 30785 1890 30825 1895
rect 31190 1895 31230 1900
rect 31190 1865 31195 1895
rect 31225 1890 31230 1895
rect 31410 1895 31450 1900
rect 31410 1890 31415 1895
rect 31225 1870 31415 1890
rect 31225 1865 31230 1870
rect 31190 1860 31230 1865
rect 31410 1865 31415 1870
rect 31445 1890 31450 1895
rect 31640 1895 31680 1900
rect 31640 1890 31645 1895
rect 31445 1870 31645 1890
rect 31445 1865 31450 1870
rect 31410 1860 31450 1865
rect 31640 1865 31645 1870
rect 31675 1890 31680 1895
rect 32230 1895 32270 1900
rect 32230 1890 32235 1895
rect 31675 1870 32235 1890
rect 31675 1865 31680 1870
rect 31640 1860 31680 1865
rect 32230 1865 32235 1870
rect 32265 1890 32270 1895
rect 32450 1895 32490 1900
rect 32450 1890 32455 1895
rect 32265 1870 32455 1890
rect 32265 1865 32270 1870
rect 32230 1860 32270 1865
rect 32450 1865 32455 1870
rect 32485 1890 32490 1895
rect 32680 1895 32720 1900
rect 32680 1890 32685 1895
rect 32485 1870 32685 1890
rect 32485 1865 32490 1870
rect 32450 1860 32490 1865
rect 32680 1865 32685 1870
rect 32715 1865 32720 1895
rect 33005 1895 33010 1925
rect 33040 1920 33045 1925
rect 33200 1925 33240 1930
rect 33200 1920 33205 1925
rect 33040 1900 33205 1920
rect 33040 1895 33045 1900
rect 33005 1890 33045 1895
rect 33200 1895 33205 1900
rect 33235 1920 33240 1925
rect 33310 1925 33350 1930
rect 33310 1920 33315 1925
rect 33235 1900 33315 1920
rect 33235 1895 33240 1900
rect 33200 1890 33240 1895
rect 33310 1895 33315 1900
rect 33345 1920 33350 1925
rect 33420 1925 33460 1930
rect 33420 1920 33425 1925
rect 33345 1900 33425 1920
rect 33345 1895 33350 1900
rect 33310 1890 33350 1895
rect 33420 1895 33425 1900
rect 33455 1920 33460 1925
rect 33530 1925 33570 1930
rect 33530 1920 33535 1925
rect 33455 1900 33535 1920
rect 33455 1895 33460 1900
rect 33420 1890 33460 1895
rect 33530 1895 33535 1900
rect 33565 1920 33570 1925
rect 33640 1925 33680 1930
rect 33640 1920 33645 1925
rect 33565 1900 33645 1920
rect 33565 1895 33570 1900
rect 33530 1890 33570 1895
rect 33640 1895 33645 1900
rect 33675 1920 33680 1925
rect 33750 1925 33790 1930
rect 33750 1920 33755 1925
rect 33675 1900 33755 1920
rect 33675 1895 33680 1900
rect 33640 1890 33680 1895
rect 33750 1895 33755 1900
rect 33785 1895 33790 1925
rect 33750 1890 33790 1895
rect 33930 1925 33970 1930
rect 33930 1895 33935 1925
rect 33965 1920 33970 1925
rect 34170 1925 34210 1930
rect 34170 1920 34175 1925
rect 33965 1900 34175 1920
rect 33965 1895 33970 1900
rect 33930 1890 33970 1895
rect 34170 1895 34175 1900
rect 34205 1895 34210 1925
rect 34170 1890 34210 1895
rect 32680 1860 32720 1865
rect 31820 1850 31860 1855
rect 29470 1820 29510 1825
rect 29470 1790 29475 1820
rect 29505 1815 29510 1820
rect 30875 1820 30915 1825
rect 30875 1815 30880 1820
rect 29505 1795 30880 1815
rect 29505 1790 29510 1795
rect 29470 1785 29510 1790
rect 30875 1790 30880 1795
rect 30910 1790 30915 1820
rect 31820 1820 31825 1850
rect 31855 1845 31860 1850
rect 31940 1850 31980 1855
rect 31940 1845 31945 1850
rect 31855 1825 31945 1845
rect 31855 1820 31860 1825
rect 31820 1815 31860 1820
rect 31940 1820 31945 1825
rect 31975 1820 31980 1850
rect 31940 1815 31980 1820
rect 32870 1825 32910 1830
rect 30875 1785 30915 1790
rect 31085 1805 31125 1810
rect 31085 1775 31090 1805
rect 31120 1800 31125 1805
rect 31305 1805 31345 1810
rect 31305 1800 31310 1805
rect 31120 1780 31310 1800
rect 31120 1775 31125 1780
rect 31085 1770 31125 1775
rect 31305 1775 31310 1780
rect 31340 1800 31345 1805
rect 31525 1805 31565 1810
rect 31525 1800 31530 1805
rect 31340 1780 31530 1800
rect 31340 1775 31345 1780
rect 31305 1770 31345 1775
rect 31525 1775 31530 1780
rect 31560 1800 31565 1805
rect 32125 1805 32165 1810
rect 32125 1800 32130 1805
rect 31560 1780 32130 1800
rect 31560 1775 31565 1780
rect 31525 1770 31565 1775
rect 32125 1775 32130 1780
rect 32160 1800 32165 1805
rect 32345 1805 32385 1810
rect 32345 1800 32350 1805
rect 32160 1780 32350 1800
rect 32160 1775 32165 1780
rect 32125 1770 32165 1775
rect 32345 1775 32350 1780
rect 32380 1800 32385 1805
rect 32565 1805 32605 1810
rect 32565 1800 32570 1805
rect 32380 1780 32570 1800
rect 32380 1775 32385 1780
rect 32345 1770 32385 1775
rect 32565 1775 32570 1780
rect 32600 1775 32605 1805
rect 32870 1795 32875 1825
rect 32905 1820 32910 1825
rect 34290 1825 34330 1830
rect 34290 1820 34295 1825
rect 32905 1800 34295 1820
rect 32905 1795 32910 1800
rect 32870 1790 32910 1795
rect 34290 1795 34295 1800
rect 34325 1795 34330 1825
rect 34290 1790 34330 1795
rect 32565 1770 32605 1775
rect 29725 1760 29765 1765
rect 29725 1730 29730 1760
rect 29760 1755 29765 1760
rect 30435 1760 30475 1765
rect 30435 1755 30440 1760
rect 29760 1735 30440 1755
rect 29760 1730 29765 1735
rect 29725 1725 29765 1730
rect 30435 1730 30440 1735
rect 30470 1755 30475 1760
rect 30740 1760 30780 1765
rect 30740 1755 30745 1760
rect 30470 1735 30745 1755
rect 30470 1730 30475 1735
rect 30435 1725 30475 1730
rect 30740 1730 30745 1735
rect 30775 1730 30780 1760
rect 31237 1760 31269 1765
rect 31237 1755 31240 1760
rect 30920 1735 31240 1755
rect 30740 1725 30780 1730
rect 31237 1730 31240 1735
rect 31266 1755 31269 1760
rect 31457 1760 31489 1765
rect 31457 1755 31460 1760
rect 31266 1735 31460 1755
rect 31266 1730 31269 1735
rect 31237 1725 31269 1730
rect 31457 1730 31460 1735
rect 31486 1755 31489 1760
rect 31601 1760 31633 1765
rect 31601 1755 31604 1760
rect 31486 1735 31604 1755
rect 31486 1730 31489 1735
rect 31457 1725 31489 1730
rect 31601 1730 31604 1735
rect 31630 1755 31633 1760
rect 31867 1760 31899 1765
rect 31867 1755 31870 1760
rect 31630 1735 31870 1755
rect 31630 1730 31633 1735
rect 31601 1725 31633 1730
rect 31867 1730 31870 1735
rect 31896 1755 31899 1760
rect 32277 1760 32309 1765
rect 32277 1755 32280 1760
rect 31896 1735 32280 1755
rect 31896 1730 31899 1735
rect 31867 1725 31899 1730
rect 32277 1730 32280 1735
rect 32306 1755 32309 1760
rect 32497 1760 32529 1765
rect 32497 1755 32500 1760
rect 32306 1735 32500 1755
rect 32306 1730 32309 1735
rect 32277 1725 32309 1730
rect 32497 1730 32500 1735
rect 32526 1755 32529 1760
rect 32641 1760 32673 1765
rect 32641 1755 32644 1760
rect 32526 1735 32644 1755
rect 32526 1730 32529 1735
rect 32497 1725 32529 1730
rect 32641 1730 32644 1735
rect 32670 1730 32673 1760
rect 32641 1725 32673 1730
rect 33015 1760 33055 1765
rect 33015 1730 33020 1760
rect 33050 1755 33055 1760
rect 33325 1760 33365 1765
rect 33325 1755 33330 1760
rect 33050 1735 33330 1755
rect 33050 1730 33055 1735
rect 33015 1725 33055 1730
rect 33325 1730 33330 1735
rect 33360 1755 33365 1760
rect 34035 1760 34075 1765
rect 34035 1755 34040 1760
rect 33360 1735 34040 1755
rect 33360 1730 33365 1735
rect 33325 1725 33365 1730
rect 34035 1730 34040 1735
rect 34070 1730 34075 1760
rect 34035 1725 34075 1730
rect 29315 1705 29355 1710
rect 29315 1675 29320 1705
rect 29350 1700 29355 1705
rect 29790 1705 29830 1710
rect 29790 1700 29795 1705
rect 29350 1680 29795 1700
rect 29350 1675 29355 1680
rect 29315 1670 29355 1675
rect 29790 1675 29795 1680
rect 29825 1700 29830 1705
rect 30135 1705 30175 1710
rect 30135 1700 30140 1705
rect 29825 1680 30140 1700
rect 29825 1675 29830 1680
rect 29790 1670 29830 1675
rect 30135 1675 30140 1680
rect 30170 1700 30175 1705
rect 30335 1705 30375 1710
rect 30335 1700 30340 1705
rect 30170 1680 30340 1700
rect 30170 1675 30175 1680
rect 30135 1670 30175 1675
rect 30335 1675 30340 1680
rect 30370 1700 30375 1705
rect 30535 1705 30575 1710
rect 30535 1700 30540 1705
rect 30370 1680 30540 1700
rect 30370 1675 30375 1680
rect 30335 1670 30375 1675
rect 30535 1675 30540 1680
rect 30570 1675 30575 1705
rect 30535 1670 30575 1675
rect 33225 1705 33265 1710
rect 33225 1675 33230 1705
rect 33260 1700 33265 1705
rect 33425 1705 33465 1710
rect 33425 1700 33430 1705
rect 33260 1680 33430 1700
rect 33260 1675 33265 1680
rect 33225 1670 33265 1675
rect 33425 1675 33430 1680
rect 33460 1700 33465 1705
rect 33625 1705 33665 1710
rect 33625 1700 33630 1705
rect 33460 1680 33630 1700
rect 33460 1675 33465 1680
rect 33425 1670 33465 1675
rect 33625 1675 33630 1680
rect 33660 1700 33665 1705
rect 33970 1705 34010 1710
rect 33970 1700 33975 1705
rect 33660 1680 33975 1700
rect 33660 1675 33665 1680
rect 33625 1670 33665 1675
rect 33970 1675 33975 1680
rect 34005 1700 34010 1705
rect 34445 1705 34485 1710
rect 34445 1700 34450 1705
rect 34005 1680 34450 1700
rect 34005 1675 34010 1680
rect 33970 1670 34010 1675
rect 34445 1675 34450 1680
rect 34480 1675 34485 1705
rect 34445 1670 34485 1675
rect 30785 1650 30825 1655
rect 29730 1645 29765 1650
rect 29730 1605 29765 1610
rect 29790 1645 29825 1650
rect 30785 1620 30790 1650
rect 30820 1645 30825 1650
rect 30940 1650 30980 1655
rect 30940 1645 30945 1650
rect 30820 1625 30945 1645
rect 30820 1620 30825 1625
rect 30785 1615 30825 1620
rect 30940 1620 30945 1625
rect 30975 1620 30980 1650
rect 30940 1615 30980 1620
rect 33975 1645 34010 1650
rect 29790 1605 29825 1610
rect 33975 1605 34010 1610
rect 34035 1645 34070 1650
rect 34035 1605 34070 1610
rect 31106 1540 31138 1545
rect 31106 1535 31109 1540
rect 30920 1515 31109 1535
rect 31106 1510 31109 1515
rect 31135 1535 31138 1540
rect 31305 1540 31345 1545
rect 31305 1535 31310 1540
rect 31135 1515 31310 1535
rect 31135 1510 31138 1515
rect 31106 1505 31138 1510
rect 31305 1510 31310 1515
rect 31340 1535 31345 1540
rect 31525 1540 31565 1545
rect 31525 1535 31530 1540
rect 31340 1515 31530 1535
rect 31340 1510 31345 1515
rect 31305 1505 31345 1510
rect 31525 1510 31530 1515
rect 31560 1535 31565 1540
rect 31922 1540 31954 1545
rect 31922 1535 31925 1540
rect 31560 1515 31925 1535
rect 31560 1510 31565 1515
rect 31525 1505 31565 1510
rect 31922 1510 31925 1515
rect 31951 1535 31954 1540
rect 32146 1540 32178 1545
rect 32146 1535 32149 1540
rect 31951 1515 32149 1535
rect 31951 1510 31954 1515
rect 31922 1505 31954 1510
rect 32146 1510 32149 1515
rect 32175 1535 32178 1540
rect 32345 1540 32385 1545
rect 32345 1535 32350 1540
rect 32175 1515 32350 1535
rect 32175 1510 32178 1515
rect 32146 1505 32178 1510
rect 32345 1510 32350 1515
rect 32380 1535 32385 1540
rect 32565 1540 32605 1545
rect 32565 1535 32570 1540
rect 32380 1515 32570 1535
rect 32380 1510 32385 1515
rect 32345 1505 32385 1510
rect 32565 1510 32570 1515
rect 32600 1510 32605 1540
rect 32565 1505 32605 1510
rect 31145 1480 31185 1485
rect 31145 1450 31150 1480
rect 31180 1475 31185 1480
rect 31250 1480 31290 1485
rect 31250 1475 31255 1480
rect 31180 1455 31255 1475
rect 31180 1450 31185 1455
rect 31145 1445 31185 1450
rect 31250 1450 31255 1455
rect 31285 1475 31290 1480
rect 31360 1480 31400 1485
rect 31360 1475 31365 1480
rect 31285 1455 31365 1475
rect 31285 1450 31290 1455
rect 31250 1445 31290 1450
rect 31360 1450 31365 1455
rect 31395 1475 31400 1480
rect 31470 1480 31510 1485
rect 31470 1475 31475 1480
rect 31395 1455 31475 1475
rect 31395 1450 31400 1455
rect 31360 1445 31400 1450
rect 31470 1450 31475 1455
rect 31505 1475 31510 1480
rect 31580 1480 31620 1485
rect 31580 1475 31585 1480
rect 31505 1455 31585 1475
rect 31505 1450 31510 1455
rect 31470 1445 31510 1450
rect 31580 1450 31585 1455
rect 31615 1475 31620 1480
rect 32185 1480 32225 1485
rect 32185 1475 32190 1480
rect 31615 1455 32190 1475
rect 31615 1450 31620 1455
rect 31580 1445 31620 1450
rect 32185 1450 32190 1455
rect 32220 1475 32225 1480
rect 32290 1480 32330 1485
rect 32290 1475 32295 1480
rect 32220 1455 32295 1475
rect 32220 1450 32225 1455
rect 32185 1445 32225 1450
rect 32290 1450 32295 1455
rect 32325 1475 32330 1480
rect 32400 1480 32440 1485
rect 32400 1475 32405 1480
rect 32325 1455 32405 1475
rect 32325 1450 32330 1455
rect 32290 1445 32330 1450
rect 32400 1450 32405 1455
rect 32435 1475 32440 1480
rect 32510 1480 32550 1485
rect 32510 1475 32515 1480
rect 32435 1455 32515 1475
rect 32435 1450 32440 1455
rect 32400 1445 32440 1450
rect 32510 1450 32515 1455
rect 32545 1475 32550 1480
rect 32620 1480 32660 1485
rect 32620 1475 32625 1480
rect 32545 1455 32625 1475
rect 32545 1450 32550 1455
rect 32510 1445 32550 1450
rect 32620 1450 32625 1455
rect 32655 1450 32660 1480
rect 32620 1445 32660 1450
rect 30740 1435 30780 1440
rect 30740 1405 30745 1435
rect 30775 1430 30780 1435
rect 33015 1435 33055 1440
rect 33015 1430 33020 1435
rect 30775 1410 33020 1430
rect 30775 1405 30780 1410
rect 30740 1400 30780 1405
rect 33015 1405 33020 1410
rect 33050 1405 33055 1435
rect 33015 1400 33055 1405
rect 31005 1390 31045 1395
rect 31005 1360 31010 1390
rect 31040 1385 31045 1390
rect 31755 1390 31795 1395
rect 31755 1385 31760 1390
rect 31040 1365 31760 1385
rect 31040 1360 31045 1365
rect 31005 1355 31045 1360
rect 31755 1360 31760 1365
rect 31790 1360 31795 1390
rect 31755 1355 31795 1360
rect 32375 1365 32415 1370
rect 31315 1345 31355 1350
rect 29875 1320 29915 1325
rect 29875 1290 29880 1320
rect 29910 1315 29915 1320
rect 29965 1320 30005 1325
rect 29965 1315 29970 1320
rect 29910 1295 29970 1315
rect 29910 1290 29915 1295
rect 29875 1285 29915 1290
rect 29965 1290 29970 1295
rect 30000 1290 30005 1320
rect 31315 1315 31320 1345
rect 31350 1340 31355 1345
rect 31870 1345 31910 1350
rect 31870 1340 31875 1345
rect 31350 1320 31875 1340
rect 31350 1315 31355 1320
rect 31315 1310 31355 1315
rect 31870 1315 31875 1320
rect 31905 1315 31910 1345
rect 32375 1335 32380 1365
rect 32410 1360 32415 1365
rect 32915 1365 32955 1370
rect 32915 1360 32920 1365
rect 32410 1340 32920 1360
rect 32410 1335 32415 1340
rect 32375 1330 32415 1335
rect 32915 1335 32920 1340
rect 32950 1335 32955 1365
rect 32915 1330 32955 1335
rect 31870 1310 31910 1315
rect 33795 1320 33835 1325
rect 29965 1285 30005 1290
rect 33795 1290 33800 1320
rect 33830 1315 33835 1320
rect 33885 1320 33925 1325
rect 33885 1315 33890 1320
rect 33830 1295 33890 1315
rect 33830 1290 33835 1295
rect 33795 1285 33835 1290
rect 33885 1290 33890 1295
rect 33920 1290 33925 1320
rect 33885 1285 33925 1290
rect 31425 1255 31465 1260
rect 31425 1225 31430 1255
rect 31460 1250 31465 1255
rect 31535 1255 31575 1260
rect 31535 1250 31540 1255
rect 31460 1230 31540 1250
rect 31460 1225 31465 1230
rect 31425 1220 31465 1225
rect 31535 1225 31540 1230
rect 31570 1250 31575 1255
rect 31645 1255 31685 1260
rect 31645 1250 31650 1255
rect 31570 1230 31650 1250
rect 31570 1225 31575 1230
rect 31535 1220 31575 1225
rect 31645 1225 31650 1230
rect 31680 1250 31685 1255
rect 31755 1255 31795 1260
rect 31755 1250 31760 1255
rect 31680 1230 31760 1250
rect 31680 1225 31685 1230
rect 31645 1220 31685 1225
rect 31755 1225 31760 1230
rect 31790 1250 31795 1255
rect 31865 1255 31905 1260
rect 31865 1250 31870 1255
rect 31790 1230 31870 1250
rect 31790 1225 31795 1230
rect 31755 1220 31795 1225
rect 31865 1225 31870 1230
rect 31900 1250 31905 1255
rect 31975 1255 32015 1260
rect 31975 1250 31980 1255
rect 31900 1230 31980 1250
rect 31900 1225 31905 1230
rect 31865 1220 31905 1225
rect 31975 1225 31980 1230
rect 32010 1250 32015 1255
rect 32085 1255 32125 1260
rect 32085 1250 32090 1255
rect 32010 1230 32090 1250
rect 32010 1225 32015 1230
rect 31975 1220 32015 1225
rect 32085 1225 32090 1230
rect 32120 1250 32125 1255
rect 32195 1255 32235 1260
rect 32195 1250 32200 1255
rect 32120 1230 32200 1250
rect 32120 1225 32125 1230
rect 32085 1220 32125 1225
rect 32195 1225 32200 1230
rect 32230 1250 32235 1255
rect 32305 1255 32345 1260
rect 32305 1250 32310 1255
rect 32230 1230 32310 1250
rect 32230 1225 32235 1230
rect 32195 1220 32235 1225
rect 32305 1225 32310 1230
rect 32340 1250 32345 1255
rect 32430 1255 32470 1260
rect 32430 1250 32435 1255
rect 32340 1230 32435 1250
rect 32340 1225 32345 1230
rect 32305 1220 32345 1225
rect 32430 1225 32435 1230
rect 32465 1225 32470 1255
rect 32430 1220 32470 1225
rect 30235 935 30275 940
rect 30235 905 30240 935
rect 30270 930 30275 935
rect 30335 935 30375 940
rect 30335 930 30340 935
rect 30270 910 30340 930
rect 30270 905 30275 910
rect 30235 900 30275 905
rect 30335 905 30340 910
rect 30370 930 30375 935
rect 30435 935 30475 940
rect 30435 930 30440 935
rect 30370 910 30440 930
rect 30370 905 30375 910
rect 30335 900 30375 905
rect 30435 905 30440 910
rect 30470 930 30475 935
rect 30785 935 30825 940
rect 30785 930 30790 935
rect 30470 910 30790 930
rect 30470 905 30475 910
rect 30435 900 30475 905
rect 30785 905 30790 910
rect 30820 930 30825 935
rect 31195 935 31235 940
rect 31195 930 31200 935
rect 30820 910 31200 930
rect 30820 905 30825 910
rect 30785 900 30825 905
rect 31195 905 31200 910
rect 31230 930 31235 935
rect 31260 935 31300 940
rect 31260 930 31265 935
rect 31230 910 31265 930
rect 31230 905 31235 910
rect 31195 900 31235 905
rect 31260 905 31265 910
rect 31295 930 31300 935
rect 31370 935 31410 940
rect 31370 930 31375 935
rect 31295 910 31375 930
rect 31295 905 31300 910
rect 31260 900 31300 905
rect 31370 905 31375 910
rect 31405 930 31410 935
rect 31480 935 31520 940
rect 31480 930 31485 935
rect 31405 910 31485 930
rect 31405 905 31410 910
rect 31370 900 31410 905
rect 31480 905 31485 910
rect 31515 930 31520 935
rect 31590 935 31630 940
rect 31590 930 31595 935
rect 31515 910 31595 930
rect 31515 905 31520 910
rect 31480 900 31520 905
rect 31590 905 31595 910
rect 31625 930 31630 935
rect 31700 935 31740 940
rect 31700 930 31705 935
rect 31625 910 31705 930
rect 31625 905 31630 910
rect 31590 900 31630 905
rect 31700 905 31705 910
rect 31735 930 31740 935
rect 31810 935 31850 940
rect 31810 930 31815 935
rect 31735 910 31815 930
rect 31735 905 31740 910
rect 31700 900 31740 905
rect 31810 905 31815 910
rect 31845 930 31850 935
rect 31920 935 31960 940
rect 31920 930 31925 935
rect 31845 910 31925 930
rect 31845 905 31850 910
rect 31810 900 31850 905
rect 31920 905 31925 910
rect 31955 930 31960 935
rect 32030 935 32070 940
rect 32030 930 32035 935
rect 31955 910 32035 930
rect 31955 905 31960 910
rect 31920 900 31960 905
rect 32030 905 32035 910
rect 32065 930 32070 935
rect 32140 935 32180 940
rect 32140 930 32145 935
rect 32065 910 32145 930
rect 32065 905 32070 910
rect 32030 900 32070 905
rect 32140 905 32145 910
rect 32175 930 32180 935
rect 32250 935 32290 940
rect 32250 930 32255 935
rect 32175 910 32255 930
rect 32175 905 32180 910
rect 32140 900 32180 905
rect 32250 905 32255 910
rect 32285 930 32290 935
rect 32360 935 32400 940
rect 32360 930 32365 935
rect 32285 910 32365 930
rect 32285 905 32290 910
rect 32250 900 32290 905
rect 32360 905 32365 910
rect 32395 930 32400 935
rect 32475 935 32515 940
rect 32475 930 32480 935
rect 32395 910 32480 930
rect 32395 905 32400 910
rect 32360 900 32400 905
rect 32475 905 32480 910
rect 32510 905 32515 935
rect 32475 900 32515 905
rect 33015 935 33055 940
rect 33015 905 33020 935
rect 33050 930 33055 935
rect 33325 935 33365 940
rect 33325 930 33330 935
rect 33050 910 33330 930
rect 33050 905 33055 910
rect 33015 900 33055 905
rect 33325 905 33330 910
rect 33360 930 33365 935
rect 33425 935 33465 940
rect 33425 930 33430 935
rect 33360 910 33430 930
rect 33360 905 33365 910
rect 33325 900 33365 905
rect 33425 905 33430 910
rect 33460 930 33465 935
rect 33525 935 33565 940
rect 33525 930 33530 935
rect 33460 910 33530 930
rect 33460 905 33465 910
rect 33425 900 33465 905
rect 33525 905 33530 910
rect 33560 905 33565 935
rect 33525 900 33565 905
rect 30335 875 30375 880
rect 30335 845 30340 875
rect 30370 845 30375 875
rect 33425 875 33465 880
rect 30335 840 30375 845
rect 30785 860 30825 865
rect 30785 830 30790 860
rect 30820 830 30825 860
rect 33425 845 33430 875
rect 33460 845 33465 875
rect 30785 825 30825 830
rect 31005 840 31045 845
rect 31005 810 31010 840
rect 31040 835 31045 840
rect 31505 840 31545 845
rect 31505 835 31510 840
rect 31040 815 31510 835
rect 31040 810 31045 815
rect 31005 805 31045 810
rect 31505 810 31510 815
rect 31540 810 31545 840
rect 31505 805 31545 810
rect 31935 840 31975 845
rect 31935 810 31940 840
rect 31970 835 31975 840
rect 32155 840 32195 845
rect 32155 835 32160 840
rect 31970 815 32160 835
rect 31970 810 31975 815
rect 31935 805 31975 810
rect 32155 810 32160 815
rect 32190 835 32195 840
rect 32375 840 32415 845
rect 32375 835 32380 840
rect 32190 815 32380 835
rect 32190 810 32195 815
rect 32155 805 32195 810
rect 32375 810 32380 815
rect 32410 835 32415 840
rect 32960 840 33000 845
rect 33425 840 33465 845
rect 32960 835 32965 840
rect 32410 815 32965 835
rect 32410 810 32415 815
rect 32375 805 32415 810
rect 32960 810 32965 815
rect 32995 810 33000 840
rect 32960 805 33000 810
rect 30830 740 30870 745
rect 30830 710 30835 740
rect 30865 735 30870 740
rect 31305 740 31345 745
rect 31305 735 31310 740
rect 30865 715 31310 735
rect 30865 710 30870 715
rect 30830 705 30870 710
rect 31305 710 31310 715
rect 31340 735 31345 740
rect 31375 740 31415 745
rect 31375 735 31380 740
rect 31340 715 31380 735
rect 31340 710 31345 715
rect 31305 705 31345 710
rect 31375 710 31380 715
rect 31410 735 31415 740
rect 31445 740 31485 745
rect 31445 735 31450 740
rect 31410 715 31450 735
rect 31410 710 31415 715
rect 31375 705 31415 710
rect 31445 710 31450 715
rect 31480 710 31485 740
rect 31445 705 31485 710
rect 32045 735 32085 740
rect 32045 705 32050 735
rect 32080 730 32085 735
rect 32265 735 32305 740
rect 32265 730 32270 735
rect 32080 710 32270 730
rect 32080 705 32085 710
rect 32045 700 32085 705
rect 32265 705 32270 710
rect 32300 730 32305 735
rect 32485 735 32525 740
rect 32485 730 32490 735
rect 32300 710 32490 730
rect 32300 705 32305 710
rect 32265 700 32305 705
rect 32485 705 32490 710
rect 32520 730 32525 735
rect 32915 735 32955 740
rect 32915 730 32920 735
rect 32520 710 32920 730
rect 32520 705 32525 710
rect 32485 700 32525 705
rect 32915 705 32920 710
rect 32950 705 32955 735
rect 32915 700 32955 705
rect 31990 615 32030 620
rect 31990 585 31995 615
rect 32025 610 32030 615
rect 32100 615 32140 620
rect 32100 610 32105 615
rect 32025 590 32105 610
rect 32025 585 32030 590
rect 31990 580 32030 585
rect 32100 585 32105 590
rect 32135 610 32140 615
rect 32210 615 32250 620
rect 32210 610 32215 615
rect 32135 590 32215 610
rect 32135 585 32140 590
rect 32100 580 32140 585
rect 32210 585 32215 590
rect 32245 610 32250 615
rect 32320 615 32360 620
rect 32320 610 32325 615
rect 32245 590 32325 610
rect 32245 585 32250 590
rect 32210 580 32250 585
rect 32320 585 32325 590
rect 32355 610 32360 615
rect 32430 615 32470 620
rect 32430 610 32435 615
rect 32355 590 32435 610
rect 32355 585 32360 590
rect 32320 580 32360 585
rect 32430 585 32435 590
rect 32465 585 32470 615
rect 32430 580 32470 585
rect 29265 495 29305 500
rect 29265 465 29270 495
rect 29300 490 29305 495
rect 30785 495 30825 500
rect 30785 490 30790 495
rect 29300 470 30790 490
rect 29300 465 29305 470
rect 29265 460 29305 465
rect 30785 465 30790 470
rect 30820 490 30825 495
rect 31375 495 31415 500
rect 31375 490 31380 495
rect 30820 470 31380 490
rect 30820 465 30825 470
rect 30785 460 30825 465
rect 31375 465 31380 470
rect 31410 490 31415 495
rect 32210 495 32250 500
rect 32210 490 32215 495
rect 31410 470 32215 490
rect 31410 465 31415 470
rect 31375 460 31415 465
rect 32210 465 32215 470
rect 32245 490 32250 495
rect 33015 495 33055 500
rect 33015 490 33020 495
rect 32245 470 33020 490
rect 32245 465 32250 470
rect 32210 460 32250 465
rect 33015 465 33020 470
rect 33050 490 33055 495
rect 34495 495 34535 500
rect 34495 490 34500 495
rect 33050 470 34500 490
rect 33050 465 33055 470
rect 33015 460 33055 465
rect 34495 465 34500 470
rect 34530 465 34535 495
rect 34495 460 34535 465
rect 30785 -515 30825 -510
rect 30785 -545 30790 -515
rect 30820 -545 30825 -515
rect 30785 -550 30825 -545
<< via2 >>
rect 30790 6155 30820 6185
rect 29610 3705 29640 3735
rect 34160 3705 34190 3735
rect 29320 2230 29350 2260
rect 34450 2230 34480 2260
rect 30790 -545 30820 -515
<< metal3 >>
rect 30780 6190 30830 6195
rect 30780 6150 30785 6190
rect 30825 6150 30830 6190
rect 30780 6145 30830 6150
rect 27410 5770 27640 5855
rect 27760 5770 27990 5855
rect 28110 5770 28340 5855
rect 27410 5720 28340 5770
rect 27410 5625 27640 5720
rect 27760 5625 27990 5720
rect 28110 5625 28340 5720
rect 28460 5625 28690 5855
rect 28810 5625 29040 5855
rect 29160 5625 29390 5855
rect 29510 5625 29740 5855
rect 29860 5625 30090 5855
rect 30210 5625 30440 5855
rect 30560 5625 30790 5855
rect 30910 5625 31140 5855
rect 31260 5625 31490 5855
rect 31610 5625 31840 5855
rect 31960 5625 32190 5855
rect 32310 5625 32540 5855
rect 32660 5625 32890 5855
rect 33010 5625 33240 5855
rect 33360 5625 33590 5855
rect 33710 5625 33940 5855
rect 34060 5625 34290 5855
rect 34410 5625 34640 5855
rect 34760 5625 34990 5855
rect 35110 5625 35340 5855
rect 35460 5770 35690 5855
rect 35810 5770 36040 5855
rect 36160 5770 36390 5855
rect 35460 5720 36390 5770
rect 35460 5625 35690 5720
rect 35810 5625 36040 5720
rect 36160 5625 36390 5720
rect 28200 5505 28250 5625
rect 28550 5505 28600 5625
rect 28900 5505 28950 5625
rect 29250 5505 29300 5625
rect 29600 5505 29650 5625
rect 29950 5505 30000 5625
rect 30300 5505 30350 5625
rect 30650 5505 30700 5625
rect 31000 5505 31050 5625
rect 31350 5505 31400 5625
rect 31700 5505 31750 5625
rect 32050 5505 32100 5625
rect 32400 5505 32450 5625
rect 32750 5505 32800 5625
rect 33100 5505 33150 5625
rect 33450 5505 33500 5625
rect 33800 5505 33850 5625
rect 34150 5505 34200 5625
rect 34500 5505 34550 5625
rect 34850 5505 34900 5625
rect 35200 5505 35250 5625
rect 35550 5505 35600 5625
rect 27410 5420 27640 5505
rect 27760 5420 27990 5505
rect 28110 5420 28340 5505
rect 28460 5420 28690 5505
rect 28810 5420 29040 5505
rect 29160 5420 29390 5505
rect 29510 5420 29740 5505
rect 29860 5420 30090 5505
rect 30210 5420 30440 5505
rect 30560 5420 30790 5505
rect 30910 5420 31140 5505
rect 31260 5420 31490 5505
rect 31610 5420 31840 5505
rect 27410 5370 31840 5420
rect 27410 5275 27640 5370
rect 27760 5275 27990 5370
rect 28110 5275 28340 5370
rect 28460 5275 28690 5370
rect 28810 5275 29040 5370
rect 29160 5275 29390 5370
rect 29510 5275 29740 5370
rect 29860 5275 30090 5370
rect 30210 5275 30440 5370
rect 30560 5275 30790 5370
rect 30910 5275 31140 5370
rect 31260 5275 31490 5370
rect 31610 5275 31840 5370
rect 31960 5420 32190 5505
rect 32310 5420 32540 5505
rect 32660 5420 32890 5505
rect 33010 5420 33240 5505
rect 33360 5420 33590 5505
rect 33710 5420 33940 5505
rect 34060 5420 34290 5505
rect 34410 5420 34640 5505
rect 34760 5420 34990 5505
rect 35110 5420 35340 5505
rect 35460 5420 35690 5505
rect 35810 5420 36040 5505
rect 36160 5420 36390 5505
rect 31960 5370 36390 5420
rect 31960 5275 32190 5370
rect 32310 5275 32540 5370
rect 32660 5275 32890 5370
rect 33010 5275 33240 5370
rect 33360 5275 33590 5370
rect 33710 5275 33940 5370
rect 34060 5275 34290 5370
rect 34410 5275 34640 5370
rect 34760 5275 34990 5370
rect 35110 5275 35340 5370
rect 35460 5275 35690 5370
rect 35810 5275 36040 5370
rect 36160 5275 36390 5370
rect 28200 5155 28250 5275
rect 29250 5155 29300 5275
rect 29600 5155 29650 5275
rect 29950 5155 30000 5275
rect 30300 5155 30350 5275
rect 33450 5155 33500 5275
rect 33800 5155 33850 5275
rect 34150 5155 34200 5275
rect 34500 5155 34550 5275
rect 35550 5155 35600 5275
rect 27410 5070 27640 5155
rect 27760 5070 27990 5155
rect 28110 5070 28340 5155
rect 28460 5070 28690 5155
rect 28810 5070 29040 5155
rect 27410 5020 29040 5070
rect 27410 4925 27640 5020
rect 27760 4925 27990 5020
rect 28110 4925 28340 5020
rect 28460 4925 28690 5020
rect 28810 4925 29040 5020
rect 29160 4925 29390 5155
rect 29510 4925 29740 5155
rect 29860 4925 30090 5155
rect 30210 4925 30440 5155
rect 33360 4925 33590 5155
rect 33710 4925 33940 5155
rect 34060 4925 34290 5155
rect 34410 4925 34640 5155
rect 34760 5070 34990 5155
rect 35110 5070 35340 5155
rect 35460 5070 35690 5155
rect 35810 5070 36040 5155
rect 36160 5070 36390 5155
rect 34760 5020 36390 5070
rect 34760 4925 34990 5020
rect 35110 4925 35340 5020
rect 35460 4925 35690 5020
rect 35810 4925 36040 5020
rect 36160 4925 36390 5020
rect 28200 4805 28250 4925
rect 29250 4805 29300 4925
rect 29600 4805 29650 4925
rect 29950 4805 30000 4925
rect 30300 4805 30350 4925
rect 33450 4805 33500 4925
rect 33800 4805 33850 4925
rect 34150 4805 34200 4925
rect 34500 4805 34550 4925
rect 35550 4805 35600 4925
rect 27410 4720 27640 4805
rect 27760 4720 27990 4805
rect 28110 4720 28340 4805
rect 28460 4720 28690 4805
rect 28810 4720 29040 4805
rect 27410 4670 29040 4720
rect 27410 4575 27640 4670
rect 27760 4575 27990 4670
rect 28110 4575 28340 4670
rect 28460 4575 28690 4670
rect 28810 4575 29040 4670
rect 29160 4575 29390 4805
rect 29510 4575 29740 4805
rect 29860 4575 30090 4805
rect 30210 4575 30440 4805
rect 33360 4575 33590 4805
rect 33710 4575 33940 4805
rect 34060 4575 34290 4805
rect 34410 4575 34640 4805
rect 34760 4720 34990 4805
rect 35110 4720 35340 4805
rect 35460 4720 35690 4805
rect 35810 4720 36040 4805
rect 36160 4720 36390 4805
rect 34760 4670 36390 4720
rect 34760 4575 34990 4670
rect 35110 4575 35340 4670
rect 35460 4575 35690 4670
rect 35810 4575 36040 4670
rect 36160 4575 36390 4670
rect 28200 4455 28250 4575
rect 29250 4455 29300 4575
rect 29600 4455 29650 4575
rect 29950 4455 30000 4575
rect 30300 4455 30350 4575
rect 33450 4455 33500 4575
rect 33800 4455 33850 4575
rect 34150 4455 34200 4575
rect 34500 4455 34550 4575
rect 35550 4455 35600 4575
rect 27410 4370 27640 4455
rect 27760 4370 27990 4455
rect 28110 4370 28340 4455
rect 28460 4370 28690 4455
rect 28810 4370 29040 4455
rect 27410 4320 29040 4370
rect 27410 4225 27640 4320
rect 27760 4225 27990 4320
rect 28110 4225 28340 4320
rect 28460 4225 28690 4320
rect 28810 4225 29040 4320
rect 29160 4225 29390 4455
rect 29510 4225 29740 4455
rect 29860 4225 30090 4455
rect 30210 4225 30440 4455
rect 33360 4225 33590 4455
rect 33710 4225 33940 4455
rect 34060 4225 34290 4455
rect 34410 4225 34640 4455
rect 34760 4370 34990 4455
rect 35110 4370 35340 4455
rect 35460 4370 35690 4455
rect 35810 4370 36040 4455
rect 36160 4370 36390 4455
rect 34760 4320 36390 4370
rect 34760 4225 34990 4320
rect 35110 4225 35340 4320
rect 35460 4225 35690 4320
rect 35810 4225 36040 4320
rect 36160 4225 36390 4320
rect 28200 4105 28250 4225
rect 29250 4105 29300 4225
rect 29600 4105 29650 4225
rect 29950 4105 30000 4225
rect 30300 4105 30350 4225
rect 33450 4105 33500 4225
rect 33800 4105 33850 4225
rect 34150 4105 34200 4225
rect 34500 4105 34550 4225
rect 35550 4105 35600 4225
rect 27410 4020 27640 4105
rect 27760 4020 27990 4105
rect 28110 4020 28340 4105
rect 28460 4020 28690 4105
rect 28810 4020 29040 4105
rect 27410 3970 29040 4020
rect 27410 3875 27640 3970
rect 27760 3875 27990 3970
rect 28110 3875 28340 3970
rect 28460 3875 28690 3970
rect 28810 3875 29040 3970
rect 29160 3875 29390 4105
rect 29510 3875 29740 4105
rect 29860 3875 30090 4105
rect 30210 3875 30440 4105
rect 33360 3875 33590 4105
rect 33710 3875 33940 4105
rect 34060 3875 34290 4105
rect 34410 3875 34640 4105
rect 34760 4020 34990 4105
rect 35110 4020 35340 4105
rect 35460 4020 35690 4105
rect 35810 4020 36040 4105
rect 36160 4020 36390 4105
rect 34760 3970 36390 4020
rect 34760 3875 34990 3970
rect 35110 3875 35340 3970
rect 35460 3875 35690 3970
rect 35810 3875 36040 3970
rect 36160 3875 36390 3970
rect 28200 3755 28250 3875
rect 27410 3670 27640 3755
rect 27760 3670 27990 3755
rect 28110 3670 28340 3755
rect 28460 3670 28690 3755
rect 28810 3670 29040 3755
rect 29605 3735 29645 3875
rect 29605 3705 29610 3735
rect 29640 3705 29645 3735
rect 29605 3700 29645 3705
rect 34155 3735 34195 3875
rect 35550 3755 35600 3875
rect 34155 3705 34160 3735
rect 34190 3705 34195 3735
rect 34155 3700 34195 3705
rect 27410 3620 29040 3670
rect 27410 3525 27640 3620
rect 27760 3525 27990 3620
rect 28110 3525 28340 3620
rect 28460 3525 28690 3620
rect 28810 3525 29040 3620
rect 34760 3670 34990 3755
rect 35110 3670 35340 3755
rect 35460 3670 35690 3755
rect 35810 3670 36040 3755
rect 36160 3670 36390 3755
rect 34760 3620 36390 3670
rect 34760 3525 34990 3620
rect 35110 3525 35340 3620
rect 35460 3525 35690 3620
rect 35810 3525 36040 3620
rect 36160 3525 36390 3620
rect 28200 3405 28250 3525
rect 35550 3405 35600 3525
rect 27410 3320 27640 3405
rect 27760 3320 27990 3405
rect 28110 3320 28340 3405
rect 28460 3320 28690 3405
rect 28810 3320 29040 3405
rect 27410 3270 29040 3320
rect 27410 3175 27640 3270
rect 27760 3175 27990 3270
rect 28110 3175 28340 3270
rect 28460 3175 28690 3270
rect 28810 3175 29040 3270
rect 34760 3320 34990 3405
rect 35110 3320 35340 3405
rect 35460 3320 35690 3405
rect 35810 3320 36040 3405
rect 36160 3320 36390 3405
rect 34760 3270 36390 3320
rect 34760 3175 34990 3270
rect 35110 3175 35340 3270
rect 35460 3175 35690 3270
rect 35810 3175 36040 3270
rect 36160 3175 36390 3270
rect 28200 3055 28250 3175
rect 35550 3055 35600 3175
rect 27410 2970 27640 3055
rect 27760 2970 27990 3055
rect 28110 2970 28340 3055
rect 28460 2970 28690 3055
rect 28810 2970 29040 3055
rect 27410 2920 29040 2970
rect 27410 2825 27640 2920
rect 27760 2825 27990 2920
rect 28110 2825 28340 2920
rect 28460 2825 28690 2920
rect 28810 2825 29040 2920
rect 34760 2970 34990 3055
rect 35110 2970 35340 3055
rect 35460 2970 35690 3055
rect 35810 2970 36040 3055
rect 36160 2970 36390 3055
rect 34760 2920 36390 2970
rect 34760 2825 34990 2920
rect 35110 2825 35340 2920
rect 35460 2825 35690 2920
rect 35810 2825 36040 2920
rect 36160 2825 36390 2920
rect 28200 2705 28250 2825
rect 35550 2705 35600 2825
rect 27410 2620 27640 2705
rect 27760 2620 27990 2705
rect 28110 2620 28340 2705
rect 28460 2620 28690 2705
rect 28810 2620 29040 2705
rect 27410 2570 29040 2620
rect 27410 2475 27640 2570
rect 27760 2475 27990 2570
rect 28110 2475 28340 2570
rect 28460 2475 28690 2570
rect 28810 2475 29040 2570
rect 34760 2620 34990 2705
rect 35110 2620 35340 2705
rect 35460 2620 35690 2705
rect 35810 2620 36040 2705
rect 36160 2620 36390 2705
rect 34760 2570 36390 2620
rect 34760 2475 34990 2570
rect 35110 2475 35340 2570
rect 35460 2475 35690 2570
rect 35810 2475 36040 2570
rect 36160 2475 36390 2570
rect 28200 2355 28250 2475
rect 35550 2355 35600 2475
rect 27410 2270 27640 2355
rect 27760 2270 27990 2355
rect 28110 2270 28340 2355
rect 28460 2270 28690 2355
rect 28810 2270 29040 2355
rect 34760 2270 34990 2355
rect 35110 2270 35340 2355
rect 35460 2270 35690 2355
rect 35810 2270 36040 2355
rect 36160 2270 36390 2355
rect 27410 2220 29040 2270
rect 29310 2265 29360 2270
rect 29310 2225 29315 2265
rect 29355 2225 29360 2265
rect 29310 2220 29360 2225
rect 34440 2265 34490 2270
rect 34440 2225 34445 2265
rect 34485 2225 34490 2265
rect 34440 2220 34490 2225
rect 34760 2220 36390 2270
rect 27410 2125 27640 2220
rect 27760 2125 27990 2220
rect 28110 2125 28340 2220
rect 28460 2125 28690 2220
rect 28810 2125 29040 2220
rect 34760 2125 34990 2220
rect 35110 2125 35340 2220
rect 35460 2125 35690 2220
rect 35810 2125 36040 2220
rect 36160 2125 36390 2220
rect 28200 2005 28250 2125
rect 35550 2005 35600 2125
rect 27410 1920 27640 2005
rect 27760 1920 27990 2005
rect 28110 1920 28340 2005
rect 28460 1920 28690 2005
rect 28810 1920 29040 2005
rect 27410 1870 29040 1920
rect 27410 1775 27640 1870
rect 27760 1775 27990 1870
rect 28110 1775 28340 1870
rect 28460 1775 28690 1870
rect 28810 1775 29040 1870
rect 34760 1920 34990 2005
rect 35110 1920 35340 2005
rect 35460 1920 35690 2005
rect 35810 1920 36040 2005
rect 36160 1920 36390 2005
rect 34760 1870 36390 1920
rect 34760 1775 34990 1870
rect 35110 1775 35340 1870
rect 35460 1775 35690 1870
rect 35810 1775 36040 1870
rect 36160 1775 36390 1870
rect 28200 1655 28250 1775
rect 35550 1655 35600 1775
rect 27410 1570 27640 1655
rect 27760 1570 27990 1655
rect 28110 1570 28340 1655
rect 28460 1570 28690 1655
rect 28810 1570 29040 1655
rect 27410 1520 29040 1570
rect 27410 1425 27640 1520
rect 27760 1425 27990 1520
rect 28110 1425 28340 1520
rect 28460 1425 28690 1520
rect 28810 1425 29040 1520
rect 34760 1570 34990 1655
rect 35110 1570 35340 1655
rect 35460 1570 35690 1655
rect 35810 1570 36040 1655
rect 36160 1570 36390 1655
rect 34760 1520 36390 1570
rect 34760 1425 34990 1520
rect 35110 1425 35340 1520
rect 35460 1425 35690 1520
rect 35810 1425 36040 1520
rect 36160 1425 36390 1520
rect 28200 1305 28250 1425
rect 35550 1305 35600 1425
rect 27410 1220 27640 1305
rect 27760 1220 27990 1305
rect 28110 1220 28340 1305
rect 28460 1220 28690 1305
rect 28810 1220 29040 1305
rect 27410 1170 29040 1220
rect 27410 1075 27640 1170
rect 27760 1075 27990 1170
rect 28110 1075 28340 1170
rect 28460 1075 28690 1170
rect 28810 1075 29040 1170
rect 34760 1220 34990 1305
rect 35110 1220 35340 1305
rect 35460 1220 35690 1305
rect 35810 1220 36040 1305
rect 36160 1220 36390 1305
rect 34760 1170 36390 1220
rect 34760 1075 34990 1170
rect 35110 1075 35340 1170
rect 35460 1075 35690 1170
rect 35810 1075 36040 1170
rect 36160 1075 36390 1170
rect 28200 955 28250 1075
rect 35550 955 35600 1075
rect 27410 870 27640 955
rect 27760 870 27990 955
rect 28110 870 28340 955
rect 28460 870 28690 955
rect 28810 870 29040 955
rect 27410 820 29040 870
rect 27410 725 27640 820
rect 27760 725 27990 820
rect 28110 725 28340 820
rect 28460 725 28690 820
rect 28810 725 29040 820
rect 34760 870 34990 955
rect 35110 870 35340 955
rect 35460 870 35690 955
rect 35810 870 36040 955
rect 36160 870 36390 955
rect 34760 820 36390 870
rect 34760 725 34990 820
rect 35110 725 35340 820
rect 35460 725 35690 820
rect 35810 725 36040 820
rect 36160 725 36390 820
rect 28200 605 28250 725
rect 35550 605 35600 725
rect 27410 520 27640 605
rect 27760 520 27990 605
rect 28110 520 28340 605
rect 28460 520 28690 605
rect 28810 520 29040 605
rect 27410 470 29040 520
rect 27410 375 27640 470
rect 27760 375 27990 470
rect 28110 375 28340 470
rect 28460 375 28690 470
rect 28810 375 29040 470
rect 34760 520 34990 605
rect 35110 520 35340 605
rect 35460 520 35690 605
rect 35810 520 36040 605
rect 36160 520 36390 605
rect 34760 470 36390 520
rect 34760 375 34990 470
rect 35110 375 35340 470
rect 35460 375 35690 470
rect 35810 375 36040 470
rect 36160 375 36390 470
rect 28200 255 28250 375
rect 35550 255 35600 375
rect 27410 170 27640 255
rect 27760 170 27990 255
rect 28110 170 28340 255
rect 28460 170 28690 255
rect 28810 170 29040 255
rect 29160 170 29390 255
rect 29510 170 29740 255
rect 29860 170 30090 255
rect 30210 170 30440 255
rect 30560 170 30790 255
rect 30910 170 31140 255
rect 31260 170 31490 255
rect 31610 170 31840 255
rect 27410 120 31840 170
rect 27410 25 27640 120
rect 27760 25 27990 120
rect 28110 25 28340 120
rect 28460 25 28690 120
rect 28810 25 29040 120
rect 29160 25 29390 120
rect 29510 25 29740 120
rect 29860 25 30090 120
rect 30210 25 30440 120
rect 30560 25 30790 120
rect 30910 25 31140 120
rect 31260 25 31490 120
rect 31610 25 31840 120
rect 31960 170 32190 255
rect 32310 170 32540 255
rect 32660 170 32890 255
rect 33010 170 33240 255
rect 33360 170 33590 255
rect 33710 170 33940 255
rect 34060 170 34290 255
rect 34410 170 34640 255
rect 34760 170 34990 255
rect 35110 170 35340 255
rect 35460 170 35690 255
rect 35810 170 36040 255
rect 36160 170 36390 255
rect 31960 120 36390 170
rect 31960 25 32190 120
rect 32310 25 32540 120
rect 32660 25 32890 120
rect 33010 25 33240 120
rect 33360 25 33590 120
rect 33710 25 33940 120
rect 34060 25 34290 120
rect 34410 25 34640 120
rect 34760 25 34990 120
rect 35110 25 35340 120
rect 35460 25 35690 120
rect 35810 25 36040 120
rect 36160 25 36390 120
rect 28200 -95 28250 25
rect 28550 -95 28600 25
rect 28900 -95 28950 25
rect 29250 -95 29300 25
rect 29600 -95 29650 25
rect 29950 -95 30000 25
rect 30300 -95 30350 25
rect 30650 -95 30700 25
rect 31000 -95 31050 25
rect 31350 -95 31400 25
rect 31700 -95 31750 25
rect 32050 -95 32100 25
rect 32400 -95 32450 25
rect 32750 -95 32800 25
rect 33100 -95 33150 25
rect 33450 -95 33500 25
rect 33800 -95 33850 25
rect 34150 -95 34200 25
rect 34500 -95 34550 25
rect 34850 -95 34900 25
rect 35200 -95 35250 25
rect 35550 -95 35600 25
rect 27410 -180 27640 -95
rect 27760 -180 27990 -95
rect 28110 -180 28340 -95
rect 27410 -230 28340 -180
rect 27410 -325 27640 -230
rect 27760 -325 27990 -230
rect 28110 -325 28340 -230
rect 28460 -325 28690 -95
rect 28810 -325 29040 -95
rect 29160 -325 29390 -95
rect 29510 -325 29740 -95
rect 29860 -325 30090 -95
rect 30210 -325 30440 -95
rect 30560 -325 30790 -95
rect 30910 -325 31140 -95
rect 31260 -325 31490 -95
rect 31610 -325 31840 -95
rect 31960 -325 32190 -95
rect 32310 -325 32540 -95
rect 32660 -325 32890 -95
rect 33010 -325 33240 -95
rect 33360 -325 33590 -95
rect 33710 -325 33940 -95
rect 34060 -325 34290 -95
rect 34410 -325 34640 -95
rect 34760 -325 34990 -95
rect 35110 -325 35340 -95
rect 35460 -180 35690 -95
rect 35810 -180 36040 -95
rect 36160 -180 36390 -95
rect 35460 -230 36390 -180
rect 35460 -325 35690 -230
rect 35810 -325 36040 -230
rect 36160 -325 36390 -230
rect 30780 -510 30830 -505
rect 30780 -550 30785 -510
rect 30825 -550 30830 -510
rect 30780 -555 30830 -550
<< via3 >>
rect 30785 6185 30825 6190
rect 30785 6155 30790 6185
rect 30790 6155 30820 6185
rect 30820 6155 30825 6185
rect 30785 6150 30825 6155
rect 29315 2260 29355 2265
rect 29315 2230 29320 2260
rect 29320 2230 29350 2260
rect 29350 2230 29355 2260
rect 29315 2225 29355 2230
rect 34445 2260 34485 2265
rect 34445 2230 34450 2260
rect 34450 2230 34480 2260
rect 34480 2230 34485 2260
rect 34445 2225 34485 2230
rect 30785 -515 30825 -510
rect 30785 -545 30790 -515
rect 30790 -545 30820 -515
rect 30820 -545 30825 -515
rect 30785 -550 30825 -545
<< mimcap >>
rect 27425 5765 27625 5840
rect 27425 5725 27505 5765
rect 27545 5725 27625 5765
rect 27425 5640 27625 5725
rect 27775 5765 27975 5840
rect 27775 5725 27855 5765
rect 27895 5725 27975 5765
rect 27775 5640 27975 5725
rect 28125 5765 28325 5840
rect 28125 5725 28205 5765
rect 28245 5725 28325 5765
rect 28125 5640 28325 5725
rect 28475 5765 28675 5840
rect 28475 5725 28555 5765
rect 28595 5725 28675 5765
rect 28475 5640 28675 5725
rect 28825 5765 29025 5840
rect 28825 5725 28905 5765
rect 28945 5725 29025 5765
rect 28825 5640 29025 5725
rect 29175 5765 29375 5840
rect 29175 5725 29255 5765
rect 29295 5725 29375 5765
rect 29175 5640 29375 5725
rect 29525 5765 29725 5840
rect 29525 5725 29605 5765
rect 29645 5725 29725 5765
rect 29525 5640 29725 5725
rect 29875 5765 30075 5840
rect 29875 5725 29955 5765
rect 29995 5725 30075 5765
rect 29875 5640 30075 5725
rect 30225 5765 30425 5840
rect 30225 5725 30305 5765
rect 30345 5725 30425 5765
rect 30225 5640 30425 5725
rect 30575 5765 30775 5840
rect 30575 5725 30655 5765
rect 30695 5725 30775 5765
rect 30575 5640 30775 5725
rect 30925 5765 31125 5840
rect 30925 5725 31005 5765
rect 31045 5725 31125 5765
rect 30925 5640 31125 5725
rect 31275 5765 31475 5840
rect 31275 5725 31355 5765
rect 31395 5725 31475 5765
rect 31275 5640 31475 5725
rect 31625 5765 31825 5840
rect 31625 5725 31705 5765
rect 31745 5725 31825 5765
rect 31625 5640 31825 5725
rect 31975 5765 32175 5840
rect 31975 5725 32055 5765
rect 32095 5725 32175 5765
rect 31975 5640 32175 5725
rect 32325 5765 32525 5840
rect 32325 5725 32405 5765
rect 32445 5725 32525 5765
rect 32325 5640 32525 5725
rect 32675 5765 32875 5840
rect 32675 5725 32755 5765
rect 32795 5725 32875 5765
rect 32675 5640 32875 5725
rect 33025 5765 33225 5840
rect 33025 5725 33105 5765
rect 33145 5725 33225 5765
rect 33025 5640 33225 5725
rect 33375 5765 33575 5840
rect 33375 5725 33455 5765
rect 33495 5725 33575 5765
rect 33375 5640 33575 5725
rect 33725 5765 33925 5840
rect 33725 5725 33805 5765
rect 33845 5725 33925 5765
rect 33725 5640 33925 5725
rect 34075 5765 34275 5840
rect 34075 5725 34155 5765
rect 34195 5725 34275 5765
rect 34075 5640 34275 5725
rect 34425 5765 34625 5840
rect 34425 5725 34505 5765
rect 34545 5725 34625 5765
rect 34425 5640 34625 5725
rect 34775 5765 34975 5840
rect 34775 5725 34855 5765
rect 34895 5725 34975 5765
rect 34775 5640 34975 5725
rect 35125 5765 35325 5840
rect 35125 5725 35205 5765
rect 35245 5725 35325 5765
rect 35125 5640 35325 5725
rect 35475 5765 35675 5840
rect 35475 5725 35555 5765
rect 35595 5725 35675 5765
rect 35475 5640 35675 5725
rect 35825 5765 36025 5840
rect 35825 5725 35905 5765
rect 35945 5725 36025 5765
rect 35825 5640 36025 5725
rect 36175 5765 36375 5840
rect 36175 5725 36255 5765
rect 36295 5725 36375 5765
rect 36175 5640 36375 5725
rect 27425 5415 27625 5490
rect 27425 5375 27505 5415
rect 27545 5375 27625 5415
rect 27425 5290 27625 5375
rect 27775 5415 27975 5490
rect 27775 5375 27855 5415
rect 27895 5375 27975 5415
rect 27775 5290 27975 5375
rect 28125 5415 28325 5490
rect 28125 5375 28205 5415
rect 28245 5375 28325 5415
rect 28125 5290 28325 5375
rect 28475 5415 28675 5490
rect 28475 5375 28555 5415
rect 28595 5375 28675 5415
rect 28475 5290 28675 5375
rect 28825 5415 29025 5490
rect 28825 5375 28905 5415
rect 28945 5375 29025 5415
rect 28825 5290 29025 5375
rect 29175 5415 29375 5490
rect 29175 5375 29255 5415
rect 29295 5375 29375 5415
rect 29175 5290 29375 5375
rect 29525 5415 29725 5490
rect 29525 5375 29605 5415
rect 29645 5375 29725 5415
rect 29525 5290 29725 5375
rect 29875 5415 30075 5490
rect 29875 5375 29955 5415
rect 29995 5375 30075 5415
rect 29875 5290 30075 5375
rect 30225 5415 30425 5490
rect 30225 5375 30305 5415
rect 30345 5375 30425 5415
rect 30225 5290 30425 5375
rect 30575 5415 30775 5490
rect 30575 5375 30655 5415
rect 30695 5375 30775 5415
rect 30575 5290 30775 5375
rect 30925 5415 31125 5490
rect 30925 5375 31005 5415
rect 31045 5375 31125 5415
rect 30925 5290 31125 5375
rect 31275 5415 31475 5490
rect 31275 5375 31355 5415
rect 31395 5375 31475 5415
rect 31275 5290 31475 5375
rect 31625 5415 31825 5490
rect 31625 5375 31705 5415
rect 31745 5375 31825 5415
rect 31625 5290 31825 5375
rect 31975 5415 32175 5490
rect 31975 5375 32055 5415
rect 32095 5375 32175 5415
rect 31975 5290 32175 5375
rect 32325 5415 32525 5490
rect 32325 5375 32405 5415
rect 32445 5375 32525 5415
rect 32325 5290 32525 5375
rect 32675 5415 32875 5490
rect 32675 5375 32755 5415
rect 32795 5375 32875 5415
rect 32675 5290 32875 5375
rect 33025 5415 33225 5490
rect 33025 5375 33105 5415
rect 33145 5375 33225 5415
rect 33025 5290 33225 5375
rect 33375 5415 33575 5490
rect 33375 5375 33455 5415
rect 33495 5375 33575 5415
rect 33375 5290 33575 5375
rect 33725 5415 33925 5490
rect 33725 5375 33805 5415
rect 33845 5375 33925 5415
rect 33725 5290 33925 5375
rect 34075 5415 34275 5490
rect 34075 5375 34155 5415
rect 34195 5375 34275 5415
rect 34075 5290 34275 5375
rect 34425 5415 34625 5490
rect 34425 5375 34505 5415
rect 34545 5375 34625 5415
rect 34425 5290 34625 5375
rect 34775 5415 34975 5490
rect 34775 5375 34855 5415
rect 34895 5375 34975 5415
rect 34775 5290 34975 5375
rect 35125 5415 35325 5490
rect 35125 5375 35205 5415
rect 35245 5375 35325 5415
rect 35125 5290 35325 5375
rect 35475 5415 35675 5490
rect 35475 5375 35555 5415
rect 35595 5375 35675 5415
rect 35475 5290 35675 5375
rect 35825 5415 36025 5490
rect 35825 5375 35905 5415
rect 35945 5375 36025 5415
rect 35825 5290 36025 5375
rect 36175 5415 36375 5490
rect 36175 5375 36255 5415
rect 36295 5375 36375 5415
rect 36175 5290 36375 5375
rect 27425 5065 27625 5140
rect 27425 5025 27505 5065
rect 27545 5025 27625 5065
rect 27425 4940 27625 5025
rect 27775 5065 27975 5140
rect 27775 5025 27855 5065
rect 27895 5025 27975 5065
rect 27775 4940 27975 5025
rect 28125 5065 28325 5140
rect 28125 5025 28205 5065
rect 28245 5025 28325 5065
rect 28125 4940 28325 5025
rect 28475 5065 28675 5140
rect 28475 5025 28555 5065
rect 28595 5025 28675 5065
rect 28475 4940 28675 5025
rect 28825 5065 29025 5140
rect 28825 5025 28905 5065
rect 28945 5025 29025 5065
rect 28825 4940 29025 5025
rect 29175 5065 29375 5140
rect 29175 5025 29255 5065
rect 29295 5025 29375 5065
rect 29175 4940 29375 5025
rect 29525 5065 29725 5140
rect 29525 5025 29605 5065
rect 29645 5025 29725 5065
rect 29525 4940 29725 5025
rect 29875 5065 30075 5140
rect 29875 5025 29955 5065
rect 29995 5025 30075 5065
rect 29875 4940 30075 5025
rect 30225 5065 30425 5140
rect 30225 5025 30305 5065
rect 30345 5025 30425 5065
rect 30225 4940 30425 5025
rect 33375 5065 33575 5140
rect 33375 5025 33455 5065
rect 33495 5025 33575 5065
rect 33375 4940 33575 5025
rect 33725 5065 33925 5140
rect 33725 5025 33805 5065
rect 33845 5025 33925 5065
rect 33725 4940 33925 5025
rect 34075 5065 34275 5140
rect 34075 5025 34155 5065
rect 34195 5025 34275 5065
rect 34075 4940 34275 5025
rect 34425 5065 34625 5140
rect 34425 5025 34505 5065
rect 34545 5025 34625 5065
rect 34425 4940 34625 5025
rect 34775 5065 34975 5140
rect 34775 5025 34855 5065
rect 34895 5025 34975 5065
rect 34775 4940 34975 5025
rect 35125 5065 35325 5140
rect 35125 5025 35205 5065
rect 35245 5025 35325 5065
rect 35125 4940 35325 5025
rect 35475 5065 35675 5140
rect 35475 5025 35555 5065
rect 35595 5025 35675 5065
rect 35475 4940 35675 5025
rect 35825 5065 36025 5140
rect 35825 5025 35905 5065
rect 35945 5025 36025 5065
rect 35825 4940 36025 5025
rect 36175 5065 36375 5140
rect 36175 5025 36255 5065
rect 36295 5025 36375 5065
rect 36175 4940 36375 5025
rect 27425 4715 27625 4790
rect 27425 4675 27505 4715
rect 27545 4675 27625 4715
rect 27425 4590 27625 4675
rect 27775 4715 27975 4790
rect 27775 4675 27855 4715
rect 27895 4675 27975 4715
rect 27775 4590 27975 4675
rect 28125 4715 28325 4790
rect 28125 4675 28205 4715
rect 28245 4675 28325 4715
rect 28125 4590 28325 4675
rect 28475 4715 28675 4790
rect 28475 4675 28555 4715
rect 28595 4675 28675 4715
rect 28475 4590 28675 4675
rect 28825 4715 29025 4790
rect 28825 4675 28905 4715
rect 28945 4675 29025 4715
rect 28825 4590 29025 4675
rect 29175 4715 29375 4790
rect 29175 4675 29255 4715
rect 29295 4675 29375 4715
rect 29175 4590 29375 4675
rect 29525 4715 29725 4790
rect 29525 4675 29605 4715
rect 29645 4675 29725 4715
rect 29525 4590 29725 4675
rect 29875 4715 30075 4790
rect 29875 4675 29955 4715
rect 29995 4675 30075 4715
rect 29875 4590 30075 4675
rect 30225 4715 30425 4790
rect 30225 4675 30305 4715
rect 30345 4675 30425 4715
rect 30225 4590 30425 4675
rect 33375 4715 33575 4790
rect 33375 4675 33455 4715
rect 33495 4675 33575 4715
rect 33375 4590 33575 4675
rect 33725 4715 33925 4790
rect 33725 4675 33805 4715
rect 33845 4675 33925 4715
rect 33725 4590 33925 4675
rect 34075 4715 34275 4790
rect 34075 4675 34155 4715
rect 34195 4675 34275 4715
rect 34075 4590 34275 4675
rect 34425 4715 34625 4790
rect 34425 4675 34505 4715
rect 34545 4675 34625 4715
rect 34425 4590 34625 4675
rect 34775 4715 34975 4790
rect 34775 4675 34855 4715
rect 34895 4675 34975 4715
rect 34775 4590 34975 4675
rect 35125 4715 35325 4790
rect 35125 4675 35205 4715
rect 35245 4675 35325 4715
rect 35125 4590 35325 4675
rect 35475 4715 35675 4790
rect 35475 4675 35555 4715
rect 35595 4675 35675 4715
rect 35475 4590 35675 4675
rect 35825 4715 36025 4790
rect 35825 4675 35905 4715
rect 35945 4675 36025 4715
rect 35825 4590 36025 4675
rect 36175 4715 36375 4790
rect 36175 4675 36255 4715
rect 36295 4675 36375 4715
rect 36175 4590 36375 4675
rect 27425 4365 27625 4440
rect 27425 4325 27505 4365
rect 27545 4325 27625 4365
rect 27425 4240 27625 4325
rect 27775 4365 27975 4440
rect 27775 4325 27855 4365
rect 27895 4325 27975 4365
rect 27775 4240 27975 4325
rect 28125 4365 28325 4440
rect 28125 4325 28205 4365
rect 28245 4325 28325 4365
rect 28125 4240 28325 4325
rect 28475 4365 28675 4440
rect 28475 4325 28555 4365
rect 28595 4325 28675 4365
rect 28475 4240 28675 4325
rect 28825 4365 29025 4440
rect 28825 4325 28905 4365
rect 28945 4325 29025 4365
rect 28825 4240 29025 4325
rect 29175 4365 29375 4440
rect 29175 4325 29255 4365
rect 29295 4325 29375 4365
rect 29175 4240 29375 4325
rect 29525 4365 29725 4440
rect 29525 4325 29605 4365
rect 29645 4325 29725 4365
rect 29525 4240 29725 4325
rect 29875 4365 30075 4440
rect 29875 4325 29955 4365
rect 29995 4325 30075 4365
rect 29875 4240 30075 4325
rect 30225 4365 30425 4440
rect 30225 4325 30305 4365
rect 30345 4325 30425 4365
rect 30225 4240 30425 4325
rect 33375 4365 33575 4440
rect 33375 4325 33455 4365
rect 33495 4325 33575 4365
rect 33375 4240 33575 4325
rect 33725 4365 33925 4440
rect 33725 4325 33805 4365
rect 33845 4325 33925 4365
rect 33725 4240 33925 4325
rect 34075 4365 34275 4440
rect 34075 4325 34155 4365
rect 34195 4325 34275 4365
rect 34075 4240 34275 4325
rect 34425 4365 34625 4440
rect 34425 4325 34505 4365
rect 34545 4325 34625 4365
rect 34425 4240 34625 4325
rect 34775 4365 34975 4440
rect 34775 4325 34855 4365
rect 34895 4325 34975 4365
rect 34775 4240 34975 4325
rect 35125 4365 35325 4440
rect 35125 4325 35205 4365
rect 35245 4325 35325 4365
rect 35125 4240 35325 4325
rect 35475 4365 35675 4440
rect 35475 4325 35555 4365
rect 35595 4325 35675 4365
rect 35475 4240 35675 4325
rect 35825 4365 36025 4440
rect 35825 4325 35905 4365
rect 35945 4325 36025 4365
rect 35825 4240 36025 4325
rect 36175 4365 36375 4440
rect 36175 4325 36255 4365
rect 36295 4325 36375 4365
rect 36175 4240 36375 4325
rect 27425 4015 27625 4090
rect 27425 3975 27505 4015
rect 27545 3975 27625 4015
rect 27425 3890 27625 3975
rect 27775 4015 27975 4090
rect 27775 3975 27855 4015
rect 27895 3975 27975 4015
rect 27775 3890 27975 3975
rect 28125 4015 28325 4090
rect 28125 3975 28205 4015
rect 28245 3975 28325 4015
rect 28125 3890 28325 3975
rect 28475 4015 28675 4090
rect 28475 3975 28555 4015
rect 28595 3975 28675 4015
rect 28475 3890 28675 3975
rect 28825 4015 29025 4090
rect 28825 3975 28905 4015
rect 28945 3975 29025 4015
rect 28825 3890 29025 3975
rect 29175 4015 29375 4090
rect 29175 3975 29255 4015
rect 29295 3975 29375 4015
rect 29175 3890 29375 3975
rect 29525 4015 29725 4090
rect 29525 3975 29605 4015
rect 29645 3975 29725 4015
rect 29525 3890 29725 3975
rect 29875 4015 30075 4090
rect 29875 3975 29955 4015
rect 29995 3975 30075 4015
rect 29875 3890 30075 3975
rect 30225 4015 30425 4090
rect 30225 3975 30305 4015
rect 30345 3975 30425 4015
rect 30225 3890 30425 3975
rect 33375 4015 33575 4090
rect 33375 3975 33455 4015
rect 33495 3975 33575 4015
rect 33375 3890 33575 3975
rect 33725 4015 33925 4090
rect 33725 3975 33805 4015
rect 33845 3975 33925 4015
rect 33725 3890 33925 3975
rect 34075 4015 34275 4090
rect 34075 3975 34155 4015
rect 34195 3975 34275 4015
rect 34075 3890 34275 3975
rect 34425 4015 34625 4090
rect 34425 3975 34505 4015
rect 34545 3975 34625 4015
rect 34425 3890 34625 3975
rect 34775 4015 34975 4090
rect 34775 3975 34855 4015
rect 34895 3975 34975 4015
rect 34775 3890 34975 3975
rect 35125 4015 35325 4090
rect 35125 3975 35205 4015
rect 35245 3975 35325 4015
rect 35125 3890 35325 3975
rect 35475 4015 35675 4090
rect 35475 3975 35555 4015
rect 35595 3975 35675 4015
rect 35475 3890 35675 3975
rect 35825 4015 36025 4090
rect 35825 3975 35905 4015
rect 35945 3975 36025 4015
rect 35825 3890 36025 3975
rect 36175 4015 36375 4090
rect 36175 3975 36255 4015
rect 36295 3975 36375 4015
rect 36175 3890 36375 3975
rect 27425 3665 27625 3740
rect 27425 3625 27505 3665
rect 27545 3625 27625 3665
rect 27425 3540 27625 3625
rect 27775 3665 27975 3740
rect 27775 3625 27855 3665
rect 27895 3625 27975 3665
rect 27775 3540 27975 3625
rect 28125 3665 28325 3740
rect 28125 3625 28205 3665
rect 28245 3625 28325 3665
rect 28125 3540 28325 3625
rect 28475 3665 28675 3740
rect 28475 3625 28555 3665
rect 28595 3625 28675 3665
rect 28475 3540 28675 3625
rect 28825 3665 29025 3740
rect 28825 3625 28905 3665
rect 28945 3625 29025 3665
rect 28825 3540 29025 3625
rect 34775 3665 34975 3740
rect 34775 3625 34855 3665
rect 34895 3625 34975 3665
rect 34775 3540 34975 3625
rect 35125 3665 35325 3740
rect 35125 3625 35205 3665
rect 35245 3625 35325 3665
rect 35125 3540 35325 3625
rect 35475 3665 35675 3740
rect 35475 3625 35555 3665
rect 35595 3625 35675 3665
rect 35475 3540 35675 3625
rect 35825 3665 36025 3740
rect 35825 3625 35905 3665
rect 35945 3625 36025 3665
rect 35825 3540 36025 3625
rect 36175 3665 36375 3740
rect 36175 3625 36255 3665
rect 36295 3625 36375 3665
rect 36175 3540 36375 3625
rect 27425 3315 27625 3390
rect 27425 3275 27505 3315
rect 27545 3275 27625 3315
rect 27425 3190 27625 3275
rect 27775 3315 27975 3390
rect 27775 3275 27855 3315
rect 27895 3275 27975 3315
rect 27775 3190 27975 3275
rect 28125 3315 28325 3390
rect 28125 3275 28205 3315
rect 28245 3275 28325 3315
rect 28125 3190 28325 3275
rect 28475 3315 28675 3390
rect 28475 3275 28555 3315
rect 28595 3275 28675 3315
rect 28475 3190 28675 3275
rect 28825 3315 29025 3390
rect 28825 3275 28905 3315
rect 28945 3275 29025 3315
rect 28825 3190 29025 3275
rect 34775 3315 34975 3390
rect 34775 3275 34855 3315
rect 34895 3275 34975 3315
rect 34775 3190 34975 3275
rect 35125 3315 35325 3390
rect 35125 3275 35205 3315
rect 35245 3275 35325 3315
rect 35125 3190 35325 3275
rect 35475 3315 35675 3390
rect 35475 3275 35555 3315
rect 35595 3275 35675 3315
rect 35475 3190 35675 3275
rect 35825 3315 36025 3390
rect 35825 3275 35905 3315
rect 35945 3275 36025 3315
rect 35825 3190 36025 3275
rect 36175 3315 36375 3390
rect 36175 3275 36255 3315
rect 36295 3275 36375 3315
rect 36175 3190 36375 3275
rect 27425 2965 27625 3040
rect 27425 2925 27505 2965
rect 27545 2925 27625 2965
rect 27425 2840 27625 2925
rect 27775 2965 27975 3040
rect 27775 2925 27855 2965
rect 27895 2925 27975 2965
rect 27775 2840 27975 2925
rect 28125 2965 28325 3040
rect 28125 2925 28205 2965
rect 28245 2925 28325 2965
rect 28125 2840 28325 2925
rect 28475 2965 28675 3040
rect 28475 2925 28555 2965
rect 28595 2925 28675 2965
rect 28475 2840 28675 2925
rect 28825 2965 29025 3040
rect 28825 2925 28905 2965
rect 28945 2925 29025 2965
rect 28825 2840 29025 2925
rect 34775 2965 34975 3040
rect 34775 2925 34855 2965
rect 34895 2925 34975 2965
rect 34775 2840 34975 2925
rect 35125 2965 35325 3040
rect 35125 2925 35205 2965
rect 35245 2925 35325 2965
rect 35125 2840 35325 2925
rect 35475 2965 35675 3040
rect 35475 2925 35555 2965
rect 35595 2925 35675 2965
rect 35475 2840 35675 2925
rect 35825 2965 36025 3040
rect 35825 2925 35905 2965
rect 35945 2925 36025 2965
rect 35825 2840 36025 2925
rect 36175 2965 36375 3040
rect 36175 2925 36255 2965
rect 36295 2925 36375 2965
rect 36175 2840 36375 2925
rect 27425 2615 27625 2690
rect 27425 2575 27505 2615
rect 27545 2575 27625 2615
rect 27425 2490 27625 2575
rect 27775 2615 27975 2690
rect 27775 2575 27855 2615
rect 27895 2575 27975 2615
rect 27775 2490 27975 2575
rect 28125 2615 28325 2690
rect 28125 2575 28205 2615
rect 28245 2575 28325 2615
rect 28125 2490 28325 2575
rect 28475 2615 28675 2690
rect 28475 2575 28555 2615
rect 28595 2575 28675 2615
rect 28475 2490 28675 2575
rect 28825 2615 29025 2690
rect 28825 2575 28905 2615
rect 28945 2575 29025 2615
rect 28825 2490 29025 2575
rect 34775 2615 34975 2690
rect 34775 2575 34855 2615
rect 34895 2575 34975 2615
rect 34775 2490 34975 2575
rect 35125 2615 35325 2690
rect 35125 2575 35205 2615
rect 35245 2575 35325 2615
rect 35125 2490 35325 2575
rect 35475 2615 35675 2690
rect 35475 2575 35555 2615
rect 35595 2575 35675 2615
rect 35475 2490 35675 2575
rect 35825 2615 36025 2690
rect 35825 2575 35905 2615
rect 35945 2575 36025 2615
rect 35825 2490 36025 2575
rect 36175 2615 36375 2690
rect 36175 2575 36255 2615
rect 36295 2575 36375 2615
rect 36175 2490 36375 2575
rect 27425 2265 27625 2340
rect 27425 2225 27505 2265
rect 27545 2225 27625 2265
rect 27425 2140 27625 2225
rect 27775 2265 27975 2340
rect 27775 2225 27855 2265
rect 27895 2225 27975 2265
rect 27775 2140 27975 2225
rect 28125 2265 28325 2340
rect 28125 2225 28205 2265
rect 28245 2225 28325 2265
rect 28125 2140 28325 2225
rect 28475 2265 28675 2340
rect 28475 2225 28555 2265
rect 28595 2225 28675 2265
rect 28475 2140 28675 2225
rect 28825 2265 29025 2340
rect 28825 2225 28905 2265
rect 28945 2225 29025 2265
rect 28825 2140 29025 2225
rect 34775 2265 34975 2340
rect 34775 2225 34855 2265
rect 34895 2225 34975 2265
rect 34775 2140 34975 2225
rect 35125 2265 35325 2340
rect 35125 2225 35205 2265
rect 35245 2225 35325 2265
rect 35125 2140 35325 2225
rect 35475 2265 35675 2340
rect 35475 2225 35555 2265
rect 35595 2225 35675 2265
rect 35475 2140 35675 2225
rect 35825 2265 36025 2340
rect 35825 2225 35905 2265
rect 35945 2225 36025 2265
rect 35825 2140 36025 2225
rect 36175 2265 36375 2340
rect 36175 2225 36255 2265
rect 36295 2225 36375 2265
rect 36175 2140 36375 2225
rect 27425 1915 27625 1990
rect 27425 1875 27505 1915
rect 27545 1875 27625 1915
rect 27425 1790 27625 1875
rect 27775 1915 27975 1990
rect 27775 1875 27855 1915
rect 27895 1875 27975 1915
rect 27775 1790 27975 1875
rect 28125 1915 28325 1990
rect 28125 1875 28205 1915
rect 28245 1875 28325 1915
rect 28125 1790 28325 1875
rect 28475 1915 28675 1990
rect 28475 1875 28555 1915
rect 28595 1875 28675 1915
rect 28475 1790 28675 1875
rect 28825 1915 29025 1990
rect 28825 1875 28905 1915
rect 28945 1875 29025 1915
rect 28825 1790 29025 1875
rect 34775 1915 34975 1990
rect 34775 1875 34855 1915
rect 34895 1875 34975 1915
rect 34775 1790 34975 1875
rect 35125 1915 35325 1990
rect 35125 1875 35205 1915
rect 35245 1875 35325 1915
rect 35125 1790 35325 1875
rect 35475 1915 35675 1990
rect 35475 1875 35555 1915
rect 35595 1875 35675 1915
rect 35475 1790 35675 1875
rect 35825 1915 36025 1990
rect 35825 1875 35905 1915
rect 35945 1875 36025 1915
rect 35825 1790 36025 1875
rect 36175 1915 36375 1990
rect 36175 1875 36255 1915
rect 36295 1875 36375 1915
rect 36175 1790 36375 1875
rect 27425 1565 27625 1640
rect 27425 1525 27505 1565
rect 27545 1525 27625 1565
rect 27425 1440 27625 1525
rect 27775 1565 27975 1640
rect 27775 1525 27855 1565
rect 27895 1525 27975 1565
rect 27775 1440 27975 1525
rect 28125 1565 28325 1640
rect 28125 1525 28205 1565
rect 28245 1525 28325 1565
rect 28125 1440 28325 1525
rect 28475 1565 28675 1640
rect 28475 1525 28555 1565
rect 28595 1525 28675 1565
rect 28475 1440 28675 1525
rect 28825 1565 29025 1640
rect 28825 1525 28905 1565
rect 28945 1525 29025 1565
rect 28825 1440 29025 1525
rect 34775 1565 34975 1640
rect 34775 1525 34855 1565
rect 34895 1525 34975 1565
rect 34775 1440 34975 1525
rect 35125 1565 35325 1640
rect 35125 1525 35205 1565
rect 35245 1525 35325 1565
rect 35125 1440 35325 1525
rect 35475 1565 35675 1640
rect 35475 1525 35555 1565
rect 35595 1525 35675 1565
rect 35475 1440 35675 1525
rect 35825 1565 36025 1640
rect 35825 1525 35905 1565
rect 35945 1525 36025 1565
rect 35825 1440 36025 1525
rect 36175 1565 36375 1640
rect 36175 1525 36255 1565
rect 36295 1525 36375 1565
rect 36175 1440 36375 1525
rect 27425 1215 27625 1290
rect 27425 1175 27505 1215
rect 27545 1175 27625 1215
rect 27425 1090 27625 1175
rect 27775 1215 27975 1290
rect 27775 1175 27855 1215
rect 27895 1175 27975 1215
rect 27775 1090 27975 1175
rect 28125 1215 28325 1290
rect 28125 1175 28205 1215
rect 28245 1175 28325 1215
rect 28125 1090 28325 1175
rect 28475 1215 28675 1290
rect 28475 1175 28555 1215
rect 28595 1175 28675 1215
rect 28475 1090 28675 1175
rect 28825 1215 29025 1290
rect 28825 1175 28905 1215
rect 28945 1175 29025 1215
rect 28825 1090 29025 1175
rect 34775 1215 34975 1290
rect 34775 1175 34855 1215
rect 34895 1175 34975 1215
rect 34775 1090 34975 1175
rect 35125 1215 35325 1290
rect 35125 1175 35205 1215
rect 35245 1175 35325 1215
rect 35125 1090 35325 1175
rect 35475 1215 35675 1290
rect 35475 1175 35555 1215
rect 35595 1175 35675 1215
rect 35475 1090 35675 1175
rect 35825 1215 36025 1290
rect 35825 1175 35905 1215
rect 35945 1175 36025 1215
rect 35825 1090 36025 1175
rect 36175 1215 36375 1290
rect 36175 1175 36255 1215
rect 36295 1175 36375 1215
rect 36175 1090 36375 1175
rect 27425 865 27625 940
rect 27425 825 27505 865
rect 27545 825 27625 865
rect 27425 740 27625 825
rect 27775 865 27975 940
rect 27775 825 27855 865
rect 27895 825 27975 865
rect 27775 740 27975 825
rect 28125 865 28325 940
rect 28125 825 28205 865
rect 28245 825 28325 865
rect 28125 740 28325 825
rect 28475 865 28675 940
rect 28475 825 28555 865
rect 28595 825 28675 865
rect 28475 740 28675 825
rect 28825 865 29025 940
rect 28825 825 28905 865
rect 28945 825 29025 865
rect 28825 740 29025 825
rect 34775 865 34975 940
rect 34775 825 34855 865
rect 34895 825 34975 865
rect 34775 740 34975 825
rect 35125 865 35325 940
rect 35125 825 35205 865
rect 35245 825 35325 865
rect 35125 740 35325 825
rect 35475 865 35675 940
rect 35475 825 35555 865
rect 35595 825 35675 865
rect 35475 740 35675 825
rect 35825 865 36025 940
rect 35825 825 35905 865
rect 35945 825 36025 865
rect 35825 740 36025 825
rect 36175 865 36375 940
rect 36175 825 36255 865
rect 36295 825 36375 865
rect 36175 740 36375 825
rect 27425 515 27625 590
rect 27425 475 27505 515
rect 27545 475 27625 515
rect 27425 390 27625 475
rect 27775 515 27975 590
rect 27775 475 27855 515
rect 27895 475 27975 515
rect 27775 390 27975 475
rect 28125 515 28325 590
rect 28125 475 28205 515
rect 28245 475 28325 515
rect 28125 390 28325 475
rect 28475 515 28675 590
rect 28475 475 28555 515
rect 28595 475 28675 515
rect 28475 390 28675 475
rect 28825 515 29025 590
rect 28825 475 28905 515
rect 28945 475 29025 515
rect 28825 390 29025 475
rect 34775 515 34975 590
rect 34775 475 34855 515
rect 34895 475 34975 515
rect 34775 390 34975 475
rect 35125 515 35325 590
rect 35125 475 35205 515
rect 35245 475 35325 515
rect 35125 390 35325 475
rect 35475 515 35675 590
rect 35475 475 35555 515
rect 35595 475 35675 515
rect 35475 390 35675 475
rect 35825 515 36025 590
rect 35825 475 35905 515
rect 35945 475 36025 515
rect 35825 390 36025 475
rect 36175 515 36375 590
rect 36175 475 36255 515
rect 36295 475 36375 515
rect 36175 390 36375 475
rect 27425 165 27625 240
rect 27425 125 27505 165
rect 27545 125 27625 165
rect 27425 40 27625 125
rect 27775 165 27975 240
rect 27775 125 27855 165
rect 27895 125 27975 165
rect 27775 40 27975 125
rect 28125 165 28325 240
rect 28125 125 28205 165
rect 28245 125 28325 165
rect 28125 40 28325 125
rect 28475 165 28675 240
rect 28475 125 28555 165
rect 28595 125 28675 165
rect 28475 40 28675 125
rect 28825 165 29025 240
rect 28825 125 28905 165
rect 28945 125 29025 165
rect 28825 40 29025 125
rect 29175 165 29375 240
rect 29175 125 29255 165
rect 29295 125 29375 165
rect 29175 40 29375 125
rect 29525 165 29725 240
rect 29525 125 29605 165
rect 29645 125 29725 165
rect 29525 40 29725 125
rect 29875 165 30075 240
rect 29875 125 29955 165
rect 29995 125 30075 165
rect 29875 40 30075 125
rect 30225 165 30425 240
rect 30225 125 30305 165
rect 30345 125 30425 165
rect 30225 40 30425 125
rect 30575 165 30775 240
rect 30575 125 30655 165
rect 30695 125 30775 165
rect 30575 40 30775 125
rect 30925 165 31125 240
rect 30925 125 31005 165
rect 31045 125 31125 165
rect 30925 40 31125 125
rect 31275 165 31475 240
rect 31275 125 31355 165
rect 31395 125 31475 165
rect 31275 40 31475 125
rect 31625 165 31825 240
rect 31625 125 31705 165
rect 31745 125 31825 165
rect 31625 40 31825 125
rect 31975 165 32175 240
rect 31975 125 32055 165
rect 32095 125 32175 165
rect 31975 40 32175 125
rect 32325 165 32525 240
rect 32325 125 32405 165
rect 32445 125 32525 165
rect 32325 40 32525 125
rect 32675 165 32875 240
rect 32675 125 32755 165
rect 32795 125 32875 165
rect 32675 40 32875 125
rect 33025 165 33225 240
rect 33025 125 33105 165
rect 33145 125 33225 165
rect 33025 40 33225 125
rect 33375 165 33575 240
rect 33375 125 33455 165
rect 33495 125 33575 165
rect 33375 40 33575 125
rect 33725 165 33925 240
rect 33725 125 33805 165
rect 33845 125 33925 165
rect 33725 40 33925 125
rect 34075 165 34275 240
rect 34075 125 34155 165
rect 34195 125 34275 165
rect 34075 40 34275 125
rect 34425 165 34625 240
rect 34425 125 34505 165
rect 34545 125 34625 165
rect 34425 40 34625 125
rect 34775 165 34975 240
rect 34775 125 34855 165
rect 34895 125 34975 165
rect 34775 40 34975 125
rect 35125 165 35325 240
rect 35125 125 35205 165
rect 35245 125 35325 165
rect 35125 40 35325 125
rect 35475 165 35675 240
rect 35475 125 35555 165
rect 35595 125 35675 165
rect 35475 40 35675 125
rect 35825 165 36025 240
rect 35825 125 35905 165
rect 35945 125 36025 165
rect 35825 40 36025 125
rect 36175 165 36375 240
rect 36175 125 36255 165
rect 36295 125 36375 165
rect 36175 40 36375 125
rect 27425 -185 27625 -110
rect 27425 -225 27505 -185
rect 27545 -225 27625 -185
rect 27425 -310 27625 -225
rect 27775 -185 27975 -110
rect 27775 -225 27855 -185
rect 27895 -225 27975 -185
rect 27775 -310 27975 -225
rect 28125 -185 28325 -110
rect 28125 -225 28205 -185
rect 28245 -225 28325 -185
rect 28125 -310 28325 -225
rect 28475 -185 28675 -110
rect 28475 -225 28555 -185
rect 28595 -225 28675 -185
rect 28475 -310 28675 -225
rect 28825 -185 29025 -110
rect 28825 -225 28905 -185
rect 28945 -225 29025 -185
rect 28825 -310 29025 -225
rect 29175 -185 29375 -110
rect 29175 -225 29255 -185
rect 29295 -225 29375 -185
rect 29175 -310 29375 -225
rect 29525 -185 29725 -110
rect 29525 -225 29605 -185
rect 29645 -225 29725 -185
rect 29525 -310 29725 -225
rect 29875 -185 30075 -110
rect 29875 -225 29955 -185
rect 29995 -225 30075 -185
rect 29875 -310 30075 -225
rect 30225 -185 30425 -110
rect 30225 -225 30305 -185
rect 30345 -225 30425 -185
rect 30225 -310 30425 -225
rect 30575 -185 30775 -110
rect 30575 -225 30655 -185
rect 30695 -225 30775 -185
rect 30575 -310 30775 -225
rect 30925 -185 31125 -110
rect 30925 -225 31005 -185
rect 31045 -225 31125 -185
rect 30925 -310 31125 -225
rect 31275 -185 31475 -110
rect 31275 -225 31355 -185
rect 31395 -225 31475 -185
rect 31275 -310 31475 -225
rect 31625 -185 31825 -110
rect 31625 -225 31705 -185
rect 31745 -225 31825 -185
rect 31625 -310 31825 -225
rect 31975 -185 32175 -110
rect 31975 -225 32055 -185
rect 32095 -225 32175 -185
rect 31975 -310 32175 -225
rect 32325 -185 32525 -110
rect 32325 -225 32405 -185
rect 32445 -225 32525 -185
rect 32325 -310 32525 -225
rect 32675 -185 32875 -110
rect 32675 -225 32755 -185
rect 32795 -225 32875 -185
rect 32675 -310 32875 -225
rect 33025 -185 33225 -110
rect 33025 -225 33105 -185
rect 33145 -225 33225 -185
rect 33025 -310 33225 -225
rect 33375 -185 33575 -110
rect 33375 -225 33455 -185
rect 33495 -225 33575 -185
rect 33375 -310 33575 -225
rect 33725 -185 33925 -110
rect 33725 -225 33805 -185
rect 33845 -225 33925 -185
rect 33725 -310 33925 -225
rect 34075 -185 34275 -110
rect 34075 -225 34155 -185
rect 34195 -225 34275 -185
rect 34075 -310 34275 -225
rect 34425 -185 34625 -110
rect 34425 -225 34505 -185
rect 34545 -225 34625 -185
rect 34425 -310 34625 -225
rect 34775 -185 34975 -110
rect 34775 -225 34855 -185
rect 34895 -225 34975 -185
rect 34775 -310 34975 -225
rect 35125 -185 35325 -110
rect 35125 -225 35205 -185
rect 35245 -225 35325 -185
rect 35125 -310 35325 -225
rect 35475 -185 35675 -110
rect 35475 -225 35555 -185
rect 35595 -225 35675 -185
rect 35475 -310 35675 -225
rect 35825 -185 36025 -110
rect 35825 -225 35905 -185
rect 35945 -225 36025 -185
rect 35825 -310 36025 -225
rect 36175 -185 36375 -110
rect 36175 -225 36255 -185
rect 36295 -225 36375 -185
rect 36175 -310 36375 -225
<< mimcapcontact >>
rect 27505 5725 27545 5765
rect 27855 5725 27895 5765
rect 28205 5725 28245 5765
rect 28555 5725 28595 5765
rect 28905 5725 28945 5765
rect 29255 5725 29295 5765
rect 29605 5725 29645 5765
rect 29955 5725 29995 5765
rect 30305 5725 30345 5765
rect 30655 5725 30695 5765
rect 31005 5725 31045 5765
rect 31355 5725 31395 5765
rect 31705 5725 31745 5765
rect 32055 5725 32095 5765
rect 32405 5725 32445 5765
rect 32755 5725 32795 5765
rect 33105 5725 33145 5765
rect 33455 5725 33495 5765
rect 33805 5725 33845 5765
rect 34155 5725 34195 5765
rect 34505 5725 34545 5765
rect 34855 5725 34895 5765
rect 35205 5725 35245 5765
rect 35555 5725 35595 5765
rect 35905 5725 35945 5765
rect 36255 5725 36295 5765
rect 27505 5375 27545 5415
rect 27855 5375 27895 5415
rect 28205 5375 28245 5415
rect 28555 5375 28595 5415
rect 28905 5375 28945 5415
rect 29255 5375 29295 5415
rect 29605 5375 29645 5415
rect 29955 5375 29995 5415
rect 30305 5375 30345 5415
rect 30655 5375 30695 5415
rect 31005 5375 31045 5415
rect 31355 5375 31395 5415
rect 31705 5375 31745 5415
rect 32055 5375 32095 5415
rect 32405 5375 32445 5415
rect 32755 5375 32795 5415
rect 33105 5375 33145 5415
rect 33455 5375 33495 5415
rect 33805 5375 33845 5415
rect 34155 5375 34195 5415
rect 34505 5375 34545 5415
rect 34855 5375 34895 5415
rect 35205 5375 35245 5415
rect 35555 5375 35595 5415
rect 35905 5375 35945 5415
rect 36255 5375 36295 5415
rect 27505 5025 27545 5065
rect 27855 5025 27895 5065
rect 28205 5025 28245 5065
rect 28555 5025 28595 5065
rect 28905 5025 28945 5065
rect 29255 5025 29295 5065
rect 29605 5025 29645 5065
rect 29955 5025 29995 5065
rect 30305 5025 30345 5065
rect 33455 5025 33495 5065
rect 33805 5025 33845 5065
rect 34155 5025 34195 5065
rect 34505 5025 34545 5065
rect 34855 5025 34895 5065
rect 35205 5025 35245 5065
rect 35555 5025 35595 5065
rect 35905 5025 35945 5065
rect 36255 5025 36295 5065
rect 27505 4675 27545 4715
rect 27855 4675 27895 4715
rect 28205 4675 28245 4715
rect 28555 4675 28595 4715
rect 28905 4675 28945 4715
rect 29255 4675 29295 4715
rect 29605 4675 29645 4715
rect 29955 4675 29995 4715
rect 30305 4675 30345 4715
rect 33455 4675 33495 4715
rect 33805 4675 33845 4715
rect 34155 4675 34195 4715
rect 34505 4675 34545 4715
rect 34855 4675 34895 4715
rect 35205 4675 35245 4715
rect 35555 4675 35595 4715
rect 35905 4675 35945 4715
rect 36255 4675 36295 4715
rect 27505 4325 27545 4365
rect 27855 4325 27895 4365
rect 28205 4325 28245 4365
rect 28555 4325 28595 4365
rect 28905 4325 28945 4365
rect 29255 4325 29295 4365
rect 29605 4325 29645 4365
rect 29955 4325 29995 4365
rect 30305 4325 30345 4365
rect 33455 4325 33495 4365
rect 33805 4325 33845 4365
rect 34155 4325 34195 4365
rect 34505 4325 34545 4365
rect 34855 4325 34895 4365
rect 35205 4325 35245 4365
rect 35555 4325 35595 4365
rect 35905 4325 35945 4365
rect 36255 4325 36295 4365
rect 27505 3975 27545 4015
rect 27855 3975 27895 4015
rect 28205 3975 28245 4015
rect 28555 3975 28595 4015
rect 28905 3975 28945 4015
rect 29255 3975 29295 4015
rect 29605 3975 29645 4015
rect 29955 3975 29995 4015
rect 30305 3975 30345 4015
rect 33455 3975 33495 4015
rect 33805 3975 33845 4015
rect 34155 3975 34195 4015
rect 34505 3975 34545 4015
rect 34855 3975 34895 4015
rect 35205 3975 35245 4015
rect 35555 3975 35595 4015
rect 35905 3975 35945 4015
rect 36255 3975 36295 4015
rect 27505 3625 27545 3665
rect 27855 3625 27895 3665
rect 28205 3625 28245 3665
rect 28555 3625 28595 3665
rect 28905 3625 28945 3665
rect 34855 3625 34895 3665
rect 35205 3625 35245 3665
rect 35555 3625 35595 3665
rect 35905 3625 35945 3665
rect 36255 3625 36295 3665
rect 27505 3275 27545 3315
rect 27855 3275 27895 3315
rect 28205 3275 28245 3315
rect 28555 3275 28595 3315
rect 28905 3275 28945 3315
rect 34855 3275 34895 3315
rect 35205 3275 35245 3315
rect 35555 3275 35595 3315
rect 35905 3275 35945 3315
rect 36255 3275 36295 3315
rect 27505 2925 27545 2965
rect 27855 2925 27895 2965
rect 28205 2925 28245 2965
rect 28555 2925 28595 2965
rect 28905 2925 28945 2965
rect 34855 2925 34895 2965
rect 35205 2925 35245 2965
rect 35555 2925 35595 2965
rect 35905 2925 35945 2965
rect 36255 2925 36295 2965
rect 27505 2575 27545 2615
rect 27855 2575 27895 2615
rect 28205 2575 28245 2615
rect 28555 2575 28595 2615
rect 28905 2575 28945 2615
rect 34855 2575 34895 2615
rect 35205 2575 35245 2615
rect 35555 2575 35595 2615
rect 35905 2575 35945 2615
rect 36255 2575 36295 2615
rect 27505 2225 27545 2265
rect 27855 2225 27895 2265
rect 28205 2225 28245 2265
rect 28555 2225 28595 2265
rect 28905 2225 28945 2265
rect 34855 2225 34895 2265
rect 35205 2225 35245 2265
rect 35555 2225 35595 2265
rect 35905 2225 35945 2265
rect 36255 2225 36295 2265
rect 27505 1875 27545 1915
rect 27855 1875 27895 1915
rect 28205 1875 28245 1915
rect 28555 1875 28595 1915
rect 28905 1875 28945 1915
rect 34855 1875 34895 1915
rect 35205 1875 35245 1915
rect 35555 1875 35595 1915
rect 35905 1875 35945 1915
rect 36255 1875 36295 1915
rect 27505 1525 27545 1565
rect 27855 1525 27895 1565
rect 28205 1525 28245 1565
rect 28555 1525 28595 1565
rect 28905 1525 28945 1565
rect 34855 1525 34895 1565
rect 35205 1525 35245 1565
rect 35555 1525 35595 1565
rect 35905 1525 35945 1565
rect 36255 1525 36295 1565
rect 27505 1175 27545 1215
rect 27855 1175 27895 1215
rect 28205 1175 28245 1215
rect 28555 1175 28595 1215
rect 28905 1175 28945 1215
rect 34855 1175 34895 1215
rect 35205 1175 35245 1215
rect 35555 1175 35595 1215
rect 35905 1175 35945 1215
rect 36255 1175 36295 1215
rect 27505 825 27545 865
rect 27855 825 27895 865
rect 28205 825 28245 865
rect 28555 825 28595 865
rect 28905 825 28945 865
rect 34855 825 34895 865
rect 35205 825 35245 865
rect 35555 825 35595 865
rect 35905 825 35945 865
rect 36255 825 36295 865
rect 27505 475 27545 515
rect 27855 475 27895 515
rect 28205 475 28245 515
rect 28555 475 28595 515
rect 28905 475 28945 515
rect 34855 475 34895 515
rect 35205 475 35245 515
rect 35555 475 35595 515
rect 35905 475 35945 515
rect 36255 475 36295 515
rect 27505 125 27545 165
rect 27855 125 27895 165
rect 28205 125 28245 165
rect 28555 125 28595 165
rect 28905 125 28945 165
rect 29255 125 29295 165
rect 29605 125 29645 165
rect 29955 125 29995 165
rect 30305 125 30345 165
rect 30655 125 30695 165
rect 31005 125 31045 165
rect 31355 125 31395 165
rect 31705 125 31745 165
rect 32055 125 32095 165
rect 32405 125 32445 165
rect 32755 125 32795 165
rect 33105 125 33145 165
rect 33455 125 33495 165
rect 33805 125 33845 165
rect 34155 125 34195 165
rect 34505 125 34545 165
rect 34855 125 34895 165
rect 35205 125 35245 165
rect 35555 125 35595 165
rect 35905 125 35945 165
rect 36255 125 36295 165
rect 27505 -225 27545 -185
rect 27855 -225 27895 -185
rect 28205 -225 28245 -185
rect 28555 -225 28595 -185
rect 28905 -225 28945 -185
rect 29255 -225 29295 -185
rect 29605 -225 29645 -185
rect 29955 -225 29995 -185
rect 30305 -225 30345 -185
rect 30655 -225 30695 -185
rect 31005 -225 31045 -185
rect 31355 -225 31395 -185
rect 31705 -225 31745 -185
rect 32055 -225 32095 -185
rect 32405 -225 32445 -185
rect 32755 -225 32795 -185
rect 33105 -225 33145 -185
rect 33455 -225 33495 -185
rect 33805 -225 33845 -185
rect 34155 -225 34195 -185
rect 34505 -225 34545 -185
rect 34855 -225 34895 -185
rect 35205 -225 35245 -185
rect 35555 -225 35595 -185
rect 35905 -225 35945 -185
rect 36255 -225 36295 -185
<< metal4 >>
rect 26855 6190 36545 6195
rect 26855 6150 30785 6190
rect 30825 6150 36545 6190
rect 26855 6145 36545 6150
rect 27500 5765 28250 5770
rect 27500 5725 27505 5765
rect 27545 5725 27855 5765
rect 27895 5725 28205 5765
rect 28245 5725 28250 5765
rect 27500 5720 28250 5725
rect 28200 5420 28250 5720
rect 28550 5765 28600 5770
rect 28550 5725 28555 5765
rect 28595 5725 28600 5765
rect 28550 5420 28600 5725
rect 28900 5765 28950 5770
rect 28900 5725 28905 5765
rect 28945 5725 28950 5765
rect 28900 5420 28950 5725
rect 29250 5765 29300 5770
rect 29250 5725 29255 5765
rect 29295 5725 29300 5765
rect 29250 5420 29300 5725
rect 29600 5765 29650 5770
rect 29600 5725 29605 5765
rect 29645 5725 29650 5765
rect 29600 5420 29650 5725
rect 29950 5765 30000 5770
rect 29950 5725 29955 5765
rect 29995 5725 30000 5765
rect 29950 5420 30000 5725
rect 30300 5765 30350 5770
rect 30300 5725 30305 5765
rect 30345 5725 30350 5765
rect 30300 5420 30350 5725
rect 30650 5765 30700 5770
rect 30650 5725 30655 5765
rect 30695 5725 30700 5765
rect 30650 5420 30700 5725
rect 31000 5765 31050 5770
rect 31000 5725 31005 5765
rect 31045 5725 31050 5765
rect 31000 5420 31050 5725
rect 31350 5765 31400 5770
rect 31350 5725 31355 5765
rect 31395 5725 31400 5765
rect 31350 5420 31400 5725
rect 31700 5765 31750 5770
rect 31700 5725 31705 5765
rect 31745 5725 31750 5765
rect 31700 5420 31750 5725
rect 27500 5415 31750 5420
rect 27500 5375 27505 5415
rect 27545 5375 27855 5415
rect 27895 5375 28205 5415
rect 28245 5375 28555 5415
rect 28595 5375 28905 5415
rect 28945 5375 29255 5415
rect 29295 5375 29605 5415
rect 29645 5375 29955 5415
rect 29995 5375 30305 5415
rect 30345 5375 30655 5415
rect 30695 5375 31005 5415
rect 31045 5375 31355 5415
rect 31395 5375 31705 5415
rect 31745 5375 31750 5415
rect 27500 5370 31750 5375
rect 32050 5765 32100 5770
rect 32050 5725 32055 5765
rect 32095 5725 32100 5765
rect 32050 5420 32100 5725
rect 32400 5765 32450 5770
rect 32400 5725 32405 5765
rect 32445 5725 32450 5765
rect 32400 5420 32450 5725
rect 32750 5765 32800 5770
rect 32750 5725 32755 5765
rect 32795 5725 32800 5765
rect 32750 5420 32800 5725
rect 33100 5765 33150 5770
rect 33100 5725 33105 5765
rect 33145 5725 33150 5765
rect 33100 5420 33150 5725
rect 33450 5765 33500 5770
rect 33450 5725 33455 5765
rect 33495 5725 33500 5765
rect 33450 5420 33500 5725
rect 33800 5765 33850 5770
rect 33800 5725 33805 5765
rect 33845 5725 33850 5765
rect 33800 5420 33850 5725
rect 34150 5765 34200 5770
rect 34150 5725 34155 5765
rect 34195 5725 34200 5765
rect 34150 5420 34200 5725
rect 34500 5765 34550 5770
rect 34500 5725 34505 5765
rect 34545 5725 34550 5765
rect 34500 5420 34550 5725
rect 34850 5765 34900 5770
rect 34850 5725 34855 5765
rect 34895 5725 34900 5765
rect 34850 5420 34900 5725
rect 35200 5765 35250 5770
rect 35200 5725 35205 5765
rect 35245 5725 35250 5765
rect 35200 5420 35250 5725
rect 35550 5765 36300 5770
rect 35550 5725 35555 5765
rect 35595 5725 35905 5765
rect 35945 5725 36255 5765
rect 36295 5725 36300 5765
rect 35550 5720 36300 5725
rect 35550 5420 35600 5720
rect 32050 5415 36300 5420
rect 32050 5375 32055 5415
rect 32095 5375 32405 5415
rect 32445 5375 32755 5415
rect 32795 5375 33105 5415
rect 33145 5375 33455 5415
rect 33495 5375 33805 5415
rect 33845 5375 34155 5415
rect 34195 5375 34505 5415
rect 34545 5375 34855 5415
rect 34895 5375 35205 5415
rect 35245 5375 35555 5415
rect 35595 5375 35905 5415
rect 35945 5375 36255 5415
rect 36295 5375 36300 5415
rect 32050 5370 36300 5375
rect 28200 5070 28250 5370
rect 27500 5065 28950 5070
rect 27500 5025 27505 5065
rect 27545 5025 27855 5065
rect 27895 5025 28205 5065
rect 28245 5025 28555 5065
rect 28595 5025 28905 5065
rect 28945 5025 28950 5065
rect 27500 5020 28950 5025
rect 29250 5065 29300 5370
rect 29250 5025 29255 5065
rect 29295 5025 29300 5065
rect 28200 4720 28250 5020
rect 27500 4715 28950 4720
rect 27500 4675 27505 4715
rect 27545 4675 27855 4715
rect 27895 4675 28205 4715
rect 28245 4675 28555 4715
rect 28595 4675 28905 4715
rect 28945 4675 28950 4715
rect 27500 4670 28950 4675
rect 29250 4715 29300 5025
rect 29250 4675 29255 4715
rect 29295 4675 29300 4715
rect 28200 4370 28250 4670
rect 27500 4365 28950 4370
rect 27500 4325 27505 4365
rect 27545 4325 27855 4365
rect 27895 4325 28205 4365
rect 28245 4325 28555 4365
rect 28595 4325 28905 4365
rect 28945 4325 28950 4365
rect 27500 4320 28950 4325
rect 29250 4365 29300 4675
rect 29250 4325 29255 4365
rect 29295 4325 29300 4365
rect 28200 4020 28250 4320
rect 27500 4015 28950 4020
rect 27500 3975 27505 4015
rect 27545 3975 27855 4015
rect 27895 3975 28205 4015
rect 28245 3975 28555 4015
rect 28595 3975 28905 4015
rect 28945 3975 28950 4015
rect 27500 3970 28950 3975
rect 29250 4015 29300 4325
rect 29250 3975 29255 4015
rect 29295 3975 29300 4015
rect 29250 3970 29300 3975
rect 29600 5065 29650 5370
rect 29600 5025 29605 5065
rect 29645 5025 29650 5065
rect 29600 4715 29650 5025
rect 29600 4675 29605 4715
rect 29645 4675 29650 4715
rect 29600 4365 29650 4675
rect 29600 4325 29605 4365
rect 29645 4325 29650 4365
rect 29600 4015 29650 4325
rect 29600 3975 29605 4015
rect 29645 3975 29650 4015
rect 29600 3970 29650 3975
rect 29950 5065 30000 5370
rect 29950 5025 29955 5065
rect 29995 5025 30000 5065
rect 29950 4715 30000 5025
rect 29950 4675 29955 4715
rect 29995 4675 30000 4715
rect 29950 4365 30000 4675
rect 29950 4325 29955 4365
rect 29995 4325 30000 4365
rect 29950 4015 30000 4325
rect 29950 3975 29955 4015
rect 29995 3975 30000 4015
rect 29950 3970 30000 3975
rect 30300 5065 30350 5370
rect 30300 5025 30305 5065
rect 30345 5025 30350 5065
rect 30300 4715 30350 5025
rect 30300 4675 30305 4715
rect 30345 4675 30350 4715
rect 30300 4365 30350 4675
rect 30300 4325 30305 4365
rect 30345 4325 30350 4365
rect 30300 4015 30350 4325
rect 30300 3975 30305 4015
rect 30345 3975 30350 4015
rect 30300 3970 30350 3975
rect 33450 5065 33500 5370
rect 33450 5025 33455 5065
rect 33495 5025 33500 5065
rect 33450 4715 33500 5025
rect 33450 4675 33455 4715
rect 33495 4675 33500 4715
rect 33450 4365 33500 4675
rect 33450 4325 33455 4365
rect 33495 4325 33500 4365
rect 33450 4015 33500 4325
rect 33450 3975 33455 4015
rect 33495 3975 33500 4015
rect 33450 3970 33500 3975
rect 33800 5065 33850 5370
rect 33800 5025 33805 5065
rect 33845 5025 33850 5065
rect 33800 4715 33850 5025
rect 33800 4675 33805 4715
rect 33845 4675 33850 4715
rect 33800 4365 33850 4675
rect 33800 4325 33805 4365
rect 33845 4325 33850 4365
rect 33800 4015 33850 4325
rect 33800 3975 33805 4015
rect 33845 3975 33850 4015
rect 33800 3970 33850 3975
rect 34150 5065 34200 5370
rect 34150 5025 34155 5065
rect 34195 5025 34200 5065
rect 34150 4715 34200 5025
rect 34150 4675 34155 4715
rect 34195 4675 34200 4715
rect 34150 4365 34200 4675
rect 34150 4325 34155 4365
rect 34195 4325 34200 4365
rect 34150 4015 34200 4325
rect 34150 3975 34155 4015
rect 34195 3975 34200 4015
rect 34150 3970 34200 3975
rect 34500 5065 34550 5370
rect 35550 5070 35600 5370
rect 34500 5025 34505 5065
rect 34545 5025 34550 5065
rect 34500 4715 34550 5025
rect 34850 5065 36300 5070
rect 34850 5025 34855 5065
rect 34895 5025 35205 5065
rect 35245 5025 35555 5065
rect 35595 5025 35905 5065
rect 35945 5025 36255 5065
rect 36295 5025 36300 5065
rect 34850 5020 36300 5025
rect 35550 4720 35600 5020
rect 34500 4675 34505 4715
rect 34545 4675 34550 4715
rect 34500 4365 34550 4675
rect 34850 4715 36300 4720
rect 34850 4675 34855 4715
rect 34895 4675 35205 4715
rect 35245 4675 35555 4715
rect 35595 4675 35905 4715
rect 35945 4675 36255 4715
rect 36295 4675 36300 4715
rect 34850 4670 36300 4675
rect 35550 4370 35600 4670
rect 34500 4325 34505 4365
rect 34545 4325 34550 4365
rect 34500 4015 34550 4325
rect 34850 4365 36300 4370
rect 34850 4325 34855 4365
rect 34895 4325 35205 4365
rect 35245 4325 35555 4365
rect 35595 4325 35905 4365
rect 35945 4325 36255 4365
rect 36295 4325 36300 4365
rect 34850 4320 36300 4325
rect 35550 4020 35600 4320
rect 34500 3975 34505 4015
rect 34545 3975 34550 4015
rect 34500 3970 34550 3975
rect 34850 4015 36300 4020
rect 34850 3975 34855 4015
rect 34895 3975 35205 4015
rect 35245 3975 35555 4015
rect 35595 3975 35905 4015
rect 35945 3975 36255 4015
rect 36295 3975 36300 4015
rect 34850 3970 36300 3975
rect 28200 3670 28250 3970
rect 35550 3670 35600 3970
rect 27500 3665 28950 3670
rect 27500 3625 27505 3665
rect 27545 3625 27855 3665
rect 27895 3625 28205 3665
rect 28245 3625 28555 3665
rect 28595 3625 28905 3665
rect 28945 3625 28950 3665
rect 27500 3620 28950 3625
rect 34850 3665 36300 3670
rect 34850 3625 34855 3665
rect 34895 3625 35205 3665
rect 35245 3625 35555 3665
rect 35595 3625 35905 3665
rect 35945 3625 36255 3665
rect 36295 3625 36300 3665
rect 34850 3620 36300 3625
rect 28200 3320 28250 3620
rect 35550 3320 35600 3620
rect 27500 3315 28950 3320
rect 27500 3275 27505 3315
rect 27545 3275 27855 3315
rect 27895 3275 28205 3315
rect 28245 3275 28555 3315
rect 28595 3275 28905 3315
rect 28945 3275 28950 3315
rect 27500 3270 28950 3275
rect 34850 3315 36300 3320
rect 34850 3275 34855 3315
rect 34895 3275 35205 3315
rect 35245 3275 35555 3315
rect 35595 3275 35905 3315
rect 35945 3275 36255 3315
rect 36295 3275 36300 3315
rect 34850 3270 36300 3275
rect 28200 2970 28250 3270
rect 35550 2970 35600 3270
rect 27500 2965 28950 2970
rect 27500 2925 27505 2965
rect 27545 2925 27855 2965
rect 27895 2925 28205 2965
rect 28245 2925 28555 2965
rect 28595 2925 28905 2965
rect 28945 2925 28950 2965
rect 27500 2920 28950 2925
rect 34850 2965 36300 2970
rect 34850 2925 34855 2965
rect 34895 2925 35205 2965
rect 35245 2925 35555 2965
rect 35595 2925 35905 2965
rect 35945 2925 36255 2965
rect 36295 2925 36300 2965
rect 34850 2920 36300 2925
rect 28200 2620 28250 2920
rect 35550 2620 35600 2920
rect 27500 2615 28950 2620
rect 27500 2575 27505 2615
rect 27545 2575 27855 2615
rect 27895 2575 28205 2615
rect 28245 2575 28555 2615
rect 28595 2575 28905 2615
rect 28945 2575 28950 2615
rect 27500 2570 28950 2575
rect 34850 2615 36300 2620
rect 34850 2575 34855 2615
rect 34895 2575 35205 2615
rect 35245 2575 35555 2615
rect 35595 2575 35905 2615
rect 35945 2575 36255 2615
rect 36295 2575 36300 2615
rect 34850 2570 36300 2575
rect 28200 2270 28250 2570
rect 35550 2270 35600 2570
rect 27500 2265 29360 2270
rect 27500 2225 27505 2265
rect 27545 2225 27855 2265
rect 27895 2225 28205 2265
rect 28245 2225 28555 2265
rect 28595 2225 28905 2265
rect 28945 2225 29315 2265
rect 29355 2225 29360 2265
rect 27500 2220 29360 2225
rect 34440 2265 36300 2270
rect 34440 2225 34445 2265
rect 34485 2225 34855 2265
rect 34895 2225 35205 2265
rect 35245 2225 35555 2265
rect 35595 2225 35905 2265
rect 35945 2225 36255 2265
rect 36295 2225 36300 2265
rect 34440 2220 36300 2225
rect 28200 1920 28250 2220
rect 35550 1920 35600 2220
rect 27500 1915 28950 1920
rect 27500 1875 27505 1915
rect 27545 1875 27855 1915
rect 27895 1875 28205 1915
rect 28245 1875 28555 1915
rect 28595 1875 28905 1915
rect 28945 1875 28950 1915
rect 27500 1870 28950 1875
rect 34855 1915 36300 1920
rect 34895 1875 35205 1915
rect 35245 1875 35555 1915
rect 35595 1875 35905 1915
rect 35945 1875 36255 1915
rect 36295 1875 36300 1915
rect 34855 1870 36300 1875
rect 28200 1570 28250 1870
rect 35550 1570 35600 1870
rect 27500 1565 28950 1570
rect 27500 1525 27505 1565
rect 27545 1525 27855 1565
rect 27895 1525 28205 1565
rect 28245 1525 28555 1565
rect 28595 1525 28905 1565
rect 28945 1525 28950 1565
rect 27500 1520 28950 1525
rect 34850 1565 36300 1570
rect 34850 1525 34855 1565
rect 34895 1525 35205 1565
rect 35245 1525 35555 1565
rect 35595 1525 35905 1565
rect 35945 1525 36255 1565
rect 36295 1525 36300 1565
rect 34850 1520 36300 1525
rect 28200 1220 28250 1520
rect 35550 1220 35600 1520
rect 27500 1215 28950 1220
rect 27500 1175 27505 1215
rect 27545 1175 27855 1215
rect 27895 1175 28205 1215
rect 28245 1175 28555 1215
rect 28595 1175 28905 1215
rect 28945 1175 28950 1215
rect 27500 1170 28950 1175
rect 34850 1215 36300 1220
rect 34850 1175 34855 1215
rect 34895 1175 35205 1215
rect 35245 1175 35555 1215
rect 35595 1175 35905 1215
rect 35945 1175 36255 1215
rect 36295 1175 36300 1215
rect 34850 1170 36300 1175
rect 28200 870 28250 1170
rect 35550 870 35600 1170
rect 27500 865 28950 870
rect 27500 825 27505 865
rect 27545 825 27855 865
rect 27895 825 28205 865
rect 28245 825 28555 865
rect 28595 825 28905 865
rect 28945 825 28950 865
rect 27500 820 28950 825
rect 34850 865 36300 870
rect 34850 825 34855 865
rect 34895 825 35205 865
rect 35245 825 35555 865
rect 35595 825 35905 865
rect 35945 825 36255 865
rect 36295 825 36300 865
rect 34850 820 36300 825
rect 28200 520 28250 820
rect 35550 520 35600 820
rect 27500 515 28950 520
rect 27500 475 27505 515
rect 27545 475 27855 515
rect 27895 475 28205 515
rect 28245 475 28555 515
rect 28595 475 28905 515
rect 28945 475 28950 515
rect 27500 470 28950 475
rect 34850 515 36300 520
rect 34850 475 34855 515
rect 34895 475 35205 515
rect 35245 475 35555 515
rect 35595 475 35905 515
rect 35945 475 36255 515
rect 36295 475 36300 515
rect 34850 470 36300 475
rect 28200 170 28250 470
rect 35550 170 35600 470
rect 27500 165 31750 170
rect 27500 125 27505 165
rect 27545 125 27855 165
rect 27895 125 28205 165
rect 28245 125 28555 165
rect 28595 125 28905 165
rect 28945 125 29255 165
rect 29295 125 29605 165
rect 29645 125 29955 165
rect 29995 125 30305 165
rect 30345 125 30655 165
rect 30695 125 31005 165
rect 31045 125 31355 165
rect 31395 125 31705 165
rect 31745 125 31750 165
rect 27500 120 31750 125
rect 28200 -180 28250 120
rect 27500 -185 28250 -180
rect 27500 -225 27505 -185
rect 27545 -225 27855 -185
rect 27895 -225 28205 -185
rect 28245 -225 28250 -185
rect 27500 -230 28250 -225
rect 28550 -185 28600 120
rect 28550 -225 28555 -185
rect 28595 -225 28600 -185
rect 28550 -230 28600 -225
rect 28900 -185 28950 120
rect 28900 -225 28905 -185
rect 28945 -225 28950 -185
rect 28900 -230 28950 -225
rect 29250 -185 29300 120
rect 29250 -225 29255 -185
rect 29295 -225 29300 -185
rect 29250 -230 29300 -225
rect 29600 -185 29650 120
rect 29600 -225 29605 -185
rect 29645 -225 29650 -185
rect 29600 -230 29650 -225
rect 29950 -185 30000 120
rect 29950 -225 29955 -185
rect 29995 -225 30000 -185
rect 29950 -230 30000 -225
rect 30300 -185 30350 120
rect 30300 -225 30305 -185
rect 30345 -225 30350 -185
rect 30300 -230 30350 -225
rect 30650 -185 30700 120
rect 30650 -225 30655 -185
rect 30695 -225 30700 -185
rect 30650 -230 30700 -225
rect 31000 -185 31050 120
rect 31000 -225 31005 -185
rect 31045 -225 31050 -185
rect 31000 -230 31050 -225
rect 31350 -185 31400 120
rect 31350 -225 31355 -185
rect 31395 -225 31400 -185
rect 31350 -230 31400 -225
rect 31700 -185 31750 120
rect 31700 -225 31705 -185
rect 31745 -225 31750 -185
rect 31700 -230 31750 -225
rect 32050 165 36300 170
rect 32050 125 32055 165
rect 32095 125 32405 165
rect 32445 125 32755 165
rect 32795 125 33105 165
rect 33145 125 33455 165
rect 33495 125 33805 165
rect 33845 125 34155 165
rect 34195 125 34505 165
rect 34545 125 34855 165
rect 34895 125 35205 165
rect 35245 125 35555 165
rect 35595 125 35905 165
rect 35945 125 36255 165
rect 36295 125 36300 165
rect 32050 120 36300 125
rect 32050 -185 32100 120
rect 32050 -225 32055 -185
rect 32095 -225 32100 -185
rect 32050 -230 32100 -225
rect 32400 -185 32450 120
rect 32400 -225 32405 -185
rect 32445 -225 32450 -185
rect 32400 -230 32450 -225
rect 32750 -185 32800 120
rect 32750 -225 32755 -185
rect 32795 -225 32800 -185
rect 32750 -230 32800 -225
rect 33100 -185 33150 120
rect 33100 -225 33105 -185
rect 33145 -225 33150 -185
rect 33100 -230 33150 -225
rect 33450 -185 33500 120
rect 33450 -225 33455 -185
rect 33495 -225 33500 -185
rect 33450 -230 33500 -225
rect 33800 -185 33850 120
rect 33800 -225 33805 -185
rect 33845 -225 33850 -185
rect 33800 -230 33850 -225
rect 34150 -185 34200 120
rect 34150 -225 34155 -185
rect 34195 -225 34200 -185
rect 34150 -230 34200 -225
rect 34500 -185 34550 120
rect 34500 -225 34505 -185
rect 34545 -225 34550 -185
rect 34500 -230 34550 -225
rect 34850 -185 34900 120
rect 34850 -225 34855 -185
rect 34895 -225 34900 -185
rect 34850 -230 34900 -225
rect 35200 -185 35250 120
rect 35200 -225 35205 -185
rect 35245 -225 35250 -185
rect 35200 -230 35250 -225
rect 35550 -180 35600 120
rect 35550 -185 36300 -180
rect 35550 -225 35555 -185
rect 35595 -225 35905 -185
rect 35945 -225 36255 -185
rect 36295 -225 36300 -185
rect 35550 -230 36300 -225
rect 26855 -510 36545 -505
rect 26855 -550 30785 -510
rect 30825 -550 36545 -510
rect 26855 -555 36545 -550
<< labels >>
flabel metal2 29335 1670 29335 1670 5 FreeSans 200 0 0 -80 VOUT-
flabel metal2 34465 1670 34465 1670 5 FreeSans 200 0 0 -80 VOUT+
flabel metal3 29605 3795 29605 3795 7 FreeSans 200 0 -80 0 cap_res_X
flabel metal3 34195 3795 34195 3795 3 FreeSans 200 0 80 0 cap_res_Y
flabel metal2 33950 2300 33950 2300 1 FreeSans 200 0 0 80 V_CMFB_S4
flabel metal2 33995 2490 33995 2490 1 FreeSans 200 0 0 80 V_CMFB_S3
flabel metal2 29855 2300 29855 2300 1 FreeSans 200 0 0 80 V_CMFB_S2
flabel metal2 29810 2490 29810 2490 1 FreeSans 200 0 0 80 V_CMFB_S1
flabel metal1 31900 2385 31900 2385 5 FreeSans 200 0 0 -80 Vb2
flabel metal4 26855 6170 26855 6170 7 FreeSans 800 0 -400 0 VDDA
flabel metal4 26855 -530 26855 -530 7 FreeSans 800 0 -400 0 GNDA
flabel metal1 31710 2360 31710 2360 3 FreeSans 200 0 80 0 X
flabel metal1 32090 2360 32090 2360 7 FreeSans 200 0 -80 0 Y
flabel metal1 30850 2235 30850 2235 1 FreeSans 200 0 0 80 Vb1
flabel metal2 31190 1880 31190 1880 7 FreeSans 200 0 -80 0 VD1
flabel metal2 30920 1745 30920 1745 7 FreeSans 200 0 -80 0 VIN-
flabel metal2 30920 1525 30920 1525 7 FreeSans 200 0 -80 0 VIN+
flabel metal1 31555 1840 31555 1840 3 FreeSans 200 0 80 0 VD2
flabel metal2 32720 1410 32720 1410 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal1 31900 1375 31900 1375 3 FreeSans 200 0 80 0 V_p_mir
flabel metal1 31845 1300 31845 1300 3 FreeSans 200 0 80 0 V_tail_gate
flabel metal1 32215 1360 32215 1360 3 FreeSans 200 0 80 0 V_p
flabel metal1 31840 3150 31840 3150 5 FreeSans 200 0 0 -80 Vb3
flabel metal1 32415 3005 32415 3005 3 FreeSans 200 0 80 0 VD4
flabel metal1 31260 3035 31260 3035 7 FreeSans 200 0 -80 0 VD3
flabel metal2 32080 3745 32080 3745 7 FreeSans 200 0 -80 0 err_amp_out
flabel metal2 33000 3835 33000 3835 3 FreeSans 200 0 80 0 err_amp_mir
flabel metal1 32910 4015 32910 4015 3 FreeSans 200 0 80 0 V_tot
flabel metal2 30950 3895 30950 3895 7 FreeSans 200 0 -80 0 V_err_amp_ref
flabel metal1 31450 4135 31450 4135 3 FreeSans 200 0 80 0 V_err_mir_p
flabel metal2 32070 4925 32070 4925 1 FreeSans 200 0 0 80 Vb2_Vb3
flabel metal1 32410 4170 32410 4170 3 FreeSans 200 0 80 0 V_err_p
flabel metal1 31375 4180 31375 4180 7 FreeSans 200 0 -80 0 V_err_gate
<< end >>
