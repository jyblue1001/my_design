magic
tech sky130A
timestamp 1739381150
<< nmos >>
rect 3460 1925 3475 1975
rect 3525 1925 3540 1975
rect 3590 1925 3605 1975
rect 3655 1925 3670 1975
rect 3720 1925 3735 1975
rect 3785 1925 3800 1975
<< ndiff >>
rect 3410 1960 3460 1975
rect 3410 1940 3425 1960
rect 3445 1940 3460 1960
rect 3410 1925 3460 1940
rect 3475 1960 3525 1975
rect 3475 1940 3490 1960
rect 3510 1940 3525 1960
rect 3475 1925 3525 1940
rect 3540 1960 3590 1975
rect 3540 1940 3555 1960
rect 3575 1940 3590 1960
rect 3540 1925 3590 1940
rect 3605 1960 3655 1975
rect 3605 1940 3620 1960
rect 3640 1940 3655 1960
rect 3605 1925 3655 1940
rect 3670 1960 3720 1975
rect 3670 1940 3685 1960
rect 3705 1940 3720 1960
rect 3670 1925 3720 1940
rect 3735 1960 3785 1975
rect 3735 1940 3750 1960
rect 3770 1940 3785 1960
rect 3735 1925 3785 1940
rect 3800 1960 3850 1975
rect 3800 1940 3815 1960
rect 3835 1940 3850 1960
rect 3800 1925 3850 1940
<< ndiffc >>
rect 3425 1940 3445 1960
rect 3490 1940 3510 1960
rect 3555 1940 3575 1960
rect 3620 1940 3640 1960
rect 3685 1940 3705 1960
rect 3750 1940 3770 1960
rect 3815 1940 3835 1960
<< psubdiff >>
rect 3360 1960 3410 1975
rect 3360 1940 3375 1960
rect 3395 1940 3410 1960
rect 3360 1925 3410 1940
rect 3850 1960 3900 1975
rect 3850 1940 3865 1960
rect 3885 1940 3900 1960
rect 3850 1925 3900 1940
<< psubdiffcont >>
rect 3375 1940 3395 1960
rect 3865 1940 3885 1960
<< poly >>
rect 3545 2020 3585 2030
rect 3545 2000 3555 2020
rect 3575 2000 3585 2020
rect 3460 1975 3475 1990
rect 3525 1985 3735 2000
rect 3525 1975 3540 1985
rect 3590 1975 3605 1985
rect 3655 1975 3670 1985
rect 3720 1975 3735 1985
rect 3785 1975 3800 1990
rect 3460 1910 3475 1925
rect 3525 1910 3540 1925
rect 3590 1910 3605 1925
rect 3655 1910 3670 1925
rect 3720 1910 3735 1925
rect 3785 1910 3800 1925
rect 3445 1900 3485 1910
rect 3445 1880 3455 1900
rect 3475 1880 3485 1900
rect 3445 1870 3485 1880
rect 3775 1900 3815 1910
rect 3775 1880 3785 1900
rect 3805 1880 3815 1900
rect 3775 1870 3815 1880
<< polycont >>
rect 3555 2000 3575 2020
rect 3455 1880 3475 1900
rect 3785 1880 3805 1900
<< locali >>
rect 3545 2020 3585 2030
rect 3545 2000 3555 2020
rect 3575 2000 3585 2020
rect 3545 1990 3585 2000
rect 3555 1970 3575 1990
rect 3685 1970 3705 2100
rect 3365 1960 3455 1970
rect 3365 1940 3375 1960
rect 3395 1940 3425 1960
rect 3445 1940 3455 1960
rect 3365 1930 3455 1940
rect 3480 1960 3520 1970
rect 3480 1940 3490 1960
rect 3510 1940 3520 1960
rect 3480 1930 3520 1940
rect 3545 1960 3585 1970
rect 3545 1940 3555 1960
rect 3575 1940 3585 1960
rect 3545 1930 3585 1940
rect 3610 1960 3650 1970
rect 3610 1940 3620 1960
rect 3640 1940 3650 1960
rect 3610 1930 3650 1940
rect 3675 1960 3715 1970
rect 3675 1940 3685 1960
rect 3705 1940 3715 1960
rect 3675 1930 3715 1940
rect 3740 1960 3780 1970
rect 3740 1940 3750 1960
rect 3770 1940 3780 1960
rect 3740 1930 3780 1940
rect 3805 1960 3895 1970
rect 3805 1940 3815 1960
rect 3835 1940 3865 1960
rect 3885 1940 3895 1960
rect 3805 1930 3895 1940
rect 3425 1910 3445 1930
rect 3490 1910 3510 1930
rect 3620 1910 3640 1930
rect 3750 1910 3770 1930
rect 3815 1910 3835 1930
rect 3425 1900 3835 1910
rect 3425 1890 3455 1900
rect 3445 1880 3455 1890
rect 3475 1890 3785 1900
rect 3475 1880 3485 1890
rect 3445 1870 3485 1880
rect 3620 1810 3640 1890
rect 3775 1880 3785 1890
rect 3805 1890 3835 1900
rect 3805 1880 3815 1890
rect 3775 1870 3815 1880
rect 3250 1790 3280 1810
rect 3300 1790 3330 1810
rect 3350 1790 3380 1810
rect 3400 1790 3430 1810
rect 3450 1790 3480 1810
rect 3500 1790 3530 1810
rect 3550 1790 3580 1810
rect 3600 1790 3630 1810
rect 3650 1790 3680 1810
rect 3700 1790 3730 1810
rect 3750 1790 3780 1810
rect 3800 1790 3830 1810
rect 3850 1790 3880 1810
rect 3900 1790 3920 1810
<< viali >>
rect 3280 1790 3300 1810
rect 3330 1790 3350 1810
rect 3380 1790 3400 1810
rect 3430 1790 3450 1810
rect 3480 1790 3500 1810
rect 3530 1790 3550 1810
rect 3580 1790 3600 1810
rect 3630 1790 3650 1810
rect 3680 1790 3700 1810
rect 3730 1790 3750 1810
rect 3780 1790 3800 1810
rect 3830 1790 3850 1810
rect 3880 1790 3900 1810
<< metal1 >>
rect 3250 1810 3920 1820
rect 3250 1790 3280 1810
rect 3300 1790 3330 1810
rect 3350 1790 3380 1810
rect 3400 1790 3430 1810
rect 3450 1790 3480 1810
rect 3500 1790 3530 1810
rect 3550 1790 3580 1810
rect 3600 1790 3630 1810
rect 3650 1790 3680 1810
rect 3700 1790 3730 1810
rect 3750 1790 3780 1810
rect 3800 1790 3830 1810
rect 3850 1790 3880 1810
rect 3900 1790 3920 1810
rect 3250 1780 3920 1790
<< labels >>
flabel locali 3250 1800 3250 1800 7 FreeSans 400 0 -200 0 GNDA
flabel poly 3665 2000 3665 2000 1 FreeSans 400 0 0 200 GATE
flabel locali 3705 2100 3705 2100 1 FreeSans 400 0 0 200 OTHER
<< end >>
