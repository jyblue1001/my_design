* PEX produced on Sat Feb  1 08:49:04 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from div8.ext - technology: sky130A

.subckt div8 VOUT VIN VDDA GNDA
X0 VDDA.t21 div2.t2 div2_3_1.A.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1 div2_3_0.C.t2 div2_3_0.CLK.t3 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 div2.t1 div2_3_1.C.t4 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X3 div2_3_0.A.t1 div2_3_0.CLK.t4 div2_3_0.B.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 GNDA.t27 div2_3_0.CLK.t5 div2_3_0.C.t1 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X5 VDDA.t19 div2.t3 div2_3_2.CLK.t1 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 div2_3_0.CLK.t1 div4.t2 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X7 div2_3_0.B.t0 VOUT.t2 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X8 GNDA.t9 div2_3_1.CLK.t3 div2_3_1.C.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X9 GNDA.t15 div4.t3 div2_3_0.CLK.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 div2_3_1.C.t0 div2_3_1.CLK.t4 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VDDA.t15 VOUT.t3 div2_3_0.A.t0 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 div2_3_2.C.t3 div2_3_2.A.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 GNDA.t17 div2_3_1.CLK.t5 div2_3_1.C.t2 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 VDDA.t5 VIN.t0 div2_3_1.CLK.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X15 div2_3_1.C.t3 div2_3_1.A.t2 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X16 GNDA.t11 div2_3_2.CLK.t3 div2_3_2.C.t2 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 div4.t0 div2_3_2.C.t4 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 div4.t1 div2_3_2.CLK.t4 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X19 GNDA.t35 div2_3_2.CLK.t5 div2_3_2.C.t1 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X20 div2_3_1.A.t1 div2_3_1.CLK.t6 div2_3_1.B.t0 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 div2_3_2.C.t0 div2_3_2.CLK.t6 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X22 div2_3_2.A.t0 div2_3_2.CLK.t7 div2_3_2.B.t0 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 div2_3_1.B.t1 div2.t4 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X24 VDDA.t25 div4.t4 div2_3_0.CLK.t2 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X25 div2_3_2.B.t1 div4.t5 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X26 div2.t0 div2_3_1.CLK.t7 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X27 div2_3_0.C.t3 div2_3_0.A.t2 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X28 GNDA.t7 VIN.t1 div2_3_1.CLK.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X29 div2_3_2.CLK.t0 div2.t5 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X30 VOUT.t1 div2_3_0.CLK.t6 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X31 GNDA.t21 div2.t6 div2_3_2.CLK.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X32 VOUT.t0 div2_3_0.C.t4 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X33 div2_3_1.CLK.t2 VIN.t2 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X34 GNDA.t25 div2_3_0.CLK.t7 div2_3_0.C.t0 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X35 VDDA.t11 div4.t6 div2_3_2.A.t1 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 div2.t2 div2.t4 819.4
R1 div2.n0 div2.t0 663.801
R2 div2.n0 div2.t2 489.168
R3 div2.t3 div2.t5 401.668
R4 div2.n1 div2.t1 270.12
R5 div2.n2 div2.t3 257.067
R6 div2_3_2.VIN div2.n2 216.9
R7 div2.n2 div2.t6 208.868
R8 div2.n3 div2_3_2.VIN 192.167
R9 div2.n1 div2.n0 67.2005
R10 div2.n3 div2.n1 25.6005
R11 div2_3_1.VOUT div2.n3 4.8005
R12 div2_3_1.A.n0 div2_3_1.A.t0 713.933
R13 div2_3_1.A.n0 div2_3_1.A.t2 314.233
R14 div2_3_1.A.t1 div2_3_1.A.n0 308.2
R15 VDDA.t24 VDDA.t8 2080.95
R16 VDDA.t6 VDDA.t18 2080.95
R17 VDDA.t14 VDDA.t12 1130.95
R18 VDDA.t16 VDDA.t10 1130.95
R19 VDDA.t20 VDDA.t26 1130.95
R20 VDDA.n3 VDDA.t28 927.381
R21 VDDA.t2 VDDA.n16 927.381
R22 VDDA.n17 VDDA.t22 927.381
R23 VDDA.n4 VDDA.t1 667.62
R24 VDDA.n1 VDDA.t7 663.801
R25 VDDA.n2 VDDA.t9 663.801
R26 VDDA.n3 VDDA.t0 610.715
R27 VDDA.n16 VDDA.t8 610.715
R28 VDDA.n17 VDDA.t6 610.715
R29 VDDA.n23 VDDA.n22 594.301
R30 VDDA.n21 VDDA.n20 594.301
R31 VDDA.n11 VDDA.n10 594.301
R32 VDDA.n13 VDDA.n12 594.301
R33 VDDA.n8 VDDA.n7 594.301
R34 VDDA.n6 VDDA.n5 594.301
R35 VDDA.t28 VDDA.t14 497.62
R36 VDDA.t12 VDDA.t24 497.62
R37 VDDA.t10 VDDA.t2 497.62
R38 VDDA.t18 VDDA.t16 497.62
R39 VDDA.t22 VDDA.t20 497.62
R40 VDDA.t26 VDDA.t4 497.62
R41 VDDA.n4 VDDA.n3 373.781
R42 VDDA.n16 VDDA.n15 370
R43 VDDA.n18 VDDA.n17 370
R44 VDDA.n22 VDDA.t27 78.8005
R45 VDDA.n22 VDDA.t5 78.8005
R46 VDDA.n20 VDDA.t23 78.8005
R47 VDDA.n20 VDDA.t21 78.8005
R48 VDDA.n10 VDDA.t17 78.8005
R49 VDDA.n10 VDDA.t19 78.8005
R50 VDDA.n12 VDDA.t3 78.8005
R51 VDDA.n12 VDDA.t11 78.8005
R52 VDDA.n7 VDDA.t13 78.8005
R53 VDDA.n7 VDDA.t25 78.8005
R54 VDDA.n5 VDDA.t29 78.8005
R55 VDDA.n5 VDDA.t15 78.8005
R56 VDDA.n18 VDDA.n1 12.8005
R57 VDDA.n15 VDDA.n2 12.8005
R58 VDDA.n9 VDDA.n2 9.3005
R59 VDDA.n15 VDDA.n14 9.3005
R60 VDDA.n1 VDDA.n0 9.3005
R61 VDDA.n19 VDDA.n18 9.3005
R62 VDDA.n6 VDDA.n4 3.10124
R63 VDDA.n9 VDDA 0.4755
R64 VDDA VDDA.n0 0.4755
R65 VDDA.n8 VDDA.n6 0.4505
R66 VDDA.n13 VDDA.n11 0.4505
R67 VDDA.n23 VDDA.n21 0.4505
R68 VDDA.n14 VDDA.n13 0.3255
R69 VDDA.n21 VDDA.n19 0.3255
R70 VDDA VDDA.n8 0.238
R71 VDDA.n11 VDDA 0.238
R72 VDDA VDDA.n23 0.238
R73 VDDA.n14 VDDA.n9 0.1005
R74 VDDA.n19 VDDA.n0 0.1005
R75 div2_3_0.CLK.n5 div2_3_0.CLK.t2 723.534
R76 div2_3_0.CLK.n4 div2_3_0.CLK.t1 723.534
R77 div2_3_0.CLK.n0 div2_3_0.CLK.t6 369.534
R78 div2_3_0.CLK.n3 div2_3_0.CLK.n2 366.856
R79 div2_3_0.CLK.t0 div2_3_0.CLK.n5 254.333
R80 div2_3_0.CLK.n3 div2_3_0.CLK.t4 190.123
R81 div2_3_0.CLK.n4 div2_3_0.CLK.n3 187.201
R82 div2_3_0.CLK.n1 div2_3_0.CLK.n0 176.733
R83 div2_3_0.CLK.n2 div2_3_0.CLK.n1 176.733
R84 div2_3_0.CLK.n0 div2_3_0.CLK.t7 112.468
R85 div2_3_0.CLK.n2 div2_3_0.CLK.t5 112.468
R86 div2_3_0.CLK.n1 div2_3_0.CLK.t3 112.468
R87 div2_3_0.CLK.n5 div2_3_0.CLK.n4 70.4005
R88 GNDA.t26 GNDA.t28 4683.87
R89 GNDA.t36 GNDA.t10 4683.87
R90 GNDA.t16 GNDA.t31 4683.87
R91 GNDA.n1 GNDA.t18 3947.35
R92 GNDA.n13 GNDA.t14 2767.74
R93 GNDA.t2 GNDA.n13 2767.74
R94 GNDA.n14 GNDA.t20 2767.74
R95 GNDA.n14 GNDA.t32 2767.74
R96 GNDA.t18 GNDA.t24 1561.29
R97 GNDA.t24 GNDA.t29 1561.29
R98 GNDA.t29 GNDA.t26 1561.29
R99 GNDA.t28 GNDA.t0 1561.29
R100 GNDA.t0 GNDA.t14 1561.29
R101 GNDA.t34 GNDA.t2 1561.29
R102 GNDA.t37 GNDA.t34 1561.29
R103 GNDA.t10 GNDA.t37 1561.29
R104 GNDA.t12 GNDA.t36 1561.29
R105 GNDA.t20 GNDA.t12 1561.29
R106 GNDA.t32 GNDA.t8 1561.29
R107 GNDA.t8 GNDA.t4 1561.29
R108 GNDA.t4 GNDA.t16 1561.29
R109 GNDA.t31 GNDA.t22 1561.29
R110 GNDA.t22 GNDA.t6 1561.29
R111 GNDA.n13 GNDA.n12 1179.3
R112 GNDA.n15 GNDA.n14 1179.3
R113 GNDA.n21 GNDA.n20 194.3
R114 GNDA.n19 GNDA.n18 194.3
R115 GNDA.n17 GNDA.n16 194.3
R116 GNDA.n7 GNDA.n6 194.3
R117 GNDA.n9 GNDA.n8 194.3
R118 GNDA.n11 GNDA.n10 194.3
R119 GNDA.n5 GNDA.n4 194.3
R120 GNDA.n3 GNDA.n2 194.3
R121 GNDA.n1 GNDA.n0 194.3
R122 GNDA.n20 GNDA.t23 48.0005
R123 GNDA.n20 GNDA.t7 48.0005
R124 GNDA.n18 GNDA.t5 48.0005
R125 GNDA.n18 GNDA.t17 48.0005
R126 GNDA.n16 GNDA.t33 48.0005
R127 GNDA.n16 GNDA.t9 48.0005
R128 GNDA.n6 GNDA.t13 48.0005
R129 GNDA.n6 GNDA.t21 48.0005
R130 GNDA.n8 GNDA.t38 48.0005
R131 GNDA.n8 GNDA.t11 48.0005
R132 GNDA.n10 GNDA.t3 48.0005
R133 GNDA.n10 GNDA.t35 48.0005
R134 GNDA.n4 GNDA.t1 48.0005
R135 GNDA.n4 GNDA.t15 48.0005
R136 GNDA.n2 GNDA.t30 48.0005
R137 GNDA.n2 GNDA.t27 48.0005
R138 GNDA.n0 GNDA.t19 48.0005
R139 GNDA.n0 GNDA.t25 48.0005
R140 GNDA.n5 GNDA.n3 0.688
R141 GNDA.n9 GNDA.n7 0.688
R142 GNDA.n21 GNDA.n19 0.688
R143 GNDA.n12 GNDA.n11 0.313
R144 GNDA.n17 GNDA.n15 0.313
R145 GNDA.n3 GNDA.n1 0.2755
R146 GNDA.n11 GNDA.n9 0.2755
R147 GNDA.n19 GNDA.n17 0.2755
R148 GNDA GNDA.n5 0.238
R149 GNDA.n7 GNDA 0.238
R150 GNDA GNDA.n21 0.238
R151 GNDA.n12 GNDA 0.0755
R152 GNDA.n15 GNDA 0.0755
R153 div2_3_0.C.n0 div2_3_0.C.t3 721.4
R154 div2_3_0.C.n1 div2_3_0.C.t4 349.433
R155 div2_3_0.C.n0 div2_3_0.C.t1 276.733
R156 div2_3_0.C.n2 div2_3_0.C.n1 206.333
R157 div2_3_0.C.n1 div2_3_0.C.n0 48.0005
R158 div2_3_0.C.n2 div2_3_0.C.t0 48.0005
R159 div2_3_0.C.t2 div2_3_0.C.n2 48.0005
R160 div2_3_1.C.n0 div2_3_1.C.t3 721.4
R161 div2_3_1.C.n1 div2_3_1.C.t4 349.433
R162 div2_3_1.C.n0 div2_3_1.C.t2 276.733
R163 div2_3_1.C.n2 div2_3_1.C.n1 206.333
R164 div2_3_1.C.n1 div2_3_1.C.n0 48.0005
R165 div2_3_1.C.n2 div2_3_1.C.t1 48.0005
R166 div2_3_1.C.t0 div2_3_1.C.n2 48.0005
R167 div2_3_0.B.t0 div2_3_0.B.t1 96.0005
R168 div2_3_0.A.n0 div2_3_0.A.t0 713.933
R169 div2_3_0.A.n0 div2_3_0.A.t2 314.233
R170 div2_3_0.A.t1 div2_3_0.A.n0 308.2
R171 div2_3_2.CLK.n4 div2_3_2.CLK.t0 723.534
R172 div2_3_2.CLK.t1 div2_3_2.CLK.n5 723.534
R173 div2_3_2.CLK.n0 div2_3_2.CLK.t4 369.534
R174 div2_3_2.CLK.n3 div2_3_2.CLK.n2 366.856
R175 div2_3_2.CLK.n5 div2_3_2.CLK.t2 254.333
R176 div2_3_2.CLK.n3 div2_3_2.CLK.t7 190.123
R177 div2_3_2.CLK.n4 div2_3_2.CLK.n3 187.201
R178 div2_3_2.CLK.n1 div2_3_2.CLK.n0 176.733
R179 div2_3_2.CLK.n2 div2_3_2.CLK.n1 176.733
R180 div2_3_2.CLK.n0 div2_3_2.CLK.t5 112.468
R181 div2_3_2.CLK.n2 div2_3_2.CLK.t3 112.468
R182 div2_3_2.CLK.n1 div2_3_2.CLK.t6 112.468
R183 div2_3_2.CLK.n5 div2_3_2.CLK.n4 70.4005
R184 div4.t6 div4.t5 819.4
R185 div4.n0 div4.t1 663.801
R186 div4.n0 div4.t6 489.168
R187 div4.t4 div4.t2 401.668
R188 div4.n1 div4.t0 270.12
R189 div4.n2 div4.t4 257.067
R190 div2_3_0.VIN div4.n2 216.9
R191 div4.n2 div4.t3 208.868
R192 div4.n3 div2_3_0.VIN 192.167
R193 div4.n1 div4.n0 67.2005
R194 div4.n3 div4.n1 25.6005
R195 div2_3_2.VOUT div4.n3 4.8005
R196 VOUT.t3 VOUT.t2 819.4
R197 VOUT.n0 VOUT.t1 663.801
R198 VOUT.n0 VOUT.t3 489.168
R199 VOUT.n1 VOUT.t0 270.12
R200 VOUT.n2 VOUT 208.233
R201 VOUT.n1 VOUT.n0 67.2005
R202 VOUT.n2 VOUT.n1 25.6005
R203 VOUT VOUT.n2 4.8005
R204 div2_3_1.CLK.n5 div2_3_1.CLK.t1 723.534
R205 div2_3_1.CLK.n4 div2_3_1.CLK.t2 723.534
R206 div2_3_1.CLK.n0 div2_3_1.CLK.t7 369.534
R207 div2_3_1.CLK.n3 div2_3_1.CLK.n2 366.856
R208 div2_3_1.CLK.t0 div2_3_1.CLK.n5 254.333
R209 div2_3_1.CLK.n3 div2_3_1.CLK.t6 190.123
R210 div2_3_1.CLK.n4 div2_3_1.CLK.n3 187.201
R211 div2_3_1.CLK.n1 div2_3_1.CLK.n0 176.733
R212 div2_3_1.CLK.n2 div2_3_1.CLK.n1 176.733
R213 div2_3_1.CLK.n0 div2_3_1.CLK.t3 112.468
R214 div2_3_1.CLK.n2 div2_3_1.CLK.t5 112.468
R215 div2_3_1.CLK.n1 div2_3_1.CLK.t4 112.468
R216 div2_3_1.CLK.n5 div2_3_1.CLK.n4 70.4005
R217 div2_3_2.A.n0 div2_3_2.A.t1 713.933
R218 div2_3_2.A.n0 div2_3_2.A.t2 314.233
R219 div2_3_2.A.t0 div2_3_2.A.n0 308.2
R220 div2_3_2.C.n2 div2_3_2.C.t3 721.4
R221 div2_3_2.C.n1 div2_3_2.C.t4 349.433
R222 div2_3_2.C.t2 div2_3_2.C.n2 276.733
R223 div2_3_2.C.n1 div2_3_2.C.n0 206.333
R224 div2_3_2.C.n0 div2_3_2.C.t1 48.0005
R225 div2_3_2.C.n0 div2_3_2.C.t0 48.0005
R226 div2_3_2.C.n2 div2_3_2.C.n1 48.0005
R227 VIN.t0 VIN.t2 401.668
R228 VIN.n0 VIN.t0 257.067
R229 VIN VIN.n0 216.9
R230 VIN.n0 VIN.t1 208.868
R231 div2_3_1.B.t0 div2_3_1.B.t1 96.0005
R232 div2_3_2.B.t0 div2_3_2.B.t1 96.0005
C0 VIN VDDA 0.125773f
C1 VOUT VDDA 0.488104f
C2 VIN GNDA 0.304628f
C3 VOUT GNDA 0.792323f
C4 VDDA GNDA 3.90136f
.ends

