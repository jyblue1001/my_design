magic
tech sky130A
timestamp 1754062532
<< error_s >>
rect 6305 11350 6335 11405
rect 4305 10210 4345 10214
rect 4415 10210 4455 10214
rect 4525 10210 4565 10214
rect 4635 10210 4675 10214
rect 4310 10196 4340 10200
rect 4420 10196 4450 10200
rect 4530 10196 4560 10200
rect 4640 10196 4670 10200
rect 4515 4540 4579 4544
rect 4525 4526 4565 4530
rect 5166 4525 5196 4570
rect 5191 4524 5196 4525
rect 5166 4520 5196 4524
rect 5205 4510 5210 4520
rect 5152 4506 5210 4510
rect 2160 1755 2190 1760
rect 2160 1730 2210 1755
rect 3625 1745 3634 1759
rect 6790 1755 6820 1760
rect 2180 1725 2210 1730
rect 6770 1730 6820 1755
rect 6770 1725 6800 1730
rect 1500 1394 1510 1470
rect 1486 1380 1524 1394
rect 1486 1370 1600 1380
rect 1486 1356 1524 1370
rect 2196 1330 2205 1540
rect 2210 1316 2219 1540
rect 6761 1316 6770 1540
rect 6775 1330 6784 1540
<< metal1 >>
rect 2320 20910 2380 20925
rect 2320 20880 2335 20910
rect 2365 20880 2380 20910
rect 2320 20845 2380 20880
rect 2320 20815 2335 20845
rect 2365 20815 2380 20845
rect 2320 20775 2380 20815
rect 2320 20745 2335 20775
rect 2365 20745 2380 20775
rect 2320 20705 2380 20745
rect 2320 20675 2335 20705
rect 2365 20675 2380 20705
rect 2320 20635 2380 20675
rect 2320 20605 2335 20635
rect 2365 20605 2380 20635
rect 2320 20570 2380 20605
rect 2320 20540 2335 20570
rect 2365 20540 2380 20570
rect 2320 20510 2380 20540
rect 2320 20480 2335 20510
rect 2365 20480 2380 20510
rect 2320 20445 2380 20480
rect 2320 20415 2335 20445
rect 2365 20415 2380 20445
rect 2320 20375 2380 20415
rect 2320 20345 2335 20375
rect 2365 20345 2380 20375
rect 2320 20305 2380 20345
rect 2320 20275 2335 20305
rect 2365 20275 2380 20305
rect 2320 20235 2380 20275
rect 2320 20205 2335 20235
rect 2365 20205 2380 20235
rect 2320 20170 2380 20205
rect 2320 20140 2335 20170
rect 2365 20140 2380 20170
rect 2320 20110 2380 20140
rect 2320 20080 2335 20110
rect 2365 20080 2380 20110
rect 2320 20045 2380 20080
rect 2320 20015 2335 20045
rect 2365 20015 2380 20045
rect 2320 19975 2380 20015
rect 2320 19945 2335 19975
rect 2365 19945 2380 19975
rect 2320 19905 2380 19945
rect 2320 19875 2335 19905
rect 2365 19875 2380 19905
rect 2320 19835 2380 19875
rect 2320 19805 2335 19835
rect 2365 19805 2380 19835
rect 2320 19770 2380 19805
rect 2320 19740 2335 19770
rect 2365 19740 2380 19770
rect 2320 19710 2380 19740
rect 2320 19680 2335 19710
rect 2365 19680 2380 19710
rect 2320 19645 2380 19680
rect 2320 19615 2335 19645
rect 2365 19615 2380 19645
rect 2320 19575 2380 19615
rect 2320 19545 2335 19575
rect 2365 19545 2380 19575
rect 2320 19505 2380 19545
rect 2320 19475 2335 19505
rect 2365 19475 2380 19505
rect 2320 19435 2380 19475
rect 2320 19405 2335 19435
rect 2365 19405 2380 19435
rect 2320 19370 2380 19405
rect 2320 19340 2335 19370
rect 2365 19340 2380 19370
rect 2320 19310 2380 19340
rect 2320 19280 2335 19310
rect 2365 19280 2380 19310
rect 2320 19245 2380 19280
rect 2320 19215 2335 19245
rect 2365 19215 2380 19245
rect 2320 19175 2380 19215
rect 2320 19145 2335 19175
rect 2365 19145 2380 19175
rect 2320 19105 2380 19145
rect 2320 19075 2335 19105
rect 2365 19075 2380 19105
rect 2320 19035 2380 19075
rect 2320 19005 2335 19035
rect 2365 19005 2380 19035
rect 2320 18970 2380 19005
rect 2320 18940 2335 18970
rect 2365 18940 2380 18970
rect 2320 18910 2380 18940
rect 2320 18880 2335 18910
rect 2365 18880 2380 18910
rect 2320 18845 2380 18880
rect 2320 18815 2335 18845
rect 2365 18815 2380 18845
rect 2320 18775 2380 18815
rect 2320 18745 2335 18775
rect 2365 18745 2380 18775
rect 2320 18705 2380 18745
rect 2320 18675 2335 18705
rect 2365 18675 2380 18705
rect 2320 18635 2380 18675
rect 2320 18605 2335 18635
rect 2365 18605 2380 18635
rect 2320 18570 2380 18605
rect 2320 18540 2335 18570
rect 2365 18540 2380 18570
rect 2320 18510 2380 18540
rect 2320 18480 2335 18510
rect 2365 18480 2380 18510
rect 2320 18445 2380 18480
rect 2320 18415 2335 18445
rect 2365 18415 2380 18445
rect 2320 18375 2380 18415
rect 2320 18345 2335 18375
rect 2365 18345 2380 18375
rect 2320 18305 2380 18345
rect 2320 18275 2335 18305
rect 2365 18275 2380 18305
rect 2320 18235 2380 18275
rect 2320 18205 2335 18235
rect 2365 18205 2380 18235
rect 2320 18170 2380 18205
rect 2320 18140 2335 18170
rect 2365 18140 2380 18170
rect 2320 18110 2380 18140
rect 2320 18080 2335 18110
rect 2365 18080 2380 18110
rect 2320 18045 2380 18080
rect 2320 18015 2335 18045
rect 2365 18015 2380 18045
rect 2320 17975 2380 18015
rect 2320 17945 2335 17975
rect 2365 17945 2380 17975
rect 2320 17905 2380 17945
rect 2320 17875 2335 17905
rect 2365 17875 2380 17905
rect 2320 17835 2380 17875
rect 2320 17805 2335 17835
rect 2365 17805 2380 17835
rect 2320 17770 2380 17805
rect 2320 17740 2335 17770
rect 2365 17740 2380 17770
rect 2320 17725 2380 17740
rect 6690 20910 6750 20925
rect 6690 20880 6705 20910
rect 6735 20880 6750 20910
rect 6690 20845 6750 20880
rect 6690 20815 6705 20845
rect 6735 20815 6750 20845
rect 6690 20775 6750 20815
rect 6690 20745 6705 20775
rect 6735 20745 6750 20775
rect 6690 20705 6750 20745
rect 6690 20675 6705 20705
rect 6735 20675 6750 20705
rect 6690 20635 6750 20675
rect 6690 20605 6705 20635
rect 6735 20605 6750 20635
rect 6690 20570 6750 20605
rect 6690 20540 6705 20570
rect 6735 20540 6750 20570
rect 6690 20510 6750 20540
rect 6690 20480 6705 20510
rect 6735 20480 6750 20510
rect 6690 20445 6750 20480
rect 6690 20415 6705 20445
rect 6735 20415 6750 20445
rect 6690 20375 6750 20415
rect 6690 20345 6705 20375
rect 6735 20345 6750 20375
rect 6690 20305 6750 20345
rect 6690 20275 6705 20305
rect 6735 20275 6750 20305
rect 6690 20235 6750 20275
rect 6690 20205 6705 20235
rect 6735 20205 6750 20235
rect 6690 20170 6750 20205
rect 6690 20140 6705 20170
rect 6735 20140 6750 20170
rect 6690 20110 6750 20140
rect 6690 20080 6705 20110
rect 6735 20080 6750 20110
rect 6690 20045 6750 20080
rect 6690 20015 6705 20045
rect 6735 20015 6750 20045
rect 6690 19975 6750 20015
rect 6690 19945 6705 19975
rect 6735 19945 6750 19975
rect 6690 19905 6750 19945
rect 6690 19875 6705 19905
rect 6735 19875 6750 19905
rect 6690 19835 6750 19875
rect 6690 19805 6705 19835
rect 6735 19805 6750 19835
rect 6690 19770 6750 19805
rect 6690 19740 6705 19770
rect 6735 19740 6750 19770
rect 6690 19710 6750 19740
rect 6690 19680 6705 19710
rect 6735 19680 6750 19710
rect 6690 19645 6750 19680
rect 6690 19615 6705 19645
rect 6735 19615 6750 19645
rect 6690 19575 6750 19615
rect 6690 19545 6705 19575
rect 6735 19545 6750 19575
rect 6690 19505 6750 19545
rect 6690 19475 6705 19505
rect 6735 19475 6750 19505
rect 6690 19435 6750 19475
rect 6690 19405 6705 19435
rect 6735 19405 6750 19435
rect 6690 19370 6750 19405
rect 6690 19340 6705 19370
rect 6735 19340 6750 19370
rect 6690 19310 6750 19340
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2330 15780 2370 17725
rect 2330 15750 2335 15780
rect 2365 15750 2370 15780
rect 2330 12760 2370 15750
rect 2330 12730 2335 12760
rect 2365 12730 2370 12760
rect 2330 12720 2370 12730
rect 2330 12690 2335 12720
rect 2365 12690 2370 12720
rect 2330 12600 2370 12690
rect 2330 12570 2335 12600
rect 2365 12570 2370 12600
rect 2330 12560 2370 12570
rect 2330 12530 2335 12560
rect 2365 12530 2370 12560
rect 2330 12520 2370 12530
rect 2330 12490 2335 12520
rect 2365 12490 2370 12520
rect 2330 12485 2370 12490
rect 2385 15925 2425 15930
rect 2385 15895 2390 15925
rect 2420 15895 2425 15925
rect 2385 9650 2425 15895
rect 6700 15705 6740 17725
rect 6700 15675 6705 15705
rect 6735 15675 6740 15705
rect 6700 13005 6740 15675
rect 6700 12975 6705 13005
rect 6735 12975 6740 13005
rect 6700 12965 6740 12975
rect 6700 12935 6705 12965
rect 6735 12935 6740 12965
rect 6700 12925 6740 12935
rect 6700 12895 6705 12925
rect 6735 12895 6740 12925
rect 6700 12890 6740 12895
rect 2475 12725 2515 12765
rect 2540 12725 2560 12765
rect 2650 12725 2670 12765
rect 2725 12725 2745 12765
rect 2790 12725 2830 12765
rect 2855 12725 2875 12765
rect 2935 12725 2955 12765
rect 2475 12525 2515 12605
rect 2540 12525 2560 12605
rect 2650 12525 2670 12605
rect 2725 12525 2745 12605
rect 2790 12525 2830 12605
rect 2855 12525 2875 12605
rect 2935 12525 2955 12605
rect 6590 12200 6630 12205
rect 6590 12170 6595 12200
rect 6625 12170 6630 12200
rect 5725 12085 5755 12165
rect 6000 12085 6020 12165
rect 6055 12085 6075 12165
rect 6100 12085 6120 12165
rect 6155 12085 6175 12165
rect 6230 12085 6250 12165
rect 6310 12085 6330 12165
rect 6465 12085 6505 12165
rect 6535 12085 6555 12165
rect 6590 12160 6630 12170
rect 6590 12130 6595 12160
rect 6625 12130 6630 12160
rect 6590 12120 6630 12130
rect 6590 12090 6595 12120
rect 6625 12090 6630 12120
rect 6300 11485 6340 11490
rect 6300 11455 6305 11485
rect 6335 11455 6340 11485
rect 6300 11445 6340 11455
rect 6300 11415 6305 11445
rect 6335 11415 6340 11445
rect 6300 11405 6340 11415
rect 6300 11375 6305 11405
rect 6335 11375 6340 11405
rect 2990 10085 3030 10090
rect 2990 10055 2995 10085
rect 3025 10055 3030 10085
rect 2990 10050 3030 10055
rect -120 9635 0 9650
rect -120 9605 -75 9635
rect -45 9605 0 9635
rect -120 9570 0 9605
rect -120 9540 -75 9570
rect -45 9540 0 9570
rect -120 9500 0 9540
rect -120 9470 -75 9500
rect -45 9470 0 9500
rect -120 9430 0 9470
rect -120 9400 -75 9430
rect -45 9400 0 9430
rect -120 9360 0 9400
rect -120 9330 -75 9360
rect -45 9330 0 9360
rect -120 9295 0 9330
rect -120 9265 -75 9295
rect -45 9265 0 9295
rect -120 9235 0 9265
rect -120 9205 -75 9235
rect -45 9205 0 9235
rect -120 9170 0 9205
rect -120 9140 -75 9170
rect -45 9140 0 9170
rect -120 9100 0 9140
rect -120 9070 -75 9100
rect -45 9070 0 9100
rect -120 9030 0 9070
rect -120 9000 -75 9030
rect -45 9000 0 9030
rect -120 8960 0 9000
rect -120 8930 -75 8960
rect -45 8930 0 8960
rect -120 8895 0 8930
rect -120 8865 -75 8895
rect -45 8865 0 8895
rect -120 8835 0 8865
rect -120 8805 -75 8835
rect -45 8805 0 8835
rect -120 8770 0 8805
rect -120 8740 -75 8770
rect -45 8740 0 8770
rect -120 8700 0 8740
rect -120 8670 -75 8700
rect -45 8670 0 8700
rect -120 8630 0 8670
rect -120 8600 -75 8630
rect -45 8600 0 8630
rect -120 8560 0 8600
rect -120 8530 -75 8560
rect -45 8530 0 8560
rect -120 8495 0 8530
rect -120 8465 -75 8495
rect -45 8465 0 8495
rect -120 8435 0 8465
rect -120 8405 -75 8435
rect -45 8405 0 8435
rect -120 8370 0 8405
rect -120 8340 -75 8370
rect -45 8340 0 8370
rect -120 8300 0 8340
rect -120 8270 -75 8300
rect -45 8270 0 8300
rect -120 8230 0 8270
rect -120 8200 -75 8230
rect -45 8200 0 8230
rect -120 8160 0 8200
rect -120 8130 -75 8160
rect -45 8130 0 8160
rect -120 8095 0 8130
rect -120 8065 -75 8095
rect -45 8065 0 8095
rect -120 8035 0 8065
rect -120 8005 -75 8035
rect -45 8005 0 8035
rect -120 7970 0 8005
rect -120 7940 -75 7970
rect -45 7940 0 7970
rect -120 7900 0 7940
rect -120 7870 -75 7900
rect -45 7870 0 7900
rect -120 7830 0 7870
rect -120 7800 -75 7830
rect -45 7800 0 7830
rect -120 7760 0 7800
rect -120 7730 -75 7760
rect -45 7730 0 7760
rect -120 7695 0 7730
rect -120 7665 -75 7695
rect -45 7665 0 7695
rect -120 7635 0 7665
rect -120 7605 -75 7635
rect -45 7605 0 7635
rect -120 7570 0 7605
rect -120 7540 -75 7570
rect -45 7540 0 7570
rect -120 7500 0 7540
rect -120 7470 -75 7500
rect -45 7470 0 7500
rect -120 7430 0 7470
rect -120 7400 -75 7430
rect -45 7400 0 7430
rect -120 7360 0 7400
rect -120 7330 -75 7360
rect -45 7330 0 7360
rect -120 7295 0 7330
rect -120 7265 -75 7295
rect -45 7265 0 7295
rect -120 7235 0 7265
rect -120 7205 -75 7235
rect -45 7205 0 7235
rect -120 7170 0 7205
rect -120 7140 -75 7170
rect -45 7140 0 7170
rect -120 7100 0 7140
rect -120 7070 -75 7100
rect -45 7070 0 7100
rect -120 7030 0 7070
rect -120 7000 -75 7030
rect -45 7000 0 7030
rect -120 6960 0 7000
rect -120 6930 -75 6960
rect -45 6930 0 6960
rect -120 6895 0 6930
rect -120 6865 -75 6895
rect -45 6865 0 6895
rect -120 6835 0 6865
rect -120 6805 -75 6835
rect -45 6805 0 6835
rect -120 6770 0 6805
rect -120 6740 -75 6770
rect -45 6740 0 6770
rect -120 6700 0 6740
rect -120 6670 -75 6700
rect -45 6670 0 6700
rect -120 6630 0 6670
rect -120 6600 -75 6630
rect -45 6600 0 6630
rect -120 6560 0 6600
rect -120 6530 -75 6560
rect -45 6530 0 6560
rect -120 6495 0 6530
rect -120 6465 -75 6495
rect -45 6465 0 6495
rect -120 6210 0 6465
rect 230 9635 350 9650
rect 230 9605 275 9635
rect 305 9605 350 9635
rect 230 9570 350 9605
rect 230 9540 275 9570
rect 305 9540 350 9570
rect 230 9500 350 9540
rect 230 9470 275 9500
rect 305 9470 350 9500
rect 230 9430 350 9470
rect 230 9400 275 9430
rect 305 9400 350 9430
rect 230 9360 350 9400
rect 230 9330 275 9360
rect 305 9330 350 9360
rect 230 9295 350 9330
rect 230 9265 275 9295
rect 305 9265 350 9295
rect 230 9235 350 9265
rect 230 9205 275 9235
rect 305 9205 350 9235
rect 230 9170 350 9205
rect 230 9140 275 9170
rect 305 9140 350 9170
rect 230 9100 350 9140
rect 230 9070 275 9100
rect 305 9070 350 9100
rect 230 9030 350 9070
rect 230 9000 275 9030
rect 305 9000 350 9030
rect 230 8960 350 9000
rect 230 8930 275 8960
rect 305 8930 350 8960
rect 230 8895 350 8930
rect 230 8865 275 8895
rect 305 8865 350 8895
rect 230 8835 350 8865
rect 230 8805 275 8835
rect 305 8805 350 8835
rect 230 8770 350 8805
rect 230 8740 275 8770
rect 305 8740 350 8770
rect 230 8700 350 8740
rect 230 8670 275 8700
rect 305 8670 350 8700
rect 230 8630 350 8670
rect 230 8600 275 8630
rect 305 8600 350 8630
rect 230 8560 350 8600
rect 230 8530 275 8560
rect 305 8530 350 8560
rect 230 8495 350 8530
rect 230 8465 275 8495
rect 305 8465 350 8495
rect 230 8435 350 8465
rect 230 8405 275 8435
rect 305 8405 350 8435
rect 230 8370 350 8405
rect 230 8340 275 8370
rect 305 8340 350 8370
rect 230 8300 350 8340
rect 230 8270 275 8300
rect 305 8270 350 8300
rect 230 8230 350 8270
rect 230 8200 275 8230
rect 305 8200 350 8230
rect 230 8160 350 8200
rect 230 8130 275 8160
rect 305 8130 350 8160
rect 230 8095 350 8130
rect 230 8065 275 8095
rect 305 8065 350 8095
rect 230 8035 350 8065
rect 230 8005 275 8035
rect 305 8005 350 8035
rect 230 7970 350 8005
rect 230 7940 275 7970
rect 305 7940 350 7970
rect 230 7900 350 7940
rect 230 7870 275 7900
rect 305 7870 350 7900
rect 230 7830 350 7870
rect 230 7800 275 7830
rect 305 7800 350 7830
rect 230 7760 350 7800
rect 230 7730 275 7760
rect 305 7730 350 7760
rect 230 7695 350 7730
rect 230 7665 275 7695
rect 305 7665 350 7695
rect 230 7635 350 7665
rect 230 7605 275 7635
rect 305 7605 350 7635
rect 230 7570 350 7605
rect 230 7540 275 7570
rect 305 7540 350 7570
rect 230 7500 350 7540
rect 230 7470 275 7500
rect 305 7470 350 7500
rect 230 7430 350 7470
rect 230 7400 275 7430
rect 305 7400 350 7430
rect 230 7360 350 7400
rect 230 7330 275 7360
rect 305 7330 350 7360
rect 230 7295 350 7330
rect 230 7265 275 7295
rect 305 7265 350 7295
rect 230 7235 350 7265
rect 230 7205 275 7235
rect 305 7205 350 7235
rect 230 7170 350 7205
rect 230 7140 275 7170
rect 305 7140 350 7170
rect 230 7100 350 7140
rect 230 7070 275 7100
rect 305 7070 350 7100
rect 230 7030 350 7070
rect 230 7000 275 7030
rect 305 7000 350 7030
rect 230 6960 350 7000
rect 230 6930 275 6960
rect 305 6930 350 6960
rect 230 6895 350 6930
rect 230 6865 275 6895
rect 305 6865 350 6895
rect 230 6835 350 6865
rect 230 6805 275 6835
rect 305 6805 350 6835
rect 230 6770 350 6805
rect 230 6740 275 6770
rect 305 6740 350 6770
rect 230 6700 350 6740
rect 230 6670 275 6700
rect 305 6670 350 6700
rect 230 6630 350 6670
rect 230 6600 275 6630
rect 305 6600 350 6630
rect 230 6560 350 6600
rect 230 6530 275 6560
rect 305 6530 350 6560
rect 230 6495 350 6530
rect 230 6465 275 6495
rect 305 6465 350 6495
rect 230 6210 350 6465
rect 580 9635 700 9650
rect 580 9605 625 9635
rect 655 9605 700 9635
rect 580 9570 700 9605
rect 580 9540 625 9570
rect 655 9540 700 9570
rect 580 9500 700 9540
rect 580 9470 625 9500
rect 655 9470 700 9500
rect 580 9430 700 9470
rect 580 9400 625 9430
rect 655 9400 700 9430
rect 580 9360 700 9400
rect 580 9330 625 9360
rect 655 9330 700 9360
rect 580 9295 700 9330
rect 580 9265 625 9295
rect 655 9265 700 9295
rect 580 9235 700 9265
rect 580 9205 625 9235
rect 655 9205 700 9235
rect 580 9170 700 9205
rect 580 9140 625 9170
rect 655 9140 700 9170
rect 580 9100 700 9140
rect 580 9070 625 9100
rect 655 9070 700 9100
rect 580 9030 700 9070
rect 580 9000 625 9030
rect 655 9000 700 9030
rect 580 8960 700 9000
rect 580 8930 625 8960
rect 655 8930 700 8960
rect 580 8895 700 8930
rect 580 8865 625 8895
rect 655 8865 700 8895
rect 580 8835 700 8865
rect 580 8805 625 8835
rect 655 8805 700 8835
rect 580 8770 700 8805
rect 580 8740 625 8770
rect 655 8740 700 8770
rect 580 8700 700 8740
rect 580 8670 625 8700
rect 655 8670 700 8700
rect 580 8630 700 8670
rect 580 8600 625 8630
rect 655 8600 700 8630
rect 580 8560 700 8600
rect 580 8530 625 8560
rect 655 8530 700 8560
rect 580 8495 700 8530
rect 580 8465 625 8495
rect 655 8465 700 8495
rect 580 8435 700 8465
rect 580 8405 625 8435
rect 655 8405 700 8435
rect 580 8370 700 8405
rect 580 8340 625 8370
rect 655 8340 700 8370
rect 580 8300 700 8340
rect 580 8270 625 8300
rect 655 8270 700 8300
rect 580 8230 700 8270
rect 580 8200 625 8230
rect 655 8200 700 8230
rect 580 8160 700 8200
rect 580 8130 625 8160
rect 655 8130 700 8160
rect 580 8095 700 8130
rect 580 8065 625 8095
rect 655 8065 700 8095
rect 580 8035 700 8065
rect 580 8005 625 8035
rect 655 8005 700 8035
rect 580 7970 700 8005
rect 580 7940 625 7970
rect 655 7940 700 7970
rect 580 7900 700 7940
rect 580 7870 625 7900
rect 655 7870 700 7900
rect 580 7830 700 7870
rect 580 7800 625 7830
rect 655 7800 700 7830
rect 580 7760 700 7800
rect 580 7730 625 7760
rect 655 7730 700 7760
rect 580 7695 700 7730
rect 580 7665 625 7695
rect 655 7665 700 7695
rect 580 7635 700 7665
rect 580 7605 625 7635
rect 655 7605 700 7635
rect 580 7570 700 7605
rect 580 7540 625 7570
rect 655 7540 700 7570
rect 580 7500 700 7540
rect 580 7470 625 7500
rect 655 7470 700 7500
rect 580 7430 700 7470
rect 580 7400 625 7430
rect 655 7400 700 7430
rect 580 7360 700 7400
rect 580 7330 625 7360
rect 655 7330 700 7360
rect 580 7295 700 7330
rect 580 7265 625 7295
rect 655 7265 700 7295
rect 580 7235 700 7265
rect 580 7205 625 7235
rect 655 7205 700 7235
rect 580 7170 700 7205
rect 580 7140 625 7170
rect 655 7140 700 7170
rect 580 7100 700 7140
rect 580 7070 625 7100
rect 655 7070 700 7100
rect 580 7030 700 7070
rect 580 7000 625 7030
rect 655 7000 700 7030
rect 580 6960 700 7000
rect 580 6930 625 6960
rect 655 6930 700 6960
rect 580 6895 700 6930
rect 580 6865 625 6895
rect 655 6865 700 6895
rect 580 6835 700 6865
rect 580 6805 625 6835
rect 655 6805 700 6835
rect 580 6770 700 6805
rect 580 6740 625 6770
rect 655 6740 700 6770
rect 580 6700 700 6740
rect 580 6670 625 6700
rect 655 6670 700 6700
rect 580 6630 700 6670
rect 580 6600 625 6630
rect 655 6600 700 6630
rect 580 6560 700 6600
rect 580 6530 625 6560
rect 655 6530 700 6560
rect 580 6495 700 6530
rect 580 6465 625 6495
rect 655 6465 700 6495
rect 580 6210 700 6465
rect 1280 9635 1400 9650
rect 1280 9605 1325 9635
rect 1355 9605 1400 9635
rect 1280 9570 1400 9605
rect 1280 9540 1325 9570
rect 1355 9540 1400 9570
rect 1280 9500 1400 9540
rect 1280 9470 1325 9500
rect 1355 9470 1400 9500
rect 1280 9430 1400 9470
rect 1280 9400 1325 9430
rect 1355 9400 1400 9430
rect 1280 9360 1400 9400
rect 1280 9330 1325 9360
rect 1355 9330 1400 9360
rect 1280 9295 1400 9330
rect 1280 9265 1325 9295
rect 1355 9265 1400 9295
rect 1280 9235 1400 9265
rect 1280 9205 1325 9235
rect 1355 9205 1400 9235
rect 1280 9170 1400 9205
rect 1280 9140 1325 9170
rect 1355 9140 1400 9170
rect 1280 9100 1400 9140
rect 1280 9070 1325 9100
rect 1355 9070 1400 9100
rect 1280 9030 1400 9070
rect 1280 9000 1325 9030
rect 1355 9000 1400 9030
rect 1280 8960 1400 9000
rect 1280 8930 1325 8960
rect 1355 8930 1400 8960
rect 1280 8895 1400 8930
rect 1280 8865 1325 8895
rect 1355 8865 1400 8895
rect 1280 8835 1400 8865
rect 1280 8805 1325 8835
rect 1355 8805 1400 8835
rect 1280 8770 1400 8805
rect 1280 8740 1325 8770
rect 1355 8740 1400 8770
rect 1280 8700 1400 8740
rect 1280 8670 1325 8700
rect 1355 8670 1400 8700
rect 1280 8630 1400 8670
rect 1280 8600 1325 8630
rect 1355 8600 1400 8630
rect 1280 8560 1400 8600
rect 1280 8530 1325 8560
rect 1355 8530 1400 8560
rect 1280 8495 1400 8530
rect 1280 8465 1325 8495
rect 1355 8465 1400 8495
rect 1280 8435 1400 8465
rect 1280 8405 1325 8435
rect 1355 8405 1400 8435
rect 1280 8370 1400 8405
rect 1280 8340 1325 8370
rect 1355 8340 1400 8370
rect 1280 8300 1400 8340
rect 1280 8270 1325 8300
rect 1355 8270 1400 8300
rect 1280 8230 1400 8270
rect 1280 8200 1325 8230
rect 1355 8200 1400 8230
rect 1280 8160 1400 8200
rect 1280 8130 1325 8160
rect 1355 8130 1400 8160
rect 1280 8095 1400 8130
rect 1280 8065 1325 8095
rect 1355 8065 1400 8095
rect 1280 8035 1400 8065
rect 1280 8005 1325 8035
rect 1355 8005 1400 8035
rect 1280 7970 1400 8005
rect 1280 7940 1325 7970
rect 1355 7940 1400 7970
rect 1280 7900 1400 7940
rect 1280 7870 1325 7900
rect 1355 7870 1400 7900
rect 1280 7830 1400 7870
rect 1280 7800 1325 7830
rect 1355 7800 1400 7830
rect 1280 7760 1400 7800
rect 1280 7730 1325 7760
rect 1355 7730 1400 7760
rect 1280 7695 1400 7730
rect 1280 7665 1325 7695
rect 1355 7665 1400 7695
rect 1280 7635 1400 7665
rect 1280 7605 1325 7635
rect 1355 7605 1400 7635
rect 1280 7570 1400 7605
rect 1280 7540 1325 7570
rect 1355 7540 1400 7570
rect 1280 7500 1400 7540
rect 1280 7470 1325 7500
rect 1355 7470 1400 7500
rect 1280 7430 1400 7470
rect 1280 7400 1325 7430
rect 1355 7400 1400 7430
rect 1280 7360 1400 7400
rect 1280 7330 1325 7360
rect 1355 7330 1400 7360
rect 1280 7295 1400 7330
rect 1280 7265 1325 7295
rect 1355 7265 1400 7295
rect 1280 7235 1400 7265
rect 1280 7205 1325 7235
rect 1355 7205 1400 7235
rect 1280 7170 1400 7205
rect 1280 7140 1325 7170
rect 1355 7140 1400 7170
rect 1280 7100 1400 7140
rect 1280 7070 1325 7100
rect 1355 7070 1400 7100
rect 1280 7030 1400 7070
rect 1280 7000 1325 7030
rect 1355 7000 1400 7030
rect 1280 6960 1400 7000
rect 1280 6930 1325 6960
rect 1355 6930 1400 6960
rect 1280 6895 1400 6930
rect 1280 6865 1325 6895
rect 1355 6865 1400 6895
rect 1280 6835 1400 6865
rect 1280 6805 1325 6835
rect 1355 6805 1400 6835
rect 1280 6770 1400 6805
rect 1280 6740 1325 6770
rect 1355 6740 1400 6770
rect 1280 6700 1400 6740
rect 1280 6670 1325 6700
rect 1355 6670 1400 6700
rect 1280 6630 1400 6670
rect 1280 6600 1325 6630
rect 1355 6600 1400 6630
rect 1280 6560 1400 6600
rect 1280 6530 1325 6560
rect 1355 6530 1400 6560
rect 1280 6495 1400 6530
rect 1280 6465 1325 6495
rect 1355 6465 1400 6495
rect 1280 6205 1400 6465
rect 1630 9635 1750 9650
rect 1630 9605 1675 9635
rect 1705 9605 1750 9635
rect 1630 9570 1750 9605
rect 1630 9540 1675 9570
rect 1705 9540 1750 9570
rect 1630 9500 1750 9540
rect 1630 9470 1675 9500
rect 1705 9470 1750 9500
rect 1630 9430 1750 9470
rect 1630 9400 1675 9430
rect 1705 9400 1750 9430
rect 1630 9360 1750 9400
rect 1630 9330 1675 9360
rect 1705 9330 1750 9360
rect 1630 9295 1750 9330
rect 1630 9265 1675 9295
rect 1705 9265 1750 9295
rect 1630 9235 1750 9265
rect 1630 9205 1675 9235
rect 1705 9205 1750 9235
rect 1630 9170 1750 9205
rect 1630 9140 1675 9170
rect 1705 9140 1750 9170
rect 1630 9100 1750 9140
rect 1630 9070 1675 9100
rect 1705 9070 1750 9100
rect 1630 9030 1750 9070
rect 1630 9000 1675 9030
rect 1705 9000 1750 9030
rect 1630 8960 1750 9000
rect 1630 8930 1675 8960
rect 1705 8930 1750 8960
rect 1630 8895 1750 8930
rect 1630 8865 1675 8895
rect 1705 8865 1750 8895
rect 1630 8835 1750 8865
rect 1630 8805 1675 8835
rect 1705 8805 1750 8835
rect 1630 8770 1750 8805
rect 1630 8740 1675 8770
rect 1705 8740 1750 8770
rect 1630 8700 1750 8740
rect 1630 8670 1675 8700
rect 1705 8670 1750 8700
rect 1630 8630 1750 8670
rect 1630 8600 1675 8630
rect 1705 8600 1750 8630
rect 1630 8560 1750 8600
rect 1630 8530 1675 8560
rect 1705 8530 1750 8560
rect 1630 8495 1750 8530
rect 1630 8465 1675 8495
rect 1705 8465 1750 8495
rect 1630 8435 1750 8465
rect 1630 8405 1675 8435
rect 1705 8405 1750 8435
rect 1630 8370 1750 8405
rect 1630 8340 1675 8370
rect 1705 8340 1750 8370
rect 1630 8300 1750 8340
rect 1630 8270 1675 8300
rect 1705 8270 1750 8300
rect 1630 8230 1750 8270
rect 1630 8200 1675 8230
rect 1705 8200 1750 8230
rect 1630 8160 1750 8200
rect 1630 8130 1675 8160
rect 1705 8130 1750 8160
rect 1630 8095 1750 8130
rect 1630 8065 1675 8095
rect 1705 8065 1750 8095
rect 1630 8035 1750 8065
rect 1630 8005 1675 8035
rect 1705 8005 1750 8035
rect 1630 7970 1750 8005
rect 1630 7940 1675 7970
rect 1705 7940 1750 7970
rect 1630 7900 1750 7940
rect 1630 7870 1675 7900
rect 1705 7870 1750 7900
rect 1630 7830 1750 7870
rect 1630 7800 1675 7830
rect 1705 7800 1750 7830
rect 1630 7760 1750 7800
rect 1630 7730 1675 7760
rect 1705 7730 1750 7760
rect 1630 7695 1750 7730
rect 1630 7665 1675 7695
rect 1705 7665 1750 7695
rect 1630 7635 1750 7665
rect 1630 7605 1675 7635
rect 1705 7605 1750 7635
rect 1630 7570 1750 7605
rect 1630 7540 1675 7570
rect 1705 7540 1750 7570
rect 1630 7500 1750 7540
rect 1630 7470 1675 7500
rect 1705 7470 1750 7500
rect 1630 7430 1750 7470
rect 1630 7400 1675 7430
rect 1705 7400 1750 7430
rect 1630 7360 1750 7400
rect 1630 7330 1675 7360
rect 1705 7330 1750 7360
rect 1630 7295 1750 7330
rect 1630 7265 1675 7295
rect 1705 7265 1750 7295
rect 1630 7235 1750 7265
rect 1630 7205 1675 7235
rect 1705 7205 1750 7235
rect 1630 7170 1750 7205
rect 1630 7140 1675 7170
rect 1705 7140 1750 7170
rect 1630 7100 1750 7140
rect 1630 7070 1675 7100
rect 1705 7070 1750 7100
rect 1630 7030 1750 7070
rect 1630 7000 1675 7030
rect 1705 7000 1750 7030
rect 1630 6960 1750 7000
rect 1630 6930 1675 6960
rect 1705 6930 1750 6960
rect 1630 6895 1750 6930
rect 1630 6865 1675 6895
rect 1705 6865 1750 6895
rect 1630 6835 1750 6865
rect 1630 6805 1675 6835
rect 1705 6805 1750 6835
rect 1630 6770 1750 6805
rect 1630 6740 1675 6770
rect 1705 6740 1750 6770
rect 1630 6700 1750 6740
rect 1630 6670 1675 6700
rect 1705 6670 1750 6700
rect 1630 6630 1750 6670
rect 1630 6600 1675 6630
rect 1705 6600 1750 6630
rect 1630 6560 1750 6600
rect 1630 6530 1675 6560
rect 1705 6530 1750 6560
rect 1630 6495 1750 6530
rect 1630 6465 1675 6495
rect 1705 6465 1750 6495
rect 1630 6210 1750 6465
rect 2375 9635 2435 9650
rect 2375 9605 2390 9635
rect 2420 9605 2435 9635
rect 2375 9570 2435 9605
rect 2375 9540 2390 9570
rect 2420 9540 2435 9570
rect 2375 9500 2435 9540
rect 2375 9470 2390 9500
rect 2420 9470 2435 9500
rect 2375 9430 2435 9470
rect 2375 9400 2390 9430
rect 2420 9400 2435 9430
rect 2375 9360 2435 9400
rect 2375 9330 2390 9360
rect 2420 9330 2435 9360
rect 2375 9295 2435 9330
rect 2375 9265 2390 9295
rect 2420 9265 2435 9295
rect 2375 9235 2435 9265
rect 2375 9205 2390 9235
rect 2420 9205 2435 9235
rect 2375 9170 2435 9205
rect 2375 9140 2390 9170
rect 2420 9140 2435 9170
rect 2375 9100 2435 9140
rect 2375 9070 2390 9100
rect 2420 9070 2435 9100
rect 2375 9030 2435 9070
rect 2375 9000 2390 9030
rect 2420 9000 2435 9030
rect 2375 8960 2435 9000
rect 2375 8930 2390 8960
rect 2420 8930 2435 8960
rect 2375 8895 2435 8930
rect 2375 8865 2390 8895
rect 2420 8865 2435 8895
rect 2375 8835 2435 8865
rect 2375 8805 2390 8835
rect 2420 8805 2435 8835
rect 2375 8770 2435 8805
rect 2375 8740 2390 8770
rect 2420 8740 2435 8770
rect 2375 8700 2435 8740
rect 2375 8670 2390 8700
rect 2420 8670 2435 8700
rect 2375 8630 2435 8670
rect 2375 8600 2390 8630
rect 2420 8600 2435 8630
rect 2375 8560 2435 8600
rect 2375 8530 2390 8560
rect 2420 8530 2435 8560
rect 2375 8495 2435 8530
rect 2375 8465 2390 8495
rect 2420 8465 2435 8495
rect 2375 8435 2435 8465
rect 2375 8405 2390 8435
rect 2420 8405 2435 8435
rect 2375 8370 2435 8405
rect 2375 8340 2390 8370
rect 2420 8340 2435 8370
rect 2375 8300 2435 8340
rect 2375 8270 2390 8300
rect 2420 8270 2435 8300
rect 2375 8230 2435 8270
rect 2375 8200 2390 8230
rect 2420 8200 2435 8230
rect 2375 8160 2435 8200
rect 2375 8130 2390 8160
rect 2420 8130 2435 8160
rect 2375 8095 2435 8130
rect 2375 8065 2390 8095
rect 2420 8065 2435 8095
rect 2375 8035 2435 8065
rect 2375 8005 2390 8035
rect 2420 8005 2435 8035
rect 2375 7970 2435 8005
rect 2375 7940 2390 7970
rect 2420 7940 2435 7970
rect 2375 7900 2435 7940
rect 2375 7870 2390 7900
rect 2420 7870 2435 7900
rect 2375 7830 2435 7870
rect 2375 7800 2390 7830
rect 2420 7800 2435 7830
rect 2375 7760 2435 7800
rect 2375 7730 2390 7760
rect 2420 7730 2435 7760
rect 2375 7695 2435 7730
rect 2375 7665 2390 7695
rect 2420 7665 2435 7695
rect 2375 7635 2435 7665
rect 2375 7605 2390 7635
rect 2420 7605 2435 7635
rect 2375 7570 2435 7605
rect 2375 7540 2390 7570
rect 2420 7540 2435 7570
rect 2375 7500 2435 7540
rect 2375 7470 2390 7500
rect 2420 7470 2435 7500
rect 2375 7430 2435 7470
rect 2375 7400 2390 7430
rect 2420 7400 2435 7430
rect 2375 7360 2435 7400
rect 2375 7330 2390 7360
rect 2420 7330 2435 7360
rect 2375 7295 2435 7330
rect 2375 7265 2390 7295
rect 2420 7265 2435 7295
rect 2375 7235 2435 7265
rect 2375 7205 2390 7235
rect 2420 7205 2435 7235
rect 2375 7170 2435 7205
rect 2375 7140 2390 7170
rect 2420 7140 2435 7170
rect 2375 7100 2435 7140
rect 2375 7070 2390 7100
rect 2420 7070 2435 7100
rect 2375 7030 2435 7070
rect 2375 7000 2390 7030
rect 2420 7000 2435 7030
rect 2375 6960 2435 7000
rect 2375 6930 2390 6960
rect 2420 6930 2435 6960
rect 2375 6895 2435 6930
rect 2375 6865 2390 6895
rect 2420 6865 2435 6895
rect 2375 6835 2435 6865
rect 2375 6805 2390 6835
rect 2420 6805 2435 6835
rect 2375 6770 2435 6805
rect 2375 6740 2390 6770
rect 2420 6740 2435 6770
rect 2375 6700 2435 6740
rect 2375 6670 2390 6700
rect 2420 6670 2435 6700
rect 2375 6630 2435 6670
rect 2375 6600 2390 6630
rect 2420 6600 2435 6630
rect 2375 6560 2435 6600
rect 2375 6530 2390 6560
rect 2420 6530 2435 6560
rect 2375 6495 2435 6530
rect 2375 6465 2390 6495
rect 2420 6465 2435 6495
rect 2375 6450 2435 6465
rect 2045 6430 2085 6435
rect 2045 6400 2050 6430
rect 2080 6400 2085 6430
rect 2045 6395 2085 6400
rect 2475 6430 2515 9890
rect 2475 6400 2480 6430
rect 2510 6400 2515 6430
rect 2475 6395 2515 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6345 2040 6375
rect 2000 6340 2040 6345
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 1400 6205
rect 1280 6165 1400 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 1400 6165
rect 1280 6125 1400 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 1400 6125
rect 1280 850 1400 6095
rect 2010 1705 2030 6340
rect 2055 1760 2075 6395
rect 2725 6335 2745 9890
rect 2855 6445 2875 9890
rect 2845 6440 2885 6445
rect 2845 6410 2850 6440
rect 2880 6410 2885 6440
rect 2845 6405 2885 6410
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6300 2755 6330
rect 2715 6295 2755 6300
rect 3000 6290 3020 9890
rect 3235 9650 3275 10545
rect 3225 9635 3285 9650
rect 3225 9605 3240 9635
rect 3270 9605 3285 9635
rect 3225 9570 3285 9605
rect 3225 9540 3240 9570
rect 3270 9540 3285 9570
rect 3225 9500 3285 9540
rect 3225 9470 3240 9500
rect 3270 9470 3285 9500
rect 3225 9430 3285 9470
rect 3225 9400 3240 9430
rect 3270 9400 3285 9430
rect 3225 9360 3285 9400
rect 3225 9330 3240 9360
rect 3270 9330 3285 9360
rect 3225 9295 3285 9330
rect 3225 9265 3240 9295
rect 3270 9265 3285 9295
rect 3225 9235 3285 9265
rect 3225 9205 3240 9235
rect 3270 9205 3285 9235
rect 3225 9170 3285 9205
rect 3225 9140 3240 9170
rect 3270 9140 3285 9170
rect 3225 9100 3285 9140
rect 3225 9070 3240 9100
rect 3270 9070 3285 9100
rect 3225 9030 3285 9070
rect 3225 9000 3240 9030
rect 3270 9000 3285 9030
rect 3225 8960 3285 9000
rect 3225 8930 3240 8960
rect 3270 8930 3285 8960
rect 3225 8895 3285 8930
rect 3225 8865 3240 8895
rect 3270 8865 3285 8895
rect 3225 8835 3285 8865
rect 3225 8805 3240 8835
rect 3270 8805 3285 8835
rect 3225 8770 3285 8805
rect 3225 8740 3240 8770
rect 3270 8740 3285 8770
rect 3225 8700 3285 8740
rect 3225 8670 3240 8700
rect 3270 8670 3285 8700
rect 3225 8630 3285 8670
rect 3225 8600 3240 8630
rect 3270 8600 3285 8630
rect 3225 8560 3285 8600
rect 3225 8530 3240 8560
rect 3270 8530 3285 8560
rect 3225 8495 3285 8530
rect 3225 8465 3240 8495
rect 3270 8465 3285 8495
rect 3225 8435 3285 8465
rect 3225 8405 3240 8435
rect 3270 8405 3285 8435
rect 3225 8370 3285 8405
rect 3225 8340 3240 8370
rect 3270 8340 3285 8370
rect 3225 8300 3285 8340
rect 3225 8270 3240 8300
rect 3270 8270 3285 8300
rect 3225 8230 3285 8270
rect 3225 8200 3240 8230
rect 3270 8200 3285 8230
rect 3225 8160 3285 8200
rect 3225 8130 3240 8160
rect 3270 8130 3285 8160
rect 3225 8095 3285 8130
rect 3225 8065 3240 8095
rect 3270 8065 3285 8095
rect 3225 8035 3285 8065
rect 3225 8005 3240 8035
rect 3270 8005 3285 8035
rect 3225 7970 3285 8005
rect 3225 7940 3240 7970
rect 3270 7940 3285 7970
rect 3225 7900 3285 7940
rect 3225 7870 3240 7900
rect 3270 7870 3285 7900
rect 3225 7830 3285 7870
rect 3225 7800 3240 7830
rect 3270 7800 3285 7830
rect 3225 7760 3285 7800
rect 3225 7730 3240 7760
rect 3270 7730 3285 7760
rect 3225 7695 3285 7730
rect 3225 7665 3240 7695
rect 3270 7665 3285 7695
rect 3225 7635 3285 7665
rect 3225 7605 3240 7635
rect 3270 7605 3285 7635
rect 3225 7570 3285 7605
rect 3225 7540 3240 7570
rect 3270 7540 3285 7570
rect 3225 7500 3285 7540
rect 3225 7470 3240 7500
rect 3270 7470 3285 7500
rect 3225 7430 3285 7470
rect 3225 7400 3240 7430
rect 3270 7400 3285 7430
rect 3225 7360 3285 7400
rect 3225 7330 3240 7360
rect 3270 7330 3285 7360
rect 3225 7295 3285 7330
rect 3225 7265 3240 7295
rect 3270 7265 3285 7295
rect 3225 7235 3285 7265
rect 3225 7205 3240 7235
rect 3270 7205 3285 7235
rect 3225 7170 3285 7205
rect 3225 7140 3240 7170
rect 3270 7140 3285 7170
rect 3225 7100 3285 7140
rect 3225 7070 3240 7100
rect 3270 7070 3285 7100
rect 3225 7030 3285 7070
rect 3225 7000 3240 7030
rect 3270 7000 3285 7030
rect 3225 6960 3285 7000
rect 3225 6930 3240 6960
rect 3270 6930 3285 6960
rect 3225 6895 3285 6930
rect 3225 6865 3240 6895
rect 3270 6865 3285 6895
rect 3225 6835 3285 6865
rect 3225 6805 3240 6835
rect 3270 6805 3285 6835
rect 3225 6770 3285 6805
rect 3225 6740 3240 6770
rect 3270 6740 3285 6770
rect 3225 6700 3285 6740
rect 3225 6670 3240 6700
rect 3270 6670 3285 6700
rect 3225 6630 3285 6670
rect 3225 6600 3240 6630
rect 3270 6600 3285 6630
rect 3225 6560 3285 6600
rect 3225 6530 3240 6560
rect 3270 6530 3285 6560
rect 3225 6495 3285 6530
rect 3225 6465 3240 6495
rect 3270 6465 3285 6495
rect 3225 6450 3285 6465
rect 3400 6440 3440 6445
rect 3400 6410 3405 6440
rect 3435 6410 3440 6440
rect 3400 6405 3440 6410
rect 2990 6285 3030 6290
rect 2990 6255 2995 6285
rect 3025 6255 3030 6285
rect 2990 6250 3030 6255
rect 3410 3060 3430 6405
rect 3640 6380 3660 9890
rect 3630 6375 3670 6380
rect 3630 6345 3635 6375
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 3455 6285 3495 6290
rect 3455 6255 3460 6285
rect 3490 6255 3495 6285
rect 3455 6250 3495 6255
rect 3400 3055 3440 3060
rect 3400 3025 3405 3055
rect 3435 3025 3440 3055
rect 3400 3020 3440 3025
rect 3465 2335 3485 6250
rect 4310 6205 4340 10200
rect 4310 6165 4340 6175
rect 4310 6125 4340 6135
rect 4310 6090 4340 6095
rect 4420 6205 4450 10200
rect 4420 6165 4450 6175
rect 4420 6125 4450 6135
rect 4420 6090 4450 6095
rect 4530 6205 4560 10200
rect 4530 6165 4560 6175
rect 4530 6125 4560 6135
rect 4530 6090 4560 6095
rect 4640 6205 4670 10200
rect 5320 6380 5340 9890
rect 5645 9650 5685 10120
rect 5635 9635 5695 9650
rect 5635 9605 5650 9635
rect 5680 9605 5695 9635
rect 5635 9570 5695 9605
rect 5635 9540 5650 9570
rect 5680 9540 5695 9570
rect 5635 9500 5695 9540
rect 5635 9470 5650 9500
rect 5680 9470 5695 9500
rect 5635 9430 5695 9470
rect 5635 9400 5650 9430
rect 5680 9400 5695 9430
rect 5635 9360 5695 9400
rect 5635 9330 5650 9360
rect 5680 9330 5695 9360
rect 5635 9295 5695 9330
rect 5635 9265 5650 9295
rect 5680 9265 5695 9295
rect 5635 9235 5695 9265
rect 5635 9205 5650 9235
rect 5680 9205 5695 9235
rect 5635 9170 5695 9205
rect 5635 9140 5650 9170
rect 5680 9140 5695 9170
rect 5635 9100 5695 9140
rect 5635 9070 5650 9100
rect 5680 9070 5695 9100
rect 5635 9030 5695 9070
rect 5635 9000 5650 9030
rect 5680 9000 5695 9030
rect 5635 8960 5695 9000
rect 5635 8930 5650 8960
rect 5680 8930 5695 8960
rect 5635 8895 5695 8930
rect 5635 8865 5650 8895
rect 5680 8865 5695 8895
rect 5635 8835 5695 8865
rect 5635 8805 5650 8835
rect 5680 8805 5695 8835
rect 5635 8770 5695 8805
rect 5635 8740 5650 8770
rect 5680 8740 5695 8770
rect 5635 8700 5695 8740
rect 5635 8670 5650 8700
rect 5680 8670 5695 8700
rect 5635 8630 5695 8670
rect 5635 8600 5650 8630
rect 5680 8600 5695 8630
rect 5635 8560 5695 8600
rect 5635 8530 5650 8560
rect 5680 8530 5695 8560
rect 5635 8495 5695 8530
rect 5635 8465 5650 8495
rect 5680 8465 5695 8495
rect 5635 8435 5695 8465
rect 5635 8405 5650 8435
rect 5680 8405 5695 8435
rect 5635 8370 5695 8405
rect 5635 8340 5650 8370
rect 5680 8340 5695 8370
rect 5635 8300 5695 8340
rect 5635 8270 5650 8300
rect 5680 8270 5695 8300
rect 5635 8230 5695 8270
rect 5635 8200 5650 8230
rect 5680 8200 5695 8230
rect 5635 8160 5695 8200
rect 5635 8130 5650 8160
rect 5680 8130 5695 8160
rect 5635 8095 5695 8130
rect 5635 8065 5650 8095
rect 5680 8065 5695 8095
rect 5635 8035 5695 8065
rect 5635 8005 5650 8035
rect 5680 8005 5695 8035
rect 5635 7970 5695 8005
rect 5635 7940 5650 7970
rect 5680 7940 5695 7970
rect 5635 7900 5695 7940
rect 5635 7870 5650 7900
rect 5680 7870 5695 7900
rect 5635 7830 5695 7870
rect 5635 7800 5650 7830
rect 5680 7800 5695 7830
rect 5635 7760 5695 7800
rect 5635 7730 5650 7760
rect 5680 7730 5695 7760
rect 5635 7695 5695 7730
rect 5635 7665 5650 7695
rect 5680 7665 5695 7695
rect 5635 7635 5695 7665
rect 5635 7605 5650 7635
rect 5680 7605 5695 7635
rect 5635 7570 5695 7605
rect 5635 7540 5650 7570
rect 5680 7540 5695 7570
rect 5635 7500 5695 7540
rect 5635 7470 5650 7500
rect 5680 7470 5695 7500
rect 5635 7430 5695 7470
rect 5635 7400 5650 7430
rect 5680 7400 5695 7430
rect 5635 7360 5695 7400
rect 5635 7330 5650 7360
rect 5680 7330 5695 7360
rect 5635 7295 5695 7330
rect 5635 7265 5650 7295
rect 5680 7265 5695 7295
rect 5635 7235 5695 7265
rect 5635 7205 5650 7235
rect 5680 7205 5695 7235
rect 5635 7170 5695 7205
rect 5635 7140 5650 7170
rect 5680 7140 5695 7170
rect 5635 7100 5695 7140
rect 5635 7070 5650 7100
rect 5680 7070 5695 7100
rect 5635 7030 5695 7070
rect 5635 7000 5650 7030
rect 5680 7000 5695 7030
rect 5635 6960 5695 7000
rect 5635 6930 5650 6960
rect 5680 6930 5695 6960
rect 5635 6895 5695 6930
rect 5635 6865 5650 6895
rect 5680 6865 5695 6895
rect 5635 6835 5695 6865
rect 5635 6805 5650 6835
rect 5680 6805 5695 6835
rect 5635 6770 5695 6805
rect 5635 6740 5650 6770
rect 5680 6740 5695 6770
rect 5635 6700 5695 6740
rect 5635 6670 5650 6700
rect 5680 6670 5695 6700
rect 5635 6630 5695 6670
rect 5635 6600 5650 6630
rect 5680 6600 5695 6630
rect 5635 6560 5695 6600
rect 5635 6530 5650 6560
rect 5680 6530 5695 6560
rect 5635 6495 5695 6530
rect 5635 6465 5650 6495
rect 5680 6465 5695 6495
rect 5635 6450 5695 6465
rect 6155 6435 6175 9890
rect 5490 6430 5530 6435
rect 5490 6400 5495 6430
rect 5525 6400 5530 6430
rect 5490 6395 5530 6400
rect 6145 6430 6185 6435
rect 6145 6400 6150 6430
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6345 5350 6375
rect 5310 6340 5350 6345
rect 4850 6330 4890 6335
rect 4850 6300 4855 6330
rect 4885 6300 4890 6330
rect 4850 6295 4890 6300
rect 4640 6165 4670 6175
rect 4640 6125 4670 6135
rect 4640 6090 4670 6095
rect 4860 5020 4880 6295
rect 4850 5015 4890 5020
rect 4850 4985 4855 5015
rect 4885 4985 4890 5015
rect 4850 4980 4890 4985
rect 4940 5015 4980 5020
rect 4940 4985 4945 5015
rect 4975 4985 4980 5015
rect 4940 4980 4980 4985
rect 4950 4505 4970 4980
rect 5166 4555 5196 4560
rect 5166 4520 5196 4525
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 5500 3125 5520 6395
rect 6230 5140 6250 9890
rect 6300 9650 6340 11375
rect 6290 9635 6350 9650
rect 6290 9605 6305 9635
rect 6335 9605 6350 9635
rect 6290 9570 6350 9605
rect 6290 9540 6305 9570
rect 6335 9540 6350 9570
rect 6290 9500 6350 9540
rect 6290 9470 6305 9500
rect 6335 9470 6350 9500
rect 6290 9430 6350 9470
rect 6290 9400 6305 9430
rect 6335 9400 6350 9430
rect 6290 9360 6350 9400
rect 6290 9330 6305 9360
rect 6335 9330 6350 9360
rect 6290 9295 6350 9330
rect 6290 9265 6305 9295
rect 6335 9265 6350 9295
rect 6290 9235 6350 9265
rect 6290 9205 6305 9235
rect 6335 9205 6350 9235
rect 6290 9170 6350 9205
rect 6290 9140 6305 9170
rect 6335 9140 6350 9170
rect 6290 9100 6350 9140
rect 6290 9070 6305 9100
rect 6335 9070 6350 9100
rect 6290 9030 6350 9070
rect 6290 9000 6305 9030
rect 6335 9000 6350 9030
rect 6290 8960 6350 9000
rect 6290 8930 6305 8960
rect 6335 8930 6350 8960
rect 6290 8895 6350 8930
rect 6290 8865 6305 8895
rect 6335 8865 6350 8895
rect 6290 8835 6350 8865
rect 6290 8805 6305 8835
rect 6335 8805 6350 8835
rect 6290 8770 6350 8805
rect 6290 8740 6305 8770
rect 6335 8740 6350 8770
rect 6290 8700 6350 8740
rect 6290 8670 6305 8700
rect 6335 8670 6350 8700
rect 6290 8630 6350 8670
rect 6290 8600 6305 8630
rect 6335 8600 6350 8630
rect 6290 8560 6350 8600
rect 6290 8530 6305 8560
rect 6335 8530 6350 8560
rect 6290 8495 6350 8530
rect 6290 8465 6305 8495
rect 6335 8465 6350 8495
rect 6290 8435 6350 8465
rect 6290 8405 6305 8435
rect 6335 8405 6350 8435
rect 6290 8370 6350 8405
rect 6290 8340 6305 8370
rect 6335 8340 6350 8370
rect 6290 8300 6350 8340
rect 6290 8270 6305 8300
rect 6335 8270 6350 8300
rect 6290 8230 6350 8270
rect 6290 8200 6305 8230
rect 6335 8200 6350 8230
rect 6290 8160 6350 8200
rect 6290 8130 6305 8160
rect 6335 8130 6350 8160
rect 6290 8095 6350 8130
rect 6290 8065 6305 8095
rect 6335 8065 6350 8095
rect 6290 8035 6350 8065
rect 6290 8005 6305 8035
rect 6335 8005 6350 8035
rect 6290 7970 6350 8005
rect 6290 7940 6305 7970
rect 6335 7940 6350 7970
rect 6290 7900 6350 7940
rect 6290 7870 6305 7900
rect 6335 7870 6350 7900
rect 6290 7830 6350 7870
rect 6290 7800 6305 7830
rect 6335 7800 6350 7830
rect 6290 7760 6350 7800
rect 6290 7730 6305 7760
rect 6335 7730 6350 7760
rect 6290 7695 6350 7730
rect 6290 7665 6305 7695
rect 6335 7665 6350 7695
rect 6290 7635 6350 7665
rect 6290 7605 6305 7635
rect 6335 7605 6350 7635
rect 6290 7570 6350 7605
rect 6290 7540 6305 7570
rect 6335 7540 6350 7570
rect 6290 7500 6350 7540
rect 6290 7470 6305 7500
rect 6335 7470 6350 7500
rect 6290 7430 6350 7470
rect 6290 7400 6305 7430
rect 6335 7400 6350 7430
rect 6290 7360 6350 7400
rect 6290 7330 6305 7360
rect 6335 7330 6350 7360
rect 6290 7295 6350 7330
rect 6290 7265 6305 7295
rect 6335 7265 6350 7295
rect 6290 7235 6350 7265
rect 6290 7205 6305 7235
rect 6335 7205 6350 7235
rect 6290 7170 6350 7205
rect 6290 7140 6305 7170
rect 6335 7140 6350 7170
rect 6290 7100 6350 7140
rect 6290 7070 6305 7100
rect 6335 7070 6350 7100
rect 6290 7030 6350 7070
rect 6290 7000 6305 7030
rect 6335 7000 6350 7030
rect 6290 6960 6350 7000
rect 6290 6930 6305 6960
rect 6335 6930 6350 6960
rect 6290 6895 6350 6930
rect 6290 6865 6305 6895
rect 6335 6865 6350 6895
rect 6290 6835 6350 6865
rect 6290 6805 6305 6835
rect 6335 6805 6350 6835
rect 6290 6770 6350 6805
rect 6290 6740 6305 6770
rect 6335 6740 6350 6770
rect 6290 6700 6350 6740
rect 6290 6670 6305 6700
rect 6335 6670 6350 6700
rect 6290 6630 6350 6670
rect 6290 6600 6305 6630
rect 6335 6600 6350 6630
rect 6290 6560 6350 6600
rect 6290 6530 6305 6560
rect 6335 6530 6350 6560
rect 6290 6495 6350 6530
rect 6290 6465 6305 6495
rect 6335 6465 6350 6495
rect 6290 6450 6350 6465
rect 6465 6430 6505 9890
rect 6590 9650 6630 12090
rect 6580 9635 6640 9650
rect 6580 9605 6595 9635
rect 6625 9605 6640 9635
rect 6580 9570 6640 9605
rect 6580 9540 6595 9570
rect 6625 9540 6640 9570
rect 6580 9500 6640 9540
rect 6580 9470 6595 9500
rect 6625 9470 6640 9500
rect 6580 9430 6640 9470
rect 6580 9400 6595 9430
rect 6625 9400 6640 9430
rect 6580 9360 6640 9400
rect 6580 9330 6595 9360
rect 6625 9330 6640 9360
rect 6580 9295 6640 9330
rect 6580 9265 6595 9295
rect 6625 9265 6640 9295
rect 6580 9235 6640 9265
rect 6580 9205 6595 9235
rect 6625 9205 6640 9235
rect 6580 9170 6640 9205
rect 6580 9140 6595 9170
rect 6625 9140 6640 9170
rect 6580 9100 6640 9140
rect 6580 9070 6595 9100
rect 6625 9070 6640 9100
rect 6580 9030 6640 9070
rect 6580 9000 6595 9030
rect 6625 9000 6640 9030
rect 6580 8960 6640 9000
rect 6580 8930 6595 8960
rect 6625 8930 6640 8960
rect 6580 8895 6640 8930
rect 6580 8865 6595 8895
rect 6625 8865 6640 8895
rect 6580 8835 6640 8865
rect 6580 8805 6595 8835
rect 6625 8805 6640 8835
rect 6580 8770 6640 8805
rect 6580 8740 6595 8770
rect 6625 8740 6640 8770
rect 6580 8700 6640 8740
rect 6580 8670 6595 8700
rect 6625 8670 6640 8700
rect 6580 8630 6640 8670
rect 6580 8600 6595 8630
rect 6625 8600 6640 8630
rect 6580 8560 6640 8600
rect 6580 8530 6595 8560
rect 6625 8530 6640 8560
rect 6580 8495 6640 8530
rect 6580 8465 6595 8495
rect 6625 8465 6640 8495
rect 6580 8435 6640 8465
rect 6580 8405 6595 8435
rect 6625 8405 6640 8435
rect 6580 8370 6640 8405
rect 6580 8340 6595 8370
rect 6625 8340 6640 8370
rect 6580 8300 6640 8340
rect 6580 8270 6595 8300
rect 6625 8270 6640 8300
rect 6580 8230 6640 8270
rect 6580 8200 6595 8230
rect 6625 8200 6640 8230
rect 6580 8160 6640 8200
rect 6580 8130 6595 8160
rect 6625 8130 6640 8160
rect 6580 8095 6640 8130
rect 6580 8065 6595 8095
rect 6625 8065 6640 8095
rect 6580 8035 6640 8065
rect 6580 8005 6595 8035
rect 6625 8005 6640 8035
rect 6580 7970 6640 8005
rect 6580 7940 6595 7970
rect 6625 7940 6640 7970
rect 6580 7900 6640 7940
rect 6580 7870 6595 7900
rect 6625 7870 6640 7900
rect 6580 7830 6640 7870
rect 6580 7800 6595 7830
rect 6625 7800 6640 7830
rect 6580 7760 6640 7800
rect 6580 7730 6595 7760
rect 6625 7730 6640 7760
rect 6580 7695 6640 7730
rect 6580 7665 6595 7695
rect 6625 7665 6640 7695
rect 6580 7635 6640 7665
rect 6580 7605 6595 7635
rect 6625 7605 6640 7635
rect 6580 7570 6640 7605
rect 6580 7540 6595 7570
rect 6625 7540 6640 7570
rect 6580 7500 6640 7540
rect 6580 7470 6595 7500
rect 6625 7470 6640 7500
rect 6580 7430 6640 7470
rect 6580 7400 6595 7430
rect 6625 7400 6640 7430
rect 6580 7360 6640 7400
rect 6580 7330 6595 7360
rect 6625 7330 6640 7360
rect 6580 7295 6640 7330
rect 6580 7265 6595 7295
rect 6625 7265 6640 7295
rect 6580 7235 6640 7265
rect 6580 7205 6595 7235
rect 6625 7205 6640 7235
rect 6580 7170 6640 7205
rect 6580 7140 6595 7170
rect 6625 7140 6640 7170
rect 6580 7100 6640 7140
rect 6580 7070 6595 7100
rect 6625 7070 6640 7100
rect 6580 7030 6640 7070
rect 6580 7000 6595 7030
rect 6625 7000 6640 7030
rect 6580 6960 6640 7000
rect 6580 6930 6595 6960
rect 6625 6930 6640 6960
rect 6580 6895 6640 6930
rect 6580 6865 6595 6895
rect 6625 6865 6640 6895
rect 6580 6835 6640 6865
rect 6580 6805 6595 6835
rect 6625 6805 6640 6835
rect 6580 6770 6640 6805
rect 6580 6740 6595 6770
rect 6625 6740 6640 6770
rect 6580 6700 6640 6740
rect 6580 6670 6595 6700
rect 6625 6670 6640 6700
rect 6580 6630 6640 6670
rect 6580 6600 6595 6630
rect 6625 6600 6640 6630
rect 6580 6560 6640 6600
rect 6580 6530 6595 6560
rect 6625 6530 6640 6560
rect 6580 6495 6640 6530
rect 6580 6465 6595 6495
rect 6625 6465 6640 6495
rect 6580 6450 6640 6465
rect 7230 9635 7350 9650
rect 7230 9605 7275 9635
rect 7305 9605 7350 9635
rect 7230 9570 7350 9605
rect 7230 9540 7275 9570
rect 7305 9540 7350 9570
rect 7230 9500 7350 9540
rect 7230 9470 7275 9500
rect 7305 9470 7350 9500
rect 7230 9430 7350 9470
rect 7230 9400 7275 9430
rect 7305 9400 7350 9430
rect 7230 9360 7350 9400
rect 7230 9330 7275 9360
rect 7305 9330 7350 9360
rect 7230 9295 7350 9330
rect 7230 9265 7275 9295
rect 7305 9265 7350 9295
rect 7230 9235 7350 9265
rect 7230 9205 7275 9235
rect 7305 9205 7350 9235
rect 7230 9170 7350 9205
rect 7230 9140 7275 9170
rect 7305 9140 7350 9170
rect 7230 9100 7350 9140
rect 7230 9070 7275 9100
rect 7305 9070 7350 9100
rect 7230 9030 7350 9070
rect 7230 9000 7275 9030
rect 7305 9000 7350 9030
rect 7230 8960 7350 9000
rect 7230 8930 7275 8960
rect 7305 8930 7350 8960
rect 7230 8895 7350 8930
rect 7230 8865 7275 8895
rect 7305 8865 7350 8895
rect 7230 8835 7350 8865
rect 7230 8805 7275 8835
rect 7305 8805 7350 8835
rect 7230 8770 7350 8805
rect 7230 8740 7275 8770
rect 7305 8740 7350 8770
rect 7230 8700 7350 8740
rect 7230 8670 7275 8700
rect 7305 8670 7350 8700
rect 7230 8630 7350 8670
rect 7230 8600 7275 8630
rect 7305 8600 7350 8630
rect 7230 8560 7350 8600
rect 7230 8530 7275 8560
rect 7305 8530 7350 8560
rect 7230 8495 7350 8530
rect 7230 8465 7275 8495
rect 7305 8465 7350 8495
rect 7230 8435 7350 8465
rect 7230 8405 7275 8435
rect 7305 8405 7350 8435
rect 7230 8370 7350 8405
rect 7230 8340 7275 8370
rect 7305 8340 7350 8370
rect 7230 8300 7350 8340
rect 7230 8270 7275 8300
rect 7305 8270 7350 8300
rect 7230 8230 7350 8270
rect 7230 8200 7275 8230
rect 7305 8200 7350 8230
rect 7230 8160 7350 8200
rect 7230 8130 7275 8160
rect 7305 8130 7350 8160
rect 7230 8095 7350 8130
rect 7230 8065 7275 8095
rect 7305 8065 7350 8095
rect 7230 8035 7350 8065
rect 7230 8005 7275 8035
rect 7305 8005 7350 8035
rect 7230 7970 7350 8005
rect 7230 7940 7275 7970
rect 7305 7940 7350 7970
rect 7230 7900 7350 7940
rect 7230 7870 7275 7900
rect 7305 7870 7350 7900
rect 7230 7830 7350 7870
rect 7230 7800 7275 7830
rect 7305 7800 7350 7830
rect 7230 7760 7350 7800
rect 7230 7730 7275 7760
rect 7305 7730 7350 7760
rect 7230 7695 7350 7730
rect 7230 7665 7275 7695
rect 7305 7665 7350 7695
rect 7230 7635 7350 7665
rect 7230 7605 7275 7635
rect 7305 7605 7350 7635
rect 7230 7570 7350 7605
rect 7230 7540 7275 7570
rect 7305 7540 7350 7570
rect 7230 7500 7350 7540
rect 7230 7470 7275 7500
rect 7305 7470 7350 7500
rect 7230 7430 7350 7470
rect 7230 7400 7275 7430
rect 7305 7400 7350 7430
rect 7230 7360 7350 7400
rect 7230 7330 7275 7360
rect 7305 7330 7350 7360
rect 7230 7295 7350 7330
rect 7230 7265 7275 7295
rect 7305 7265 7350 7295
rect 7230 7235 7350 7265
rect 7230 7205 7275 7235
rect 7305 7205 7350 7235
rect 7230 7170 7350 7205
rect 7230 7140 7275 7170
rect 7305 7140 7350 7170
rect 7230 7100 7350 7140
rect 7230 7070 7275 7100
rect 7305 7070 7350 7100
rect 7230 7030 7350 7070
rect 7230 7000 7275 7030
rect 7305 7000 7350 7030
rect 7230 6960 7350 7000
rect 7230 6930 7275 6960
rect 7305 6930 7350 6960
rect 7230 6895 7350 6930
rect 7230 6865 7275 6895
rect 7305 6865 7350 6895
rect 7230 6835 7350 6865
rect 7230 6805 7275 6835
rect 7305 6805 7350 6835
rect 7230 6770 7350 6805
rect 7230 6740 7275 6770
rect 7305 6740 7350 6770
rect 7230 6700 7350 6740
rect 7230 6670 7275 6700
rect 7305 6670 7350 6700
rect 7230 6630 7350 6670
rect 7230 6600 7275 6630
rect 7305 6600 7350 6630
rect 7230 6560 7350 6600
rect 7230 6530 7275 6560
rect 7305 6530 7350 6560
rect 7230 6495 7350 6530
rect 7230 6465 7275 6495
rect 7305 6465 7350 6495
rect 6465 6400 6470 6430
rect 6500 6400 6505 6430
rect 6465 6395 6505 6400
rect 6895 6430 6935 6435
rect 6895 6400 6900 6430
rect 6930 6400 6935 6430
rect 6895 6395 6935 6400
rect 5870 5135 5910 5140
rect 5870 5105 5875 5135
rect 5905 5105 5910 5135
rect 5870 5100 5910 5105
rect 6220 5135 6260 5140
rect 6220 5105 6225 5135
rect 6255 5105 6260 5135
rect 6220 5100 6260 5105
rect 5880 4570 5900 5100
rect 5870 4565 5910 4570
rect 5870 4535 5875 4565
rect 5905 4535 5910 4565
rect 5870 4530 5910 4535
rect 5490 3120 5530 3125
rect 5490 3090 5495 3120
rect 5525 3090 5530 3120
rect 5490 3085 5530 3090
rect 6905 1760 6925 6395
rect 6940 6375 6980 6380
rect 6940 6345 6945 6375
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2045 1755 2085 1760
rect 2045 1725 2050 1755
rect 2080 1725 2085 1755
rect 2045 1720 2085 1725
rect 2175 1755 2215 1760
rect 2175 1725 2180 1755
rect 2210 1725 2215 1755
rect 2175 1720 2215 1725
rect 6765 1755 6805 1760
rect 6765 1725 6770 1755
rect 6800 1725 6805 1755
rect 6765 1720 6805 1725
rect 6895 1755 6935 1760
rect 6895 1725 6900 1755
rect 6930 1725 6935 1755
rect 6895 1720 6935 1725
rect 2000 1700 2040 1705
rect 2000 1670 2005 1700
rect 2035 1670 2040 1700
rect 2000 1665 2040 1670
rect 2100 1700 2140 1705
rect 2100 1670 2105 1700
rect 2135 1670 2140 1700
rect 2100 1665 2140 1670
rect 2110 1515 2130 1665
rect 2185 1330 2205 1720
rect 6775 1330 6795 1720
rect 6950 1705 6970 6340
rect 7230 6210 7350 6465
rect 7580 9635 7700 9650
rect 7580 9605 7625 9635
rect 7655 9605 7700 9635
rect 7580 9570 7700 9605
rect 7580 9540 7625 9570
rect 7655 9540 7700 9570
rect 7580 9500 7700 9540
rect 7580 9470 7625 9500
rect 7655 9470 7700 9500
rect 7580 9430 7700 9470
rect 7580 9400 7625 9430
rect 7655 9400 7700 9430
rect 7580 9360 7700 9400
rect 7580 9330 7625 9360
rect 7655 9330 7700 9360
rect 7580 9295 7700 9330
rect 7580 9265 7625 9295
rect 7655 9265 7700 9295
rect 7580 9235 7700 9265
rect 7580 9205 7625 9235
rect 7655 9205 7700 9235
rect 7580 9170 7700 9205
rect 7580 9140 7625 9170
rect 7655 9140 7700 9170
rect 7580 9100 7700 9140
rect 7580 9070 7625 9100
rect 7655 9070 7700 9100
rect 7580 9030 7700 9070
rect 7580 9000 7625 9030
rect 7655 9000 7700 9030
rect 7580 8960 7700 9000
rect 7580 8930 7625 8960
rect 7655 8930 7700 8960
rect 7580 8895 7700 8930
rect 7580 8865 7625 8895
rect 7655 8865 7700 8895
rect 7580 8835 7700 8865
rect 7580 8805 7625 8835
rect 7655 8805 7700 8835
rect 7580 8770 7700 8805
rect 7580 8740 7625 8770
rect 7655 8740 7700 8770
rect 7580 8700 7700 8740
rect 7580 8670 7625 8700
rect 7655 8670 7700 8700
rect 7580 8630 7700 8670
rect 7580 8600 7625 8630
rect 7655 8600 7700 8630
rect 7580 8560 7700 8600
rect 7580 8530 7625 8560
rect 7655 8530 7700 8560
rect 7580 8495 7700 8530
rect 7580 8465 7625 8495
rect 7655 8465 7700 8495
rect 7580 8435 7700 8465
rect 7580 8405 7625 8435
rect 7655 8405 7700 8435
rect 7580 8370 7700 8405
rect 7580 8340 7625 8370
rect 7655 8340 7700 8370
rect 7580 8300 7700 8340
rect 7580 8270 7625 8300
rect 7655 8270 7700 8300
rect 7580 8230 7700 8270
rect 7580 8200 7625 8230
rect 7655 8200 7700 8230
rect 7580 8160 7700 8200
rect 7580 8130 7625 8160
rect 7655 8130 7700 8160
rect 7580 8095 7700 8130
rect 7580 8065 7625 8095
rect 7655 8065 7700 8095
rect 7580 8035 7700 8065
rect 7580 8005 7625 8035
rect 7655 8005 7700 8035
rect 7580 7970 7700 8005
rect 7580 7940 7625 7970
rect 7655 7940 7700 7970
rect 7580 7900 7700 7940
rect 7580 7870 7625 7900
rect 7655 7870 7700 7900
rect 7580 7830 7700 7870
rect 7580 7800 7625 7830
rect 7655 7800 7700 7830
rect 7580 7760 7700 7800
rect 7580 7730 7625 7760
rect 7655 7730 7700 7760
rect 7580 7695 7700 7730
rect 7580 7665 7625 7695
rect 7655 7665 7700 7695
rect 7580 7635 7700 7665
rect 7580 7605 7625 7635
rect 7655 7605 7700 7635
rect 7580 7570 7700 7605
rect 7580 7540 7625 7570
rect 7655 7540 7700 7570
rect 7580 7500 7700 7540
rect 7580 7470 7625 7500
rect 7655 7470 7700 7500
rect 7580 7430 7700 7470
rect 7580 7400 7625 7430
rect 7655 7400 7700 7430
rect 7580 7360 7700 7400
rect 7580 7330 7625 7360
rect 7655 7330 7700 7360
rect 7580 7295 7700 7330
rect 7580 7265 7625 7295
rect 7655 7265 7700 7295
rect 7580 7235 7700 7265
rect 7580 7205 7625 7235
rect 7655 7205 7700 7235
rect 7580 7170 7700 7205
rect 7580 7140 7625 7170
rect 7655 7140 7700 7170
rect 7580 7100 7700 7140
rect 7580 7070 7625 7100
rect 7655 7070 7700 7100
rect 7580 7030 7700 7070
rect 7580 7000 7625 7030
rect 7655 7000 7700 7030
rect 7580 6960 7700 7000
rect 7580 6930 7625 6960
rect 7655 6930 7700 6960
rect 7580 6895 7700 6930
rect 7580 6865 7625 6895
rect 7655 6865 7700 6895
rect 7580 6835 7700 6865
rect 7580 6805 7625 6835
rect 7655 6805 7700 6835
rect 7580 6770 7700 6805
rect 7580 6740 7625 6770
rect 7655 6740 7700 6770
rect 7580 6700 7700 6740
rect 7580 6670 7625 6700
rect 7655 6670 7700 6700
rect 7580 6630 7700 6670
rect 7580 6600 7625 6630
rect 7655 6600 7700 6630
rect 7580 6560 7700 6600
rect 7580 6530 7625 6560
rect 7655 6530 7700 6560
rect 7580 6495 7700 6530
rect 7580 6465 7625 6495
rect 7655 6465 7700 6495
rect 7580 6205 7700 6465
rect 8280 9635 8400 9650
rect 8280 9605 8325 9635
rect 8355 9605 8400 9635
rect 8280 9570 8400 9605
rect 8280 9540 8325 9570
rect 8355 9540 8400 9570
rect 8280 9500 8400 9540
rect 8280 9470 8325 9500
rect 8355 9470 8400 9500
rect 8280 9430 8400 9470
rect 8280 9400 8325 9430
rect 8355 9400 8400 9430
rect 8280 9360 8400 9400
rect 8280 9330 8325 9360
rect 8355 9330 8400 9360
rect 8280 9295 8400 9330
rect 8280 9265 8325 9295
rect 8355 9265 8400 9295
rect 8280 9235 8400 9265
rect 8280 9205 8325 9235
rect 8355 9205 8400 9235
rect 8280 9170 8400 9205
rect 8280 9140 8325 9170
rect 8355 9140 8400 9170
rect 8280 9100 8400 9140
rect 8280 9070 8325 9100
rect 8355 9070 8400 9100
rect 8280 9030 8400 9070
rect 8280 9000 8325 9030
rect 8355 9000 8400 9030
rect 8280 8960 8400 9000
rect 8280 8930 8325 8960
rect 8355 8930 8400 8960
rect 8280 8895 8400 8930
rect 8280 8865 8325 8895
rect 8355 8865 8400 8895
rect 8280 8835 8400 8865
rect 8280 8805 8325 8835
rect 8355 8805 8400 8835
rect 8280 8770 8400 8805
rect 8280 8740 8325 8770
rect 8355 8740 8400 8770
rect 8280 8700 8400 8740
rect 8280 8670 8325 8700
rect 8355 8670 8400 8700
rect 8280 8630 8400 8670
rect 8280 8600 8325 8630
rect 8355 8600 8400 8630
rect 8280 8560 8400 8600
rect 8280 8530 8325 8560
rect 8355 8530 8400 8560
rect 8280 8495 8400 8530
rect 8280 8465 8325 8495
rect 8355 8465 8400 8495
rect 8280 8435 8400 8465
rect 8280 8405 8325 8435
rect 8355 8405 8400 8435
rect 8280 8370 8400 8405
rect 8280 8340 8325 8370
rect 8355 8340 8400 8370
rect 8280 8300 8400 8340
rect 8280 8270 8325 8300
rect 8355 8270 8400 8300
rect 8280 8230 8400 8270
rect 8280 8200 8325 8230
rect 8355 8200 8400 8230
rect 8280 8160 8400 8200
rect 8280 8130 8325 8160
rect 8355 8130 8400 8160
rect 8280 8095 8400 8130
rect 8280 8065 8325 8095
rect 8355 8065 8400 8095
rect 8280 8035 8400 8065
rect 8280 8005 8325 8035
rect 8355 8005 8400 8035
rect 8280 7970 8400 8005
rect 8280 7940 8325 7970
rect 8355 7940 8400 7970
rect 8280 7900 8400 7940
rect 8280 7870 8325 7900
rect 8355 7870 8400 7900
rect 8280 7830 8400 7870
rect 8280 7800 8325 7830
rect 8355 7800 8400 7830
rect 8280 7760 8400 7800
rect 8280 7730 8325 7760
rect 8355 7730 8400 7760
rect 8280 7695 8400 7730
rect 8280 7665 8325 7695
rect 8355 7665 8400 7695
rect 8280 7635 8400 7665
rect 8280 7605 8325 7635
rect 8355 7605 8400 7635
rect 8280 7570 8400 7605
rect 8280 7540 8325 7570
rect 8355 7540 8400 7570
rect 8280 7500 8400 7540
rect 8280 7470 8325 7500
rect 8355 7470 8400 7500
rect 8280 7430 8400 7470
rect 8280 7400 8325 7430
rect 8355 7400 8400 7430
rect 8280 7360 8400 7400
rect 8280 7330 8325 7360
rect 8355 7330 8400 7360
rect 8280 7295 8400 7330
rect 8280 7265 8325 7295
rect 8355 7265 8400 7295
rect 8280 7235 8400 7265
rect 8280 7205 8325 7235
rect 8355 7205 8400 7235
rect 8280 7170 8400 7205
rect 8280 7140 8325 7170
rect 8355 7140 8400 7170
rect 8280 7100 8400 7140
rect 8280 7070 8325 7100
rect 8355 7070 8400 7100
rect 8280 7030 8400 7070
rect 8280 7000 8325 7030
rect 8355 7000 8400 7030
rect 8280 6960 8400 7000
rect 8280 6930 8325 6960
rect 8355 6930 8400 6960
rect 8280 6895 8400 6930
rect 8280 6865 8325 6895
rect 8355 6865 8400 6895
rect 8280 6835 8400 6865
rect 8280 6805 8325 6835
rect 8355 6805 8400 6835
rect 8280 6770 8400 6805
rect 8280 6740 8325 6770
rect 8355 6740 8400 6770
rect 8280 6700 8400 6740
rect 8280 6670 8325 6700
rect 8355 6670 8400 6700
rect 8280 6630 8400 6670
rect 8280 6600 8325 6630
rect 8355 6600 8400 6630
rect 8280 6560 8400 6600
rect 8280 6530 8325 6560
rect 8355 6530 8400 6560
rect 8280 6495 8400 6530
rect 8280 6465 8325 6495
rect 8355 6465 8400 6495
rect 8280 6210 8400 6465
rect 8630 9635 8750 9650
rect 8630 9605 8675 9635
rect 8705 9605 8750 9635
rect 8630 9570 8750 9605
rect 8630 9540 8675 9570
rect 8705 9540 8750 9570
rect 8630 9500 8750 9540
rect 8630 9470 8675 9500
rect 8705 9470 8750 9500
rect 8630 9430 8750 9470
rect 8630 9400 8675 9430
rect 8705 9400 8750 9430
rect 8630 9360 8750 9400
rect 8630 9330 8675 9360
rect 8705 9330 8750 9360
rect 8630 9295 8750 9330
rect 8630 9265 8675 9295
rect 8705 9265 8750 9295
rect 8630 9235 8750 9265
rect 8630 9205 8675 9235
rect 8705 9205 8750 9235
rect 8630 9170 8750 9205
rect 8630 9140 8675 9170
rect 8705 9140 8750 9170
rect 8630 9100 8750 9140
rect 8630 9070 8675 9100
rect 8705 9070 8750 9100
rect 8630 9030 8750 9070
rect 8630 9000 8675 9030
rect 8705 9000 8750 9030
rect 8630 8960 8750 9000
rect 8630 8930 8675 8960
rect 8705 8930 8750 8960
rect 8630 8895 8750 8930
rect 8630 8865 8675 8895
rect 8705 8865 8750 8895
rect 8630 8835 8750 8865
rect 8630 8805 8675 8835
rect 8705 8805 8750 8835
rect 8630 8770 8750 8805
rect 8630 8740 8675 8770
rect 8705 8740 8750 8770
rect 8630 8700 8750 8740
rect 8630 8670 8675 8700
rect 8705 8670 8750 8700
rect 8630 8630 8750 8670
rect 8630 8600 8675 8630
rect 8705 8600 8750 8630
rect 8630 8560 8750 8600
rect 8630 8530 8675 8560
rect 8705 8530 8750 8560
rect 8630 8495 8750 8530
rect 8630 8465 8675 8495
rect 8705 8465 8750 8495
rect 8630 8435 8750 8465
rect 8630 8405 8675 8435
rect 8705 8405 8750 8435
rect 8630 8370 8750 8405
rect 8630 8340 8675 8370
rect 8705 8340 8750 8370
rect 8630 8300 8750 8340
rect 8630 8270 8675 8300
rect 8705 8270 8750 8300
rect 8630 8230 8750 8270
rect 8630 8200 8675 8230
rect 8705 8200 8750 8230
rect 8630 8160 8750 8200
rect 8630 8130 8675 8160
rect 8705 8130 8750 8160
rect 8630 8095 8750 8130
rect 8630 8065 8675 8095
rect 8705 8065 8750 8095
rect 8630 8035 8750 8065
rect 8630 8005 8675 8035
rect 8705 8005 8750 8035
rect 8630 7970 8750 8005
rect 8630 7940 8675 7970
rect 8705 7940 8750 7970
rect 8630 7900 8750 7940
rect 8630 7870 8675 7900
rect 8705 7870 8750 7900
rect 8630 7830 8750 7870
rect 8630 7800 8675 7830
rect 8705 7800 8750 7830
rect 8630 7760 8750 7800
rect 8630 7730 8675 7760
rect 8705 7730 8750 7760
rect 8630 7695 8750 7730
rect 8630 7665 8675 7695
rect 8705 7665 8750 7695
rect 8630 7635 8750 7665
rect 8630 7605 8675 7635
rect 8705 7605 8750 7635
rect 8630 7570 8750 7605
rect 8630 7540 8675 7570
rect 8705 7540 8750 7570
rect 8630 7500 8750 7540
rect 8630 7470 8675 7500
rect 8705 7470 8750 7500
rect 8630 7430 8750 7470
rect 8630 7400 8675 7430
rect 8705 7400 8750 7430
rect 8630 7360 8750 7400
rect 8630 7330 8675 7360
rect 8705 7330 8750 7360
rect 8630 7295 8750 7330
rect 8630 7265 8675 7295
rect 8705 7265 8750 7295
rect 8630 7235 8750 7265
rect 8630 7205 8675 7235
rect 8705 7205 8750 7235
rect 8630 7170 8750 7205
rect 8630 7140 8675 7170
rect 8705 7140 8750 7170
rect 8630 7100 8750 7140
rect 8630 7070 8675 7100
rect 8705 7070 8750 7100
rect 8630 7030 8750 7070
rect 8630 7000 8675 7030
rect 8705 7000 8750 7030
rect 8630 6960 8750 7000
rect 8630 6930 8675 6960
rect 8705 6930 8750 6960
rect 8630 6895 8750 6930
rect 8630 6865 8675 6895
rect 8705 6865 8750 6895
rect 8630 6835 8750 6865
rect 8630 6805 8675 6835
rect 8705 6805 8750 6835
rect 8630 6770 8750 6805
rect 8630 6740 8675 6770
rect 8705 6740 8750 6770
rect 8630 6700 8750 6740
rect 8630 6670 8675 6700
rect 8705 6670 8750 6700
rect 8630 6630 8750 6670
rect 8630 6600 8675 6630
rect 8705 6600 8750 6630
rect 8630 6560 8750 6600
rect 8630 6530 8675 6560
rect 8705 6530 8750 6560
rect 8630 6495 8750 6530
rect 8630 6465 8675 6495
rect 8705 6465 8750 6495
rect 8630 6210 8750 6465
rect 8980 9635 9100 9650
rect 8980 9605 9025 9635
rect 9055 9605 9100 9635
rect 8980 9570 9100 9605
rect 8980 9540 9025 9570
rect 9055 9540 9100 9570
rect 8980 9500 9100 9540
rect 8980 9470 9025 9500
rect 9055 9470 9100 9500
rect 8980 9430 9100 9470
rect 8980 9400 9025 9430
rect 9055 9400 9100 9430
rect 8980 9360 9100 9400
rect 8980 9330 9025 9360
rect 9055 9330 9100 9360
rect 8980 9295 9100 9330
rect 8980 9265 9025 9295
rect 9055 9265 9100 9295
rect 8980 9235 9100 9265
rect 8980 9205 9025 9235
rect 9055 9205 9100 9235
rect 8980 9170 9100 9205
rect 8980 9140 9025 9170
rect 9055 9140 9100 9170
rect 8980 9100 9100 9140
rect 8980 9070 9025 9100
rect 9055 9070 9100 9100
rect 8980 9030 9100 9070
rect 8980 9000 9025 9030
rect 9055 9000 9100 9030
rect 8980 8960 9100 9000
rect 8980 8930 9025 8960
rect 9055 8930 9100 8960
rect 8980 8895 9100 8930
rect 8980 8865 9025 8895
rect 9055 8865 9100 8895
rect 8980 8835 9100 8865
rect 8980 8805 9025 8835
rect 9055 8805 9100 8835
rect 8980 8770 9100 8805
rect 8980 8740 9025 8770
rect 9055 8740 9100 8770
rect 8980 8700 9100 8740
rect 8980 8670 9025 8700
rect 9055 8670 9100 8700
rect 8980 8630 9100 8670
rect 8980 8600 9025 8630
rect 9055 8600 9100 8630
rect 8980 8560 9100 8600
rect 8980 8530 9025 8560
rect 9055 8530 9100 8560
rect 8980 8495 9100 8530
rect 8980 8465 9025 8495
rect 9055 8465 9100 8495
rect 8980 8435 9100 8465
rect 8980 8405 9025 8435
rect 9055 8405 9100 8435
rect 8980 8370 9100 8405
rect 8980 8340 9025 8370
rect 9055 8340 9100 8370
rect 8980 8300 9100 8340
rect 8980 8270 9025 8300
rect 9055 8270 9100 8300
rect 8980 8230 9100 8270
rect 8980 8200 9025 8230
rect 9055 8200 9100 8230
rect 8980 8160 9100 8200
rect 8980 8130 9025 8160
rect 9055 8130 9100 8160
rect 8980 8095 9100 8130
rect 8980 8065 9025 8095
rect 9055 8065 9100 8095
rect 8980 8035 9100 8065
rect 8980 8005 9025 8035
rect 9055 8005 9100 8035
rect 8980 7970 9100 8005
rect 8980 7940 9025 7970
rect 9055 7940 9100 7970
rect 8980 7900 9100 7940
rect 8980 7870 9025 7900
rect 9055 7870 9100 7900
rect 8980 7830 9100 7870
rect 8980 7800 9025 7830
rect 9055 7800 9100 7830
rect 8980 7760 9100 7800
rect 8980 7730 9025 7760
rect 9055 7730 9100 7760
rect 8980 7695 9100 7730
rect 8980 7665 9025 7695
rect 9055 7665 9100 7695
rect 8980 7635 9100 7665
rect 8980 7605 9025 7635
rect 9055 7605 9100 7635
rect 8980 7570 9100 7605
rect 8980 7540 9025 7570
rect 9055 7540 9100 7570
rect 8980 7500 9100 7540
rect 8980 7470 9025 7500
rect 9055 7470 9100 7500
rect 8980 7430 9100 7470
rect 8980 7400 9025 7430
rect 9055 7400 9100 7430
rect 8980 7360 9100 7400
rect 8980 7330 9025 7360
rect 9055 7330 9100 7360
rect 8980 7295 9100 7330
rect 8980 7265 9025 7295
rect 9055 7265 9100 7295
rect 8980 7235 9100 7265
rect 8980 7205 9025 7235
rect 9055 7205 9100 7235
rect 8980 7170 9100 7205
rect 8980 7140 9025 7170
rect 9055 7140 9100 7170
rect 8980 7100 9100 7140
rect 8980 7070 9025 7100
rect 9055 7070 9100 7100
rect 8980 7030 9100 7070
rect 8980 7000 9025 7030
rect 9055 7000 9100 7030
rect 8980 6960 9100 7000
rect 8980 6930 9025 6960
rect 9055 6930 9100 6960
rect 8980 6895 9100 6930
rect 8980 6865 9025 6895
rect 9055 6865 9100 6895
rect 8980 6835 9100 6865
rect 8980 6805 9025 6835
rect 9055 6805 9100 6835
rect 8980 6770 9100 6805
rect 8980 6740 9025 6770
rect 9055 6740 9100 6770
rect 8980 6700 9100 6740
rect 8980 6670 9025 6700
rect 9055 6670 9100 6700
rect 8980 6630 9100 6670
rect 8980 6600 9025 6630
rect 9055 6600 9100 6630
rect 8980 6560 9100 6600
rect 8980 6530 9025 6560
rect 9055 6530 9100 6560
rect 8980 6495 9100 6530
rect 8980 6465 9025 6495
rect 9055 6465 9100 6495
rect 8980 6210 9100 6465
rect 7580 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 7580 6165 7700 6175
rect 7580 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 7580 6125 7700 6135
rect 7580 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 6830 1700 6870 1705
rect 6830 1670 6835 1700
rect 6865 1670 6870 1700
rect 6830 1665 6870 1670
rect 6940 1700 6980 1705
rect 6940 1670 6945 1700
rect 6975 1670 6980 1700
rect 6940 1665 6980 1670
rect 6840 1515 6860 1665
rect 1280 820 1285 850
rect 1315 820 1325 850
rect 1355 820 1365 850
rect 1395 820 1400 850
rect 1280 810 1400 820
rect 1280 780 1285 810
rect 1315 780 1325 810
rect 1355 780 1365 810
rect 1395 780 1400 810
rect 1280 770 1400 780
rect 1280 740 1285 770
rect 1315 740 1325 770
rect 1355 740 1365 770
rect 1395 740 1400 770
rect 1280 735 1400 740
rect 4415 850 4565 855
rect 4415 820 4420 850
rect 4450 820 4475 850
rect 4505 820 4530 850
rect 4560 820 4565 850
rect 4415 810 4565 820
rect 4415 780 4420 810
rect 4450 780 4475 810
rect 4505 780 4530 810
rect 4560 780 4565 810
rect 4415 770 4565 780
rect 4415 740 4420 770
rect 4450 740 4475 770
rect 4505 740 4530 770
rect 4560 740 4565 770
rect 4415 735 4565 740
rect 7580 850 7700 6095
rect 7580 820 7585 850
rect 7615 820 7625 850
rect 7655 820 7665 850
rect 7695 820 7700 850
rect 7580 810 7700 820
rect 7580 780 7585 810
rect 7615 780 7625 810
rect 7655 780 7665 810
rect 7695 780 7700 810
rect 7580 770 7700 780
rect 7580 740 7585 770
rect 7615 740 7625 770
rect 7655 740 7665 770
rect 7695 740 7700 770
rect 7580 735 7700 740
rect -120 -1305 0 -1240
rect -120 -1335 -75 -1305
rect -45 -1335 0 -1305
rect -120 -1370 0 -1335
rect -120 -1400 -75 -1370
rect -45 -1400 0 -1370
rect -120 -1440 0 -1400
rect -120 -1470 -75 -1440
rect -45 -1470 0 -1440
rect -120 -1510 0 -1470
rect -120 -1540 -75 -1510
rect -45 -1540 0 -1510
rect -120 -1580 0 -1540
rect -120 -1610 -75 -1580
rect -45 -1610 0 -1580
rect -120 -1645 0 -1610
rect -120 -1675 -75 -1645
rect -45 -1675 0 -1645
rect -120 -1705 0 -1675
rect -120 -1735 -75 -1705
rect -45 -1735 0 -1705
rect -120 -1770 0 -1735
rect -120 -1800 -75 -1770
rect -45 -1800 0 -1770
rect -120 -1840 0 -1800
rect -120 -1870 -75 -1840
rect -45 -1870 0 -1840
rect -120 -1910 0 -1870
rect -120 -1940 -75 -1910
rect -45 -1940 0 -1910
rect -120 -1980 0 -1940
rect -120 -2010 -75 -1980
rect -45 -2010 0 -1980
rect -120 -2045 0 -2010
rect -120 -2075 -75 -2045
rect -45 -2075 0 -2045
rect -120 -2105 0 -2075
rect -120 -2135 -75 -2105
rect -45 -2135 0 -2105
rect -120 -2170 0 -2135
rect -120 -2200 -75 -2170
rect -45 -2200 0 -2170
rect -120 -2240 0 -2200
rect -120 -2270 -75 -2240
rect -45 -2270 0 -2240
rect -120 -2310 0 -2270
rect -120 -2340 -75 -2310
rect -45 -2340 0 -2310
rect -120 -2380 0 -2340
rect -120 -2410 -75 -2380
rect -45 -2410 0 -2380
rect -120 -2445 0 -2410
rect -120 -2475 -75 -2445
rect -45 -2475 0 -2445
rect -120 -2505 0 -2475
rect -120 -2535 -75 -2505
rect -45 -2535 0 -2505
rect -120 -2570 0 -2535
rect -120 -2600 -75 -2570
rect -45 -2600 0 -2570
rect -120 -2640 0 -2600
rect -120 -2670 -75 -2640
rect -45 -2670 0 -2640
rect -120 -2710 0 -2670
rect -120 -2740 -75 -2710
rect -45 -2740 0 -2710
rect -120 -2780 0 -2740
rect -120 -2810 -75 -2780
rect -45 -2810 0 -2780
rect -120 -2845 0 -2810
rect -120 -2875 -75 -2845
rect -45 -2875 0 -2845
rect -120 -2905 0 -2875
rect -120 -2935 -75 -2905
rect -45 -2935 0 -2905
rect -120 -2970 0 -2935
rect -120 -3000 -75 -2970
rect -45 -3000 0 -2970
rect -120 -3040 0 -3000
rect -120 -3070 -75 -3040
rect -45 -3070 0 -3040
rect -120 -3110 0 -3070
rect -120 -3140 -75 -3110
rect -45 -3140 0 -3110
rect -120 -3180 0 -3140
rect -120 -3210 -75 -3180
rect -45 -3210 0 -3180
rect -120 -3245 0 -3210
rect -120 -3275 -75 -3245
rect -45 -3275 0 -3245
rect -120 -3305 0 -3275
rect -120 -3335 -75 -3305
rect -45 -3335 0 -3305
rect -120 -3370 0 -3335
rect -120 -3400 -75 -3370
rect -45 -3400 0 -3370
rect -120 -3440 0 -3400
rect -120 -3470 -75 -3440
rect -45 -3470 0 -3440
rect -120 -3510 0 -3470
rect -120 -3540 -75 -3510
rect -45 -3540 0 -3510
rect -120 -3580 0 -3540
rect -120 -3610 -75 -3580
rect -45 -3610 0 -3580
rect -120 -3645 0 -3610
rect -120 -3675 -75 -3645
rect -45 -3675 0 -3645
rect -120 -3705 0 -3675
rect -120 -3735 -75 -3705
rect -45 -3735 0 -3705
rect -120 -3770 0 -3735
rect -120 -3800 -75 -3770
rect -45 -3800 0 -3770
rect -120 -3840 0 -3800
rect -120 -3870 -75 -3840
rect -45 -3870 0 -3840
rect -120 -3910 0 -3870
rect -120 -3940 -75 -3910
rect -45 -3940 0 -3910
rect -120 -3980 0 -3940
rect -120 -4010 -75 -3980
rect -45 -4010 0 -3980
rect -120 -4045 0 -4010
rect -120 -4075 -75 -4045
rect -45 -4075 0 -4045
rect -120 -4105 0 -4075
rect -120 -4135 -75 -4105
rect -45 -4135 0 -4105
rect -120 -4170 0 -4135
rect -120 -4200 -75 -4170
rect -45 -4200 0 -4170
rect -120 -4240 0 -4200
rect -120 -4270 -75 -4240
rect -45 -4270 0 -4240
rect -120 -4310 0 -4270
rect -120 -4340 -75 -4310
rect -45 -4340 0 -4310
rect -120 -4380 0 -4340
rect -120 -4410 -75 -4380
rect -45 -4410 0 -4380
rect -120 -4445 0 -4410
rect -120 -4475 -75 -4445
rect -45 -4475 0 -4445
rect -120 -4490 0 -4475
rect 230 -1305 350 -1240
rect 230 -1335 275 -1305
rect 305 -1335 350 -1305
rect 230 -1370 350 -1335
rect 230 -1400 275 -1370
rect 305 -1400 350 -1370
rect 230 -1440 350 -1400
rect 230 -1470 275 -1440
rect 305 -1470 350 -1440
rect 230 -1510 350 -1470
rect 230 -1540 275 -1510
rect 305 -1540 350 -1510
rect 230 -1580 350 -1540
rect 230 -1610 275 -1580
rect 305 -1610 350 -1580
rect 230 -1645 350 -1610
rect 230 -1675 275 -1645
rect 305 -1675 350 -1645
rect 230 -1705 350 -1675
rect 230 -1735 275 -1705
rect 305 -1735 350 -1705
rect 230 -1770 350 -1735
rect 230 -1800 275 -1770
rect 305 -1800 350 -1770
rect 230 -1840 350 -1800
rect 230 -1870 275 -1840
rect 305 -1870 350 -1840
rect 230 -1910 350 -1870
rect 230 -1940 275 -1910
rect 305 -1940 350 -1910
rect 230 -1980 350 -1940
rect 230 -2010 275 -1980
rect 305 -2010 350 -1980
rect 230 -2045 350 -2010
rect 230 -2075 275 -2045
rect 305 -2075 350 -2045
rect 230 -2105 350 -2075
rect 230 -2135 275 -2105
rect 305 -2135 350 -2105
rect 230 -2170 350 -2135
rect 230 -2200 275 -2170
rect 305 -2200 350 -2170
rect 230 -2240 350 -2200
rect 230 -2270 275 -2240
rect 305 -2270 350 -2240
rect 230 -2310 350 -2270
rect 230 -2340 275 -2310
rect 305 -2340 350 -2310
rect 230 -2380 350 -2340
rect 230 -2410 275 -2380
rect 305 -2410 350 -2380
rect 230 -2445 350 -2410
rect 230 -2475 275 -2445
rect 305 -2475 350 -2445
rect 230 -2505 350 -2475
rect 230 -2535 275 -2505
rect 305 -2535 350 -2505
rect 230 -2570 350 -2535
rect 230 -2600 275 -2570
rect 305 -2600 350 -2570
rect 230 -2640 350 -2600
rect 230 -2670 275 -2640
rect 305 -2670 350 -2640
rect 230 -2710 350 -2670
rect 230 -2740 275 -2710
rect 305 -2740 350 -2710
rect 230 -2780 350 -2740
rect 230 -2810 275 -2780
rect 305 -2810 350 -2780
rect 230 -2845 350 -2810
rect 230 -2875 275 -2845
rect 305 -2875 350 -2845
rect 230 -2905 350 -2875
rect 230 -2935 275 -2905
rect 305 -2935 350 -2905
rect 230 -2970 350 -2935
rect 230 -3000 275 -2970
rect 305 -3000 350 -2970
rect 230 -3040 350 -3000
rect 230 -3070 275 -3040
rect 305 -3070 350 -3040
rect 230 -3110 350 -3070
rect 230 -3140 275 -3110
rect 305 -3140 350 -3110
rect 230 -3180 350 -3140
rect 230 -3210 275 -3180
rect 305 -3210 350 -3180
rect 230 -3245 350 -3210
rect 230 -3275 275 -3245
rect 305 -3275 350 -3245
rect 230 -3305 350 -3275
rect 230 -3335 275 -3305
rect 305 -3335 350 -3305
rect 230 -3370 350 -3335
rect 230 -3400 275 -3370
rect 305 -3400 350 -3370
rect 230 -3440 350 -3400
rect 230 -3470 275 -3440
rect 305 -3470 350 -3440
rect 230 -3510 350 -3470
rect 230 -3540 275 -3510
rect 305 -3540 350 -3510
rect 230 -3580 350 -3540
rect 230 -3610 275 -3580
rect 305 -3610 350 -3580
rect 230 -3645 350 -3610
rect 230 -3675 275 -3645
rect 305 -3675 350 -3645
rect 230 -3705 350 -3675
rect 230 -3735 275 -3705
rect 305 -3735 350 -3705
rect 230 -3770 350 -3735
rect 230 -3800 275 -3770
rect 305 -3800 350 -3770
rect 230 -3840 350 -3800
rect 230 -3870 275 -3840
rect 305 -3870 350 -3840
rect 230 -3910 350 -3870
rect 230 -3940 275 -3910
rect 305 -3940 350 -3910
rect 230 -3980 350 -3940
rect 230 -4010 275 -3980
rect 305 -4010 350 -3980
rect 230 -4045 350 -4010
rect 230 -4075 275 -4045
rect 305 -4075 350 -4045
rect 230 -4105 350 -4075
rect 230 -4135 275 -4105
rect 305 -4135 350 -4105
rect 230 -4170 350 -4135
rect 230 -4200 275 -4170
rect 305 -4200 350 -4170
rect 230 -4240 350 -4200
rect 230 -4270 275 -4240
rect 305 -4270 350 -4240
rect 230 -4310 350 -4270
rect 230 -4340 275 -4310
rect 305 -4340 350 -4310
rect 230 -4380 350 -4340
rect 230 -4410 275 -4380
rect 305 -4410 350 -4380
rect 230 -4445 350 -4410
rect 230 -4475 275 -4445
rect 305 -4475 350 -4445
rect 230 -4490 350 -4475
rect 580 -1305 700 -1240
rect 580 -1335 625 -1305
rect 655 -1335 700 -1305
rect 580 -1370 700 -1335
rect 580 -1400 625 -1370
rect 655 -1400 700 -1370
rect 580 -1440 700 -1400
rect 580 -1470 625 -1440
rect 655 -1470 700 -1440
rect 580 -1510 700 -1470
rect 580 -1540 625 -1510
rect 655 -1540 700 -1510
rect 580 -1580 700 -1540
rect 580 -1610 625 -1580
rect 655 -1610 700 -1580
rect 580 -1645 700 -1610
rect 580 -1675 625 -1645
rect 655 -1675 700 -1645
rect 580 -1705 700 -1675
rect 580 -1735 625 -1705
rect 655 -1735 700 -1705
rect 580 -1770 700 -1735
rect 580 -1800 625 -1770
rect 655 -1800 700 -1770
rect 580 -1840 700 -1800
rect 580 -1870 625 -1840
rect 655 -1870 700 -1840
rect 580 -1910 700 -1870
rect 580 -1940 625 -1910
rect 655 -1940 700 -1910
rect 580 -1980 700 -1940
rect 580 -2010 625 -1980
rect 655 -2010 700 -1980
rect 580 -2045 700 -2010
rect 580 -2075 625 -2045
rect 655 -2075 700 -2045
rect 580 -2105 700 -2075
rect 580 -2135 625 -2105
rect 655 -2135 700 -2105
rect 580 -2170 700 -2135
rect 580 -2200 625 -2170
rect 655 -2200 700 -2170
rect 580 -2240 700 -2200
rect 580 -2270 625 -2240
rect 655 -2270 700 -2240
rect 580 -2310 700 -2270
rect 580 -2340 625 -2310
rect 655 -2340 700 -2310
rect 580 -2380 700 -2340
rect 580 -2410 625 -2380
rect 655 -2410 700 -2380
rect 580 -2445 700 -2410
rect 580 -2475 625 -2445
rect 655 -2475 700 -2445
rect 580 -2505 700 -2475
rect 580 -2535 625 -2505
rect 655 -2535 700 -2505
rect 580 -2570 700 -2535
rect 580 -2600 625 -2570
rect 655 -2600 700 -2570
rect 580 -2640 700 -2600
rect 580 -2670 625 -2640
rect 655 -2670 700 -2640
rect 580 -2710 700 -2670
rect 580 -2740 625 -2710
rect 655 -2740 700 -2710
rect 580 -2780 700 -2740
rect 580 -2810 625 -2780
rect 655 -2810 700 -2780
rect 580 -2845 700 -2810
rect 580 -2875 625 -2845
rect 655 -2875 700 -2845
rect 580 -2905 700 -2875
rect 580 -2935 625 -2905
rect 655 -2935 700 -2905
rect 580 -2970 700 -2935
rect 580 -3000 625 -2970
rect 655 -3000 700 -2970
rect 580 -3040 700 -3000
rect 580 -3070 625 -3040
rect 655 -3070 700 -3040
rect 580 -3110 700 -3070
rect 580 -3140 625 -3110
rect 655 -3140 700 -3110
rect 580 -3180 700 -3140
rect 580 -3210 625 -3180
rect 655 -3210 700 -3180
rect 580 -3245 700 -3210
rect 580 -3275 625 -3245
rect 655 -3275 700 -3245
rect 580 -3305 700 -3275
rect 580 -3335 625 -3305
rect 655 -3335 700 -3305
rect 580 -3370 700 -3335
rect 580 -3400 625 -3370
rect 655 -3400 700 -3370
rect 580 -3440 700 -3400
rect 580 -3470 625 -3440
rect 655 -3470 700 -3440
rect 580 -3510 700 -3470
rect 580 -3540 625 -3510
rect 655 -3540 700 -3510
rect 580 -3580 700 -3540
rect 580 -3610 625 -3580
rect 655 -3610 700 -3580
rect 580 -3645 700 -3610
rect 580 -3675 625 -3645
rect 655 -3675 700 -3645
rect 580 -3705 700 -3675
rect 580 -3735 625 -3705
rect 655 -3735 700 -3705
rect 580 -3770 700 -3735
rect 580 -3800 625 -3770
rect 655 -3800 700 -3770
rect 580 -3840 700 -3800
rect 580 -3870 625 -3840
rect 655 -3870 700 -3840
rect 580 -3910 700 -3870
rect 580 -3940 625 -3910
rect 655 -3940 700 -3910
rect 580 -3980 700 -3940
rect 580 -4010 625 -3980
rect 655 -4010 700 -3980
rect 580 -4045 700 -4010
rect 580 -4075 625 -4045
rect 655 -4075 700 -4045
rect 580 -4105 700 -4075
rect 580 -4135 625 -4105
rect 655 -4135 700 -4105
rect 580 -4170 700 -4135
rect 580 -4200 625 -4170
rect 655 -4200 700 -4170
rect 580 -4240 700 -4200
rect 580 -4270 625 -4240
rect 655 -4270 700 -4240
rect 580 -4310 700 -4270
rect 580 -4340 625 -4310
rect 655 -4340 700 -4310
rect 580 -4380 700 -4340
rect 580 -4410 625 -4380
rect 655 -4410 700 -4380
rect 580 -4445 700 -4410
rect 580 -4475 625 -4445
rect 655 -4475 700 -4445
rect 580 -4490 700 -4475
rect 930 -1305 1050 -1240
rect 930 -1335 975 -1305
rect 1005 -1335 1050 -1305
rect 930 -1370 1050 -1335
rect 930 -1400 975 -1370
rect 1005 -1400 1050 -1370
rect 930 -1440 1050 -1400
rect 930 -1470 975 -1440
rect 1005 -1470 1050 -1440
rect 930 -1510 1050 -1470
rect 930 -1540 975 -1510
rect 1005 -1540 1050 -1510
rect 930 -1580 1050 -1540
rect 930 -1610 975 -1580
rect 1005 -1610 1050 -1580
rect 930 -1645 1050 -1610
rect 930 -1675 975 -1645
rect 1005 -1675 1050 -1645
rect 930 -1705 1050 -1675
rect 930 -1735 975 -1705
rect 1005 -1735 1050 -1705
rect 930 -1770 1050 -1735
rect 930 -1800 975 -1770
rect 1005 -1800 1050 -1770
rect 930 -1840 1050 -1800
rect 930 -1870 975 -1840
rect 1005 -1870 1050 -1840
rect 930 -1910 1050 -1870
rect 930 -1940 975 -1910
rect 1005 -1940 1050 -1910
rect 930 -1980 1050 -1940
rect 930 -2010 975 -1980
rect 1005 -2010 1050 -1980
rect 930 -2045 1050 -2010
rect 930 -2075 975 -2045
rect 1005 -2075 1050 -2045
rect 930 -2105 1050 -2075
rect 930 -2135 975 -2105
rect 1005 -2135 1050 -2105
rect 930 -2170 1050 -2135
rect 930 -2200 975 -2170
rect 1005 -2200 1050 -2170
rect 930 -2240 1050 -2200
rect 930 -2270 975 -2240
rect 1005 -2270 1050 -2240
rect 930 -2310 1050 -2270
rect 930 -2340 975 -2310
rect 1005 -2340 1050 -2310
rect 930 -2380 1050 -2340
rect 930 -2410 975 -2380
rect 1005 -2410 1050 -2380
rect 930 -2445 1050 -2410
rect 930 -2475 975 -2445
rect 1005 -2475 1050 -2445
rect 930 -2505 1050 -2475
rect 930 -2535 975 -2505
rect 1005 -2535 1050 -2505
rect 930 -2570 1050 -2535
rect 930 -2600 975 -2570
rect 1005 -2600 1050 -2570
rect 930 -2640 1050 -2600
rect 930 -2670 975 -2640
rect 1005 -2670 1050 -2640
rect 930 -2710 1050 -2670
rect 930 -2740 975 -2710
rect 1005 -2740 1050 -2710
rect 930 -2780 1050 -2740
rect 930 -2810 975 -2780
rect 1005 -2810 1050 -2780
rect 930 -2845 1050 -2810
rect 930 -2875 975 -2845
rect 1005 -2875 1050 -2845
rect 930 -2905 1050 -2875
rect 930 -2935 975 -2905
rect 1005 -2935 1050 -2905
rect 930 -2970 1050 -2935
rect 930 -3000 975 -2970
rect 1005 -3000 1050 -2970
rect 930 -3040 1050 -3000
rect 930 -3070 975 -3040
rect 1005 -3070 1050 -3040
rect 930 -3110 1050 -3070
rect 930 -3140 975 -3110
rect 1005 -3140 1050 -3110
rect 930 -3180 1050 -3140
rect 930 -3210 975 -3180
rect 1005 -3210 1050 -3180
rect 930 -3245 1050 -3210
rect 930 -3275 975 -3245
rect 1005 -3275 1050 -3245
rect 930 -3305 1050 -3275
rect 930 -3335 975 -3305
rect 1005 -3335 1050 -3305
rect 930 -3370 1050 -3335
rect 930 -3400 975 -3370
rect 1005 -3400 1050 -3370
rect 930 -3440 1050 -3400
rect 930 -3470 975 -3440
rect 1005 -3470 1050 -3440
rect 930 -3510 1050 -3470
rect 930 -3540 975 -3510
rect 1005 -3540 1050 -3510
rect 930 -3580 1050 -3540
rect 930 -3610 975 -3580
rect 1005 -3610 1050 -3580
rect 930 -3645 1050 -3610
rect 930 -3675 975 -3645
rect 1005 -3675 1050 -3645
rect 930 -3705 1050 -3675
rect 930 -3735 975 -3705
rect 1005 -3735 1050 -3705
rect 930 -3770 1050 -3735
rect 930 -3800 975 -3770
rect 1005 -3800 1050 -3770
rect 930 -3840 1050 -3800
rect 930 -3870 975 -3840
rect 1005 -3870 1050 -3840
rect 930 -3910 1050 -3870
rect 930 -3940 975 -3910
rect 1005 -3940 1050 -3910
rect 930 -3980 1050 -3940
rect 930 -4010 975 -3980
rect 1005 -4010 1050 -3980
rect 930 -4045 1050 -4010
rect 930 -4075 975 -4045
rect 1005 -4075 1050 -4045
rect 930 -4105 1050 -4075
rect 930 -4135 975 -4105
rect 1005 -4135 1050 -4105
rect 930 -4170 1050 -4135
rect 930 -4200 975 -4170
rect 1005 -4200 1050 -4170
rect 930 -4240 1050 -4200
rect 930 -4270 975 -4240
rect 1005 -4270 1050 -4240
rect 930 -4310 1050 -4270
rect 930 -4340 975 -4310
rect 1005 -4340 1050 -4310
rect 930 -4380 1050 -4340
rect 930 -4410 975 -4380
rect 1005 -4410 1050 -4380
rect 930 -4445 1050 -4410
rect 930 -4475 975 -4445
rect 1005 -4475 1050 -4445
rect 930 -4490 1050 -4475
rect 1280 -1305 1400 -1240
rect 1280 -1335 1325 -1305
rect 1355 -1335 1400 -1305
rect 1280 -1370 1400 -1335
rect 1280 -1400 1325 -1370
rect 1355 -1400 1400 -1370
rect 1280 -1440 1400 -1400
rect 1280 -1470 1325 -1440
rect 1355 -1470 1400 -1440
rect 1280 -1510 1400 -1470
rect 1280 -1540 1325 -1510
rect 1355 -1540 1400 -1510
rect 1280 -1580 1400 -1540
rect 1280 -1610 1325 -1580
rect 1355 -1610 1400 -1580
rect 1280 -1645 1400 -1610
rect 1280 -1675 1325 -1645
rect 1355 -1675 1400 -1645
rect 1280 -1705 1400 -1675
rect 1280 -1735 1325 -1705
rect 1355 -1735 1400 -1705
rect 1280 -1770 1400 -1735
rect 1280 -1800 1325 -1770
rect 1355 -1800 1400 -1770
rect 1280 -1840 1400 -1800
rect 1280 -1870 1325 -1840
rect 1355 -1870 1400 -1840
rect 1280 -1910 1400 -1870
rect 1280 -1940 1325 -1910
rect 1355 -1940 1400 -1910
rect 1280 -1980 1400 -1940
rect 1280 -2010 1325 -1980
rect 1355 -2010 1400 -1980
rect 1280 -2045 1400 -2010
rect 1280 -2075 1325 -2045
rect 1355 -2075 1400 -2045
rect 1280 -2105 1400 -2075
rect 1280 -2135 1325 -2105
rect 1355 -2135 1400 -2105
rect 1280 -2170 1400 -2135
rect 1280 -2200 1325 -2170
rect 1355 -2200 1400 -2170
rect 1280 -2240 1400 -2200
rect 1280 -2270 1325 -2240
rect 1355 -2270 1400 -2240
rect 1280 -2310 1400 -2270
rect 1280 -2340 1325 -2310
rect 1355 -2340 1400 -2310
rect 1280 -2380 1400 -2340
rect 1280 -2410 1325 -2380
rect 1355 -2410 1400 -2380
rect 1280 -2445 1400 -2410
rect 1280 -2475 1325 -2445
rect 1355 -2475 1400 -2445
rect 1280 -2505 1400 -2475
rect 1280 -2535 1325 -2505
rect 1355 -2535 1400 -2505
rect 1280 -2570 1400 -2535
rect 1280 -2600 1325 -2570
rect 1355 -2600 1400 -2570
rect 1280 -2640 1400 -2600
rect 1280 -2670 1325 -2640
rect 1355 -2670 1400 -2640
rect 1280 -2710 1400 -2670
rect 1280 -2740 1325 -2710
rect 1355 -2740 1400 -2710
rect 1280 -2780 1400 -2740
rect 1280 -2810 1325 -2780
rect 1355 -2810 1400 -2780
rect 1280 -2845 1400 -2810
rect 1280 -2875 1325 -2845
rect 1355 -2875 1400 -2845
rect 1280 -2905 1400 -2875
rect 1280 -2935 1325 -2905
rect 1355 -2935 1400 -2905
rect 1280 -2970 1400 -2935
rect 1280 -3000 1325 -2970
rect 1355 -3000 1400 -2970
rect 1280 -3040 1400 -3000
rect 1280 -3070 1325 -3040
rect 1355 -3070 1400 -3040
rect 1280 -3110 1400 -3070
rect 1280 -3140 1325 -3110
rect 1355 -3140 1400 -3110
rect 1280 -3180 1400 -3140
rect 1280 -3210 1325 -3180
rect 1355 -3210 1400 -3180
rect 1280 -3245 1400 -3210
rect 1280 -3275 1325 -3245
rect 1355 -3275 1400 -3245
rect 1280 -3305 1400 -3275
rect 1280 -3335 1325 -3305
rect 1355 -3335 1400 -3305
rect 1280 -3370 1400 -3335
rect 1280 -3400 1325 -3370
rect 1355 -3400 1400 -3370
rect 1280 -3440 1400 -3400
rect 1280 -3470 1325 -3440
rect 1355 -3470 1400 -3440
rect 1280 -3510 1400 -3470
rect 1280 -3540 1325 -3510
rect 1355 -3540 1400 -3510
rect 1280 -3580 1400 -3540
rect 1280 -3610 1325 -3580
rect 1355 -3610 1400 -3580
rect 1280 -3645 1400 -3610
rect 1280 -3675 1325 -3645
rect 1355 -3675 1400 -3645
rect 1280 -3705 1400 -3675
rect 1280 -3735 1325 -3705
rect 1355 -3735 1400 -3705
rect 1280 -3770 1400 -3735
rect 1280 -3800 1325 -3770
rect 1355 -3800 1400 -3770
rect 1280 -3840 1400 -3800
rect 1280 -3870 1325 -3840
rect 1355 -3870 1400 -3840
rect 1280 -3910 1400 -3870
rect 1280 -3940 1325 -3910
rect 1355 -3940 1400 -3910
rect 1280 -3980 1400 -3940
rect 1280 -4010 1325 -3980
rect 1355 -4010 1400 -3980
rect 1280 -4045 1400 -4010
rect 1280 -4075 1325 -4045
rect 1355 -4075 1400 -4045
rect 1280 -4105 1400 -4075
rect 1280 -4135 1325 -4105
rect 1355 -4135 1400 -4105
rect 1280 -4170 1400 -4135
rect 1280 -4200 1325 -4170
rect 1355 -4200 1400 -4170
rect 1280 -4240 1400 -4200
rect 1280 -4270 1325 -4240
rect 1355 -4270 1400 -4240
rect 1280 -4310 1400 -4270
rect 1280 -4340 1325 -4310
rect 1355 -4340 1400 -4310
rect 1280 -4380 1400 -4340
rect 1280 -4410 1325 -4380
rect 1355 -4410 1400 -4380
rect 1280 -4445 1400 -4410
rect 1280 -4475 1325 -4445
rect 1355 -4475 1400 -4445
rect 1280 -4490 1400 -4475
rect 1630 -1305 1750 -1240
rect 1630 -1335 1675 -1305
rect 1705 -1335 1750 -1305
rect 1630 -1370 1750 -1335
rect 1630 -1400 1675 -1370
rect 1705 -1400 1750 -1370
rect 1630 -1440 1750 -1400
rect 1630 -1470 1675 -1440
rect 1705 -1470 1750 -1440
rect 1630 -1510 1750 -1470
rect 1630 -1540 1675 -1510
rect 1705 -1540 1750 -1510
rect 1630 -1580 1750 -1540
rect 1630 -1610 1675 -1580
rect 1705 -1610 1750 -1580
rect 1630 -1645 1750 -1610
rect 1630 -1675 1675 -1645
rect 1705 -1675 1750 -1645
rect 1630 -1705 1750 -1675
rect 1630 -1735 1675 -1705
rect 1705 -1735 1750 -1705
rect 1630 -1770 1750 -1735
rect 1630 -1800 1675 -1770
rect 1705 -1800 1750 -1770
rect 1630 -1840 1750 -1800
rect 1630 -1870 1675 -1840
rect 1705 -1870 1750 -1840
rect 1630 -1910 1750 -1870
rect 1630 -1940 1675 -1910
rect 1705 -1940 1750 -1910
rect 1630 -1980 1750 -1940
rect 1630 -2010 1675 -1980
rect 1705 -2010 1750 -1980
rect 1630 -2045 1750 -2010
rect 1630 -2075 1675 -2045
rect 1705 -2075 1750 -2045
rect 1630 -2105 1750 -2075
rect 1630 -2135 1675 -2105
rect 1705 -2135 1750 -2105
rect 1630 -2170 1750 -2135
rect 1630 -2200 1675 -2170
rect 1705 -2200 1750 -2170
rect 1630 -2240 1750 -2200
rect 1630 -2270 1675 -2240
rect 1705 -2270 1750 -2240
rect 1630 -2310 1750 -2270
rect 1630 -2340 1675 -2310
rect 1705 -2340 1750 -2310
rect 1630 -2380 1750 -2340
rect 1630 -2410 1675 -2380
rect 1705 -2410 1750 -2380
rect 1630 -2445 1750 -2410
rect 1630 -2475 1675 -2445
rect 1705 -2475 1750 -2445
rect 1630 -2505 1750 -2475
rect 1630 -2535 1675 -2505
rect 1705 -2535 1750 -2505
rect 1630 -2570 1750 -2535
rect 1630 -2600 1675 -2570
rect 1705 -2600 1750 -2570
rect 1630 -2640 1750 -2600
rect 1630 -2670 1675 -2640
rect 1705 -2670 1750 -2640
rect 1630 -2710 1750 -2670
rect 1630 -2740 1675 -2710
rect 1705 -2740 1750 -2710
rect 1630 -2780 1750 -2740
rect 1630 -2810 1675 -2780
rect 1705 -2810 1750 -2780
rect 1630 -2845 1750 -2810
rect 1630 -2875 1675 -2845
rect 1705 -2875 1750 -2845
rect 1630 -2905 1750 -2875
rect 1630 -2935 1675 -2905
rect 1705 -2935 1750 -2905
rect 1630 -2970 1750 -2935
rect 1630 -3000 1675 -2970
rect 1705 -3000 1750 -2970
rect 1630 -3040 1750 -3000
rect 1630 -3070 1675 -3040
rect 1705 -3070 1750 -3040
rect 1630 -3110 1750 -3070
rect 1630 -3140 1675 -3110
rect 1705 -3140 1750 -3110
rect 1630 -3180 1750 -3140
rect 1630 -3210 1675 -3180
rect 1705 -3210 1750 -3180
rect 1630 -3245 1750 -3210
rect 1630 -3275 1675 -3245
rect 1705 -3275 1750 -3245
rect 1630 -3305 1750 -3275
rect 1630 -3335 1675 -3305
rect 1705 -3335 1750 -3305
rect 1630 -3370 1750 -3335
rect 1630 -3400 1675 -3370
rect 1705 -3400 1750 -3370
rect 1630 -3440 1750 -3400
rect 1630 -3470 1675 -3440
rect 1705 -3470 1750 -3440
rect 1630 -3510 1750 -3470
rect 1630 -3540 1675 -3510
rect 1705 -3540 1750 -3510
rect 1630 -3580 1750 -3540
rect 1630 -3610 1675 -3580
rect 1705 -3610 1750 -3580
rect 1630 -3645 1750 -3610
rect 1630 -3675 1675 -3645
rect 1705 -3675 1750 -3645
rect 1630 -3705 1750 -3675
rect 1630 -3735 1675 -3705
rect 1705 -3735 1750 -3705
rect 1630 -3770 1750 -3735
rect 1630 -3800 1675 -3770
rect 1705 -3800 1750 -3770
rect 1630 -3840 1750 -3800
rect 1630 -3870 1675 -3840
rect 1705 -3870 1750 -3840
rect 1630 -3910 1750 -3870
rect 1630 -3940 1675 -3910
rect 1705 -3940 1750 -3910
rect 1630 -3980 1750 -3940
rect 1630 -4010 1675 -3980
rect 1705 -4010 1750 -3980
rect 1630 -4045 1750 -4010
rect 1630 -4075 1675 -4045
rect 1705 -4075 1750 -4045
rect 1630 -4105 1750 -4075
rect 1630 -4135 1675 -4105
rect 1705 -4135 1750 -4105
rect 1630 -4170 1750 -4135
rect 1630 -4200 1675 -4170
rect 1705 -4200 1750 -4170
rect 1630 -4240 1750 -4200
rect 1630 -4270 1675 -4240
rect 1705 -4270 1750 -4240
rect 1630 -4310 1750 -4270
rect 1630 -4340 1675 -4310
rect 1705 -4340 1750 -4310
rect 1630 -4380 1750 -4340
rect 1630 -4410 1675 -4380
rect 1705 -4410 1750 -4380
rect 1630 -4445 1750 -4410
rect 1630 -4475 1675 -4445
rect 1705 -4475 1750 -4445
rect 1630 -4490 1750 -4475
rect 1980 -1305 2100 -1240
rect 1980 -1335 2025 -1305
rect 2055 -1335 2100 -1305
rect 1980 -1370 2100 -1335
rect 1980 -1400 2025 -1370
rect 2055 -1400 2100 -1370
rect 1980 -1440 2100 -1400
rect 1980 -1470 2025 -1440
rect 2055 -1470 2100 -1440
rect 1980 -1510 2100 -1470
rect 1980 -1540 2025 -1510
rect 2055 -1540 2100 -1510
rect 1980 -1580 2100 -1540
rect 1980 -1610 2025 -1580
rect 2055 -1610 2100 -1580
rect 1980 -1645 2100 -1610
rect 1980 -1675 2025 -1645
rect 2055 -1675 2100 -1645
rect 1980 -1705 2100 -1675
rect 1980 -1735 2025 -1705
rect 2055 -1735 2100 -1705
rect 1980 -1770 2100 -1735
rect 1980 -1800 2025 -1770
rect 2055 -1800 2100 -1770
rect 1980 -1840 2100 -1800
rect 1980 -1870 2025 -1840
rect 2055 -1870 2100 -1840
rect 1980 -1910 2100 -1870
rect 1980 -1940 2025 -1910
rect 2055 -1940 2100 -1910
rect 1980 -1980 2100 -1940
rect 1980 -2010 2025 -1980
rect 2055 -2010 2100 -1980
rect 1980 -2045 2100 -2010
rect 1980 -2075 2025 -2045
rect 2055 -2075 2100 -2045
rect 1980 -2105 2100 -2075
rect 1980 -2135 2025 -2105
rect 2055 -2135 2100 -2105
rect 1980 -2170 2100 -2135
rect 1980 -2200 2025 -2170
rect 2055 -2200 2100 -2170
rect 1980 -2240 2100 -2200
rect 1980 -2270 2025 -2240
rect 2055 -2270 2100 -2240
rect 1980 -2310 2100 -2270
rect 1980 -2340 2025 -2310
rect 2055 -2340 2100 -2310
rect 1980 -2380 2100 -2340
rect 1980 -2410 2025 -2380
rect 2055 -2410 2100 -2380
rect 1980 -2445 2100 -2410
rect 1980 -2475 2025 -2445
rect 2055 -2475 2100 -2445
rect 1980 -2505 2100 -2475
rect 1980 -2535 2025 -2505
rect 2055 -2535 2100 -2505
rect 1980 -2570 2100 -2535
rect 1980 -2600 2025 -2570
rect 2055 -2600 2100 -2570
rect 1980 -2640 2100 -2600
rect 1980 -2670 2025 -2640
rect 2055 -2670 2100 -2640
rect 1980 -2710 2100 -2670
rect 1980 -2740 2025 -2710
rect 2055 -2740 2100 -2710
rect 1980 -2780 2100 -2740
rect 1980 -2810 2025 -2780
rect 2055 -2810 2100 -2780
rect 1980 -2845 2100 -2810
rect 1980 -2875 2025 -2845
rect 2055 -2875 2100 -2845
rect 1980 -2905 2100 -2875
rect 1980 -2935 2025 -2905
rect 2055 -2935 2100 -2905
rect 1980 -2970 2100 -2935
rect 1980 -3000 2025 -2970
rect 2055 -3000 2100 -2970
rect 1980 -3040 2100 -3000
rect 1980 -3070 2025 -3040
rect 2055 -3070 2100 -3040
rect 1980 -3110 2100 -3070
rect 1980 -3140 2025 -3110
rect 2055 -3140 2100 -3110
rect 1980 -3180 2100 -3140
rect 1980 -3210 2025 -3180
rect 2055 -3210 2100 -3180
rect 1980 -3245 2100 -3210
rect 1980 -3275 2025 -3245
rect 2055 -3275 2100 -3245
rect 1980 -3305 2100 -3275
rect 1980 -3335 2025 -3305
rect 2055 -3335 2100 -3305
rect 1980 -3370 2100 -3335
rect 1980 -3400 2025 -3370
rect 2055 -3400 2100 -3370
rect 1980 -3440 2100 -3400
rect 1980 -3470 2025 -3440
rect 2055 -3470 2100 -3440
rect 1980 -3510 2100 -3470
rect 1980 -3540 2025 -3510
rect 2055 -3540 2100 -3510
rect 1980 -3580 2100 -3540
rect 1980 -3610 2025 -3580
rect 2055 -3610 2100 -3580
rect 1980 -3645 2100 -3610
rect 1980 -3675 2025 -3645
rect 2055 -3675 2100 -3645
rect 1980 -3705 2100 -3675
rect 1980 -3735 2025 -3705
rect 2055 -3735 2100 -3705
rect 1980 -3770 2100 -3735
rect 1980 -3800 2025 -3770
rect 2055 -3800 2100 -3770
rect 1980 -3840 2100 -3800
rect 1980 -3870 2025 -3840
rect 2055 -3870 2100 -3840
rect 1980 -3910 2100 -3870
rect 1980 -3940 2025 -3910
rect 2055 -3940 2100 -3910
rect 1980 -3980 2100 -3940
rect 1980 -4010 2025 -3980
rect 2055 -4010 2100 -3980
rect 1980 -4045 2100 -4010
rect 1980 -4075 2025 -4045
rect 2055 -4075 2100 -4045
rect 1980 -4105 2100 -4075
rect 1980 -4135 2025 -4105
rect 2055 -4135 2100 -4105
rect 1980 -4170 2100 -4135
rect 1980 -4200 2025 -4170
rect 2055 -4200 2100 -4170
rect 1980 -4240 2100 -4200
rect 1980 -4270 2025 -4240
rect 2055 -4270 2100 -4240
rect 1980 -4310 2100 -4270
rect 1980 -4340 2025 -4310
rect 2055 -4340 2100 -4310
rect 1980 -4380 2100 -4340
rect 1980 -4410 2025 -4380
rect 2055 -4410 2100 -4380
rect 1980 -4445 2100 -4410
rect 1980 -4475 2025 -4445
rect 2055 -4475 2100 -4445
rect 1980 -4490 2100 -4475
rect 2330 -1305 2450 -1240
rect 2330 -1335 2375 -1305
rect 2405 -1335 2450 -1305
rect 2330 -1370 2450 -1335
rect 2330 -1400 2375 -1370
rect 2405 -1400 2450 -1370
rect 2330 -1440 2450 -1400
rect 2330 -1470 2375 -1440
rect 2405 -1470 2450 -1440
rect 2330 -1510 2450 -1470
rect 2330 -1540 2375 -1510
rect 2405 -1540 2450 -1510
rect 2330 -1580 2450 -1540
rect 2330 -1610 2375 -1580
rect 2405 -1610 2450 -1580
rect 2330 -1645 2450 -1610
rect 2330 -1675 2375 -1645
rect 2405 -1675 2450 -1645
rect 2330 -1705 2450 -1675
rect 2330 -1735 2375 -1705
rect 2405 -1735 2450 -1705
rect 2330 -1770 2450 -1735
rect 2330 -1800 2375 -1770
rect 2405 -1800 2450 -1770
rect 2330 -1840 2450 -1800
rect 2330 -1870 2375 -1840
rect 2405 -1870 2450 -1840
rect 2330 -1910 2450 -1870
rect 2330 -1940 2375 -1910
rect 2405 -1940 2450 -1910
rect 2330 -1980 2450 -1940
rect 2330 -2010 2375 -1980
rect 2405 -2010 2450 -1980
rect 2330 -2045 2450 -2010
rect 2330 -2075 2375 -2045
rect 2405 -2075 2450 -2045
rect 2330 -2105 2450 -2075
rect 2330 -2135 2375 -2105
rect 2405 -2135 2450 -2105
rect 2330 -2170 2450 -2135
rect 2330 -2200 2375 -2170
rect 2405 -2200 2450 -2170
rect 2330 -2240 2450 -2200
rect 2330 -2270 2375 -2240
rect 2405 -2270 2450 -2240
rect 2330 -2310 2450 -2270
rect 2330 -2340 2375 -2310
rect 2405 -2340 2450 -2310
rect 2330 -2380 2450 -2340
rect 2330 -2410 2375 -2380
rect 2405 -2410 2450 -2380
rect 2330 -2445 2450 -2410
rect 2330 -2475 2375 -2445
rect 2405 -2475 2450 -2445
rect 2330 -2505 2450 -2475
rect 2330 -2535 2375 -2505
rect 2405 -2535 2450 -2505
rect 2330 -2570 2450 -2535
rect 2330 -2600 2375 -2570
rect 2405 -2600 2450 -2570
rect 2330 -2640 2450 -2600
rect 2330 -2670 2375 -2640
rect 2405 -2670 2450 -2640
rect 2330 -2710 2450 -2670
rect 2330 -2740 2375 -2710
rect 2405 -2740 2450 -2710
rect 2330 -2780 2450 -2740
rect 2330 -2810 2375 -2780
rect 2405 -2810 2450 -2780
rect 2330 -2845 2450 -2810
rect 2330 -2875 2375 -2845
rect 2405 -2875 2450 -2845
rect 2330 -2905 2450 -2875
rect 2330 -2935 2375 -2905
rect 2405 -2935 2450 -2905
rect 2330 -2970 2450 -2935
rect 2330 -3000 2375 -2970
rect 2405 -3000 2450 -2970
rect 2330 -3040 2450 -3000
rect 2330 -3070 2375 -3040
rect 2405 -3070 2450 -3040
rect 2330 -3110 2450 -3070
rect 2330 -3140 2375 -3110
rect 2405 -3140 2450 -3110
rect 2330 -3180 2450 -3140
rect 2330 -3210 2375 -3180
rect 2405 -3210 2450 -3180
rect 2330 -3245 2450 -3210
rect 2330 -3275 2375 -3245
rect 2405 -3275 2450 -3245
rect 2330 -3305 2450 -3275
rect 2330 -3335 2375 -3305
rect 2405 -3335 2450 -3305
rect 2330 -3370 2450 -3335
rect 2330 -3400 2375 -3370
rect 2405 -3400 2450 -3370
rect 2330 -3440 2450 -3400
rect 2330 -3470 2375 -3440
rect 2405 -3470 2450 -3440
rect 2330 -3510 2450 -3470
rect 2330 -3540 2375 -3510
rect 2405 -3540 2450 -3510
rect 2330 -3580 2450 -3540
rect 2330 -3610 2375 -3580
rect 2405 -3610 2450 -3580
rect 2330 -3645 2450 -3610
rect 2330 -3675 2375 -3645
rect 2405 -3675 2450 -3645
rect 2330 -3705 2450 -3675
rect 2330 -3735 2375 -3705
rect 2405 -3735 2450 -3705
rect 2330 -3770 2450 -3735
rect 2330 -3800 2375 -3770
rect 2405 -3800 2450 -3770
rect 2330 -3840 2450 -3800
rect 2330 -3870 2375 -3840
rect 2405 -3870 2450 -3840
rect 2330 -3910 2450 -3870
rect 2330 -3940 2375 -3910
rect 2405 -3940 2450 -3910
rect 2330 -3980 2450 -3940
rect 2330 -4010 2375 -3980
rect 2405 -4010 2450 -3980
rect 2330 -4045 2450 -4010
rect 2330 -4075 2375 -4045
rect 2405 -4075 2450 -4045
rect 2330 -4105 2450 -4075
rect 2330 -4135 2375 -4105
rect 2405 -4135 2450 -4105
rect 2330 -4170 2450 -4135
rect 2330 -4200 2375 -4170
rect 2405 -4200 2450 -4170
rect 2330 -4240 2450 -4200
rect 2330 -4270 2375 -4240
rect 2405 -4270 2450 -4240
rect 2330 -4310 2450 -4270
rect 2330 -4340 2375 -4310
rect 2405 -4340 2450 -4310
rect 2330 -4380 2450 -4340
rect 2330 -4410 2375 -4380
rect 2405 -4410 2450 -4380
rect 2330 -4445 2450 -4410
rect 2330 -4475 2375 -4445
rect 2405 -4475 2450 -4445
rect 2330 -4490 2450 -4475
rect 2680 -1305 2800 -1240
rect 2680 -1335 2725 -1305
rect 2755 -1335 2800 -1305
rect 2680 -1370 2800 -1335
rect 2680 -1400 2725 -1370
rect 2755 -1400 2800 -1370
rect 2680 -1440 2800 -1400
rect 2680 -1470 2725 -1440
rect 2755 -1470 2800 -1440
rect 2680 -1510 2800 -1470
rect 2680 -1540 2725 -1510
rect 2755 -1540 2800 -1510
rect 2680 -1580 2800 -1540
rect 2680 -1610 2725 -1580
rect 2755 -1610 2800 -1580
rect 2680 -1645 2800 -1610
rect 2680 -1675 2725 -1645
rect 2755 -1675 2800 -1645
rect 2680 -1705 2800 -1675
rect 2680 -1735 2725 -1705
rect 2755 -1735 2800 -1705
rect 2680 -1770 2800 -1735
rect 2680 -1800 2725 -1770
rect 2755 -1800 2800 -1770
rect 2680 -1840 2800 -1800
rect 2680 -1870 2725 -1840
rect 2755 -1870 2800 -1840
rect 2680 -1910 2800 -1870
rect 2680 -1940 2725 -1910
rect 2755 -1940 2800 -1910
rect 2680 -1980 2800 -1940
rect 2680 -2010 2725 -1980
rect 2755 -2010 2800 -1980
rect 2680 -2045 2800 -2010
rect 2680 -2075 2725 -2045
rect 2755 -2075 2800 -2045
rect 2680 -2105 2800 -2075
rect 2680 -2135 2725 -2105
rect 2755 -2135 2800 -2105
rect 2680 -2170 2800 -2135
rect 2680 -2200 2725 -2170
rect 2755 -2200 2800 -2170
rect 2680 -2240 2800 -2200
rect 2680 -2270 2725 -2240
rect 2755 -2270 2800 -2240
rect 2680 -2310 2800 -2270
rect 2680 -2340 2725 -2310
rect 2755 -2340 2800 -2310
rect 2680 -2380 2800 -2340
rect 2680 -2410 2725 -2380
rect 2755 -2410 2800 -2380
rect 2680 -2445 2800 -2410
rect 2680 -2475 2725 -2445
rect 2755 -2475 2800 -2445
rect 2680 -2505 2800 -2475
rect 2680 -2535 2725 -2505
rect 2755 -2535 2800 -2505
rect 2680 -2570 2800 -2535
rect 2680 -2600 2725 -2570
rect 2755 -2600 2800 -2570
rect 2680 -2640 2800 -2600
rect 2680 -2670 2725 -2640
rect 2755 -2670 2800 -2640
rect 2680 -2710 2800 -2670
rect 2680 -2740 2725 -2710
rect 2755 -2740 2800 -2710
rect 2680 -2780 2800 -2740
rect 2680 -2810 2725 -2780
rect 2755 -2810 2800 -2780
rect 2680 -2845 2800 -2810
rect 2680 -2875 2725 -2845
rect 2755 -2875 2800 -2845
rect 2680 -2905 2800 -2875
rect 2680 -2935 2725 -2905
rect 2755 -2935 2800 -2905
rect 2680 -2970 2800 -2935
rect 2680 -3000 2725 -2970
rect 2755 -3000 2800 -2970
rect 2680 -3040 2800 -3000
rect 2680 -3070 2725 -3040
rect 2755 -3070 2800 -3040
rect 2680 -3110 2800 -3070
rect 2680 -3140 2725 -3110
rect 2755 -3140 2800 -3110
rect 2680 -3180 2800 -3140
rect 2680 -3210 2725 -3180
rect 2755 -3210 2800 -3180
rect 2680 -3245 2800 -3210
rect 2680 -3275 2725 -3245
rect 2755 -3275 2800 -3245
rect 2680 -3305 2800 -3275
rect 2680 -3335 2725 -3305
rect 2755 -3335 2800 -3305
rect 2680 -3370 2800 -3335
rect 2680 -3400 2725 -3370
rect 2755 -3400 2800 -3370
rect 2680 -3440 2800 -3400
rect 2680 -3470 2725 -3440
rect 2755 -3470 2800 -3440
rect 2680 -3510 2800 -3470
rect 2680 -3540 2725 -3510
rect 2755 -3540 2800 -3510
rect 2680 -3580 2800 -3540
rect 2680 -3610 2725 -3580
rect 2755 -3610 2800 -3580
rect 2680 -3645 2800 -3610
rect 2680 -3675 2725 -3645
rect 2755 -3675 2800 -3645
rect 2680 -3705 2800 -3675
rect 2680 -3735 2725 -3705
rect 2755 -3735 2800 -3705
rect 2680 -3770 2800 -3735
rect 2680 -3800 2725 -3770
rect 2755 -3800 2800 -3770
rect 2680 -3840 2800 -3800
rect 2680 -3870 2725 -3840
rect 2755 -3870 2800 -3840
rect 2680 -3910 2800 -3870
rect 2680 -3940 2725 -3910
rect 2755 -3940 2800 -3910
rect 2680 -3980 2800 -3940
rect 2680 -4010 2725 -3980
rect 2755 -4010 2800 -3980
rect 2680 -4045 2800 -4010
rect 2680 -4075 2725 -4045
rect 2755 -4075 2800 -4045
rect 2680 -4105 2800 -4075
rect 2680 -4135 2725 -4105
rect 2755 -4135 2800 -4105
rect 2680 -4170 2800 -4135
rect 2680 -4200 2725 -4170
rect 2755 -4200 2800 -4170
rect 2680 -4240 2800 -4200
rect 2680 -4270 2725 -4240
rect 2755 -4270 2800 -4240
rect 2680 -4310 2800 -4270
rect 2680 -4340 2725 -4310
rect 2755 -4340 2800 -4310
rect 2680 -4380 2800 -4340
rect 2680 -4410 2725 -4380
rect 2755 -4410 2800 -4380
rect 2680 -4445 2800 -4410
rect 2680 -4475 2725 -4445
rect 2755 -4475 2800 -4445
rect 2680 -4490 2800 -4475
rect 3030 -1305 3150 -1240
rect 3030 -1335 3075 -1305
rect 3105 -1335 3150 -1305
rect 3030 -1370 3150 -1335
rect 3030 -1400 3075 -1370
rect 3105 -1400 3150 -1370
rect 3030 -1440 3150 -1400
rect 3030 -1470 3075 -1440
rect 3105 -1470 3150 -1440
rect 3030 -1510 3150 -1470
rect 3030 -1540 3075 -1510
rect 3105 -1540 3150 -1510
rect 3030 -1580 3150 -1540
rect 3030 -1610 3075 -1580
rect 3105 -1610 3150 -1580
rect 3030 -1645 3150 -1610
rect 3030 -1675 3075 -1645
rect 3105 -1675 3150 -1645
rect 3030 -1705 3150 -1675
rect 3030 -1735 3075 -1705
rect 3105 -1735 3150 -1705
rect 3030 -1770 3150 -1735
rect 3030 -1800 3075 -1770
rect 3105 -1800 3150 -1770
rect 3030 -1840 3150 -1800
rect 3030 -1870 3075 -1840
rect 3105 -1870 3150 -1840
rect 3030 -1910 3150 -1870
rect 3030 -1940 3075 -1910
rect 3105 -1940 3150 -1910
rect 3030 -1980 3150 -1940
rect 3030 -2010 3075 -1980
rect 3105 -2010 3150 -1980
rect 3030 -2045 3150 -2010
rect 3030 -2075 3075 -2045
rect 3105 -2075 3150 -2045
rect 3030 -2105 3150 -2075
rect 3030 -2135 3075 -2105
rect 3105 -2135 3150 -2105
rect 3030 -2170 3150 -2135
rect 3030 -2200 3075 -2170
rect 3105 -2200 3150 -2170
rect 3030 -2240 3150 -2200
rect 3030 -2270 3075 -2240
rect 3105 -2270 3150 -2240
rect 3030 -2310 3150 -2270
rect 3030 -2340 3075 -2310
rect 3105 -2340 3150 -2310
rect 3030 -2380 3150 -2340
rect 3030 -2410 3075 -2380
rect 3105 -2410 3150 -2380
rect 3030 -2445 3150 -2410
rect 3030 -2475 3075 -2445
rect 3105 -2475 3150 -2445
rect 3030 -2505 3150 -2475
rect 3030 -2535 3075 -2505
rect 3105 -2535 3150 -2505
rect 3030 -2570 3150 -2535
rect 3030 -2600 3075 -2570
rect 3105 -2600 3150 -2570
rect 3030 -2640 3150 -2600
rect 3030 -2670 3075 -2640
rect 3105 -2670 3150 -2640
rect 3030 -2710 3150 -2670
rect 3030 -2740 3075 -2710
rect 3105 -2740 3150 -2710
rect 3030 -2780 3150 -2740
rect 3030 -2810 3075 -2780
rect 3105 -2810 3150 -2780
rect 3030 -2845 3150 -2810
rect 3030 -2875 3075 -2845
rect 3105 -2875 3150 -2845
rect 3030 -2905 3150 -2875
rect 3030 -2935 3075 -2905
rect 3105 -2935 3150 -2905
rect 3030 -2970 3150 -2935
rect 3030 -3000 3075 -2970
rect 3105 -3000 3150 -2970
rect 3030 -3040 3150 -3000
rect 3030 -3070 3075 -3040
rect 3105 -3070 3150 -3040
rect 3030 -3110 3150 -3070
rect 3030 -3140 3075 -3110
rect 3105 -3140 3150 -3110
rect 3030 -3180 3150 -3140
rect 3030 -3210 3075 -3180
rect 3105 -3210 3150 -3180
rect 3030 -3245 3150 -3210
rect 3030 -3275 3075 -3245
rect 3105 -3275 3150 -3245
rect 3030 -3305 3150 -3275
rect 3030 -3335 3075 -3305
rect 3105 -3335 3150 -3305
rect 3030 -3370 3150 -3335
rect 3030 -3400 3075 -3370
rect 3105 -3400 3150 -3370
rect 3030 -3440 3150 -3400
rect 3030 -3470 3075 -3440
rect 3105 -3470 3150 -3440
rect 3030 -3510 3150 -3470
rect 3030 -3540 3075 -3510
rect 3105 -3540 3150 -3510
rect 3030 -3580 3150 -3540
rect 3030 -3610 3075 -3580
rect 3105 -3610 3150 -3580
rect 3030 -3645 3150 -3610
rect 3030 -3675 3075 -3645
rect 3105 -3675 3150 -3645
rect 3030 -3705 3150 -3675
rect 3030 -3735 3075 -3705
rect 3105 -3735 3150 -3705
rect 3030 -3770 3150 -3735
rect 3030 -3800 3075 -3770
rect 3105 -3800 3150 -3770
rect 3030 -3840 3150 -3800
rect 3030 -3870 3075 -3840
rect 3105 -3870 3150 -3840
rect 3030 -3910 3150 -3870
rect 3030 -3940 3075 -3910
rect 3105 -3940 3150 -3910
rect 3030 -3980 3150 -3940
rect 3030 -4010 3075 -3980
rect 3105 -4010 3150 -3980
rect 3030 -4045 3150 -4010
rect 3030 -4075 3075 -4045
rect 3105 -4075 3150 -4045
rect 3030 -4105 3150 -4075
rect 3030 -4135 3075 -4105
rect 3105 -4135 3150 -4105
rect 3030 -4170 3150 -4135
rect 3030 -4200 3075 -4170
rect 3105 -4200 3150 -4170
rect 3030 -4240 3150 -4200
rect 3030 -4270 3075 -4240
rect 3105 -4270 3150 -4240
rect 3030 -4310 3150 -4270
rect 3030 -4340 3075 -4310
rect 3105 -4340 3150 -4310
rect 3030 -4380 3150 -4340
rect 3030 -4410 3075 -4380
rect 3105 -4410 3150 -4380
rect 3030 -4445 3150 -4410
rect 3030 -4475 3075 -4445
rect 3105 -4475 3150 -4445
rect 3030 -4490 3150 -4475
rect 3380 -1305 3500 -1240
rect 3380 -1335 3425 -1305
rect 3455 -1335 3500 -1305
rect 3380 -1370 3500 -1335
rect 3380 -1400 3425 -1370
rect 3455 -1400 3500 -1370
rect 3380 -1440 3500 -1400
rect 3380 -1470 3425 -1440
rect 3455 -1470 3500 -1440
rect 3380 -1510 3500 -1470
rect 3380 -1540 3425 -1510
rect 3455 -1540 3500 -1510
rect 3380 -1580 3500 -1540
rect 3380 -1610 3425 -1580
rect 3455 -1610 3500 -1580
rect 3380 -1645 3500 -1610
rect 3380 -1675 3425 -1645
rect 3455 -1675 3500 -1645
rect 3380 -1705 3500 -1675
rect 3380 -1735 3425 -1705
rect 3455 -1735 3500 -1705
rect 3380 -1770 3500 -1735
rect 3380 -1800 3425 -1770
rect 3455 -1800 3500 -1770
rect 3380 -1840 3500 -1800
rect 3380 -1870 3425 -1840
rect 3455 -1870 3500 -1840
rect 3380 -1910 3500 -1870
rect 3380 -1940 3425 -1910
rect 3455 -1940 3500 -1910
rect 3380 -1980 3500 -1940
rect 3380 -2010 3425 -1980
rect 3455 -2010 3500 -1980
rect 3380 -2045 3500 -2010
rect 3380 -2075 3425 -2045
rect 3455 -2075 3500 -2045
rect 3380 -2105 3500 -2075
rect 3380 -2135 3425 -2105
rect 3455 -2135 3500 -2105
rect 3380 -2170 3500 -2135
rect 3380 -2200 3425 -2170
rect 3455 -2200 3500 -2170
rect 3380 -2240 3500 -2200
rect 3380 -2270 3425 -2240
rect 3455 -2270 3500 -2240
rect 3380 -2310 3500 -2270
rect 3380 -2340 3425 -2310
rect 3455 -2340 3500 -2310
rect 3380 -2380 3500 -2340
rect 3380 -2410 3425 -2380
rect 3455 -2410 3500 -2380
rect 3380 -2445 3500 -2410
rect 3380 -2475 3425 -2445
rect 3455 -2475 3500 -2445
rect 3380 -2505 3500 -2475
rect 3380 -2535 3425 -2505
rect 3455 -2535 3500 -2505
rect 3380 -2570 3500 -2535
rect 3380 -2600 3425 -2570
rect 3455 -2600 3500 -2570
rect 3380 -2640 3500 -2600
rect 3380 -2670 3425 -2640
rect 3455 -2670 3500 -2640
rect 3380 -2710 3500 -2670
rect 3380 -2740 3425 -2710
rect 3455 -2740 3500 -2710
rect 3380 -2780 3500 -2740
rect 3380 -2810 3425 -2780
rect 3455 -2810 3500 -2780
rect 3380 -2845 3500 -2810
rect 3380 -2875 3425 -2845
rect 3455 -2875 3500 -2845
rect 3380 -2905 3500 -2875
rect 3380 -2935 3425 -2905
rect 3455 -2935 3500 -2905
rect 3380 -2970 3500 -2935
rect 3380 -3000 3425 -2970
rect 3455 -3000 3500 -2970
rect 3380 -3040 3500 -3000
rect 3380 -3070 3425 -3040
rect 3455 -3070 3500 -3040
rect 3380 -3110 3500 -3070
rect 3380 -3140 3425 -3110
rect 3455 -3140 3500 -3110
rect 3380 -3180 3500 -3140
rect 3380 -3210 3425 -3180
rect 3455 -3210 3500 -3180
rect 3380 -3245 3500 -3210
rect 3380 -3275 3425 -3245
rect 3455 -3275 3500 -3245
rect 3380 -3305 3500 -3275
rect 3380 -3335 3425 -3305
rect 3455 -3335 3500 -3305
rect 3380 -3370 3500 -3335
rect 3380 -3400 3425 -3370
rect 3455 -3400 3500 -3370
rect 3380 -3440 3500 -3400
rect 3380 -3470 3425 -3440
rect 3455 -3470 3500 -3440
rect 3380 -3510 3500 -3470
rect 3380 -3540 3425 -3510
rect 3455 -3540 3500 -3510
rect 3380 -3580 3500 -3540
rect 3380 -3610 3425 -3580
rect 3455 -3610 3500 -3580
rect 3380 -3645 3500 -3610
rect 3380 -3675 3425 -3645
rect 3455 -3675 3500 -3645
rect 3380 -3705 3500 -3675
rect 3380 -3735 3425 -3705
rect 3455 -3735 3500 -3705
rect 3380 -3770 3500 -3735
rect 3380 -3800 3425 -3770
rect 3455 -3800 3500 -3770
rect 3380 -3840 3500 -3800
rect 3380 -3870 3425 -3840
rect 3455 -3870 3500 -3840
rect 3380 -3910 3500 -3870
rect 3380 -3940 3425 -3910
rect 3455 -3940 3500 -3910
rect 3380 -3980 3500 -3940
rect 3380 -4010 3425 -3980
rect 3455 -4010 3500 -3980
rect 3380 -4045 3500 -4010
rect 3380 -4075 3425 -4045
rect 3455 -4075 3500 -4045
rect 3380 -4105 3500 -4075
rect 3380 -4135 3425 -4105
rect 3455 -4135 3500 -4105
rect 3380 -4170 3500 -4135
rect 3380 -4200 3425 -4170
rect 3455 -4200 3500 -4170
rect 3380 -4240 3500 -4200
rect 3380 -4270 3425 -4240
rect 3455 -4270 3500 -4240
rect 3380 -4310 3500 -4270
rect 3380 -4340 3425 -4310
rect 3455 -4340 3500 -4310
rect 3380 -4380 3500 -4340
rect 3380 -4410 3425 -4380
rect 3455 -4410 3500 -4380
rect 3380 -4445 3500 -4410
rect 3380 -4475 3425 -4445
rect 3455 -4475 3500 -4445
rect 3380 -4490 3500 -4475
rect 3730 -1305 3850 -1240
rect 3730 -1335 3775 -1305
rect 3805 -1335 3850 -1305
rect 3730 -1370 3850 -1335
rect 3730 -1400 3775 -1370
rect 3805 -1400 3850 -1370
rect 3730 -1440 3850 -1400
rect 3730 -1470 3775 -1440
rect 3805 -1470 3850 -1440
rect 3730 -1510 3850 -1470
rect 3730 -1540 3775 -1510
rect 3805 -1540 3850 -1510
rect 3730 -1580 3850 -1540
rect 3730 -1610 3775 -1580
rect 3805 -1610 3850 -1580
rect 3730 -1645 3850 -1610
rect 3730 -1675 3775 -1645
rect 3805 -1675 3850 -1645
rect 3730 -1705 3850 -1675
rect 3730 -1735 3775 -1705
rect 3805 -1735 3850 -1705
rect 3730 -1770 3850 -1735
rect 3730 -1800 3775 -1770
rect 3805 -1800 3850 -1770
rect 3730 -1840 3850 -1800
rect 3730 -1870 3775 -1840
rect 3805 -1870 3850 -1840
rect 3730 -1910 3850 -1870
rect 3730 -1940 3775 -1910
rect 3805 -1940 3850 -1910
rect 3730 -1980 3850 -1940
rect 3730 -2010 3775 -1980
rect 3805 -2010 3850 -1980
rect 3730 -2045 3850 -2010
rect 3730 -2075 3775 -2045
rect 3805 -2075 3850 -2045
rect 3730 -2105 3850 -2075
rect 3730 -2135 3775 -2105
rect 3805 -2135 3850 -2105
rect 3730 -2170 3850 -2135
rect 3730 -2200 3775 -2170
rect 3805 -2200 3850 -2170
rect 3730 -2240 3850 -2200
rect 3730 -2270 3775 -2240
rect 3805 -2270 3850 -2240
rect 3730 -2310 3850 -2270
rect 3730 -2340 3775 -2310
rect 3805 -2340 3850 -2310
rect 3730 -2380 3850 -2340
rect 3730 -2410 3775 -2380
rect 3805 -2410 3850 -2380
rect 3730 -2445 3850 -2410
rect 3730 -2475 3775 -2445
rect 3805 -2475 3850 -2445
rect 3730 -2505 3850 -2475
rect 3730 -2535 3775 -2505
rect 3805 -2535 3850 -2505
rect 3730 -2570 3850 -2535
rect 3730 -2600 3775 -2570
rect 3805 -2600 3850 -2570
rect 3730 -2640 3850 -2600
rect 3730 -2670 3775 -2640
rect 3805 -2670 3850 -2640
rect 3730 -2710 3850 -2670
rect 3730 -2740 3775 -2710
rect 3805 -2740 3850 -2710
rect 3730 -2780 3850 -2740
rect 3730 -2810 3775 -2780
rect 3805 -2810 3850 -2780
rect 3730 -2845 3850 -2810
rect 3730 -2875 3775 -2845
rect 3805 -2875 3850 -2845
rect 3730 -2905 3850 -2875
rect 3730 -2935 3775 -2905
rect 3805 -2935 3850 -2905
rect 3730 -2970 3850 -2935
rect 3730 -3000 3775 -2970
rect 3805 -3000 3850 -2970
rect 3730 -3040 3850 -3000
rect 3730 -3070 3775 -3040
rect 3805 -3070 3850 -3040
rect 3730 -3110 3850 -3070
rect 3730 -3140 3775 -3110
rect 3805 -3140 3850 -3110
rect 3730 -3180 3850 -3140
rect 3730 -3210 3775 -3180
rect 3805 -3210 3850 -3180
rect 3730 -3245 3850 -3210
rect 3730 -3275 3775 -3245
rect 3805 -3275 3850 -3245
rect 3730 -3305 3850 -3275
rect 3730 -3335 3775 -3305
rect 3805 -3335 3850 -3305
rect 3730 -3370 3850 -3335
rect 3730 -3400 3775 -3370
rect 3805 -3400 3850 -3370
rect 3730 -3440 3850 -3400
rect 3730 -3470 3775 -3440
rect 3805 -3470 3850 -3440
rect 3730 -3510 3850 -3470
rect 3730 -3540 3775 -3510
rect 3805 -3540 3850 -3510
rect 3730 -3580 3850 -3540
rect 3730 -3610 3775 -3580
rect 3805 -3610 3850 -3580
rect 3730 -3645 3850 -3610
rect 3730 -3675 3775 -3645
rect 3805 -3675 3850 -3645
rect 3730 -3705 3850 -3675
rect 3730 -3735 3775 -3705
rect 3805 -3735 3850 -3705
rect 3730 -3770 3850 -3735
rect 3730 -3800 3775 -3770
rect 3805 -3800 3850 -3770
rect 3730 -3840 3850 -3800
rect 3730 -3870 3775 -3840
rect 3805 -3870 3850 -3840
rect 3730 -3910 3850 -3870
rect 3730 -3940 3775 -3910
rect 3805 -3940 3850 -3910
rect 3730 -3980 3850 -3940
rect 3730 -4010 3775 -3980
rect 3805 -4010 3850 -3980
rect 3730 -4045 3850 -4010
rect 3730 -4075 3775 -4045
rect 3805 -4075 3850 -4045
rect 3730 -4105 3850 -4075
rect 3730 -4135 3775 -4105
rect 3805 -4135 3850 -4105
rect 3730 -4170 3850 -4135
rect 3730 -4200 3775 -4170
rect 3805 -4200 3850 -4170
rect 3730 -4240 3850 -4200
rect 3730 -4270 3775 -4240
rect 3805 -4270 3850 -4240
rect 3730 -4310 3850 -4270
rect 3730 -4340 3775 -4310
rect 3805 -4340 3850 -4310
rect 3730 -4380 3850 -4340
rect 3730 -4410 3775 -4380
rect 3805 -4410 3850 -4380
rect 3730 -4445 3850 -4410
rect 3730 -4475 3775 -4445
rect 3805 -4475 3850 -4445
rect 3730 -4490 3850 -4475
rect 4080 -1305 4200 -1240
rect 4080 -1335 4125 -1305
rect 4155 -1335 4200 -1305
rect 4080 -1370 4200 -1335
rect 4080 -1400 4125 -1370
rect 4155 -1400 4200 -1370
rect 4080 -1440 4200 -1400
rect 4080 -1470 4125 -1440
rect 4155 -1470 4200 -1440
rect 4080 -1510 4200 -1470
rect 4080 -1540 4125 -1510
rect 4155 -1540 4200 -1510
rect 4080 -1580 4200 -1540
rect 4080 -1610 4125 -1580
rect 4155 -1610 4200 -1580
rect 4080 -1645 4200 -1610
rect 4080 -1675 4125 -1645
rect 4155 -1675 4200 -1645
rect 4080 -1705 4200 -1675
rect 4080 -1735 4125 -1705
rect 4155 -1735 4200 -1705
rect 4080 -1770 4200 -1735
rect 4080 -1800 4125 -1770
rect 4155 -1800 4200 -1770
rect 4080 -1840 4200 -1800
rect 4080 -1870 4125 -1840
rect 4155 -1870 4200 -1840
rect 4080 -1910 4200 -1870
rect 4080 -1940 4125 -1910
rect 4155 -1940 4200 -1910
rect 4080 -1980 4200 -1940
rect 4080 -2010 4125 -1980
rect 4155 -2010 4200 -1980
rect 4080 -2045 4200 -2010
rect 4080 -2075 4125 -2045
rect 4155 -2075 4200 -2045
rect 4080 -2105 4200 -2075
rect 4080 -2135 4125 -2105
rect 4155 -2135 4200 -2105
rect 4080 -2170 4200 -2135
rect 4080 -2200 4125 -2170
rect 4155 -2200 4200 -2170
rect 4080 -2240 4200 -2200
rect 4080 -2270 4125 -2240
rect 4155 -2270 4200 -2240
rect 4080 -2310 4200 -2270
rect 4080 -2340 4125 -2310
rect 4155 -2340 4200 -2310
rect 4080 -2380 4200 -2340
rect 4080 -2410 4125 -2380
rect 4155 -2410 4200 -2380
rect 4080 -2445 4200 -2410
rect 4080 -2475 4125 -2445
rect 4155 -2475 4200 -2445
rect 4080 -2505 4200 -2475
rect 4080 -2535 4125 -2505
rect 4155 -2535 4200 -2505
rect 4080 -2570 4200 -2535
rect 4080 -2600 4125 -2570
rect 4155 -2600 4200 -2570
rect 4080 -2640 4200 -2600
rect 4080 -2670 4125 -2640
rect 4155 -2670 4200 -2640
rect 4080 -2710 4200 -2670
rect 4080 -2740 4125 -2710
rect 4155 -2740 4200 -2710
rect 4080 -2780 4200 -2740
rect 4080 -2810 4125 -2780
rect 4155 -2810 4200 -2780
rect 4080 -2845 4200 -2810
rect 4080 -2875 4125 -2845
rect 4155 -2875 4200 -2845
rect 4080 -2905 4200 -2875
rect 4080 -2935 4125 -2905
rect 4155 -2935 4200 -2905
rect 4080 -2970 4200 -2935
rect 4080 -3000 4125 -2970
rect 4155 -3000 4200 -2970
rect 4080 -3040 4200 -3000
rect 4080 -3070 4125 -3040
rect 4155 -3070 4200 -3040
rect 4080 -3110 4200 -3070
rect 4080 -3140 4125 -3110
rect 4155 -3140 4200 -3110
rect 4080 -3180 4200 -3140
rect 4080 -3210 4125 -3180
rect 4155 -3210 4200 -3180
rect 4080 -3245 4200 -3210
rect 4080 -3275 4125 -3245
rect 4155 -3275 4200 -3245
rect 4080 -3305 4200 -3275
rect 4080 -3335 4125 -3305
rect 4155 -3335 4200 -3305
rect 4080 -3370 4200 -3335
rect 4080 -3400 4125 -3370
rect 4155 -3400 4200 -3370
rect 4080 -3440 4200 -3400
rect 4080 -3470 4125 -3440
rect 4155 -3470 4200 -3440
rect 4080 -3510 4200 -3470
rect 4080 -3540 4125 -3510
rect 4155 -3540 4200 -3510
rect 4080 -3580 4200 -3540
rect 4080 -3610 4125 -3580
rect 4155 -3610 4200 -3580
rect 4080 -3645 4200 -3610
rect 4080 -3675 4125 -3645
rect 4155 -3675 4200 -3645
rect 4080 -3705 4200 -3675
rect 4080 -3735 4125 -3705
rect 4155 -3735 4200 -3705
rect 4080 -3770 4200 -3735
rect 4080 -3800 4125 -3770
rect 4155 -3800 4200 -3770
rect 4080 -3840 4200 -3800
rect 4080 -3870 4125 -3840
rect 4155 -3870 4200 -3840
rect 4080 -3910 4200 -3870
rect 4080 -3940 4125 -3910
rect 4155 -3940 4200 -3910
rect 4080 -3980 4200 -3940
rect 4080 -4010 4125 -3980
rect 4155 -4010 4200 -3980
rect 4080 -4045 4200 -4010
rect 4080 -4075 4125 -4045
rect 4155 -4075 4200 -4045
rect 4080 -4105 4200 -4075
rect 4080 -4135 4125 -4105
rect 4155 -4135 4200 -4105
rect 4080 -4170 4200 -4135
rect 4080 -4200 4125 -4170
rect 4155 -4200 4200 -4170
rect 4080 -4240 4200 -4200
rect 4080 -4270 4125 -4240
rect 4155 -4270 4200 -4240
rect 4080 -4310 4200 -4270
rect 4080 -4340 4125 -4310
rect 4155 -4340 4200 -4310
rect 4080 -4380 4200 -4340
rect 4080 -4410 4125 -4380
rect 4155 -4410 4200 -4380
rect 4080 -4445 4200 -4410
rect 4080 -4475 4125 -4445
rect 4155 -4475 4200 -4445
rect 4080 -4490 4200 -4475
rect 4430 -1305 4550 -1240
rect 4430 -1335 4475 -1305
rect 4505 -1335 4550 -1305
rect 4430 -1370 4550 -1335
rect 4430 -1400 4475 -1370
rect 4505 -1400 4550 -1370
rect 4430 -1440 4550 -1400
rect 4430 -1470 4475 -1440
rect 4505 -1470 4550 -1440
rect 4430 -1510 4550 -1470
rect 4430 -1540 4475 -1510
rect 4505 -1540 4550 -1510
rect 4430 -1580 4550 -1540
rect 4430 -1610 4475 -1580
rect 4505 -1610 4550 -1580
rect 4430 -1645 4550 -1610
rect 4430 -1675 4475 -1645
rect 4505 -1675 4550 -1645
rect 4430 -1705 4550 -1675
rect 4430 -1735 4475 -1705
rect 4505 -1735 4550 -1705
rect 4430 -1770 4550 -1735
rect 4430 -1800 4475 -1770
rect 4505 -1800 4550 -1770
rect 4430 -1840 4550 -1800
rect 4430 -1870 4475 -1840
rect 4505 -1870 4550 -1840
rect 4430 -1910 4550 -1870
rect 4430 -1940 4475 -1910
rect 4505 -1940 4550 -1910
rect 4430 -1980 4550 -1940
rect 4430 -2010 4475 -1980
rect 4505 -2010 4550 -1980
rect 4430 -2045 4550 -2010
rect 4430 -2075 4475 -2045
rect 4505 -2075 4550 -2045
rect 4430 -2105 4550 -2075
rect 4430 -2135 4475 -2105
rect 4505 -2135 4550 -2105
rect 4430 -2170 4550 -2135
rect 4430 -2200 4475 -2170
rect 4505 -2200 4550 -2170
rect 4430 -2240 4550 -2200
rect 4430 -2270 4475 -2240
rect 4505 -2270 4550 -2240
rect 4430 -2310 4550 -2270
rect 4430 -2340 4475 -2310
rect 4505 -2340 4550 -2310
rect 4430 -2380 4550 -2340
rect 4430 -2410 4475 -2380
rect 4505 -2410 4550 -2380
rect 4430 -2445 4550 -2410
rect 4430 -2475 4475 -2445
rect 4505 -2475 4550 -2445
rect 4430 -2505 4550 -2475
rect 4430 -2535 4475 -2505
rect 4505 -2535 4550 -2505
rect 4430 -2570 4550 -2535
rect 4430 -2600 4475 -2570
rect 4505 -2600 4550 -2570
rect 4430 -2640 4550 -2600
rect 4430 -2670 4475 -2640
rect 4505 -2670 4550 -2640
rect 4430 -2710 4550 -2670
rect 4430 -2740 4475 -2710
rect 4505 -2740 4550 -2710
rect 4430 -2780 4550 -2740
rect 4430 -2810 4475 -2780
rect 4505 -2810 4550 -2780
rect 4430 -2845 4550 -2810
rect 4430 -2875 4475 -2845
rect 4505 -2875 4550 -2845
rect 4430 -2905 4550 -2875
rect 4430 -2935 4475 -2905
rect 4505 -2935 4550 -2905
rect 4430 -2970 4550 -2935
rect 4430 -3000 4475 -2970
rect 4505 -3000 4550 -2970
rect 4430 -3040 4550 -3000
rect 4430 -3070 4475 -3040
rect 4505 -3070 4550 -3040
rect 4430 -3110 4550 -3070
rect 4430 -3140 4475 -3110
rect 4505 -3140 4550 -3110
rect 4430 -3180 4550 -3140
rect 4430 -3210 4475 -3180
rect 4505 -3210 4550 -3180
rect 4430 -3245 4550 -3210
rect 4430 -3275 4475 -3245
rect 4505 -3275 4550 -3245
rect 4430 -3305 4550 -3275
rect 4430 -3335 4475 -3305
rect 4505 -3335 4550 -3305
rect 4430 -3370 4550 -3335
rect 4430 -3400 4475 -3370
rect 4505 -3400 4550 -3370
rect 4430 -3440 4550 -3400
rect 4430 -3470 4475 -3440
rect 4505 -3470 4550 -3440
rect 4430 -3510 4550 -3470
rect 4430 -3540 4475 -3510
rect 4505 -3540 4550 -3510
rect 4430 -3580 4550 -3540
rect 4430 -3610 4475 -3580
rect 4505 -3610 4550 -3580
rect 4430 -3645 4550 -3610
rect 4430 -3675 4475 -3645
rect 4505 -3675 4550 -3645
rect 4430 -3705 4550 -3675
rect 4430 -3735 4475 -3705
rect 4505 -3735 4550 -3705
rect 4430 -3770 4550 -3735
rect 4430 -3800 4475 -3770
rect 4505 -3800 4550 -3770
rect 4430 -3840 4550 -3800
rect 4430 -3870 4475 -3840
rect 4505 -3870 4550 -3840
rect 4430 -3910 4550 -3870
rect 4430 -3940 4475 -3910
rect 4505 -3940 4550 -3910
rect 4430 -3980 4550 -3940
rect 4430 -4010 4475 -3980
rect 4505 -4010 4550 -3980
rect 4430 -4045 4550 -4010
rect 4430 -4075 4475 -4045
rect 4505 -4075 4550 -4045
rect 4430 -4105 4550 -4075
rect 4430 -4135 4475 -4105
rect 4505 -4135 4550 -4105
rect 4430 -4170 4550 -4135
rect 4430 -4200 4475 -4170
rect 4505 -4200 4550 -4170
rect 4430 -4240 4550 -4200
rect 4430 -4270 4475 -4240
rect 4505 -4270 4550 -4240
rect 4430 -4310 4550 -4270
rect 4430 -4340 4475 -4310
rect 4505 -4340 4550 -4310
rect 4430 -4380 4550 -4340
rect 4430 -4410 4475 -4380
rect 4505 -4410 4550 -4380
rect 4430 -4445 4550 -4410
rect 4430 -4475 4475 -4445
rect 4505 -4475 4550 -4445
rect 4430 -4490 4550 -4475
rect 4780 -1305 4900 -1240
rect 4780 -1335 4825 -1305
rect 4855 -1335 4900 -1305
rect 4780 -1370 4900 -1335
rect 4780 -1400 4825 -1370
rect 4855 -1400 4900 -1370
rect 4780 -1440 4900 -1400
rect 4780 -1470 4825 -1440
rect 4855 -1470 4900 -1440
rect 4780 -1510 4900 -1470
rect 4780 -1540 4825 -1510
rect 4855 -1540 4900 -1510
rect 4780 -1580 4900 -1540
rect 4780 -1610 4825 -1580
rect 4855 -1610 4900 -1580
rect 4780 -1645 4900 -1610
rect 4780 -1675 4825 -1645
rect 4855 -1675 4900 -1645
rect 4780 -1705 4900 -1675
rect 4780 -1735 4825 -1705
rect 4855 -1735 4900 -1705
rect 4780 -1770 4900 -1735
rect 4780 -1800 4825 -1770
rect 4855 -1800 4900 -1770
rect 4780 -1840 4900 -1800
rect 4780 -1870 4825 -1840
rect 4855 -1870 4900 -1840
rect 4780 -1910 4900 -1870
rect 4780 -1940 4825 -1910
rect 4855 -1940 4900 -1910
rect 4780 -1980 4900 -1940
rect 4780 -2010 4825 -1980
rect 4855 -2010 4900 -1980
rect 4780 -2045 4900 -2010
rect 4780 -2075 4825 -2045
rect 4855 -2075 4900 -2045
rect 4780 -2105 4900 -2075
rect 4780 -2135 4825 -2105
rect 4855 -2135 4900 -2105
rect 4780 -2170 4900 -2135
rect 4780 -2200 4825 -2170
rect 4855 -2200 4900 -2170
rect 4780 -2240 4900 -2200
rect 4780 -2270 4825 -2240
rect 4855 -2270 4900 -2240
rect 4780 -2310 4900 -2270
rect 4780 -2340 4825 -2310
rect 4855 -2340 4900 -2310
rect 4780 -2380 4900 -2340
rect 4780 -2410 4825 -2380
rect 4855 -2410 4900 -2380
rect 4780 -2445 4900 -2410
rect 4780 -2475 4825 -2445
rect 4855 -2475 4900 -2445
rect 4780 -2505 4900 -2475
rect 4780 -2535 4825 -2505
rect 4855 -2535 4900 -2505
rect 4780 -2570 4900 -2535
rect 4780 -2600 4825 -2570
rect 4855 -2600 4900 -2570
rect 4780 -2640 4900 -2600
rect 4780 -2670 4825 -2640
rect 4855 -2670 4900 -2640
rect 4780 -2710 4900 -2670
rect 4780 -2740 4825 -2710
rect 4855 -2740 4900 -2710
rect 4780 -2780 4900 -2740
rect 4780 -2810 4825 -2780
rect 4855 -2810 4900 -2780
rect 4780 -2845 4900 -2810
rect 4780 -2875 4825 -2845
rect 4855 -2875 4900 -2845
rect 4780 -2905 4900 -2875
rect 4780 -2935 4825 -2905
rect 4855 -2935 4900 -2905
rect 4780 -2970 4900 -2935
rect 4780 -3000 4825 -2970
rect 4855 -3000 4900 -2970
rect 4780 -3040 4900 -3000
rect 4780 -3070 4825 -3040
rect 4855 -3070 4900 -3040
rect 4780 -3110 4900 -3070
rect 4780 -3140 4825 -3110
rect 4855 -3140 4900 -3110
rect 4780 -3180 4900 -3140
rect 4780 -3210 4825 -3180
rect 4855 -3210 4900 -3180
rect 4780 -3245 4900 -3210
rect 4780 -3275 4825 -3245
rect 4855 -3275 4900 -3245
rect 4780 -3305 4900 -3275
rect 4780 -3335 4825 -3305
rect 4855 -3335 4900 -3305
rect 4780 -3370 4900 -3335
rect 4780 -3400 4825 -3370
rect 4855 -3400 4900 -3370
rect 4780 -3440 4900 -3400
rect 4780 -3470 4825 -3440
rect 4855 -3470 4900 -3440
rect 4780 -3510 4900 -3470
rect 4780 -3540 4825 -3510
rect 4855 -3540 4900 -3510
rect 4780 -3580 4900 -3540
rect 4780 -3610 4825 -3580
rect 4855 -3610 4900 -3580
rect 4780 -3645 4900 -3610
rect 4780 -3675 4825 -3645
rect 4855 -3675 4900 -3645
rect 4780 -3705 4900 -3675
rect 4780 -3735 4825 -3705
rect 4855 -3735 4900 -3705
rect 4780 -3770 4900 -3735
rect 4780 -3800 4825 -3770
rect 4855 -3800 4900 -3770
rect 4780 -3840 4900 -3800
rect 4780 -3870 4825 -3840
rect 4855 -3870 4900 -3840
rect 4780 -3910 4900 -3870
rect 4780 -3940 4825 -3910
rect 4855 -3940 4900 -3910
rect 4780 -3980 4900 -3940
rect 4780 -4010 4825 -3980
rect 4855 -4010 4900 -3980
rect 4780 -4045 4900 -4010
rect 4780 -4075 4825 -4045
rect 4855 -4075 4900 -4045
rect 4780 -4105 4900 -4075
rect 4780 -4135 4825 -4105
rect 4855 -4135 4900 -4105
rect 4780 -4170 4900 -4135
rect 4780 -4200 4825 -4170
rect 4855 -4200 4900 -4170
rect 4780 -4240 4900 -4200
rect 4780 -4270 4825 -4240
rect 4855 -4270 4900 -4240
rect 4780 -4310 4900 -4270
rect 4780 -4340 4825 -4310
rect 4855 -4340 4900 -4310
rect 4780 -4380 4900 -4340
rect 4780 -4410 4825 -4380
rect 4855 -4410 4900 -4380
rect 4780 -4445 4900 -4410
rect 4780 -4475 4825 -4445
rect 4855 -4475 4900 -4445
rect 4780 -4490 4900 -4475
rect 5130 -1305 5250 -1240
rect 5130 -1335 5175 -1305
rect 5205 -1335 5250 -1305
rect 5130 -1370 5250 -1335
rect 5130 -1400 5175 -1370
rect 5205 -1400 5250 -1370
rect 5130 -1440 5250 -1400
rect 5130 -1470 5175 -1440
rect 5205 -1470 5250 -1440
rect 5130 -1510 5250 -1470
rect 5130 -1540 5175 -1510
rect 5205 -1540 5250 -1510
rect 5130 -1580 5250 -1540
rect 5130 -1610 5175 -1580
rect 5205 -1610 5250 -1580
rect 5130 -1645 5250 -1610
rect 5130 -1675 5175 -1645
rect 5205 -1675 5250 -1645
rect 5130 -1705 5250 -1675
rect 5130 -1735 5175 -1705
rect 5205 -1735 5250 -1705
rect 5130 -1770 5250 -1735
rect 5130 -1800 5175 -1770
rect 5205 -1800 5250 -1770
rect 5130 -1840 5250 -1800
rect 5130 -1870 5175 -1840
rect 5205 -1870 5250 -1840
rect 5130 -1910 5250 -1870
rect 5130 -1940 5175 -1910
rect 5205 -1940 5250 -1910
rect 5130 -1980 5250 -1940
rect 5130 -2010 5175 -1980
rect 5205 -2010 5250 -1980
rect 5130 -2045 5250 -2010
rect 5130 -2075 5175 -2045
rect 5205 -2075 5250 -2045
rect 5130 -2105 5250 -2075
rect 5130 -2135 5175 -2105
rect 5205 -2135 5250 -2105
rect 5130 -2170 5250 -2135
rect 5130 -2200 5175 -2170
rect 5205 -2200 5250 -2170
rect 5130 -2240 5250 -2200
rect 5130 -2270 5175 -2240
rect 5205 -2270 5250 -2240
rect 5130 -2310 5250 -2270
rect 5130 -2340 5175 -2310
rect 5205 -2340 5250 -2310
rect 5130 -2380 5250 -2340
rect 5130 -2410 5175 -2380
rect 5205 -2410 5250 -2380
rect 5130 -2445 5250 -2410
rect 5130 -2475 5175 -2445
rect 5205 -2475 5250 -2445
rect 5130 -2505 5250 -2475
rect 5130 -2535 5175 -2505
rect 5205 -2535 5250 -2505
rect 5130 -2570 5250 -2535
rect 5130 -2600 5175 -2570
rect 5205 -2600 5250 -2570
rect 5130 -2640 5250 -2600
rect 5130 -2670 5175 -2640
rect 5205 -2670 5250 -2640
rect 5130 -2710 5250 -2670
rect 5130 -2740 5175 -2710
rect 5205 -2740 5250 -2710
rect 5130 -2780 5250 -2740
rect 5130 -2810 5175 -2780
rect 5205 -2810 5250 -2780
rect 5130 -2845 5250 -2810
rect 5130 -2875 5175 -2845
rect 5205 -2875 5250 -2845
rect 5130 -2905 5250 -2875
rect 5130 -2935 5175 -2905
rect 5205 -2935 5250 -2905
rect 5130 -2970 5250 -2935
rect 5130 -3000 5175 -2970
rect 5205 -3000 5250 -2970
rect 5130 -3040 5250 -3000
rect 5130 -3070 5175 -3040
rect 5205 -3070 5250 -3040
rect 5130 -3110 5250 -3070
rect 5130 -3140 5175 -3110
rect 5205 -3140 5250 -3110
rect 5130 -3180 5250 -3140
rect 5130 -3210 5175 -3180
rect 5205 -3210 5250 -3180
rect 5130 -3245 5250 -3210
rect 5130 -3275 5175 -3245
rect 5205 -3275 5250 -3245
rect 5130 -3305 5250 -3275
rect 5130 -3335 5175 -3305
rect 5205 -3335 5250 -3305
rect 5130 -3370 5250 -3335
rect 5130 -3400 5175 -3370
rect 5205 -3400 5250 -3370
rect 5130 -3440 5250 -3400
rect 5130 -3470 5175 -3440
rect 5205 -3470 5250 -3440
rect 5130 -3510 5250 -3470
rect 5130 -3540 5175 -3510
rect 5205 -3540 5250 -3510
rect 5130 -3580 5250 -3540
rect 5130 -3610 5175 -3580
rect 5205 -3610 5250 -3580
rect 5130 -3645 5250 -3610
rect 5130 -3675 5175 -3645
rect 5205 -3675 5250 -3645
rect 5130 -3705 5250 -3675
rect 5130 -3735 5175 -3705
rect 5205 -3735 5250 -3705
rect 5130 -3770 5250 -3735
rect 5130 -3800 5175 -3770
rect 5205 -3800 5250 -3770
rect 5130 -3840 5250 -3800
rect 5130 -3870 5175 -3840
rect 5205 -3870 5250 -3840
rect 5130 -3910 5250 -3870
rect 5130 -3940 5175 -3910
rect 5205 -3940 5250 -3910
rect 5130 -3980 5250 -3940
rect 5130 -4010 5175 -3980
rect 5205 -4010 5250 -3980
rect 5130 -4045 5250 -4010
rect 5130 -4075 5175 -4045
rect 5205 -4075 5250 -4045
rect 5130 -4105 5250 -4075
rect 5130 -4135 5175 -4105
rect 5205 -4135 5250 -4105
rect 5130 -4170 5250 -4135
rect 5130 -4200 5175 -4170
rect 5205 -4200 5250 -4170
rect 5130 -4240 5250 -4200
rect 5130 -4270 5175 -4240
rect 5205 -4270 5250 -4240
rect 5130 -4310 5250 -4270
rect 5130 -4340 5175 -4310
rect 5205 -4340 5250 -4310
rect 5130 -4380 5250 -4340
rect 5130 -4410 5175 -4380
rect 5205 -4410 5250 -4380
rect 5130 -4445 5250 -4410
rect 5130 -4475 5175 -4445
rect 5205 -4475 5250 -4445
rect 5130 -4490 5250 -4475
rect 5480 -1305 5600 -1240
rect 5480 -1335 5525 -1305
rect 5555 -1335 5600 -1305
rect 5480 -1370 5600 -1335
rect 5480 -1400 5525 -1370
rect 5555 -1400 5600 -1370
rect 5480 -1440 5600 -1400
rect 5480 -1470 5525 -1440
rect 5555 -1470 5600 -1440
rect 5480 -1510 5600 -1470
rect 5480 -1540 5525 -1510
rect 5555 -1540 5600 -1510
rect 5480 -1580 5600 -1540
rect 5480 -1610 5525 -1580
rect 5555 -1610 5600 -1580
rect 5480 -1645 5600 -1610
rect 5480 -1675 5525 -1645
rect 5555 -1675 5600 -1645
rect 5480 -1705 5600 -1675
rect 5480 -1735 5525 -1705
rect 5555 -1735 5600 -1705
rect 5480 -1770 5600 -1735
rect 5480 -1800 5525 -1770
rect 5555 -1800 5600 -1770
rect 5480 -1840 5600 -1800
rect 5480 -1870 5525 -1840
rect 5555 -1870 5600 -1840
rect 5480 -1910 5600 -1870
rect 5480 -1940 5525 -1910
rect 5555 -1940 5600 -1910
rect 5480 -1980 5600 -1940
rect 5480 -2010 5525 -1980
rect 5555 -2010 5600 -1980
rect 5480 -2045 5600 -2010
rect 5480 -2075 5525 -2045
rect 5555 -2075 5600 -2045
rect 5480 -2105 5600 -2075
rect 5480 -2135 5525 -2105
rect 5555 -2135 5600 -2105
rect 5480 -2170 5600 -2135
rect 5480 -2200 5525 -2170
rect 5555 -2200 5600 -2170
rect 5480 -2240 5600 -2200
rect 5480 -2270 5525 -2240
rect 5555 -2270 5600 -2240
rect 5480 -2310 5600 -2270
rect 5480 -2340 5525 -2310
rect 5555 -2340 5600 -2310
rect 5480 -2380 5600 -2340
rect 5480 -2410 5525 -2380
rect 5555 -2410 5600 -2380
rect 5480 -2445 5600 -2410
rect 5480 -2475 5525 -2445
rect 5555 -2475 5600 -2445
rect 5480 -2505 5600 -2475
rect 5480 -2535 5525 -2505
rect 5555 -2535 5600 -2505
rect 5480 -2570 5600 -2535
rect 5480 -2600 5525 -2570
rect 5555 -2600 5600 -2570
rect 5480 -2640 5600 -2600
rect 5480 -2670 5525 -2640
rect 5555 -2670 5600 -2640
rect 5480 -2710 5600 -2670
rect 5480 -2740 5525 -2710
rect 5555 -2740 5600 -2710
rect 5480 -2780 5600 -2740
rect 5480 -2810 5525 -2780
rect 5555 -2810 5600 -2780
rect 5480 -2845 5600 -2810
rect 5480 -2875 5525 -2845
rect 5555 -2875 5600 -2845
rect 5480 -2905 5600 -2875
rect 5480 -2935 5525 -2905
rect 5555 -2935 5600 -2905
rect 5480 -2970 5600 -2935
rect 5480 -3000 5525 -2970
rect 5555 -3000 5600 -2970
rect 5480 -3040 5600 -3000
rect 5480 -3070 5525 -3040
rect 5555 -3070 5600 -3040
rect 5480 -3110 5600 -3070
rect 5480 -3140 5525 -3110
rect 5555 -3140 5600 -3110
rect 5480 -3180 5600 -3140
rect 5480 -3210 5525 -3180
rect 5555 -3210 5600 -3180
rect 5480 -3245 5600 -3210
rect 5480 -3275 5525 -3245
rect 5555 -3275 5600 -3245
rect 5480 -3305 5600 -3275
rect 5480 -3335 5525 -3305
rect 5555 -3335 5600 -3305
rect 5480 -3370 5600 -3335
rect 5480 -3400 5525 -3370
rect 5555 -3400 5600 -3370
rect 5480 -3440 5600 -3400
rect 5480 -3470 5525 -3440
rect 5555 -3470 5600 -3440
rect 5480 -3510 5600 -3470
rect 5480 -3540 5525 -3510
rect 5555 -3540 5600 -3510
rect 5480 -3580 5600 -3540
rect 5480 -3610 5525 -3580
rect 5555 -3610 5600 -3580
rect 5480 -3645 5600 -3610
rect 5480 -3675 5525 -3645
rect 5555 -3675 5600 -3645
rect 5480 -3705 5600 -3675
rect 5480 -3735 5525 -3705
rect 5555 -3735 5600 -3705
rect 5480 -3770 5600 -3735
rect 5480 -3800 5525 -3770
rect 5555 -3800 5600 -3770
rect 5480 -3840 5600 -3800
rect 5480 -3870 5525 -3840
rect 5555 -3870 5600 -3840
rect 5480 -3910 5600 -3870
rect 5480 -3940 5525 -3910
rect 5555 -3940 5600 -3910
rect 5480 -3980 5600 -3940
rect 5480 -4010 5525 -3980
rect 5555 -4010 5600 -3980
rect 5480 -4045 5600 -4010
rect 5480 -4075 5525 -4045
rect 5555 -4075 5600 -4045
rect 5480 -4105 5600 -4075
rect 5480 -4135 5525 -4105
rect 5555 -4135 5600 -4105
rect 5480 -4170 5600 -4135
rect 5480 -4200 5525 -4170
rect 5555 -4200 5600 -4170
rect 5480 -4240 5600 -4200
rect 5480 -4270 5525 -4240
rect 5555 -4270 5600 -4240
rect 5480 -4310 5600 -4270
rect 5480 -4340 5525 -4310
rect 5555 -4340 5600 -4310
rect 5480 -4380 5600 -4340
rect 5480 -4410 5525 -4380
rect 5555 -4410 5600 -4380
rect 5480 -4445 5600 -4410
rect 5480 -4475 5525 -4445
rect 5555 -4475 5600 -4445
rect 5480 -4490 5600 -4475
rect 5830 -1305 5950 -1240
rect 5830 -1335 5875 -1305
rect 5905 -1335 5950 -1305
rect 5830 -1370 5950 -1335
rect 5830 -1400 5875 -1370
rect 5905 -1400 5950 -1370
rect 5830 -1440 5950 -1400
rect 5830 -1470 5875 -1440
rect 5905 -1470 5950 -1440
rect 5830 -1510 5950 -1470
rect 5830 -1540 5875 -1510
rect 5905 -1540 5950 -1510
rect 5830 -1580 5950 -1540
rect 5830 -1610 5875 -1580
rect 5905 -1610 5950 -1580
rect 5830 -1645 5950 -1610
rect 5830 -1675 5875 -1645
rect 5905 -1675 5950 -1645
rect 5830 -1705 5950 -1675
rect 5830 -1735 5875 -1705
rect 5905 -1735 5950 -1705
rect 5830 -1770 5950 -1735
rect 5830 -1800 5875 -1770
rect 5905 -1800 5950 -1770
rect 5830 -1840 5950 -1800
rect 5830 -1870 5875 -1840
rect 5905 -1870 5950 -1840
rect 5830 -1910 5950 -1870
rect 5830 -1940 5875 -1910
rect 5905 -1940 5950 -1910
rect 5830 -1980 5950 -1940
rect 5830 -2010 5875 -1980
rect 5905 -2010 5950 -1980
rect 5830 -2045 5950 -2010
rect 5830 -2075 5875 -2045
rect 5905 -2075 5950 -2045
rect 5830 -2105 5950 -2075
rect 5830 -2135 5875 -2105
rect 5905 -2135 5950 -2105
rect 5830 -2170 5950 -2135
rect 5830 -2200 5875 -2170
rect 5905 -2200 5950 -2170
rect 5830 -2240 5950 -2200
rect 5830 -2270 5875 -2240
rect 5905 -2270 5950 -2240
rect 5830 -2310 5950 -2270
rect 5830 -2340 5875 -2310
rect 5905 -2340 5950 -2310
rect 5830 -2380 5950 -2340
rect 5830 -2410 5875 -2380
rect 5905 -2410 5950 -2380
rect 5830 -2445 5950 -2410
rect 5830 -2475 5875 -2445
rect 5905 -2475 5950 -2445
rect 5830 -2505 5950 -2475
rect 5830 -2535 5875 -2505
rect 5905 -2535 5950 -2505
rect 5830 -2570 5950 -2535
rect 5830 -2600 5875 -2570
rect 5905 -2600 5950 -2570
rect 5830 -2640 5950 -2600
rect 5830 -2670 5875 -2640
rect 5905 -2670 5950 -2640
rect 5830 -2710 5950 -2670
rect 5830 -2740 5875 -2710
rect 5905 -2740 5950 -2710
rect 5830 -2780 5950 -2740
rect 5830 -2810 5875 -2780
rect 5905 -2810 5950 -2780
rect 5830 -2845 5950 -2810
rect 5830 -2875 5875 -2845
rect 5905 -2875 5950 -2845
rect 5830 -2905 5950 -2875
rect 5830 -2935 5875 -2905
rect 5905 -2935 5950 -2905
rect 5830 -2970 5950 -2935
rect 5830 -3000 5875 -2970
rect 5905 -3000 5950 -2970
rect 5830 -3040 5950 -3000
rect 5830 -3070 5875 -3040
rect 5905 -3070 5950 -3040
rect 5830 -3110 5950 -3070
rect 5830 -3140 5875 -3110
rect 5905 -3140 5950 -3110
rect 5830 -3180 5950 -3140
rect 5830 -3210 5875 -3180
rect 5905 -3210 5950 -3180
rect 5830 -3245 5950 -3210
rect 5830 -3275 5875 -3245
rect 5905 -3275 5950 -3245
rect 5830 -3305 5950 -3275
rect 5830 -3335 5875 -3305
rect 5905 -3335 5950 -3305
rect 5830 -3370 5950 -3335
rect 5830 -3400 5875 -3370
rect 5905 -3400 5950 -3370
rect 5830 -3440 5950 -3400
rect 5830 -3470 5875 -3440
rect 5905 -3470 5950 -3440
rect 5830 -3510 5950 -3470
rect 5830 -3540 5875 -3510
rect 5905 -3540 5950 -3510
rect 5830 -3580 5950 -3540
rect 5830 -3610 5875 -3580
rect 5905 -3610 5950 -3580
rect 5830 -3645 5950 -3610
rect 5830 -3675 5875 -3645
rect 5905 -3675 5950 -3645
rect 5830 -3705 5950 -3675
rect 5830 -3735 5875 -3705
rect 5905 -3735 5950 -3705
rect 5830 -3770 5950 -3735
rect 5830 -3800 5875 -3770
rect 5905 -3800 5950 -3770
rect 5830 -3840 5950 -3800
rect 5830 -3870 5875 -3840
rect 5905 -3870 5950 -3840
rect 5830 -3910 5950 -3870
rect 5830 -3940 5875 -3910
rect 5905 -3940 5950 -3910
rect 5830 -3980 5950 -3940
rect 5830 -4010 5875 -3980
rect 5905 -4010 5950 -3980
rect 5830 -4045 5950 -4010
rect 5830 -4075 5875 -4045
rect 5905 -4075 5950 -4045
rect 5830 -4105 5950 -4075
rect 5830 -4135 5875 -4105
rect 5905 -4135 5950 -4105
rect 5830 -4170 5950 -4135
rect 5830 -4200 5875 -4170
rect 5905 -4200 5950 -4170
rect 5830 -4240 5950 -4200
rect 5830 -4270 5875 -4240
rect 5905 -4270 5950 -4240
rect 5830 -4310 5950 -4270
rect 5830 -4340 5875 -4310
rect 5905 -4340 5950 -4310
rect 5830 -4380 5950 -4340
rect 5830 -4410 5875 -4380
rect 5905 -4410 5950 -4380
rect 5830 -4445 5950 -4410
rect 5830 -4475 5875 -4445
rect 5905 -4475 5950 -4445
rect 5830 -4490 5950 -4475
rect 6180 -1305 6300 -1240
rect 6180 -1335 6225 -1305
rect 6255 -1335 6300 -1305
rect 6180 -1370 6300 -1335
rect 6180 -1400 6225 -1370
rect 6255 -1400 6300 -1370
rect 6180 -1440 6300 -1400
rect 6180 -1470 6225 -1440
rect 6255 -1470 6300 -1440
rect 6180 -1510 6300 -1470
rect 6180 -1540 6225 -1510
rect 6255 -1540 6300 -1510
rect 6180 -1580 6300 -1540
rect 6180 -1610 6225 -1580
rect 6255 -1610 6300 -1580
rect 6180 -1645 6300 -1610
rect 6180 -1675 6225 -1645
rect 6255 -1675 6300 -1645
rect 6180 -1705 6300 -1675
rect 6180 -1735 6225 -1705
rect 6255 -1735 6300 -1705
rect 6180 -1770 6300 -1735
rect 6180 -1800 6225 -1770
rect 6255 -1800 6300 -1770
rect 6180 -1840 6300 -1800
rect 6180 -1870 6225 -1840
rect 6255 -1870 6300 -1840
rect 6180 -1910 6300 -1870
rect 6180 -1940 6225 -1910
rect 6255 -1940 6300 -1910
rect 6180 -1980 6300 -1940
rect 6180 -2010 6225 -1980
rect 6255 -2010 6300 -1980
rect 6180 -2045 6300 -2010
rect 6180 -2075 6225 -2045
rect 6255 -2075 6300 -2045
rect 6180 -2105 6300 -2075
rect 6180 -2135 6225 -2105
rect 6255 -2135 6300 -2105
rect 6180 -2170 6300 -2135
rect 6180 -2200 6225 -2170
rect 6255 -2200 6300 -2170
rect 6180 -2240 6300 -2200
rect 6180 -2270 6225 -2240
rect 6255 -2270 6300 -2240
rect 6180 -2310 6300 -2270
rect 6180 -2340 6225 -2310
rect 6255 -2340 6300 -2310
rect 6180 -2380 6300 -2340
rect 6180 -2410 6225 -2380
rect 6255 -2410 6300 -2380
rect 6180 -2445 6300 -2410
rect 6180 -2475 6225 -2445
rect 6255 -2475 6300 -2445
rect 6180 -2505 6300 -2475
rect 6180 -2535 6225 -2505
rect 6255 -2535 6300 -2505
rect 6180 -2570 6300 -2535
rect 6180 -2600 6225 -2570
rect 6255 -2600 6300 -2570
rect 6180 -2640 6300 -2600
rect 6180 -2670 6225 -2640
rect 6255 -2670 6300 -2640
rect 6180 -2710 6300 -2670
rect 6180 -2740 6225 -2710
rect 6255 -2740 6300 -2710
rect 6180 -2780 6300 -2740
rect 6180 -2810 6225 -2780
rect 6255 -2810 6300 -2780
rect 6180 -2845 6300 -2810
rect 6180 -2875 6225 -2845
rect 6255 -2875 6300 -2845
rect 6180 -2905 6300 -2875
rect 6180 -2935 6225 -2905
rect 6255 -2935 6300 -2905
rect 6180 -2970 6300 -2935
rect 6180 -3000 6225 -2970
rect 6255 -3000 6300 -2970
rect 6180 -3040 6300 -3000
rect 6180 -3070 6225 -3040
rect 6255 -3070 6300 -3040
rect 6180 -3110 6300 -3070
rect 6180 -3140 6225 -3110
rect 6255 -3140 6300 -3110
rect 6180 -3180 6300 -3140
rect 6180 -3210 6225 -3180
rect 6255 -3210 6300 -3180
rect 6180 -3245 6300 -3210
rect 6180 -3275 6225 -3245
rect 6255 -3275 6300 -3245
rect 6180 -3305 6300 -3275
rect 6180 -3335 6225 -3305
rect 6255 -3335 6300 -3305
rect 6180 -3370 6300 -3335
rect 6180 -3400 6225 -3370
rect 6255 -3400 6300 -3370
rect 6180 -3440 6300 -3400
rect 6180 -3470 6225 -3440
rect 6255 -3470 6300 -3440
rect 6180 -3510 6300 -3470
rect 6180 -3540 6225 -3510
rect 6255 -3540 6300 -3510
rect 6180 -3580 6300 -3540
rect 6180 -3610 6225 -3580
rect 6255 -3610 6300 -3580
rect 6180 -3645 6300 -3610
rect 6180 -3675 6225 -3645
rect 6255 -3675 6300 -3645
rect 6180 -3705 6300 -3675
rect 6180 -3735 6225 -3705
rect 6255 -3735 6300 -3705
rect 6180 -3770 6300 -3735
rect 6180 -3800 6225 -3770
rect 6255 -3800 6300 -3770
rect 6180 -3840 6300 -3800
rect 6180 -3870 6225 -3840
rect 6255 -3870 6300 -3840
rect 6180 -3910 6300 -3870
rect 6180 -3940 6225 -3910
rect 6255 -3940 6300 -3910
rect 6180 -3980 6300 -3940
rect 6180 -4010 6225 -3980
rect 6255 -4010 6300 -3980
rect 6180 -4045 6300 -4010
rect 6180 -4075 6225 -4045
rect 6255 -4075 6300 -4045
rect 6180 -4105 6300 -4075
rect 6180 -4135 6225 -4105
rect 6255 -4135 6300 -4105
rect 6180 -4170 6300 -4135
rect 6180 -4200 6225 -4170
rect 6255 -4200 6300 -4170
rect 6180 -4240 6300 -4200
rect 6180 -4270 6225 -4240
rect 6255 -4270 6300 -4240
rect 6180 -4310 6300 -4270
rect 6180 -4340 6225 -4310
rect 6255 -4340 6300 -4310
rect 6180 -4380 6300 -4340
rect 6180 -4410 6225 -4380
rect 6255 -4410 6300 -4380
rect 6180 -4445 6300 -4410
rect 6180 -4475 6225 -4445
rect 6255 -4475 6300 -4445
rect 6180 -4490 6300 -4475
rect 6530 -1305 6650 -1240
rect 6530 -1335 6575 -1305
rect 6605 -1335 6650 -1305
rect 6530 -1370 6650 -1335
rect 6530 -1400 6575 -1370
rect 6605 -1400 6650 -1370
rect 6530 -1440 6650 -1400
rect 6530 -1470 6575 -1440
rect 6605 -1470 6650 -1440
rect 6530 -1510 6650 -1470
rect 6530 -1540 6575 -1510
rect 6605 -1540 6650 -1510
rect 6530 -1580 6650 -1540
rect 6530 -1610 6575 -1580
rect 6605 -1610 6650 -1580
rect 6530 -1645 6650 -1610
rect 6530 -1675 6575 -1645
rect 6605 -1675 6650 -1645
rect 6530 -1705 6650 -1675
rect 6530 -1735 6575 -1705
rect 6605 -1735 6650 -1705
rect 6530 -1770 6650 -1735
rect 6530 -1800 6575 -1770
rect 6605 -1800 6650 -1770
rect 6530 -1840 6650 -1800
rect 6530 -1870 6575 -1840
rect 6605 -1870 6650 -1840
rect 6530 -1910 6650 -1870
rect 6530 -1940 6575 -1910
rect 6605 -1940 6650 -1910
rect 6530 -1980 6650 -1940
rect 6530 -2010 6575 -1980
rect 6605 -2010 6650 -1980
rect 6530 -2045 6650 -2010
rect 6530 -2075 6575 -2045
rect 6605 -2075 6650 -2045
rect 6530 -2105 6650 -2075
rect 6530 -2135 6575 -2105
rect 6605 -2135 6650 -2105
rect 6530 -2170 6650 -2135
rect 6530 -2200 6575 -2170
rect 6605 -2200 6650 -2170
rect 6530 -2240 6650 -2200
rect 6530 -2270 6575 -2240
rect 6605 -2270 6650 -2240
rect 6530 -2310 6650 -2270
rect 6530 -2340 6575 -2310
rect 6605 -2340 6650 -2310
rect 6530 -2380 6650 -2340
rect 6530 -2410 6575 -2380
rect 6605 -2410 6650 -2380
rect 6530 -2445 6650 -2410
rect 6530 -2475 6575 -2445
rect 6605 -2475 6650 -2445
rect 6530 -2505 6650 -2475
rect 6530 -2535 6575 -2505
rect 6605 -2535 6650 -2505
rect 6530 -2570 6650 -2535
rect 6530 -2600 6575 -2570
rect 6605 -2600 6650 -2570
rect 6530 -2640 6650 -2600
rect 6530 -2670 6575 -2640
rect 6605 -2670 6650 -2640
rect 6530 -2710 6650 -2670
rect 6530 -2740 6575 -2710
rect 6605 -2740 6650 -2710
rect 6530 -2780 6650 -2740
rect 6530 -2810 6575 -2780
rect 6605 -2810 6650 -2780
rect 6530 -2845 6650 -2810
rect 6530 -2875 6575 -2845
rect 6605 -2875 6650 -2845
rect 6530 -2905 6650 -2875
rect 6530 -2935 6575 -2905
rect 6605 -2935 6650 -2905
rect 6530 -2970 6650 -2935
rect 6530 -3000 6575 -2970
rect 6605 -3000 6650 -2970
rect 6530 -3040 6650 -3000
rect 6530 -3070 6575 -3040
rect 6605 -3070 6650 -3040
rect 6530 -3110 6650 -3070
rect 6530 -3140 6575 -3110
rect 6605 -3140 6650 -3110
rect 6530 -3180 6650 -3140
rect 6530 -3210 6575 -3180
rect 6605 -3210 6650 -3180
rect 6530 -3245 6650 -3210
rect 6530 -3275 6575 -3245
rect 6605 -3275 6650 -3245
rect 6530 -3305 6650 -3275
rect 6530 -3335 6575 -3305
rect 6605 -3335 6650 -3305
rect 6530 -3370 6650 -3335
rect 6530 -3400 6575 -3370
rect 6605 -3400 6650 -3370
rect 6530 -3440 6650 -3400
rect 6530 -3470 6575 -3440
rect 6605 -3470 6650 -3440
rect 6530 -3510 6650 -3470
rect 6530 -3540 6575 -3510
rect 6605 -3540 6650 -3510
rect 6530 -3580 6650 -3540
rect 6530 -3610 6575 -3580
rect 6605 -3610 6650 -3580
rect 6530 -3645 6650 -3610
rect 6530 -3675 6575 -3645
rect 6605 -3675 6650 -3645
rect 6530 -3705 6650 -3675
rect 6530 -3735 6575 -3705
rect 6605 -3735 6650 -3705
rect 6530 -3770 6650 -3735
rect 6530 -3800 6575 -3770
rect 6605 -3800 6650 -3770
rect 6530 -3840 6650 -3800
rect 6530 -3870 6575 -3840
rect 6605 -3870 6650 -3840
rect 6530 -3910 6650 -3870
rect 6530 -3940 6575 -3910
rect 6605 -3940 6650 -3910
rect 6530 -3980 6650 -3940
rect 6530 -4010 6575 -3980
rect 6605 -4010 6650 -3980
rect 6530 -4045 6650 -4010
rect 6530 -4075 6575 -4045
rect 6605 -4075 6650 -4045
rect 6530 -4105 6650 -4075
rect 6530 -4135 6575 -4105
rect 6605 -4135 6650 -4105
rect 6530 -4170 6650 -4135
rect 6530 -4200 6575 -4170
rect 6605 -4200 6650 -4170
rect 6530 -4240 6650 -4200
rect 6530 -4270 6575 -4240
rect 6605 -4270 6650 -4240
rect 6530 -4310 6650 -4270
rect 6530 -4340 6575 -4310
rect 6605 -4340 6650 -4310
rect 6530 -4380 6650 -4340
rect 6530 -4410 6575 -4380
rect 6605 -4410 6650 -4380
rect 6530 -4445 6650 -4410
rect 6530 -4475 6575 -4445
rect 6605 -4475 6650 -4445
rect 6530 -4490 6650 -4475
rect 6880 -1305 7000 -1240
rect 6880 -1335 6925 -1305
rect 6955 -1335 7000 -1305
rect 6880 -1370 7000 -1335
rect 6880 -1400 6925 -1370
rect 6955 -1400 7000 -1370
rect 6880 -1440 7000 -1400
rect 6880 -1470 6925 -1440
rect 6955 -1470 7000 -1440
rect 6880 -1510 7000 -1470
rect 6880 -1540 6925 -1510
rect 6955 -1540 7000 -1510
rect 6880 -1580 7000 -1540
rect 6880 -1610 6925 -1580
rect 6955 -1610 7000 -1580
rect 6880 -1645 7000 -1610
rect 6880 -1675 6925 -1645
rect 6955 -1675 7000 -1645
rect 6880 -1705 7000 -1675
rect 6880 -1735 6925 -1705
rect 6955 -1735 7000 -1705
rect 6880 -1770 7000 -1735
rect 6880 -1800 6925 -1770
rect 6955 -1800 7000 -1770
rect 6880 -1840 7000 -1800
rect 6880 -1870 6925 -1840
rect 6955 -1870 7000 -1840
rect 6880 -1910 7000 -1870
rect 6880 -1940 6925 -1910
rect 6955 -1940 7000 -1910
rect 6880 -1980 7000 -1940
rect 6880 -2010 6925 -1980
rect 6955 -2010 7000 -1980
rect 6880 -2045 7000 -2010
rect 6880 -2075 6925 -2045
rect 6955 -2075 7000 -2045
rect 6880 -2105 7000 -2075
rect 6880 -2135 6925 -2105
rect 6955 -2135 7000 -2105
rect 6880 -2170 7000 -2135
rect 6880 -2200 6925 -2170
rect 6955 -2200 7000 -2170
rect 6880 -2240 7000 -2200
rect 6880 -2270 6925 -2240
rect 6955 -2270 7000 -2240
rect 6880 -2310 7000 -2270
rect 6880 -2340 6925 -2310
rect 6955 -2340 7000 -2310
rect 6880 -2380 7000 -2340
rect 6880 -2410 6925 -2380
rect 6955 -2410 7000 -2380
rect 6880 -2445 7000 -2410
rect 6880 -2475 6925 -2445
rect 6955 -2475 7000 -2445
rect 6880 -2505 7000 -2475
rect 6880 -2535 6925 -2505
rect 6955 -2535 7000 -2505
rect 6880 -2570 7000 -2535
rect 6880 -2600 6925 -2570
rect 6955 -2600 7000 -2570
rect 6880 -2640 7000 -2600
rect 6880 -2670 6925 -2640
rect 6955 -2670 7000 -2640
rect 6880 -2710 7000 -2670
rect 6880 -2740 6925 -2710
rect 6955 -2740 7000 -2710
rect 6880 -2780 7000 -2740
rect 6880 -2810 6925 -2780
rect 6955 -2810 7000 -2780
rect 6880 -2845 7000 -2810
rect 6880 -2875 6925 -2845
rect 6955 -2875 7000 -2845
rect 6880 -2905 7000 -2875
rect 6880 -2935 6925 -2905
rect 6955 -2935 7000 -2905
rect 6880 -2970 7000 -2935
rect 6880 -3000 6925 -2970
rect 6955 -3000 7000 -2970
rect 6880 -3040 7000 -3000
rect 6880 -3070 6925 -3040
rect 6955 -3070 7000 -3040
rect 6880 -3110 7000 -3070
rect 6880 -3140 6925 -3110
rect 6955 -3140 7000 -3110
rect 6880 -3180 7000 -3140
rect 6880 -3210 6925 -3180
rect 6955 -3210 7000 -3180
rect 6880 -3245 7000 -3210
rect 6880 -3275 6925 -3245
rect 6955 -3275 7000 -3245
rect 6880 -3305 7000 -3275
rect 6880 -3335 6925 -3305
rect 6955 -3335 7000 -3305
rect 6880 -3370 7000 -3335
rect 6880 -3400 6925 -3370
rect 6955 -3400 7000 -3370
rect 6880 -3440 7000 -3400
rect 6880 -3470 6925 -3440
rect 6955 -3470 7000 -3440
rect 6880 -3510 7000 -3470
rect 6880 -3540 6925 -3510
rect 6955 -3540 7000 -3510
rect 6880 -3580 7000 -3540
rect 6880 -3610 6925 -3580
rect 6955 -3610 7000 -3580
rect 6880 -3645 7000 -3610
rect 6880 -3675 6925 -3645
rect 6955 -3675 7000 -3645
rect 6880 -3705 7000 -3675
rect 6880 -3735 6925 -3705
rect 6955 -3735 7000 -3705
rect 6880 -3770 7000 -3735
rect 6880 -3800 6925 -3770
rect 6955 -3800 7000 -3770
rect 6880 -3840 7000 -3800
rect 6880 -3870 6925 -3840
rect 6955 -3870 7000 -3840
rect 6880 -3910 7000 -3870
rect 6880 -3940 6925 -3910
rect 6955 -3940 7000 -3910
rect 6880 -3980 7000 -3940
rect 6880 -4010 6925 -3980
rect 6955 -4010 7000 -3980
rect 6880 -4045 7000 -4010
rect 6880 -4075 6925 -4045
rect 6955 -4075 7000 -4045
rect 6880 -4105 7000 -4075
rect 6880 -4135 6925 -4105
rect 6955 -4135 7000 -4105
rect 6880 -4170 7000 -4135
rect 6880 -4200 6925 -4170
rect 6955 -4200 7000 -4170
rect 6880 -4240 7000 -4200
rect 6880 -4270 6925 -4240
rect 6955 -4270 7000 -4240
rect 6880 -4310 7000 -4270
rect 6880 -4340 6925 -4310
rect 6955 -4340 7000 -4310
rect 6880 -4380 7000 -4340
rect 6880 -4410 6925 -4380
rect 6955 -4410 7000 -4380
rect 6880 -4445 7000 -4410
rect 6880 -4475 6925 -4445
rect 6955 -4475 7000 -4445
rect 6880 -4490 7000 -4475
rect 7230 -1305 7350 -1240
rect 7230 -1335 7275 -1305
rect 7305 -1335 7350 -1305
rect 7230 -1370 7350 -1335
rect 7230 -1400 7275 -1370
rect 7305 -1400 7350 -1370
rect 7230 -1440 7350 -1400
rect 7230 -1470 7275 -1440
rect 7305 -1470 7350 -1440
rect 7230 -1510 7350 -1470
rect 7230 -1540 7275 -1510
rect 7305 -1540 7350 -1510
rect 7230 -1580 7350 -1540
rect 7230 -1610 7275 -1580
rect 7305 -1610 7350 -1580
rect 7230 -1645 7350 -1610
rect 7230 -1675 7275 -1645
rect 7305 -1675 7350 -1645
rect 7230 -1705 7350 -1675
rect 7230 -1735 7275 -1705
rect 7305 -1735 7350 -1705
rect 7230 -1770 7350 -1735
rect 7230 -1800 7275 -1770
rect 7305 -1800 7350 -1770
rect 7230 -1840 7350 -1800
rect 7230 -1870 7275 -1840
rect 7305 -1870 7350 -1840
rect 7230 -1910 7350 -1870
rect 7230 -1940 7275 -1910
rect 7305 -1940 7350 -1910
rect 7230 -1980 7350 -1940
rect 7230 -2010 7275 -1980
rect 7305 -2010 7350 -1980
rect 7230 -2045 7350 -2010
rect 7230 -2075 7275 -2045
rect 7305 -2075 7350 -2045
rect 7230 -2105 7350 -2075
rect 7230 -2135 7275 -2105
rect 7305 -2135 7350 -2105
rect 7230 -2170 7350 -2135
rect 7230 -2200 7275 -2170
rect 7305 -2200 7350 -2170
rect 7230 -2240 7350 -2200
rect 7230 -2270 7275 -2240
rect 7305 -2270 7350 -2240
rect 7230 -2310 7350 -2270
rect 7230 -2340 7275 -2310
rect 7305 -2340 7350 -2310
rect 7230 -2380 7350 -2340
rect 7230 -2410 7275 -2380
rect 7305 -2410 7350 -2380
rect 7230 -2445 7350 -2410
rect 7230 -2475 7275 -2445
rect 7305 -2475 7350 -2445
rect 7230 -2505 7350 -2475
rect 7230 -2535 7275 -2505
rect 7305 -2535 7350 -2505
rect 7230 -2570 7350 -2535
rect 7230 -2600 7275 -2570
rect 7305 -2600 7350 -2570
rect 7230 -2640 7350 -2600
rect 7230 -2670 7275 -2640
rect 7305 -2670 7350 -2640
rect 7230 -2710 7350 -2670
rect 7230 -2740 7275 -2710
rect 7305 -2740 7350 -2710
rect 7230 -2780 7350 -2740
rect 7230 -2810 7275 -2780
rect 7305 -2810 7350 -2780
rect 7230 -2845 7350 -2810
rect 7230 -2875 7275 -2845
rect 7305 -2875 7350 -2845
rect 7230 -2905 7350 -2875
rect 7230 -2935 7275 -2905
rect 7305 -2935 7350 -2905
rect 7230 -2970 7350 -2935
rect 7230 -3000 7275 -2970
rect 7305 -3000 7350 -2970
rect 7230 -3040 7350 -3000
rect 7230 -3070 7275 -3040
rect 7305 -3070 7350 -3040
rect 7230 -3110 7350 -3070
rect 7230 -3140 7275 -3110
rect 7305 -3140 7350 -3110
rect 7230 -3180 7350 -3140
rect 7230 -3210 7275 -3180
rect 7305 -3210 7350 -3180
rect 7230 -3245 7350 -3210
rect 7230 -3275 7275 -3245
rect 7305 -3275 7350 -3245
rect 7230 -3305 7350 -3275
rect 7230 -3335 7275 -3305
rect 7305 -3335 7350 -3305
rect 7230 -3370 7350 -3335
rect 7230 -3400 7275 -3370
rect 7305 -3400 7350 -3370
rect 7230 -3440 7350 -3400
rect 7230 -3470 7275 -3440
rect 7305 -3470 7350 -3440
rect 7230 -3510 7350 -3470
rect 7230 -3540 7275 -3510
rect 7305 -3540 7350 -3510
rect 7230 -3580 7350 -3540
rect 7230 -3610 7275 -3580
rect 7305 -3610 7350 -3580
rect 7230 -3645 7350 -3610
rect 7230 -3675 7275 -3645
rect 7305 -3675 7350 -3645
rect 7230 -3705 7350 -3675
rect 7230 -3735 7275 -3705
rect 7305 -3735 7350 -3705
rect 7230 -3770 7350 -3735
rect 7230 -3800 7275 -3770
rect 7305 -3800 7350 -3770
rect 7230 -3840 7350 -3800
rect 7230 -3870 7275 -3840
rect 7305 -3870 7350 -3840
rect 7230 -3910 7350 -3870
rect 7230 -3940 7275 -3910
rect 7305 -3940 7350 -3910
rect 7230 -3980 7350 -3940
rect 7230 -4010 7275 -3980
rect 7305 -4010 7350 -3980
rect 7230 -4045 7350 -4010
rect 7230 -4075 7275 -4045
rect 7305 -4075 7350 -4045
rect 7230 -4105 7350 -4075
rect 7230 -4135 7275 -4105
rect 7305 -4135 7350 -4105
rect 7230 -4170 7350 -4135
rect 7230 -4200 7275 -4170
rect 7305 -4200 7350 -4170
rect 7230 -4240 7350 -4200
rect 7230 -4270 7275 -4240
rect 7305 -4270 7350 -4240
rect 7230 -4310 7350 -4270
rect 7230 -4340 7275 -4310
rect 7305 -4340 7350 -4310
rect 7230 -4380 7350 -4340
rect 7230 -4410 7275 -4380
rect 7305 -4410 7350 -4380
rect 7230 -4445 7350 -4410
rect 7230 -4475 7275 -4445
rect 7305 -4475 7350 -4445
rect 7230 -4490 7350 -4475
rect 7580 -1305 7700 -1240
rect 7580 -1335 7625 -1305
rect 7655 -1335 7700 -1305
rect 7580 -1370 7700 -1335
rect 7580 -1400 7625 -1370
rect 7655 -1400 7700 -1370
rect 7580 -1440 7700 -1400
rect 7580 -1470 7625 -1440
rect 7655 -1470 7700 -1440
rect 7580 -1510 7700 -1470
rect 7580 -1540 7625 -1510
rect 7655 -1540 7700 -1510
rect 7580 -1580 7700 -1540
rect 7580 -1610 7625 -1580
rect 7655 -1610 7700 -1580
rect 7580 -1645 7700 -1610
rect 7580 -1675 7625 -1645
rect 7655 -1675 7700 -1645
rect 7580 -1705 7700 -1675
rect 7580 -1735 7625 -1705
rect 7655 -1735 7700 -1705
rect 7580 -1770 7700 -1735
rect 7580 -1800 7625 -1770
rect 7655 -1800 7700 -1770
rect 7580 -1840 7700 -1800
rect 7580 -1870 7625 -1840
rect 7655 -1870 7700 -1840
rect 7580 -1910 7700 -1870
rect 7580 -1940 7625 -1910
rect 7655 -1940 7700 -1910
rect 7580 -1980 7700 -1940
rect 7580 -2010 7625 -1980
rect 7655 -2010 7700 -1980
rect 7580 -2045 7700 -2010
rect 7580 -2075 7625 -2045
rect 7655 -2075 7700 -2045
rect 7580 -2105 7700 -2075
rect 7580 -2135 7625 -2105
rect 7655 -2135 7700 -2105
rect 7580 -2170 7700 -2135
rect 7580 -2200 7625 -2170
rect 7655 -2200 7700 -2170
rect 7580 -2240 7700 -2200
rect 7580 -2270 7625 -2240
rect 7655 -2270 7700 -2240
rect 7580 -2310 7700 -2270
rect 7580 -2340 7625 -2310
rect 7655 -2340 7700 -2310
rect 7580 -2380 7700 -2340
rect 7580 -2410 7625 -2380
rect 7655 -2410 7700 -2380
rect 7580 -2445 7700 -2410
rect 7580 -2475 7625 -2445
rect 7655 -2475 7700 -2445
rect 7580 -2505 7700 -2475
rect 7580 -2535 7625 -2505
rect 7655 -2535 7700 -2505
rect 7580 -2570 7700 -2535
rect 7580 -2600 7625 -2570
rect 7655 -2600 7700 -2570
rect 7580 -2640 7700 -2600
rect 7580 -2670 7625 -2640
rect 7655 -2670 7700 -2640
rect 7580 -2710 7700 -2670
rect 7580 -2740 7625 -2710
rect 7655 -2740 7700 -2710
rect 7580 -2780 7700 -2740
rect 7580 -2810 7625 -2780
rect 7655 -2810 7700 -2780
rect 7580 -2845 7700 -2810
rect 7580 -2875 7625 -2845
rect 7655 -2875 7700 -2845
rect 7580 -2905 7700 -2875
rect 7580 -2935 7625 -2905
rect 7655 -2935 7700 -2905
rect 7580 -2970 7700 -2935
rect 7580 -3000 7625 -2970
rect 7655 -3000 7700 -2970
rect 7580 -3040 7700 -3000
rect 7580 -3070 7625 -3040
rect 7655 -3070 7700 -3040
rect 7580 -3110 7700 -3070
rect 7580 -3140 7625 -3110
rect 7655 -3140 7700 -3110
rect 7580 -3180 7700 -3140
rect 7580 -3210 7625 -3180
rect 7655 -3210 7700 -3180
rect 7580 -3245 7700 -3210
rect 7580 -3275 7625 -3245
rect 7655 -3275 7700 -3245
rect 7580 -3305 7700 -3275
rect 7580 -3335 7625 -3305
rect 7655 -3335 7700 -3305
rect 7580 -3370 7700 -3335
rect 7580 -3400 7625 -3370
rect 7655 -3400 7700 -3370
rect 7580 -3440 7700 -3400
rect 7580 -3470 7625 -3440
rect 7655 -3470 7700 -3440
rect 7580 -3510 7700 -3470
rect 7580 -3540 7625 -3510
rect 7655 -3540 7700 -3510
rect 7580 -3580 7700 -3540
rect 7580 -3610 7625 -3580
rect 7655 -3610 7700 -3580
rect 7580 -3645 7700 -3610
rect 7580 -3675 7625 -3645
rect 7655 -3675 7700 -3645
rect 7580 -3705 7700 -3675
rect 7580 -3735 7625 -3705
rect 7655 -3735 7700 -3705
rect 7580 -3770 7700 -3735
rect 7580 -3800 7625 -3770
rect 7655 -3800 7700 -3770
rect 7580 -3840 7700 -3800
rect 7580 -3870 7625 -3840
rect 7655 -3870 7700 -3840
rect 7580 -3910 7700 -3870
rect 7580 -3940 7625 -3910
rect 7655 -3940 7700 -3910
rect 7580 -3980 7700 -3940
rect 7580 -4010 7625 -3980
rect 7655 -4010 7700 -3980
rect 7580 -4045 7700 -4010
rect 7580 -4075 7625 -4045
rect 7655 -4075 7700 -4045
rect 7580 -4105 7700 -4075
rect 7580 -4135 7625 -4105
rect 7655 -4135 7700 -4105
rect 7580 -4170 7700 -4135
rect 7580 -4200 7625 -4170
rect 7655 -4200 7700 -4170
rect 7580 -4240 7700 -4200
rect 7580 -4270 7625 -4240
rect 7655 -4270 7700 -4240
rect 7580 -4310 7700 -4270
rect 7580 -4340 7625 -4310
rect 7655 -4340 7700 -4310
rect 7580 -4380 7700 -4340
rect 7580 -4410 7625 -4380
rect 7655 -4410 7700 -4380
rect 7580 -4445 7700 -4410
rect 7580 -4475 7625 -4445
rect 7655 -4475 7700 -4445
rect 7580 -4490 7700 -4475
rect 7930 -1305 8050 -1240
rect 7930 -1335 7975 -1305
rect 8005 -1335 8050 -1305
rect 7930 -1370 8050 -1335
rect 7930 -1400 7975 -1370
rect 8005 -1400 8050 -1370
rect 7930 -1440 8050 -1400
rect 7930 -1470 7975 -1440
rect 8005 -1470 8050 -1440
rect 7930 -1510 8050 -1470
rect 7930 -1540 7975 -1510
rect 8005 -1540 8050 -1510
rect 7930 -1580 8050 -1540
rect 7930 -1610 7975 -1580
rect 8005 -1610 8050 -1580
rect 7930 -1645 8050 -1610
rect 7930 -1675 7975 -1645
rect 8005 -1675 8050 -1645
rect 7930 -1705 8050 -1675
rect 7930 -1735 7975 -1705
rect 8005 -1735 8050 -1705
rect 7930 -1770 8050 -1735
rect 7930 -1800 7975 -1770
rect 8005 -1800 8050 -1770
rect 7930 -1840 8050 -1800
rect 7930 -1870 7975 -1840
rect 8005 -1870 8050 -1840
rect 7930 -1910 8050 -1870
rect 7930 -1940 7975 -1910
rect 8005 -1940 8050 -1910
rect 7930 -1980 8050 -1940
rect 7930 -2010 7975 -1980
rect 8005 -2010 8050 -1980
rect 7930 -2045 8050 -2010
rect 7930 -2075 7975 -2045
rect 8005 -2075 8050 -2045
rect 7930 -2105 8050 -2075
rect 7930 -2135 7975 -2105
rect 8005 -2135 8050 -2105
rect 7930 -2170 8050 -2135
rect 7930 -2200 7975 -2170
rect 8005 -2200 8050 -2170
rect 7930 -2240 8050 -2200
rect 7930 -2270 7975 -2240
rect 8005 -2270 8050 -2240
rect 7930 -2310 8050 -2270
rect 7930 -2340 7975 -2310
rect 8005 -2340 8050 -2310
rect 7930 -2380 8050 -2340
rect 7930 -2410 7975 -2380
rect 8005 -2410 8050 -2380
rect 7930 -2445 8050 -2410
rect 7930 -2475 7975 -2445
rect 8005 -2475 8050 -2445
rect 7930 -2505 8050 -2475
rect 7930 -2535 7975 -2505
rect 8005 -2535 8050 -2505
rect 7930 -2570 8050 -2535
rect 7930 -2600 7975 -2570
rect 8005 -2600 8050 -2570
rect 7930 -2640 8050 -2600
rect 7930 -2670 7975 -2640
rect 8005 -2670 8050 -2640
rect 7930 -2710 8050 -2670
rect 7930 -2740 7975 -2710
rect 8005 -2740 8050 -2710
rect 7930 -2780 8050 -2740
rect 7930 -2810 7975 -2780
rect 8005 -2810 8050 -2780
rect 7930 -2845 8050 -2810
rect 7930 -2875 7975 -2845
rect 8005 -2875 8050 -2845
rect 7930 -2905 8050 -2875
rect 7930 -2935 7975 -2905
rect 8005 -2935 8050 -2905
rect 7930 -2970 8050 -2935
rect 7930 -3000 7975 -2970
rect 8005 -3000 8050 -2970
rect 7930 -3040 8050 -3000
rect 7930 -3070 7975 -3040
rect 8005 -3070 8050 -3040
rect 7930 -3110 8050 -3070
rect 7930 -3140 7975 -3110
rect 8005 -3140 8050 -3110
rect 7930 -3180 8050 -3140
rect 7930 -3210 7975 -3180
rect 8005 -3210 8050 -3180
rect 7930 -3245 8050 -3210
rect 7930 -3275 7975 -3245
rect 8005 -3275 8050 -3245
rect 7930 -3305 8050 -3275
rect 7930 -3335 7975 -3305
rect 8005 -3335 8050 -3305
rect 7930 -3370 8050 -3335
rect 7930 -3400 7975 -3370
rect 8005 -3400 8050 -3370
rect 7930 -3440 8050 -3400
rect 7930 -3470 7975 -3440
rect 8005 -3470 8050 -3440
rect 7930 -3510 8050 -3470
rect 7930 -3540 7975 -3510
rect 8005 -3540 8050 -3510
rect 7930 -3580 8050 -3540
rect 7930 -3610 7975 -3580
rect 8005 -3610 8050 -3580
rect 7930 -3645 8050 -3610
rect 7930 -3675 7975 -3645
rect 8005 -3675 8050 -3645
rect 7930 -3705 8050 -3675
rect 7930 -3735 7975 -3705
rect 8005 -3735 8050 -3705
rect 7930 -3770 8050 -3735
rect 7930 -3800 7975 -3770
rect 8005 -3800 8050 -3770
rect 7930 -3840 8050 -3800
rect 7930 -3870 7975 -3840
rect 8005 -3870 8050 -3840
rect 7930 -3910 8050 -3870
rect 7930 -3940 7975 -3910
rect 8005 -3940 8050 -3910
rect 7930 -3980 8050 -3940
rect 7930 -4010 7975 -3980
rect 8005 -4010 8050 -3980
rect 7930 -4045 8050 -4010
rect 7930 -4075 7975 -4045
rect 8005 -4075 8050 -4045
rect 7930 -4105 8050 -4075
rect 7930 -4135 7975 -4105
rect 8005 -4135 8050 -4105
rect 7930 -4170 8050 -4135
rect 7930 -4200 7975 -4170
rect 8005 -4200 8050 -4170
rect 7930 -4240 8050 -4200
rect 7930 -4270 7975 -4240
rect 8005 -4270 8050 -4240
rect 7930 -4310 8050 -4270
rect 7930 -4340 7975 -4310
rect 8005 -4340 8050 -4310
rect 7930 -4380 8050 -4340
rect 7930 -4410 7975 -4380
rect 8005 -4410 8050 -4380
rect 7930 -4445 8050 -4410
rect 7930 -4475 7975 -4445
rect 8005 -4475 8050 -4445
rect 7930 -4490 8050 -4475
rect 8280 -1305 8400 -1240
rect 8280 -1335 8325 -1305
rect 8355 -1335 8400 -1305
rect 8280 -1370 8400 -1335
rect 8280 -1400 8325 -1370
rect 8355 -1400 8400 -1370
rect 8280 -1440 8400 -1400
rect 8280 -1470 8325 -1440
rect 8355 -1470 8400 -1440
rect 8280 -1510 8400 -1470
rect 8280 -1540 8325 -1510
rect 8355 -1540 8400 -1510
rect 8280 -1580 8400 -1540
rect 8280 -1610 8325 -1580
rect 8355 -1610 8400 -1580
rect 8280 -1645 8400 -1610
rect 8280 -1675 8325 -1645
rect 8355 -1675 8400 -1645
rect 8280 -1705 8400 -1675
rect 8280 -1735 8325 -1705
rect 8355 -1735 8400 -1705
rect 8280 -1770 8400 -1735
rect 8280 -1800 8325 -1770
rect 8355 -1800 8400 -1770
rect 8280 -1840 8400 -1800
rect 8280 -1870 8325 -1840
rect 8355 -1870 8400 -1840
rect 8280 -1910 8400 -1870
rect 8280 -1940 8325 -1910
rect 8355 -1940 8400 -1910
rect 8280 -1980 8400 -1940
rect 8280 -2010 8325 -1980
rect 8355 -2010 8400 -1980
rect 8280 -2045 8400 -2010
rect 8280 -2075 8325 -2045
rect 8355 -2075 8400 -2045
rect 8280 -2105 8400 -2075
rect 8280 -2135 8325 -2105
rect 8355 -2135 8400 -2105
rect 8280 -2170 8400 -2135
rect 8280 -2200 8325 -2170
rect 8355 -2200 8400 -2170
rect 8280 -2240 8400 -2200
rect 8280 -2270 8325 -2240
rect 8355 -2270 8400 -2240
rect 8280 -2310 8400 -2270
rect 8280 -2340 8325 -2310
rect 8355 -2340 8400 -2310
rect 8280 -2380 8400 -2340
rect 8280 -2410 8325 -2380
rect 8355 -2410 8400 -2380
rect 8280 -2445 8400 -2410
rect 8280 -2475 8325 -2445
rect 8355 -2475 8400 -2445
rect 8280 -2505 8400 -2475
rect 8280 -2535 8325 -2505
rect 8355 -2535 8400 -2505
rect 8280 -2570 8400 -2535
rect 8280 -2600 8325 -2570
rect 8355 -2600 8400 -2570
rect 8280 -2640 8400 -2600
rect 8280 -2670 8325 -2640
rect 8355 -2670 8400 -2640
rect 8280 -2710 8400 -2670
rect 8280 -2740 8325 -2710
rect 8355 -2740 8400 -2710
rect 8280 -2780 8400 -2740
rect 8280 -2810 8325 -2780
rect 8355 -2810 8400 -2780
rect 8280 -2845 8400 -2810
rect 8280 -2875 8325 -2845
rect 8355 -2875 8400 -2845
rect 8280 -2905 8400 -2875
rect 8280 -2935 8325 -2905
rect 8355 -2935 8400 -2905
rect 8280 -2970 8400 -2935
rect 8280 -3000 8325 -2970
rect 8355 -3000 8400 -2970
rect 8280 -3040 8400 -3000
rect 8280 -3070 8325 -3040
rect 8355 -3070 8400 -3040
rect 8280 -3110 8400 -3070
rect 8280 -3140 8325 -3110
rect 8355 -3140 8400 -3110
rect 8280 -3180 8400 -3140
rect 8280 -3210 8325 -3180
rect 8355 -3210 8400 -3180
rect 8280 -3245 8400 -3210
rect 8280 -3275 8325 -3245
rect 8355 -3275 8400 -3245
rect 8280 -3305 8400 -3275
rect 8280 -3335 8325 -3305
rect 8355 -3335 8400 -3305
rect 8280 -3370 8400 -3335
rect 8280 -3400 8325 -3370
rect 8355 -3400 8400 -3370
rect 8280 -3440 8400 -3400
rect 8280 -3470 8325 -3440
rect 8355 -3470 8400 -3440
rect 8280 -3510 8400 -3470
rect 8280 -3540 8325 -3510
rect 8355 -3540 8400 -3510
rect 8280 -3580 8400 -3540
rect 8280 -3610 8325 -3580
rect 8355 -3610 8400 -3580
rect 8280 -3645 8400 -3610
rect 8280 -3675 8325 -3645
rect 8355 -3675 8400 -3645
rect 8280 -3705 8400 -3675
rect 8280 -3735 8325 -3705
rect 8355 -3735 8400 -3705
rect 8280 -3770 8400 -3735
rect 8280 -3800 8325 -3770
rect 8355 -3800 8400 -3770
rect 8280 -3840 8400 -3800
rect 8280 -3870 8325 -3840
rect 8355 -3870 8400 -3840
rect 8280 -3910 8400 -3870
rect 8280 -3940 8325 -3910
rect 8355 -3940 8400 -3910
rect 8280 -3980 8400 -3940
rect 8280 -4010 8325 -3980
rect 8355 -4010 8400 -3980
rect 8280 -4045 8400 -4010
rect 8280 -4075 8325 -4045
rect 8355 -4075 8400 -4045
rect 8280 -4105 8400 -4075
rect 8280 -4135 8325 -4105
rect 8355 -4135 8400 -4105
rect 8280 -4170 8400 -4135
rect 8280 -4200 8325 -4170
rect 8355 -4200 8400 -4170
rect 8280 -4240 8400 -4200
rect 8280 -4270 8325 -4240
rect 8355 -4270 8400 -4240
rect 8280 -4310 8400 -4270
rect 8280 -4340 8325 -4310
rect 8355 -4340 8400 -4310
rect 8280 -4380 8400 -4340
rect 8280 -4410 8325 -4380
rect 8355 -4410 8400 -4380
rect 8280 -4445 8400 -4410
rect 8280 -4475 8325 -4445
rect 8355 -4475 8400 -4445
rect 8280 -4490 8400 -4475
rect 8630 -1305 8750 -1240
rect 8630 -1335 8675 -1305
rect 8705 -1335 8750 -1305
rect 8630 -1370 8750 -1335
rect 8630 -1400 8675 -1370
rect 8705 -1400 8750 -1370
rect 8630 -1440 8750 -1400
rect 8630 -1470 8675 -1440
rect 8705 -1470 8750 -1440
rect 8630 -1510 8750 -1470
rect 8630 -1540 8675 -1510
rect 8705 -1540 8750 -1510
rect 8630 -1580 8750 -1540
rect 8630 -1610 8675 -1580
rect 8705 -1610 8750 -1580
rect 8630 -1645 8750 -1610
rect 8630 -1675 8675 -1645
rect 8705 -1675 8750 -1645
rect 8630 -1705 8750 -1675
rect 8630 -1735 8675 -1705
rect 8705 -1735 8750 -1705
rect 8630 -1770 8750 -1735
rect 8630 -1800 8675 -1770
rect 8705 -1800 8750 -1770
rect 8630 -1840 8750 -1800
rect 8630 -1870 8675 -1840
rect 8705 -1870 8750 -1840
rect 8630 -1910 8750 -1870
rect 8630 -1940 8675 -1910
rect 8705 -1940 8750 -1910
rect 8630 -1980 8750 -1940
rect 8630 -2010 8675 -1980
rect 8705 -2010 8750 -1980
rect 8630 -2045 8750 -2010
rect 8630 -2075 8675 -2045
rect 8705 -2075 8750 -2045
rect 8630 -2105 8750 -2075
rect 8630 -2135 8675 -2105
rect 8705 -2135 8750 -2105
rect 8630 -2170 8750 -2135
rect 8630 -2200 8675 -2170
rect 8705 -2200 8750 -2170
rect 8630 -2240 8750 -2200
rect 8630 -2270 8675 -2240
rect 8705 -2270 8750 -2240
rect 8630 -2310 8750 -2270
rect 8630 -2340 8675 -2310
rect 8705 -2340 8750 -2310
rect 8630 -2380 8750 -2340
rect 8630 -2410 8675 -2380
rect 8705 -2410 8750 -2380
rect 8630 -2445 8750 -2410
rect 8630 -2475 8675 -2445
rect 8705 -2475 8750 -2445
rect 8630 -2505 8750 -2475
rect 8630 -2535 8675 -2505
rect 8705 -2535 8750 -2505
rect 8630 -2570 8750 -2535
rect 8630 -2600 8675 -2570
rect 8705 -2600 8750 -2570
rect 8630 -2640 8750 -2600
rect 8630 -2670 8675 -2640
rect 8705 -2670 8750 -2640
rect 8630 -2710 8750 -2670
rect 8630 -2740 8675 -2710
rect 8705 -2740 8750 -2710
rect 8630 -2780 8750 -2740
rect 8630 -2810 8675 -2780
rect 8705 -2810 8750 -2780
rect 8630 -2845 8750 -2810
rect 8630 -2875 8675 -2845
rect 8705 -2875 8750 -2845
rect 8630 -2905 8750 -2875
rect 8630 -2935 8675 -2905
rect 8705 -2935 8750 -2905
rect 8630 -2970 8750 -2935
rect 8630 -3000 8675 -2970
rect 8705 -3000 8750 -2970
rect 8630 -3040 8750 -3000
rect 8630 -3070 8675 -3040
rect 8705 -3070 8750 -3040
rect 8630 -3110 8750 -3070
rect 8630 -3140 8675 -3110
rect 8705 -3140 8750 -3110
rect 8630 -3180 8750 -3140
rect 8630 -3210 8675 -3180
rect 8705 -3210 8750 -3180
rect 8630 -3245 8750 -3210
rect 8630 -3275 8675 -3245
rect 8705 -3275 8750 -3245
rect 8630 -3305 8750 -3275
rect 8630 -3335 8675 -3305
rect 8705 -3335 8750 -3305
rect 8630 -3370 8750 -3335
rect 8630 -3400 8675 -3370
rect 8705 -3400 8750 -3370
rect 8630 -3440 8750 -3400
rect 8630 -3470 8675 -3440
rect 8705 -3470 8750 -3440
rect 8630 -3510 8750 -3470
rect 8630 -3540 8675 -3510
rect 8705 -3540 8750 -3510
rect 8630 -3580 8750 -3540
rect 8630 -3610 8675 -3580
rect 8705 -3610 8750 -3580
rect 8630 -3645 8750 -3610
rect 8630 -3675 8675 -3645
rect 8705 -3675 8750 -3645
rect 8630 -3705 8750 -3675
rect 8630 -3735 8675 -3705
rect 8705 -3735 8750 -3705
rect 8630 -3770 8750 -3735
rect 8630 -3800 8675 -3770
rect 8705 -3800 8750 -3770
rect 8630 -3840 8750 -3800
rect 8630 -3870 8675 -3840
rect 8705 -3870 8750 -3840
rect 8630 -3910 8750 -3870
rect 8630 -3940 8675 -3910
rect 8705 -3940 8750 -3910
rect 8630 -3980 8750 -3940
rect 8630 -4010 8675 -3980
rect 8705 -4010 8750 -3980
rect 8630 -4045 8750 -4010
rect 8630 -4075 8675 -4045
rect 8705 -4075 8750 -4045
rect 8630 -4105 8750 -4075
rect 8630 -4135 8675 -4105
rect 8705 -4135 8750 -4105
rect 8630 -4170 8750 -4135
rect 8630 -4200 8675 -4170
rect 8705 -4200 8750 -4170
rect 8630 -4240 8750 -4200
rect 8630 -4270 8675 -4240
rect 8705 -4270 8750 -4240
rect 8630 -4310 8750 -4270
rect 8630 -4340 8675 -4310
rect 8705 -4340 8750 -4310
rect 8630 -4380 8750 -4340
rect 8630 -4410 8675 -4380
rect 8705 -4410 8750 -4380
rect 8630 -4445 8750 -4410
rect 8630 -4475 8675 -4445
rect 8705 -4475 8750 -4445
rect 8630 -4490 8750 -4475
<< via1 >>
rect 2335 20880 2365 20910
rect 2335 20815 2365 20845
rect 2335 20745 2365 20775
rect 2335 20675 2365 20705
rect 2335 20605 2365 20635
rect 2335 20540 2365 20570
rect 2335 20480 2365 20510
rect 2335 20415 2365 20445
rect 2335 20345 2365 20375
rect 2335 20275 2365 20305
rect 2335 20205 2365 20235
rect 2335 20140 2365 20170
rect 2335 20080 2365 20110
rect 2335 20015 2365 20045
rect 2335 19945 2365 19975
rect 2335 19875 2365 19905
rect 2335 19805 2365 19835
rect 2335 19740 2365 19770
rect 2335 19680 2365 19710
rect 2335 19615 2365 19645
rect 2335 19545 2365 19575
rect 2335 19475 2365 19505
rect 2335 19405 2365 19435
rect 2335 19340 2365 19370
rect 2335 19280 2365 19310
rect 2335 19215 2365 19245
rect 2335 19145 2365 19175
rect 2335 19075 2365 19105
rect 2335 19005 2365 19035
rect 2335 18940 2365 18970
rect 2335 18880 2365 18910
rect 2335 18815 2365 18845
rect 2335 18745 2365 18775
rect 2335 18675 2365 18705
rect 2335 18605 2365 18635
rect 2335 18540 2365 18570
rect 2335 18480 2365 18510
rect 2335 18415 2365 18445
rect 2335 18345 2365 18375
rect 2335 18275 2365 18305
rect 2335 18205 2365 18235
rect 2335 18140 2365 18170
rect 2335 18080 2365 18110
rect 2335 18015 2365 18045
rect 2335 17945 2365 17975
rect 2335 17875 2365 17905
rect 2335 17805 2365 17835
rect 2335 17740 2365 17770
rect 6705 20880 6735 20910
rect 6705 20815 6735 20845
rect 6705 20745 6735 20775
rect 6705 20675 6735 20705
rect 6705 20605 6735 20635
rect 6705 20540 6735 20570
rect 6705 20480 6735 20510
rect 6705 20415 6735 20445
rect 6705 20345 6735 20375
rect 6705 20275 6735 20305
rect 6705 20205 6735 20235
rect 6705 20140 6735 20170
rect 6705 20080 6735 20110
rect 6705 20015 6735 20045
rect 6705 19945 6735 19975
rect 6705 19875 6735 19905
rect 6705 19805 6735 19835
rect 6705 19740 6735 19770
rect 6705 19680 6735 19710
rect 6705 19615 6735 19645
rect 6705 19545 6735 19575
rect 6705 19475 6735 19505
rect 6705 19405 6735 19435
rect 6705 19340 6735 19370
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 2335 15750 2365 15780
rect 2335 12730 2365 12760
rect 2335 12690 2365 12720
rect 2335 12570 2365 12600
rect 2335 12530 2365 12560
rect 2335 12490 2365 12520
rect 2390 15895 2420 15925
rect 6705 15675 6735 15705
rect 6705 12975 6735 13005
rect 6705 12935 6735 12965
rect 6705 12895 6735 12925
rect 6595 12170 6625 12200
rect 6595 12130 6625 12160
rect 6595 12090 6625 12120
rect 6305 11455 6335 11485
rect 6305 11415 6335 11445
rect 6305 11375 6335 11405
rect 2995 10055 3025 10085
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 1325 8065 1355 8095
rect 1325 8005 1355 8035
rect 1325 7940 1355 7970
rect 1325 7870 1355 7900
rect 1325 7800 1355 7830
rect 1325 7730 1355 7760
rect 1325 7665 1355 7695
rect 1325 7605 1355 7635
rect 1325 7540 1355 7570
rect 1325 7470 1355 7500
rect 1325 7400 1355 7430
rect 1325 7330 1355 7360
rect 1325 7265 1355 7295
rect 1325 7205 1355 7235
rect 1325 7140 1355 7170
rect 1325 7070 1355 7100
rect 1325 7000 1355 7030
rect 1325 6930 1355 6960
rect 1325 6865 1355 6895
rect 1325 6805 1355 6835
rect 1325 6740 1355 6770
rect 1325 6670 1355 6700
rect 1325 6600 1355 6630
rect 1325 6530 1355 6560
rect 1325 6465 1355 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 2390 9605 2420 9635
rect 2390 9540 2420 9570
rect 2390 9470 2420 9500
rect 2390 9400 2420 9430
rect 2390 9330 2420 9360
rect 2390 9265 2420 9295
rect 2390 9205 2420 9235
rect 2390 9140 2420 9170
rect 2390 9070 2420 9100
rect 2390 9000 2420 9030
rect 2390 8930 2420 8960
rect 2390 8865 2420 8895
rect 2390 8805 2420 8835
rect 2390 8740 2420 8770
rect 2390 8670 2420 8700
rect 2390 8600 2420 8630
rect 2390 8530 2420 8560
rect 2390 8465 2420 8495
rect 2390 8405 2420 8435
rect 2390 8340 2420 8370
rect 2390 8270 2420 8300
rect 2390 8200 2420 8230
rect 2390 8130 2420 8160
rect 2390 8065 2420 8095
rect 2390 8005 2420 8035
rect 2390 7940 2420 7970
rect 2390 7870 2420 7900
rect 2390 7800 2420 7830
rect 2390 7730 2420 7760
rect 2390 7665 2420 7695
rect 2390 7605 2420 7635
rect 2390 7540 2420 7570
rect 2390 7470 2420 7500
rect 2390 7400 2420 7430
rect 2390 7330 2420 7360
rect 2390 7265 2420 7295
rect 2390 7205 2420 7235
rect 2390 7140 2420 7170
rect 2390 7070 2420 7100
rect 2390 7000 2420 7030
rect 2390 6930 2420 6960
rect 2390 6865 2420 6895
rect 2390 6805 2420 6835
rect 2390 6740 2420 6770
rect 2390 6670 2420 6700
rect 2390 6600 2420 6630
rect 2390 6530 2420 6560
rect 2390 6465 2420 6495
rect 2050 6400 2080 6430
rect 2480 6400 2510 6430
rect 2005 6345 2035 6375
rect 1285 6175 1315 6205
rect 1325 6175 1355 6205
rect 1365 6175 1395 6205
rect 1285 6135 1315 6165
rect 1325 6135 1355 6165
rect 1365 6135 1395 6165
rect 1285 6095 1315 6125
rect 1325 6095 1355 6125
rect 1365 6095 1395 6125
rect 2850 6410 2880 6440
rect 2720 6300 2750 6330
rect 3240 9605 3270 9635
rect 3240 9540 3270 9570
rect 3240 9470 3270 9500
rect 3240 9400 3270 9430
rect 3240 9330 3270 9360
rect 3240 9265 3270 9295
rect 3240 9205 3270 9235
rect 3240 9140 3270 9170
rect 3240 9070 3270 9100
rect 3240 9000 3270 9030
rect 3240 8930 3270 8960
rect 3240 8865 3270 8895
rect 3240 8805 3270 8835
rect 3240 8740 3270 8770
rect 3240 8670 3270 8700
rect 3240 8600 3270 8630
rect 3240 8530 3270 8560
rect 3240 8465 3270 8495
rect 3240 8405 3270 8435
rect 3240 8340 3270 8370
rect 3240 8270 3270 8300
rect 3240 8200 3270 8230
rect 3240 8130 3270 8160
rect 3240 8065 3270 8095
rect 3240 8005 3270 8035
rect 3240 7940 3270 7970
rect 3240 7870 3270 7900
rect 3240 7800 3270 7830
rect 3240 7730 3270 7760
rect 3240 7665 3270 7695
rect 3240 7605 3270 7635
rect 3240 7540 3270 7570
rect 3240 7470 3270 7500
rect 3240 7400 3270 7430
rect 3240 7330 3270 7360
rect 3240 7265 3270 7295
rect 3240 7205 3270 7235
rect 3240 7140 3270 7170
rect 3240 7070 3270 7100
rect 3240 7000 3270 7030
rect 3240 6930 3270 6960
rect 3240 6865 3270 6895
rect 3240 6805 3270 6835
rect 3240 6740 3270 6770
rect 3240 6670 3270 6700
rect 3240 6600 3270 6630
rect 3240 6530 3270 6560
rect 3240 6465 3270 6495
rect 3405 6410 3435 6440
rect 2995 6255 3025 6285
rect 3635 6345 3665 6375
rect 3460 6255 3490 6285
rect 3405 3025 3435 3055
rect 4310 6175 4340 6205
rect 4310 6135 4340 6165
rect 4310 6095 4340 6125
rect 4420 6175 4450 6205
rect 4420 6135 4450 6165
rect 4420 6095 4450 6125
rect 4530 6175 4560 6205
rect 4530 6135 4560 6165
rect 4530 6095 4560 6125
rect 5650 9605 5680 9635
rect 5650 9540 5680 9570
rect 5650 9470 5680 9500
rect 5650 9400 5680 9430
rect 5650 9330 5680 9360
rect 5650 9265 5680 9295
rect 5650 9205 5680 9235
rect 5650 9140 5680 9170
rect 5650 9070 5680 9100
rect 5650 9000 5680 9030
rect 5650 8930 5680 8960
rect 5650 8865 5680 8895
rect 5650 8805 5680 8835
rect 5650 8740 5680 8770
rect 5650 8670 5680 8700
rect 5650 8600 5680 8630
rect 5650 8530 5680 8560
rect 5650 8465 5680 8495
rect 5650 8405 5680 8435
rect 5650 8340 5680 8370
rect 5650 8270 5680 8300
rect 5650 8200 5680 8230
rect 5650 8130 5680 8160
rect 5650 8065 5680 8095
rect 5650 8005 5680 8035
rect 5650 7940 5680 7970
rect 5650 7870 5680 7900
rect 5650 7800 5680 7830
rect 5650 7730 5680 7760
rect 5650 7665 5680 7695
rect 5650 7605 5680 7635
rect 5650 7540 5680 7570
rect 5650 7470 5680 7500
rect 5650 7400 5680 7430
rect 5650 7330 5680 7360
rect 5650 7265 5680 7295
rect 5650 7205 5680 7235
rect 5650 7140 5680 7170
rect 5650 7070 5680 7100
rect 5650 7000 5680 7030
rect 5650 6930 5680 6960
rect 5650 6865 5680 6895
rect 5650 6805 5680 6835
rect 5650 6740 5680 6770
rect 5650 6670 5680 6700
rect 5650 6600 5680 6630
rect 5650 6530 5680 6560
rect 5650 6465 5680 6495
rect 5495 6400 5525 6430
rect 6150 6400 6180 6430
rect 5315 6345 5345 6375
rect 4855 6300 4885 6330
rect 4640 6175 4670 6205
rect 4640 6135 4670 6165
rect 4640 6095 4670 6125
rect 4855 4985 4885 5015
rect 4945 4985 4975 5015
rect 5166 4525 5196 4555
rect 4945 4470 4975 4500
rect 6305 9605 6335 9635
rect 6305 9540 6335 9570
rect 6305 9470 6335 9500
rect 6305 9400 6335 9430
rect 6305 9330 6335 9360
rect 6305 9265 6335 9295
rect 6305 9205 6335 9235
rect 6305 9140 6335 9170
rect 6305 9070 6335 9100
rect 6305 9000 6335 9030
rect 6305 8930 6335 8960
rect 6305 8865 6335 8895
rect 6305 8805 6335 8835
rect 6305 8740 6335 8770
rect 6305 8670 6335 8700
rect 6305 8600 6335 8630
rect 6305 8530 6335 8560
rect 6305 8465 6335 8495
rect 6305 8405 6335 8435
rect 6305 8340 6335 8370
rect 6305 8270 6335 8300
rect 6305 8200 6335 8230
rect 6305 8130 6335 8160
rect 6305 8065 6335 8095
rect 6305 8005 6335 8035
rect 6305 7940 6335 7970
rect 6305 7870 6335 7900
rect 6305 7800 6335 7830
rect 6305 7730 6335 7760
rect 6305 7665 6335 7695
rect 6305 7605 6335 7635
rect 6305 7540 6335 7570
rect 6305 7470 6335 7500
rect 6305 7400 6335 7430
rect 6305 7330 6335 7360
rect 6305 7265 6335 7295
rect 6305 7205 6335 7235
rect 6305 7140 6335 7170
rect 6305 7070 6335 7100
rect 6305 7000 6335 7030
rect 6305 6930 6335 6960
rect 6305 6865 6335 6895
rect 6305 6805 6335 6835
rect 6305 6740 6335 6770
rect 6305 6670 6335 6700
rect 6305 6600 6335 6630
rect 6305 6530 6335 6560
rect 6305 6465 6335 6495
rect 6595 9605 6625 9635
rect 6595 9540 6625 9570
rect 6595 9470 6625 9500
rect 6595 9400 6625 9430
rect 6595 9330 6625 9360
rect 6595 9265 6625 9295
rect 6595 9205 6625 9235
rect 6595 9140 6625 9170
rect 6595 9070 6625 9100
rect 6595 9000 6625 9030
rect 6595 8930 6625 8960
rect 6595 8865 6625 8895
rect 6595 8805 6625 8835
rect 6595 8740 6625 8770
rect 6595 8670 6625 8700
rect 6595 8600 6625 8630
rect 6595 8530 6625 8560
rect 6595 8465 6625 8495
rect 6595 8405 6625 8435
rect 6595 8340 6625 8370
rect 6595 8270 6625 8300
rect 6595 8200 6625 8230
rect 6595 8130 6625 8160
rect 6595 8065 6625 8095
rect 6595 8005 6625 8035
rect 6595 7940 6625 7970
rect 6595 7870 6625 7900
rect 6595 7800 6625 7830
rect 6595 7730 6625 7760
rect 6595 7665 6625 7695
rect 6595 7605 6625 7635
rect 6595 7540 6625 7570
rect 6595 7470 6625 7500
rect 6595 7400 6625 7430
rect 6595 7330 6625 7360
rect 6595 7265 6625 7295
rect 6595 7205 6625 7235
rect 6595 7140 6625 7170
rect 6595 7070 6625 7100
rect 6595 7000 6625 7030
rect 6595 6930 6625 6960
rect 6595 6865 6625 6895
rect 6595 6805 6625 6835
rect 6595 6740 6625 6770
rect 6595 6670 6625 6700
rect 6595 6600 6625 6630
rect 6595 6530 6625 6560
rect 6595 6465 6625 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 6470 6400 6500 6430
rect 6900 6400 6930 6430
rect 5875 5105 5905 5135
rect 6225 5105 6255 5135
rect 5875 4535 5905 4565
rect 5495 3090 5525 3120
rect 6945 6345 6975 6375
rect 2050 1725 2080 1755
rect 2180 1725 2210 1755
rect 6770 1725 6800 1755
rect 6900 1725 6930 1755
rect 2005 1670 2035 1700
rect 2105 1670 2135 1700
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect 7625 8065 7655 8095
rect 7625 8005 7655 8035
rect 7625 7940 7655 7970
rect 7625 7870 7655 7900
rect 7625 7800 7655 7830
rect 7625 7730 7655 7760
rect 7625 7665 7655 7695
rect 7625 7605 7655 7635
rect 7625 7540 7655 7570
rect 7625 7470 7655 7500
rect 7625 7400 7655 7430
rect 7625 7330 7655 7360
rect 7625 7265 7655 7295
rect 7625 7205 7655 7235
rect 7625 7140 7655 7170
rect 7625 7070 7655 7100
rect 7625 7000 7655 7030
rect 7625 6930 7655 6960
rect 7625 6865 7655 6895
rect 7625 6805 7655 6835
rect 7625 6740 7655 6770
rect 7625 6670 7655 6700
rect 7625 6600 7655 6630
rect 7625 6530 7655 6560
rect 7625 6465 7655 6495
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect 7585 6175 7615 6205
rect 7625 6175 7655 6205
rect 7665 6175 7695 6205
rect 7585 6135 7615 6165
rect 7625 6135 7655 6165
rect 7665 6135 7695 6165
rect 7585 6095 7615 6125
rect 7625 6095 7655 6125
rect 7665 6095 7695 6125
rect 6835 1670 6865 1700
rect 6945 1670 6975 1700
rect 1285 820 1315 850
rect 1325 820 1355 850
rect 1365 820 1395 850
rect 1285 780 1315 810
rect 1325 780 1355 810
rect 1365 780 1395 810
rect 1285 740 1315 770
rect 1325 740 1355 770
rect 1365 740 1395 770
rect 4420 820 4450 850
rect 4475 820 4505 850
rect 4530 820 4560 850
rect 4420 780 4450 810
rect 4475 780 4505 810
rect 4530 780 4560 810
rect 4420 740 4450 770
rect 4475 740 4505 770
rect 4530 740 4560 770
rect 7585 820 7615 850
rect 7625 820 7655 850
rect 7665 820 7695 850
rect 7585 780 7615 810
rect 7625 780 7655 810
rect 7665 780 7695 810
rect 7585 740 7615 770
rect 7625 740 7655 770
rect 7665 740 7695 770
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect -75 -2935 -45 -2905
rect -75 -3000 -45 -2970
rect -75 -3070 -45 -3040
rect -75 -3140 -45 -3110
rect -75 -3210 -45 -3180
rect -75 -3275 -45 -3245
rect -75 -3335 -45 -3305
rect -75 -3400 -45 -3370
rect -75 -3470 -45 -3440
rect -75 -3540 -45 -3510
rect -75 -3610 -45 -3580
rect -75 -3675 -45 -3645
rect -75 -3735 -45 -3705
rect -75 -3800 -45 -3770
rect -75 -3870 -45 -3840
rect -75 -3940 -45 -3910
rect -75 -4010 -45 -3980
rect -75 -4075 -45 -4045
rect -75 -4135 -45 -4105
rect -75 -4200 -45 -4170
rect -75 -4270 -45 -4240
rect -75 -4340 -45 -4310
rect -75 -4410 -45 -4380
rect -75 -4475 -45 -4445
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 275 -2935 305 -2905
rect 275 -3000 305 -2970
rect 275 -3070 305 -3040
rect 275 -3140 305 -3110
rect 275 -3210 305 -3180
rect 275 -3275 305 -3245
rect 275 -3335 305 -3305
rect 275 -3400 305 -3370
rect 275 -3470 305 -3440
rect 275 -3540 305 -3510
rect 275 -3610 305 -3580
rect 275 -3675 305 -3645
rect 275 -3735 305 -3705
rect 275 -3800 305 -3770
rect 275 -3870 305 -3840
rect 275 -3940 305 -3910
rect 275 -4010 305 -3980
rect 275 -4075 305 -4045
rect 275 -4135 305 -4105
rect 275 -4200 305 -4170
rect 275 -4270 305 -4240
rect 275 -4340 305 -4310
rect 275 -4410 305 -4380
rect 275 -4475 305 -4445
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 625 -2935 655 -2905
rect 625 -3000 655 -2970
rect 625 -3070 655 -3040
rect 625 -3140 655 -3110
rect 625 -3210 655 -3180
rect 625 -3275 655 -3245
rect 625 -3335 655 -3305
rect 625 -3400 655 -3370
rect 625 -3470 655 -3440
rect 625 -3540 655 -3510
rect 625 -3610 655 -3580
rect 625 -3675 655 -3645
rect 625 -3735 655 -3705
rect 625 -3800 655 -3770
rect 625 -3870 655 -3840
rect 625 -3940 655 -3910
rect 625 -4010 655 -3980
rect 625 -4075 655 -4045
rect 625 -4135 655 -4105
rect 625 -4200 655 -4170
rect 625 -4270 655 -4240
rect 625 -4340 655 -4310
rect 625 -4410 655 -4380
rect 625 -4475 655 -4445
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 975 -2935 1005 -2905
rect 975 -3000 1005 -2970
rect 975 -3070 1005 -3040
rect 975 -3140 1005 -3110
rect 975 -3210 1005 -3180
rect 975 -3275 1005 -3245
rect 975 -3335 1005 -3305
rect 975 -3400 1005 -3370
rect 975 -3470 1005 -3440
rect 975 -3540 1005 -3510
rect 975 -3610 1005 -3580
rect 975 -3675 1005 -3645
rect 975 -3735 1005 -3705
rect 975 -3800 1005 -3770
rect 975 -3870 1005 -3840
rect 975 -3940 1005 -3910
rect 975 -4010 1005 -3980
rect 975 -4075 1005 -4045
rect 975 -4135 1005 -4105
rect 975 -4200 1005 -4170
rect 975 -4270 1005 -4240
rect 975 -4340 1005 -4310
rect 975 -4410 1005 -4380
rect 975 -4475 1005 -4445
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1325 -2935 1355 -2905
rect 1325 -3000 1355 -2970
rect 1325 -3070 1355 -3040
rect 1325 -3140 1355 -3110
rect 1325 -3210 1355 -3180
rect 1325 -3275 1355 -3245
rect 1325 -3335 1355 -3305
rect 1325 -3400 1355 -3370
rect 1325 -3470 1355 -3440
rect 1325 -3540 1355 -3510
rect 1325 -3610 1355 -3580
rect 1325 -3675 1355 -3645
rect 1325 -3735 1355 -3705
rect 1325 -3800 1355 -3770
rect 1325 -3870 1355 -3840
rect 1325 -3940 1355 -3910
rect 1325 -4010 1355 -3980
rect 1325 -4075 1355 -4045
rect 1325 -4135 1355 -4105
rect 1325 -4200 1355 -4170
rect 1325 -4270 1355 -4240
rect 1325 -4340 1355 -4310
rect 1325 -4410 1355 -4380
rect 1325 -4475 1355 -4445
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 1675 -2935 1705 -2905
rect 1675 -3000 1705 -2970
rect 1675 -3070 1705 -3040
rect 1675 -3140 1705 -3110
rect 1675 -3210 1705 -3180
rect 1675 -3275 1705 -3245
rect 1675 -3335 1705 -3305
rect 1675 -3400 1705 -3370
rect 1675 -3470 1705 -3440
rect 1675 -3540 1705 -3510
rect 1675 -3610 1705 -3580
rect 1675 -3675 1705 -3645
rect 1675 -3735 1705 -3705
rect 1675 -3800 1705 -3770
rect 1675 -3870 1705 -3840
rect 1675 -3940 1705 -3910
rect 1675 -4010 1705 -3980
rect 1675 -4075 1705 -4045
rect 1675 -4135 1705 -4105
rect 1675 -4200 1705 -4170
rect 1675 -4270 1705 -4240
rect 1675 -4340 1705 -4310
rect 1675 -4410 1705 -4380
rect 1675 -4475 1705 -4445
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2025 -2935 2055 -2905
rect 2025 -3000 2055 -2970
rect 2025 -3070 2055 -3040
rect 2025 -3140 2055 -3110
rect 2025 -3210 2055 -3180
rect 2025 -3275 2055 -3245
rect 2025 -3335 2055 -3305
rect 2025 -3400 2055 -3370
rect 2025 -3470 2055 -3440
rect 2025 -3540 2055 -3510
rect 2025 -3610 2055 -3580
rect 2025 -3675 2055 -3645
rect 2025 -3735 2055 -3705
rect 2025 -3800 2055 -3770
rect 2025 -3870 2055 -3840
rect 2025 -3940 2055 -3910
rect 2025 -4010 2055 -3980
rect 2025 -4075 2055 -4045
rect 2025 -4135 2055 -4105
rect 2025 -4200 2055 -4170
rect 2025 -4270 2055 -4240
rect 2025 -4340 2055 -4310
rect 2025 -4410 2055 -4380
rect 2025 -4475 2055 -4445
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2375 -2935 2405 -2905
rect 2375 -3000 2405 -2970
rect 2375 -3070 2405 -3040
rect 2375 -3140 2405 -3110
rect 2375 -3210 2405 -3180
rect 2375 -3275 2405 -3245
rect 2375 -3335 2405 -3305
rect 2375 -3400 2405 -3370
rect 2375 -3470 2405 -3440
rect 2375 -3540 2405 -3510
rect 2375 -3610 2405 -3580
rect 2375 -3675 2405 -3645
rect 2375 -3735 2405 -3705
rect 2375 -3800 2405 -3770
rect 2375 -3870 2405 -3840
rect 2375 -3940 2405 -3910
rect 2375 -4010 2405 -3980
rect 2375 -4075 2405 -4045
rect 2375 -4135 2405 -4105
rect 2375 -4200 2405 -4170
rect 2375 -4270 2405 -4240
rect 2375 -4340 2405 -4310
rect 2375 -4410 2405 -4380
rect 2375 -4475 2405 -4445
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 2725 -2935 2755 -2905
rect 2725 -3000 2755 -2970
rect 2725 -3070 2755 -3040
rect 2725 -3140 2755 -3110
rect 2725 -3210 2755 -3180
rect 2725 -3275 2755 -3245
rect 2725 -3335 2755 -3305
rect 2725 -3400 2755 -3370
rect 2725 -3470 2755 -3440
rect 2725 -3540 2755 -3510
rect 2725 -3610 2755 -3580
rect 2725 -3675 2755 -3645
rect 2725 -3735 2755 -3705
rect 2725 -3800 2755 -3770
rect 2725 -3870 2755 -3840
rect 2725 -3940 2755 -3910
rect 2725 -4010 2755 -3980
rect 2725 -4075 2755 -4045
rect 2725 -4135 2755 -4105
rect 2725 -4200 2755 -4170
rect 2725 -4270 2755 -4240
rect 2725 -4340 2755 -4310
rect 2725 -4410 2755 -4380
rect 2725 -4475 2755 -4445
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3075 -2935 3105 -2905
rect 3075 -3000 3105 -2970
rect 3075 -3070 3105 -3040
rect 3075 -3140 3105 -3110
rect 3075 -3210 3105 -3180
rect 3075 -3275 3105 -3245
rect 3075 -3335 3105 -3305
rect 3075 -3400 3105 -3370
rect 3075 -3470 3105 -3440
rect 3075 -3540 3105 -3510
rect 3075 -3610 3105 -3580
rect 3075 -3675 3105 -3645
rect 3075 -3735 3105 -3705
rect 3075 -3800 3105 -3770
rect 3075 -3870 3105 -3840
rect 3075 -3940 3105 -3910
rect 3075 -4010 3105 -3980
rect 3075 -4075 3105 -4045
rect 3075 -4135 3105 -4105
rect 3075 -4200 3105 -4170
rect 3075 -4270 3105 -4240
rect 3075 -4340 3105 -4310
rect 3075 -4410 3105 -4380
rect 3075 -4475 3105 -4445
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3425 -2935 3455 -2905
rect 3425 -3000 3455 -2970
rect 3425 -3070 3455 -3040
rect 3425 -3140 3455 -3110
rect 3425 -3210 3455 -3180
rect 3425 -3275 3455 -3245
rect 3425 -3335 3455 -3305
rect 3425 -3400 3455 -3370
rect 3425 -3470 3455 -3440
rect 3425 -3540 3455 -3510
rect 3425 -3610 3455 -3580
rect 3425 -3675 3455 -3645
rect 3425 -3735 3455 -3705
rect 3425 -3800 3455 -3770
rect 3425 -3870 3455 -3840
rect 3425 -3940 3455 -3910
rect 3425 -4010 3455 -3980
rect 3425 -4075 3455 -4045
rect 3425 -4135 3455 -4105
rect 3425 -4200 3455 -4170
rect 3425 -4270 3455 -4240
rect 3425 -4340 3455 -4310
rect 3425 -4410 3455 -4380
rect 3425 -4475 3455 -4445
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 3775 -2935 3805 -2905
rect 3775 -3000 3805 -2970
rect 3775 -3070 3805 -3040
rect 3775 -3140 3805 -3110
rect 3775 -3210 3805 -3180
rect 3775 -3275 3805 -3245
rect 3775 -3335 3805 -3305
rect 3775 -3400 3805 -3370
rect 3775 -3470 3805 -3440
rect 3775 -3540 3805 -3510
rect 3775 -3610 3805 -3580
rect 3775 -3675 3805 -3645
rect 3775 -3735 3805 -3705
rect 3775 -3800 3805 -3770
rect 3775 -3870 3805 -3840
rect 3775 -3940 3805 -3910
rect 3775 -4010 3805 -3980
rect 3775 -4075 3805 -4045
rect 3775 -4135 3805 -4105
rect 3775 -4200 3805 -4170
rect 3775 -4270 3805 -4240
rect 3775 -4340 3805 -4310
rect 3775 -4410 3805 -4380
rect 3775 -4475 3805 -4445
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4125 -2935 4155 -2905
rect 4125 -3000 4155 -2970
rect 4125 -3070 4155 -3040
rect 4125 -3140 4155 -3110
rect 4125 -3210 4155 -3180
rect 4125 -3275 4155 -3245
rect 4125 -3335 4155 -3305
rect 4125 -3400 4155 -3370
rect 4125 -3470 4155 -3440
rect 4125 -3540 4155 -3510
rect 4125 -3610 4155 -3580
rect 4125 -3675 4155 -3645
rect 4125 -3735 4155 -3705
rect 4125 -3800 4155 -3770
rect 4125 -3870 4155 -3840
rect 4125 -3940 4155 -3910
rect 4125 -4010 4155 -3980
rect 4125 -4075 4155 -4045
rect 4125 -4135 4155 -4105
rect 4125 -4200 4155 -4170
rect 4125 -4270 4155 -4240
rect 4125 -4340 4155 -4310
rect 4125 -4410 4155 -4380
rect 4125 -4475 4155 -4445
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4475 -2935 4505 -2905
rect 4475 -3000 4505 -2970
rect 4475 -3070 4505 -3040
rect 4475 -3140 4505 -3110
rect 4475 -3210 4505 -3180
rect 4475 -3275 4505 -3245
rect 4475 -3335 4505 -3305
rect 4475 -3400 4505 -3370
rect 4475 -3470 4505 -3440
rect 4475 -3540 4505 -3510
rect 4475 -3610 4505 -3580
rect 4475 -3675 4505 -3645
rect 4475 -3735 4505 -3705
rect 4475 -3800 4505 -3770
rect 4475 -3870 4505 -3840
rect 4475 -3940 4505 -3910
rect 4475 -4010 4505 -3980
rect 4475 -4075 4505 -4045
rect 4475 -4135 4505 -4105
rect 4475 -4200 4505 -4170
rect 4475 -4270 4505 -4240
rect 4475 -4340 4505 -4310
rect 4475 -4410 4505 -4380
rect 4475 -4475 4505 -4445
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 4825 -2935 4855 -2905
rect 4825 -3000 4855 -2970
rect 4825 -3070 4855 -3040
rect 4825 -3140 4855 -3110
rect 4825 -3210 4855 -3180
rect 4825 -3275 4855 -3245
rect 4825 -3335 4855 -3305
rect 4825 -3400 4855 -3370
rect 4825 -3470 4855 -3440
rect 4825 -3540 4855 -3510
rect 4825 -3610 4855 -3580
rect 4825 -3675 4855 -3645
rect 4825 -3735 4855 -3705
rect 4825 -3800 4855 -3770
rect 4825 -3870 4855 -3840
rect 4825 -3940 4855 -3910
rect 4825 -4010 4855 -3980
rect 4825 -4075 4855 -4045
rect 4825 -4135 4855 -4105
rect 4825 -4200 4855 -4170
rect 4825 -4270 4855 -4240
rect 4825 -4340 4855 -4310
rect 4825 -4410 4855 -4380
rect 4825 -4475 4855 -4445
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5175 -2935 5205 -2905
rect 5175 -3000 5205 -2970
rect 5175 -3070 5205 -3040
rect 5175 -3140 5205 -3110
rect 5175 -3210 5205 -3180
rect 5175 -3275 5205 -3245
rect 5175 -3335 5205 -3305
rect 5175 -3400 5205 -3370
rect 5175 -3470 5205 -3440
rect 5175 -3540 5205 -3510
rect 5175 -3610 5205 -3580
rect 5175 -3675 5205 -3645
rect 5175 -3735 5205 -3705
rect 5175 -3800 5205 -3770
rect 5175 -3870 5205 -3840
rect 5175 -3940 5205 -3910
rect 5175 -4010 5205 -3980
rect 5175 -4075 5205 -4045
rect 5175 -4135 5205 -4105
rect 5175 -4200 5205 -4170
rect 5175 -4270 5205 -4240
rect 5175 -4340 5205 -4310
rect 5175 -4410 5205 -4380
rect 5175 -4475 5205 -4445
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5525 -2935 5555 -2905
rect 5525 -3000 5555 -2970
rect 5525 -3070 5555 -3040
rect 5525 -3140 5555 -3110
rect 5525 -3210 5555 -3180
rect 5525 -3275 5555 -3245
rect 5525 -3335 5555 -3305
rect 5525 -3400 5555 -3370
rect 5525 -3470 5555 -3440
rect 5525 -3540 5555 -3510
rect 5525 -3610 5555 -3580
rect 5525 -3675 5555 -3645
rect 5525 -3735 5555 -3705
rect 5525 -3800 5555 -3770
rect 5525 -3870 5555 -3840
rect 5525 -3940 5555 -3910
rect 5525 -4010 5555 -3980
rect 5525 -4075 5555 -4045
rect 5525 -4135 5555 -4105
rect 5525 -4200 5555 -4170
rect 5525 -4270 5555 -4240
rect 5525 -4340 5555 -4310
rect 5525 -4410 5555 -4380
rect 5525 -4475 5555 -4445
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 5875 -2935 5905 -2905
rect 5875 -3000 5905 -2970
rect 5875 -3070 5905 -3040
rect 5875 -3140 5905 -3110
rect 5875 -3210 5905 -3180
rect 5875 -3275 5905 -3245
rect 5875 -3335 5905 -3305
rect 5875 -3400 5905 -3370
rect 5875 -3470 5905 -3440
rect 5875 -3540 5905 -3510
rect 5875 -3610 5905 -3580
rect 5875 -3675 5905 -3645
rect 5875 -3735 5905 -3705
rect 5875 -3800 5905 -3770
rect 5875 -3870 5905 -3840
rect 5875 -3940 5905 -3910
rect 5875 -4010 5905 -3980
rect 5875 -4075 5905 -4045
rect 5875 -4135 5905 -4105
rect 5875 -4200 5905 -4170
rect 5875 -4270 5905 -4240
rect 5875 -4340 5905 -4310
rect 5875 -4410 5905 -4380
rect 5875 -4475 5905 -4445
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6225 -2935 6255 -2905
rect 6225 -3000 6255 -2970
rect 6225 -3070 6255 -3040
rect 6225 -3140 6255 -3110
rect 6225 -3210 6255 -3180
rect 6225 -3275 6255 -3245
rect 6225 -3335 6255 -3305
rect 6225 -3400 6255 -3370
rect 6225 -3470 6255 -3440
rect 6225 -3540 6255 -3510
rect 6225 -3610 6255 -3580
rect 6225 -3675 6255 -3645
rect 6225 -3735 6255 -3705
rect 6225 -3800 6255 -3770
rect 6225 -3870 6255 -3840
rect 6225 -3940 6255 -3910
rect 6225 -4010 6255 -3980
rect 6225 -4075 6255 -4045
rect 6225 -4135 6255 -4105
rect 6225 -4200 6255 -4170
rect 6225 -4270 6255 -4240
rect 6225 -4340 6255 -4310
rect 6225 -4410 6255 -4380
rect 6225 -4475 6255 -4445
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6575 -2935 6605 -2905
rect 6575 -3000 6605 -2970
rect 6575 -3070 6605 -3040
rect 6575 -3140 6605 -3110
rect 6575 -3210 6605 -3180
rect 6575 -3275 6605 -3245
rect 6575 -3335 6605 -3305
rect 6575 -3400 6605 -3370
rect 6575 -3470 6605 -3440
rect 6575 -3540 6605 -3510
rect 6575 -3610 6605 -3580
rect 6575 -3675 6605 -3645
rect 6575 -3735 6605 -3705
rect 6575 -3800 6605 -3770
rect 6575 -3870 6605 -3840
rect 6575 -3940 6605 -3910
rect 6575 -4010 6605 -3980
rect 6575 -4075 6605 -4045
rect 6575 -4135 6605 -4105
rect 6575 -4200 6605 -4170
rect 6575 -4270 6605 -4240
rect 6575 -4340 6605 -4310
rect 6575 -4410 6605 -4380
rect 6575 -4475 6605 -4445
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 6925 -2935 6955 -2905
rect 6925 -3000 6955 -2970
rect 6925 -3070 6955 -3040
rect 6925 -3140 6955 -3110
rect 6925 -3210 6955 -3180
rect 6925 -3275 6955 -3245
rect 6925 -3335 6955 -3305
rect 6925 -3400 6955 -3370
rect 6925 -3470 6955 -3440
rect 6925 -3540 6955 -3510
rect 6925 -3610 6955 -3580
rect 6925 -3675 6955 -3645
rect 6925 -3735 6955 -3705
rect 6925 -3800 6955 -3770
rect 6925 -3870 6955 -3840
rect 6925 -3940 6955 -3910
rect 6925 -4010 6955 -3980
rect 6925 -4075 6955 -4045
rect 6925 -4135 6955 -4105
rect 6925 -4200 6955 -4170
rect 6925 -4270 6955 -4240
rect 6925 -4340 6955 -4310
rect 6925 -4410 6955 -4380
rect 6925 -4475 6955 -4445
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7275 -2935 7305 -2905
rect 7275 -3000 7305 -2970
rect 7275 -3070 7305 -3040
rect 7275 -3140 7305 -3110
rect 7275 -3210 7305 -3180
rect 7275 -3275 7305 -3245
rect 7275 -3335 7305 -3305
rect 7275 -3400 7305 -3370
rect 7275 -3470 7305 -3440
rect 7275 -3540 7305 -3510
rect 7275 -3610 7305 -3580
rect 7275 -3675 7305 -3645
rect 7275 -3735 7305 -3705
rect 7275 -3800 7305 -3770
rect 7275 -3870 7305 -3840
rect 7275 -3940 7305 -3910
rect 7275 -4010 7305 -3980
rect 7275 -4075 7305 -4045
rect 7275 -4135 7305 -4105
rect 7275 -4200 7305 -4170
rect 7275 -4270 7305 -4240
rect 7275 -4340 7305 -4310
rect 7275 -4410 7305 -4380
rect 7275 -4475 7305 -4445
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7625 -2935 7655 -2905
rect 7625 -3000 7655 -2970
rect 7625 -3070 7655 -3040
rect 7625 -3140 7655 -3110
rect 7625 -3210 7655 -3180
rect 7625 -3275 7655 -3245
rect 7625 -3335 7655 -3305
rect 7625 -3400 7655 -3370
rect 7625 -3470 7655 -3440
rect 7625 -3540 7655 -3510
rect 7625 -3610 7655 -3580
rect 7625 -3675 7655 -3645
rect 7625 -3735 7655 -3705
rect 7625 -3800 7655 -3770
rect 7625 -3870 7655 -3840
rect 7625 -3940 7655 -3910
rect 7625 -4010 7655 -3980
rect 7625 -4075 7655 -4045
rect 7625 -4135 7655 -4105
rect 7625 -4200 7655 -4170
rect 7625 -4270 7655 -4240
rect 7625 -4340 7655 -4310
rect 7625 -4410 7655 -4380
rect 7625 -4475 7655 -4445
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 7975 -2935 8005 -2905
rect 7975 -3000 8005 -2970
rect 7975 -3070 8005 -3040
rect 7975 -3140 8005 -3110
rect 7975 -3210 8005 -3180
rect 7975 -3275 8005 -3245
rect 7975 -3335 8005 -3305
rect 7975 -3400 8005 -3370
rect 7975 -3470 8005 -3440
rect 7975 -3540 8005 -3510
rect 7975 -3610 8005 -3580
rect 7975 -3675 8005 -3645
rect 7975 -3735 8005 -3705
rect 7975 -3800 8005 -3770
rect 7975 -3870 8005 -3840
rect 7975 -3940 8005 -3910
rect 7975 -4010 8005 -3980
rect 7975 -4075 8005 -4045
rect 7975 -4135 8005 -4105
rect 7975 -4200 8005 -4170
rect 7975 -4270 8005 -4240
rect 7975 -4340 8005 -4310
rect 7975 -4410 8005 -4380
rect 7975 -4475 8005 -4445
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8325 -2935 8355 -2905
rect 8325 -3000 8355 -2970
rect 8325 -3070 8355 -3040
rect 8325 -3140 8355 -3110
rect 8325 -3210 8355 -3180
rect 8325 -3275 8355 -3245
rect 8325 -3335 8355 -3305
rect 8325 -3400 8355 -3370
rect 8325 -3470 8355 -3440
rect 8325 -3540 8355 -3510
rect 8325 -3610 8355 -3580
rect 8325 -3675 8355 -3645
rect 8325 -3735 8355 -3705
rect 8325 -3800 8355 -3770
rect 8325 -3870 8355 -3840
rect 8325 -3940 8355 -3910
rect 8325 -4010 8355 -3980
rect 8325 -4075 8355 -4045
rect 8325 -4135 8355 -4105
rect 8325 -4200 8355 -4170
rect 8325 -4270 8355 -4240
rect 8325 -4340 8355 -4310
rect 8325 -4410 8355 -4380
rect 8325 -4475 8355 -4445
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 8675 -2935 8705 -2905
rect 8675 -3000 8705 -2970
rect 8675 -3070 8705 -3040
rect 8675 -3140 8705 -3110
rect 8675 -3210 8705 -3180
rect 8675 -3275 8705 -3245
rect 8675 -3335 8705 -3305
rect 8675 -3400 8705 -3370
rect 8675 -3470 8705 -3440
rect 8675 -3540 8705 -3510
rect 8675 -3610 8705 -3580
rect 8675 -3675 8705 -3645
rect 8675 -3735 8705 -3705
rect 8675 -3800 8705 -3770
rect 8675 -3870 8705 -3840
rect 8675 -3940 8705 -3910
rect 8675 -4010 8705 -3980
rect 8675 -4075 8705 -4045
rect 8675 -4135 8705 -4105
rect 8675 -4200 8705 -4170
rect 8675 -4270 8705 -4240
rect 8675 -4340 8705 -4310
rect 8675 -4410 8705 -4380
rect 8675 -4475 8705 -4445
<< metal2 >>
rect 2320 20910 2380 20925
rect 2320 20880 2335 20910
rect 2365 20880 2380 20910
rect 2320 20845 2380 20880
rect 2320 20815 2335 20845
rect 2365 20815 2380 20845
rect 2320 20775 2380 20815
rect 2320 20745 2335 20775
rect 2365 20745 2380 20775
rect 2320 20705 2380 20745
rect 2320 20675 2335 20705
rect 2365 20675 2380 20705
rect 2320 20635 2380 20675
rect 2320 20605 2335 20635
rect 2365 20605 2380 20635
rect 2320 20570 2380 20605
rect 2320 20540 2335 20570
rect 2365 20540 2380 20570
rect 2320 20510 2380 20540
rect 2320 20480 2335 20510
rect 2365 20480 2380 20510
rect 2320 20445 2380 20480
rect 2320 20415 2335 20445
rect 2365 20415 2380 20445
rect 2320 20375 2380 20415
rect 2320 20345 2335 20375
rect 2365 20345 2380 20375
rect 2320 20305 2380 20345
rect 2320 20275 2335 20305
rect 2365 20275 2380 20305
rect 2320 20235 2380 20275
rect 2320 20205 2335 20235
rect 2365 20205 2380 20235
rect 2320 20170 2380 20205
rect 2320 20140 2335 20170
rect 2365 20140 2380 20170
rect 2320 20110 2380 20140
rect 2320 20080 2335 20110
rect 2365 20080 2380 20110
rect 2320 20045 2380 20080
rect 2320 20015 2335 20045
rect 2365 20015 2380 20045
rect 2320 19975 2380 20015
rect 2320 19945 2335 19975
rect 2365 19945 2380 19975
rect 2320 19905 2380 19945
rect 2320 19875 2335 19905
rect 2365 19875 2380 19905
rect 2320 19835 2380 19875
rect 2320 19805 2335 19835
rect 2365 19805 2380 19835
rect 2320 19770 2380 19805
rect 2320 19740 2335 19770
rect 2365 19740 2380 19770
rect 2320 19710 2380 19740
rect 2320 19680 2335 19710
rect 2365 19680 2380 19710
rect 2320 19645 2380 19680
rect 2320 19615 2335 19645
rect 2365 19615 2380 19645
rect 2320 19575 2380 19615
rect 2320 19545 2335 19575
rect 2365 19545 2380 19575
rect 2320 19505 2380 19545
rect 2320 19475 2335 19505
rect 2365 19475 2380 19505
rect 2320 19435 2380 19475
rect 2320 19405 2335 19435
rect 2365 19405 2380 19435
rect 2320 19370 2380 19405
rect 2320 19340 2335 19370
rect 2365 19340 2380 19370
rect 2320 19310 2380 19340
rect 2320 19280 2335 19310
rect 2365 19280 2380 19310
rect 2320 19245 2380 19280
rect 2320 19215 2335 19245
rect 2365 19215 2380 19245
rect 2320 19175 2380 19215
rect 2320 19145 2335 19175
rect 2365 19145 2380 19175
rect 2320 19105 2380 19145
rect 2320 19075 2335 19105
rect 2365 19075 2380 19105
rect 2320 19035 2380 19075
rect 2320 19005 2335 19035
rect 2365 19005 2380 19035
rect 2320 18970 2380 19005
rect 2320 18940 2335 18970
rect 2365 18940 2380 18970
rect 2320 18910 2380 18940
rect 2320 18880 2335 18910
rect 2365 18880 2380 18910
rect 2320 18845 2380 18880
rect 2320 18815 2335 18845
rect 2365 18815 2380 18845
rect 2320 18775 2380 18815
rect 2320 18745 2335 18775
rect 2365 18745 2380 18775
rect 2320 18705 2380 18745
rect 2320 18675 2335 18705
rect 2365 18675 2380 18705
rect 2320 18635 2380 18675
rect 2320 18605 2335 18635
rect 2365 18605 2380 18635
rect 2320 18570 2380 18605
rect 2320 18540 2335 18570
rect 2365 18540 2380 18570
rect 2320 18510 2380 18540
rect 2320 18480 2335 18510
rect 2365 18480 2380 18510
rect 2320 18445 2380 18480
rect 2320 18415 2335 18445
rect 2365 18415 2380 18445
rect 2320 18375 2380 18415
rect 2320 18345 2335 18375
rect 2365 18345 2380 18375
rect 2320 18305 2380 18345
rect 2320 18275 2335 18305
rect 2365 18275 2380 18305
rect 2320 18235 2380 18275
rect 2320 18205 2335 18235
rect 2365 18205 2380 18235
rect 2320 18170 2380 18205
rect 2320 18140 2335 18170
rect 2365 18140 2380 18170
rect 2320 18110 2380 18140
rect 2320 18080 2335 18110
rect 2365 18080 2380 18110
rect 2320 18045 2380 18080
rect 2320 18015 2335 18045
rect 2365 18015 2380 18045
rect 2320 17975 2380 18015
rect 2320 17945 2335 17975
rect 2365 17945 2380 17975
rect 2320 17905 2380 17945
rect 2320 17875 2335 17905
rect 2365 17875 2380 17905
rect 2320 17835 2380 17875
rect 2320 17805 2335 17835
rect 2365 17805 2380 17835
rect 2320 17770 2380 17805
rect 2320 17740 2335 17770
rect 2365 17740 2380 17770
rect 2320 17725 2380 17740
rect 6690 20910 6750 20925
rect 6690 20880 6705 20910
rect 6735 20880 6750 20910
rect 6690 20845 6750 20880
rect 6690 20815 6705 20845
rect 6735 20815 6750 20845
rect 6690 20775 6750 20815
rect 6690 20745 6705 20775
rect 6735 20745 6750 20775
rect 6690 20705 6750 20745
rect 6690 20675 6705 20705
rect 6735 20675 6750 20705
rect 6690 20635 6750 20675
rect 6690 20605 6705 20635
rect 6735 20605 6750 20635
rect 6690 20570 6750 20605
rect 6690 20540 6705 20570
rect 6735 20540 6750 20570
rect 6690 20510 6750 20540
rect 6690 20480 6705 20510
rect 6735 20480 6750 20510
rect 6690 20445 6750 20480
rect 6690 20415 6705 20445
rect 6735 20415 6750 20445
rect 6690 20375 6750 20415
rect 6690 20345 6705 20375
rect 6735 20345 6750 20375
rect 6690 20305 6750 20345
rect 6690 20275 6705 20305
rect 6735 20275 6750 20305
rect 6690 20235 6750 20275
rect 6690 20205 6705 20235
rect 6735 20205 6750 20235
rect 6690 20170 6750 20205
rect 6690 20140 6705 20170
rect 6735 20140 6750 20170
rect 6690 20110 6750 20140
rect 6690 20080 6705 20110
rect 6735 20080 6750 20110
rect 6690 20045 6750 20080
rect 6690 20015 6705 20045
rect 6735 20015 6750 20045
rect 6690 19975 6750 20015
rect 6690 19945 6705 19975
rect 6735 19945 6750 19975
rect 6690 19905 6750 19945
rect 6690 19875 6705 19905
rect 6735 19875 6750 19905
rect 6690 19835 6750 19875
rect 6690 19805 6705 19835
rect 6735 19805 6750 19835
rect 6690 19770 6750 19805
rect 6690 19740 6705 19770
rect 6735 19740 6750 19770
rect 6690 19710 6750 19740
rect 6690 19680 6705 19710
rect 6735 19680 6750 19710
rect 6690 19645 6750 19680
rect 6690 19615 6705 19645
rect 6735 19615 6750 19645
rect 6690 19575 6750 19615
rect 6690 19545 6705 19575
rect 6735 19545 6750 19575
rect 6690 19505 6750 19545
rect 6690 19475 6705 19505
rect 6735 19475 6750 19505
rect 6690 19435 6750 19475
rect 6690 19405 6705 19435
rect 6735 19405 6750 19435
rect 6690 19370 6750 19405
rect 6690 19340 6705 19370
rect 6735 19340 6750 19370
rect 6690 19310 6750 19340
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2385 15925 2425 15930
rect 2385 15895 2390 15925
rect 2420 15895 2425 15925
rect 2385 15890 2425 15895
rect 2330 15780 2370 15785
rect 2330 15750 2335 15780
rect 2365 15775 2370 15780
rect 2365 15755 2970 15775
rect 2365 15750 2370 15755
rect 2330 15745 2370 15750
rect 6700 15705 6740 15710
rect 6700 15700 6705 15705
rect 6625 15680 6705 15700
rect 6700 15675 6705 15680
rect 6735 15675 6740 15705
rect 6700 15670 6740 15675
rect 5750 13005 6740 13010
rect 5750 12975 6705 13005
rect 6735 12975 6740 13005
rect 5750 12965 6740 12975
rect 5750 12935 6705 12965
rect 6735 12935 6740 12965
rect 5750 12925 6740 12935
rect 5750 12895 6705 12925
rect 6735 12895 6740 12925
rect 5750 12890 6740 12895
rect 2330 12760 3355 12765
rect 2330 12730 2335 12760
rect 2365 12730 3355 12760
rect 2330 12720 3355 12730
rect 2330 12690 2335 12720
rect 2365 12690 3355 12720
rect 2330 12685 3355 12690
rect 2330 12600 3800 12605
rect 2330 12570 2335 12600
rect 2365 12570 3800 12600
rect 2330 12560 3800 12570
rect 2330 12530 2335 12560
rect 2365 12530 3800 12560
rect 2330 12520 3800 12530
rect 2330 12490 2335 12520
rect 2365 12490 3800 12520
rect 2330 12485 3800 12490
rect 5670 12200 6630 12205
rect 5670 12170 6595 12200
rect 6625 12170 6630 12200
rect 5670 12160 6630 12170
rect 5670 12130 6595 12160
rect 6625 12130 6630 12160
rect 5670 12120 6630 12130
rect 5670 12090 6595 12120
rect 6625 12090 6630 12120
rect 5670 12085 6630 12090
rect 5870 11485 6340 11490
rect 5870 11455 6305 11485
rect 6335 11455 6340 11485
rect 5870 11445 6340 11455
rect 5870 11415 6305 11445
rect 6335 11415 6340 11445
rect 5870 11405 6340 11415
rect 5870 11375 6305 11405
rect 6335 11375 6340 11405
rect 5870 11370 6340 11375
rect 2055 10085 3030 10090
rect 2055 10055 2060 10085
rect 2090 10055 2995 10085
rect 3025 10055 3030 10085
rect 2055 10050 3030 10055
rect -90 9635 -30 9650
rect -90 9605 -75 9635
rect -45 9605 -30 9635
rect -90 9570 -30 9605
rect -90 9540 -75 9570
rect -45 9540 -30 9570
rect -90 9500 -30 9540
rect -90 9470 -75 9500
rect -45 9470 -30 9500
rect -90 9430 -30 9470
rect -90 9400 -75 9430
rect -45 9400 -30 9430
rect -90 9360 -30 9400
rect -90 9330 -75 9360
rect -45 9330 -30 9360
rect -90 9295 -30 9330
rect -90 9265 -75 9295
rect -45 9265 -30 9295
rect -90 9235 -30 9265
rect -90 9205 -75 9235
rect -45 9205 -30 9235
rect -90 9170 -30 9205
rect -90 9140 -75 9170
rect -45 9140 -30 9170
rect -90 9100 -30 9140
rect -90 9070 -75 9100
rect -45 9070 -30 9100
rect -90 9030 -30 9070
rect -90 9000 -75 9030
rect -45 9000 -30 9030
rect -90 8960 -30 9000
rect -90 8930 -75 8960
rect -45 8930 -30 8960
rect -90 8895 -30 8930
rect -90 8865 -75 8895
rect -45 8865 -30 8895
rect -90 8835 -30 8865
rect -90 8805 -75 8835
rect -45 8805 -30 8835
rect -90 8770 -30 8805
rect -90 8740 -75 8770
rect -45 8740 -30 8770
rect -90 8700 -30 8740
rect -90 8670 -75 8700
rect -45 8670 -30 8700
rect -90 8630 -30 8670
rect -90 8600 -75 8630
rect -45 8600 -30 8630
rect -90 8560 -30 8600
rect -90 8530 -75 8560
rect -45 8530 -30 8560
rect -90 8495 -30 8530
rect -90 8465 -75 8495
rect -45 8465 -30 8495
rect -90 8435 -30 8465
rect -90 8405 -75 8435
rect -45 8405 -30 8435
rect -90 8370 -30 8405
rect -90 8340 -75 8370
rect -45 8340 -30 8370
rect -90 8300 -30 8340
rect -90 8270 -75 8300
rect -45 8270 -30 8300
rect -90 8230 -30 8270
rect -90 8200 -75 8230
rect -45 8200 -30 8230
rect -90 8160 -30 8200
rect -90 8130 -75 8160
rect -45 8130 -30 8160
rect -90 8095 -30 8130
rect -90 8065 -75 8095
rect -45 8065 -30 8095
rect -90 8035 -30 8065
rect -90 8005 -75 8035
rect -45 8005 -30 8035
rect -90 7970 -30 8005
rect -90 7940 -75 7970
rect -45 7940 -30 7970
rect -90 7900 -30 7940
rect -90 7870 -75 7900
rect -45 7870 -30 7900
rect -90 7830 -30 7870
rect -90 7800 -75 7830
rect -45 7800 -30 7830
rect -90 7760 -30 7800
rect -90 7730 -75 7760
rect -45 7730 -30 7760
rect -90 7695 -30 7730
rect -90 7665 -75 7695
rect -45 7665 -30 7695
rect -90 7635 -30 7665
rect -90 7605 -75 7635
rect -45 7605 -30 7635
rect -90 7570 -30 7605
rect -90 7540 -75 7570
rect -45 7540 -30 7570
rect -90 7500 -30 7540
rect -90 7470 -75 7500
rect -45 7470 -30 7500
rect -90 7430 -30 7470
rect -90 7400 -75 7430
rect -45 7400 -30 7430
rect -90 7360 -30 7400
rect -90 7330 -75 7360
rect -45 7330 -30 7360
rect -90 7295 -30 7330
rect -90 7265 -75 7295
rect -45 7265 -30 7295
rect -90 7235 -30 7265
rect -90 7205 -75 7235
rect -45 7205 -30 7235
rect -90 7170 -30 7205
rect -90 7140 -75 7170
rect -45 7140 -30 7170
rect -90 7100 -30 7140
rect -90 7070 -75 7100
rect -45 7070 -30 7100
rect -90 7030 -30 7070
rect -90 7000 -75 7030
rect -45 7000 -30 7030
rect -90 6960 -30 7000
rect -90 6930 -75 6960
rect -45 6930 -30 6960
rect -90 6895 -30 6930
rect -90 6865 -75 6895
rect -45 6865 -30 6895
rect -90 6835 -30 6865
rect -90 6805 -75 6835
rect -45 6805 -30 6835
rect -90 6770 -30 6805
rect -90 6740 -75 6770
rect -45 6740 -30 6770
rect -90 6700 -30 6740
rect -90 6670 -75 6700
rect -45 6670 -30 6700
rect -90 6630 -30 6670
rect -90 6600 -75 6630
rect -45 6600 -30 6630
rect -90 6560 -30 6600
rect -90 6530 -75 6560
rect -45 6530 -30 6560
rect -90 6495 -30 6530
rect -90 6465 -75 6495
rect -45 6465 -30 6495
rect -90 6450 -30 6465
rect 260 9635 320 9650
rect 260 9605 275 9635
rect 305 9605 320 9635
rect 260 9570 320 9605
rect 260 9540 275 9570
rect 305 9540 320 9570
rect 260 9500 320 9540
rect 260 9470 275 9500
rect 305 9470 320 9500
rect 260 9430 320 9470
rect 260 9400 275 9430
rect 305 9400 320 9430
rect 260 9360 320 9400
rect 260 9330 275 9360
rect 305 9330 320 9360
rect 260 9295 320 9330
rect 260 9265 275 9295
rect 305 9265 320 9295
rect 260 9235 320 9265
rect 260 9205 275 9235
rect 305 9205 320 9235
rect 260 9170 320 9205
rect 260 9140 275 9170
rect 305 9140 320 9170
rect 260 9100 320 9140
rect 260 9070 275 9100
rect 305 9070 320 9100
rect 260 9030 320 9070
rect 260 9000 275 9030
rect 305 9000 320 9030
rect 260 8960 320 9000
rect 260 8930 275 8960
rect 305 8930 320 8960
rect 260 8895 320 8930
rect 260 8865 275 8895
rect 305 8865 320 8895
rect 260 8835 320 8865
rect 260 8805 275 8835
rect 305 8805 320 8835
rect 260 8770 320 8805
rect 260 8740 275 8770
rect 305 8740 320 8770
rect 260 8700 320 8740
rect 260 8670 275 8700
rect 305 8670 320 8700
rect 260 8630 320 8670
rect 260 8600 275 8630
rect 305 8600 320 8630
rect 260 8560 320 8600
rect 260 8530 275 8560
rect 305 8530 320 8560
rect 260 8495 320 8530
rect 260 8465 275 8495
rect 305 8465 320 8495
rect 260 8435 320 8465
rect 260 8405 275 8435
rect 305 8405 320 8435
rect 260 8370 320 8405
rect 260 8340 275 8370
rect 305 8340 320 8370
rect 260 8300 320 8340
rect 260 8270 275 8300
rect 305 8270 320 8300
rect 260 8230 320 8270
rect 260 8200 275 8230
rect 305 8200 320 8230
rect 260 8160 320 8200
rect 260 8130 275 8160
rect 305 8130 320 8160
rect 260 8095 320 8130
rect 260 8065 275 8095
rect 305 8065 320 8095
rect 260 8035 320 8065
rect 260 8005 275 8035
rect 305 8005 320 8035
rect 260 7970 320 8005
rect 260 7940 275 7970
rect 305 7940 320 7970
rect 260 7900 320 7940
rect 260 7870 275 7900
rect 305 7870 320 7900
rect 260 7830 320 7870
rect 260 7800 275 7830
rect 305 7800 320 7830
rect 260 7760 320 7800
rect 260 7730 275 7760
rect 305 7730 320 7760
rect 260 7695 320 7730
rect 260 7665 275 7695
rect 305 7665 320 7695
rect 260 7635 320 7665
rect 260 7605 275 7635
rect 305 7605 320 7635
rect 260 7570 320 7605
rect 260 7540 275 7570
rect 305 7540 320 7570
rect 260 7500 320 7540
rect 260 7470 275 7500
rect 305 7470 320 7500
rect 260 7430 320 7470
rect 260 7400 275 7430
rect 305 7400 320 7430
rect 260 7360 320 7400
rect 260 7330 275 7360
rect 305 7330 320 7360
rect 260 7295 320 7330
rect 260 7265 275 7295
rect 305 7265 320 7295
rect 260 7235 320 7265
rect 260 7205 275 7235
rect 305 7205 320 7235
rect 260 7170 320 7205
rect 260 7140 275 7170
rect 305 7140 320 7170
rect 260 7100 320 7140
rect 260 7070 275 7100
rect 305 7070 320 7100
rect 260 7030 320 7070
rect 260 7000 275 7030
rect 305 7000 320 7030
rect 260 6960 320 7000
rect 260 6930 275 6960
rect 305 6930 320 6960
rect 260 6895 320 6930
rect 260 6865 275 6895
rect 305 6865 320 6895
rect 260 6835 320 6865
rect 260 6805 275 6835
rect 305 6805 320 6835
rect 260 6770 320 6805
rect 260 6740 275 6770
rect 305 6740 320 6770
rect 260 6700 320 6740
rect 260 6670 275 6700
rect 305 6670 320 6700
rect 260 6630 320 6670
rect 260 6600 275 6630
rect 305 6600 320 6630
rect 260 6560 320 6600
rect 260 6530 275 6560
rect 305 6530 320 6560
rect 260 6495 320 6530
rect 260 6465 275 6495
rect 305 6465 320 6495
rect 260 6450 320 6465
rect 610 9635 670 9650
rect 610 9605 625 9635
rect 655 9605 670 9635
rect 610 9570 670 9605
rect 610 9540 625 9570
rect 655 9540 670 9570
rect 610 9500 670 9540
rect 610 9470 625 9500
rect 655 9470 670 9500
rect 610 9430 670 9470
rect 610 9400 625 9430
rect 655 9400 670 9430
rect 610 9360 670 9400
rect 610 9330 625 9360
rect 655 9330 670 9360
rect 610 9295 670 9330
rect 610 9265 625 9295
rect 655 9265 670 9295
rect 610 9235 670 9265
rect 610 9205 625 9235
rect 655 9205 670 9235
rect 610 9170 670 9205
rect 610 9140 625 9170
rect 655 9140 670 9170
rect 610 9100 670 9140
rect 610 9070 625 9100
rect 655 9070 670 9100
rect 610 9030 670 9070
rect 610 9000 625 9030
rect 655 9000 670 9030
rect 610 8960 670 9000
rect 610 8930 625 8960
rect 655 8930 670 8960
rect 610 8895 670 8930
rect 610 8865 625 8895
rect 655 8865 670 8895
rect 610 8835 670 8865
rect 610 8805 625 8835
rect 655 8805 670 8835
rect 610 8770 670 8805
rect 610 8740 625 8770
rect 655 8740 670 8770
rect 610 8700 670 8740
rect 610 8670 625 8700
rect 655 8670 670 8700
rect 610 8630 670 8670
rect 610 8600 625 8630
rect 655 8600 670 8630
rect 610 8560 670 8600
rect 610 8530 625 8560
rect 655 8530 670 8560
rect 610 8495 670 8530
rect 610 8465 625 8495
rect 655 8465 670 8495
rect 610 8435 670 8465
rect 610 8405 625 8435
rect 655 8405 670 8435
rect 610 8370 670 8405
rect 610 8340 625 8370
rect 655 8340 670 8370
rect 610 8300 670 8340
rect 610 8270 625 8300
rect 655 8270 670 8300
rect 610 8230 670 8270
rect 610 8200 625 8230
rect 655 8200 670 8230
rect 610 8160 670 8200
rect 610 8130 625 8160
rect 655 8130 670 8160
rect 610 8095 670 8130
rect 610 8065 625 8095
rect 655 8065 670 8095
rect 610 8035 670 8065
rect 610 8005 625 8035
rect 655 8005 670 8035
rect 610 7970 670 8005
rect 610 7940 625 7970
rect 655 7940 670 7970
rect 610 7900 670 7940
rect 610 7870 625 7900
rect 655 7870 670 7900
rect 610 7830 670 7870
rect 610 7800 625 7830
rect 655 7800 670 7830
rect 610 7760 670 7800
rect 610 7730 625 7760
rect 655 7730 670 7760
rect 610 7695 670 7730
rect 610 7665 625 7695
rect 655 7665 670 7695
rect 610 7635 670 7665
rect 610 7605 625 7635
rect 655 7605 670 7635
rect 610 7570 670 7605
rect 610 7540 625 7570
rect 655 7540 670 7570
rect 610 7500 670 7540
rect 610 7470 625 7500
rect 655 7470 670 7500
rect 610 7430 670 7470
rect 610 7400 625 7430
rect 655 7400 670 7430
rect 610 7360 670 7400
rect 610 7330 625 7360
rect 655 7330 670 7360
rect 610 7295 670 7330
rect 610 7265 625 7295
rect 655 7265 670 7295
rect 610 7235 670 7265
rect 610 7205 625 7235
rect 655 7205 670 7235
rect 610 7170 670 7205
rect 610 7140 625 7170
rect 655 7140 670 7170
rect 610 7100 670 7140
rect 610 7070 625 7100
rect 655 7070 670 7100
rect 610 7030 670 7070
rect 610 7000 625 7030
rect 655 7000 670 7030
rect 610 6960 670 7000
rect 610 6930 625 6960
rect 655 6930 670 6960
rect 610 6895 670 6930
rect 610 6865 625 6895
rect 655 6865 670 6895
rect 610 6835 670 6865
rect 610 6805 625 6835
rect 655 6805 670 6835
rect 610 6770 670 6805
rect 610 6740 625 6770
rect 655 6740 670 6770
rect 610 6700 670 6740
rect 610 6670 625 6700
rect 655 6670 670 6700
rect 610 6630 670 6670
rect 610 6600 625 6630
rect 655 6600 670 6630
rect 610 6560 670 6600
rect 610 6530 625 6560
rect 655 6530 670 6560
rect 610 6495 670 6530
rect 610 6465 625 6495
rect 655 6465 670 6495
rect 610 6450 670 6465
rect 1310 9635 1370 9650
rect 1310 9605 1325 9635
rect 1355 9605 1370 9635
rect 1310 9570 1370 9605
rect 1310 9540 1325 9570
rect 1355 9540 1370 9570
rect 1310 9500 1370 9540
rect 1310 9470 1325 9500
rect 1355 9470 1370 9500
rect 1310 9430 1370 9470
rect 1310 9400 1325 9430
rect 1355 9400 1370 9430
rect 1310 9360 1370 9400
rect 1310 9330 1325 9360
rect 1355 9330 1370 9360
rect 1310 9295 1370 9330
rect 1310 9265 1325 9295
rect 1355 9265 1370 9295
rect 1310 9235 1370 9265
rect 1310 9205 1325 9235
rect 1355 9205 1370 9235
rect 1310 9170 1370 9205
rect 1310 9140 1325 9170
rect 1355 9140 1370 9170
rect 1310 9100 1370 9140
rect 1310 9070 1325 9100
rect 1355 9070 1370 9100
rect 1310 9030 1370 9070
rect 1310 9000 1325 9030
rect 1355 9000 1370 9030
rect 1310 8960 1370 9000
rect 1310 8930 1325 8960
rect 1355 8930 1370 8960
rect 1310 8895 1370 8930
rect 1310 8865 1325 8895
rect 1355 8865 1370 8895
rect 1310 8835 1370 8865
rect 1310 8805 1325 8835
rect 1355 8805 1370 8835
rect 1310 8770 1370 8805
rect 1310 8740 1325 8770
rect 1355 8740 1370 8770
rect 1310 8700 1370 8740
rect 1310 8670 1325 8700
rect 1355 8670 1370 8700
rect 1310 8630 1370 8670
rect 1310 8600 1325 8630
rect 1355 8600 1370 8630
rect 1310 8560 1370 8600
rect 1310 8530 1325 8560
rect 1355 8530 1370 8560
rect 1310 8495 1370 8530
rect 1310 8465 1325 8495
rect 1355 8465 1370 8495
rect 1310 8435 1370 8465
rect 1310 8405 1325 8435
rect 1355 8405 1370 8435
rect 1310 8370 1370 8405
rect 1310 8340 1325 8370
rect 1355 8340 1370 8370
rect 1310 8300 1370 8340
rect 1310 8270 1325 8300
rect 1355 8270 1370 8300
rect 1310 8230 1370 8270
rect 1310 8200 1325 8230
rect 1355 8200 1370 8230
rect 1310 8160 1370 8200
rect 1310 8130 1325 8160
rect 1355 8130 1370 8160
rect 1310 8095 1370 8130
rect 1310 8065 1325 8095
rect 1355 8065 1370 8095
rect 1310 8035 1370 8065
rect 1310 8005 1325 8035
rect 1355 8005 1370 8035
rect 1310 7970 1370 8005
rect 1310 7940 1325 7970
rect 1355 7940 1370 7970
rect 1310 7900 1370 7940
rect 1310 7870 1325 7900
rect 1355 7870 1370 7900
rect 1310 7830 1370 7870
rect 1310 7800 1325 7830
rect 1355 7800 1370 7830
rect 1310 7760 1370 7800
rect 1310 7730 1325 7760
rect 1355 7730 1370 7760
rect 1310 7695 1370 7730
rect 1310 7665 1325 7695
rect 1355 7665 1370 7695
rect 1310 7635 1370 7665
rect 1310 7605 1325 7635
rect 1355 7605 1370 7635
rect 1310 7570 1370 7605
rect 1310 7540 1325 7570
rect 1355 7540 1370 7570
rect 1310 7500 1370 7540
rect 1310 7470 1325 7500
rect 1355 7470 1370 7500
rect 1310 7430 1370 7470
rect 1310 7400 1325 7430
rect 1355 7400 1370 7430
rect 1310 7360 1370 7400
rect 1310 7330 1325 7360
rect 1355 7330 1370 7360
rect 1310 7295 1370 7330
rect 1310 7265 1325 7295
rect 1355 7265 1370 7295
rect 1310 7235 1370 7265
rect 1310 7205 1325 7235
rect 1355 7205 1370 7235
rect 1310 7170 1370 7205
rect 1310 7140 1325 7170
rect 1355 7140 1370 7170
rect 1310 7100 1370 7140
rect 1310 7070 1325 7100
rect 1355 7070 1370 7100
rect 1310 7030 1370 7070
rect 1310 7000 1325 7030
rect 1355 7000 1370 7030
rect 1310 6960 1370 7000
rect 1310 6930 1325 6960
rect 1355 6930 1370 6960
rect 1310 6895 1370 6930
rect 1310 6865 1325 6895
rect 1355 6865 1370 6895
rect 1310 6835 1370 6865
rect 1310 6805 1325 6835
rect 1355 6805 1370 6835
rect 1310 6770 1370 6805
rect 1310 6740 1325 6770
rect 1355 6740 1370 6770
rect 1310 6700 1370 6740
rect 1310 6670 1325 6700
rect 1355 6670 1370 6700
rect 1310 6630 1370 6670
rect 1310 6600 1325 6630
rect 1355 6600 1370 6630
rect 1310 6560 1370 6600
rect 1310 6530 1325 6560
rect 1355 6530 1370 6560
rect 1310 6495 1370 6530
rect 1310 6465 1325 6495
rect 1355 6465 1370 6495
rect 1310 6450 1370 6465
rect 1660 9635 1720 9650
rect 1660 9605 1675 9635
rect 1705 9605 1720 9635
rect 1660 9570 1720 9605
rect 1660 9540 1675 9570
rect 1705 9540 1720 9570
rect 1660 9500 1720 9540
rect 1660 9470 1675 9500
rect 1705 9470 1720 9500
rect 1660 9430 1720 9470
rect 1660 9400 1675 9430
rect 1705 9400 1720 9430
rect 1660 9360 1720 9400
rect 1660 9330 1675 9360
rect 1705 9330 1720 9360
rect 1660 9295 1720 9330
rect 1660 9265 1675 9295
rect 1705 9265 1720 9295
rect 1660 9235 1720 9265
rect 1660 9205 1675 9235
rect 1705 9205 1720 9235
rect 1660 9170 1720 9205
rect 1660 9140 1675 9170
rect 1705 9140 1720 9170
rect 1660 9100 1720 9140
rect 1660 9070 1675 9100
rect 1705 9070 1720 9100
rect 1660 9030 1720 9070
rect 1660 9000 1675 9030
rect 1705 9000 1720 9030
rect 1660 8960 1720 9000
rect 1660 8930 1675 8960
rect 1705 8930 1720 8960
rect 1660 8895 1720 8930
rect 1660 8865 1675 8895
rect 1705 8865 1720 8895
rect 1660 8835 1720 8865
rect 1660 8805 1675 8835
rect 1705 8805 1720 8835
rect 1660 8770 1720 8805
rect 1660 8740 1675 8770
rect 1705 8740 1720 8770
rect 1660 8700 1720 8740
rect 1660 8670 1675 8700
rect 1705 8670 1720 8700
rect 1660 8630 1720 8670
rect 1660 8600 1675 8630
rect 1705 8600 1720 8630
rect 1660 8560 1720 8600
rect 1660 8530 1675 8560
rect 1705 8530 1720 8560
rect 1660 8495 1720 8530
rect 1660 8465 1675 8495
rect 1705 8465 1720 8495
rect 1660 8435 1720 8465
rect 1660 8405 1675 8435
rect 1705 8405 1720 8435
rect 1660 8370 1720 8405
rect 1660 8340 1675 8370
rect 1705 8340 1720 8370
rect 1660 8300 1720 8340
rect 1660 8270 1675 8300
rect 1705 8270 1720 8300
rect 1660 8230 1720 8270
rect 1660 8200 1675 8230
rect 1705 8200 1720 8230
rect 1660 8160 1720 8200
rect 1660 8130 1675 8160
rect 1705 8130 1720 8160
rect 1660 8095 1720 8130
rect 1660 8065 1675 8095
rect 1705 8065 1720 8095
rect 1660 8035 1720 8065
rect 1660 8005 1675 8035
rect 1705 8005 1720 8035
rect 1660 7970 1720 8005
rect 1660 7940 1675 7970
rect 1705 7940 1720 7970
rect 1660 7900 1720 7940
rect 1660 7870 1675 7900
rect 1705 7870 1720 7900
rect 1660 7830 1720 7870
rect 1660 7800 1675 7830
rect 1705 7800 1720 7830
rect 1660 7760 1720 7800
rect 1660 7730 1675 7760
rect 1705 7730 1720 7760
rect 1660 7695 1720 7730
rect 1660 7665 1675 7695
rect 1705 7665 1720 7695
rect 1660 7635 1720 7665
rect 1660 7605 1675 7635
rect 1705 7605 1720 7635
rect 1660 7570 1720 7605
rect 1660 7540 1675 7570
rect 1705 7540 1720 7570
rect 1660 7500 1720 7540
rect 1660 7470 1675 7500
rect 1705 7470 1720 7500
rect 1660 7430 1720 7470
rect 1660 7400 1675 7430
rect 1705 7400 1720 7430
rect 1660 7360 1720 7400
rect 1660 7330 1675 7360
rect 1705 7330 1720 7360
rect 1660 7295 1720 7330
rect 1660 7265 1675 7295
rect 1705 7265 1720 7295
rect 1660 7235 1720 7265
rect 1660 7205 1675 7235
rect 1705 7205 1720 7235
rect 1660 7170 1720 7205
rect 1660 7140 1675 7170
rect 1705 7140 1720 7170
rect 1660 7100 1720 7140
rect 1660 7070 1675 7100
rect 1705 7070 1720 7100
rect 1660 7030 1720 7070
rect 1660 7000 1675 7030
rect 1705 7000 1720 7030
rect 1660 6960 1720 7000
rect 1660 6930 1675 6960
rect 1705 6930 1720 6960
rect 1660 6895 1720 6930
rect 1660 6865 1675 6895
rect 1705 6865 1720 6895
rect 1660 6835 1720 6865
rect 1660 6805 1675 6835
rect 1705 6805 1720 6835
rect 1660 6770 1720 6805
rect 1660 6740 1675 6770
rect 1705 6740 1720 6770
rect 1660 6700 1720 6740
rect 1660 6670 1675 6700
rect 1705 6670 1720 6700
rect 1660 6630 1720 6670
rect 1660 6600 1675 6630
rect 1705 6600 1720 6630
rect 1660 6560 1720 6600
rect 1660 6530 1675 6560
rect 1705 6530 1720 6560
rect 1660 6495 1720 6530
rect 1660 6465 1675 6495
rect 1705 6465 1720 6495
rect 1660 6450 1720 6465
rect 2375 9635 2435 9650
rect 2375 9605 2390 9635
rect 2420 9605 2435 9635
rect 2375 9570 2435 9605
rect 2375 9540 2390 9570
rect 2420 9540 2435 9570
rect 2375 9500 2435 9540
rect 2375 9470 2390 9500
rect 2420 9470 2435 9500
rect 2375 9430 2435 9470
rect 2375 9400 2390 9430
rect 2420 9400 2435 9430
rect 2375 9360 2435 9400
rect 2375 9330 2390 9360
rect 2420 9330 2435 9360
rect 2375 9295 2435 9330
rect 2375 9265 2390 9295
rect 2420 9265 2435 9295
rect 2375 9235 2435 9265
rect 2375 9205 2390 9235
rect 2420 9205 2435 9235
rect 2375 9170 2435 9205
rect 2375 9140 2390 9170
rect 2420 9140 2435 9170
rect 2375 9100 2435 9140
rect 2375 9070 2390 9100
rect 2420 9070 2435 9100
rect 2375 9030 2435 9070
rect 2375 9000 2390 9030
rect 2420 9000 2435 9030
rect 2375 8960 2435 9000
rect 2375 8930 2390 8960
rect 2420 8930 2435 8960
rect 2375 8895 2435 8930
rect 2375 8865 2390 8895
rect 2420 8865 2435 8895
rect 2375 8835 2435 8865
rect 2375 8805 2390 8835
rect 2420 8805 2435 8835
rect 2375 8770 2435 8805
rect 2375 8740 2390 8770
rect 2420 8740 2435 8770
rect 2375 8700 2435 8740
rect 2375 8670 2390 8700
rect 2420 8670 2435 8700
rect 2375 8630 2435 8670
rect 2375 8600 2390 8630
rect 2420 8600 2435 8630
rect 2375 8560 2435 8600
rect 2375 8530 2390 8560
rect 2420 8530 2435 8560
rect 2375 8495 2435 8530
rect 2375 8465 2390 8495
rect 2420 8465 2435 8495
rect 2375 8435 2435 8465
rect 2375 8405 2390 8435
rect 2420 8405 2435 8435
rect 2375 8370 2435 8405
rect 2375 8340 2390 8370
rect 2420 8340 2435 8370
rect 2375 8300 2435 8340
rect 2375 8270 2390 8300
rect 2420 8270 2435 8300
rect 2375 8230 2435 8270
rect 2375 8200 2390 8230
rect 2420 8200 2435 8230
rect 2375 8160 2435 8200
rect 2375 8130 2390 8160
rect 2420 8130 2435 8160
rect 2375 8095 2435 8130
rect 2375 8065 2390 8095
rect 2420 8065 2435 8095
rect 2375 8035 2435 8065
rect 2375 8005 2390 8035
rect 2420 8005 2435 8035
rect 2375 7970 2435 8005
rect 2375 7940 2390 7970
rect 2420 7940 2435 7970
rect 2375 7900 2435 7940
rect 2375 7870 2390 7900
rect 2420 7870 2435 7900
rect 2375 7830 2435 7870
rect 2375 7800 2390 7830
rect 2420 7800 2435 7830
rect 2375 7760 2435 7800
rect 2375 7730 2390 7760
rect 2420 7730 2435 7760
rect 2375 7695 2435 7730
rect 2375 7665 2390 7695
rect 2420 7665 2435 7695
rect 2375 7635 2435 7665
rect 2375 7605 2390 7635
rect 2420 7605 2435 7635
rect 2375 7570 2435 7605
rect 2375 7540 2390 7570
rect 2420 7540 2435 7570
rect 2375 7500 2435 7540
rect 2375 7470 2390 7500
rect 2420 7470 2435 7500
rect 2375 7430 2435 7470
rect 2375 7400 2390 7430
rect 2420 7400 2435 7430
rect 2375 7360 2435 7400
rect 2375 7330 2390 7360
rect 2420 7330 2435 7360
rect 2375 7295 2435 7330
rect 2375 7265 2390 7295
rect 2420 7265 2435 7295
rect 2375 7235 2435 7265
rect 2375 7205 2390 7235
rect 2420 7205 2435 7235
rect 2375 7170 2435 7205
rect 2375 7140 2390 7170
rect 2420 7140 2435 7170
rect 2375 7100 2435 7140
rect 2375 7070 2390 7100
rect 2420 7070 2435 7100
rect 2375 7030 2435 7070
rect 2375 7000 2390 7030
rect 2420 7000 2435 7030
rect 2375 6960 2435 7000
rect 2375 6930 2390 6960
rect 2420 6930 2435 6960
rect 2375 6895 2435 6930
rect 2375 6865 2390 6895
rect 2420 6865 2435 6895
rect 2375 6835 2435 6865
rect 2375 6805 2390 6835
rect 2420 6805 2435 6835
rect 2375 6770 2435 6805
rect 2375 6740 2390 6770
rect 2420 6740 2435 6770
rect 2375 6700 2435 6740
rect 2375 6670 2390 6700
rect 2420 6670 2435 6700
rect 2375 6630 2435 6670
rect 2375 6600 2390 6630
rect 2420 6600 2435 6630
rect 2375 6560 2435 6600
rect 2375 6530 2390 6560
rect 2420 6530 2435 6560
rect 2375 6495 2435 6530
rect 2375 6465 2390 6495
rect 2420 6465 2435 6495
rect 2375 6450 2435 6465
rect 3225 9635 3285 9650
rect 3225 9605 3240 9635
rect 3270 9605 3285 9635
rect 3225 9570 3285 9605
rect 3225 9540 3240 9570
rect 3270 9540 3285 9570
rect 3225 9500 3285 9540
rect 3225 9470 3240 9500
rect 3270 9470 3285 9500
rect 3225 9430 3285 9470
rect 3225 9400 3240 9430
rect 3270 9400 3285 9430
rect 3225 9360 3285 9400
rect 3225 9330 3240 9360
rect 3270 9330 3285 9360
rect 3225 9295 3285 9330
rect 3225 9265 3240 9295
rect 3270 9265 3285 9295
rect 3225 9235 3285 9265
rect 3225 9205 3240 9235
rect 3270 9205 3285 9235
rect 3225 9170 3285 9205
rect 3225 9140 3240 9170
rect 3270 9140 3285 9170
rect 3225 9100 3285 9140
rect 3225 9070 3240 9100
rect 3270 9070 3285 9100
rect 3225 9030 3285 9070
rect 3225 9000 3240 9030
rect 3270 9000 3285 9030
rect 3225 8960 3285 9000
rect 3225 8930 3240 8960
rect 3270 8930 3285 8960
rect 3225 8895 3285 8930
rect 3225 8865 3240 8895
rect 3270 8865 3285 8895
rect 3225 8835 3285 8865
rect 3225 8805 3240 8835
rect 3270 8805 3285 8835
rect 3225 8770 3285 8805
rect 3225 8740 3240 8770
rect 3270 8740 3285 8770
rect 3225 8700 3285 8740
rect 3225 8670 3240 8700
rect 3270 8670 3285 8700
rect 3225 8630 3285 8670
rect 3225 8600 3240 8630
rect 3270 8600 3285 8630
rect 3225 8560 3285 8600
rect 3225 8530 3240 8560
rect 3270 8530 3285 8560
rect 3225 8495 3285 8530
rect 3225 8465 3240 8495
rect 3270 8465 3285 8495
rect 3225 8435 3285 8465
rect 3225 8405 3240 8435
rect 3270 8405 3285 8435
rect 3225 8370 3285 8405
rect 3225 8340 3240 8370
rect 3270 8340 3285 8370
rect 3225 8300 3285 8340
rect 3225 8270 3240 8300
rect 3270 8270 3285 8300
rect 3225 8230 3285 8270
rect 3225 8200 3240 8230
rect 3270 8200 3285 8230
rect 3225 8160 3285 8200
rect 3225 8130 3240 8160
rect 3270 8130 3285 8160
rect 3225 8095 3285 8130
rect 3225 8065 3240 8095
rect 3270 8065 3285 8095
rect 3225 8035 3285 8065
rect 3225 8005 3240 8035
rect 3270 8005 3285 8035
rect 3225 7970 3285 8005
rect 3225 7940 3240 7970
rect 3270 7940 3285 7970
rect 3225 7900 3285 7940
rect 3225 7870 3240 7900
rect 3270 7870 3285 7900
rect 3225 7830 3285 7870
rect 3225 7800 3240 7830
rect 3270 7800 3285 7830
rect 3225 7760 3285 7800
rect 3225 7730 3240 7760
rect 3270 7730 3285 7760
rect 3225 7695 3285 7730
rect 3225 7665 3240 7695
rect 3270 7665 3285 7695
rect 3225 7635 3285 7665
rect 3225 7605 3240 7635
rect 3270 7605 3285 7635
rect 3225 7570 3285 7605
rect 3225 7540 3240 7570
rect 3270 7540 3285 7570
rect 3225 7500 3285 7540
rect 3225 7470 3240 7500
rect 3270 7470 3285 7500
rect 3225 7430 3285 7470
rect 3225 7400 3240 7430
rect 3270 7400 3285 7430
rect 3225 7360 3285 7400
rect 3225 7330 3240 7360
rect 3270 7330 3285 7360
rect 3225 7295 3285 7330
rect 3225 7265 3240 7295
rect 3270 7265 3285 7295
rect 3225 7235 3285 7265
rect 3225 7205 3240 7235
rect 3270 7205 3285 7235
rect 3225 7170 3285 7205
rect 3225 7140 3240 7170
rect 3270 7140 3285 7170
rect 3225 7100 3285 7140
rect 3225 7070 3240 7100
rect 3270 7070 3285 7100
rect 3225 7030 3285 7070
rect 3225 7000 3240 7030
rect 3270 7000 3285 7030
rect 3225 6960 3285 7000
rect 3225 6930 3240 6960
rect 3270 6930 3285 6960
rect 3225 6895 3285 6930
rect 3225 6865 3240 6895
rect 3270 6865 3285 6895
rect 3225 6835 3285 6865
rect 3225 6805 3240 6835
rect 3270 6805 3285 6835
rect 3225 6770 3285 6805
rect 3225 6740 3240 6770
rect 3270 6740 3285 6770
rect 3225 6700 3285 6740
rect 3225 6670 3240 6700
rect 3270 6670 3285 6700
rect 3225 6630 3285 6670
rect 3225 6600 3240 6630
rect 3270 6600 3285 6630
rect 3225 6560 3285 6600
rect 3225 6530 3240 6560
rect 3270 6530 3285 6560
rect 3225 6495 3285 6530
rect 3225 6465 3240 6495
rect 3270 6465 3285 6495
rect 3225 6450 3285 6465
rect 5635 9635 5695 9650
rect 5635 9605 5650 9635
rect 5680 9605 5695 9635
rect 5635 9570 5695 9605
rect 5635 9540 5650 9570
rect 5680 9540 5695 9570
rect 5635 9500 5695 9540
rect 5635 9470 5650 9500
rect 5680 9470 5695 9500
rect 5635 9430 5695 9470
rect 5635 9400 5650 9430
rect 5680 9400 5695 9430
rect 5635 9360 5695 9400
rect 5635 9330 5650 9360
rect 5680 9330 5695 9360
rect 5635 9295 5695 9330
rect 5635 9265 5650 9295
rect 5680 9265 5695 9295
rect 5635 9235 5695 9265
rect 5635 9205 5650 9235
rect 5680 9205 5695 9235
rect 5635 9170 5695 9205
rect 5635 9140 5650 9170
rect 5680 9140 5695 9170
rect 5635 9100 5695 9140
rect 5635 9070 5650 9100
rect 5680 9070 5695 9100
rect 5635 9030 5695 9070
rect 5635 9000 5650 9030
rect 5680 9000 5695 9030
rect 5635 8960 5695 9000
rect 5635 8930 5650 8960
rect 5680 8930 5695 8960
rect 5635 8895 5695 8930
rect 5635 8865 5650 8895
rect 5680 8865 5695 8895
rect 5635 8835 5695 8865
rect 5635 8805 5650 8835
rect 5680 8805 5695 8835
rect 5635 8770 5695 8805
rect 5635 8740 5650 8770
rect 5680 8740 5695 8770
rect 5635 8700 5695 8740
rect 5635 8670 5650 8700
rect 5680 8670 5695 8700
rect 5635 8630 5695 8670
rect 5635 8600 5650 8630
rect 5680 8600 5695 8630
rect 5635 8560 5695 8600
rect 5635 8530 5650 8560
rect 5680 8530 5695 8560
rect 5635 8495 5695 8530
rect 5635 8465 5650 8495
rect 5680 8465 5695 8495
rect 5635 8435 5695 8465
rect 5635 8405 5650 8435
rect 5680 8405 5695 8435
rect 5635 8370 5695 8405
rect 5635 8340 5650 8370
rect 5680 8340 5695 8370
rect 5635 8300 5695 8340
rect 5635 8270 5650 8300
rect 5680 8270 5695 8300
rect 5635 8230 5695 8270
rect 5635 8200 5650 8230
rect 5680 8200 5695 8230
rect 5635 8160 5695 8200
rect 5635 8130 5650 8160
rect 5680 8130 5695 8160
rect 5635 8095 5695 8130
rect 5635 8065 5650 8095
rect 5680 8065 5695 8095
rect 5635 8035 5695 8065
rect 5635 8005 5650 8035
rect 5680 8005 5695 8035
rect 5635 7970 5695 8005
rect 5635 7940 5650 7970
rect 5680 7940 5695 7970
rect 5635 7900 5695 7940
rect 5635 7870 5650 7900
rect 5680 7870 5695 7900
rect 5635 7830 5695 7870
rect 5635 7800 5650 7830
rect 5680 7800 5695 7830
rect 5635 7760 5695 7800
rect 5635 7730 5650 7760
rect 5680 7730 5695 7760
rect 5635 7695 5695 7730
rect 5635 7665 5650 7695
rect 5680 7665 5695 7695
rect 5635 7635 5695 7665
rect 5635 7605 5650 7635
rect 5680 7605 5695 7635
rect 5635 7570 5695 7605
rect 5635 7540 5650 7570
rect 5680 7540 5695 7570
rect 5635 7500 5695 7540
rect 5635 7470 5650 7500
rect 5680 7470 5695 7500
rect 5635 7430 5695 7470
rect 5635 7400 5650 7430
rect 5680 7400 5695 7430
rect 5635 7360 5695 7400
rect 5635 7330 5650 7360
rect 5680 7330 5695 7360
rect 5635 7295 5695 7330
rect 5635 7265 5650 7295
rect 5680 7265 5695 7295
rect 5635 7235 5695 7265
rect 5635 7205 5650 7235
rect 5680 7205 5695 7235
rect 5635 7170 5695 7205
rect 5635 7140 5650 7170
rect 5680 7140 5695 7170
rect 5635 7100 5695 7140
rect 5635 7070 5650 7100
rect 5680 7070 5695 7100
rect 5635 7030 5695 7070
rect 5635 7000 5650 7030
rect 5680 7000 5695 7030
rect 5635 6960 5695 7000
rect 5635 6930 5650 6960
rect 5680 6930 5695 6960
rect 5635 6895 5695 6930
rect 5635 6865 5650 6895
rect 5680 6865 5695 6895
rect 5635 6835 5695 6865
rect 5635 6805 5650 6835
rect 5680 6805 5695 6835
rect 5635 6770 5695 6805
rect 5635 6740 5650 6770
rect 5680 6740 5695 6770
rect 5635 6700 5695 6740
rect 5635 6670 5650 6700
rect 5680 6670 5695 6700
rect 5635 6630 5695 6670
rect 5635 6600 5650 6630
rect 5680 6600 5695 6630
rect 5635 6560 5695 6600
rect 5635 6530 5650 6560
rect 5680 6530 5695 6560
rect 5635 6495 5695 6530
rect 5635 6465 5650 6495
rect 5680 6465 5695 6495
rect 5635 6450 5695 6465
rect 6290 9635 6350 9650
rect 6290 9605 6305 9635
rect 6335 9605 6350 9635
rect 6290 9570 6350 9605
rect 6290 9540 6305 9570
rect 6335 9540 6350 9570
rect 6290 9500 6350 9540
rect 6290 9470 6305 9500
rect 6335 9470 6350 9500
rect 6290 9430 6350 9470
rect 6290 9400 6305 9430
rect 6335 9400 6350 9430
rect 6290 9360 6350 9400
rect 6290 9330 6305 9360
rect 6335 9330 6350 9360
rect 6290 9295 6350 9330
rect 6290 9265 6305 9295
rect 6335 9265 6350 9295
rect 6290 9235 6350 9265
rect 6290 9205 6305 9235
rect 6335 9205 6350 9235
rect 6290 9170 6350 9205
rect 6290 9140 6305 9170
rect 6335 9140 6350 9170
rect 6290 9100 6350 9140
rect 6290 9070 6305 9100
rect 6335 9070 6350 9100
rect 6290 9030 6350 9070
rect 6290 9000 6305 9030
rect 6335 9000 6350 9030
rect 6290 8960 6350 9000
rect 6290 8930 6305 8960
rect 6335 8930 6350 8960
rect 6290 8895 6350 8930
rect 6290 8865 6305 8895
rect 6335 8865 6350 8895
rect 6290 8835 6350 8865
rect 6290 8805 6305 8835
rect 6335 8805 6350 8835
rect 6290 8770 6350 8805
rect 6290 8740 6305 8770
rect 6335 8740 6350 8770
rect 6290 8700 6350 8740
rect 6290 8670 6305 8700
rect 6335 8670 6350 8700
rect 6290 8630 6350 8670
rect 6290 8600 6305 8630
rect 6335 8600 6350 8630
rect 6290 8560 6350 8600
rect 6290 8530 6305 8560
rect 6335 8530 6350 8560
rect 6290 8495 6350 8530
rect 6290 8465 6305 8495
rect 6335 8465 6350 8495
rect 6290 8435 6350 8465
rect 6290 8405 6305 8435
rect 6335 8405 6350 8435
rect 6290 8370 6350 8405
rect 6290 8340 6305 8370
rect 6335 8340 6350 8370
rect 6290 8300 6350 8340
rect 6290 8270 6305 8300
rect 6335 8270 6350 8300
rect 6290 8230 6350 8270
rect 6290 8200 6305 8230
rect 6335 8200 6350 8230
rect 6290 8160 6350 8200
rect 6290 8130 6305 8160
rect 6335 8130 6350 8160
rect 6290 8095 6350 8130
rect 6290 8065 6305 8095
rect 6335 8065 6350 8095
rect 6290 8035 6350 8065
rect 6290 8005 6305 8035
rect 6335 8005 6350 8035
rect 6290 7970 6350 8005
rect 6290 7940 6305 7970
rect 6335 7940 6350 7970
rect 6290 7900 6350 7940
rect 6290 7870 6305 7900
rect 6335 7870 6350 7900
rect 6290 7830 6350 7870
rect 6290 7800 6305 7830
rect 6335 7800 6350 7830
rect 6290 7760 6350 7800
rect 6290 7730 6305 7760
rect 6335 7730 6350 7760
rect 6290 7695 6350 7730
rect 6290 7665 6305 7695
rect 6335 7665 6350 7695
rect 6290 7635 6350 7665
rect 6290 7605 6305 7635
rect 6335 7605 6350 7635
rect 6290 7570 6350 7605
rect 6290 7540 6305 7570
rect 6335 7540 6350 7570
rect 6290 7500 6350 7540
rect 6290 7470 6305 7500
rect 6335 7470 6350 7500
rect 6290 7430 6350 7470
rect 6290 7400 6305 7430
rect 6335 7400 6350 7430
rect 6290 7360 6350 7400
rect 6290 7330 6305 7360
rect 6335 7330 6350 7360
rect 6290 7295 6350 7330
rect 6290 7265 6305 7295
rect 6335 7265 6350 7295
rect 6290 7235 6350 7265
rect 6290 7205 6305 7235
rect 6335 7205 6350 7235
rect 6290 7170 6350 7205
rect 6290 7140 6305 7170
rect 6335 7140 6350 7170
rect 6290 7100 6350 7140
rect 6290 7070 6305 7100
rect 6335 7070 6350 7100
rect 6290 7030 6350 7070
rect 6290 7000 6305 7030
rect 6335 7000 6350 7030
rect 6290 6960 6350 7000
rect 6290 6930 6305 6960
rect 6335 6930 6350 6960
rect 6290 6895 6350 6930
rect 6290 6865 6305 6895
rect 6335 6865 6350 6895
rect 6290 6835 6350 6865
rect 6290 6805 6305 6835
rect 6335 6805 6350 6835
rect 6290 6770 6350 6805
rect 6290 6740 6305 6770
rect 6335 6740 6350 6770
rect 6290 6700 6350 6740
rect 6290 6670 6305 6700
rect 6335 6670 6350 6700
rect 6290 6630 6350 6670
rect 6290 6600 6305 6630
rect 6335 6600 6350 6630
rect 6290 6560 6350 6600
rect 6290 6530 6305 6560
rect 6335 6530 6350 6560
rect 6290 6495 6350 6530
rect 6290 6465 6305 6495
rect 6335 6465 6350 6495
rect 6290 6450 6350 6465
rect 6580 9635 6640 9650
rect 6580 9605 6595 9635
rect 6625 9605 6640 9635
rect 6580 9570 6640 9605
rect 6580 9540 6595 9570
rect 6625 9540 6640 9570
rect 6580 9500 6640 9540
rect 6580 9470 6595 9500
rect 6625 9470 6640 9500
rect 6580 9430 6640 9470
rect 6580 9400 6595 9430
rect 6625 9400 6640 9430
rect 6580 9360 6640 9400
rect 6580 9330 6595 9360
rect 6625 9330 6640 9360
rect 6580 9295 6640 9330
rect 6580 9265 6595 9295
rect 6625 9265 6640 9295
rect 6580 9235 6640 9265
rect 6580 9205 6595 9235
rect 6625 9205 6640 9235
rect 6580 9170 6640 9205
rect 6580 9140 6595 9170
rect 6625 9140 6640 9170
rect 6580 9100 6640 9140
rect 6580 9070 6595 9100
rect 6625 9070 6640 9100
rect 6580 9030 6640 9070
rect 6580 9000 6595 9030
rect 6625 9000 6640 9030
rect 6580 8960 6640 9000
rect 6580 8930 6595 8960
rect 6625 8930 6640 8960
rect 6580 8895 6640 8930
rect 6580 8865 6595 8895
rect 6625 8865 6640 8895
rect 6580 8835 6640 8865
rect 6580 8805 6595 8835
rect 6625 8805 6640 8835
rect 6580 8770 6640 8805
rect 6580 8740 6595 8770
rect 6625 8740 6640 8770
rect 6580 8700 6640 8740
rect 6580 8670 6595 8700
rect 6625 8670 6640 8700
rect 6580 8630 6640 8670
rect 6580 8600 6595 8630
rect 6625 8600 6640 8630
rect 6580 8560 6640 8600
rect 6580 8530 6595 8560
rect 6625 8530 6640 8560
rect 6580 8495 6640 8530
rect 6580 8465 6595 8495
rect 6625 8465 6640 8495
rect 6580 8435 6640 8465
rect 6580 8405 6595 8435
rect 6625 8405 6640 8435
rect 6580 8370 6640 8405
rect 6580 8340 6595 8370
rect 6625 8340 6640 8370
rect 6580 8300 6640 8340
rect 6580 8270 6595 8300
rect 6625 8270 6640 8300
rect 6580 8230 6640 8270
rect 6580 8200 6595 8230
rect 6625 8200 6640 8230
rect 6580 8160 6640 8200
rect 6580 8130 6595 8160
rect 6625 8130 6640 8160
rect 6580 8095 6640 8130
rect 6580 8065 6595 8095
rect 6625 8065 6640 8095
rect 6580 8035 6640 8065
rect 6580 8005 6595 8035
rect 6625 8005 6640 8035
rect 6580 7970 6640 8005
rect 6580 7940 6595 7970
rect 6625 7940 6640 7970
rect 6580 7900 6640 7940
rect 6580 7870 6595 7900
rect 6625 7870 6640 7900
rect 6580 7830 6640 7870
rect 6580 7800 6595 7830
rect 6625 7800 6640 7830
rect 6580 7760 6640 7800
rect 6580 7730 6595 7760
rect 6625 7730 6640 7760
rect 6580 7695 6640 7730
rect 6580 7665 6595 7695
rect 6625 7665 6640 7695
rect 6580 7635 6640 7665
rect 6580 7605 6595 7635
rect 6625 7605 6640 7635
rect 6580 7570 6640 7605
rect 6580 7540 6595 7570
rect 6625 7540 6640 7570
rect 6580 7500 6640 7540
rect 6580 7470 6595 7500
rect 6625 7470 6640 7500
rect 6580 7430 6640 7470
rect 6580 7400 6595 7430
rect 6625 7400 6640 7430
rect 6580 7360 6640 7400
rect 6580 7330 6595 7360
rect 6625 7330 6640 7360
rect 6580 7295 6640 7330
rect 6580 7265 6595 7295
rect 6625 7265 6640 7295
rect 6580 7235 6640 7265
rect 6580 7205 6595 7235
rect 6625 7205 6640 7235
rect 6580 7170 6640 7205
rect 6580 7140 6595 7170
rect 6625 7140 6640 7170
rect 6580 7100 6640 7140
rect 6580 7070 6595 7100
rect 6625 7070 6640 7100
rect 6580 7030 6640 7070
rect 6580 7000 6595 7030
rect 6625 7000 6640 7030
rect 6580 6960 6640 7000
rect 6580 6930 6595 6960
rect 6625 6930 6640 6960
rect 6580 6895 6640 6930
rect 6580 6865 6595 6895
rect 6625 6865 6640 6895
rect 6580 6835 6640 6865
rect 6580 6805 6595 6835
rect 6625 6805 6640 6835
rect 6580 6770 6640 6805
rect 6580 6740 6595 6770
rect 6625 6740 6640 6770
rect 6580 6700 6640 6740
rect 6580 6670 6595 6700
rect 6625 6670 6640 6700
rect 6580 6630 6640 6670
rect 6580 6600 6595 6630
rect 6625 6600 6640 6630
rect 6580 6560 6640 6600
rect 6580 6530 6595 6560
rect 6625 6530 6640 6560
rect 6580 6495 6640 6530
rect 6580 6465 6595 6495
rect 6625 6465 6640 6495
rect 6580 6450 6640 6465
rect 7260 9635 7320 9650
rect 7260 9605 7275 9635
rect 7305 9605 7320 9635
rect 7260 9570 7320 9605
rect 7260 9540 7275 9570
rect 7305 9540 7320 9570
rect 7260 9500 7320 9540
rect 7260 9470 7275 9500
rect 7305 9470 7320 9500
rect 7260 9430 7320 9470
rect 7260 9400 7275 9430
rect 7305 9400 7320 9430
rect 7260 9360 7320 9400
rect 7260 9330 7275 9360
rect 7305 9330 7320 9360
rect 7260 9295 7320 9330
rect 7260 9265 7275 9295
rect 7305 9265 7320 9295
rect 7260 9235 7320 9265
rect 7260 9205 7275 9235
rect 7305 9205 7320 9235
rect 7260 9170 7320 9205
rect 7260 9140 7275 9170
rect 7305 9140 7320 9170
rect 7260 9100 7320 9140
rect 7260 9070 7275 9100
rect 7305 9070 7320 9100
rect 7260 9030 7320 9070
rect 7260 9000 7275 9030
rect 7305 9000 7320 9030
rect 7260 8960 7320 9000
rect 7260 8930 7275 8960
rect 7305 8930 7320 8960
rect 7260 8895 7320 8930
rect 7260 8865 7275 8895
rect 7305 8865 7320 8895
rect 7260 8835 7320 8865
rect 7260 8805 7275 8835
rect 7305 8805 7320 8835
rect 7260 8770 7320 8805
rect 7260 8740 7275 8770
rect 7305 8740 7320 8770
rect 7260 8700 7320 8740
rect 7260 8670 7275 8700
rect 7305 8670 7320 8700
rect 7260 8630 7320 8670
rect 7260 8600 7275 8630
rect 7305 8600 7320 8630
rect 7260 8560 7320 8600
rect 7260 8530 7275 8560
rect 7305 8530 7320 8560
rect 7260 8495 7320 8530
rect 7260 8465 7275 8495
rect 7305 8465 7320 8495
rect 7260 8435 7320 8465
rect 7260 8405 7275 8435
rect 7305 8405 7320 8435
rect 7260 8370 7320 8405
rect 7260 8340 7275 8370
rect 7305 8340 7320 8370
rect 7260 8300 7320 8340
rect 7260 8270 7275 8300
rect 7305 8270 7320 8300
rect 7260 8230 7320 8270
rect 7260 8200 7275 8230
rect 7305 8200 7320 8230
rect 7260 8160 7320 8200
rect 7260 8130 7275 8160
rect 7305 8130 7320 8160
rect 7260 8095 7320 8130
rect 7260 8065 7275 8095
rect 7305 8065 7320 8095
rect 7260 8035 7320 8065
rect 7260 8005 7275 8035
rect 7305 8005 7320 8035
rect 7260 7970 7320 8005
rect 7260 7940 7275 7970
rect 7305 7940 7320 7970
rect 7260 7900 7320 7940
rect 7260 7870 7275 7900
rect 7305 7870 7320 7900
rect 7260 7830 7320 7870
rect 7260 7800 7275 7830
rect 7305 7800 7320 7830
rect 7260 7760 7320 7800
rect 7260 7730 7275 7760
rect 7305 7730 7320 7760
rect 7260 7695 7320 7730
rect 7260 7665 7275 7695
rect 7305 7665 7320 7695
rect 7260 7635 7320 7665
rect 7260 7605 7275 7635
rect 7305 7605 7320 7635
rect 7260 7570 7320 7605
rect 7260 7540 7275 7570
rect 7305 7540 7320 7570
rect 7260 7500 7320 7540
rect 7260 7470 7275 7500
rect 7305 7470 7320 7500
rect 7260 7430 7320 7470
rect 7260 7400 7275 7430
rect 7305 7400 7320 7430
rect 7260 7360 7320 7400
rect 7260 7330 7275 7360
rect 7305 7330 7320 7360
rect 7260 7295 7320 7330
rect 7260 7265 7275 7295
rect 7305 7265 7320 7295
rect 7260 7235 7320 7265
rect 7260 7205 7275 7235
rect 7305 7205 7320 7235
rect 7260 7170 7320 7205
rect 7260 7140 7275 7170
rect 7305 7140 7320 7170
rect 7260 7100 7320 7140
rect 7260 7070 7275 7100
rect 7305 7070 7320 7100
rect 7260 7030 7320 7070
rect 7260 7000 7275 7030
rect 7305 7000 7320 7030
rect 7260 6960 7320 7000
rect 7260 6930 7275 6960
rect 7305 6930 7320 6960
rect 7260 6895 7320 6930
rect 7260 6865 7275 6895
rect 7305 6865 7320 6895
rect 7260 6835 7320 6865
rect 7260 6805 7275 6835
rect 7305 6805 7320 6835
rect 7260 6770 7320 6805
rect 7260 6740 7275 6770
rect 7305 6740 7320 6770
rect 7260 6700 7320 6740
rect 7260 6670 7275 6700
rect 7305 6670 7320 6700
rect 7260 6630 7320 6670
rect 7260 6600 7275 6630
rect 7305 6600 7320 6630
rect 7260 6560 7320 6600
rect 7260 6530 7275 6560
rect 7305 6530 7320 6560
rect 7260 6495 7320 6530
rect 7260 6465 7275 6495
rect 7305 6465 7320 6495
rect 7260 6450 7320 6465
rect 7610 9635 7670 9650
rect 7610 9605 7625 9635
rect 7655 9605 7670 9635
rect 7610 9570 7670 9605
rect 7610 9540 7625 9570
rect 7655 9540 7670 9570
rect 7610 9500 7670 9540
rect 7610 9470 7625 9500
rect 7655 9470 7670 9500
rect 7610 9430 7670 9470
rect 7610 9400 7625 9430
rect 7655 9400 7670 9430
rect 7610 9360 7670 9400
rect 7610 9330 7625 9360
rect 7655 9330 7670 9360
rect 7610 9295 7670 9330
rect 7610 9265 7625 9295
rect 7655 9265 7670 9295
rect 7610 9235 7670 9265
rect 7610 9205 7625 9235
rect 7655 9205 7670 9235
rect 7610 9170 7670 9205
rect 7610 9140 7625 9170
rect 7655 9140 7670 9170
rect 7610 9100 7670 9140
rect 7610 9070 7625 9100
rect 7655 9070 7670 9100
rect 7610 9030 7670 9070
rect 7610 9000 7625 9030
rect 7655 9000 7670 9030
rect 7610 8960 7670 9000
rect 7610 8930 7625 8960
rect 7655 8930 7670 8960
rect 7610 8895 7670 8930
rect 7610 8865 7625 8895
rect 7655 8865 7670 8895
rect 7610 8835 7670 8865
rect 7610 8805 7625 8835
rect 7655 8805 7670 8835
rect 7610 8770 7670 8805
rect 7610 8740 7625 8770
rect 7655 8740 7670 8770
rect 7610 8700 7670 8740
rect 7610 8670 7625 8700
rect 7655 8670 7670 8700
rect 7610 8630 7670 8670
rect 7610 8600 7625 8630
rect 7655 8600 7670 8630
rect 7610 8560 7670 8600
rect 7610 8530 7625 8560
rect 7655 8530 7670 8560
rect 7610 8495 7670 8530
rect 7610 8465 7625 8495
rect 7655 8465 7670 8495
rect 7610 8435 7670 8465
rect 7610 8405 7625 8435
rect 7655 8405 7670 8435
rect 7610 8370 7670 8405
rect 7610 8340 7625 8370
rect 7655 8340 7670 8370
rect 7610 8300 7670 8340
rect 7610 8270 7625 8300
rect 7655 8270 7670 8300
rect 7610 8230 7670 8270
rect 7610 8200 7625 8230
rect 7655 8200 7670 8230
rect 7610 8160 7670 8200
rect 7610 8130 7625 8160
rect 7655 8130 7670 8160
rect 7610 8095 7670 8130
rect 7610 8065 7625 8095
rect 7655 8065 7670 8095
rect 7610 8035 7670 8065
rect 7610 8005 7625 8035
rect 7655 8005 7670 8035
rect 7610 7970 7670 8005
rect 7610 7940 7625 7970
rect 7655 7940 7670 7970
rect 7610 7900 7670 7940
rect 7610 7870 7625 7900
rect 7655 7870 7670 7900
rect 7610 7830 7670 7870
rect 7610 7800 7625 7830
rect 7655 7800 7670 7830
rect 7610 7760 7670 7800
rect 7610 7730 7625 7760
rect 7655 7730 7670 7760
rect 7610 7695 7670 7730
rect 7610 7665 7625 7695
rect 7655 7665 7670 7695
rect 7610 7635 7670 7665
rect 7610 7605 7625 7635
rect 7655 7605 7670 7635
rect 7610 7570 7670 7605
rect 7610 7540 7625 7570
rect 7655 7540 7670 7570
rect 7610 7500 7670 7540
rect 7610 7470 7625 7500
rect 7655 7470 7670 7500
rect 7610 7430 7670 7470
rect 7610 7400 7625 7430
rect 7655 7400 7670 7430
rect 7610 7360 7670 7400
rect 7610 7330 7625 7360
rect 7655 7330 7670 7360
rect 7610 7295 7670 7330
rect 7610 7265 7625 7295
rect 7655 7265 7670 7295
rect 7610 7235 7670 7265
rect 7610 7205 7625 7235
rect 7655 7205 7670 7235
rect 7610 7170 7670 7205
rect 7610 7140 7625 7170
rect 7655 7140 7670 7170
rect 7610 7100 7670 7140
rect 7610 7070 7625 7100
rect 7655 7070 7670 7100
rect 7610 7030 7670 7070
rect 7610 7000 7625 7030
rect 7655 7000 7670 7030
rect 7610 6960 7670 7000
rect 7610 6930 7625 6960
rect 7655 6930 7670 6960
rect 7610 6895 7670 6930
rect 7610 6865 7625 6895
rect 7655 6865 7670 6895
rect 7610 6835 7670 6865
rect 7610 6805 7625 6835
rect 7655 6805 7670 6835
rect 7610 6770 7670 6805
rect 7610 6740 7625 6770
rect 7655 6740 7670 6770
rect 7610 6700 7670 6740
rect 7610 6670 7625 6700
rect 7655 6670 7670 6700
rect 7610 6630 7670 6670
rect 7610 6600 7625 6630
rect 7655 6600 7670 6630
rect 7610 6560 7670 6600
rect 7610 6530 7625 6560
rect 7655 6530 7670 6560
rect 7610 6495 7670 6530
rect 7610 6465 7625 6495
rect 7655 6465 7670 6495
rect 7610 6450 7670 6465
rect 8310 9635 8370 9650
rect 8310 9605 8325 9635
rect 8355 9605 8370 9635
rect 8310 9570 8370 9605
rect 8310 9540 8325 9570
rect 8355 9540 8370 9570
rect 8310 9500 8370 9540
rect 8310 9470 8325 9500
rect 8355 9470 8370 9500
rect 8310 9430 8370 9470
rect 8310 9400 8325 9430
rect 8355 9400 8370 9430
rect 8310 9360 8370 9400
rect 8310 9330 8325 9360
rect 8355 9330 8370 9360
rect 8310 9295 8370 9330
rect 8310 9265 8325 9295
rect 8355 9265 8370 9295
rect 8310 9235 8370 9265
rect 8310 9205 8325 9235
rect 8355 9205 8370 9235
rect 8310 9170 8370 9205
rect 8310 9140 8325 9170
rect 8355 9140 8370 9170
rect 8310 9100 8370 9140
rect 8310 9070 8325 9100
rect 8355 9070 8370 9100
rect 8310 9030 8370 9070
rect 8310 9000 8325 9030
rect 8355 9000 8370 9030
rect 8310 8960 8370 9000
rect 8310 8930 8325 8960
rect 8355 8930 8370 8960
rect 8310 8895 8370 8930
rect 8310 8865 8325 8895
rect 8355 8865 8370 8895
rect 8310 8835 8370 8865
rect 8310 8805 8325 8835
rect 8355 8805 8370 8835
rect 8310 8770 8370 8805
rect 8310 8740 8325 8770
rect 8355 8740 8370 8770
rect 8310 8700 8370 8740
rect 8310 8670 8325 8700
rect 8355 8670 8370 8700
rect 8310 8630 8370 8670
rect 8310 8600 8325 8630
rect 8355 8600 8370 8630
rect 8310 8560 8370 8600
rect 8310 8530 8325 8560
rect 8355 8530 8370 8560
rect 8310 8495 8370 8530
rect 8310 8465 8325 8495
rect 8355 8465 8370 8495
rect 8310 8435 8370 8465
rect 8310 8405 8325 8435
rect 8355 8405 8370 8435
rect 8310 8370 8370 8405
rect 8310 8340 8325 8370
rect 8355 8340 8370 8370
rect 8310 8300 8370 8340
rect 8310 8270 8325 8300
rect 8355 8270 8370 8300
rect 8310 8230 8370 8270
rect 8310 8200 8325 8230
rect 8355 8200 8370 8230
rect 8310 8160 8370 8200
rect 8310 8130 8325 8160
rect 8355 8130 8370 8160
rect 8310 8095 8370 8130
rect 8310 8065 8325 8095
rect 8355 8065 8370 8095
rect 8310 8035 8370 8065
rect 8310 8005 8325 8035
rect 8355 8005 8370 8035
rect 8310 7970 8370 8005
rect 8310 7940 8325 7970
rect 8355 7940 8370 7970
rect 8310 7900 8370 7940
rect 8310 7870 8325 7900
rect 8355 7870 8370 7900
rect 8310 7830 8370 7870
rect 8310 7800 8325 7830
rect 8355 7800 8370 7830
rect 8310 7760 8370 7800
rect 8310 7730 8325 7760
rect 8355 7730 8370 7760
rect 8310 7695 8370 7730
rect 8310 7665 8325 7695
rect 8355 7665 8370 7695
rect 8310 7635 8370 7665
rect 8310 7605 8325 7635
rect 8355 7605 8370 7635
rect 8310 7570 8370 7605
rect 8310 7540 8325 7570
rect 8355 7540 8370 7570
rect 8310 7500 8370 7540
rect 8310 7470 8325 7500
rect 8355 7470 8370 7500
rect 8310 7430 8370 7470
rect 8310 7400 8325 7430
rect 8355 7400 8370 7430
rect 8310 7360 8370 7400
rect 8310 7330 8325 7360
rect 8355 7330 8370 7360
rect 8310 7295 8370 7330
rect 8310 7265 8325 7295
rect 8355 7265 8370 7295
rect 8310 7235 8370 7265
rect 8310 7205 8325 7235
rect 8355 7205 8370 7235
rect 8310 7170 8370 7205
rect 8310 7140 8325 7170
rect 8355 7140 8370 7170
rect 8310 7100 8370 7140
rect 8310 7070 8325 7100
rect 8355 7070 8370 7100
rect 8310 7030 8370 7070
rect 8310 7000 8325 7030
rect 8355 7000 8370 7030
rect 8310 6960 8370 7000
rect 8310 6930 8325 6960
rect 8355 6930 8370 6960
rect 8310 6895 8370 6930
rect 8310 6865 8325 6895
rect 8355 6865 8370 6895
rect 8310 6835 8370 6865
rect 8310 6805 8325 6835
rect 8355 6805 8370 6835
rect 8310 6770 8370 6805
rect 8310 6740 8325 6770
rect 8355 6740 8370 6770
rect 8310 6700 8370 6740
rect 8310 6670 8325 6700
rect 8355 6670 8370 6700
rect 8310 6630 8370 6670
rect 8310 6600 8325 6630
rect 8355 6600 8370 6630
rect 8310 6560 8370 6600
rect 8310 6530 8325 6560
rect 8355 6530 8370 6560
rect 8310 6495 8370 6530
rect 8310 6465 8325 6495
rect 8355 6465 8370 6495
rect 8310 6450 8370 6465
rect 8660 9635 8720 9650
rect 8660 9605 8675 9635
rect 8705 9605 8720 9635
rect 8660 9570 8720 9605
rect 8660 9540 8675 9570
rect 8705 9540 8720 9570
rect 8660 9500 8720 9540
rect 8660 9470 8675 9500
rect 8705 9470 8720 9500
rect 8660 9430 8720 9470
rect 8660 9400 8675 9430
rect 8705 9400 8720 9430
rect 8660 9360 8720 9400
rect 8660 9330 8675 9360
rect 8705 9330 8720 9360
rect 8660 9295 8720 9330
rect 8660 9265 8675 9295
rect 8705 9265 8720 9295
rect 8660 9235 8720 9265
rect 8660 9205 8675 9235
rect 8705 9205 8720 9235
rect 8660 9170 8720 9205
rect 8660 9140 8675 9170
rect 8705 9140 8720 9170
rect 8660 9100 8720 9140
rect 8660 9070 8675 9100
rect 8705 9070 8720 9100
rect 8660 9030 8720 9070
rect 8660 9000 8675 9030
rect 8705 9000 8720 9030
rect 8660 8960 8720 9000
rect 8660 8930 8675 8960
rect 8705 8930 8720 8960
rect 8660 8895 8720 8930
rect 8660 8865 8675 8895
rect 8705 8865 8720 8895
rect 8660 8835 8720 8865
rect 8660 8805 8675 8835
rect 8705 8805 8720 8835
rect 8660 8770 8720 8805
rect 8660 8740 8675 8770
rect 8705 8740 8720 8770
rect 8660 8700 8720 8740
rect 8660 8670 8675 8700
rect 8705 8670 8720 8700
rect 8660 8630 8720 8670
rect 8660 8600 8675 8630
rect 8705 8600 8720 8630
rect 8660 8560 8720 8600
rect 8660 8530 8675 8560
rect 8705 8530 8720 8560
rect 8660 8495 8720 8530
rect 8660 8465 8675 8495
rect 8705 8465 8720 8495
rect 8660 8435 8720 8465
rect 8660 8405 8675 8435
rect 8705 8405 8720 8435
rect 8660 8370 8720 8405
rect 8660 8340 8675 8370
rect 8705 8340 8720 8370
rect 8660 8300 8720 8340
rect 8660 8270 8675 8300
rect 8705 8270 8720 8300
rect 8660 8230 8720 8270
rect 8660 8200 8675 8230
rect 8705 8200 8720 8230
rect 8660 8160 8720 8200
rect 8660 8130 8675 8160
rect 8705 8130 8720 8160
rect 8660 8095 8720 8130
rect 8660 8065 8675 8095
rect 8705 8065 8720 8095
rect 8660 8035 8720 8065
rect 8660 8005 8675 8035
rect 8705 8005 8720 8035
rect 8660 7970 8720 8005
rect 8660 7940 8675 7970
rect 8705 7940 8720 7970
rect 8660 7900 8720 7940
rect 8660 7870 8675 7900
rect 8705 7870 8720 7900
rect 8660 7830 8720 7870
rect 8660 7800 8675 7830
rect 8705 7800 8720 7830
rect 8660 7760 8720 7800
rect 8660 7730 8675 7760
rect 8705 7730 8720 7760
rect 8660 7695 8720 7730
rect 8660 7665 8675 7695
rect 8705 7665 8720 7695
rect 8660 7635 8720 7665
rect 8660 7605 8675 7635
rect 8705 7605 8720 7635
rect 8660 7570 8720 7605
rect 8660 7540 8675 7570
rect 8705 7540 8720 7570
rect 8660 7500 8720 7540
rect 8660 7470 8675 7500
rect 8705 7470 8720 7500
rect 8660 7430 8720 7470
rect 8660 7400 8675 7430
rect 8705 7400 8720 7430
rect 8660 7360 8720 7400
rect 8660 7330 8675 7360
rect 8705 7330 8720 7360
rect 8660 7295 8720 7330
rect 8660 7265 8675 7295
rect 8705 7265 8720 7295
rect 8660 7235 8720 7265
rect 8660 7205 8675 7235
rect 8705 7205 8720 7235
rect 8660 7170 8720 7205
rect 8660 7140 8675 7170
rect 8705 7140 8720 7170
rect 8660 7100 8720 7140
rect 8660 7070 8675 7100
rect 8705 7070 8720 7100
rect 8660 7030 8720 7070
rect 8660 7000 8675 7030
rect 8705 7000 8720 7030
rect 8660 6960 8720 7000
rect 8660 6930 8675 6960
rect 8705 6930 8720 6960
rect 8660 6895 8720 6930
rect 8660 6865 8675 6895
rect 8705 6865 8720 6895
rect 8660 6835 8720 6865
rect 8660 6805 8675 6835
rect 8705 6805 8720 6835
rect 8660 6770 8720 6805
rect 8660 6740 8675 6770
rect 8705 6740 8720 6770
rect 8660 6700 8720 6740
rect 8660 6670 8675 6700
rect 8705 6670 8720 6700
rect 8660 6630 8720 6670
rect 8660 6600 8675 6630
rect 8705 6600 8720 6630
rect 8660 6560 8720 6600
rect 8660 6530 8675 6560
rect 8705 6530 8720 6560
rect 8660 6495 8720 6530
rect 8660 6465 8675 6495
rect 8705 6465 8720 6495
rect 8660 6450 8720 6465
rect 9010 9635 9070 9650
rect 9010 9605 9025 9635
rect 9055 9605 9070 9635
rect 9010 9570 9070 9605
rect 9010 9540 9025 9570
rect 9055 9540 9070 9570
rect 9010 9500 9070 9540
rect 9010 9470 9025 9500
rect 9055 9470 9070 9500
rect 9010 9430 9070 9470
rect 9010 9400 9025 9430
rect 9055 9400 9070 9430
rect 9010 9360 9070 9400
rect 9010 9330 9025 9360
rect 9055 9330 9070 9360
rect 9010 9295 9070 9330
rect 9010 9265 9025 9295
rect 9055 9265 9070 9295
rect 9010 9235 9070 9265
rect 9010 9205 9025 9235
rect 9055 9205 9070 9235
rect 9010 9170 9070 9205
rect 9010 9140 9025 9170
rect 9055 9140 9070 9170
rect 9010 9100 9070 9140
rect 9010 9070 9025 9100
rect 9055 9070 9070 9100
rect 9010 9030 9070 9070
rect 9010 9000 9025 9030
rect 9055 9000 9070 9030
rect 9010 8960 9070 9000
rect 9010 8930 9025 8960
rect 9055 8930 9070 8960
rect 9010 8895 9070 8930
rect 9010 8865 9025 8895
rect 9055 8865 9070 8895
rect 9010 8835 9070 8865
rect 9010 8805 9025 8835
rect 9055 8805 9070 8835
rect 9010 8770 9070 8805
rect 9010 8740 9025 8770
rect 9055 8740 9070 8770
rect 9010 8700 9070 8740
rect 9010 8670 9025 8700
rect 9055 8670 9070 8700
rect 9010 8630 9070 8670
rect 9010 8600 9025 8630
rect 9055 8600 9070 8630
rect 9010 8560 9070 8600
rect 9010 8530 9025 8560
rect 9055 8530 9070 8560
rect 9010 8495 9070 8530
rect 9010 8465 9025 8495
rect 9055 8465 9070 8495
rect 9010 8435 9070 8465
rect 9010 8405 9025 8435
rect 9055 8405 9070 8435
rect 9010 8370 9070 8405
rect 9010 8340 9025 8370
rect 9055 8340 9070 8370
rect 9010 8300 9070 8340
rect 9010 8270 9025 8300
rect 9055 8270 9070 8300
rect 9010 8230 9070 8270
rect 9010 8200 9025 8230
rect 9055 8200 9070 8230
rect 9010 8160 9070 8200
rect 9010 8130 9025 8160
rect 9055 8130 9070 8160
rect 9010 8095 9070 8130
rect 9010 8065 9025 8095
rect 9055 8065 9070 8095
rect 9010 8035 9070 8065
rect 9010 8005 9025 8035
rect 9055 8005 9070 8035
rect 9010 7970 9070 8005
rect 9010 7940 9025 7970
rect 9055 7940 9070 7970
rect 9010 7900 9070 7940
rect 9010 7870 9025 7900
rect 9055 7870 9070 7900
rect 9010 7830 9070 7870
rect 9010 7800 9025 7830
rect 9055 7800 9070 7830
rect 9010 7760 9070 7800
rect 9010 7730 9025 7760
rect 9055 7730 9070 7760
rect 9010 7695 9070 7730
rect 9010 7665 9025 7695
rect 9055 7665 9070 7695
rect 9010 7635 9070 7665
rect 9010 7605 9025 7635
rect 9055 7605 9070 7635
rect 9010 7570 9070 7605
rect 9010 7540 9025 7570
rect 9055 7540 9070 7570
rect 9010 7500 9070 7540
rect 9010 7470 9025 7500
rect 9055 7470 9070 7500
rect 9010 7430 9070 7470
rect 9010 7400 9025 7430
rect 9055 7400 9070 7430
rect 9010 7360 9070 7400
rect 9010 7330 9025 7360
rect 9055 7330 9070 7360
rect 9010 7295 9070 7330
rect 9010 7265 9025 7295
rect 9055 7265 9070 7295
rect 9010 7235 9070 7265
rect 9010 7205 9025 7235
rect 9055 7205 9070 7235
rect 9010 7170 9070 7205
rect 9010 7140 9025 7170
rect 9055 7140 9070 7170
rect 9010 7100 9070 7140
rect 9010 7070 9025 7100
rect 9055 7070 9070 7100
rect 9010 7030 9070 7070
rect 9010 7000 9025 7030
rect 9055 7000 9070 7030
rect 9010 6960 9070 7000
rect 9010 6930 9025 6960
rect 9055 6930 9070 6960
rect 9010 6895 9070 6930
rect 9010 6865 9025 6895
rect 9055 6865 9070 6895
rect 9010 6835 9070 6865
rect 9010 6805 9025 6835
rect 9055 6805 9070 6835
rect 9010 6770 9070 6805
rect 9010 6740 9025 6770
rect 9055 6740 9070 6770
rect 9010 6700 9070 6740
rect 9010 6670 9025 6700
rect 9055 6670 9070 6700
rect 9010 6630 9070 6670
rect 9010 6600 9025 6630
rect 9055 6600 9070 6630
rect 9010 6560 9070 6600
rect 9010 6530 9025 6560
rect 9055 6530 9070 6560
rect 9010 6495 9070 6530
rect 9010 6465 9025 6495
rect 9055 6465 9070 6495
rect 9010 6450 9070 6465
rect 2845 6440 2885 6445
rect 2045 6430 2515 6435
rect 2045 6400 2050 6430
rect 2080 6400 2480 6430
rect 2510 6400 2515 6430
rect 2845 6410 2850 6440
rect 2880 6435 2885 6440
rect 3400 6440 3440 6445
rect 3400 6435 3405 6440
rect 2880 6415 3405 6435
rect 2880 6410 2885 6415
rect 2845 6405 2885 6410
rect 3400 6410 3405 6415
rect 3435 6410 3440 6440
rect 3400 6405 3440 6410
rect 5490 6430 5530 6435
rect 2045 6395 2515 6400
rect 5490 6400 5495 6430
rect 5525 6425 5530 6430
rect 6145 6430 6185 6435
rect 6145 6425 6150 6430
rect 5525 6405 6150 6425
rect 5525 6400 5530 6405
rect 5490 6395 5530 6400
rect 6145 6400 6150 6405
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 6465 6430 6935 6435
rect 6465 6400 6470 6430
rect 6500 6400 6900 6430
rect 6930 6400 6935 6430
rect 6465 6395 6935 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6370 2040 6375
rect 3630 6375 3670 6380
rect 3630 6370 3635 6375
rect 2035 6350 3635 6370
rect 2035 6345 2040 6350
rect 2000 6340 2040 6345
rect 3630 6345 3635 6350
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6370 5350 6375
rect 6940 6375 6980 6380
rect 6940 6370 6945 6375
rect 5345 6350 6945 6370
rect 5345 6345 5350 6350
rect 5310 6340 5350 6345
rect 6940 6345 6945 6350
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6325 2755 6330
rect 4850 6330 4890 6335
rect 4850 6325 4855 6330
rect 2750 6305 4855 6325
rect 2750 6300 2755 6305
rect 2715 6295 2755 6300
rect 4850 6300 4855 6305
rect 4885 6300 4890 6330
rect 4850 6295 4890 6300
rect 2990 6285 3030 6290
rect 2990 6255 2995 6285
rect 3025 6280 3030 6285
rect 3455 6285 3495 6290
rect 3455 6280 3460 6285
rect 3025 6260 3460 6280
rect 3025 6255 3030 6260
rect 2990 6250 3030 6255
rect 3455 6255 3460 6260
rect 3490 6255 3495 6285
rect 3455 6250 3495 6255
rect 1280 6205 7700 6210
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 4310 6205
rect 4340 6175 4420 6205
rect 4450 6175 4530 6205
rect 4560 6175 4640 6205
rect 4670 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 1280 6165 7700 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 4310 6165
rect 4340 6135 4420 6165
rect 4450 6135 4530 6165
rect 4560 6135 4640 6165
rect 4670 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 1280 6125 7700 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 4310 6125
rect 4340 6095 4420 6125
rect 4450 6095 4530 6125
rect 4560 6095 4640 6125
rect 4670 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 1280 6090 7700 6095
rect 5870 5135 5910 5140
rect 5870 5105 5875 5135
rect 5905 5130 5910 5135
rect 6220 5135 6260 5140
rect 6220 5130 6225 5135
rect 5905 5110 6225 5130
rect 5905 5105 5910 5110
rect 5870 5100 5910 5105
rect 6220 5105 6225 5110
rect 6255 5105 6260 5135
rect 6220 5100 6260 5105
rect 4850 5015 4890 5020
rect 4940 5015 4980 5020
rect 4850 4985 4855 5015
rect 4885 4990 4945 5015
rect 4885 4985 4890 4990
rect 4850 4980 4890 4985
rect 4940 4985 4945 4990
rect 4975 4985 4980 5015
rect 4940 4980 4980 4985
rect 5870 4565 5910 4570
rect 5870 4560 5875 4565
rect 4515 4555 5875 4560
rect 4515 4540 5166 4555
rect 5196 4540 5875 4555
rect 5870 4535 5875 4540
rect 5905 4535 5910 4565
rect 5870 4530 5910 4535
rect 5166 4520 5196 4525
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 5490 3120 5530 3125
rect 5490 3110 5495 3120
rect 4720 3090 5495 3110
rect 5525 3090 5530 3120
rect 5490 3085 5530 3090
rect 3400 3055 3440 3060
rect 3400 3025 3405 3055
rect 3435 3050 3440 3055
rect 3435 3030 3955 3050
rect 3435 3025 3440 3030
rect 3400 3020 3440 3025
rect 2045 1755 2085 1760
rect 2045 1725 2050 1755
rect 2080 1750 2085 1755
rect 2175 1755 2215 1760
rect 2175 1750 2180 1755
rect 2080 1730 2180 1750
rect 2080 1725 2085 1730
rect 2045 1720 2085 1725
rect 2175 1725 2180 1730
rect 2210 1725 2215 1755
rect 3605 1745 3625 1765
rect 5355 1745 5375 1765
rect 6765 1755 6805 1760
rect 2175 1720 2215 1725
rect 6765 1725 6770 1755
rect 6800 1750 6805 1755
rect 6895 1755 6935 1760
rect 6895 1750 6900 1755
rect 6800 1730 6900 1750
rect 6800 1725 6805 1730
rect 6765 1720 6805 1725
rect 6895 1725 6900 1730
rect 6930 1725 6935 1755
rect 6895 1720 6935 1725
rect 2000 1700 2040 1705
rect 2000 1670 2005 1700
rect 2035 1695 2040 1700
rect 2100 1700 2140 1705
rect 2100 1695 2105 1700
rect 2035 1675 2105 1695
rect 2035 1670 2040 1675
rect 2000 1665 2040 1670
rect 2100 1670 2105 1675
rect 2135 1670 2140 1700
rect 2100 1665 2140 1670
rect 6830 1700 6870 1705
rect 6830 1670 6835 1700
rect 6865 1695 6870 1700
rect 6940 1700 6980 1705
rect 6940 1695 6945 1700
rect 6865 1675 6945 1695
rect 6865 1670 6870 1675
rect 6830 1665 6870 1670
rect 6940 1670 6945 1675
rect 6975 1670 6980 1700
rect 6940 1665 6980 1670
rect 1280 850 7700 855
rect 1280 820 1285 850
rect 1315 820 1325 850
rect 1355 820 1365 850
rect 1395 820 4420 850
rect 4450 820 4475 850
rect 4505 820 4530 850
rect 4560 820 7585 850
rect 7615 820 7625 850
rect 7655 820 7665 850
rect 7695 820 7700 850
rect 1280 810 7700 820
rect 1280 780 1285 810
rect 1315 780 1325 810
rect 1355 780 1365 810
rect 1395 780 4420 810
rect 4450 780 4475 810
rect 4505 780 4530 810
rect 4560 780 7585 810
rect 7615 780 7625 810
rect 7655 780 7665 810
rect 7695 780 7700 810
rect 1280 770 7700 780
rect 1280 740 1285 770
rect 1315 740 1325 770
rect 1355 740 1365 770
rect 1395 740 4420 770
rect 4450 740 4475 770
rect 4505 740 4530 770
rect 4560 740 7585 770
rect 7615 740 7625 770
rect 7655 740 7665 770
rect 7695 740 7700 770
rect 1280 735 7700 740
rect -90 -1305 -30 -1290
rect -90 -1335 -75 -1305
rect -45 -1335 -30 -1305
rect -90 -1370 -30 -1335
rect -90 -1400 -75 -1370
rect -45 -1400 -30 -1370
rect -90 -1440 -30 -1400
rect -90 -1470 -75 -1440
rect -45 -1470 -30 -1440
rect -90 -1510 -30 -1470
rect -90 -1540 -75 -1510
rect -45 -1540 -30 -1510
rect -90 -1580 -30 -1540
rect -90 -1610 -75 -1580
rect -45 -1610 -30 -1580
rect -90 -1645 -30 -1610
rect -90 -1675 -75 -1645
rect -45 -1675 -30 -1645
rect -90 -1705 -30 -1675
rect -90 -1735 -75 -1705
rect -45 -1735 -30 -1705
rect -90 -1770 -30 -1735
rect -90 -1800 -75 -1770
rect -45 -1800 -30 -1770
rect -90 -1840 -30 -1800
rect -90 -1870 -75 -1840
rect -45 -1870 -30 -1840
rect -90 -1910 -30 -1870
rect -90 -1940 -75 -1910
rect -45 -1940 -30 -1910
rect -90 -1980 -30 -1940
rect -90 -2010 -75 -1980
rect -45 -2010 -30 -1980
rect -90 -2045 -30 -2010
rect -90 -2075 -75 -2045
rect -45 -2075 -30 -2045
rect -90 -2105 -30 -2075
rect -90 -2135 -75 -2105
rect -45 -2135 -30 -2105
rect -90 -2170 -30 -2135
rect -90 -2200 -75 -2170
rect -45 -2200 -30 -2170
rect -90 -2240 -30 -2200
rect -90 -2270 -75 -2240
rect -45 -2270 -30 -2240
rect -90 -2310 -30 -2270
rect -90 -2340 -75 -2310
rect -45 -2340 -30 -2310
rect -90 -2380 -30 -2340
rect -90 -2410 -75 -2380
rect -45 -2410 -30 -2380
rect -90 -2445 -30 -2410
rect -90 -2475 -75 -2445
rect -45 -2475 -30 -2445
rect -90 -2505 -30 -2475
rect -90 -2535 -75 -2505
rect -45 -2535 -30 -2505
rect -90 -2570 -30 -2535
rect -90 -2600 -75 -2570
rect -45 -2600 -30 -2570
rect -90 -2640 -30 -2600
rect -90 -2670 -75 -2640
rect -45 -2670 -30 -2640
rect -90 -2710 -30 -2670
rect -90 -2740 -75 -2710
rect -45 -2740 -30 -2710
rect -90 -2780 -30 -2740
rect -90 -2810 -75 -2780
rect -45 -2810 -30 -2780
rect -90 -2845 -30 -2810
rect -90 -2875 -75 -2845
rect -45 -2875 -30 -2845
rect -90 -2905 -30 -2875
rect -90 -2935 -75 -2905
rect -45 -2935 -30 -2905
rect -90 -2970 -30 -2935
rect -90 -3000 -75 -2970
rect -45 -3000 -30 -2970
rect -90 -3040 -30 -3000
rect -90 -3070 -75 -3040
rect -45 -3070 -30 -3040
rect -90 -3110 -30 -3070
rect -90 -3140 -75 -3110
rect -45 -3140 -30 -3110
rect -90 -3180 -30 -3140
rect -90 -3210 -75 -3180
rect -45 -3210 -30 -3180
rect -90 -3245 -30 -3210
rect -90 -3275 -75 -3245
rect -45 -3275 -30 -3245
rect -90 -3305 -30 -3275
rect -90 -3335 -75 -3305
rect -45 -3335 -30 -3305
rect -90 -3370 -30 -3335
rect -90 -3400 -75 -3370
rect -45 -3400 -30 -3370
rect -90 -3440 -30 -3400
rect -90 -3470 -75 -3440
rect -45 -3470 -30 -3440
rect -90 -3510 -30 -3470
rect -90 -3540 -75 -3510
rect -45 -3540 -30 -3510
rect -90 -3580 -30 -3540
rect -90 -3610 -75 -3580
rect -45 -3610 -30 -3580
rect -90 -3645 -30 -3610
rect -90 -3675 -75 -3645
rect -45 -3675 -30 -3645
rect -90 -3705 -30 -3675
rect -90 -3735 -75 -3705
rect -45 -3735 -30 -3705
rect -90 -3770 -30 -3735
rect -90 -3800 -75 -3770
rect -45 -3800 -30 -3770
rect -90 -3840 -30 -3800
rect -90 -3870 -75 -3840
rect -45 -3870 -30 -3840
rect -90 -3910 -30 -3870
rect -90 -3940 -75 -3910
rect -45 -3940 -30 -3910
rect -90 -3980 -30 -3940
rect -90 -4010 -75 -3980
rect -45 -4010 -30 -3980
rect -90 -4045 -30 -4010
rect -90 -4075 -75 -4045
rect -45 -4075 -30 -4045
rect -90 -4105 -30 -4075
rect -90 -4135 -75 -4105
rect -45 -4135 -30 -4105
rect -90 -4170 -30 -4135
rect -90 -4200 -75 -4170
rect -45 -4200 -30 -4170
rect -90 -4240 -30 -4200
rect -90 -4270 -75 -4240
rect -45 -4270 -30 -4240
rect -90 -4310 -30 -4270
rect -90 -4340 -75 -4310
rect -45 -4340 -30 -4310
rect -90 -4380 -30 -4340
rect -90 -4410 -75 -4380
rect -45 -4410 -30 -4380
rect -90 -4445 -30 -4410
rect -90 -4475 -75 -4445
rect -45 -4475 -30 -4445
rect -90 -4490 -30 -4475
rect 260 -1305 320 -1290
rect 260 -1335 275 -1305
rect 305 -1335 320 -1305
rect 260 -1370 320 -1335
rect 260 -1400 275 -1370
rect 305 -1400 320 -1370
rect 260 -1440 320 -1400
rect 260 -1470 275 -1440
rect 305 -1470 320 -1440
rect 260 -1510 320 -1470
rect 260 -1540 275 -1510
rect 305 -1540 320 -1510
rect 260 -1580 320 -1540
rect 260 -1610 275 -1580
rect 305 -1610 320 -1580
rect 260 -1645 320 -1610
rect 260 -1675 275 -1645
rect 305 -1675 320 -1645
rect 260 -1705 320 -1675
rect 260 -1735 275 -1705
rect 305 -1735 320 -1705
rect 260 -1770 320 -1735
rect 260 -1800 275 -1770
rect 305 -1800 320 -1770
rect 260 -1840 320 -1800
rect 260 -1870 275 -1840
rect 305 -1870 320 -1840
rect 260 -1910 320 -1870
rect 260 -1940 275 -1910
rect 305 -1940 320 -1910
rect 260 -1980 320 -1940
rect 260 -2010 275 -1980
rect 305 -2010 320 -1980
rect 260 -2045 320 -2010
rect 260 -2075 275 -2045
rect 305 -2075 320 -2045
rect 260 -2105 320 -2075
rect 260 -2135 275 -2105
rect 305 -2135 320 -2105
rect 260 -2170 320 -2135
rect 260 -2200 275 -2170
rect 305 -2200 320 -2170
rect 260 -2240 320 -2200
rect 260 -2270 275 -2240
rect 305 -2270 320 -2240
rect 260 -2310 320 -2270
rect 260 -2340 275 -2310
rect 305 -2340 320 -2310
rect 260 -2380 320 -2340
rect 260 -2410 275 -2380
rect 305 -2410 320 -2380
rect 260 -2445 320 -2410
rect 260 -2475 275 -2445
rect 305 -2475 320 -2445
rect 260 -2505 320 -2475
rect 260 -2535 275 -2505
rect 305 -2535 320 -2505
rect 260 -2570 320 -2535
rect 260 -2600 275 -2570
rect 305 -2600 320 -2570
rect 260 -2640 320 -2600
rect 260 -2670 275 -2640
rect 305 -2670 320 -2640
rect 260 -2710 320 -2670
rect 260 -2740 275 -2710
rect 305 -2740 320 -2710
rect 260 -2780 320 -2740
rect 260 -2810 275 -2780
rect 305 -2810 320 -2780
rect 260 -2845 320 -2810
rect 260 -2875 275 -2845
rect 305 -2875 320 -2845
rect 260 -2905 320 -2875
rect 260 -2935 275 -2905
rect 305 -2935 320 -2905
rect 260 -2970 320 -2935
rect 260 -3000 275 -2970
rect 305 -3000 320 -2970
rect 260 -3040 320 -3000
rect 260 -3070 275 -3040
rect 305 -3070 320 -3040
rect 260 -3110 320 -3070
rect 260 -3140 275 -3110
rect 305 -3140 320 -3110
rect 260 -3180 320 -3140
rect 260 -3210 275 -3180
rect 305 -3210 320 -3180
rect 260 -3245 320 -3210
rect 260 -3275 275 -3245
rect 305 -3275 320 -3245
rect 260 -3305 320 -3275
rect 260 -3335 275 -3305
rect 305 -3335 320 -3305
rect 260 -3370 320 -3335
rect 260 -3400 275 -3370
rect 305 -3400 320 -3370
rect 260 -3440 320 -3400
rect 260 -3470 275 -3440
rect 305 -3470 320 -3440
rect 260 -3510 320 -3470
rect 260 -3540 275 -3510
rect 305 -3540 320 -3510
rect 260 -3580 320 -3540
rect 260 -3610 275 -3580
rect 305 -3610 320 -3580
rect 260 -3645 320 -3610
rect 260 -3675 275 -3645
rect 305 -3675 320 -3645
rect 260 -3705 320 -3675
rect 260 -3735 275 -3705
rect 305 -3735 320 -3705
rect 260 -3770 320 -3735
rect 260 -3800 275 -3770
rect 305 -3800 320 -3770
rect 260 -3840 320 -3800
rect 260 -3870 275 -3840
rect 305 -3870 320 -3840
rect 260 -3910 320 -3870
rect 260 -3940 275 -3910
rect 305 -3940 320 -3910
rect 260 -3980 320 -3940
rect 260 -4010 275 -3980
rect 305 -4010 320 -3980
rect 260 -4045 320 -4010
rect 260 -4075 275 -4045
rect 305 -4075 320 -4045
rect 260 -4105 320 -4075
rect 260 -4135 275 -4105
rect 305 -4135 320 -4105
rect 260 -4170 320 -4135
rect 260 -4200 275 -4170
rect 305 -4200 320 -4170
rect 260 -4240 320 -4200
rect 260 -4270 275 -4240
rect 305 -4270 320 -4240
rect 260 -4310 320 -4270
rect 260 -4340 275 -4310
rect 305 -4340 320 -4310
rect 260 -4380 320 -4340
rect 260 -4410 275 -4380
rect 305 -4410 320 -4380
rect 260 -4445 320 -4410
rect 260 -4475 275 -4445
rect 305 -4475 320 -4445
rect 260 -4490 320 -4475
rect 610 -1305 670 -1290
rect 610 -1335 625 -1305
rect 655 -1335 670 -1305
rect 610 -1370 670 -1335
rect 610 -1400 625 -1370
rect 655 -1400 670 -1370
rect 610 -1440 670 -1400
rect 610 -1470 625 -1440
rect 655 -1470 670 -1440
rect 610 -1510 670 -1470
rect 610 -1540 625 -1510
rect 655 -1540 670 -1510
rect 610 -1580 670 -1540
rect 610 -1610 625 -1580
rect 655 -1610 670 -1580
rect 610 -1645 670 -1610
rect 610 -1675 625 -1645
rect 655 -1675 670 -1645
rect 610 -1705 670 -1675
rect 610 -1735 625 -1705
rect 655 -1735 670 -1705
rect 610 -1770 670 -1735
rect 610 -1800 625 -1770
rect 655 -1800 670 -1770
rect 610 -1840 670 -1800
rect 610 -1870 625 -1840
rect 655 -1870 670 -1840
rect 610 -1910 670 -1870
rect 610 -1940 625 -1910
rect 655 -1940 670 -1910
rect 610 -1980 670 -1940
rect 610 -2010 625 -1980
rect 655 -2010 670 -1980
rect 610 -2045 670 -2010
rect 610 -2075 625 -2045
rect 655 -2075 670 -2045
rect 610 -2105 670 -2075
rect 610 -2135 625 -2105
rect 655 -2135 670 -2105
rect 610 -2170 670 -2135
rect 610 -2200 625 -2170
rect 655 -2200 670 -2170
rect 610 -2240 670 -2200
rect 610 -2270 625 -2240
rect 655 -2270 670 -2240
rect 610 -2310 670 -2270
rect 610 -2340 625 -2310
rect 655 -2340 670 -2310
rect 610 -2380 670 -2340
rect 610 -2410 625 -2380
rect 655 -2410 670 -2380
rect 610 -2445 670 -2410
rect 610 -2475 625 -2445
rect 655 -2475 670 -2445
rect 610 -2505 670 -2475
rect 610 -2535 625 -2505
rect 655 -2535 670 -2505
rect 610 -2570 670 -2535
rect 610 -2600 625 -2570
rect 655 -2600 670 -2570
rect 610 -2640 670 -2600
rect 610 -2670 625 -2640
rect 655 -2670 670 -2640
rect 610 -2710 670 -2670
rect 610 -2740 625 -2710
rect 655 -2740 670 -2710
rect 610 -2780 670 -2740
rect 610 -2810 625 -2780
rect 655 -2810 670 -2780
rect 610 -2845 670 -2810
rect 610 -2875 625 -2845
rect 655 -2875 670 -2845
rect 610 -2905 670 -2875
rect 610 -2935 625 -2905
rect 655 -2935 670 -2905
rect 610 -2970 670 -2935
rect 610 -3000 625 -2970
rect 655 -3000 670 -2970
rect 610 -3040 670 -3000
rect 610 -3070 625 -3040
rect 655 -3070 670 -3040
rect 610 -3110 670 -3070
rect 610 -3140 625 -3110
rect 655 -3140 670 -3110
rect 610 -3180 670 -3140
rect 610 -3210 625 -3180
rect 655 -3210 670 -3180
rect 610 -3245 670 -3210
rect 610 -3275 625 -3245
rect 655 -3275 670 -3245
rect 610 -3305 670 -3275
rect 610 -3335 625 -3305
rect 655 -3335 670 -3305
rect 610 -3370 670 -3335
rect 610 -3400 625 -3370
rect 655 -3400 670 -3370
rect 610 -3440 670 -3400
rect 610 -3470 625 -3440
rect 655 -3470 670 -3440
rect 610 -3510 670 -3470
rect 610 -3540 625 -3510
rect 655 -3540 670 -3510
rect 610 -3580 670 -3540
rect 610 -3610 625 -3580
rect 655 -3610 670 -3580
rect 610 -3645 670 -3610
rect 610 -3675 625 -3645
rect 655 -3675 670 -3645
rect 610 -3705 670 -3675
rect 610 -3735 625 -3705
rect 655 -3735 670 -3705
rect 610 -3770 670 -3735
rect 610 -3800 625 -3770
rect 655 -3800 670 -3770
rect 610 -3840 670 -3800
rect 610 -3870 625 -3840
rect 655 -3870 670 -3840
rect 610 -3910 670 -3870
rect 610 -3940 625 -3910
rect 655 -3940 670 -3910
rect 610 -3980 670 -3940
rect 610 -4010 625 -3980
rect 655 -4010 670 -3980
rect 610 -4045 670 -4010
rect 610 -4075 625 -4045
rect 655 -4075 670 -4045
rect 610 -4105 670 -4075
rect 610 -4135 625 -4105
rect 655 -4135 670 -4105
rect 610 -4170 670 -4135
rect 610 -4200 625 -4170
rect 655 -4200 670 -4170
rect 610 -4240 670 -4200
rect 610 -4270 625 -4240
rect 655 -4270 670 -4240
rect 610 -4310 670 -4270
rect 610 -4340 625 -4310
rect 655 -4340 670 -4310
rect 610 -4380 670 -4340
rect 610 -4410 625 -4380
rect 655 -4410 670 -4380
rect 610 -4445 670 -4410
rect 610 -4475 625 -4445
rect 655 -4475 670 -4445
rect 610 -4490 670 -4475
rect 960 -1305 1020 -1290
rect 960 -1335 975 -1305
rect 1005 -1335 1020 -1305
rect 960 -1370 1020 -1335
rect 960 -1400 975 -1370
rect 1005 -1400 1020 -1370
rect 960 -1440 1020 -1400
rect 960 -1470 975 -1440
rect 1005 -1470 1020 -1440
rect 960 -1510 1020 -1470
rect 960 -1540 975 -1510
rect 1005 -1540 1020 -1510
rect 960 -1580 1020 -1540
rect 960 -1610 975 -1580
rect 1005 -1610 1020 -1580
rect 960 -1645 1020 -1610
rect 960 -1675 975 -1645
rect 1005 -1675 1020 -1645
rect 960 -1705 1020 -1675
rect 960 -1735 975 -1705
rect 1005 -1735 1020 -1705
rect 960 -1770 1020 -1735
rect 960 -1800 975 -1770
rect 1005 -1800 1020 -1770
rect 960 -1840 1020 -1800
rect 960 -1870 975 -1840
rect 1005 -1870 1020 -1840
rect 960 -1910 1020 -1870
rect 960 -1940 975 -1910
rect 1005 -1940 1020 -1910
rect 960 -1980 1020 -1940
rect 960 -2010 975 -1980
rect 1005 -2010 1020 -1980
rect 960 -2045 1020 -2010
rect 960 -2075 975 -2045
rect 1005 -2075 1020 -2045
rect 960 -2105 1020 -2075
rect 960 -2135 975 -2105
rect 1005 -2135 1020 -2105
rect 960 -2170 1020 -2135
rect 960 -2200 975 -2170
rect 1005 -2200 1020 -2170
rect 960 -2240 1020 -2200
rect 960 -2270 975 -2240
rect 1005 -2270 1020 -2240
rect 960 -2310 1020 -2270
rect 960 -2340 975 -2310
rect 1005 -2340 1020 -2310
rect 960 -2380 1020 -2340
rect 960 -2410 975 -2380
rect 1005 -2410 1020 -2380
rect 960 -2445 1020 -2410
rect 960 -2475 975 -2445
rect 1005 -2475 1020 -2445
rect 960 -2505 1020 -2475
rect 960 -2535 975 -2505
rect 1005 -2535 1020 -2505
rect 960 -2570 1020 -2535
rect 960 -2600 975 -2570
rect 1005 -2600 1020 -2570
rect 960 -2640 1020 -2600
rect 960 -2670 975 -2640
rect 1005 -2670 1020 -2640
rect 960 -2710 1020 -2670
rect 960 -2740 975 -2710
rect 1005 -2740 1020 -2710
rect 960 -2780 1020 -2740
rect 960 -2810 975 -2780
rect 1005 -2810 1020 -2780
rect 960 -2845 1020 -2810
rect 960 -2875 975 -2845
rect 1005 -2875 1020 -2845
rect 960 -2905 1020 -2875
rect 960 -2935 975 -2905
rect 1005 -2935 1020 -2905
rect 960 -2970 1020 -2935
rect 960 -3000 975 -2970
rect 1005 -3000 1020 -2970
rect 960 -3040 1020 -3000
rect 960 -3070 975 -3040
rect 1005 -3070 1020 -3040
rect 960 -3110 1020 -3070
rect 960 -3140 975 -3110
rect 1005 -3140 1020 -3110
rect 960 -3180 1020 -3140
rect 960 -3210 975 -3180
rect 1005 -3210 1020 -3180
rect 960 -3245 1020 -3210
rect 960 -3275 975 -3245
rect 1005 -3275 1020 -3245
rect 960 -3305 1020 -3275
rect 960 -3335 975 -3305
rect 1005 -3335 1020 -3305
rect 960 -3370 1020 -3335
rect 960 -3400 975 -3370
rect 1005 -3400 1020 -3370
rect 960 -3440 1020 -3400
rect 960 -3470 975 -3440
rect 1005 -3470 1020 -3440
rect 960 -3510 1020 -3470
rect 960 -3540 975 -3510
rect 1005 -3540 1020 -3510
rect 960 -3580 1020 -3540
rect 960 -3610 975 -3580
rect 1005 -3610 1020 -3580
rect 960 -3645 1020 -3610
rect 960 -3675 975 -3645
rect 1005 -3675 1020 -3645
rect 960 -3705 1020 -3675
rect 960 -3735 975 -3705
rect 1005 -3735 1020 -3705
rect 960 -3770 1020 -3735
rect 960 -3800 975 -3770
rect 1005 -3800 1020 -3770
rect 960 -3840 1020 -3800
rect 960 -3870 975 -3840
rect 1005 -3870 1020 -3840
rect 960 -3910 1020 -3870
rect 960 -3940 975 -3910
rect 1005 -3940 1020 -3910
rect 960 -3980 1020 -3940
rect 960 -4010 975 -3980
rect 1005 -4010 1020 -3980
rect 960 -4045 1020 -4010
rect 960 -4075 975 -4045
rect 1005 -4075 1020 -4045
rect 960 -4105 1020 -4075
rect 960 -4135 975 -4105
rect 1005 -4135 1020 -4105
rect 960 -4170 1020 -4135
rect 960 -4200 975 -4170
rect 1005 -4200 1020 -4170
rect 960 -4240 1020 -4200
rect 960 -4270 975 -4240
rect 1005 -4270 1020 -4240
rect 960 -4310 1020 -4270
rect 960 -4340 975 -4310
rect 1005 -4340 1020 -4310
rect 960 -4380 1020 -4340
rect 960 -4410 975 -4380
rect 1005 -4410 1020 -4380
rect 960 -4445 1020 -4410
rect 960 -4475 975 -4445
rect 1005 -4475 1020 -4445
rect 960 -4490 1020 -4475
rect 1310 -1305 1370 -1290
rect 1310 -1335 1325 -1305
rect 1355 -1335 1370 -1305
rect 1310 -1370 1370 -1335
rect 1310 -1400 1325 -1370
rect 1355 -1400 1370 -1370
rect 1310 -1440 1370 -1400
rect 1310 -1470 1325 -1440
rect 1355 -1470 1370 -1440
rect 1310 -1510 1370 -1470
rect 1310 -1540 1325 -1510
rect 1355 -1540 1370 -1510
rect 1310 -1580 1370 -1540
rect 1310 -1610 1325 -1580
rect 1355 -1610 1370 -1580
rect 1310 -1645 1370 -1610
rect 1310 -1675 1325 -1645
rect 1355 -1675 1370 -1645
rect 1310 -1705 1370 -1675
rect 1310 -1735 1325 -1705
rect 1355 -1735 1370 -1705
rect 1310 -1770 1370 -1735
rect 1310 -1800 1325 -1770
rect 1355 -1800 1370 -1770
rect 1310 -1840 1370 -1800
rect 1310 -1870 1325 -1840
rect 1355 -1870 1370 -1840
rect 1310 -1910 1370 -1870
rect 1310 -1940 1325 -1910
rect 1355 -1940 1370 -1910
rect 1310 -1980 1370 -1940
rect 1310 -2010 1325 -1980
rect 1355 -2010 1370 -1980
rect 1310 -2045 1370 -2010
rect 1310 -2075 1325 -2045
rect 1355 -2075 1370 -2045
rect 1310 -2105 1370 -2075
rect 1310 -2135 1325 -2105
rect 1355 -2135 1370 -2105
rect 1310 -2170 1370 -2135
rect 1310 -2200 1325 -2170
rect 1355 -2200 1370 -2170
rect 1310 -2240 1370 -2200
rect 1310 -2270 1325 -2240
rect 1355 -2270 1370 -2240
rect 1310 -2310 1370 -2270
rect 1310 -2340 1325 -2310
rect 1355 -2340 1370 -2310
rect 1310 -2380 1370 -2340
rect 1310 -2410 1325 -2380
rect 1355 -2410 1370 -2380
rect 1310 -2445 1370 -2410
rect 1310 -2475 1325 -2445
rect 1355 -2475 1370 -2445
rect 1310 -2505 1370 -2475
rect 1310 -2535 1325 -2505
rect 1355 -2535 1370 -2505
rect 1310 -2570 1370 -2535
rect 1310 -2600 1325 -2570
rect 1355 -2600 1370 -2570
rect 1310 -2640 1370 -2600
rect 1310 -2670 1325 -2640
rect 1355 -2670 1370 -2640
rect 1310 -2710 1370 -2670
rect 1310 -2740 1325 -2710
rect 1355 -2740 1370 -2710
rect 1310 -2780 1370 -2740
rect 1310 -2810 1325 -2780
rect 1355 -2810 1370 -2780
rect 1310 -2845 1370 -2810
rect 1310 -2875 1325 -2845
rect 1355 -2875 1370 -2845
rect 1310 -2905 1370 -2875
rect 1310 -2935 1325 -2905
rect 1355 -2935 1370 -2905
rect 1310 -2970 1370 -2935
rect 1310 -3000 1325 -2970
rect 1355 -3000 1370 -2970
rect 1310 -3040 1370 -3000
rect 1310 -3070 1325 -3040
rect 1355 -3070 1370 -3040
rect 1310 -3110 1370 -3070
rect 1310 -3140 1325 -3110
rect 1355 -3140 1370 -3110
rect 1310 -3180 1370 -3140
rect 1310 -3210 1325 -3180
rect 1355 -3210 1370 -3180
rect 1310 -3245 1370 -3210
rect 1310 -3275 1325 -3245
rect 1355 -3275 1370 -3245
rect 1310 -3305 1370 -3275
rect 1310 -3335 1325 -3305
rect 1355 -3335 1370 -3305
rect 1310 -3370 1370 -3335
rect 1310 -3400 1325 -3370
rect 1355 -3400 1370 -3370
rect 1310 -3440 1370 -3400
rect 1310 -3470 1325 -3440
rect 1355 -3470 1370 -3440
rect 1310 -3510 1370 -3470
rect 1310 -3540 1325 -3510
rect 1355 -3540 1370 -3510
rect 1310 -3580 1370 -3540
rect 1310 -3610 1325 -3580
rect 1355 -3610 1370 -3580
rect 1310 -3645 1370 -3610
rect 1310 -3675 1325 -3645
rect 1355 -3675 1370 -3645
rect 1310 -3705 1370 -3675
rect 1310 -3735 1325 -3705
rect 1355 -3735 1370 -3705
rect 1310 -3770 1370 -3735
rect 1310 -3800 1325 -3770
rect 1355 -3800 1370 -3770
rect 1310 -3840 1370 -3800
rect 1310 -3870 1325 -3840
rect 1355 -3870 1370 -3840
rect 1310 -3910 1370 -3870
rect 1310 -3940 1325 -3910
rect 1355 -3940 1370 -3910
rect 1310 -3980 1370 -3940
rect 1310 -4010 1325 -3980
rect 1355 -4010 1370 -3980
rect 1310 -4045 1370 -4010
rect 1310 -4075 1325 -4045
rect 1355 -4075 1370 -4045
rect 1310 -4105 1370 -4075
rect 1310 -4135 1325 -4105
rect 1355 -4135 1370 -4105
rect 1310 -4170 1370 -4135
rect 1310 -4200 1325 -4170
rect 1355 -4200 1370 -4170
rect 1310 -4240 1370 -4200
rect 1310 -4270 1325 -4240
rect 1355 -4270 1370 -4240
rect 1310 -4310 1370 -4270
rect 1310 -4340 1325 -4310
rect 1355 -4340 1370 -4310
rect 1310 -4380 1370 -4340
rect 1310 -4410 1325 -4380
rect 1355 -4410 1370 -4380
rect 1310 -4445 1370 -4410
rect 1310 -4475 1325 -4445
rect 1355 -4475 1370 -4445
rect 1310 -4490 1370 -4475
rect 1660 -1305 1720 -1290
rect 1660 -1335 1675 -1305
rect 1705 -1335 1720 -1305
rect 1660 -1370 1720 -1335
rect 1660 -1400 1675 -1370
rect 1705 -1400 1720 -1370
rect 1660 -1440 1720 -1400
rect 1660 -1470 1675 -1440
rect 1705 -1470 1720 -1440
rect 1660 -1510 1720 -1470
rect 1660 -1540 1675 -1510
rect 1705 -1540 1720 -1510
rect 1660 -1580 1720 -1540
rect 1660 -1610 1675 -1580
rect 1705 -1610 1720 -1580
rect 1660 -1645 1720 -1610
rect 1660 -1675 1675 -1645
rect 1705 -1675 1720 -1645
rect 1660 -1705 1720 -1675
rect 1660 -1735 1675 -1705
rect 1705 -1735 1720 -1705
rect 1660 -1770 1720 -1735
rect 1660 -1800 1675 -1770
rect 1705 -1800 1720 -1770
rect 1660 -1840 1720 -1800
rect 1660 -1870 1675 -1840
rect 1705 -1870 1720 -1840
rect 1660 -1910 1720 -1870
rect 1660 -1940 1675 -1910
rect 1705 -1940 1720 -1910
rect 1660 -1980 1720 -1940
rect 1660 -2010 1675 -1980
rect 1705 -2010 1720 -1980
rect 1660 -2045 1720 -2010
rect 1660 -2075 1675 -2045
rect 1705 -2075 1720 -2045
rect 1660 -2105 1720 -2075
rect 1660 -2135 1675 -2105
rect 1705 -2135 1720 -2105
rect 1660 -2170 1720 -2135
rect 1660 -2200 1675 -2170
rect 1705 -2200 1720 -2170
rect 1660 -2240 1720 -2200
rect 1660 -2270 1675 -2240
rect 1705 -2270 1720 -2240
rect 1660 -2310 1720 -2270
rect 1660 -2340 1675 -2310
rect 1705 -2340 1720 -2310
rect 1660 -2380 1720 -2340
rect 1660 -2410 1675 -2380
rect 1705 -2410 1720 -2380
rect 1660 -2445 1720 -2410
rect 1660 -2475 1675 -2445
rect 1705 -2475 1720 -2445
rect 1660 -2505 1720 -2475
rect 1660 -2535 1675 -2505
rect 1705 -2535 1720 -2505
rect 1660 -2570 1720 -2535
rect 1660 -2600 1675 -2570
rect 1705 -2600 1720 -2570
rect 1660 -2640 1720 -2600
rect 1660 -2670 1675 -2640
rect 1705 -2670 1720 -2640
rect 1660 -2710 1720 -2670
rect 1660 -2740 1675 -2710
rect 1705 -2740 1720 -2710
rect 1660 -2780 1720 -2740
rect 1660 -2810 1675 -2780
rect 1705 -2810 1720 -2780
rect 1660 -2845 1720 -2810
rect 1660 -2875 1675 -2845
rect 1705 -2875 1720 -2845
rect 1660 -2905 1720 -2875
rect 1660 -2935 1675 -2905
rect 1705 -2935 1720 -2905
rect 1660 -2970 1720 -2935
rect 1660 -3000 1675 -2970
rect 1705 -3000 1720 -2970
rect 1660 -3040 1720 -3000
rect 1660 -3070 1675 -3040
rect 1705 -3070 1720 -3040
rect 1660 -3110 1720 -3070
rect 1660 -3140 1675 -3110
rect 1705 -3140 1720 -3110
rect 1660 -3180 1720 -3140
rect 1660 -3210 1675 -3180
rect 1705 -3210 1720 -3180
rect 1660 -3245 1720 -3210
rect 1660 -3275 1675 -3245
rect 1705 -3275 1720 -3245
rect 1660 -3305 1720 -3275
rect 1660 -3335 1675 -3305
rect 1705 -3335 1720 -3305
rect 1660 -3370 1720 -3335
rect 1660 -3400 1675 -3370
rect 1705 -3400 1720 -3370
rect 1660 -3440 1720 -3400
rect 1660 -3470 1675 -3440
rect 1705 -3470 1720 -3440
rect 1660 -3510 1720 -3470
rect 1660 -3540 1675 -3510
rect 1705 -3540 1720 -3510
rect 1660 -3580 1720 -3540
rect 1660 -3610 1675 -3580
rect 1705 -3610 1720 -3580
rect 1660 -3645 1720 -3610
rect 1660 -3675 1675 -3645
rect 1705 -3675 1720 -3645
rect 1660 -3705 1720 -3675
rect 1660 -3735 1675 -3705
rect 1705 -3735 1720 -3705
rect 1660 -3770 1720 -3735
rect 1660 -3800 1675 -3770
rect 1705 -3800 1720 -3770
rect 1660 -3840 1720 -3800
rect 1660 -3870 1675 -3840
rect 1705 -3870 1720 -3840
rect 1660 -3910 1720 -3870
rect 1660 -3940 1675 -3910
rect 1705 -3940 1720 -3910
rect 1660 -3980 1720 -3940
rect 1660 -4010 1675 -3980
rect 1705 -4010 1720 -3980
rect 1660 -4045 1720 -4010
rect 1660 -4075 1675 -4045
rect 1705 -4075 1720 -4045
rect 1660 -4105 1720 -4075
rect 1660 -4135 1675 -4105
rect 1705 -4135 1720 -4105
rect 1660 -4170 1720 -4135
rect 1660 -4200 1675 -4170
rect 1705 -4200 1720 -4170
rect 1660 -4240 1720 -4200
rect 1660 -4270 1675 -4240
rect 1705 -4270 1720 -4240
rect 1660 -4310 1720 -4270
rect 1660 -4340 1675 -4310
rect 1705 -4340 1720 -4310
rect 1660 -4380 1720 -4340
rect 1660 -4410 1675 -4380
rect 1705 -4410 1720 -4380
rect 1660 -4445 1720 -4410
rect 1660 -4475 1675 -4445
rect 1705 -4475 1720 -4445
rect 1660 -4490 1720 -4475
rect 2010 -1305 2070 -1290
rect 2010 -1335 2025 -1305
rect 2055 -1335 2070 -1305
rect 2010 -1370 2070 -1335
rect 2010 -1400 2025 -1370
rect 2055 -1400 2070 -1370
rect 2010 -1440 2070 -1400
rect 2010 -1470 2025 -1440
rect 2055 -1470 2070 -1440
rect 2010 -1510 2070 -1470
rect 2010 -1540 2025 -1510
rect 2055 -1540 2070 -1510
rect 2010 -1580 2070 -1540
rect 2010 -1610 2025 -1580
rect 2055 -1610 2070 -1580
rect 2010 -1645 2070 -1610
rect 2010 -1675 2025 -1645
rect 2055 -1675 2070 -1645
rect 2010 -1705 2070 -1675
rect 2010 -1735 2025 -1705
rect 2055 -1735 2070 -1705
rect 2010 -1770 2070 -1735
rect 2010 -1800 2025 -1770
rect 2055 -1800 2070 -1770
rect 2010 -1840 2070 -1800
rect 2010 -1870 2025 -1840
rect 2055 -1870 2070 -1840
rect 2010 -1910 2070 -1870
rect 2010 -1940 2025 -1910
rect 2055 -1940 2070 -1910
rect 2010 -1980 2070 -1940
rect 2010 -2010 2025 -1980
rect 2055 -2010 2070 -1980
rect 2010 -2045 2070 -2010
rect 2010 -2075 2025 -2045
rect 2055 -2075 2070 -2045
rect 2010 -2105 2070 -2075
rect 2010 -2135 2025 -2105
rect 2055 -2135 2070 -2105
rect 2010 -2170 2070 -2135
rect 2010 -2200 2025 -2170
rect 2055 -2200 2070 -2170
rect 2010 -2240 2070 -2200
rect 2010 -2270 2025 -2240
rect 2055 -2270 2070 -2240
rect 2010 -2310 2070 -2270
rect 2010 -2340 2025 -2310
rect 2055 -2340 2070 -2310
rect 2010 -2380 2070 -2340
rect 2010 -2410 2025 -2380
rect 2055 -2410 2070 -2380
rect 2010 -2445 2070 -2410
rect 2010 -2475 2025 -2445
rect 2055 -2475 2070 -2445
rect 2010 -2505 2070 -2475
rect 2010 -2535 2025 -2505
rect 2055 -2535 2070 -2505
rect 2010 -2570 2070 -2535
rect 2010 -2600 2025 -2570
rect 2055 -2600 2070 -2570
rect 2010 -2640 2070 -2600
rect 2010 -2670 2025 -2640
rect 2055 -2670 2070 -2640
rect 2010 -2710 2070 -2670
rect 2010 -2740 2025 -2710
rect 2055 -2740 2070 -2710
rect 2010 -2780 2070 -2740
rect 2010 -2810 2025 -2780
rect 2055 -2810 2070 -2780
rect 2010 -2845 2070 -2810
rect 2010 -2875 2025 -2845
rect 2055 -2875 2070 -2845
rect 2010 -2905 2070 -2875
rect 2010 -2935 2025 -2905
rect 2055 -2935 2070 -2905
rect 2010 -2970 2070 -2935
rect 2010 -3000 2025 -2970
rect 2055 -3000 2070 -2970
rect 2010 -3040 2070 -3000
rect 2010 -3070 2025 -3040
rect 2055 -3070 2070 -3040
rect 2010 -3110 2070 -3070
rect 2010 -3140 2025 -3110
rect 2055 -3140 2070 -3110
rect 2010 -3180 2070 -3140
rect 2010 -3210 2025 -3180
rect 2055 -3210 2070 -3180
rect 2010 -3245 2070 -3210
rect 2010 -3275 2025 -3245
rect 2055 -3275 2070 -3245
rect 2010 -3305 2070 -3275
rect 2010 -3335 2025 -3305
rect 2055 -3335 2070 -3305
rect 2010 -3370 2070 -3335
rect 2010 -3400 2025 -3370
rect 2055 -3400 2070 -3370
rect 2010 -3440 2070 -3400
rect 2010 -3470 2025 -3440
rect 2055 -3470 2070 -3440
rect 2010 -3510 2070 -3470
rect 2010 -3540 2025 -3510
rect 2055 -3540 2070 -3510
rect 2010 -3580 2070 -3540
rect 2010 -3610 2025 -3580
rect 2055 -3610 2070 -3580
rect 2010 -3645 2070 -3610
rect 2010 -3675 2025 -3645
rect 2055 -3675 2070 -3645
rect 2010 -3705 2070 -3675
rect 2010 -3735 2025 -3705
rect 2055 -3735 2070 -3705
rect 2010 -3770 2070 -3735
rect 2010 -3800 2025 -3770
rect 2055 -3800 2070 -3770
rect 2010 -3840 2070 -3800
rect 2010 -3870 2025 -3840
rect 2055 -3870 2070 -3840
rect 2010 -3910 2070 -3870
rect 2010 -3940 2025 -3910
rect 2055 -3940 2070 -3910
rect 2010 -3980 2070 -3940
rect 2010 -4010 2025 -3980
rect 2055 -4010 2070 -3980
rect 2010 -4045 2070 -4010
rect 2010 -4075 2025 -4045
rect 2055 -4075 2070 -4045
rect 2010 -4105 2070 -4075
rect 2010 -4135 2025 -4105
rect 2055 -4135 2070 -4105
rect 2010 -4170 2070 -4135
rect 2010 -4200 2025 -4170
rect 2055 -4200 2070 -4170
rect 2010 -4240 2070 -4200
rect 2010 -4270 2025 -4240
rect 2055 -4270 2070 -4240
rect 2010 -4310 2070 -4270
rect 2010 -4340 2025 -4310
rect 2055 -4340 2070 -4310
rect 2010 -4380 2070 -4340
rect 2010 -4410 2025 -4380
rect 2055 -4410 2070 -4380
rect 2010 -4445 2070 -4410
rect 2010 -4475 2025 -4445
rect 2055 -4475 2070 -4445
rect 2010 -4490 2070 -4475
rect 2360 -1305 2420 -1290
rect 2360 -1335 2375 -1305
rect 2405 -1335 2420 -1305
rect 2360 -1370 2420 -1335
rect 2360 -1400 2375 -1370
rect 2405 -1400 2420 -1370
rect 2360 -1440 2420 -1400
rect 2360 -1470 2375 -1440
rect 2405 -1470 2420 -1440
rect 2360 -1510 2420 -1470
rect 2360 -1540 2375 -1510
rect 2405 -1540 2420 -1510
rect 2360 -1580 2420 -1540
rect 2360 -1610 2375 -1580
rect 2405 -1610 2420 -1580
rect 2360 -1645 2420 -1610
rect 2360 -1675 2375 -1645
rect 2405 -1675 2420 -1645
rect 2360 -1705 2420 -1675
rect 2360 -1735 2375 -1705
rect 2405 -1735 2420 -1705
rect 2360 -1770 2420 -1735
rect 2360 -1800 2375 -1770
rect 2405 -1800 2420 -1770
rect 2360 -1840 2420 -1800
rect 2360 -1870 2375 -1840
rect 2405 -1870 2420 -1840
rect 2360 -1910 2420 -1870
rect 2360 -1940 2375 -1910
rect 2405 -1940 2420 -1910
rect 2360 -1980 2420 -1940
rect 2360 -2010 2375 -1980
rect 2405 -2010 2420 -1980
rect 2360 -2045 2420 -2010
rect 2360 -2075 2375 -2045
rect 2405 -2075 2420 -2045
rect 2360 -2105 2420 -2075
rect 2360 -2135 2375 -2105
rect 2405 -2135 2420 -2105
rect 2360 -2170 2420 -2135
rect 2360 -2200 2375 -2170
rect 2405 -2200 2420 -2170
rect 2360 -2240 2420 -2200
rect 2360 -2270 2375 -2240
rect 2405 -2270 2420 -2240
rect 2360 -2310 2420 -2270
rect 2360 -2340 2375 -2310
rect 2405 -2340 2420 -2310
rect 2360 -2380 2420 -2340
rect 2360 -2410 2375 -2380
rect 2405 -2410 2420 -2380
rect 2360 -2445 2420 -2410
rect 2360 -2475 2375 -2445
rect 2405 -2475 2420 -2445
rect 2360 -2505 2420 -2475
rect 2360 -2535 2375 -2505
rect 2405 -2535 2420 -2505
rect 2360 -2570 2420 -2535
rect 2360 -2600 2375 -2570
rect 2405 -2600 2420 -2570
rect 2360 -2640 2420 -2600
rect 2360 -2670 2375 -2640
rect 2405 -2670 2420 -2640
rect 2360 -2710 2420 -2670
rect 2360 -2740 2375 -2710
rect 2405 -2740 2420 -2710
rect 2360 -2780 2420 -2740
rect 2360 -2810 2375 -2780
rect 2405 -2810 2420 -2780
rect 2360 -2845 2420 -2810
rect 2360 -2875 2375 -2845
rect 2405 -2875 2420 -2845
rect 2360 -2905 2420 -2875
rect 2360 -2935 2375 -2905
rect 2405 -2935 2420 -2905
rect 2360 -2970 2420 -2935
rect 2360 -3000 2375 -2970
rect 2405 -3000 2420 -2970
rect 2360 -3040 2420 -3000
rect 2360 -3070 2375 -3040
rect 2405 -3070 2420 -3040
rect 2360 -3110 2420 -3070
rect 2360 -3140 2375 -3110
rect 2405 -3140 2420 -3110
rect 2360 -3180 2420 -3140
rect 2360 -3210 2375 -3180
rect 2405 -3210 2420 -3180
rect 2360 -3245 2420 -3210
rect 2360 -3275 2375 -3245
rect 2405 -3275 2420 -3245
rect 2360 -3305 2420 -3275
rect 2360 -3335 2375 -3305
rect 2405 -3335 2420 -3305
rect 2360 -3370 2420 -3335
rect 2360 -3400 2375 -3370
rect 2405 -3400 2420 -3370
rect 2360 -3440 2420 -3400
rect 2360 -3470 2375 -3440
rect 2405 -3470 2420 -3440
rect 2360 -3510 2420 -3470
rect 2360 -3540 2375 -3510
rect 2405 -3540 2420 -3510
rect 2360 -3580 2420 -3540
rect 2360 -3610 2375 -3580
rect 2405 -3610 2420 -3580
rect 2360 -3645 2420 -3610
rect 2360 -3675 2375 -3645
rect 2405 -3675 2420 -3645
rect 2360 -3705 2420 -3675
rect 2360 -3735 2375 -3705
rect 2405 -3735 2420 -3705
rect 2360 -3770 2420 -3735
rect 2360 -3800 2375 -3770
rect 2405 -3800 2420 -3770
rect 2360 -3840 2420 -3800
rect 2360 -3870 2375 -3840
rect 2405 -3870 2420 -3840
rect 2360 -3910 2420 -3870
rect 2360 -3940 2375 -3910
rect 2405 -3940 2420 -3910
rect 2360 -3980 2420 -3940
rect 2360 -4010 2375 -3980
rect 2405 -4010 2420 -3980
rect 2360 -4045 2420 -4010
rect 2360 -4075 2375 -4045
rect 2405 -4075 2420 -4045
rect 2360 -4105 2420 -4075
rect 2360 -4135 2375 -4105
rect 2405 -4135 2420 -4105
rect 2360 -4170 2420 -4135
rect 2360 -4200 2375 -4170
rect 2405 -4200 2420 -4170
rect 2360 -4240 2420 -4200
rect 2360 -4270 2375 -4240
rect 2405 -4270 2420 -4240
rect 2360 -4310 2420 -4270
rect 2360 -4340 2375 -4310
rect 2405 -4340 2420 -4310
rect 2360 -4380 2420 -4340
rect 2360 -4410 2375 -4380
rect 2405 -4410 2420 -4380
rect 2360 -4445 2420 -4410
rect 2360 -4475 2375 -4445
rect 2405 -4475 2420 -4445
rect 2360 -4490 2420 -4475
rect 2710 -1305 2770 -1290
rect 2710 -1335 2725 -1305
rect 2755 -1335 2770 -1305
rect 2710 -1370 2770 -1335
rect 2710 -1400 2725 -1370
rect 2755 -1400 2770 -1370
rect 2710 -1440 2770 -1400
rect 2710 -1470 2725 -1440
rect 2755 -1470 2770 -1440
rect 2710 -1510 2770 -1470
rect 2710 -1540 2725 -1510
rect 2755 -1540 2770 -1510
rect 2710 -1580 2770 -1540
rect 2710 -1610 2725 -1580
rect 2755 -1610 2770 -1580
rect 2710 -1645 2770 -1610
rect 2710 -1675 2725 -1645
rect 2755 -1675 2770 -1645
rect 2710 -1705 2770 -1675
rect 2710 -1735 2725 -1705
rect 2755 -1735 2770 -1705
rect 2710 -1770 2770 -1735
rect 2710 -1800 2725 -1770
rect 2755 -1800 2770 -1770
rect 2710 -1840 2770 -1800
rect 2710 -1870 2725 -1840
rect 2755 -1870 2770 -1840
rect 2710 -1910 2770 -1870
rect 2710 -1940 2725 -1910
rect 2755 -1940 2770 -1910
rect 2710 -1980 2770 -1940
rect 2710 -2010 2725 -1980
rect 2755 -2010 2770 -1980
rect 2710 -2045 2770 -2010
rect 2710 -2075 2725 -2045
rect 2755 -2075 2770 -2045
rect 2710 -2105 2770 -2075
rect 2710 -2135 2725 -2105
rect 2755 -2135 2770 -2105
rect 2710 -2170 2770 -2135
rect 2710 -2200 2725 -2170
rect 2755 -2200 2770 -2170
rect 2710 -2240 2770 -2200
rect 2710 -2270 2725 -2240
rect 2755 -2270 2770 -2240
rect 2710 -2310 2770 -2270
rect 2710 -2340 2725 -2310
rect 2755 -2340 2770 -2310
rect 2710 -2380 2770 -2340
rect 2710 -2410 2725 -2380
rect 2755 -2410 2770 -2380
rect 2710 -2445 2770 -2410
rect 2710 -2475 2725 -2445
rect 2755 -2475 2770 -2445
rect 2710 -2505 2770 -2475
rect 2710 -2535 2725 -2505
rect 2755 -2535 2770 -2505
rect 2710 -2570 2770 -2535
rect 2710 -2600 2725 -2570
rect 2755 -2600 2770 -2570
rect 2710 -2640 2770 -2600
rect 2710 -2670 2725 -2640
rect 2755 -2670 2770 -2640
rect 2710 -2710 2770 -2670
rect 2710 -2740 2725 -2710
rect 2755 -2740 2770 -2710
rect 2710 -2780 2770 -2740
rect 2710 -2810 2725 -2780
rect 2755 -2810 2770 -2780
rect 2710 -2845 2770 -2810
rect 2710 -2875 2725 -2845
rect 2755 -2875 2770 -2845
rect 2710 -2905 2770 -2875
rect 2710 -2935 2725 -2905
rect 2755 -2935 2770 -2905
rect 2710 -2970 2770 -2935
rect 2710 -3000 2725 -2970
rect 2755 -3000 2770 -2970
rect 2710 -3040 2770 -3000
rect 2710 -3070 2725 -3040
rect 2755 -3070 2770 -3040
rect 2710 -3110 2770 -3070
rect 2710 -3140 2725 -3110
rect 2755 -3140 2770 -3110
rect 2710 -3180 2770 -3140
rect 2710 -3210 2725 -3180
rect 2755 -3210 2770 -3180
rect 2710 -3245 2770 -3210
rect 2710 -3275 2725 -3245
rect 2755 -3275 2770 -3245
rect 2710 -3305 2770 -3275
rect 2710 -3335 2725 -3305
rect 2755 -3335 2770 -3305
rect 2710 -3370 2770 -3335
rect 2710 -3400 2725 -3370
rect 2755 -3400 2770 -3370
rect 2710 -3440 2770 -3400
rect 2710 -3470 2725 -3440
rect 2755 -3470 2770 -3440
rect 2710 -3510 2770 -3470
rect 2710 -3540 2725 -3510
rect 2755 -3540 2770 -3510
rect 2710 -3580 2770 -3540
rect 2710 -3610 2725 -3580
rect 2755 -3610 2770 -3580
rect 2710 -3645 2770 -3610
rect 2710 -3675 2725 -3645
rect 2755 -3675 2770 -3645
rect 2710 -3705 2770 -3675
rect 2710 -3735 2725 -3705
rect 2755 -3735 2770 -3705
rect 2710 -3770 2770 -3735
rect 2710 -3800 2725 -3770
rect 2755 -3800 2770 -3770
rect 2710 -3840 2770 -3800
rect 2710 -3870 2725 -3840
rect 2755 -3870 2770 -3840
rect 2710 -3910 2770 -3870
rect 2710 -3940 2725 -3910
rect 2755 -3940 2770 -3910
rect 2710 -3980 2770 -3940
rect 2710 -4010 2725 -3980
rect 2755 -4010 2770 -3980
rect 2710 -4045 2770 -4010
rect 2710 -4075 2725 -4045
rect 2755 -4075 2770 -4045
rect 2710 -4105 2770 -4075
rect 2710 -4135 2725 -4105
rect 2755 -4135 2770 -4105
rect 2710 -4170 2770 -4135
rect 2710 -4200 2725 -4170
rect 2755 -4200 2770 -4170
rect 2710 -4240 2770 -4200
rect 2710 -4270 2725 -4240
rect 2755 -4270 2770 -4240
rect 2710 -4310 2770 -4270
rect 2710 -4340 2725 -4310
rect 2755 -4340 2770 -4310
rect 2710 -4380 2770 -4340
rect 2710 -4410 2725 -4380
rect 2755 -4410 2770 -4380
rect 2710 -4445 2770 -4410
rect 2710 -4475 2725 -4445
rect 2755 -4475 2770 -4445
rect 2710 -4490 2770 -4475
rect 3060 -1305 3120 -1290
rect 3060 -1335 3075 -1305
rect 3105 -1335 3120 -1305
rect 3060 -1370 3120 -1335
rect 3060 -1400 3075 -1370
rect 3105 -1400 3120 -1370
rect 3060 -1440 3120 -1400
rect 3060 -1470 3075 -1440
rect 3105 -1470 3120 -1440
rect 3060 -1510 3120 -1470
rect 3060 -1540 3075 -1510
rect 3105 -1540 3120 -1510
rect 3060 -1580 3120 -1540
rect 3060 -1610 3075 -1580
rect 3105 -1610 3120 -1580
rect 3060 -1645 3120 -1610
rect 3060 -1675 3075 -1645
rect 3105 -1675 3120 -1645
rect 3060 -1705 3120 -1675
rect 3060 -1735 3075 -1705
rect 3105 -1735 3120 -1705
rect 3060 -1770 3120 -1735
rect 3060 -1800 3075 -1770
rect 3105 -1800 3120 -1770
rect 3060 -1840 3120 -1800
rect 3060 -1870 3075 -1840
rect 3105 -1870 3120 -1840
rect 3060 -1910 3120 -1870
rect 3060 -1940 3075 -1910
rect 3105 -1940 3120 -1910
rect 3060 -1980 3120 -1940
rect 3060 -2010 3075 -1980
rect 3105 -2010 3120 -1980
rect 3060 -2045 3120 -2010
rect 3060 -2075 3075 -2045
rect 3105 -2075 3120 -2045
rect 3060 -2105 3120 -2075
rect 3060 -2135 3075 -2105
rect 3105 -2135 3120 -2105
rect 3060 -2170 3120 -2135
rect 3060 -2200 3075 -2170
rect 3105 -2200 3120 -2170
rect 3060 -2240 3120 -2200
rect 3060 -2270 3075 -2240
rect 3105 -2270 3120 -2240
rect 3060 -2310 3120 -2270
rect 3060 -2340 3075 -2310
rect 3105 -2340 3120 -2310
rect 3060 -2380 3120 -2340
rect 3060 -2410 3075 -2380
rect 3105 -2410 3120 -2380
rect 3060 -2445 3120 -2410
rect 3060 -2475 3075 -2445
rect 3105 -2475 3120 -2445
rect 3060 -2505 3120 -2475
rect 3060 -2535 3075 -2505
rect 3105 -2535 3120 -2505
rect 3060 -2570 3120 -2535
rect 3060 -2600 3075 -2570
rect 3105 -2600 3120 -2570
rect 3060 -2640 3120 -2600
rect 3060 -2670 3075 -2640
rect 3105 -2670 3120 -2640
rect 3060 -2710 3120 -2670
rect 3060 -2740 3075 -2710
rect 3105 -2740 3120 -2710
rect 3060 -2780 3120 -2740
rect 3060 -2810 3075 -2780
rect 3105 -2810 3120 -2780
rect 3060 -2845 3120 -2810
rect 3060 -2875 3075 -2845
rect 3105 -2875 3120 -2845
rect 3060 -2905 3120 -2875
rect 3060 -2935 3075 -2905
rect 3105 -2935 3120 -2905
rect 3060 -2970 3120 -2935
rect 3060 -3000 3075 -2970
rect 3105 -3000 3120 -2970
rect 3060 -3040 3120 -3000
rect 3060 -3070 3075 -3040
rect 3105 -3070 3120 -3040
rect 3060 -3110 3120 -3070
rect 3060 -3140 3075 -3110
rect 3105 -3140 3120 -3110
rect 3060 -3180 3120 -3140
rect 3060 -3210 3075 -3180
rect 3105 -3210 3120 -3180
rect 3060 -3245 3120 -3210
rect 3060 -3275 3075 -3245
rect 3105 -3275 3120 -3245
rect 3060 -3305 3120 -3275
rect 3060 -3335 3075 -3305
rect 3105 -3335 3120 -3305
rect 3060 -3370 3120 -3335
rect 3060 -3400 3075 -3370
rect 3105 -3400 3120 -3370
rect 3060 -3440 3120 -3400
rect 3060 -3470 3075 -3440
rect 3105 -3470 3120 -3440
rect 3060 -3510 3120 -3470
rect 3060 -3540 3075 -3510
rect 3105 -3540 3120 -3510
rect 3060 -3580 3120 -3540
rect 3060 -3610 3075 -3580
rect 3105 -3610 3120 -3580
rect 3060 -3645 3120 -3610
rect 3060 -3675 3075 -3645
rect 3105 -3675 3120 -3645
rect 3060 -3705 3120 -3675
rect 3060 -3735 3075 -3705
rect 3105 -3735 3120 -3705
rect 3060 -3770 3120 -3735
rect 3060 -3800 3075 -3770
rect 3105 -3800 3120 -3770
rect 3060 -3840 3120 -3800
rect 3060 -3870 3075 -3840
rect 3105 -3870 3120 -3840
rect 3060 -3910 3120 -3870
rect 3060 -3940 3075 -3910
rect 3105 -3940 3120 -3910
rect 3060 -3980 3120 -3940
rect 3060 -4010 3075 -3980
rect 3105 -4010 3120 -3980
rect 3060 -4045 3120 -4010
rect 3060 -4075 3075 -4045
rect 3105 -4075 3120 -4045
rect 3060 -4105 3120 -4075
rect 3060 -4135 3075 -4105
rect 3105 -4135 3120 -4105
rect 3060 -4170 3120 -4135
rect 3060 -4200 3075 -4170
rect 3105 -4200 3120 -4170
rect 3060 -4240 3120 -4200
rect 3060 -4270 3075 -4240
rect 3105 -4270 3120 -4240
rect 3060 -4310 3120 -4270
rect 3060 -4340 3075 -4310
rect 3105 -4340 3120 -4310
rect 3060 -4380 3120 -4340
rect 3060 -4410 3075 -4380
rect 3105 -4410 3120 -4380
rect 3060 -4445 3120 -4410
rect 3060 -4475 3075 -4445
rect 3105 -4475 3120 -4445
rect 3060 -4490 3120 -4475
rect 3410 -1305 3470 -1290
rect 3410 -1335 3425 -1305
rect 3455 -1335 3470 -1305
rect 3410 -1370 3470 -1335
rect 3410 -1400 3425 -1370
rect 3455 -1400 3470 -1370
rect 3410 -1440 3470 -1400
rect 3410 -1470 3425 -1440
rect 3455 -1470 3470 -1440
rect 3410 -1510 3470 -1470
rect 3410 -1540 3425 -1510
rect 3455 -1540 3470 -1510
rect 3410 -1580 3470 -1540
rect 3410 -1610 3425 -1580
rect 3455 -1610 3470 -1580
rect 3410 -1645 3470 -1610
rect 3410 -1675 3425 -1645
rect 3455 -1675 3470 -1645
rect 3410 -1705 3470 -1675
rect 3410 -1735 3425 -1705
rect 3455 -1735 3470 -1705
rect 3410 -1770 3470 -1735
rect 3410 -1800 3425 -1770
rect 3455 -1800 3470 -1770
rect 3410 -1840 3470 -1800
rect 3410 -1870 3425 -1840
rect 3455 -1870 3470 -1840
rect 3410 -1910 3470 -1870
rect 3410 -1940 3425 -1910
rect 3455 -1940 3470 -1910
rect 3410 -1980 3470 -1940
rect 3410 -2010 3425 -1980
rect 3455 -2010 3470 -1980
rect 3410 -2045 3470 -2010
rect 3410 -2075 3425 -2045
rect 3455 -2075 3470 -2045
rect 3410 -2105 3470 -2075
rect 3410 -2135 3425 -2105
rect 3455 -2135 3470 -2105
rect 3410 -2170 3470 -2135
rect 3410 -2200 3425 -2170
rect 3455 -2200 3470 -2170
rect 3410 -2240 3470 -2200
rect 3410 -2270 3425 -2240
rect 3455 -2270 3470 -2240
rect 3410 -2310 3470 -2270
rect 3410 -2340 3425 -2310
rect 3455 -2340 3470 -2310
rect 3410 -2380 3470 -2340
rect 3410 -2410 3425 -2380
rect 3455 -2410 3470 -2380
rect 3410 -2445 3470 -2410
rect 3410 -2475 3425 -2445
rect 3455 -2475 3470 -2445
rect 3410 -2505 3470 -2475
rect 3410 -2535 3425 -2505
rect 3455 -2535 3470 -2505
rect 3410 -2570 3470 -2535
rect 3410 -2600 3425 -2570
rect 3455 -2600 3470 -2570
rect 3410 -2640 3470 -2600
rect 3410 -2670 3425 -2640
rect 3455 -2670 3470 -2640
rect 3410 -2710 3470 -2670
rect 3410 -2740 3425 -2710
rect 3455 -2740 3470 -2710
rect 3410 -2780 3470 -2740
rect 3410 -2810 3425 -2780
rect 3455 -2810 3470 -2780
rect 3410 -2845 3470 -2810
rect 3410 -2875 3425 -2845
rect 3455 -2875 3470 -2845
rect 3410 -2905 3470 -2875
rect 3410 -2935 3425 -2905
rect 3455 -2935 3470 -2905
rect 3410 -2970 3470 -2935
rect 3410 -3000 3425 -2970
rect 3455 -3000 3470 -2970
rect 3410 -3040 3470 -3000
rect 3410 -3070 3425 -3040
rect 3455 -3070 3470 -3040
rect 3410 -3110 3470 -3070
rect 3410 -3140 3425 -3110
rect 3455 -3140 3470 -3110
rect 3410 -3180 3470 -3140
rect 3410 -3210 3425 -3180
rect 3455 -3210 3470 -3180
rect 3410 -3245 3470 -3210
rect 3410 -3275 3425 -3245
rect 3455 -3275 3470 -3245
rect 3410 -3305 3470 -3275
rect 3410 -3335 3425 -3305
rect 3455 -3335 3470 -3305
rect 3410 -3370 3470 -3335
rect 3410 -3400 3425 -3370
rect 3455 -3400 3470 -3370
rect 3410 -3440 3470 -3400
rect 3410 -3470 3425 -3440
rect 3455 -3470 3470 -3440
rect 3410 -3510 3470 -3470
rect 3410 -3540 3425 -3510
rect 3455 -3540 3470 -3510
rect 3410 -3580 3470 -3540
rect 3410 -3610 3425 -3580
rect 3455 -3610 3470 -3580
rect 3410 -3645 3470 -3610
rect 3410 -3675 3425 -3645
rect 3455 -3675 3470 -3645
rect 3410 -3705 3470 -3675
rect 3410 -3735 3425 -3705
rect 3455 -3735 3470 -3705
rect 3410 -3770 3470 -3735
rect 3410 -3800 3425 -3770
rect 3455 -3800 3470 -3770
rect 3410 -3840 3470 -3800
rect 3410 -3870 3425 -3840
rect 3455 -3870 3470 -3840
rect 3410 -3910 3470 -3870
rect 3410 -3940 3425 -3910
rect 3455 -3940 3470 -3910
rect 3410 -3980 3470 -3940
rect 3410 -4010 3425 -3980
rect 3455 -4010 3470 -3980
rect 3410 -4045 3470 -4010
rect 3410 -4075 3425 -4045
rect 3455 -4075 3470 -4045
rect 3410 -4105 3470 -4075
rect 3410 -4135 3425 -4105
rect 3455 -4135 3470 -4105
rect 3410 -4170 3470 -4135
rect 3410 -4200 3425 -4170
rect 3455 -4200 3470 -4170
rect 3410 -4240 3470 -4200
rect 3410 -4270 3425 -4240
rect 3455 -4270 3470 -4240
rect 3410 -4310 3470 -4270
rect 3410 -4340 3425 -4310
rect 3455 -4340 3470 -4310
rect 3410 -4380 3470 -4340
rect 3410 -4410 3425 -4380
rect 3455 -4410 3470 -4380
rect 3410 -4445 3470 -4410
rect 3410 -4475 3425 -4445
rect 3455 -4475 3470 -4445
rect 3410 -4490 3470 -4475
rect 3760 -1305 3820 -1290
rect 3760 -1335 3775 -1305
rect 3805 -1335 3820 -1305
rect 3760 -1370 3820 -1335
rect 3760 -1400 3775 -1370
rect 3805 -1400 3820 -1370
rect 3760 -1440 3820 -1400
rect 3760 -1470 3775 -1440
rect 3805 -1470 3820 -1440
rect 3760 -1510 3820 -1470
rect 3760 -1540 3775 -1510
rect 3805 -1540 3820 -1510
rect 3760 -1580 3820 -1540
rect 3760 -1610 3775 -1580
rect 3805 -1610 3820 -1580
rect 3760 -1645 3820 -1610
rect 3760 -1675 3775 -1645
rect 3805 -1675 3820 -1645
rect 3760 -1705 3820 -1675
rect 3760 -1735 3775 -1705
rect 3805 -1735 3820 -1705
rect 3760 -1770 3820 -1735
rect 3760 -1800 3775 -1770
rect 3805 -1800 3820 -1770
rect 3760 -1840 3820 -1800
rect 3760 -1870 3775 -1840
rect 3805 -1870 3820 -1840
rect 3760 -1910 3820 -1870
rect 3760 -1940 3775 -1910
rect 3805 -1940 3820 -1910
rect 3760 -1980 3820 -1940
rect 3760 -2010 3775 -1980
rect 3805 -2010 3820 -1980
rect 3760 -2045 3820 -2010
rect 3760 -2075 3775 -2045
rect 3805 -2075 3820 -2045
rect 3760 -2105 3820 -2075
rect 3760 -2135 3775 -2105
rect 3805 -2135 3820 -2105
rect 3760 -2170 3820 -2135
rect 3760 -2200 3775 -2170
rect 3805 -2200 3820 -2170
rect 3760 -2240 3820 -2200
rect 3760 -2270 3775 -2240
rect 3805 -2270 3820 -2240
rect 3760 -2310 3820 -2270
rect 3760 -2340 3775 -2310
rect 3805 -2340 3820 -2310
rect 3760 -2380 3820 -2340
rect 3760 -2410 3775 -2380
rect 3805 -2410 3820 -2380
rect 3760 -2445 3820 -2410
rect 3760 -2475 3775 -2445
rect 3805 -2475 3820 -2445
rect 3760 -2505 3820 -2475
rect 3760 -2535 3775 -2505
rect 3805 -2535 3820 -2505
rect 3760 -2570 3820 -2535
rect 3760 -2600 3775 -2570
rect 3805 -2600 3820 -2570
rect 3760 -2640 3820 -2600
rect 3760 -2670 3775 -2640
rect 3805 -2670 3820 -2640
rect 3760 -2710 3820 -2670
rect 3760 -2740 3775 -2710
rect 3805 -2740 3820 -2710
rect 3760 -2780 3820 -2740
rect 3760 -2810 3775 -2780
rect 3805 -2810 3820 -2780
rect 3760 -2845 3820 -2810
rect 3760 -2875 3775 -2845
rect 3805 -2875 3820 -2845
rect 3760 -2905 3820 -2875
rect 3760 -2935 3775 -2905
rect 3805 -2935 3820 -2905
rect 3760 -2970 3820 -2935
rect 3760 -3000 3775 -2970
rect 3805 -3000 3820 -2970
rect 3760 -3040 3820 -3000
rect 3760 -3070 3775 -3040
rect 3805 -3070 3820 -3040
rect 3760 -3110 3820 -3070
rect 3760 -3140 3775 -3110
rect 3805 -3140 3820 -3110
rect 3760 -3180 3820 -3140
rect 3760 -3210 3775 -3180
rect 3805 -3210 3820 -3180
rect 3760 -3245 3820 -3210
rect 3760 -3275 3775 -3245
rect 3805 -3275 3820 -3245
rect 3760 -3305 3820 -3275
rect 3760 -3335 3775 -3305
rect 3805 -3335 3820 -3305
rect 3760 -3370 3820 -3335
rect 3760 -3400 3775 -3370
rect 3805 -3400 3820 -3370
rect 3760 -3440 3820 -3400
rect 3760 -3470 3775 -3440
rect 3805 -3470 3820 -3440
rect 3760 -3510 3820 -3470
rect 3760 -3540 3775 -3510
rect 3805 -3540 3820 -3510
rect 3760 -3580 3820 -3540
rect 3760 -3610 3775 -3580
rect 3805 -3610 3820 -3580
rect 3760 -3645 3820 -3610
rect 3760 -3675 3775 -3645
rect 3805 -3675 3820 -3645
rect 3760 -3705 3820 -3675
rect 3760 -3735 3775 -3705
rect 3805 -3735 3820 -3705
rect 3760 -3770 3820 -3735
rect 3760 -3800 3775 -3770
rect 3805 -3800 3820 -3770
rect 3760 -3840 3820 -3800
rect 3760 -3870 3775 -3840
rect 3805 -3870 3820 -3840
rect 3760 -3910 3820 -3870
rect 3760 -3940 3775 -3910
rect 3805 -3940 3820 -3910
rect 3760 -3980 3820 -3940
rect 3760 -4010 3775 -3980
rect 3805 -4010 3820 -3980
rect 3760 -4045 3820 -4010
rect 3760 -4075 3775 -4045
rect 3805 -4075 3820 -4045
rect 3760 -4105 3820 -4075
rect 3760 -4135 3775 -4105
rect 3805 -4135 3820 -4105
rect 3760 -4170 3820 -4135
rect 3760 -4200 3775 -4170
rect 3805 -4200 3820 -4170
rect 3760 -4240 3820 -4200
rect 3760 -4270 3775 -4240
rect 3805 -4270 3820 -4240
rect 3760 -4310 3820 -4270
rect 3760 -4340 3775 -4310
rect 3805 -4340 3820 -4310
rect 3760 -4380 3820 -4340
rect 3760 -4410 3775 -4380
rect 3805 -4410 3820 -4380
rect 3760 -4445 3820 -4410
rect 3760 -4475 3775 -4445
rect 3805 -4475 3820 -4445
rect 3760 -4490 3820 -4475
rect 4110 -1305 4170 -1290
rect 4110 -1335 4125 -1305
rect 4155 -1335 4170 -1305
rect 4110 -1370 4170 -1335
rect 4110 -1400 4125 -1370
rect 4155 -1400 4170 -1370
rect 4110 -1440 4170 -1400
rect 4110 -1470 4125 -1440
rect 4155 -1470 4170 -1440
rect 4110 -1510 4170 -1470
rect 4110 -1540 4125 -1510
rect 4155 -1540 4170 -1510
rect 4110 -1580 4170 -1540
rect 4110 -1610 4125 -1580
rect 4155 -1610 4170 -1580
rect 4110 -1645 4170 -1610
rect 4110 -1675 4125 -1645
rect 4155 -1675 4170 -1645
rect 4110 -1705 4170 -1675
rect 4110 -1735 4125 -1705
rect 4155 -1735 4170 -1705
rect 4110 -1770 4170 -1735
rect 4110 -1800 4125 -1770
rect 4155 -1800 4170 -1770
rect 4110 -1840 4170 -1800
rect 4110 -1870 4125 -1840
rect 4155 -1870 4170 -1840
rect 4110 -1910 4170 -1870
rect 4110 -1940 4125 -1910
rect 4155 -1940 4170 -1910
rect 4110 -1980 4170 -1940
rect 4110 -2010 4125 -1980
rect 4155 -2010 4170 -1980
rect 4110 -2045 4170 -2010
rect 4110 -2075 4125 -2045
rect 4155 -2075 4170 -2045
rect 4110 -2105 4170 -2075
rect 4110 -2135 4125 -2105
rect 4155 -2135 4170 -2105
rect 4110 -2170 4170 -2135
rect 4110 -2200 4125 -2170
rect 4155 -2200 4170 -2170
rect 4110 -2240 4170 -2200
rect 4110 -2270 4125 -2240
rect 4155 -2270 4170 -2240
rect 4110 -2310 4170 -2270
rect 4110 -2340 4125 -2310
rect 4155 -2340 4170 -2310
rect 4110 -2380 4170 -2340
rect 4110 -2410 4125 -2380
rect 4155 -2410 4170 -2380
rect 4110 -2445 4170 -2410
rect 4110 -2475 4125 -2445
rect 4155 -2475 4170 -2445
rect 4110 -2505 4170 -2475
rect 4110 -2535 4125 -2505
rect 4155 -2535 4170 -2505
rect 4110 -2570 4170 -2535
rect 4110 -2600 4125 -2570
rect 4155 -2600 4170 -2570
rect 4110 -2640 4170 -2600
rect 4110 -2670 4125 -2640
rect 4155 -2670 4170 -2640
rect 4110 -2710 4170 -2670
rect 4110 -2740 4125 -2710
rect 4155 -2740 4170 -2710
rect 4110 -2780 4170 -2740
rect 4110 -2810 4125 -2780
rect 4155 -2810 4170 -2780
rect 4110 -2845 4170 -2810
rect 4110 -2875 4125 -2845
rect 4155 -2875 4170 -2845
rect 4110 -2905 4170 -2875
rect 4110 -2935 4125 -2905
rect 4155 -2935 4170 -2905
rect 4110 -2970 4170 -2935
rect 4110 -3000 4125 -2970
rect 4155 -3000 4170 -2970
rect 4110 -3040 4170 -3000
rect 4110 -3070 4125 -3040
rect 4155 -3070 4170 -3040
rect 4110 -3110 4170 -3070
rect 4110 -3140 4125 -3110
rect 4155 -3140 4170 -3110
rect 4110 -3180 4170 -3140
rect 4110 -3210 4125 -3180
rect 4155 -3210 4170 -3180
rect 4110 -3245 4170 -3210
rect 4110 -3275 4125 -3245
rect 4155 -3275 4170 -3245
rect 4110 -3305 4170 -3275
rect 4110 -3335 4125 -3305
rect 4155 -3335 4170 -3305
rect 4110 -3370 4170 -3335
rect 4110 -3400 4125 -3370
rect 4155 -3400 4170 -3370
rect 4110 -3440 4170 -3400
rect 4110 -3470 4125 -3440
rect 4155 -3470 4170 -3440
rect 4110 -3510 4170 -3470
rect 4110 -3540 4125 -3510
rect 4155 -3540 4170 -3510
rect 4110 -3580 4170 -3540
rect 4110 -3610 4125 -3580
rect 4155 -3610 4170 -3580
rect 4110 -3645 4170 -3610
rect 4110 -3675 4125 -3645
rect 4155 -3675 4170 -3645
rect 4110 -3705 4170 -3675
rect 4110 -3735 4125 -3705
rect 4155 -3735 4170 -3705
rect 4110 -3770 4170 -3735
rect 4110 -3800 4125 -3770
rect 4155 -3800 4170 -3770
rect 4110 -3840 4170 -3800
rect 4110 -3870 4125 -3840
rect 4155 -3870 4170 -3840
rect 4110 -3910 4170 -3870
rect 4110 -3940 4125 -3910
rect 4155 -3940 4170 -3910
rect 4110 -3980 4170 -3940
rect 4110 -4010 4125 -3980
rect 4155 -4010 4170 -3980
rect 4110 -4045 4170 -4010
rect 4110 -4075 4125 -4045
rect 4155 -4075 4170 -4045
rect 4110 -4105 4170 -4075
rect 4110 -4135 4125 -4105
rect 4155 -4135 4170 -4105
rect 4110 -4170 4170 -4135
rect 4110 -4200 4125 -4170
rect 4155 -4200 4170 -4170
rect 4110 -4240 4170 -4200
rect 4110 -4270 4125 -4240
rect 4155 -4270 4170 -4240
rect 4110 -4310 4170 -4270
rect 4110 -4340 4125 -4310
rect 4155 -4340 4170 -4310
rect 4110 -4380 4170 -4340
rect 4110 -4410 4125 -4380
rect 4155 -4410 4170 -4380
rect 4110 -4445 4170 -4410
rect 4110 -4475 4125 -4445
rect 4155 -4475 4170 -4445
rect 4110 -4490 4170 -4475
rect 4460 -1305 4520 -1290
rect 4460 -1335 4475 -1305
rect 4505 -1335 4520 -1305
rect 4460 -1370 4520 -1335
rect 4460 -1400 4475 -1370
rect 4505 -1400 4520 -1370
rect 4460 -1440 4520 -1400
rect 4460 -1470 4475 -1440
rect 4505 -1470 4520 -1440
rect 4460 -1510 4520 -1470
rect 4460 -1540 4475 -1510
rect 4505 -1540 4520 -1510
rect 4460 -1580 4520 -1540
rect 4460 -1610 4475 -1580
rect 4505 -1610 4520 -1580
rect 4460 -1645 4520 -1610
rect 4460 -1675 4475 -1645
rect 4505 -1675 4520 -1645
rect 4460 -1705 4520 -1675
rect 4460 -1735 4475 -1705
rect 4505 -1735 4520 -1705
rect 4460 -1770 4520 -1735
rect 4460 -1800 4475 -1770
rect 4505 -1800 4520 -1770
rect 4460 -1840 4520 -1800
rect 4460 -1870 4475 -1840
rect 4505 -1870 4520 -1840
rect 4460 -1910 4520 -1870
rect 4460 -1940 4475 -1910
rect 4505 -1940 4520 -1910
rect 4460 -1980 4520 -1940
rect 4460 -2010 4475 -1980
rect 4505 -2010 4520 -1980
rect 4460 -2045 4520 -2010
rect 4460 -2075 4475 -2045
rect 4505 -2075 4520 -2045
rect 4460 -2105 4520 -2075
rect 4460 -2135 4475 -2105
rect 4505 -2135 4520 -2105
rect 4460 -2170 4520 -2135
rect 4460 -2200 4475 -2170
rect 4505 -2200 4520 -2170
rect 4460 -2240 4520 -2200
rect 4460 -2270 4475 -2240
rect 4505 -2270 4520 -2240
rect 4460 -2310 4520 -2270
rect 4460 -2340 4475 -2310
rect 4505 -2340 4520 -2310
rect 4460 -2380 4520 -2340
rect 4460 -2410 4475 -2380
rect 4505 -2410 4520 -2380
rect 4460 -2445 4520 -2410
rect 4460 -2475 4475 -2445
rect 4505 -2475 4520 -2445
rect 4460 -2505 4520 -2475
rect 4460 -2535 4475 -2505
rect 4505 -2535 4520 -2505
rect 4460 -2570 4520 -2535
rect 4460 -2600 4475 -2570
rect 4505 -2600 4520 -2570
rect 4460 -2640 4520 -2600
rect 4460 -2670 4475 -2640
rect 4505 -2670 4520 -2640
rect 4460 -2710 4520 -2670
rect 4460 -2740 4475 -2710
rect 4505 -2740 4520 -2710
rect 4460 -2780 4520 -2740
rect 4460 -2810 4475 -2780
rect 4505 -2810 4520 -2780
rect 4460 -2845 4520 -2810
rect 4460 -2875 4475 -2845
rect 4505 -2875 4520 -2845
rect 4460 -2905 4520 -2875
rect 4460 -2935 4475 -2905
rect 4505 -2935 4520 -2905
rect 4460 -2970 4520 -2935
rect 4460 -3000 4475 -2970
rect 4505 -3000 4520 -2970
rect 4460 -3040 4520 -3000
rect 4460 -3070 4475 -3040
rect 4505 -3070 4520 -3040
rect 4460 -3110 4520 -3070
rect 4460 -3140 4475 -3110
rect 4505 -3140 4520 -3110
rect 4460 -3180 4520 -3140
rect 4460 -3210 4475 -3180
rect 4505 -3210 4520 -3180
rect 4460 -3245 4520 -3210
rect 4460 -3275 4475 -3245
rect 4505 -3275 4520 -3245
rect 4460 -3305 4520 -3275
rect 4460 -3335 4475 -3305
rect 4505 -3335 4520 -3305
rect 4460 -3370 4520 -3335
rect 4460 -3400 4475 -3370
rect 4505 -3400 4520 -3370
rect 4460 -3440 4520 -3400
rect 4460 -3470 4475 -3440
rect 4505 -3470 4520 -3440
rect 4460 -3510 4520 -3470
rect 4460 -3540 4475 -3510
rect 4505 -3540 4520 -3510
rect 4460 -3580 4520 -3540
rect 4460 -3610 4475 -3580
rect 4505 -3610 4520 -3580
rect 4460 -3645 4520 -3610
rect 4460 -3675 4475 -3645
rect 4505 -3675 4520 -3645
rect 4460 -3705 4520 -3675
rect 4460 -3735 4475 -3705
rect 4505 -3735 4520 -3705
rect 4460 -3770 4520 -3735
rect 4460 -3800 4475 -3770
rect 4505 -3800 4520 -3770
rect 4460 -3840 4520 -3800
rect 4460 -3870 4475 -3840
rect 4505 -3870 4520 -3840
rect 4460 -3910 4520 -3870
rect 4460 -3940 4475 -3910
rect 4505 -3940 4520 -3910
rect 4460 -3980 4520 -3940
rect 4460 -4010 4475 -3980
rect 4505 -4010 4520 -3980
rect 4460 -4045 4520 -4010
rect 4460 -4075 4475 -4045
rect 4505 -4075 4520 -4045
rect 4460 -4105 4520 -4075
rect 4460 -4135 4475 -4105
rect 4505 -4135 4520 -4105
rect 4460 -4170 4520 -4135
rect 4460 -4200 4475 -4170
rect 4505 -4200 4520 -4170
rect 4460 -4240 4520 -4200
rect 4460 -4270 4475 -4240
rect 4505 -4270 4520 -4240
rect 4460 -4310 4520 -4270
rect 4460 -4340 4475 -4310
rect 4505 -4340 4520 -4310
rect 4460 -4380 4520 -4340
rect 4460 -4410 4475 -4380
rect 4505 -4410 4520 -4380
rect 4460 -4445 4520 -4410
rect 4460 -4475 4475 -4445
rect 4505 -4475 4520 -4445
rect 4460 -4490 4520 -4475
rect 4810 -1305 4870 -1290
rect 4810 -1335 4825 -1305
rect 4855 -1335 4870 -1305
rect 4810 -1370 4870 -1335
rect 4810 -1400 4825 -1370
rect 4855 -1400 4870 -1370
rect 4810 -1440 4870 -1400
rect 4810 -1470 4825 -1440
rect 4855 -1470 4870 -1440
rect 4810 -1510 4870 -1470
rect 4810 -1540 4825 -1510
rect 4855 -1540 4870 -1510
rect 4810 -1580 4870 -1540
rect 4810 -1610 4825 -1580
rect 4855 -1610 4870 -1580
rect 4810 -1645 4870 -1610
rect 4810 -1675 4825 -1645
rect 4855 -1675 4870 -1645
rect 4810 -1705 4870 -1675
rect 4810 -1735 4825 -1705
rect 4855 -1735 4870 -1705
rect 4810 -1770 4870 -1735
rect 4810 -1800 4825 -1770
rect 4855 -1800 4870 -1770
rect 4810 -1840 4870 -1800
rect 4810 -1870 4825 -1840
rect 4855 -1870 4870 -1840
rect 4810 -1910 4870 -1870
rect 4810 -1940 4825 -1910
rect 4855 -1940 4870 -1910
rect 4810 -1980 4870 -1940
rect 4810 -2010 4825 -1980
rect 4855 -2010 4870 -1980
rect 4810 -2045 4870 -2010
rect 4810 -2075 4825 -2045
rect 4855 -2075 4870 -2045
rect 4810 -2105 4870 -2075
rect 4810 -2135 4825 -2105
rect 4855 -2135 4870 -2105
rect 4810 -2170 4870 -2135
rect 4810 -2200 4825 -2170
rect 4855 -2200 4870 -2170
rect 4810 -2240 4870 -2200
rect 4810 -2270 4825 -2240
rect 4855 -2270 4870 -2240
rect 4810 -2310 4870 -2270
rect 4810 -2340 4825 -2310
rect 4855 -2340 4870 -2310
rect 4810 -2380 4870 -2340
rect 4810 -2410 4825 -2380
rect 4855 -2410 4870 -2380
rect 4810 -2445 4870 -2410
rect 4810 -2475 4825 -2445
rect 4855 -2475 4870 -2445
rect 4810 -2505 4870 -2475
rect 4810 -2535 4825 -2505
rect 4855 -2535 4870 -2505
rect 4810 -2570 4870 -2535
rect 4810 -2600 4825 -2570
rect 4855 -2600 4870 -2570
rect 4810 -2640 4870 -2600
rect 4810 -2670 4825 -2640
rect 4855 -2670 4870 -2640
rect 4810 -2710 4870 -2670
rect 4810 -2740 4825 -2710
rect 4855 -2740 4870 -2710
rect 4810 -2780 4870 -2740
rect 4810 -2810 4825 -2780
rect 4855 -2810 4870 -2780
rect 4810 -2845 4870 -2810
rect 4810 -2875 4825 -2845
rect 4855 -2875 4870 -2845
rect 4810 -2905 4870 -2875
rect 4810 -2935 4825 -2905
rect 4855 -2935 4870 -2905
rect 4810 -2970 4870 -2935
rect 4810 -3000 4825 -2970
rect 4855 -3000 4870 -2970
rect 4810 -3040 4870 -3000
rect 4810 -3070 4825 -3040
rect 4855 -3070 4870 -3040
rect 4810 -3110 4870 -3070
rect 4810 -3140 4825 -3110
rect 4855 -3140 4870 -3110
rect 4810 -3180 4870 -3140
rect 4810 -3210 4825 -3180
rect 4855 -3210 4870 -3180
rect 4810 -3245 4870 -3210
rect 4810 -3275 4825 -3245
rect 4855 -3275 4870 -3245
rect 4810 -3305 4870 -3275
rect 4810 -3335 4825 -3305
rect 4855 -3335 4870 -3305
rect 4810 -3370 4870 -3335
rect 4810 -3400 4825 -3370
rect 4855 -3400 4870 -3370
rect 4810 -3440 4870 -3400
rect 4810 -3470 4825 -3440
rect 4855 -3470 4870 -3440
rect 4810 -3510 4870 -3470
rect 4810 -3540 4825 -3510
rect 4855 -3540 4870 -3510
rect 4810 -3580 4870 -3540
rect 4810 -3610 4825 -3580
rect 4855 -3610 4870 -3580
rect 4810 -3645 4870 -3610
rect 4810 -3675 4825 -3645
rect 4855 -3675 4870 -3645
rect 4810 -3705 4870 -3675
rect 4810 -3735 4825 -3705
rect 4855 -3735 4870 -3705
rect 4810 -3770 4870 -3735
rect 4810 -3800 4825 -3770
rect 4855 -3800 4870 -3770
rect 4810 -3840 4870 -3800
rect 4810 -3870 4825 -3840
rect 4855 -3870 4870 -3840
rect 4810 -3910 4870 -3870
rect 4810 -3940 4825 -3910
rect 4855 -3940 4870 -3910
rect 4810 -3980 4870 -3940
rect 4810 -4010 4825 -3980
rect 4855 -4010 4870 -3980
rect 4810 -4045 4870 -4010
rect 4810 -4075 4825 -4045
rect 4855 -4075 4870 -4045
rect 4810 -4105 4870 -4075
rect 4810 -4135 4825 -4105
rect 4855 -4135 4870 -4105
rect 4810 -4170 4870 -4135
rect 4810 -4200 4825 -4170
rect 4855 -4200 4870 -4170
rect 4810 -4240 4870 -4200
rect 4810 -4270 4825 -4240
rect 4855 -4270 4870 -4240
rect 4810 -4310 4870 -4270
rect 4810 -4340 4825 -4310
rect 4855 -4340 4870 -4310
rect 4810 -4380 4870 -4340
rect 4810 -4410 4825 -4380
rect 4855 -4410 4870 -4380
rect 4810 -4445 4870 -4410
rect 4810 -4475 4825 -4445
rect 4855 -4475 4870 -4445
rect 4810 -4490 4870 -4475
rect 5160 -1305 5220 -1290
rect 5160 -1335 5175 -1305
rect 5205 -1335 5220 -1305
rect 5160 -1370 5220 -1335
rect 5160 -1400 5175 -1370
rect 5205 -1400 5220 -1370
rect 5160 -1440 5220 -1400
rect 5160 -1470 5175 -1440
rect 5205 -1470 5220 -1440
rect 5160 -1510 5220 -1470
rect 5160 -1540 5175 -1510
rect 5205 -1540 5220 -1510
rect 5160 -1580 5220 -1540
rect 5160 -1610 5175 -1580
rect 5205 -1610 5220 -1580
rect 5160 -1645 5220 -1610
rect 5160 -1675 5175 -1645
rect 5205 -1675 5220 -1645
rect 5160 -1705 5220 -1675
rect 5160 -1735 5175 -1705
rect 5205 -1735 5220 -1705
rect 5160 -1770 5220 -1735
rect 5160 -1800 5175 -1770
rect 5205 -1800 5220 -1770
rect 5160 -1840 5220 -1800
rect 5160 -1870 5175 -1840
rect 5205 -1870 5220 -1840
rect 5160 -1910 5220 -1870
rect 5160 -1940 5175 -1910
rect 5205 -1940 5220 -1910
rect 5160 -1980 5220 -1940
rect 5160 -2010 5175 -1980
rect 5205 -2010 5220 -1980
rect 5160 -2045 5220 -2010
rect 5160 -2075 5175 -2045
rect 5205 -2075 5220 -2045
rect 5160 -2105 5220 -2075
rect 5160 -2135 5175 -2105
rect 5205 -2135 5220 -2105
rect 5160 -2170 5220 -2135
rect 5160 -2200 5175 -2170
rect 5205 -2200 5220 -2170
rect 5160 -2240 5220 -2200
rect 5160 -2270 5175 -2240
rect 5205 -2270 5220 -2240
rect 5160 -2310 5220 -2270
rect 5160 -2340 5175 -2310
rect 5205 -2340 5220 -2310
rect 5160 -2380 5220 -2340
rect 5160 -2410 5175 -2380
rect 5205 -2410 5220 -2380
rect 5160 -2445 5220 -2410
rect 5160 -2475 5175 -2445
rect 5205 -2475 5220 -2445
rect 5160 -2505 5220 -2475
rect 5160 -2535 5175 -2505
rect 5205 -2535 5220 -2505
rect 5160 -2570 5220 -2535
rect 5160 -2600 5175 -2570
rect 5205 -2600 5220 -2570
rect 5160 -2640 5220 -2600
rect 5160 -2670 5175 -2640
rect 5205 -2670 5220 -2640
rect 5160 -2710 5220 -2670
rect 5160 -2740 5175 -2710
rect 5205 -2740 5220 -2710
rect 5160 -2780 5220 -2740
rect 5160 -2810 5175 -2780
rect 5205 -2810 5220 -2780
rect 5160 -2845 5220 -2810
rect 5160 -2875 5175 -2845
rect 5205 -2875 5220 -2845
rect 5160 -2905 5220 -2875
rect 5160 -2935 5175 -2905
rect 5205 -2935 5220 -2905
rect 5160 -2970 5220 -2935
rect 5160 -3000 5175 -2970
rect 5205 -3000 5220 -2970
rect 5160 -3040 5220 -3000
rect 5160 -3070 5175 -3040
rect 5205 -3070 5220 -3040
rect 5160 -3110 5220 -3070
rect 5160 -3140 5175 -3110
rect 5205 -3140 5220 -3110
rect 5160 -3180 5220 -3140
rect 5160 -3210 5175 -3180
rect 5205 -3210 5220 -3180
rect 5160 -3245 5220 -3210
rect 5160 -3275 5175 -3245
rect 5205 -3275 5220 -3245
rect 5160 -3305 5220 -3275
rect 5160 -3335 5175 -3305
rect 5205 -3335 5220 -3305
rect 5160 -3370 5220 -3335
rect 5160 -3400 5175 -3370
rect 5205 -3400 5220 -3370
rect 5160 -3440 5220 -3400
rect 5160 -3470 5175 -3440
rect 5205 -3470 5220 -3440
rect 5160 -3510 5220 -3470
rect 5160 -3540 5175 -3510
rect 5205 -3540 5220 -3510
rect 5160 -3580 5220 -3540
rect 5160 -3610 5175 -3580
rect 5205 -3610 5220 -3580
rect 5160 -3645 5220 -3610
rect 5160 -3675 5175 -3645
rect 5205 -3675 5220 -3645
rect 5160 -3705 5220 -3675
rect 5160 -3735 5175 -3705
rect 5205 -3735 5220 -3705
rect 5160 -3770 5220 -3735
rect 5160 -3800 5175 -3770
rect 5205 -3800 5220 -3770
rect 5160 -3840 5220 -3800
rect 5160 -3870 5175 -3840
rect 5205 -3870 5220 -3840
rect 5160 -3910 5220 -3870
rect 5160 -3940 5175 -3910
rect 5205 -3940 5220 -3910
rect 5160 -3980 5220 -3940
rect 5160 -4010 5175 -3980
rect 5205 -4010 5220 -3980
rect 5160 -4045 5220 -4010
rect 5160 -4075 5175 -4045
rect 5205 -4075 5220 -4045
rect 5160 -4105 5220 -4075
rect 5160 -4135 5175 -4105
rect 5205 -4135 5220 -4105
rect 5160 -4170 5220 -4135
rect 5160 -4200 5175 -4170
rect 5205 -4200 5220 -4170
rect 5160 -4240 5220 -4200
rect 5160 -4270 5175 -4240
rect 5205 -4270 5220 -4240
rect 5160 -4310 5220 -4270
rect 5160 -4340 5175 -4310
rect 5205 -4340 5220 -4310
rect 5160 -4380 5220 -4340
rect 5160 -4410 5175 -4380
rect 5205 -4410 5220 -4380
rect 5160 -4445 5220 -4410
rect 5160 -4475 5175 -4445
rect 5205 -4475 5220 -4445
rect 5160 -4490 5220 -4475
rect 5510 -1305 5570 -1290
rect 5510 -1335 5525 -1305
rect 5555 -1335 5570 -1305
rect 5510 -1370 5570 -1335
rect 5510 -1400 5525 -1370
rect 5555 -1400 5570 -1370
rect 5510 -1440 5570 -1400
rect 5510 -1470 5525 -1440
rect 5555 -1470 5570 -1440
rect 5510 -1510 5570 -1470
rect 5510 -1540 5525 -1510
rect 5555 -1540 5570 -1510
rect 5510 -1580 5570 -1540
rect 5510 -1610 5525 -1580
rect 5555 -1610 5570 -1580
rect 5510 -1645 5570 -1610
rect 5510 -1675 5525 -1645
rect 5555 -1675 5570 -1645
rect 5510 -1705 5570 -1675
rect 5510 -1735 5525 -1705
rect 5555 -1735 5570 -1705
rect 5510 -1770 5570 -1735
rect 5510 -1800 5525 -1770
rect 5555 -1800 5570 -1770
rect 5510 -1840 5570 -1800
rect 5510 -1870 5525 -1840
rect 5555 -1870 5570 -1840
rect 5510 -1910 5570 -1870
rect 5510 -1940 5525 -1910
rect 5555 -1940 5570 -1910
rect 5510 -1980 5570 -1940
rect 5510 -2010 5525 -1980
rect 5555 -2010 5570 -1980
rect 5510 -2045 5570 -2010
rect 5510 -2075 5525 -2045
rect 5555 -2075 5570 -2045
rect 5510 -2105 5570 -2075
rect 5510 -2135 5525 -2105
rect 5555 -2135 5570 -2105
rect 5510 -2170 5570 -2135
rect 5510 -2200 5525 -2170
rect 5555 -2200 5570 -2170
rect 5510 -2240 5570 -2200
rect 5510 -2270 5525 -2240
rect 5555 -2270 5570 -2240
rect 5510 -2310 5570 -2270
rect 5510 -2340 5525 -2310
rect 5555 -2340 5570 -2310
rect 5510 -2380 5570 -2340
rect 5510 -2410 5525 -2380
rect 5555 -2410 5570 -2380
rect 5510 -2445 5570 -2410
rect 5510 -2475 5525 -2445
rect 5555 -2475 5570 -2445
rect 5510 -2505 5570 -2475
rect 5510 -2535 5525 -2505
rect 5555 -2535 5570 -2505
rect 5510 -2570 5570 -2535
rect 5510 -2600 5525 -2570
rect 5555 -2600 5570 -2570
rect 5510 -2640 5570 -2600
rect 5510 -2670 5525 -2640
rect 5555 -2670 5570 -2640
rect 5510 -2710 5570 -2670
rect 5510 -2740 5525 -2710
rect 5555 -2740 5570 -2710
rect 5510 -2780 5570 -2740
rect 5510 -2810 5525 -2780
rect 5555 -2810 5570 -2780
rect 5510 -2845 5570 -2810
rect 5510 -2875 5525 -2845
rect 5555 -2875 5570 -2845
rect 5510 -2905 5570 -2875
rect 5510 -2935 5525 -2905
rect 5555 -2935 5570 -2905
rect 5510 -2970 5570 -2935
rect 5510 -3000 5525 -2970
rect 5555 -3000 5570 -2970
rect 5510 -3040 5570 -3000
rect 5510 -3070 5525 -3040
rect 5555 -3070 5570 -3040
rect 5510 -3110 5570 -3070
rect 5510 -3140 5525 -3110
rect 5555 -3140 5570 -3110
rect 5510 -3180 5570 -3140
rect 5510 -3210 5525 -3180
rect 5555 -3210 5570 -3180
rect 5510 -3245 5570 -3210
rect 5510 -3275 5525 -3245
rect 5555 -3275 5570 -3245
rect 5510 -3305 5570 -3275
rect 5510 -3335 5525 -3305
rect 5555 -3335 5570 -3305
rect 5510 -3370 5570 -3335
rect 5510 -3400 5525 -3370
rect 5555 -3400 5570 -3370
rect 5510 -3440 5570 -3400
rect 5510 -3470 5525 -3440
rect 5555 -3470 5570 -3440
rect 5510 -3510 5570 -3470
rect 5510 -3540 5525 -3510
rect 5555 -3540 5570 -3510
rect 5510 -3580 5570 -3540
rect 5510 -3610 5525 -3580
rect 5555 -3610 5570 -3580
rect 5510 -3645 5570 -3610
rect 5510 -3675 5525 -3645
rect 5555 -3675 5570 -3645
rect 5510 -3705 5570 -3675
rect 5510 -3735 5525 -3705
rect 5555 -3735 5570 -3705
rect 5510 -3770 5570 -3735
rect 5510 -3800 5525 -3770
rect 5555 -3800 5570 -3770
rect 5510 -3840 5570 -3800
rect 5510 -3870 5525 -3840
rect 5555 -3870 5570 -3840
rect 5510 -3910 5570 -3870
rect 5510 -3940 5525 -3910
rect 5555 -3940 5570 -3910
rect 5510 -3980 5570 -3940
rect 5510 -4010 5525 -3980
rect 5555 -4010 5570 -3980
rect 5510 -4045 5570 -4010
rect 5510 -4075 5525 -4045
rect 5555 -4075 5570 -4045
rect 5510 -4105 5570 -4075
rect 5510 -4135 5525 -4105
rect 5555 -4135 5570 -4105
rect 5510 -4170 5570 -4135
rect 5510 -4200 5525 -4170
rect 5555 -4200 5570 -4170
rect 5510 -4240 5570 -4200
rect 5510 -4270 5525 -4240
rect 5555 -4270 5570 -4240
rect 5510 -4310 5570 -4270
rect 5510 -4340 5525 -4310
rect 5555 -4340 5570 -4310
rect 5510 -4380 5570 -4340
rect 5510 -4410 5525 -4380
rect 5555 -4410 5570 -4380
rect 5510 -4445 5570 -4410
rect 5510 -4475 5525 -4445
rect 5555 -4475 5570 -4445
rect 5510 -4490 5570 -4475
rect 5860 -1305 5920 -1290
rect 5860 -1335 5875 -1305
rect 5905 -1335 5920 -1305
rect 5860 -1370 5920 -1335
rect 5860 -1400 5875 -1370
rect 5905 -1400 5920 -1370
rect 5860 -1440 5920 -1400
rect 5860 -1470 5875 -1440
rect 5905 -1470 5920 -1440
rect 5860 -1510 5920 -1470
rect 5860 -1540 5875 -1510
rect 5905 -1540 5920 -1510
rect 5860 -1580 5920 -1540
rect 5860 -1610 5875 -1580
rect 5905 -1610 5920 -1580
rect 5860 -1645 5920 -1610
rect 5860 -1675 5875 -1645
rect 5905 -1675 5920 -1645
rect 5860 -1705 5920 -1675
rect 5860 -1735 5875 -1705
rect 5905 -1735 5920 -1705
rect 5860 -1770 5920 -1735
rect 5860 -1800 5875 -1770
rect 5905 -1800 5920 -1770
rect 5860 -1840 5920 -1800
rect 5860 -1870 5875 -1840
rect 5905 -1870 5920 -1840
rect 5860 -1910 5920 -1870
rect 5860 -1940 5875 -1910
rect 5905 -1940 5920 -1910
rect 5860 -1980 5920 -1940
rect 5860 -2010 5875 -1980
rect 5905 -2010 5920 -1980
rect 5860 -2045 5920 -2010
rect 5860 -2075 5875 -2045
rect 5905 -2075 5920 -2045
rect 5860 -2105 5920 -2075
rect 5860 -2135 5875 -2105
rect 5905 -2135 5920 -2105
rect 5860 -2170 5920 -2135
rect 5860 -2200 5875 -2170
rect 5905 -2200 5920 -2170
rect 5860 -2240 5920 -2200
rect 5860 -2270 5875 -2240
rect 5905 -2270 5920 -2240
rect 5860 -2310 5920 -2270
rect 5860 -2340 5875 -2310
rect 5905 -2340 5920 -2310
rect 5860 -2380 5920 -2340
rect 5860 -2410 5875 -2380
rect 5905 -2410 5920 -2380
rect 5860 -2445 5920 -2410
rect 5860 -2475 5875 -2445
rect 5905 -2475 5920 -2445
rect 5860 -2505 5920 -2475
rect 5860 -2535 5875 -2505
rect 5905 -2535 5920 -2505
rect 5860 -2570 5920 -2535
rect 5860 -2600 5875 -2570
rect 5905 -2600 5920 -2570
rect 5860 -2640 5920 -2600
rect 5860 -2670 5875 -2640
rect 5905 -2670 5920 -2640
rect 5860 -2710 5920 -2670
rect 5860 -2740 5875 -2710
rect 5905 -2740 5920 -2710
rect 5860 -2780 5920 -2740
rect 5860 -2810 5875 -2780
rect 5905 -2810 5920 -2780
rect 5860 -2845 5920 -2810
rect 5860 -2875 5875 -2845
rect 5905 -2875 5920 -2845
rect 5860 -2905 5920 -2875
rect 5860 -2935 5875 -2905
rect 5905 -2935 5920 -2905
rect 5860 -2970 5920 -2935
rect 5860 -3000 5875 -2970
rect 5905 -3000 5920 -2970
rect 5860 -3040 5920 -3000
rect 5860 -3070 5875 -3040
rect 5905 -3070 5920 -3040
rect 5860 -3110 5920 -3070
rect 5860 -3140 5875 -3110
rect 5905 -3140 5920 -3110
rect 5860 -3180 5920 -3140
rect 5860 -3210 5875 -3180
rect 5905 -3210 5920 -3180
rect 5860 -3245 5920 -3210
rect 5860 -3275 5875 -3245
rect 5905 -3275 5920 -3245
rect 5860 -3305 5920 -3275
rect 5860 -3335 5875 -3305
rect 5905 -3335 5920 -3305
rect 5860 -3370 5920 -3335
rect 5860 -3400 5875 -3370
rect 5905 -3400 5920 -3370
rect 5860 -3440 5920 -3400
rect 5860 -3470 5875 -3440
rect 5905 -3470 5920 -3440
rect 5860 -3510 5920 -3470
rect 5860 -3540 5875 -3510
rect 5905 -3540 5920 -3510
rect 5860 -3580 5920 -3540
rect 5860 -3610 5875 -3580
rect 5905 -3610 5920 -3580
rect 5860 -3645 5920 -3610
rect 5860 -3675 5875 -3645
rect 5905 -3675 5920 -3645
rect 5860 -3705 5920 -3675
rect 5860 -3735 5875 -3705
rect 5905 -3735 5920 -3705
rect 5860 -3770 5920 -3735
rect 5860 -3800 5875 -3770
rect 5905 -3800 5920 -3770
rect 5860 -3840 5920 -3800
rect 5860 -3870 5875 -3840
rect 5905 -3870 5920 -3840
rect 5860 -3910 5920 -3870
rect 5860 -3940 5875 -3910
rect 5905 -3940 5920 -3910
rect 5860 -3980 5920 -3940
rect 5860 -4010 5875 -3980
rect 5905 -4010 5920 -3980
rect 5860 -4045 5920 -4010
rect 5860 -4075 5875 -4045
rect 5905 -4075 5920 -4045
rect 5860 -4105 5920 -4075
rect 5860 -4135 5875 -4105
rect 5905 -4135 5920 -4105
rect 5860 -4170 5920 -4135
rect 5860 -4200 5875 -4170
rect 5905 -4200 5920 -4170
rect 5860 -4240 5920 -4200
rect 5860 -4270 5875 -4240
rect 5905 -4270 5920 -4240
rect 5860 -4310 5920 -4270
rect 5860 -4340 5875 -4310
rect 5905 -4340 5920 -4310
rect 5860 -4380 5920 -4340
rect 5860 -4410 5875 -4380
rect 5905 -4410 5920 -4380
rect 5860 -4445 5920 -4410
rect 5860 -4475 5875 -4445
rect 5905 -4475 5920 -4445
rect 5860 -4490 5920 -4475
rect 6210 -1305 6270 -1290
rect 6210 -1335 6225 -1305
rect 6255 -1335 6270 -1305
rect 6210 -1370 6270 -1335
rect 6210 -1400 6225 -1370
rect 6255 -1400 6270 -1370
rect 6210 -1440 6270 -1400
rect 6210 -1470 6225 -1440
rect 6255 -1470 6270 -1440
rect 6210 -1510 6270 -1470
rect 6210 -1540 6225 -1510
rect 6255 -1540 6270 -1510
rect 6210 -1580 6270 -1540
rect 6210 -1610 6225 -1580
rect 6255 -1610 6270 -1580
rect 6210 -1645 6270 -1610
rect 6210 -1675 6225 -1645
rect 6255 -1675 6270 -1645
rect 6210 -1705 6270 -1675
rect 6210 -1735 6225 -1705
rect 6255 -1735 6270 -1705
rect 6210 -1770 6270 -1735
rect 6210 -1800 6225 -1770
rect 6255 -1800 6270 -1770
rect 6210 -1840 6270 -1800
rect 6210 -1870 6225 -1840
rect 6255 -1870 6270 -1840
rect 6210 -1910 6270 -1870
rect 6210 -1940 6225 -1910
rect 6255 -1940 6270 -1910
rect 6210 -1980 6270 -1940
rect 6210 -2010 6225 -1980
rect 6255 -2010 6270 -1980
rect 6210 -2045 6270 -2010
rect 6210 -2075 6225 -2045
rect 6255 -2075 6270 -2045
rect 6210 -2105 6270 -2075
rect 6210 -2135 6225 -2105
rect 6255 -2135 6270 -2105
rect 6210 -2170 6270 -2135
rect 6210 -2200 6225 -2170
rect 6255 -2200 6270 -2170
rect 6210 -2240 6270 -2200
rect 6210 -2270 6225 -2240
rect 6255 -2270 6270 -2240
rect 6210 -2310 6270 -2270
rect 6210 -2340 6225 -2310
rect 6255 -2340 6270 -2310
rect 6210 -2380 6270 -2340
rect 6210 -2410 6225 -2380
rect 6255 -2410 6270 -2380
rect 6210 -2445 6270 -2410
rect 6210 -2475 6225 -2445
rect 6255 -2475 6270 -2445
rect 6210 -2505 6270 -2475
rect 6210 -2535 6225 -2505
rect 6255 -2535 6270 -2505
rect 6210 -2570 6270 -2535
rect 6210 -2600 6225 -2570
rect 6255 -2600 6270 -2570
rect 6210 -2640 6270 -2600
rect 6210 -2670 6225 -2640
rect 6255 -2670 6270 -2640
rect 6210 -2710 6270 -2670
rect 6210 -2740 6225 -2710
rect 6255 -2740 6270 -2710
rect 6210 -2780 6270 -2740
rect 6210 -2810 6225 -2780
rect 6255 -2810 6270 -2780
rect 6210 -2845 6270 -2810
rect 6210 -2875 6225 -2845
rect 6255 -2875 6270 -2845
rect 6210 -2905 6270 -2875
rect 6210 -2935 6225 -2905
rect 6255 -2935 6270 -2905
rect 6210 -2970 6270 -2935
rect 6210 -3000 6225 -2970
rect 6255 -3000 6270 -2970
rect 6210 -3040 6270 -3000
rect 6210 -3070 6225 -3040
rect 6255 -3070 6270 -3040
rect 6210 -3110 6270 -3070
rect 6210 -3140 6225 -3110
rect 6255 -3140 6270 -3110
rect 6210 -3180 6270 -3140
rect 6210 -3210 6225 -3180
rect 6255 -3210 6270 -3180
rect 6210 -3245 6270 -3210
rect 6210 -3275 6225 -3245
rect 6255 -3275 6270 -3245
rect 6210 -3305 6270 -3275
rect 6210 -3335 6225 -3305
rect 6255 -3335 6270 -3305
rect 6210 -3370 6270 -3335
rect 6210 -3400 6225 -3370
rect 6255 -3400 6270 -3370
rect 6210 -3440 6270 -3400
rect 6210 -3470 6225 -3440
rect 6255 -3470 6270 -3440
rect 6210 -3510 6270 -3470
rect 6210 -3540 6225 -3510
rect 6255 -3540 6270 -3510
rect 6210 -3580 6270 -3540
rect 6210 -3610 6225 -3580
rect 6255 -3610 6270 -3580
rect 6210 -3645 6270 -3610
rect 6210 -3675 6225 -3645
rect 6255 -3675 6270 -3645
rect 6210 -3705 6270 -3675
rect 6210 -3735 6225 -3705
rect 6255 -3735 6270 -3705
rect 6210 -3770 6270 -3735
rect 6210 -3800 6225 -3770
rect 6255 -3800 6270 -3770
rect 6210 -3840 6270 -3800
rect 6210 -3870 6225 -3840
rect 6255 -3870 6270 -3840
rect 6210 -3910 6270 -3870
rect 6210 -3940 6225 -3910
rect 6255 -3940 6270 -3910
rect 6210 -3980 6270 -3940
rect 6210 -4010 6225 -3980
rect 6255 -4010 6270 -3980
rect 6210 -4045 6270 -4010
rect 6210 -4075 6225 -4045
rect 6255 -4075 6270 -4045
rect 6210 -4105 6270 -4075
rect 6210 -4135 6225 -4105
rect 6255 -4135 6270 -4105
rect 6210 -4170 6270 -4135
rect 6210 -4200 6225 -4170
rect 6255 -4200 6270 -4170
rect 6210 -4240 6270 -4200
rect 6210 -4270 6225 -4240
rect 6255 -4270 6270 -4240
rect 6210 -4310 6270 -4270
rect 6210 -4340 6225 -4310
rect 6255 -4340 6270 -4310
rect 6210 -4380 6270 -4340
rect 6210 -4410 6225 -4380
rect 6255 -4410 6270 -4380
rect 6210 -4445 6270 -4410
rect 6210 -4475 6225 -4445
rect 6255 -4475 6270 -4445
rect 6210 -4490 6270 -4475
rect 6560 -1305 6620 -1290
rect 6560 -1335 6575 -1305
rect 6605 -1335 6620 -1305
rect 6560 -1370 6620 -1335
rect 6560 -1400 6575 -1370
rect 6605 -1400 6620 -1370
rect 6560 -1440 6620 -1400
rect 6560 -1470 6575 -1440
rect 6605 -1470 6620 -1440
rect 6560 -1510 6620 -1470
rect 6560 -1540 6575 -1510
rect 6605 -1540 6620 -1510
rect 6560 -1580 6620 -1540
rect 6560 -1610 6575 -1580
rect 6605 -1610 6620 -1580
rect 6560 -1645 6620 -1610
rect 6560 -1675 6575 -1645
rect 6605 -1675 6620 -1645
rect 6560 -1705 6620 -1675
rect 6560 -1735 6575 -1705
rect 6605 -1735 6620 -1705
rect 6560 -1770 6620 -1735
rect 6560 -1800 6575 -1770
rect 6605 -1800 6620 -1770
rect 6560 -1840 6620 -1800
rect 6560 -1870 6575 -1840
rect 6605 -1870 6620 -1840
rect 6560 -1910 6620 -1870
rect 6560 -1940 6575 -1910
rect 6605 -1940 6620 -1910
rect 6560 -1980 6620 -1940
rect 6560 -2010 6575 -1980
rect 6605 -2010 6620 -1980
rect 6560 -2045 6620 -2010
rect 6560 -2075 6575 -2045
rect 6605 -2075 6620 -2045
rect 6560 -2105 6620 -2075
rect 6560 -2135 6575 -2105
rect 6605 -2135 6620 -2105
rect 6560 -2170 6620 -2135
rect 6560 -2200 6575 -2170
rect 6605 -2200 6620 -2170
rect 6560 -2240 6620 -2200
rect 6560 -2270 6575 -2240
rect 6605 -2270 6620 -2240
rect 6560 -2310 6620 -2270
rect 6560 -2340 6575 -2310
rect 6605 -2340 6620 -2310
rect 6560 -2380 6620 -2340
rect 6560 -2410 6575 -2380
rect 6605 -2410 6620 -2380
rect 6560 -2445 6620 -2410
rect 6560 -2475 6575 -2445
rect 6605 -2475 6620 -2445
rect 6560 -2505 6620 -2475
rect 6560 -2535 6575 -2505
rect 6605 -2535 6620 -2505
rect 6560 -2570 6620 -2535
rect 6560 -2600 6575 -2570
rect 6605 -2600 6620 -2570
rect 6560 -2640 6620 -2600
rect 6560 -2670 6575 -2640
rect 6605 -2670 6620 -2640
rect 6560 -2710 6620 -2670
rect 6560 -2740 6575 -2710
rect 6605 -2740 6620 -2710
rect 6560 -2780 6620 -2740
rect 6560 -2810 6575 -2780
rect 6605 -2810 6620 -2780
rect 6560 -2845 6620 -2810
rect 6560 -2875 6575 -2845
rect 6605 -2875 6620 -2845
rect 6560 -2905 6620 -2875
rect 6560 -2935 6575 -2905
rect 6605 -2935 6620 -2905
rect 6560 -2970 6620 -2935
rect 6560 -3000 6575 -2970
rect 6605 -3000 6620 -2970
rect 6560 -3040 6620 -3000
rect 6560 -3070 6575 -3040
rect 6605 -3070 6620 -3040
rect 6560 -3110 6620 -3070
rect 6560 -3140 6575 -3110
rect 6605 -3140 6620 -3110
rect 6560 -3180 6620 -3140
rect 6560 -3210 6575 -3180
rect 6605 -3210 6620 -3180
rect 6560 -3245 6620 -3210
rect 6560 -3275 6575 -3245
rect 6605 -3275 6620 -3245
rect 6560 -3305 6620 -3275
rect 6560 -3335 6575 -3305
rect 6605 -3335 6620 -3305
rect 6560 -3370 6620 -3335
rect 6560 -3400 6575 -3370
rect 6605 -3400 6620 -3370
rect 6560 -3440 6620 -3400
rect 6560 -3470 6575 -3440
rect 6605 -3470 6620 -3440
rect 6560 -3510 6620 -3470
rect 6560 -3540 6575 -3510
rect 6605 -3540 6620 -3510
rect 6560 -3580 6620 -3540
rect 6560 -3610 6575 -3580
rect 6605 -3610 6620 -3580
rect 6560 -3645 6620 -3610
rect 6560 -3675 6575 -3645
rect 6605 -3675 6620 -3645
rect 6560 -3705 6620 -3675
rect 6560 -3735 6575 -3705
rect 6605 -3735 6620 -3705
rect 6560 -3770 6620 -3735
rect 6560 -3800 6575 -3770
rect 6605 -3800 6620 -3770
rect 6560 -3840 6620 -3800
rect 6560 -3870 6575 -3840
rect 6605 -3870 6620 -3840
rect 6560 -3910 6620 -3870
rect 6560 -3940 6575 -3910
rect 6605 -3940 6620 -3910
rect 6560 -3980 6620 -3940
rect 6560 -4010 6575 -3980
rect 6605 -4010 6620 -3980
rect 6560 -4045 6620 -4010
rect 6560 -4075 6575 -4045
rect 6605 -4075 6620 -4045
rect 6560 -4105 6620 -4075
rect 6560 -4135 6575 -4105
rect 6605 -4135 6620 -4105
rect 6560 -4170 6620 -4135
rect 6560 -4200 6575 -4170
rect 6605 -4200 6620 -4170
rect 6560 -4240 6620 -4200
rect 6560 -4270 6575 -4240
rect 6605 -4270 6620 -4240
rect 6560 -4310 6620 -4270
rect 6560 -4340 6575 -4310
rect 6605 -4340 6620 -4310
rect 6560 -4380 6620 -4340
rect 6560 -4410 6575 -4380
rect 6605 -4410 6620 -4380
rect 6560 -4445 6620 -4410
rect 6560 -4475 6575 -4445
rect 6605 -4475 6620 -4445
rect 6560 -4490 6620 -4475
rect 6910 -1305 6970 -1290
rect 6910 -1335 6925 -1305
rect 6955 -1335 6970 -1305
rect 6910 -1370 6970 -1335
rect 6910 -1400 6925 -1370
rect 6955 -1400 6970 -1370
rect 6910 -1440 6970 -1400
rect 6910 -1470 6925 -1440
rect 6955 -1470 6970 -1440
rect 6910 -1510 6970 -1470
rect 6910 -1540 6925 -1510
rect 6955 -1540 6970 -1510
rect 6910 -1580 6970 -1540
rect 6910 -1610 6925 -1580
rect 6955 -1610 6970 -1580
rect 6910 -1645 6970 -1610
rect 6910 -1675 6925 -1645
rect 6955 -1675 6970 -1645
rect 6910 -1705 6970 -1675
rect 6910 -1735 6925 -1705
rect 6955 -1735 6970 -1705
rect 6910 -1770 6970 -1735
rect 6910 -1800 6925 -1770
rect 6955 -1800 6970 -1770
rect 6910 -1840 6970 -1800
rect 6910 -1870 6925 -1840
rect 6955 -1870 6970 -1840
rect 6910 -1910 6970 -1870
rect 6910 -1940 6925 -1910
rect 6955 -1940 6970 -1910
rect 6910 -1980 6970 -1940
rect 6910 -2010 6925 -1980
rect 6955 -2010 6970 -1980
rect 6910 -2045 6970 -2010
rect 6910 -2075 6925 -2045
rect 6955 -2075 6970 -2045
rect 6910 -2105 6970 -2075
rect 6910 -2135 6925 -2105
rect 6955 -2135 6970 -2105
rect 6910 -2170 6970 -2135
rect 6910 -2200 6925 -2170
rect 6955 -2200 6970 -2170
rect 6910 -2240 6970 -2200
rect 6910 -2270 6925 -2240
rect 6955 -2270 6970 -2240
rect 6910 -2310 6970 -2270
rect 6910 -2340 6925 -2310
rect 6955 -2340 6970 -2310
rect 6910 -2380 6970 -2340
rect 6910 -2410 6925 -2380
rect 6955 -2410 6970 -2380
rect 6910 -2445 6970 -2410
rect 6910 -2475 6925 -2445
rect 6955 -2475 6970 -2445
rect 6910 -2505 6970 -2475
rect 6910 -2535 6925 -2505
rect 6955 -2535 6970 -2505
rect 6910 -2570 6970 -2535
rect 6910 -2600 6925 -2570
rect 6955 -2600 6970 -2570
rect 6910 -2640 6970 -2600
rect 6910 -2670 6925 -2640
rect 6955 -2670 6970 -2640
rect 6910 -2710 6970 -2670
rect 6910 -2740 6925 -2710
rect 6955 -2740 6970 -2710
rect 6910 -2780 6970 -2740
rect 6910 -2810 6925 -2780
rect 6955 -2810 6970 -2780
rect 6910 -2845 6970 -2810
rect 6910 -2875 6925 -2845
rect 6955 -2875 6970 -2845
rect 6910 -2905 6970 -2875
rect 6910 -2935 6925 -2905
rect 6955 -2935 6970 -2905
rect 6910 -2970 6970 -2935
rect 6910 -3000 6925 -2970
rect 6955 -3000 6970 -2970
rect 6910 -3040 6970 -3000
rect 6910 -3070 6925 -3040
rect 6955 -3070 6970 -3040
rect 6910 -3110 6970 -3070
rect 6910 -3140 6925 -3110
rect 6955 -3140 6970 -3110
rect 6910 -3180 6970 -3140
rect 6910 -3210 6925 -3180
rect 6955 -3210 6970 -3180
rect 6910 -3245 6970 -3210
rect 6910 -3275 6925 -3245
rect 6955 -3275 6970 -3245
rect 6910 -3305 6970 -3275
rect 6910 -3335 6925 -3305
rect 6955 -3335 6970 -3305
rect 6910 -3370 6970 -3335
rect 6910 -3400 6925 -3370
rect 6955 -3400 6970 -3370
rect 6910 -3440 6970 -3400
rect 6910 -3470 6925 -3440
rect 6955 -3470 6970 -3440
rect 6910 -3510 6970 -3470
rect 6910 -3540 6925 -3510
rect 6955 -3540 6970 -3510
rect 6910 -3580 6970 -3540
rect 6910 -3610 6925 -3580
rect 6955 -3610 6970 -3580
rect 6910 -3645 6970 -3610
rect 6910 -3675 6925 -3645
rect 6955 -3675 6970 -3645
rect 6910 -3705 6970 -3675
rect 6910 -3735 6925 -3705
rect 6955 -3735 6970 -3705
rect 6910 -3770 6970 -3735
rect 6910 -3800 6925 -3770
rect 6955 -3800 6970 -3770
rect 6910 -3840 6970 -3800
rect 6910 -3870 6925 -3840
rect 6955 -3870 6970 -3840
rect 6910 -3910 6970 -3870
rect 6910 -3940 6925 -3910
rect 6955 -3940 6970 -3910
rect 6910 -3980 6970 -3940
rect 6910 -4010 6925 -3980
rect 6955 -4010 6970 -3980
rect 6910 -4045 6970 -4010
rect 6910 -4075 6925 -4045
rect 6955 -4075 6970 -4045
rect 6910 -4105 6970 -4075
rect 6910 -4135 6925 -4105
rect 6955 -4135 6970 -4105
rect 6910 -4170 6970 -4135
rect 6910 -4200 6925 -4170
rect 6955 -4200 6970 -4170
rect 6910 -4240 6970 -4200
rect 6910 -4270 6925 -4240
rect 6955 -4270 6970 -4240
rect 6910 -4310 6970 -4270
rect 6910 -4340 6925 -4310
rect 6955 -4340 6970 -4310
rect 6910 -4380 6970 -4340
rect 6910 -4410 6925 -4380
rect 6955 -4410 6970 -4380
rect 6910 -4445 6970 -4410
rect 6910 -4475 6925 -4445
rect 6955 -4475 6970 -4445
rect 6910 -4490 6970 -4475
rect 7260 -1305 7320 -1290
rect 7260 -1335 7275 -1305
rect 7305 -1335 7320 -1305
rect 7260 -1370 7320 -1335
rect 7260 -1400 7275 -1370
rect 7305 -1400 7320 -1370
rect 7260 -1440 7320 -1400
rect 7260 -1470 7275 -1440
rect 7305 -1470 7320 -1440
rect 7260 -1510 7320 -1470
rect 7260 -1540 7275 -1510
rect 7305 -1540 7320 -1510
rect 7260 -1580 7320 -1540
rect 7260 -1610 7275 -1580
rect 7305 -1610 7320 -1580
rect 7260 -1645 7320 -1610
rect 7260 -1675 7275 -1645
rect 7305 -1675 7320 -1645
rect 7260 -1705 7320 -1675
rect 7260 -1735 7275 -1705
rect 7305 -1735 7320 -1705
rect 7260 -1770 7320 -1735
rect 7260 -1800 7275 -1770
rect 7305 -1800 7320 -1770
rect 7260 -1840 7320 -1800
rect 7260 -1870 7275 -1840
rect 7305 -1870 7320 -1840
rect 7260 -1910 7320 -1870
rect 7260 -1940 7275 -1910
rect 7305 -1940 7320 -1910
rect 7260 -1980 7320 -1940
rect 7260 -2010 7275 -1980
rect 7305 -2010 7320 -1980
rect 7260 -2045 7320 -2010
rect 7260 -2075 7275 -2045
rect 7305 -2075 7320 -2045
rect 7260 -2105 7320 -2075
rect 7260 -2135 7275 -2105
rect 7305 -2135 7320 -2105
rect 7260 -2170 7320 -2135
rect 7260 -2200 7275 -2170
rect 7305 -2200 7320 -2170
rect 7260 -2240 7320 -2200
rect 7260 -2270 7275 -2240
rect 7305 -2270 7320 -2240
rect 7260 -2310 7320 -2270
rect 7260 -2340 7275 -2310
rect 7305 -2340 7320 -2310
rect 7260 -2380 7320 -2340
rect 7260 -2410 7275 -2380
rect 7305 -2410 7320 -2380
rect 7260 -2445 7320 -2410
rect 7260 -2475 7275 -2445
rect 7305 -2475 7320 -2445
rect 7260 -2505 7320 -2475
rect 7260 -2535 7275 -2505
rect 7305 -2535 7320 -2505
rect 7260 -2570 7320 -2535
rect 7260 -2600 7275 -2570
rect 7305 -2600 7320 -2570
rect 7260 -2640 7320 -2600
rect 7260 -2670 7275 -2640
rect 7305 -2670 7320 -2640
rect 7260 -2710 7320 -2670
rect 7260 -2740 7275 -2710
rect 7305 -2740 7320 -2710
rect 7260 -2780 7320 -2740
rect 7260 -2810 7275 -2780
rect 7305 -2810 7320 -2780
rect 7260 -2845 7320 -2810
rect 7260 -2875 7275 -2845
rect 7305 -2875 7320 -2845
rect 7260 -2905 7320 -2875
rect 7260 -2935 7275 -2905
rect 7305 -2935 7320 -2905
rect 7260 -2970 7320 -2935
rect 7260 -3000 7275 -2970
rect 7305 -3000 7320 -2970
rect 7260 -3040 7320 -3000
rect 7260 -3070 7275 -3040
rect 7305 -3070 7320 -3040
rect 7260 -3110 7320 -3070
rect 7260 -3140 7275 -3110
rect 7305 -3140 7320 -3110
rect 7260 -3180 7320 -3140
rect 7260 -3210 7275 -3180
rect 7305 -3210 7320 -3180
rect 7260 -3245 7320 -3210
rect 7260 -3275 7275 -3245
rect 7305 -3275 7320 -3245
rect 7260 -3305 7320 -3275
rect 7260 -3335 7275 -3305
rect 7305 -3335 7320 -3305
rect 7260 -3370 7320 -3335
rect 7260 -3400 7275 -3370
rect 7305 -3400 7320 -3370
rect 7260 -3440 7320 -3400
rect 7260 -3470 7275 -3440
rect 7305 -3470 7320 -3440
rect 7260 -3510 7320 -3470
rect 7260 -3540 7275 -3510
rect 7305 -3540 7320 -3510
rect 7260 -3580 7320 -3540
rect 7260 -3610 7275 -3580
rect 7305 -3610 7320 -3580
rect 7260 -3645 7320 -3610
rect 7260 -3675 7275 -3645
rect 7305 -3675 7320 -3645
rect 7260 -3705 7320 -3675
rect 7260 -3735 7275 -3705
rect 7305 -3735 7320 -3705
rect 7260 -3770 7320 -3735
rect 7260 -3800 7275 -3770
rect 7305 -3800 7320 -3770
rect 7260 -3840 7320 -3800
rect 7260 -3870 7275 -3840
rect 7305 -3870 7320 -3840
rect 7260 -3910 7320 -3870
rect 7260 -3940 7275 -3910
rect 7305 -3940 7320 -3910
rect 7260 -3980 7320 -3940
rect 7260 -4010 7275 -3980
rect 7305 -4010 7320 -3980
rect 7260 -4045 7320 -4010
rect 7260 -4075 7275 -4045
rect 7305 -4075 7320 -4045
rect 7260 -4105 7320 -4075
rect 7260 -4135 7275 -4105
rect 7305 -4135 7320 -4105
rect 7260 -4170 7320 -4135
rect 7260 -4200 7275 -4170
rect 7305 -4200 7320 -4170
rect 7260 -4240 7320 -4200
rect 7260 -4270 7275 -4240
rect 7305 -4270 7320 -4240
rect 7260 -4310 7320 -4270
rect 7260 -4340 7275 -4310
rect 7305 -4340 7320 -4310
rect 7260 -4380 7320 -4340
rect 7260 -4410 7275 -4380
rect 7305 -4410 7320 -4380
rect 7260 -4445 7320 -4410
rect 7260 -4475 7275 -4445
rect 7305 -4475 7320 -4445
rect 7260 -4490 7320 -4475
rect 7610 -1305 7670 -1290
rect 7610 -1335 7625 -1305
rect 7655 -1335 7670 -1305
rect 7610 -1370 7670 -1335
rect 7610 -1400 7625 -1370
rect 7655 -1400 7670 -1370
rect 7610 -1440 7670 -1400
rect 7610 -1470 7625 -1440
rect 7655 -1470 7670 -1440
rect 7610 -1510 7670 -1470
rect 7610 -1540 7625 -1510
rect 7655 -1540 7670 -1510
rect 7610 -1580 7670 -1540
rect 7610 -1610 7625 -1580
rect 7655 -1610 7670 -1580
rect 7610 -1645 7670 -1610
rect 7610 -1675 7625 -1645
rect 7655 -1675 7670 -1645
rect 7610 -1705 7670 -1675
rect 7610 -1735 7625 -1705
rect 7655 -1735 7670 -1705
rect 7610 -1770 7670 -1735
rect 7610 -1800 7625 -1770
rect 7655 -1800 7670 -1770
rect 7610 -1840 7670 -1800
rect 7610 -1870 7625 -1840
rect 7655 -1870 7670 -1840
rect 7610 -1910 7670 -1870
rect 7610 -1940 7625 -1910
rect 7655 -1940 7670 -1910
rect 7610 -1980 7670 -1940
rect 7610 -2010 7625 -1980
rect 7655 -2010 7670 -1980
rect 7610 -2045 7670 -2010
rect 7610 -2075 7625 -2045
rect 7655 -2075 7670 -2045
rect 7610 -2105 7670 -2075
rect 7610 -2135 7625 -2105
rect 7655 -2135 7670 -2105
rect 7610 -2170 7670 -2135
rect 7610 -2200 7625 -2170
rect 7655 -2200 7670 -2170
rect 7610 -2240 7670 -2200
rect 7610 -2270 7625 -2240
rect 7655 -2270 7670 -2240
rect 7610 -2310 7670 -2270
rect 7610 -2340 7625 -2310
rect 7655 -2340 7670 -2310
rect 7610 -2380 7670 -2340
rect 7610 -2410 7625 -2380
rect 7655 -2410 7670 -2380
rect 7610 -2445 7670 -2410
rect 7610 -2475 7625 -2445
rect 7655 -2475 7670 -2445
rect 7610 -2505 7670 -2475
rect 7610 -2535 7625 -2505
rect 7655 -2535 7670 -2505
rect 7610 -2570 7670 -2535
rect 7610 -2600 7625 -2570
rect 7655 -2600 7670 -2570
rect 7610 -2640 7670 -2600
rect 7610 -2670 7625 -2640
rect 7655 -2670 7670 -2640
rect 7610 -2710 7670 -2670
rect 7610 -2740 7625 -2710
rect 7655 -2740 7670 -2710
rect 7610 -2780 7670 -2740
rect 7610 -2810 7625 -2780
rect 7655 -2810 7670 -2780
rect 7610 -2845 7670 -2810
rect 7610 -2875 7625 -2845
rect 7655 -2875 7670 -2845
rect 7610 -2905 7670 -2875
rect 7610 -2935 7625 -2905
rect 7655 -2935 7670 -2905
rect 7610 -2970 7670 -2935
rect 7610 -3000 7625 -2970
rect 7655 -3000 7670 -2970
rect 7610 -3040 7670 -3000
rect 7610 -3070 7625 -3040
rect 7655 -3070 7670 -3040
rect 7610 -3110 7670 -3070
rect 7610 -3140 7625 -3110
rect 7655 -3140 7670 -3110
rect 7610 -3180 7670 -3140
rect 7610 -3210 7625 -3180
rect 7655 -3210 7670 -3180
rect 7610 -3245 7670 -3210
rect 7610 -3275 7625 -3245
rect 7655 -3275 7670 -3245
rect 7610 -3305 7670 -3275
rect 7610 -3335 7625 -3305
rect 7655 -3335 7670 -3305
rect 7610 -3370 7670 -3335
rect 7610 -3400 7625 -3370
rect 7655 -3400 7670 -3370
rect 7610 -3440 7670 -3400
rect 7610 -3470 7625 -3440
rect 7655 -3470 7670 -3440
rect 7610 -3510 7670 -3470
rect 7610 -3540 7625 -3510
rect 7655 -3540 7670 -3510
rect 7610 -3580 7670 -3540
rect 7610 -3610 7625 -3580
rect 7655 -3610 7670 -3580
rect 7610 -3645 7670 -3610
rect 7610 -3675 7625 -3645
rect 7655 -3675 7670 -3645
rect 7610 -3705 7670 -3675
rect 7610 -3735 7625 -3705
rect 7655 -3735 7670 -3705
rect 7610 -3770 7670 -3735
rect 7610 -3800 7625 -3770
rect 7655 -3800 7670 -3770
rect 7610 -3840 7670 -3800
rect 7610 -3870 7625 -3840
rect 7655 -3870 7670 -3840
rect 7610 -3910 7670 -3870
rect 7610 -3940 7625 -3910
rect 7655 -3940 7670 -3910
rect 7610 -3980 7670 -3940
rect 7610 -4010 7625 -3980
rect 7655 -4010 7670 -3980
rect 7610 -4045 7670 -4010
rect 7610 -4075 7625 -4045
rect 7655 -4075 7670 -4045
rect 7610 -4105 7670 -4075
rect 7610 -4135 7625 -4105
rect 7655 -4135 7670 -4105
rect 7610 -4170 7670 -4135
rect 7610 -4200 7625 -4170
rect 7655 -4200 7670 -4170
rect 7610 -4240 7670 -4200
rect 7610 -4270 7625 -4240
rect 7655 -4270 7670 -4240
rect 7610 -4310 7670 -4270
rect 7610 -4340 7625 -4310
rect 7655 -4340 7670 -4310
rect 7610 -4380 7670 -4340
rect 7610 -4410 7625 -4380
rect 7655 -4410 7670 -4380
rect 7610 -4445 7670 -4410
rect 7610 -4475 7625 -4445
rect 7655 -4475 7670 -4445
rect 7610 -4490 7670 -4475
rect 7960 -1305 8020 -1290
rect 7960 -1335 7975 -1305
rect 8005 -1335 8020 -1305
rect 7960 -1370 8020 -1335
rect 7960 -1400 7975 -1370
rect 8005 -1400 8020 -1370
rect 7960 -1440 8020 -1400
rect 7960 -1470 7975 -1440
rect 8005 -1470 8020 -1440
rect 7960 -1510 8020 -1470
rect 7960 -1540 7975 -1510
rect 8005 -1540 8020 -1510
rect 7960 -1580 8020 -1540
rect 7960 -1610 7975 -1580
rect 8005 -1610 8020 -1580
rect 7960 -1645 8020 -1610
rect 7960 -1675 7975 -1645
rect 8005 -1675 8020 -1645
rect 7960 -1705 8020 -1675
rect 7960 -1735 7975 -1705
rect 8005 -1735 8020 -1705
rect 7960 -1770 8020 -1735
rect 7960 -1800 7975 -1770
rect 8005 -1800 8020 -1770
rect 7960 -1840 8020 -1800
rect 7960 -1870 7975 -1840
rect 8005 -1870 8020 -1840
rect 7960 -1910 8020 -1870
rect 7960 -1940 7975 -1910
rect 8005 -1940 8020 -1910
rect 7960 -1980 8020 -1940
rect 7960 -2010 7975 -1980
rect 8005 -2010 8020 -1980
rect 7960 -2045 8020 -2010
rect 7960 -2075 7975 -2045
rect 8005 -2075 8020 -2045
rect 7960 -2105 8020 -2075
rect 7960 -2135 7975 -2105
rect 8005 -2135 8020 -2105
rect 7960 -2170 8020 -2135
rect 7960 -2200 7975 -2170
rect 8005 -2200 8020 -2170
rect 7960 -2240 8020 -2200
rect 7960 -2270 7975 -2240
rect 8005 -2270 8020 -2240
rect 7960 -2310 8020 -2270
rect 7960 -2340 7975 -2310
rect 8005 -2340 8020 -2310
rect 7960 -2380 8020 -2340
rect 7960 -2410 7975 -2380
rect 8005 -2410 8020 -2380
rect 7960 -2445 8020 -2410
rect 7960 -2475 7975 -2445
rect 8005 -2475 8020 -2445
rect 7960 -2505 8020 -2475
rect 7960 -2535 7975 -2505
rect 8005 -2535 8020 -2505
rect 7960 -2570 8020 -2535
rect 7960 -2600 7975 -2570
rect 8005 -2600 8020 -2570
rect 7960 -2640 8020 -2600
rect 7960 -2670 7975 -2640
rect 8005 -2670 8020 -2640
rect 7960 -2710 8020 -2670
rect 7960 -2740 7975 -2710
rect 8005 -2740 8020 -2710
rect 7960 -2780 8020 -2740
rect 7960 -2810 7975 -2780
rect 8005 -2810 8020 -2780
rect 7960 -2845 8020 -2810
rect 7960 -2875 7975 -2845
rect 8005 -2875 8020 -2845
rect 7960 -2905 8020 -2875
rect 7960 -2935 7975 -2905
rect 8005 -2935 8020 -2905
rect 7960 -2970 8020 -2935
rect 7960 -3000 7975 -2970
rect 8005 -3000 8020 -2970
rect 7960 -3040 8020 -3000
rect 7960 -3070 7975 -3040
rect 8005 -3070 8020 -3040
rect 7960 -3110 8020 -3070
rect 7960 -3140 7975 -3110
rect 8005 -3140 8020 -3110
rect 7960 -3180 8020 -3140
rect 7960 -3210 7975 -3180
rect 8005 -3210 8020 -3180
rect 7960 -3245 8020 -3210
rect 7960 -3275 7975 -3245
rect 8005 -3275 8020 -3245
rect 7960 -3305 8020 -3275
rect 7960 -3335 7975 -3305
rect 8005 -3335 8020 -3305
rect 7960 -3370 8020 -3335
rect 7960 -3400 7975 -3370
rect 8005 -3400 8020 -3370
rect 7960 -3440 8020 -3400
rect 7960 -3470 7975 -3440
rect 8005 -3470 8020 -3440
rect 7960 -3510 8020 -3470
rect 7960 -3540 7975 -3510
rect 8005 -3540 8020 -3510
rect 7960 -3580 8020 -3540
rect 7960 -3610 7975 -3580
rect 8005 -3610 8020 -3580
rect 7960 -3645 8020 -3610
rect 7960 -3675 7975 -3645
rect 8005 -3675 8020 -3645
rect 7960 -3705 8020 -3675
rect 7960 -3735 7975 -3705
rect 8005 -3735 8020 -3705
rect 7960 -3770 8020 -3735
rect 7960 -3800 7975 -3770
rect 8005 -3800 8020 -3770
rect 7960 -3840 8020 -3800
rect 7960 -3870 7975 -3840
rect 8005 -3870 8020 -3840
rect 7960 -3910 8020 -3870
rect 7960 -3940 7975 -3910
rect 8005 -3940 8020 -3910
rect 7960 -3980 8020 -3940
rect 7960 -4010 7975 -3980
rect 8005 -4010 8020 -3980
rect 7960 -4045 8020 -4010
rect 7960 -4075 7975 -4045
rect 8005 -4075 8020 -4045
rect 7960 -4105 8020 -4075
rect 7960 -4135 7975 -4105
rect 8005 -4135 8020 -4105
rect 7960 -4170 8020 -4135
rect 7960 -4200 7975 -4170
rect 8005 -4200 8020 -4170
rect 7960 -4240 8020 -4200
rect 7960 -4270 7975 -4240
rect 8005 -4270 8020 -4240
rect 7960 -4310 8020 -4270
rect 7960 -4340 7975 -4310
rect 8005 -4340 8020 -4310
rect 7960 -4380 8020 -4340
rect 7960 -4410 7975 -4380
rect 8005 -4410 8020 -4380
rect 7960 -4445 8020 -4410
rect 7960 -4475 7975 -4445
rect 8005 -4475 8020 -4445
rect 7960 -4490 8020 -4475
rect 8310 -1305 8370 -1290
rect 8310 -1335 8325 -1305
rect 8355 -1335 8370 -1305
rect 8310 -1370 8370 -1335
rect 8310 -1400 8325 -1370
rect 8355 -1400 8370 -1370
rect 8310 -1440 8370 -1400
rect 8310 -1470 8325 -1440
rect 8355 -1470 8370 -1440
rect 8310 -1510 8370 -1470
rect 8310 -1540 8325 -1510
rect 8355 -1540 8370 -1510
rect 8310 -1580 8370 -1540
rect 8310 -1610 8325 -1580
rect 8355 -1610 8370 -1580
rect 8310 -1645 8370 -1610
rect 8310 -1675 8325 -1645
rect 8355 -1675 8370 -1645
rect 8310 -1705 8370 -1675
rect 8310 -1735 8325 -1705
rect 8355 -1735 8370 -1705
rect 8310 -1770 8370 -1735
rect 8310 -1800 8325 -1770
rect 8355 -1800 8370 -1770
rect 8310 -1840 8370 -1800
rect 8310 -1870 8325 -1840
rect 8355 -1870 8370 -1840
rect 8310 -1910 8370 -1870
rect 8310 -1940 8325 -1910
rect 8355 -1940 8370 -1910
rect 8310 -1980 8370 -1940
rect 8310 -2010 8325 -1980
rect 8355 -2010 8370 -1980
rect 8310 -2045 8370 -2010
rect 8310 -2075 8325 -2045
rect 8355 -2075 8370 -2045
rect 8310 -2105 8370 -2075
rect 8310 -2135 8325 -2105
rect 8355 -2135 8370 -2105
rect 8310 -2170 8370 -2135
rect 8310 -2200 8325 -2170
rect 8355 -2200 8370 -2170
rect 8310 -2240 8370 -2200
rect 8310 -2270 8325 -2240
rect 8355 -2270 8370 -2240
rect 8310 -2310 8370 -2270
rect 8310 -2340 8325 -2310
rect 8355 -2340 8370 -2310
rect 8310 -2380 8370 -2340
rect 8310 -2410 8325 -2380
rect 8355 -2410 8370 -2380
rect 8310 -2445 8370 -2410
rect 8310 -2475 8325 -2445
rect 8355 -2475 8370 -2445
rect 8310 -2505 8370 -2475
rect 8310 -2535 8325 -2505
rect 8355 -2535 8370 -2505
rect 8310 -2570 8370 -2535
rect 8310 -2600 8325 -2570
rect 8355 -2600 8370 -2570
rect 8310 -2640 8370 -2600
rect 8310 -2670 8325 -2640
rect 8355 -2670 8370 -2640
rect 8310 -2710 8370 -2670
rect 8310 -2740 8325 -2710
rect 8355 -2740 8370 -2710
rect 8310 -2780 8370 -2740
rect 8310 -2810 8325 -2780
rect 8355 -2810 8370 -2780
rect 8310 -2845 8370 -2810
rect 8310 -2875 8325 -2845
rect 8355 -2875 8370 -2845
rect 8310 -2905 8370 -2875
rect 8310 -2935 8325 -2905
rect 8355 -2935 8370 -2905
rect 8310 -2970 8370 -2935
rect 8310 -3000 8325 -2970
rect 8355 -3000 8370 -2970
rect 8310 -3040 8370 -3000
rect 8310 -3070 8325 -3040
rect 8355 -3070 8370 -3040
rect 8310 -3110 8370 -3070
rect 8310 -3140 8325 -3110
rect 8355 -3140 8370 -3110
rect 8310 -3180 8370 -3140
rect 8310 -3210 8325 -3180
rect 8355 -3210 8370 -3180
rect 8310 -3245 8370 -3210
rect 8310 -3275 8325 -3245
rect 8355 -3275 8370 -3245
rect 8310 -3305 8370 -3275
rect 8310 -3335 8325 -3305
rect 8355 -3335 8370 -3305
rect 8310 -3370 8370 -3335
rect 8310 -3400 8325 -3370
rect 8355 -3400 8370 -3370
rect 8310 -3440 8370 -3400
rect 8310 -3470 8325 -3440
rect 8355 -3470 8370 -3440
rect 8310 -3510 8370 -3470
rect 8310 -3540 8325 -3510
rect 8355 -3540 8370 -3510
rect 8310 -3580 8370 -3540
rect 8310 -3610 8325 -3580
rect 8355 -3610 8370 -3580
rect 8310 -3645 8370 -3610
rect 8310 -3675 8325 -3645
rect 8355 -3675 8370 -3645
rect 8310 -3705 8370 -3675
rect 8310 -3735 8325 -3705
rect 8355 -3735 8370 -3705
rect 8310 -3770 8370 -3735
rect 8310 -3800 8325 -3770
rect 8355 -3800 8370 -3770
rect 8310 -3840 8370 -3800
rect 8310 -3870 8325 -3840
rect 8355 -3870 8370 -3840
rect 8310 -3910 8370 -3870
rect 8310 -3940 8325 -3910
rect 8355 -3940 8370 -3910
rect 8310 -3980 8370 -3940
rect 8310 -4010 8325 -3980
rect 8355 -4010 8370 -3980
rect 8310 -4045 8370 -4010
rect 8310 -4075 8325 -4045
rect 8355 -4075 8370 -4045
rect 8310 -4105 8370 -4075
rect 8310 -4135 8325 -4105
rect 8355 -4135 8370 -4105
rect 8310 -4170 8370 -4135
rect 8310 -4200 8325 -4170
rect 8355 -4200 8370 -4170
rect 8310 -4240 8370 -4200
rect 8310 -4270 8325 -4240
rect 8355 -4270 8370 -4240
rect 8310 -4310 8370 -4270
rect 8310 -4340 8325 -4310
rect 8355 -4340 8370 -4310
rect 8310 -4380 8370 -4340
rect 8310 -4410 8325 -4380
rect 8355 -4410 8370 -4380
rect 8310 -4445 8370 -4410
rect 8310 -4475 8325 -4445
rect 8355 -4475 8370 -4445
rect 8310 -4490 8370 -4475
rect 8660 -1305 8720 -1290
rect 8660 -1335 8675 -1305
rect 8705 -1335 8720 -1305
rect 8660 -1370 8720 -1335
rect 8660 -1400 8675 -1370
rect 8705 -1400 8720 -1370
rect 8660 -1440 8720 -1400
rect 8660 -1470 8675 -1440
rect 8705 -1470 8720 -1440
rect 8660 -1510 8720 -1470
rect 8660 -1540 8675 -1510
rect 8705 -1540 8720 -1510
rect 8660 -1580 8720 -1540
rect 8660 -1610 8675 -1580
rect 8705 -1610 8720 -1580
rect 8660 -1645 8720 -1610
rect 8660 -1675 8675 -1645
rect 8705 -1675 8720 -1645
rect 8660 -1705 8720 -1675
rect 8660 -1735 8675 -1705
rect 8705 -1735 8720 -1705
rect 8660 -1770 8720 -1735
rect 8660 -1800 8675 -1770
rect 8705 -1800 8720 -1770
rect 8660 -1840 8720 -1800
rect 8660 -1870 8675 -1840
rect 8705 -1870 8720 -1840
rect 8660 -1910 8720 -1870
rect 8660 -1940 8675 -1910
rect 8705 -1940 8720 -1910
rect 8660 -1980 8720 -1940
rect 8660 -2010 8675 -1980
rect 8705 -2010 8720 -1980
rect 8660 -2045 8720 -2010
rect 8660 -2075 8675 -2045
rect 8705 -2075 8720 -2045
rect 8660 -2105 8720 -2075
rect 8660 -2135 8675 -2105
rect 8705 -2135 8720 -2105
rect 8660 -2170 8720 -2135
rect 8660 -2200 8675 -2170
rect 8705 -2200 8720 -2170
rect 8660 -2240 8720 -2200
rect 8660 -2270 8675 -2240
rect 8705 -2270 8720 -2240
rect 8660 -2310 8720 -2270
rect 8660 -2340 8675 -2310
rect 8705 -2340 8720 -2310
rect 8660 -2380 8720 -2340
rect 8660 -2410 8675 -2380
rect 8705 -2410 8720 -2380
rect 8660 -2445 8720 -2410
rect 8660 -2475 8675 -2445
rect 8705 -2475 8720 -2445
rect 8660 -2505 8720 -2475
rect 8660 -2535 8675 -2505
rect 8705 -2535 8720 -2505
rect 8660 -2570 8720 -2535
rect 8660 -2600 8675 -2570
rect 8705 -2600 8720 -2570
rect 8660 -2640 8720 -2600
rect 8660 -2670 8675 -2640
rect 8705 -2670 8720 -2640
rect 8660 -2710 8720 -2670
rect 8660 -2740 8675 -2710
rect 8705 -2740 8720 -2710
rect 8660 -2780 8720 -2740
rect 8660 -2810 8675 -2780
rect 8705 -2810 8720 -2780
rect 8660 -2845 8720 -2810
rect 8660 -2875 8675 -2845
rect 8705 -2875 8720 -2845
rect 8660 -2905 8720 -2875
rect 8660 -2935 8675 -2905
rect 8705 -2935 8720 -2905
rect 8660 -2970 8720 -2935
rect 8660 -3000 8675 -2970
rect 8705 -3000 8720 -2970
rect 8660 -3040 8720 -3000
rect 8660 -3070 8675 -3040
rect 8705 -3070 8720 -3040
rect 8660 -3110 8720 -3070
rect 8660 -3140 8675 -3110
rect 8705 -3140 8720 -3110
rect 8660 -3180 8720 -3140
rect 8660 -3210 8675 -3180
rect 8705 -3210 8720 -3180
rect 8660 -3245 8720 -3210
rect 8660 -3275 8675 -3245
rect 8705 -3275 8720 -3245
rect 8660 -3305 8720 -3275
rect 8660 -3335 8675 -3305
rect 8705 -3335 8720 -3305
rect 8660 -3370 8720 -3335
rect 8660 -3400 8675 -3370
rect 8705 -3400 8720 -3370
rect 8660 -3440 8720 -3400
rect 8660 -3470 8675 -3440
rect 8705 -3470 8720 -3440
rect 8660 -3510 8720 -3470
rect 8660 -3540 8675 -3510
rect 8705 -3540 8720 -3510
rect 8660 -3580 8720 -3540
rect 8660 -3610 8675 -3580
rect 8705 -3610 8720 -3580
rect 8660 -3645 8720 -3610
rect 8660 -3675 8675 -3645
rect 8705 -3675 8720 -3645
rect 8660 -3705 8720 -3675
rect 8660 -3735 8675 -3705
rect 8705 -3735 8720 -3705
rect 8660 -3770 8720 -3735
rect 8660 -3800 8675 -3770
rect 8705 -3800 8720 -3770
rect 8660 -3840 8720 -3800
rect 8660 -3870 8675 -3840
rect 8705 -3870 8720 -3840
rect 8660 -3910 8720 -3870
rect 8660 -3940 8675 -3910
rect 8705 -3940 8720 -3910
rect 8660 -3980 8720 -3940
rect 8660 -4010 8675 -3980
rect 8705 -4010 8720 -3980
rect 8660 -4045 8720 -4010
rect 8660 -4075 8675 -4045
rect 8705 -4075 8720 -4045
rect 8660 -4105 8720 -4075
rect 8660 -4135 8675 -4105
rect 8705 -4135 8720 -4105
rect 8660 -4170 8720 -4135
rect 8660 -4200 8675 -4170
rect 8705 -4200 8720 -4170
rect 8660 -4240 8720 -4200
rect 8660 -4270 8675 -4240
rect 8705 -4270 8720 -4240
rect 8660 -4310 8720 -4270
rect 8660 -4340 8675 -4310
rect 8705 -4340 8720 -4310
rect 8660 -4380 8720 -4340
rect 8660 -4410 8675 -4380
rect 8705 -4410 8720 -4380
rect 8660 -4445 8720 -4410
rect 8660 -4475 8675 -4445
rect 8705 -4475 8720 -4445
rect 8660 -4490 8720 -4475
<< via2 >>
rect 2335 20880 2365 20910
rect 2335 20815 2365 20845
rect 2335 20745 2365 20775
rect 2335 20675 2365 20705
rect 2335 20605 2365 20635
rect 2335 20540 2365 20570
rect 2335 20480 2365 20510
rect 2335 20415 2365 20445
rect 2335 20345 2365 20375
rect 2335 20275 2365 20305
rect 2335 20205 2365 20235
rect 2335 20140 2365 20170
rect 2335 20080 2365 20110
rect 2335 20015 2365 20045
rect 2335 19945 2365 19975
rect 2335 19875 2365 19905
rect 2335 19805 2365 19835
rect 2335 19740 2365 19770
rect 2335 19680 2365 19710
rect 2335 19615 2365 19645
rect 2335 19545 2365 19575
rect 2335 19475 2365 19505
rect 2335 19405 2365 19435
rect 2335 19340 2365 19370
rect 2335 19280 2365 19310
rect 2335 19215 2365 19245
rect 2335 19145 2365 19175
rect 2335 19075 2365 19105
rect 2335 19005 2365 19035
rect 2335 18940 2365 18970
rect 2335 18880 2365 18910
rect 2335 18815 2365 18845
rect 2335 18745 2365 18775
rect 2335 18675 2365 18705
rect 2335 18605 2365 18635
rect 2335 18540 2365 18570
rect 2335 18480 2365 18510
rect 2335 18415 2365 18445
rect 2335 18345 2365 18375
rect 2335 18275 2365 18305
rect 2335 18205 2365 18235
rect 2335 18140 2365 18170
rect 2335 18080 2365 18110
rect 2335 18015 2365 18045
rect 2335 17945 2365 17975
rect 2335 17875 2365 17905
rect 2335 17805 2365 17835
rect 2335 17740 2365 17770
rect 6705 20880 6735 20910
rect 6705 20815 6735 20845
rect 6705 20745 6735 20775
rect 6705 20675 6735 20705
rect 6705 20605 6735 20635
rect 6705 20540 6735 20570
rect 6705 20480 6735 20510
rect 6705 20415 6735 20445
rect 6705 20345 6735 20375
rect 6705 20275 6735 20305
rect 6705 20205 6735 20235
rect 6705 20140 6735 20170
rect 6705 20080 6735 20110
rect 6705 20015 6735 20045
rect 6705 19945 6735 19975
rect 6705 19875 6735 19905
rect 6705 19805 6735 19835
rect 6705 19740 6735 19770
rect 6705 19680 6735 19710
rect 6705 19615 6735 19645
rect 6705 19545 6735 19575
rect 6705 19475 6735 19505
rect 6705 19405 6735 19435
rect 6705 19340 6735 19370
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 2060 10055 2090 10085
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 1325 8065 1355 8095
rect 1325 8005 1355 8035
rect 1325 7940 1355 7970
rect 1325 7870 1355 7900
rect 1325 7800 1355 7830
rect 1325 7730 1355 7760
rect 1325 7665 1355 7695
rect 1325 7605 1355 7635
rect 1325 7540 1355 7570
rect 1325 7470 1355 7500
rect 1325 7400 1355 7430
rect 1325 7330 1355 7360
rect 1325 7265 1355 7295
rect 1325 7205 1355 7235
rect 1325 7140 1355 7170
rect 1325 7070 1355 7100
rect 1325 7000 1355 7030
rect 1325 6930 1355 6960
rect 1325 6865 1355 6895
rect 1325 6805 1355 6835
rect 1325 6740 1355 6770
rect 1325 6670 1355 6700
rect 1325 6600 1355 6630
rect 1325 6530 1355 6560
rect 1325 6465 1355 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 2390 9605 2420 9635
rect 2390 9540 2420 9570
rect 2390 9470 2420 9500
rect 2390 9400 2420 9430
rect 2390 9330 2420 9360
rect 2390 9265 2420 9295
rect 2390 9205 2420 9235
rect 2390 9140 2420 9170
rect 2390 9070 2420 9100
rect 2390 9000 2420 9030
rect 2390 8930 2420 8960
rect 2390 8865 2420 8895
rect 2390 8805 2420 8835
rect 2390 8740 2420 8770
rect 2390 8670 2420 8700
rect 2390 8600 2420 8630
rect 2390 8530 2420 8560
rect 2390 8465 2420 8495
rect 2390 8405 2420 8435
rect 2390 8340 2420 8370
rect 2390 8270 2420 8300
rect 2390 8200 2420 8230
rect 2390 8130 2420 8160
rect 2390 8065 2420 8095
rect 2390 8005 2420 8035
rect 2390 7940 2420 7970
rect 2390 7870 2420 7900
rect 2390 7800 2420 7830
rect 2390 7730 2420 7760
rect 2390 7665 2420 7695
rect 2390 7605 2420 7635
rect 2390 7540 2420 7570
rect 2390 7470 2420 7500
rect 2390 7400 2420 7430
rect 2390 7330 2420 7360
rect 2390 7265 2420 7295
rect 2390 7205 2420 7235
rect 2390 7140 2420 7170
rect 2390 7070 2420 7100
rect 2390 7000 2420 7030
rect 2390 6930 2420 6960
rect 2390 6865 2420 6895
rect 2390 6805 2420 6835
rect 2390 6740 2420 6770
rect 2390 6670 2420 6700
rect 2390 6600 2420 6630
rect 2390 6530 2420 6560
rect 2390 6465 2420 6495
rect 3240 9605 3270 9635
rect 3240 9540 3270 9570
rect 3240 9470 3270 9500
rect 3240 9400 3270 9430
rect 3240 9330 3270 9360
rect 3240 9265 3270 9295
rect 3240 9205 3270 9235
rect 3240 9140 3270 9170
rect 3240 9070 3270 9100
rect 3240 9000 3270 9030
rect 3240 8930 3270 8960
rect 3240 8865 3270 8895
rect 3240 8805 3270 8835
rect 3240 8740 3270 8770
rect 3240 8670 3270 8700
rect 3240 8600 3270 8630
rect 3240 8530 3270 8560
rect 3240 8465 3270 8495
rect 3240 8405 3270 8435
rect 3240 8340 3270 8370
rect 3240 8270 3270 8300
rect 3240 8200 3270 8230
rect 3240 8130 3270 8160
rect 3240 8065 3270 8095
rect 3240 8005 3270 8035
rect 3240 7940 3270 7970
rect 3240 7870 3270 7900
rect 3240 7800 3270 7830
rect 3240 7730 3270 7760
rect 3240 7665 3270 7695
rect 3240 7605 3270 7635
rect 3240 7540 3270 7570
rect 3240 7470 3270 7500
rect 3240 7400 3270 7430
rect 3240 7330 3270 7360
rect 3240 7265 3270 7295
rect 3240 7205 3270 7235
rect 3240 7140 3270 7170
rect 3240 7070 3270 7100
rect 3240 7000 3270 7030
rect 3240 6930 3270 6960
rect 3240 6865 3270 6895
rect 3240 6805 3270 6835
rect 3240 6740 3270 6770
rect 3240 6670 3270 6700
rect 3240 6600 3270 6630
rect 3240 6530 3270 6560
rect 3240 6465 3270 6495
rect 5650 9605 5680 9635
rect 5650 9540 5680 9570
rect 5650 9470 5680 9500
rect 5650 9400 5680 9430
rect 5650 9330 5680 9360
rect 5650 9265 5680 9295
rect 5650 9205 5680 9235
rect 5650 9140 5680 9170
rect 5650 9070 5680 9100
rect 5650 9000 5680 9030
rect 5650 8930 5680 8960
rect 5650 8865 5680 8895
rect 5650 8805 5680 8835
rect 5650 8740 5680 8770
rect 5650 8670 5680 8700
rect 5650 8600 5680 8630
rect 5650 8530 5680 8560
rect 5650 8465 5680 8495
rect 5650 8405 5680 8435
rect 5650 8340 5680 8370
rect 5650 8270 5680 8300
rect 5650 8200 5680 8230
rect 5650 8130 5680 8160
rect 5650 8065 5680 8095
rect 5650 8005 5680 8035
rect 5650 7940 5680 7970
rect 5650 7870 5680 7900
rect 5650 7800 5680 7830
rect 5650 7730 5680 7760
rect 5650 7665 5680 7695
rect 5650 7605 5680 7635
rect 5650 7540 5680 7570
rect 5650 7470 5680 7500
rect 5650 7400 5680 7430
rect 5650 7330 5680 7360
rect 5650 7265 5680 7295
rect 5650 7205 5680 7235
rect 5650 7140 5680 7170
rect 5650 7070 5680 7100
rect 5650 7000 5680 7030
rect 5650 6930 5680 6960
rect 5650 6865 5680 6895
rect 5650 6805 5680 6835
rect 5650 6740 5680 6770
rect 5650 6670 5680 6700
rect 5650 6600 5680 6630
rect 5650 6530 5680 6560
rect 5650 6465 5680 6495
rect 6305 9605 6335 9635
rect 6305 9540 6335 9570
rect 6305 9470 6335 9500
rect 6305 9400 6335 9430
rect 6305 9330 6335 9360
rect 6305 9265 6335 9295
rect 6305 9205 6335 9235
rect 6305 9140 6335 9170
rect 6305 9070 6335 9100
rect 6305 9000 6335 9030
rect 6305 8930 6335 8960
rect 6305 8865 6335 8895
rect 6305 8805 6335 8835
rect 6305 8740 6335 8770
rect 6305 8670 6335 8700
rect 6305 8600 6335 8630
rect 6305 8530 6335 8560
rect 6305 8465 6335 8495
rect 6305 8405 6335 8435
rect 6305 8340 6335 8370
rect 6305 8270 6335 8300
rect 6305 8200 6335 8230
rect 6305 8130 6335 8160
rect 6305 8065 6335 8095
rect 6305 8005 6335 8035
rect 6305 7940 6335 7970
rect 6305 7870 6335 7900
rect 6305 7800 6335 7830
rect 6305 7730 6335 7760
rect 6305 7665 6335 7695
rect 6305 7605 6335 7635
rect 6305 7540 6335 7570
rect 6305 7470 6335 7500
rect 6305 7400 6335 7430
rect 6305 7330 6335 7360
rect 6305 7265 6335 7295
rect 6305 7205 6335 7235
rect 6305 7140 6335 7170
rect 6305 7070 6335 7100
rect 6305 7000 6335 7030
rect 6305 6930 6335 6960
rect 6305 6865 6335 6895
rect 6305 6805 6335 6835
rect 6305 6740 6335 6770
rect 6305 6670 6335 6700
rect 6305 6600 6335 6630
rect 6305 6530 6335 6560
rect 6305 6465 6335 6495
rect 6595 9605 6625 9635
rect 6595 9540 6625 9570
rect 6595 9470 6625 9500
rect 6595 9400 6625 9430
rect 6595 9330 6625 9360
rect 6595 9265 6625 9295
rect 6595 9205 6625 9235
rect 6595 9140 6625 9170
rect 6595 9070 6625 9100
rect 6595 9000 6625 9030
rect 6595 8930 6625 8960
rect 6595 8865 6625 8895
rect 6595 8805 6625 8835
rect 6595 8740 6625 8770
rect 6595 8670 6625 8700
rect 6595 8600 6625 8630
rect 6595 8530 6625 8560
rect 6595 8465 6625 8495
rect 6595 8405 6625 8435
rect 6595 8340 6625 8370
rect 6595 8270 6625 8300
rect 6595 8200 6625 8230
rect 6595 8130 6625 8160
rect 6595 8065 6625 8095
rect 6595 8005 6625 8035
rect 6595 7940 6625 7970
rect 6595 7870 6625 7900
rect 6595 7800 6625 7830
rect 6595 7730 6625 7760
rect 6595 7665 6625 7695
rect 6595 7605 6625 7635
rect 6595 7540 6625 7570
rect 6595 7470 6625 7500
rect 6595 7400 6625 7430
rect 6595 7330 6625 7360
rect 6595 7265 6625 7295
rect 6595 7205 6625 7235
rect 6595 7140 6625 7170
rect 6595 7070 6625 7100
rect 6595 7000 6625 7030
rect 6595 6930 6625 6960
rect 6595 6865 6625 6895
rect 6595 6805 6625 6835
rect 6595 6740 6625 6770
rect 6595 6670 6625 6700
rect 6595 6600 6625 6630
rect 6595 6530 6625 6560
rect 6595 6465 6625 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect 7625 8065 7655 8095
rect 7625 8005 7655 8035
rect 7625 7940 7655 7970
rect 7625 7870 7655 7900
rect 7625 7800 7655 7830
rect 7625 7730 7655 7760
rect 7625 7665 7655 7695
rect 7625 7605 7655 7635
rect 7625 7540 7655 7570
rect 7625 7470 7655 7500
rect 7625 7400 7655 7430
rect 7625 7330 7655 7360
rect 7625 7265 7655 7295
rect 7625 7205 7655 7235
rect 7625 7140 7655 7170
rect 7625 7070 7655 7100
rect 7625 7000 7655 7030
rect 7625 6930 7655 6960
rect 7625 6865 7655 6895
rect 7625 6805 7655 6835
rect 7625 6740 7655 6770
rect 7625 6670 7655 6700
rect 7625 6600 7655 6630
rect 7625 6530 7655 6560
rect 7625 6465 7655 6495
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect -75 -2935 -45 -2905
rect -75 -3000 -45 -2970
rect -75 -3070 -45 -3040
rect -75 -3140 -45 -3110
rect -75 -3210 -45 -3180
rect -75 -3275 -45 -3245
rect -75 -3335 -45 -3305
rect -75 -3400 -45 -3370
rect -75 -3470 -45 -3440
rect -75 -3540 -45 -3510
rect -75 -3610 -45 -3580
rect -75 -3675 -45 -3645
rect -75 -3735 -45 -3705
rect -75 -3800 -45 -3770
rect -75 -3870 -45 -3840
rect -75 -3940 -45 -3910
rect -75 -4010 -45 -3980
rect -75 -4075 -45 -4045
rect -75 -4135 -45 -4105
rect -75 -4200 -45 -4170
rect -75 -4270 -45 -4240
rect -75 -4340 -45 -4310
rect -75 -4410 -45 -4380
rect -75 -4475 -45 -4445
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 275 -2935 305 -2905
rect 275 -3000 305 -2970
rect 275 -3070 305 -3040
rect 275 -3140 305 -3110
rect 275 -3210 305 -3180
rect 275 -3275 305 -3245
rect 275 -3335 305 -3305
rect 275 -3400 305 -3370
rect 275 -3470 305 -3440
rect 275 -3540 305 -3510
rect 275 -3610 305 -3580
rect 275 -3675 305 -3645
rect 275 -3735 305 -3705
rect 275 -3800 305 -3770
rect 275 -3870 305 -3840
rect 275 -3940 305 -3910
rect 275 -4010 305 -3980
rect 275 -4075 305 -4045
rect 275 -4135 305 -4105
rect 275 -4200 305 -4170
rect 275 -4270 305 -4240
rect 275 -4340 305 -4310
rect 275 -4410 305 -4380
rect 275 -4475 305 -4445
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 625 -2935 655 -2905
rect 625 -3000 655 -2970
rect 625 -3070 655 -3040
rect 625 -3140 655 -3110
rect 625 -3210 655 -3180
rect 625 -3275 655 -3245
rect 625 -3335 655 -3305
rect 625 -3400 655 -3370
rect 625 -3470 655 -3440
rect 625 -3540 655 -3510
rect 625 -3610 655 -3580
rect 625 -3675 655 -3645
rect 625 -3735 655 -3705
rect 625 -3800 655 -3770
rect 625 -3870 655 -3840
rect 625 -3940 655 -3910
rect 625 -4010 655 -3980
rect 625 -4075 655 -4045
rect 625 -4135 655 -4105
rect 625 -4200 655 -4170
rect 625 -4270 655 -4240
rect 625 -4340 655 -4310
rect 625 -4410 655 -4380
rect 625 -4475 655 -4445
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 975 -2935 1005 -2905
rect 975 -3000 1005 -2970
rect 975 -3070 1005 -3040
rect 975 -3140 1005 -3110
rect 975 -3210 1005 -3180
rect 975 -3275 1005 -3245
rect 975 -3335 1005 -3305
rect 975 -3400 1005 -3370
rect 975 -3470 1005 -3440
rect 975 -3540 1005 -3510
rect 975 -3610 1005 -3580
rect 975 -3675 1005 -3645
rect 975 -3735 1005 -3705
rect 975 -3800 1005 -3770
rect 975 -3870 1005 -3840
rect 975 -3940 1005 -3910
rect 975 -4010 1005 -3980
rect 975 -4075 1005 -4045
rect 975 -4135 1005 -4105
rect 975 -4200 1005 -4170
rect 975 -4270 1005 -4240
rect 975 -4340 1005 -4310
rect 975 -4410 1005 -4380
rect 975 -4475 1005 -4445
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1325 -2935 1355 -2905
rect 1325 -3000 1355 -2970
rect 1325 -3070 1355 -3040
rect 1325 -3140 1355 -3110
rect 1325 -3210 1355 -3180
rect 1325 -3275 1355 -3245
rect 1325 -3335 1355 -3305
rect 1325 -3400 1355 -3370
rect 1325 -3470 1355 -3440
rect 1325 -3540 1355 -3510
rect 1325 -3610 1355 -3580
rect 1325 -3675 1355 -3645
rect 1325 -3735 1355 -3705
rect 1325 -3800 1355 -3770
rect 1325 -3870 1355 -3840
rect 1325 -3940 1355 -3910
rect 1325 -4010 1355 -3980
rect 1325 -4075 1355 -4045
rect 1325 -4135 1355 -4105
rect 1325 -4200 1355 -4170
rect 1325 -4270 1355 -4240
rect 1325 -4340 1355 -4310
rect 1325 -4410 1355 -4380
rect 1325 -4475 1355 -4445
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 1675 -2935 1705 -2905
rect 1675 -3000 1705 -2970
rect 1675 -3070 1705 -3040
rect 1675 -3140 1705 -3110
rect 1675 -3210 1705 -3180
rect 1675 -3275 1705 -3245
rect 1675 -3335 1705 -3305
rect 1675 -3400 1705 -3370
rect 1675 -3470 1705 -3440
rect 1675 -3540 1705 -3510
rect 1675 -3610 1705 -3580
rect 1675 -3675 1705 -3645
rect 1675 -3735 1705 -3705
rect 1675 -3800 1705 -3770
rect 1675 -3870 1705 -3840
rect 1675 -3940 1705 -3910
rect 1675 -4010 1705 -3980
rect 1675 -4075 1705 -4045
rect 1675 -4135 1705 -4105
rect 1675 -4200 1705 -4170
rect 1675 -4270 1705 -4240
rect 1675 -4340 1705 -4310
rect 1675 -4410 1705 -4380
rect 1675 -4475 1705 -4445
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2025 -2935 2055 -2905
rect 2025 -3000 2055 -2970
rect 2025 -3070 2055 -3040
rect 2025 -3140 2055 -3110
rect 2025 -3210 2055 -3180
rect 2025 -3275 2055 -3245
rect 2025 -3335 2055 -3305
rect 2025 -3400 2055 -3370
rect 2025 -3470 2055 -3440
rect 2025 -3540 2055 -3510
rect 2025 -3610 2055 -3580
rect 2025 -3675 2055 -3645
rect 2025 -3735 2055 -3705
rect 2025 -3800 2055 -3770
rect 2025 -3870 2055 -3840
rect 2025 -3940 2055 -3910
rect 2025 -4010 2055 -3980
rect 2025 -4075 2055 -4045
rect 2025 -4135 2055 -4105
rect 2025 -4200 2055 -4170
rect 2025 -4270 2055 -4240
rect 2025 -4340 2055 -4310
rect 2025 -4410 2055 -4380
rect 2025 -4475 2055 -4445
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2375 -2935 2405 -2905
rect 2375 -3000 2405 -2970
rect 2375 -3070 2405 -3040
rect 2375 -3140 2405 -3110
rect 2375 -3210 2405 -3180
rect 2375 -3275 2405 -3245
rect 2375 -3335 2405 -3305
rect 2375 -3400 2405 -3370
rect 2375 -3470 2405 -3440
rect 2375 -3540 2405 -3510
rect 2375 -3610 2405 -3580
rect 2375 -3675 2405 -3645
rect 2375 -3735 2405 -3705
rect 2375 -3800 2405 -3770
rect 2375 -3870 2405 -3840
rect 2375 -3940 2405 -3910
rect 2375 -4010 2405 -3980
rect 2375 -4075 2405 -4045
rect 2375 -4135 2405 -4105
rect 2375 -4200 2405 -4170
rect 2375 -4270 2405 -4240
rect 2375 -4340 2405 -4310
rect 2375 -4410 2405 -4380
rect 2375 -4475 2405 -4445
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 2725 -2935 2755 -2905
rect 2725 -3000 2755 -2970
rect 2725 -3070 2755 -3040
rect 2725 -3140 2755 -3110
rect 2725 -3210 2755 -3180
rect 2725 -3275 2755 -3245
rect 2725 -3335 2755 -3305
rect 2725 -3400 2755 -3370
rect 2725 -3470 2755 -3440
rect 2725 -3540 2755 -3510
rect 2725 -3610 2755 -3580
rect 2725 -3675 2755 -3645
rect 2725 -3735 2755 -3705
rect 2725 -3800 2755 -3770
rect 2725 -3870 2755 -3840
rect 2725 -3940 2755 -3910
rect 2725 -4010 2755 -3980
rect 2725 -4075 2755 -4045
rect 2725 -4135 2755 -4105
rect 2725 -4200 2755 -4170
rect 2725 -4270 2755 -4240
rect 2725 -4340 2755 -4310
rect 2725 -4410 2755 -4380
rect 2725 -4475 2755 -4445
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3075 -2935 3105 -2905
rect 3075 -3000 3105 -2970
rect 3075 -3070 3105 -3040
rect 3075 -3140 3105 -3110
rect 3075 -3210 3105 -3180
rect 3075 -3275 3105 -3245
rect 3075 -3335 3105 -3305
rect 3075 -3400 3105 -3370
rect 3075 -3470 3105 -3440
rect 3075 -3540 3105 -3510
rect 3075 -3610 3105 -3580
rect 3075 -3675 3105 -3645
rect 3075 -3735 3105 -3705
rect 3075 -3800 3105 -3770
rect 3075 -3870 3105 -3840
rect 3075 -3940 3105 -3910
rect 3075 -4010 3105 -3980
rect 3075 -4075 3105 -4045
rect 3075 -4135 3105 -4105
rect 3075 -4200 3105 -4170
rect 3075 -4270 3105 -4240
rect 3075 -4340 3105 -4310
rect 3075 -4410 3105 -4380
rect 3075 -4475 3105 -4445
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3425 -2935 3455 -2905
rect 3425 -3000 3455 -2970
rect 3425 -3070 3455 -3040
rect 3425 -3140 3455 -3110
rect 3425 -3210 3455 -3180
rect 3425 -3275 3455 -3245
rect 3425 -3335 3455 -3305
rect 3425 -3400 3455 -3370
rect 3425 -3470 3455 -3440
rect 3425 -3540 3455 -3510
rect 3425 -3610 3455 -3580
rect 3425 -3675 3455 -3645
rect 3425 -3735 3455 -3705
rect 3425 -3800 3455 -3770
rect 3425 -3870 3455 -3840
rect 3425 -3940 3455 -3910
rect 3425 -4010 3455 -3980
rect 3425 -4075 3455 -4045
rect 3425 -4135 3455 -4105
rect 3425 -4200 3455 -4170
rect 3425 -4270 3455 -4240
rect 3425 -4340 3455 -4310
rect 3425 -4410 3455 -4380
rect 3425 -4475 3455 -4445
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 3775 -2935 3805 -2905
rect 3775 -3000 3805 -2970
rect 3775 -3070 3805 -3040
rect 3775 -3140 3805 -3110
rect 3775 -3210 3805 -3180
rect 3775 -3275 3805 -3245
rect 3775 -3335 3805 -3305
rect 3775 -3400 3805 -3370
rect 3775 -3470 3805 -3440
rect 3775 -3540 3805 -3510
rect 3775 -3610 3805 -3580
rect 3775 -3675 3805 -3645
rect 3775 -3735 3805 -3705
rect 3775 -3800 3805 -3770
rect 3775 -3870 3805 -3840
rect 3775 -3940 3805 -3910
rect 3775 -4010 3805 -3980
rect 3775 -4075 3805 -4045
rect 3775 -4135 3805 -4105
rect 3775 -4200 3805 -4170
rect 3775 -4270 3805 -4240
rect 3775 -4340 3805 -4310
rect 3775 -4410 3805 -4380
rect 3775 -4475 3805 -4445
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4125 -2935 4155 -2905
rect 4125 -3000 4155 -2970
rect 4125 -3070 4155 -3040
rect 4125 -3140 4155 -3110
rect 4125 -3210 4155 -3180
rect 4125 -3275 4155 -3245
rect 4125 -3335 4155 -3305
rect 4125 -3400 4155 -3370
rect 4125 -3470 4155 -3440
rect 4125 -3540 4155 -3510
rect 4125 -3610 4155 -3580
rect 4125 -3675 4155 -3645
rect 4125 -3735 4155 -3705
rect 4125 -3800 4155 -3770
rect 4125 -3870 4155 -3840
rect 4125 -3940 4155 -3910
rect 4125 -4010 4155 -3980
rect 4125 -4075 4155 -4045
rect 4125 -4135 4155 -4105
rect 4125 -4200 4155 -4170
rect 4125 -4270 4155 -4240
rect 4125 -4340 4155 -4310
rect 4125 -4410 4155 -4380
rect 4125 -4475 4155 -4445
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4475 -2935 4505 -2905
rect 4475 -3000 4505 -2970
rect 4475 -3070 4505 -3040
rect 4475 -3140 4505 -3110
rect 4475 -3210 4505 -3180
rect 4475 -3275 4505 -3245
rect 4475 -3335 4505 -3305
rect 4475 -3400 4505 -3370
rect 4475 -3470 4505 -3440
rect 4475 -3540 4505 -3510
rect 4475 -3610 4505 -3580
rect 4475 -3675 4505 -3645
rect 4475 -3735 4505 -3705
rect 4475 -3800 4505 -3770
rect 4475 -3870 4505 -3840
rect 4475 -3940 4505 -3910
rect 4475 -4010 4505 -3980
rect 4475 -4075 4505 -4045
rect 4475 -4135 4505 -4105
rect 4475 -4200 4505 -4170
rect 4475 -4270 4505 -4240
rect 4475 -4340 4505 -4310
rect 4475 -4410 4505 -4380
rect 4475 -4475 4505 -4445
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 4825 -2935 4855 -2905
rect 4825 -3000 4855 -2970
rect 4825 -3070 4855 -3040
rect 4825 -3140 4855 -3110
rect 4825 -3210 4855 -3180
rect 4825 -3275 4855 -3245
rect 4825 -3335 4855 -3305
rect 4825 -3400 4855 -3370
rect 4825 -3470 4855 -3440
rect 4825 -3540 4855 -3510
rect 4825 -3610 4855 -3580
rect 4825 -3675 4855 -3645
rect 4825 -3735 4855 -3705
rect 4825 -3800 4855 -3770
rect 4825 -3870 4855 -3840
rect 4825 -3940 4855 -3910
rect 4825 -4010 4855 -3980
rect 4825 -4075 4855 -4045
rect 4825 -4135 4855 -4105
rect 4825 -4200 4855 -4170
rect 4825 -4270 4855 -4240
rect 4825 -4340 4855 -4310
rect 4825 -4410 4855 -4380
rect 4825 -4475 4855 -4445
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5175 -2935 5205 -2905
rect 5175 -3000 5205 -2970
rect 5175 -3070 5205 -3040
rect 5175 -3140 5205 -3110
rect 5175 -3210 5205 -3180
rect 5175 -3275 5205 -3245
rect 5175 -3335 5205 -3305
rect 5175 -3400 5205 -3370
rect 5175 -3470 5205 -3440
rect 5175 -3540 5205 -3510
rect 5175 -3610 5205 -3580
rect 5175 -3675 5205 -3645
rect 5175 -3735 5205 -3705
rect 5175 -3800 5205 -3770
rect 5175 -3870 5205 -3840
rect 5175 -3940 5205 -3910
rect 5175 -4010 5205 -3980
rect 5175 -4075 5205 -4045
rect 5175 -4135 5205 -4105
rect 5175 -4200 5205 -4170
rect 5175 -4270 5205 -4240
rect 5175 -4340 5205 -4310
rect 5175 -4410 5205 -4380
rect 5175 -4475 5205 -4445
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5525 -2935 5555 -2905
rect 5525 -3000 5555 -2970
rect 5525 -3070 5555 -3040
rect 5525 -3140 5555 -3110
rect 5525 -3210 5555 -3180
rect 5525 -3275 5555 -3245
rect 5525 -3335 5555 -3305
rect 5525 -3400 5555 -3370
rect 5525 -3470 5555 -3440
rect 5525 -3540 5555 -3510
rect 5525 -3610 5555 -3580
rect 5525 -3675 5555 -3645
rect 5525 -3735 5555 -3705
rect 5525 -3800 5555 -3770
rect 5525 -3870 5555 -3840
rect 5525 -3940 5555 -3910
rect 5525 -4010 5555 -3980
rect 5525 -4075 5555 -4045
rect 5525 -4135 5555 -4105
rect 5525 -4200 5555 -4170
rect 5525 -4270 5555 -4240
rect 5525 -4340 5555 -4310
rect 5525 -4410 5555 -4380
rect 5525 -4475 5555 -4445
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 5875 -2935 5905 -2905
rect 5875 -3000 5905 -2970
rect 5875 -3070 5905 -3040
rect 5875 -3140 5905 -3110
rect 5875 -3210 5905 -3180
rect 5875 -3275 5905 -3245
rect 5875 -3335 5905 -3305
rect 5875 -3400 5905 -3370
rect 5875 -3470 5905 -3440
rect 5875 -3540 5905 -3510
rect 5875 -3610 5905 -3580
rect 5875 -3675 5905 -3645
rect 5875 -3735 5905 -3705
rect 5875 -3800 5905 -3770
rect 5875 -3870 5905 -3840
rect 5875 -3940 5905 -3910
rect 5875 -4010 5905 -3980
rect 5875 -4075 5905 -4045
rect 5875 -4135 5905 -4105
rect 5875 -4200 5905 -4170
rect 5875 -4270 5905 -4240
rect 5875 -4340 5905 -4310
rect 5875 -4410 5905 -4380
rect 5875 -4475 5905 -4445
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6225 -2935 6255 -2905
rect 6225 -3000 6255 -2970
rect 6225 -3070 6255 -3040
rect 6225 -3140 6255 -3110
rect 6225 -3210 6255 -3180
rect 6225 -3275 6255 -3245
rect 6225 -3335 6255 -3305
rect 6225 -3400 6255 -3370
rect 6225 -3470 6255 -3440
rect 6225 -3540 6255 -3510
rect 6225 -3610 6255 -3580
rect 6225 -3675 6255 -3645
rect 6225 -3735 6255 -3705
rect 6225 -3800 6255 -3770
rect 6225 -3870 6255 -3840
rect 6225 -3940 6255 -3910
rect 6225 -4010 6255 -3980
rect 6225 -4075 6255 -4045
rect 6225 -4135 6255 -4105
rect 6225 -4200 6255 -4170
rect 6225 -4270 6255 -4240
rect 6225 -4340 6255 -4310
rect 6225 -4410 6255 -4380
rect 6225 -4475 6255 -4445
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6575 -2935 6605 -2905
rect 6575 -3000 6605 -2970
rect 6575 -3070 6605 -3040
rect 6575 -3140 6605 -3110
rect 6575 -3210 6605 -3180
rect 6575 -3275 6605 -3245
rect 6575 -3335 6605 -3305
rect 6575 -3400 6605 -3370
rect 6575 -3470 6605 -3440
rect 6575 -3540 6605 -3510
rect 6575 -3610 6605 -3580
rect 6575 -3675 6605 -3645
rect 6575 -3735 6605 -3705
rect 6575 -3800 6605 -3770
rect 6575 -3870 6605 -3840
rect 6575 -3940 6605 -3910
rect 6575 -4010 6605 -3980
rect 6575 -4075 6605 -4045
rect 6575 -4135 6605 -4105
rect 6575 -4200 6605 -4170
rect 6575 -4270 6605 -4240
rect 6575 -4340 6605 -4310
rect 6575 -4410 6605 -4380
rect 6575 -4475 6605 -4445
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 6925 -2935 6955 -2905
rect 6925 -3000 6955 -2970
rect 6925 -3070 6955 -3040
rect 6925 -3140 6955 -3110
rect 6925 -3210 6955 -3180
rect 6925 -3275 6955 -3245
rect 6925 -3335 6955 -3305
rect 6925 -3400 6955 -3370
rect 6925 -3470 6955 -3440
rect 6925 -3540 6955 -3510
rect 6925 -3610 6955 -3580
rect 6925 -3675 6955 -3645
rect 6925 -3735 6955 -3705
rect 6925 -3800 6955 -3770
rect 6925 -3870 6955 -3840
rect 6925 -3940 6955 -3910
rect 6925 -4010 6955 -3980
rect 6925 -4075 6955 -4045
rect 6925 -4135 6955 -4105
rect 6925 -4200 6955 -4170
rect 6925 -4270 6955 -4240
rect 6925 -4340 6955 -4310
rect 6925 -4410 6955 -4380
rect 6925 -4475 6955 -4445
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7275 -2935 7305 -2905
rect 7275 -3000 7305 -2970
rect 7275 -3070 7305 -3040
rect 7275 -3140 7305 -3110
rect 7275 -3210 7305 -3180
rect 7275 -3275 7305 -3245
rect 7275 -3335 7305 -3305
rect 7275 -3400 7305 -3370
rect 7275 -3470 7305 -3440
rect 7275 -3540 7305 -3510
rect 7275 -3610 7305 -3580
rect 7275 -3675 7305 -3645
rect 7275 -3735 7305 -3705
rect 7275 -3800 7305 -3770
rect 7275 -3870 7305 -3840
rect 7275 -3940 7305 -3910
rect 7275 -4010 7305 -3980
rect 7275 -4075 7305 -4045
rect 7275 -4135 7305 -4105
rect 7275 -4200 7305 -4170
rect 7275 -4270 7305 -4240
rect 7275 -4340 7305 -4310
rect 7275 -4410 7305 -4380
rect 7275 -4475 7305 -4445
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7625 -2935 7655 -2905
rect 7625 -3000 7655 -2970
rect 7625 -3070 7655 -3040
rect 7625 -3140 7655 -3110
rect 7625 -3210 7655 -3180
rect 7625 -3275 7655 -3245
rect 7625 -3335 7655 -3305
rect 7625 -3400 7655 -3370
rect 7625 -3470 7655 -3440
rect 7625 -3540 7655 -3510
rect 7625 -3610 7655 -3580
rect 7625 -3675 7655 -3645
rect 7625 -3735 7655 -3705
rect 7625 -3800 7655 -3770
rect 7625 -3870 7655 -3840
rect 7625 -3940 7655 -3910
rect 7625 -4010 7655 -3980
rect 7625 -4075 7655 -4045
rect 7625 -4135 7655 -4105
rect 7625 -4200 7655 -4170
rect 7625 -4270 7655 -4240
rect 7625 -4340 7655 -4310
rect 7625 -4410 7655 -4380
rect 7625 -4475 7655 -4445
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 7975 -2935 8005 -2905
rect 7975 -3000 8005 -2970
rect 7975 -3070 8005 -3040
rect 7975 -3140 8005 -3110
rect 7975 -3210 8005 -3180
rect 7975 -3275 8005 -3245
rect 7975 -3335 8005 -3305
rect 7975 -3400 8005 -3370
rect 7975 -3470 8005 -3440
rect 7975 -3540 8005 -3510
rect 7975 -3610 8005 -3580
rect 7975 -3675 8005 -3645
rect 7975 -3735 8005 -3705
rect 7975 -3800 8005 -3770
rect 7975 -3870 8005 -3840
rect 7975 -3940 8005 -3910
rect 7975 -4010 8005 -3980
rect 7975 -4075 8005 -4045
rect 7975 -4135 8005 -4105
rect 7975 -4200 8005 -4170
rect 7975 -4270 8005 -4240
rect 7975 -4340 8005 -4310
rect 7975 -4410 8005 -4380
rect 7975 -4475 8005 -4445
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8325 -2935 8355 -2905
rect 8325 -3000 8355 -2970
rect 8325 -3070 8355 -3040
rect 8325 -3140 8355 -3110
rect 8325 -3210 8355 -3180
rect 8325 -3275 8355 -3245
rect 8325 -3335 8355 -3305
rect 8325 -3400 8355 -3370
rect 8325 -3470 8355 -3440
rect 8325 -3540 8355 -3510
rect 8325 -3610 8355 -3580
rect 8325 -3675 8355 -3645
rect 8325 -3735 8355 -3705
rect 8325 -3800 8355 -3770
rect 8325 -3870 8355 -3840
rect 8325 -3940 8355 -3910
rect 8325 -4010 8355 -3980
rect 8325 -4075 8355 -4045
rect 8325 -4135 8355 -4105
rect 8325 -4200 8355 -4170
rect 8325 -4270 8355 -4240
rect 8325 -4340 8355 -4310
rect 8325 -4410 8355 -4380
rect 8325 -4475 8355 -4445
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 8675 -2935 8705 -2905
rect 8675 -3000 8705 -2970
rect 8675 -3070 8705 -3040
rect 8675 -3140 8705 -3110
rect 8675 -3210 8705 -3180
rect 8675 -3275 8705 -3245
rect 8675 -3335 8705 -3305
rect 8675 -3400 8705 -3370
rect 8675 -3470 8705 -3440
rect 8675 -3540 8705 -3510
rect 8675 -3610 8705 -3580
rect 8675 -3675 8705 -3645
rect 8675 -3735 8705 -3705
rect 8675 -3800 8705 -3770
rect 8675 -3870 8705 -3840
rect 8675 -3940 8705 -3910
rect 8675 -4010 8705 -3980
rect 8675 -4075 8705 -4045
rect 8675 -4135 8705 -4105
rect 8675 -4200 8705 -4170
rect 8675 -4270 8705 -4240
rect 8675 -4340 8705 -4310
rect 8675 -4410 8705 -4380
rect 8675 -4475 8705 -4445
<< metal3 >>
rect 2320 20915 2380 20925
rect 2320 20875 2330 20915
rect 2370 20875 2380 20915
rect 2320 20850 2380 20875
rect 2320 20810 2330 20850
rect 2370 20810 2380 20850
rect 2320 20780 2380 20810
rect 2320 20740 2330 20780
rect 2370 20740 2380 20780
rect 2320 20710 2380 20740
rect 2320 20670 2330 20710
rect 2370 20670 2380 20710
rect 2320 20640 2380 20670
rect 2320 20600 2330 20640
rect 2370 20600 2380 20640
rect 2320 20575 2380 20600
rect 2320 20535 2330 20575
rect 2370 20535 2380 20575
rect 2320 20515 2380 20535
rect 2320 20475 2330 20515
rect 2370 20475 2380 20515
rect 2320 20450 2380 20475
rect 2320 20410 2330 20450
rect 2370 20410 2380 20450
rect 2320 20380 2380 20410
rect 2320 20340 2330 20380
rect 2370 20340 2380 20380
rect 2320 20310 2380 20340
rect 2320 20270 2330 20310
rect 2370 20270 2380 20310
rect 2320 20240 2380 20270
rect 2320 20200 2330 20240
rect 2370 20200 2380 20240
rect 2320 20175 2380 20200
rect 2320 20135 2330 20175
rect 2370 20135 2380 20175
rect 2320 20115 2380 20135
rect 2320 20075 2330 20115
rect 2370 20075 2380 20115
rect 2320 20050 2380 20075
rect 2320 20010 2330 20050
rect 2370 20010 2380 20050
rect 2320 19980 2380 20010
rect 2320 19940 2330 19980
rect 2370 19940 2380 19980
rect 2320 19910 2380 19940
rect 2320 19870 2330 19910
rect 2370 19870 2380 19910
rect 2320 19840 2380 19870
rect 2320 19800 2330 19840
rect 2370 19800 2380 19840
rect 2320 19775 2380 19800
rect 2320 19735 2330 19775
rect 2370 19735 2380 19775
rect 2320 19715 2380 19735
rect 2320 19675 2330 19715
rect 2370 19675 2380 19715
rect 2320 19650 2380 19675
rect 2320 19610 2330 19650
rect 2370 19610 2380 19650
rect 2320 19580 2380 19610
rect 2320 19540 2330 19580
rect 2370 19540 2380 19580
rect 2320 19510 2380 19540
rect 2320 19470 2330 19510
rect 2370 19470 2380 19510
rect 2320 19440 2380 19470
rect 2320 19400 2330 19440
rect 2370 19400 2380 19440
rect 2320 19375 2380 19400
rect 2320 19335 2330 19375
rect 2370 19335 2380 19375
rect 2320 19315 2380 19335
rect 2320 19275 2330 19315
rect 2370 19275 2380 19315
rect 2320 19250 2380 19275
rect 2320 19210 2330 19250
rect 2370 19210 2380 19250
rect 2320 19180 2380 19210
rect 2320 19140 2330 19180
rect 2370 19140 2380 19180
rect 2320 19110 2380 19140
rect 2320 19070 2330 19110
rect 2370 19070 2380 19110
rect 2320 19040 2380 19070
rect 2320 19000 2330 19040
rect 2370 19000 2380 19040
rect 2320 18975 2380 19000
rect 2320 18935 2330 18975
rect 2370 18935 2380 18975
rect 2320 18915 2380 18935
rect 2320 18875 2330 18915
rect 2370 18875 2380 18915
rect 2320 18850 2380 18875
rect 2320 18810 2330 18850
rect 2370 18810 2380 18850
rect 2320 18780 2380 18810
rect 2320 18740 2330 18780
rect 2370 18740 2380 18780
rect 2320 18710 2380 18740
rect 2320 18670 2330 18710
rect 2370 18670 2380 18710
rect 2320 18640 2380 18670
rect 2320 18600 2330 18640
rect 2370 18600 2380 18640
rect 2320 18575 2380 18600
rect 2320 18535 2330 18575
rect 2370 18535 2380 18575
rect 2320 18515 2380 18535
rect 2320 18475 2330 18515
rect 2370 18475 2380 18515
rect 2320 18450 2380 18475
rect 2320 18410 2330 18450
rect 2370 18410 2380 18450
rect 2320 18380 2380 18410
rect 2320 18340 2330 18380
rect 2370 18340 2380 18380
rect 2320 18310 2380 18340
rect 2320 18270 2330 18310
rect 2370 18270 2380 18310
rect 2320 18240 2380 18270
rect -1260 18145 -1030 18230
rect -910 18145 -680 18230
rect -560 18145 -330 18230
rect -210 18145 20 18230
rect 140 18145 370 18230
rect 490 18145 720 18230
rect 840 18145 1070 18230
rect 1190 18145 1420 18230
rect 1540 18145 1770 18230
rect -1260 18095 1770 18145
rect -1260 18000 -1030 18095
rect -910 18000 -680 18095
rect -560 18000 -330 18095
rect -210 18000 20 18095
rect 140 18000 370 18095
rect 490 18000 720 18095
rect 840 18000 1070 18095
rect 1190 18000 1420 18095
rect 1540 18000 1770 18095
rect 2320 18200 2330 18240
rect 2370 18200 2380 18240
rect 2320 18175 2380 18200
rect 2320 18135 2330 18175
rect 2370 18135 2380 18175
rect 2320 18115 2380 18135
rect 2320 18075 2330 18115
rect 2370 18075 2380 18115
rect 2320 18050 2380 18075
rect 2320 18010 2330 18050
rect 2370 18010 2380 18050
rect 230 17880 280 18000
rect 2320 17980 2380 18010
rect 2320 17940 2330 17980
rect 2370 17940 2380 17980
rect 2320 17910 2380 17940
rect -1260 17795 -1030 17880
rect -910 17795 -680 17880
rect -560 17795 -330 17880
rect -210 17795 20 17880
rect 140 17795 370 17880
rect 490 17795 720 17880
rect 840 17795 1070 17880
rect 1190 17795 1420 17880
rect 1540 17795 1770 17880
rect -1260 17745 1770 17795
rect -1260 17650 -1030 17745
rect -910 17650 -680 17745
rect -560 17650 -330 17745
rect -210 17650 20 17745
rect 140 17650 370 17745
rect 490 17650 720 17745
rect 840 17650 1070 17745
rect 1190 17650 1420 17745
rect 1540 17650 1770 17745
rect 2320 17870 2330 17910
rect 2370 17870 2380 17910
rect 2320 17840 2380 17870
rect 2320 17800 2330 17840
rect 2370 17800 2380 17840
rect 2320 17775 2380 17800
rect 2320 17735 2330 17775
rect 2370 17735 2380 17775
rect 2320 17725 2380 17735
rect 6690 20915 6750 20925
rect 6690 20875 6700 20915
rect 6740 20875 6750 20915
rect 6690 20850 6750 20875
rect 6690 20810 6700 20850
rect 6740 20810 6750 20850
rect 6690 20780 6750 20810
rect 6690 20740 6700 20780
rect 6740 20740 6750 20780
rect 6690 20710 6750 20740
rect 6690 20670 6700 20710
rect 6740 20670 6750 20710
rect 6690 20640 6750 20670
rect 6690 20600 6700 20640
rect 6740 20600 6750 20640
rect 6690 20575 6750 20600
rect 6690 20535 6700 20575
rect 6740 20535 6750 20575
rect 6690 20515 6750 20535
rect 6690 20475 6700 20515
rect 6740 20475 6750 20515
rect 6690 20450 6750 20475
rect 6690 20410 6700 20450
rect 6740 20410 6750 20450
rect 6690 20380 6750 20410
rect 6690 20340 6700 20380
rect 6740 20340 6750 20380
rect 6690 20310 6750 20340
rect 6690 20270 6700 20310
rect 6740 20270 6750 20310
rect 6690 20240 6750 20270
rect 6690 20200 6700 20240
rect 6740 20200 6750 20240
rect 6690 20175 6750 20200
rect 6690 20135 6700 20175
rect 6740 20135 6750 20175
rect 6690 20115 6750 20135
rect 6690 20075 6700 20115
rect 6740 20075 6750 20115
rect 6690 20050 6750 20075
rect 6690 20010 6700 20050
rect 6740 20010 6750 20050
rect 6690 19980 6750 20010
rect 6690 19940 6700 19980
rect 6740 19940 6750 19980
rect 6690 19910 6750 19940
rect 6690 19870 6700 19910
rect 6740 19870 6750 19910
rect 6690 19840 6750 19870
rect 6690 19800 6700 19840
rect 6740 19800 6750 19840
rect 6690 19775 6750 19800
rect 6690 19735 6700 19775
rect 6740 19735 6750 19775
rect 6690 19715 6750 19735
rect 6690 19675 6700 19715
rect 6740 19675 6750 19715
rect 6690 19650 6750 19675
rect 6690 19610 6700 19650
rect 6740 19610 6750 19650
rect 6690 19580 6750 19610
rect 6690 19540 6700 19580
rect 6740 19540 6750 19580
rect 6690 19510 6750 19540
rect 6690 19470 6700 19510
rect 6740 19470 6750 19510
rect 6690 19440 6750 19470
rect 6690 19400 6700 19440
rect 6740 19400 6750 19440
rect 6690 19375 6750 19400
rect 6690 19335 6700 19375
rect 6740 19335 6750 19375
rect 6690 19315 6750 19335
rect 6690 19275 6700 19315
rect 6740 19275 6750 19315
rect 6690 19250 6750 19275
rect 6690 19210 6700 19250
rect 6740 19210 6750 19250
rect 6690 19180 6750 19210
rect 6690 19140 6700 19180
rect 6740 19140 6750 19180
rect 6690 19110 6750 19140
rect 6690 19070 6700 19110
rect 6740 19070 6750 19110
rect 6690 19040 6750 19070
rect 6690 19000 6700 19040
rect 6740 19000 6750 19040
rect 6690 18975 6750 19000
rect 6690 18935 6700 18975
rect 6740 18935 6750 18975
rect 6690 18915 6750 18935
rect 6690 18875 6700 18915
rect 6740 18875 6750 18915
rect 6690 18850 6750 18875
rect 6690 18810 6700 18850
rect 6740 18810 6750 18850
rect 6690 18780 6750 18810
rect 6690 18740 6700 18780
rect 6740 18740 6750 18780
rect 6690 18710 6750 18740
rect 6690 18670 6700 18710
rect 6740 18670 6750 18710
rect 6690 18640 6750 18670
rect 6690 18600 6700 18640
rect 6740 18600 6750 18640
rect 6690 18575 6750 18600
rect 6690 18535 6700 18575
rect 6740 18535 6750 18575
rect 6690 18515 6750 18535
rect 6690 18475 6700 18515
rect 6740 18475 6750 18515
rect 6690 18450 6750 18475
rect 6690 18410 6700 18450
rect 6740 18410 6750 18450
rect 6690 18380 6750 18410
rect 6690 18340 6700 18380
rect 6740 18340 6750 18380
rect 6690 18310 6750 18340
rect 6690 18270 6700 18310
rect 6740 18270 6750 18310
rect 6690 18240 6750 18270
rect 6690 18200 6700 18240
rect 6740 18200 6750 18240
rect 6690 18175 6750 18200
rect 6690 18135 6700 18175
rect 6740 18135 6750 18175
rect 6690 18115 6750 18135
rect 6690 18075 6700 18115
rect 6740 18075 6750 18115
rect 6690 18050 6750 18075
rect 6690 18010 6700 18050
rect 6740 18010 6750 18050
rect 6690 17980 6750 18010
rect 6690 17940 6700 17980
rect 6740 17940 6750 17980
rect 6690 17910 6750 17940
rect 6690 17870 6700 17910
rect 6740 17870 6750 17910
rect 6690 17840 6750 17870
rect 6690 17800 6700 17840
rect 6740 17800 6750 17840
rect 6690 17775 6750 17800
rect 6690 17735 6700 17775
rect 6740 17735 6750 17775
rect 6690 17725 6750 17735
rect 14790 20890 17990 20925
rect 14790 20840 14825 20890
rect 14875 20840 14920 20890
rect 14970 20840 15015 20890
rect 15065 20840 15115 20890
rect 15165 20840 15215 20890
rect 15265 20840 15315 20890
rect 15365 20840 15410 20890
rect 15460 20840 15505 20890
rect 15555 20840 15625 20890
rect 15675 20840 15720 20890
rect 15770 20840 15815 20890
rect 15865 20840 15915 20890
rect 15965 20840 16015 20890
rect 16065 20840 16115 20890
rect 16165 20840 16210 20890
rect 16260 20840 16305 20890
rect 16355 20840 16425 20890
rect 16475 20840 16520 20890
rect 16570 20840 16615 20890
rect 16665 20840 16715 20890
rect 16765 20840 16815 20890
rect 16865 20840 16915 20890
rect 16965 20840 17010 20890
rect 17060 20840 17105 20890
rect 17155 20840 17225 20890
rect 17275 20840 17320 20890
rect 17370 20840 17415 20890
rect 17465 20840 17515 20890
rect 17565 20840 17615 20890
rect 17665 20840 17715 20890
rect 17765 20840 17810 20890
rect 17860 20840 17905 20890
rect 17955 20840 17990 20890
rect 14790 20800 17990 20840
rect 14790 20750 14825 20800
rect 14875 20750 14920 20800
rect 14970 20750 15015 20800
rect 15065 20750 15115 20800
rect 15165 20750 15215 20800
rect 15265 20750 15315 20800
rect 15365 20750 15410 20800
rect 15460 20750 15505 20800
rect 15555 20750 15625 20800
rect 15675 20750 15720 20800
rect 15770 20750 15815 20800
rect 15865 20750 15915 20800
rect 15965 20750 16015 20800
rect 16065 20750 16115 20800
rect 16165 20750 16210 20800
rect 16260 20750 16305 20800
rect 16355 20750 16425 20800
rect 16475 20750 16520 20800
rect 16570 20750 16615 20800
rect 16665 20750 16715 20800
rect 16765 20750 16815 20800
rect 16865 20750 16915 20800
rect 16965 20750 17010 20800
rect 17060 20750 17105 20800
rect 17155 20750 17225 20800
rect 17275 20750 17320 20800
rect 17370 20750 17415 20800
rect 17465 20750 17515 20800
rect 17565 20750 17615 20800
rect 17665 20750 17715 20800
rect 17765 20750 17810 20800
rect 17860 20750 17905 20800
rect 17955 20750 17990 20800
rect 14790 20700 17990 20750
rect 14790 20650 14825 20700
rect 14875 20650 14920 20700
rect 14970 20650 15015 20700
rect 15065 20650 15115 20700
rect 15165 20650 15215 20700
rect 15265 20650 15315 20700
rect 15365 20650 15410 20700
rect 15460 20650 15505 20700
rect 15555 20650 15625 20700
rect 15675 20650 15720 20700
rect 15770 20650 15815 20700
rect 15865 20650 15915 20700
rect 15965 20650 16015 20700
rect 16065 20650 16115 20700
rect 16165 20650 16210 20700
rect 16260 20650 16305 20700
rect 16355 20650 16425 20700
rect 16475 20650 16520 20700
rect 16570 20650 16615 20700
rect 16665 20650 16715 20700
rect 16765 20650 16815 20700
rect 16865 20650 16915 20700
rect 16965 20650 17010 20700
rect 17060 20650 17105 20700
rect 17155 20650 17225 20700
rect 17275 20650 17320 20700
rect 17370 20650 17415 20700
rect 17465 20650 17515 20700
rect 17565 20650 17615 20700
rect 17665 20650 17715 20700
rect 17765 20650 17810 20700
rect 17860 20650 17905 20700
rect 17955 20650 17990 20700
rect 14790 20610 17990 20650
rect 14790 20560 14825 20610
rect 14875 20560 14920 20610
rect 14970 20560 15015 20610
rect 15065 20560 15115 20610
rect 15165 20560 15215 20610
rect 15265 20560 15315 20610
rect 15365 20560 15410 20610
rect 15460 20560 15505 20610
rect 15555 20560 15625 20610
rect 15675 20560 15720 20610
rect 15770 20560 15815 20610
rect 15865 20560 15915 20610
rect 15965 20560 16015 20610
rect 16065 20560 16115 20610
rect 16165 20560 16210 20610
rect 16260 20560 16305 20610
rect 16355 20560 16425 20610
rect 16475 20560 16520 20610
rect 16570 20560 16615 20610
rect 16665 20560 16715 20610
rect 16765 20560 16815 20610
rect 16865 20560 16915 20610
rect 16965 20560 17010 20610
rect 17060 20560 17105 20610
rect 17155 20560 17225 20610
rect 17275 20560 17320 20610
rect 17370 20560 17415 20610
rect 17465 20560 17515 20610
rect 17565 20560 17615 20610
rect 17665 20560 17715 20610
rect 17765 20560 17810 20610
rect 17860 20560 17905 20610
rect 17955 20560 17990 20610
rect 14790 20490 17990 20560
rect 14790 20440 14825 20490
rect 14875 20440 14920 20490
rect 14970 20440 15015 20490
rect 15065 20440 15115 20490
rect 15165 20440 15215 20490
rect 15265 20440 15315 20490
rect 15365 20440 15410 20490
rect 15460 20440 15505 20490
rect 15555 20440 15625 20490
rect 15675 20440 15720 20490
rect 15770 20440 15815 20490
rect 15865 20440 15915 20490
rect 15965 20440 16015 20490
rect 16065 20440 16115 20490
rect 16165 20440 16210 20490
rect 16260 20440 16305 20490
rect 16355 20440 16425 20490
rect 16475 20440 16520 20490
rect 16570 20440 16615 20490
rect 16665 20440 16715 20490
rect 16765 20440 16815 20490
rect 16865 20440 16915 20490
rect 16965 20440 17010 20490
rect 17060 20440 17105 20490
rect 17155 20440 17225 20490
rect 17275 20440 17320 20490
rect 17370 20440 17415 20490
rect 17465 20440 17515 20490
rect 17565 20440 17615 20490
rect 17665 20440 17715 20490
rect 17765 20440 17810 20490
rect 17860 20440 17905 20490
rect 17955 20440 17990 20490
rect 14790 20400 17990 20440
rect 14790 20350 14825 20400
rect 14875 20350 14920 20400
rect 14970 20350 15015 20400
rect 15065 20350 15115 20400
rect 15165 20350 15215 20400
rect 15265 20350 15315 20400
rect 15365 20350 15410 20400
rect 15460 20350 15505 20400
rect 15555 20350 15625 20400
rect 15675 20350 15720 20400
rect 15770 20350 15815 20400
rect 15865 20350 15915 20400
rect 15965 20350 16015 20400
rect 16065 20350 16115 20400
rect 16165 20350 16210 20400
rect 16260 20350 16305 20400
rect 16355 20350 16425 20400
rect 16475 20350 16520 20400
rect 16570 20350 16615 20400
rect 16665 20350 16715 20400
rect 16765 20350 16815 20400
rect 16865 20350 16915 20400
rect 16965 20350 17010 20400
rect 17060 20350 17105 20400
rect 17155 20350 17225 20400
rect 17275 20350 17320 20400
rect 17370 20350 17415 20400
rect 17465 20350 17515 20400
rect 17565 20350 17615 20400
rect 17665 20350 17715 20400
rect 17765 20350 17810 20400
rect 17860 20350 17905 20400
rect 17955 20350 17990 20400
rect 14790 20300 17990 20350
rect 14790 20250 14825 20300
rect 14875 20250 14920 20300
rect 14970 20250 15015 20300
rect 15065 20250 15115 20300
rect 15165 20250 15215 20300
rect 15265 20250 15315 20300
rect 15365 20250 15410 20300
rect 15460 20250 15505 20300
rect 15555 20250 15625 20300
rect 15675 20250 15720 20300
rect 15770 20250 15815 20300
rect 15865 20250 15915 20300
rect 15965 20250 16015 20300
rect 16065 20250 16115 20300
rect 16165 20250 16210 20300
rect 16260 20250 16305 20300
rect 16355 20250 16425 20300
rect 16475 20250 16520 20300
rect 16570 20250 16615 20300
rect 16665 20250 16715 20300
rect 16765 20250 16815 20300
rect 16865 20250 16915 20300
rect 16965 20250 17010 20300
rect 17060 20250 17105 20300
rect 17155 20250 17225 20300
rect 17275 20250 17320 20300
rect 17370 20250 17415 20300
rect 17465 20250 17515 20300
rect 17565 20250 17615 20300
rect 17665 20250 17715 20300
rect 17765 20250 17810 20300
rect 17860 20250 17905 20300
rect 17955 20250 17990 20300
rect 14790 20210 17990 20250
rect 14790 20160 14825 20210
rect 14875 20160 14920 20210
rect 14970 20160 15015 20210
rect 15065 20160 15115 20210
rect 15165 20160 15215 20210
rect 15265 20160 15315 20210
rect 15365 20160 15410 20210
rect 15460 20160 15505 20210
rect 15555 20160 15625 20210
rect 15675 20160 15720 20210
rect 15770 20160 15815 20210
rect 15865 20160 15915 20210
rect 15965 20160 16015 20210
rect 16065 20160 16115 20210
rect 16165 20160 16210 20210
rect 16260 20160 16305 20210
rect 16355 20160 16425 20210
rect 16475 20160 16520 20210
rect 16570 20160 16615 20210
rect 16665 20160 16715 20210
rect 16765 20160 16815 20210
rect 16865 20160 16915 20210
rect 16965 20160 17010 20210
rect 17060 20160 17105 20210
rect 17155 20160 17225 20210
rect 17275 20160 17320 20210
rect 17370 20160 17415 20210
rect 17465 20160 17515 20210
rect 17565 20160 17615 20210
rect 17665 20160 17715 20210
rect 17765 20160 17810 20210
rect 17860 20160 17905 20210
rect 17955 20160 17990 20210
rect 14790 20090 17990 20160
rect 14790 20040 14825 20090
rect 14875 20040 14920 20090
rect 14970 20040 15015 20090
rect 15065 20040 15115 20090
rect 15165 20040 15215 20090
rect 15265 20040 15315 20090
rect 15365 20040 15410 20090
rect 15460 20040 15505 20090
rect 15555 20040 15625 20090
rect 15675 20040 15720 20090
rect 15770 20040 15815 20090
rect 15865 20040 15915 20090
rect 15965 20040 16015 20090
rect 16065 20040 16115 20090
rect 16165 20040 16210 20090
rect 16260 20040 16305 20090
rect 16355 20040 16425 20090
rect 16475 20040 16520 20090
rect 16570 20040 16615 20090
rect 16665 20040 16715 20090
rect 16765 20040 16815 20090
rect 16865 20040 16915 20090
rect 16965 20040 17010 20090
rect 17060 20040 17105 20090
rect 17155 20040 17225 20090
rect 17275 20040 17320 20090
rect 17370 20040 17415 20090
rect 17465 20040 17515 20090
rect 17565 20040 17615 20090
rect 17665 20040 17715 20090
rect 17765 20040 17810 20090
rect 17860 20040 17905 20090
rect 17955 20040 17990 20090
rect 14790 20000 17990 20040
rect 14790 19950 14825 20000
rect 14875 19950 14920 20000
rect 14970 19950 15015 20000
rect 15065 19950 15115 20000
rect 15165 19950 15215 20000
rect 15265 19950 15315 20000
rect 15365 19950 15410 20000
rect 15460 19950 15505 20000
rect 15555 19950 15625 20000
rect 15675 19950 15720 20000
rect 15770 19950 15815 20000
rect 15865 19950 15915 20000
rect 15965 19950 16015 20000
rect 16065 19950 16115 20000
rect 16165 19950 16210 20000
rect 16260 19950 16305 20000
rect 16355 19950 16425 20000
rect 16475 19950 16520 20000
rect 16570 19950 16615 20000
rect 16665 19950 16715 20000
rect 16765 19950 16815 20000
rect 16865 19950 16915 20000
rect 16965 19950 17010 20000
rect 17060 19950 17105 20000
rect 17155 19950 17225 20000
rect 17275 19950 17320 20000
rect 17370 19950 17415 20000
rect 17465 19950 17515 20000
rect 17565 19950 17615 20000
rect 17665 19950 17715 20000
rect 17765 19950 17810 20000
rect 17860 19950 17905 20000
rect 17955 19950 17990 20000
rect 14790 19900 17990 19950
rect 14790 19850 14825 19900
rect 14875 19850 14920 19900
rect 14970 19850 15015 19900
rect 15065 19850 15115 19900
rect 15165 19850 15215 19900
rect 15265 19850 15315 19900
rect 15365 19850 15410 19900
rect 15460 19850 15505 19900
rect 15555 19850 15625 19900
rect 15675 19850 15720 19900
rect 15770 19850 15815 19900
rect 15865 19850 15915 19900
rect 15965 19850 16015 19900
rect 16065 19850 16115 19900
rect 16165 19850 16210 19900
rect 16260 19850 16305 19900
rect 16355 19850 16425 19900
rect 16475 19850 16520 19900
rect 16570 19850 16615 19900
rect 16665 19850 16715 19900
rect 16765 19850 16815 19900
rect 16865 19850 16915 19900
rect 16965 19850 17010 19900
rect 17060 19850 17105 19900
rect 17155 19850 17225 19900
rect 17275 19850 17320 19900
rect 17370 19850 17415 19900
rect 17465 19850 17515 19900
rect 17565 19850 17615 19900
rect 17665 19850 17715 19900
rect 17765 19850 17810 19900
rect 17860 19850 17905 19900
rect 17955 19850 17990 19900
rect 14790 19810 17990 19850
rect 14790 19760 14825 19810
rect 14875 19760 14920 19810
rect 14970 19760 15015 19810
rect 15065 19760 15115 19810
rect 15165 19760 15215 19810
rect 15265 19760 15315 19810
rect 15365 19760 15410 19810
rect 15460 19760 15505 19810
rect 15555 19760 15625 19810
rect 15675 19760 15720 19810
rect 15770 19760 15815 19810
rect 15865 19760 15915 19810
rect 15965 19760 16015 19810
rect 16065 19760 16115 19810
rect 16165 19760 16210 19810
rect 16260 19760 16305 19810
rect 16355 19760 16425 19810
rect 16475 19760 16520 19810
rect 16570 19760 16615 19810
rect 16665 19760 16715 19810
rect 16765 19760 16815 19810
rect 16865 19760 16915 19810
rect 16965 19760 17010 19810
rect 17060 19760 17105 19810
rect 17155 19760 17225 19810
rect 17275 19760 17320 19810
rect 17370 19760 17415 19810
rect 17465 19760 17515 19810
rect 17565 19760 17615 19810
rect 17665 19760 17715 19810
rect 17765 19760 17810 19810
rect 17860 19760 17905 19810
rect 17955 19760 17990 19810
rect 14790 19690 17990 19760
rect 14790 19640 14825 19690
rect 14875 19640 14920 19690
rect 14970 19640 15015 19690
rect 15065 19640 15115 19690
rect 15165 19640 15215 19690
rect 15265 19640 15315 19690
rect 15365 19640 15410 19690
rect 15460 19640 15505 19690
rect 15555 19640 15625 19690
rect 15675 19640 15720 19690
rect 15770 19640 15815 19690
rect 15865 19640 15915 19690
rect 15965 19640 16015 19690
rect 16065 19640 16115 19690
rect 16165 19640 16210 19690
rect 16260 19640 16305 19690
rect 16355 19640 16425 19690
rect 16475 19640 16520 19690
rect 16570 19640 16615 19690
rect 16665 19640 16715 19690
rect 16765 19640 16815 19690
rect 16865 19640 16915 19690
rect 16965 19640 17010 19690
rect 17060 19640 17105 19690
rect 17155 19640 17225 19690
rect 17275 19640 17320 19690
rect 17370 19640 17415 19690
rect 17465 19640 17515 19690
rect 17565 19640 17615 19690
rect 17665 19640 17715 19690
rect 17765 19640 17810 19690
rect 17860 19640 17905 19690
rect 17955 19640 17990 19690
rect 14790 19600 17990 19640
rect 14790 19550 14825 19600
rect 14875 19550 14920 19600
rect 14970 19550 15015 19600
rect 15065 19550 15115 19600
rect 15165 19550 15215 19600
rect 15265 19550 15315 19600
rect 15365 19550 15410 19600
rect 15460 19550 15505 19600
rect 15555 19550 15625 19600
rect 15675 19550 15720 19600
rect 15770 19550 15815 19600
rect 15865 19550 15915 19600
rect 15965 19550 16015 19600
rect 16065 19550 16115 19600
rect 16165 19550 16210 19600
rect 16260 19550 16305 19600
rect 16355 19550 16425 19600
rect 16475 19550 16520 19600
rect 16570 19550 16615 19600
rect 16665 19550 16715 19600
rect 16765 19550 16815 19600
rect 16865 19550 16915 19600
rect 16965 19550 17010 19600
rect 17060 19550 17105 19600
rect 17155 19550 17225 19600
rect 17275 19550 17320 19600
rect 17370 19550 17415 19600
rect 17465 19550 17515 19600
rect 17565 19550 17615 19600
rect 17665 19550 17715 19600
rect 17765 19550 17810 19600
rect 17860 19550 17905 19600
rect 17955 19550 17990 19600
rect 14790 19500 17990 19550
rect 14790 19450 14825 19500
rect 14875 19450 14920 19500
rect 14970 19450 15015 19500
rect 15065 19450 15115 19500
rect 15165 19450 15215 19500
rect 15265 19450 15315 19500
rect 15365 19450 15410 19500
rect 15460 19450 15505 19500
rect 15555 19450 15625 19500
rect 15675 19450 15720 19500
rect 15770 19450 15815 19500
rect 15865 19450 15915 19500
rect 15965 19450 16015 19500
rect 16065 19450 16115 19500
rect 16165 19450 16210 19500
rect 16260 19450 16305 19500
rect 16355 19450 16425 19500
rect 16475 19450 16520 19500
rect 16570 19450 16615 19500
rect 16665 19450 16715 19500
rect 16765 19450 16815 19500
rect 16865 19450 16915 19500
rect 16965 19450 17010 19500
rect 17060 19450 17105 19500
rect 17155 19450 17225 19500
rect 17275 19450 17320 19500
rect 17370 19450 17415 19500
rect 17465 19450 17515 19500
rect 17565 19450 17615 19500
rect 17665 19450 17715 19500
rect 17765 19450 17810 19500
rect 17860 19450 17905 19500
rect 17955 19450 17990 19500
rect 14790 19410 17990 19450
rect 14790 19360 14825 19410
rect 14875 19360 14920 19410
rect 14970 19360 15015 19410
rect 15065 19360 15115 19410
rect 15165 19360 15215 19410
rect 15265 19360 15315 19410
rect 15365 19360 15410 19410
rect 15460 19360 15505 19410
rect 15555 19360 15625 19410
rect 15675 19360 15720 19410
rect 15770 19360 15815 19410
rect 15865 19360 15915 19410
rect 15965 19360 16015 19410
rect 16065 19360 16115 19410
rect 16165 19360 16210 19410
rect 16260 19360 16305 19410
rect 16355 19360 16425 19410
rect 16475 19360 16520 19410
rect 16570 19360 16615 19410
rect 16665 19360 16715 19410
rect 16765 19360 16815 19410
rect 16865 19360 16915 19410
rect 16965 19360 17010 19410
rect 17060 19360 17105 19410
rect 17155 19360 17225 19410
rect 17275 19360 17320 19410
rect 17370 19360 17415 19410
rect 17465 19360 17515 19410
rect 17565 19360 17615 19410
rect 17665 19360 17715 19410
rect 17765 19360 17810 19410
rect 17860 19360 17905 19410
rect 17955 19360 17990 19410
rect 14790 19290 17990 19360
rect 14790 19240 14825 19290
rect 14875 19240 14920 19290
rect 14970 19240 15015 19290
rect 15065 19240 15115 19290
rect 15165 19240 15215 19290
rect 15265 19240 15315 19290
rect 15365 19240 15410 19290
rect 15460 19240 15505 19290
rect 15555 19240 15625 19290
rect 15675 19240 15720 19290
rect 15770 19240 15815 19290
rect 15865 19240 15915 19290
rect 15965 19240 16015 19290
rect 16065 19240 16115 19290
rect 16165 19240 16210 19290
rect 16260 19240 16305 19290
rect 16355 19240 16425 19290
rect 16475 19240 16520 19290
rect 16570 19240 16615 19290
rect 16665 19240 16715 19290
rect 16765 19240 16815 19290
rect 16865 19240 16915 19290
rect 16965 19240 17010 19290
rect 17060 19240 17105 19290
rect 17155 19240 17225 19290
rect 17275 19240 17320 19290
rect 17370 19240 17415 19290
rect 17465 19240 17515 19290
rect 17565 19240 17615 19290
rect 17665 19240 17715 19290
rect 17765 19240 17810 19290
rect 17860 19240 17905 19290
rect 17955 19240 17990 19290
rect 14790 19200 17990 19240
rect 14790 19150 14825 19200
rect 14875 19150 14920 19200
rect 14970 19150 15015 19200
rect 15065 19150 15115 19200
rect 15165 19150 15215 19200
rect 15265 19150 15315 19200
rect 15365 19150 15410 19200
rect 15460 19150 15505 19200
rect 15555 19150 15625 19200
rect 15675 19150 15720 19200
rect 15770 19150 15815 19200
rect 15865 19150 15915 19200
rect 15965 19150 16015 19200
rect 16065 19150 16115 19200
rect 16165 19150 16210 19200
rect 16260 19150 16305 19200
rect 16355 19150 16425 19200
rect 16475 19150 16520 19200
rect 16570 19150 16615 19200
rect 16665 19150 16715 19200
rect 16765 19150 16815 19200
rect 16865 19150 16915 19200
rect 16965 19150 17010 19200
rect 17060 19150 17105 19200
rect 17155 19150 17225 19200
rect 17275 19150 17320 19200
rect 17370 19150 17415 19200
rect 17465 19150 17515 19200
rect 17565 19150 17615 19200
rect 17665 19150 17715 19200
rect 17765 19150 17810 19200
rect 17860 19150 17905 19200
rect 17955 19150 17990 19200
rect 14790 19100 17990 19150
rect 14790 19050 14825 19100
rect 14875 19050 14920 19100
rect 14970 19050 15015 19100
rect 15065 19050 15115 19100
rect 15165 19050 15215 19100
rect 15265 19050 15315 19100
rect 15365 19050 15410 19100
rect 15460 19050 15505 19100
rect 15555 19050 15625 19100
rect 15675 19050 15720 19100
rect 15770 19050 15815 19100
rect 15865 19050 15915 19100
rect 15965 19050 16015 19100
rect 16065 19050 16115 19100
rect 16165 19050 16210 19100
rect 16260 19050 16305 19100
rect 16355 19050 16425 19100
rect 16475 19050 16520 19100
rect 16570 19050 16615 19100
rect 16665 19050 16715 19100
rect 16765 19050 16815 19100
rect 16865 19050 16915 19100
rect 16965 19050 17010 19100
rect 17060 19050 17105 19100
rect 17155 19050 17225 19100
rect 17275 19050 17320 19100
rect 17370 19050 17415 19100
rect 17465 19050 17515 19100
rect 17565 19050 17615 19100
rect 17665 19050 17715 19100
rect 17765 19050 17810 19100
rect 17860 19050 17905 19100
rect 17955 19050 17990 19100
rect 14790 19010 17990 19050
rect 14790 18960 14825 19010
rect 14875 18960 14920 19010
rect 14970 18960 15015 19010
rect 15065 18960 15115 19010
rect 15165 18960 15215 19010
rect 15265 18960 15315 19010
rect 15365 18960 15410 19010
rect 15460 18960 15505 19010
rect 15555 18960 15625 19010
rect 15675 18960 15720 19010
rect 15770 18960 15815 19010
rect 15865 18960 15915 19010
rect 15965 18960 16015 19010
rect 16065 18960 16115 19010
rect 16165 18960 16210 19010
rect 16260 18960 16305 19010
rect 16355 18960 16425 19010
rect 16475 18960 16520 19010
rect 16570 18960 16615 19010
rect 16665 18960 16715 19010
rect 16765 18960 16815 19010
rect 16865 18960 16915 19010
rect 16965 18960 17010 19010
rect 17060 18960 17105 19010
rect 17155 18960 17225 19010
rect 17275 18960 17320 19010
rect 17370 18960 17415 19010
rect 17465 18960 17515 19010
rect 17565 18960 17615 19010
rect 17665 18960 17715 19010
rect 17765 18960 17810 19010
rect 17860 18960 17905 19010
rect 17955 18960 17990 19010
rect 14790 18890 17990 18960
rect 14790 18840 14825 18890
rect 14875 18840 14920 18890
rect 14970 18840 15015 18890
rect 15065 18840 15115 18890
rect 15165 18840 15215 18890
rect 15265 18840 15315 18890
rect 15365 18840 15410 18890
rect 15460 18840 15505 18890
rect 15555 18840 15625 18890
rect 15675 18840 15720 18890
rect 15770 18840 15815 18890
rect 15865 18840 15915 18890
rect 15965 18840 16015 18890
rect 16065 18840 16115 18890
rect 16165 18840 16210 18890
rect 16260 18840 16305 18890
rect 16355 18840 16425 18890
rect 16475 18840 16520 18890
rect 16570 18840 16615 18890
rect 16665 18840 16715 18890
rect 16765 18840 16815 18890
rect 16865 18840 16915 18890
rect 16965 18840 17010 18890
rect 17060 18840 17105 18890
rect 17155 18840 17225 18890
rect 17275 18840 17320 18890
rect 17370 18840 17415 18890
rect 17465 18840 17515 18890
rect 17565 18840 17615 18890
rect 17665 18840 17715 18890
rect 17765 18840 17810 18890
rect 17860 18840 17905 18890
rect 17955 18840 17990 18890
rect 14790 18800 17990 18840
rect 14790 18750 14825 18800
rect 14875 18750 14920 18800
rect 14970 18750 15015 18800
rect 15065 18750 15115 18800
rect 15165 18750 15215 18800
rect 15265 18750 15315 18800
rect 15365 18750 15410 18800
rect 15460 18750 15505 18800
rect 15555 18750 15625 18800
rect 15675 18750 15720 18800
rect 15770 18750 15815 18800
rect 15865 18750 15915 18800
rect 15965 18750 16015 18800
rect 16065 18750 16115 18800
rect 16165 18750 16210 18800
rect 16260 18750 16305 18800
rect 16355 18750 16425 18800
rect 16475 18750 16520 18800
rect 16570 18750 16615 18800
rect 16665 18750 16715 18800
rect 16765 18750 16815 18800
rect 16865 18750 16915 18800
rect 16965 18750 17010 18800
rect 17060 18750 17105 18800
rect 17155 18750 17225 18800
rect 17275 18750 17320 18800
rect 17370 18750 17415 18800
rect 17465 18750 17515 18800
rect 17565 18750 17615 18800
rect 17665 18750 17715 18800
rect 17765 18750 17810 18800
rect 17860 18750 17905 18800
rect 17955 18750 17990 18800
rect 14790 18700 17990 18750
rect 14790 18650 14825 18700
rect 14875 18650 14920 18700
rect 14970 18650 15015 18700
rect 15065 18650 15115 18700
rect 15165 18650 15215 18700
rect 15265 18650 15315 18700
rect 15365 18650 15410 18700
rect 15460 18650 15505 18700
rect 15555 18650 15625 18700
rect 15675 18650 15720 18700
rect 15770 18650 15815 18700
rect 15865 18650 15915 18700
rect 15965 18650 16015 18700
rect 16065 18650 16115 18700
rect 16165 18650 16210 18700
rect 16260 18650 16305 18700
rect 16355 18650 16425 18700
rect 16475 18650 16520 18700
rect 16570 18650 16615 18700
rect 16665 18650 16715 18700
rect 16765 18650 16815 18700
rect 16865 18650 16915 18700
rect 16965 18650 17010 18700
rect 17060 18650 17105 18700
rect 17155 18650 17225 18700
rect 17275 18650 17320 18700
rect 17370 18650 17415 18700
rect 17465 18650 17515 18700
rect 17565 18650 17615 18700
rect 17665 18650 17715 18700
rect 17765 18650 17810 18700
rect 17860 18650 17905 18700
rect 17955 18650 17990 18700
rect 14790 18610 17990 18650
rect 14790 18560 14825 18610
rect 14875 18560 14920 18610
rect 14970 18560 15015 18610
rect 15065 18560 15115 18610
rect 15165 18560 15215 18610
rect 15265 18560 15315 18610
rect 15365 18560 15410 18610
rect 15460 18560 15505 18610
rect 15555 18560 15625 18610
rect 15675 18560 15720 18610
rect 15770 18560 15815 18610
rect 15865 18560 15915 18610
rect 15965 18560 16015 18610
rect 16065 18560 16115 18610
rect 16165 18560 16210 18610
rect 16260 18560 16305 18610
rect 16355 18560 16425 18610
rect 16475 18560 16520 18610
rect 16570 18560 16615 18610
rect 16665 18560 16715 18610
rect 16765 18560 16815 18610
rect 16865 18560 16915 18610
rect 16965 18560 17010 18610
rect 17060 18560 17105 18610
rect 17155 18560 17225 18610
rect 17275 18560 17320 18610
rect 17370 18560 17415 18610
rect 17465 18560 17515 18610
rect 17565 18560 17615 18610
rect 17665 18560 17715 18610
rect 17765 18560 17810 18610
rect 17860 18560 17905 18610
rect 17955 18560 17990 18610
rect 14790 18490 17990 18560
rect 14790 18440 14825 18490
rect 14875 18440 14920 18490
rect 14970 18440 15015 18490
rect 15065 18440 15115 18490
rect 15165 18440 15215 18490
rect 15265 18440 15315 18490
rect 15365 18440 15410 18490
rect 15460 18440 15505 18490
rect 15555 18440 15625 18490
rect 15675 18440 15720 18490
rect 15770 18440 15815 18490
rect 15865 18440 15915 18490
rect 15965 18440 16015 18490
rect 16065 18440 16115 18490
rect 16165 18440 16210 18490
rect 16260 18440 16305 18490
rect 16355 18440 16425 18490
rect 16475 18440 16520 18490
rect 16570 18440 16615 18490
rect 16665 18440 16715 18490
rect 16765 18440 16815 18490
rect 16865 18440 16915 18490
rect 16965 18440 17010 18490
rect 17060 18440 17105 18490
rect 17155 18440 17225 18490
rect 17275 18440 17320 18490
rect 17370 18440 17415 18490
rect 17465 18440 17515 18490
rect 17565 18440 17615 18490
rect 17665 18440 17715 18490
rect 17765 18440 17810 18490
rect 17860 18440 17905 18490
rect 17955 18440 17990 18490
rect 14790 18400 17990 18440
rect 14790 18350 14825 18400
rect 14875 18350 14920 18400
rect 14970 18350 15015 18400
rect 15065 18350 15115 18400
rect 15165 18350 15215 18400
rect 15265 18350 15315 18400
rect 15365 18350 15410 18400
rect 15460 18350 15505 18400
rect 15555 18350 15625 18400
rect 15675 18350 15720 18400
rect 15770 18350 15815 18400
rect 15865 18350 15915 18400
rect 15965 18350 16015 18400
rect 16065 18350 16115 18400
rect 16165 18350 16210 18400
rect 16260 18350 16305 18400
rect 16355 18350 16425 18400
rect 16475 18350 16520 18400
rect 16570 18350 16615 18400
rect 16665 18350 16715 18400
rect 16765 18350 16815 18400
rect 16865 18350 16915 18400
rect 16965 18350 17010 18400
rect 17060 18350 17105 18400
rect 17155 18350 17225 18400
rect 17275 18350 17320 18400
rect 17370 18350 17415 18400
rect 17465 18350 17515 18400
rect 17565 18350 17615 18400
rect 17665 18350 17715 18400
rect 17765 18350 17810 18400
rect 17860 18350 17905 18400
rect 17955 18350 17990 18400
rect 14790 18300 17990 18350
rect 14790 18250 14825 18300
rect 14875 18250 14920 18300
rect 14970 18250 15015 18300
rect 15065 18250 15115 18300
rect 15165 18250 15215 18300
rect 15265 18250 15315 18300
rect 15365 18250 15410 18300
rect 15460 18250 15505 18300
rect 15555 18250 15625 18300
rect 15675 18250 15720 18300
rect 15770 18250 15815 18300
rect 15865 18250 15915 18300
rect 15965 18250 16015 18300
rect 16065 18250 16115 18300
rect 16165 18250 16210 18300
rect 16260 18250 16305 18300
rect 16355 18250 16425 18300
rect 16475 18250 16520 18300
rect 16570 18250 16615 18300
rect 16665 18250 16715 18300
rect 16765 18250 16815 18300
rect 16865 18250 16915 18300
rect 16965 18250 17010 18300
rect 17060 18250 17105 18300
rect 17155 18250 17225 18300
rect 17275 18250 17320 18300
rect 17370 18250 17415 18300
rect 17465 18250 17515 18300
rect 17565 18250 17615 18300
rect 17665 18250 17715 18300
rect 17765 18250 17810 18300
rect 17860 18250 17905 18300
rect 17955 18250 17990 18300
rect 14790 18210 17990 18250
rect 14790 18160 14825 18210
rect 14875 18160 14920 18210
rect 14970 18160 15015 18210
rect 15065 18160 15115 18210
rect 15165 18160 15215 18210
rect 15265 18160 15315 18210
rect 15365 18160 15410 18210
rect 15460 18160 15505 18210
rect 15555 18160 15625 18210
rect 15675 18160 15720 18210
rect 15770 18160 15815 18210
rect 15865 18160 15915 18210
rect 15965 18160 16015 18210
rect 16065 18160 16115 18210
rect 16165 18160 16210 18210
rect 16260 18160 16305 18210
rect 16355 18160 16425 18210
rect 16475 18160 16520 18210
rect 16570 18160 16615 18210
rect 16665 18160 16715 18210
rect 16765 18160 16815 18210
rect 16865 18160 16915 18210
rect 16965 18160 17010 18210
rect 17060 18160 17105 18210
rect 17155 18160 17225 18210
rect 17275 18160 17320 18210
rect 17370 18160 17415 18210
rect 17465 18160 17515 18210
rect 17565 18160 17615 18210
rect 17665 18160 17715 18210
rect 17765 18160 17810 18210
rect 17860 18160 17905 18210
rect 17955 18160 17990 18210
rect 14790 18090 17990 18160
rect 14790 18040 14825 18090
rect 14875 18040 14920 18090
rect 14970 18040 15015 18090
rect 15065 18040 15115 18090
rect 15165 18040 15215 18090
rect 15265 18040 15315 18090
rect 15365 18040 15410 18090
rect 15460 18040 15505 18090
rect 15555 18040 15625 18090
rect 15675 18040 15720 18090
rect 15770 18040 15815 18090
rect 15865 18040 15915 18090
rect 15965 18040 16015 18090
rect 16065 18040 16115 18090
rect 16165 18040 16210 18090
rect 16260 18040 16305 18090
rect 16355 18040 16425 18090
rect 16475 18040 16520 18090
rect 16570 18040 16615 18090
rect 16665 18040 16715 18090
rect 16765 18040 16815 18090
rect 16865 18040 16915 18090
rect 16965 18040 17010 18090
rect 17060 18040 17105 18090
rect 17155 18040 17225 18090
rect 17275 18040 17320 18090
rect 17370 18040 17415 18090
rect 17465 18040 17515 18090
rect 17565 18040 17615 18090
rect 17665 18040 17715 18090
rect 17765 18040 17810 18090
rect 17860 18040 17905 18090
rect 17955 18040 17990 18090
rect 14790 18000 17990 18040
rect 14790 17950 14825 18000
rect 14875 17950 14920 18000
rect 14970 17950 15015 18000
rect 15065 17950 15115 18000
rect 15165 17950 15215 18000
rect 15265 17950 15315 18000
rect 15365 17950 15410 18000
rect 15460 17950 15505 18000
rect 15555 17950 15625 18000
rect 15675 17950 15720 18000
rect 15770 17950 15815 18000
rect 15865 17950 15915 18000
rect 15965 17950 16015 18000
rect 16065 17950 16115 18000
rect 16165 17950 16210 18000
rect 16260 17950 16305 18000
rect 16355 17950 16425 18000
rect 16475 17950 16520 18000
rect 16570 17950 16615 18000
rect 16665 17950 16715 18000
rect 16765 17950 16815 18000
rect 16865 17950 16915 18000
rect 16965 17950 17010 18000
rect 17060 17950 17105 18000
rect 17155 17950 17225 18000
rect 17275 17950 17320 18000
rect 17370 17950 17415 18000
rect 17465 17950 17515 18000
rect 17565 17950 17615 18000
rect 17665 17950 17715 18000
rect 17765 17950 17810 18000
rect 17860 17950 17905 18000
rect 17955 17950 17990 18000
rect 14790 17900 17990 17950
rect 14790 17850 14825 17900
rect 14875 17850 14920 17900
rect 14970 17850 15015 17900
rect 15065 17850 15115 17900
rect 15165 17850 15215 17900
rect 15265 17850 15315 17900
rect 15365 17850 15410 17900
rect 15460 17850 15505 17900
rect 15555 17850 15625 17900
rect 15675 17850 15720 17900
rect 15770 17850 15815 17900
rect 15865 17850 15915 17900
rect 15965 17850 16015 17900
rect 16065 17850 16115 17900
rect 16165 17850 16210 17900
rect 16260 17850 16305 17900
rect 16355 17850 16425 17900
rect 16475 17850 16520 17900
rect 16570 17850 16615 17900
rect 16665 17850 16715 17900
rect 16765 17850 16815 17900
rect 16865 17850 16915 17900
rect 16965 17850 17010 17900
rect 17060 17850 17105 17900
rect 17155 17850 17225 17900
rect 17275 17850 17320 17900
rect 17370 17850 17415 17900
rect 17465 17850 17515 17900
rect 17565 17850 17615 17900
rect 17665 17850 17715 17900
rect 17765 17850 17810 17900
rect 17860 17850 17905 17900
rect 17955 17850 17990 17900
rect 14790 17810 17990 17850
rect 14790 17760 14825 17810
rect 14875 17760 14920 17810
rect 14970 17760 15015 17810
rect 15065 17760 15115 17810
rect 15165 17760 15215 17810
rect 15265 17760 15315 17810
rect 15365 17760 15410 17810
rect 15460 17760 15505 17810
rect 15555 17760 15625 17810
rect 15675 17760 15720 17810
rect 15770 17760 15815 17810
rect 15865 17760 15915 17810
rect 15965 17760 16015 17810
rect 16065 17760 16115 17810
rect 16165 17760 16210 17810
rect 16260 17760 16305 17810
rect 16355 17760 16425 17810
rect 16475 17760 16520 17810
rect 16570 17760 16615 17810
rect 16665 17760 16715 17810
rect 16765 17760 16815 17810
rect 16865 17760 16915 17810
rect 16965 17760 17010 17810
rect 17060 17760 17105 17810
rect 17155 17760 17225 17810
rect 17275 17760 17320 17810
rect 17370 17760 17415 17810
rect 17465 17760 17515 17810
rect 17565 17760 17615 17810
rect 17665 17760 17715 17810
rect 17765 17760 17810 17810
rect 17860 17760 17905 17810
rect 17955 17760 17990 17810
rect 230 17530 280 17650
rect -1260 17445 -1030 17530
rect -910 17445 -680 17530
rect -560 17445 -330 17530
rect -210 17445 20 17530
rect 140 17445 370 17530
rect 490 17445 720 17530
rect 840 17445 1070 17530
rect 1190 17445 1420 17530
rect 1540 17445 1770 17530
rect -1260 17395 1770 17445
rect -1260 17300 -1030 17395
rect -910 17300 -680 17395
rect -560 17300 -330 17395
rect -210 17300 20 17395
rect 140 17300 370 17395
rect 490 17300 720 17395
rect 840 17300 1070 17395
rect 1190 17300 1420 17395
rect 1540 17300 1770 17395
rect 9540 17445 9770 17530
rect 9890 17445 10120 17530
rect 10240 17445 10470 17530
rect 10590 17445 10820 17530
rect 10940 17445 11170 17530
rect 11290 17445 11520 17530
rect 11640 17445 11870 17530
rect 11990 17445 12220 17530
rect 12340 17445 12570 17530
rect 12690 17445 12920 17530
rect 13040 17445 13270 17530
rect 13390 17445 13620 17530
rect 13740 17445 13970 17530
rect 14090 17445 14320 17530
rect 14440 17445 14670 17530
rect 14790 17445 17990 17760
rect 9540 17395 17990 17445
rect 9540 17300 9770 17395
rect 9890 17300 10120 17395
rect 10240 17300 10470 17395
rect 10590 17300 10820 17395
rect 10940 17300 11170 17395
rect 11290 17300 11520 17395
rect 11640 17300 11870 17395
rect 11990 17300 12220 17395
rect 12340 17300 12570 17395
rect 12690 17300 12920 17395
rect 13040 17300 13270 17395
rect 13390 17300 13620 17395
rect 13740 17300 13970 17395
rect 14090 17300 14320 17395
rect 14440 17300 14670 17395
rect 230 17180 280 17300
rect 12080 17180 12130 17300
rect -1260 17095 -1030 17180
rect -910 17095 -680 17180
rect -560 17095 -330 17180
rect -210 17095 20 17180
rect 140 17095 370 17180
rect 490 17095 720 17180
rect 840 17095 1070 17180
rect 1190 17095 1420 17180
rect 1540 17095 1770 17180
rect -1260 17045 1770 17095
rect -1260 16950 -1030 17045
rect -910 16950 -680 17045
rect -560 16950 -330 17045
rect -210 16950 20 17045
rect 140 16950 370 17045
rect 490 16950 720 17045
rect 840 16950 1070 17045
rect 1190 16950 1420 17045
rect 1540 16950 1770 17045
rect 9540 17095 9770 17180
rect 9890 17095 10120 17180
rect 10240 17095 10470 17180
rect 10590 17095 10820 17180
rect 10940 17095 11170 17180
rect 11290 17095 11520 17180
rect 11640 17095 11870 17180
rect 11990 17095 12220 17180
rect 12340 17095 12570 17180
rect 12690 17095 12920 17180
rect 13040 17095 13270 17180
rect 13390 17095 13620 17180
rect 13740 17095 13970 17180
rect 14090 17095 14320 17180
rect 14440 17095 14670 17180
rect 9540 17045 14670 17095
rect 9540 16950 9770 17045
rect 9890 16950 10120 17045
rect 10240 16950 10470 17045
rect 10590 16950 10820 17045
rect 10940 16950 11170 17045
rect 11290 16950 11520 17045
rect 11640 16950 11870 17045
rect 11990 16950 12220 17045
rect 12340 16950 12570 17045
rect 12690 16950 12920 17045
rect 13040 16950 13270 17045
rect 13390 16950 13620 17045
rect 13740 16950 13970 17045
rect 14090 16950 14320 17045
rect 14440 16950 14670 17045
rect 230 16830 280 16950
rect 12080 16830 12130 16950
rect -1260 16745 -1030 16830
rect -910 16745 -680 16830
rect -560 16745 -330 16830
rect -210 16745 20 16830
rect 140 16745 370 16830
rect 490 16745 720 16830
rect 840 16745 1070 16830
rect 1190 16745 1420 16830
rect 1540 16745 1770 16830
rect -1260 16695 1770 16745
rect -1260 16600 -1030 16695
rect -910 16600 -680 16695
rect -560 16600 -330 16695
rect -210 16600 20 16695
rect 140 16600 370 16695
rect 490 16600 720 16695
rect 840 16600 1070 16695
rect 1190 16600 1420 16695
rect 1540 16600 1770 16695
rect 9540 16745 9770 16830
rect 9890 16745 10120 16830
rect 10240 16745 10470 16830
rect 10590 16745 10820 16830
rect 10940 16745 11170 16830
rect 11290 16745 11520 16830
rect 11640 16745 11870 16830
rect 11990 16745 12220 16830
rect 12340 16745 12570 16830
rect 12690 16745 12920 16830
rect 13040 16745 13270 16830
rect 13390 16745 13620 16830
rect 13740 16745 13970 16830
rect 14090 16745 14320 16830
rect 14440 16745 14670 16830
rect 9540 16695 14670 16745
rect 9540 16600 9770 16695
rect 9890 16600 10120 16695
rect 10240 16600 10470 16695
rect 10590 16600 10820 16695
rect 10940 16600 11170 16695
rect 11290 16600 11520 16695
rect 11640 16600 11870 16695
rect 11990 16600 12220 16695
rect 12340 16600 12570 16695
rect 12690 16600 12920 16695
rect 13040 16600 13270 16695
rect 13390 16600 13620 16695
rect 13740 16600 13970 16695
rect 14090 16600 14320 16695
rect 14440 16600 14670 16695
rect 230 16480 280 16600
rect 12080 16480 12130 16600
rect -1260 16395 -1030 16480
rect -910 16395 -680 16480
rect -560 16395 -330 16480
rect -210 16395 20 16480
rect 140 16395 370 16480
rect 490 16395 720 16480
rect 840 16395 1070 16480
rect 1190 16395 1420 16480
rect 1540 16395 1770 16480
rect -1260 16345 1770 16395
rect -1260 16250 -1030 16345
rect -910 16250 -680 16345
rect -560 16250 -330 16345
rect -210 16250 20 16345
rect 140 16250 370 16345
rect 490 16250 720 16345
rect 840 16250 1070 16345
rect 1190 16250 1420 16345
rect 1540 16250 1770 16345
rect 9540 16395 9770 16480
rect 9890 16395 10120 16480
rect 10240 16395 10470 16480
rect 10590 16395 10820 16480
rect 10940 16395 11170 16480
rect 11290 16395 11520 16480
rect 11640 16395 11870 16480
rect 11990 16395 12220 16480
rect 12340 16395 12570 16480
rect 12690 16395 12920 16480
rect 13040 16395 13270 16480
rect 13390 16395 13620 16480
rect 13740 16395 13970 16480
rect 14090 16395 14320 16480
rect 14440 16395 14670 16480
rect 9540 16345 14670 16395
rect 9540 16250 9770 16345
rect 9890 16250 10120 16345
rect 10240 16250 10470 16345
rect 10590 16250 10820 16345
rect 10940 16250 11170 16345
rect 11290 16250 11520 16345
rect 11640 16250 11870 16345
rect 11990 16250 12220 16345
rect 12340 16250 12570 16345
rect 12690 16250 12920 16345
rect 13040 16250 13270 16345
rect 13390 16250 13620 16345
rect 13740 16250 13970 16345
rect 14090 16250 14320 16345
rect 14440 16250 14670 16345
rect 230 16130 280 16250
rect 12080 16130 12130 16250
rect -1260 16045 -1030 16130
rect -910 16045 -680 16130
rect -560 16045 -330 16130
rect -210 16045 20 16130
rect 140 16045 370 16130
rect 490 16045 720 16130
rect 840 16045 1070 16130
rect 1190 16045 1420 16130
rect 1540 16045 1770 16130
rect -1260 15995 1770 16045
rect -1260 15900 -1030 15995
rect -910 15900 -680 15995
rect -560 15900 -330 15995
rect -210 15900 20 15995
rect 140 15900 370 15995
rect 490 15900 720 15995
rect 840 15900 1070 15995
rect 1190 15900 1420 15995
rect 1540 15900 1770 15995
rect 9540 16045 9770 16130
rect 9890 16045 10120 16130
rect 10240 16045 10470 16130
rect 10590 16045 10820 16130
rect 10940 16045 11170 16130
rect 11290 16045 11520 16130
rect 11640 16045 11870 16130
rect 11990 16045 12220 16130
rect 12340 16045 12570 16130
rect 12690 16045 12920 16130
rect 13040 16045 13270 16130
rect 13390 16045 13620 16130
rect 13740 16045 13970 16130
rect 14090 16045 14320 16130
rect 14440 16045 14670 16130
rect 9540 15995 14670 16045
rect 9540 15900 9770 15995
rect 9890 15900 10120 15995
rect 10240 15900 10470 15995
rect 10590 15900 10820 15995
rect 10940 15900 11170 15995
rect 11290 15900 11520 15995
rect 11640 15900 11870 15995
rect 11990 15900 12220 15995
rect 12340 15900 12570 15995
rect 12690 15900 12920 15995
rect 13040 15900 13270 15995
rect 13390 15900 13620 15995
rect 13740 15900 13970 15995
rect 14090 15900 14320 15995
rect 14440 15900 14670 15995
rect 230 15780 280 15900
rect 12080 15780 12130 15900
rect -1260 15695 -1030 15780
rect -910 15695 -680 15780
rect -560 15695 -330 15780
rect -210 15695 20 15780
rect 140 15695 370 15780
rect 490 15695 720 15780
rect 840 15695 1070 15780
rect 1190 15695 1420 15780
rect 1540 15695 1770 15780
rect -1260 15645 1770 15695
rect -1260 15550 -1030 15645
rect -910 15550 -680 15645
rect -560 15550 -330 15645
rect -210 15550 20 15645
rect 140 15550 370 15645
rect 490 15550 720 15645
rect 840 15550 1070 15645
rect 1190 15550 1420 15645
rect 1540 15550 1770 15645
rect 9540 15695 9770 15780
rect 9890 15695 10120 15780
rect 10240 15695 10470 15780
rect 10590 15695 10820 15780
rect 10940 15695 11170 15780
rect 11290 15695 11520 15780
rect 11640 15695 11870 15780
rect 11990 15695 12220 15780
rect 12340 15695 12570 15780
rect 12690 15695 12920 15780
rect 13040 15695 13270 15780
rect 13390 15695 13620 15780
rect 13740 15695 13970 15780
rect 14090 15695 14320 15780
rect 14440 15695 14670 15780
rect 9540 15645 14670 15695
rect 9540 15550 9770 15645
rect 9890 15550 10120 15645
rect 10240 15550 10470 15645
rect 10590 15550 10820 15645
rect 10940 15550 11170 15645
rect 11290 15550 11520 15645
rect 11640 15550 11870 15645
rect 11990 15550 12220 15645
rect 12340 15550 12570 15645
rect 12690 15550 12920 15645
rect 13040 15550 13270 15645
rect 13390 15550 13620 15645
rect 13740 15550 13970 15645
rect 14090 15550 14320 15645
rect 14440 15550 14670 15645
rect 230 15430 280 15550
rect 12080 15430 12130 15550
rect -1260 15345 -1030 15430
rect -910 15345 -680 15430
rect -560 15345 -330 15430
rect -210 15345 20 15430
rect 140 15345 370 15430
rect 490 15345 720 15430
rect 840 15345 1070 15430
rect 1190 15345 1420 15430
rect 1540 15345 1770 15430
rect -1260 15295 1770 15345
rect -1260 15200 -1030 15295
rect -910 15200 -680 15295
rect -560 15200 -330 15295
rect -210 15200 20 15295
rect 140 15200 370 15295
rect 490 15200 720 15295
rect 840 15200 1070 15295
rect 1190 15200 1420 15295
rect 1540 15200 1770 15295
rect 9540 15345 9770 15430
rect 9890 15345 10120 15430
rect 10240 15345 10470 15430
rect 10590 15345 10820 15430
rect 10940 15345 11170 15430
rect 11290 15345 11520 15430
rect 11640 15345 11870 15430
rect 11990 15345 12220 15430
rect 12340 15345 12570 15430
rect 12690 15345 12920 15430
rect 13040 15345 13270 15430
rect 13390 15345 13620 15430
rect 13740 15345 13970 15430
rect 14090 15345 14320 15430
rect 14440 15345 14670 15430
rect 9540 15295 14670 15345
rect 9540 15200 9770 15295
rect 9890 15200 10120 15295
rect 10240 15200 10470 15295
rect 10590 15200 10820 15295
rect 10940 15200 11170 15295
rect 11290 15200 11520 15295
rect 11640 15200 11870 15295
rect 11990 15200 12220 15295
rect 12340 15200 12570 15295
rect 12690 15200 12920 15295
rect 13040 15200 13270 15295
rect 13390 15200 13620 15295
rect 13740 15200 13970 15295
rect 14090 15200 14320 15295
rect 14440 15200 14670 15295
rect 230 15080 280 15200
rect 12080 15080 12130 15200
rect -1260 14995 -1030 15080
rect -910 14995 -680 15080
rect -560 14995 -330 15080
rect -210 14995 20 15080
rect 140 14995 370 15080
rect 490 14995 720 15080
rect 840 14995 1070 15080
rect 1190 14995 1420 15080
rect 1540 14995 1770 15080
rect -1260 14945 1770 14995
rect -1260 14850 -1030 14945
rect -910 14850 -680 14945
rect -560 14850 -330 14945
rect -210 14850 20 14945
rect 140 14850 370 14945
rect 490 14850 720 14945
rect 840 14850 1070 14945
rect 1190 14850 1420 14945
rect 1540 14850 1770 14945
rect 9540 14995 9770 15080
rect 9890 14995 10120 15080
rect 10240 14995 10470 15080
rect 10590 14995 10820 15080
rect 10940 14995 11170 15080
rect 11290 14995 11520 15080
rect 11640 14995 11870 15080
rect 11990 14995 12220 15080
rect 12340 14995 12570 15080
rect 12690 14995 12920 15080
rect 13040 14995 13270 15080
rect 13390 14995 13620 15080
rect 13740 14995 13970 15080
rect 14090 14995 14320 15080
rect 14440 14995 14670 15080
rect 9540 14945 14670 14995
rect 9540 14850 9770 14945
rect 9890 14850 10120 14945
rect 10240 14850 10470 14945
rect 10590 14850 10820 14945
rect 10940 14850 11170 14945
rect 11290 14850 11520 14945
rect 11640 14850 11870 14945
rect 11990 14850 12220 14945
rect 12340 14850 12570 14945
rect 12690 14850 12920 14945
rect 13040 14850 13270 14945
rect 13390 14850 13620 14945
rect 13740 14850 13970 14945
rect 14090 14850 14320 14945
rect 14440 14850 14670 14945
rect 230 14730 280 14850
rect 12080 14730 12130 14850
rect -1260 14645 -1030 14730
rect -910 14645 -680 14730
rect -560 14645 -330 14730
rect -210 14645 20 14730
rect 140 14645 370 14730
rect 490 14645 720 14730
rect 840 14645 1070 14730
rect 1190 14645 1420 14730
rect 1540 14645 1770 14730
rect -1260 14595 1770 14645
rect -1260 14500 -1030 14595
rect -910 14500 -680 14595
rect -560 14500 -330 14595
rect -210 14500 20 14595
rect 140 14500 370 14595
rect 490 14500 720 14595
rect 840 14500 1070 14595
rect 1190 14500 1420 14595
rect 1540 14500 1770 14595
rect 9540 14645 9770 14730
rect 9890 14645 10120 14730
rect 10240 14645 10470 14730
rect 10590 14645 10820 14730
rect 10940 14645 11170 14730
rect 11290 14645 11520 14730
rect 11640 14645 11870 14730
rect 11990 14645 12220 14730
rect 12340 14645 12570 14730
rect 12690 14645 12920 14730
rect 13040 14645 13270 14730
rect 13390 14645 13620 14730
rect 13740 14645 13970 14730
rect 14090 14645 14320 14730
rect 14440 14645 14670 14730
rect 9540 14595 14670 14645
rect 9540 14500 9770 14595
rect 9890 14500 10120 14595
rect 10240 14500 10470 14595
rect 10590 14500 10820 14595
rect 10940 14500 11170 14595
rect 11290 14500 11520 14595
rect 11640 14500 11870 14595
rect 11990 14500 12220 14595
rect 12340 14500 12570 14595
rect 12690 14500 12920 14595
rect 13040 14500 13270 14595
rect 13390 14500 13620 14595
rect 13740 14500 13970 14595
rect 14090 14500 14320 14595
rect 14440 14500 14670 14595
rect 230 14380 280 14500
rect 12080 14380 12130 14500
rect -1260 14295 -1030 14380
rect -910 14295 -680 14380
rect -560 14295 -330 14380
rect -210 14295 20 14380
rect 140 14295 370 14380
rect 490 14295 720 14380
rect 840 14295 1070 14380
rect 1190 14295 1420 14380
rect 1540 14295 1770 14380
rect -1260 14245 1770 14295
rect -1260 14150 -1030 14245
rect -910 14150 -680 14245
rect -560 14150 -330 14245
rect -210 14150 20 14245
rect 140 14150 370 14245
rect 490 14150 720 14245
rect 840 14150 1070 14245
rect 1190 14150 1420 14245
rect 1540 14150 1770 14245
rect 9540 14295 9770 14380
rect 9890 14295 10120 14380
rect 10240 14295 10470 14380
rect 10590 14295 10820 14380
rect 10940 14295 11170 14380
rect 11290 14295 11520 14380
rect 11640 14295 11870 14380
rect 11990 14295 12220 14380
rect 12340 14295 12570 14380
rect 12690 14295 12920 14380
rect 13040 14295 13270 14380
rect 13390 14295 13620 14380
rect 13740 14295 13970 14380
rect 14090 14295 14320 14380
rect 14440 14295 14670 14380
rect 9540 14245 14670 14295
rect 9540 14150 9770 14245
rect 9890 14150 10120 14245
rect 10240 14150 10470 14245
rect 10590 14150 10820 14245
rect 10940 14150 11170 14245
rect 11290 14150 11520 14245
rect 11640 14150 11870 14245
rect 11990 14150 12220 14245
rect 12340 14150 12570 14245
rect 12690 14150 12920 14245
rect 13040 14150 13270 14245
rect 13390 14150 13620 14245
rect 13740 14150 13970 14245
rect 14090 14150 14320 14245
rect 14440 14150 14670 14245
rect 230 14030 280 14150
rect 12080 14030 12130 14150
rect -1260 13945 -1030 14030
rect -910 13945 -680 14030
rect -560 13945 -330 14030
rect -210 13945 20 14030
rect 140 13945 370 14030
rect 490 13945 720 14030
rect 840 13945 1070 14030
rect 1190 13945 1420 14030
rect 1540 13945 1770 14030
rect -1260 13895 1770 13945
rect -1260 13800 -1030 13895
rect -910 13800 -680 13895
rect -560 13800 -330 13895
rect -210 13800 20 13895
rect 140 13800 370 13895
rect 490 13800 720 13895
rect 840 13800 1070 13895
rect 1190 13800 1420 13895
rect 1540 13800 1770 13895
rect 9540 13945 9770 14030
rect 9890 13945 10120 14030
rect 10240 13945 10470 14030
rect 10590 13945 10820 14030
rect 10940 13945 11170 14030
rect 11290 13945 11520 14030
rect 11640 13945 11870 14030
rect 11990 13945 12220 14030
rect 12340 13945 12570 14030
rect 12690 13945 12920 14030
rect 13040 13945 13270 14030
rect 13390 13945 13620 14030
rect 13740 13945 13970 14030
rect 14090 13945 14320 14030
rect 14440 13945 14670 14030
rect 9540 13895 14670 13945
rect 9540 13800 9770 13895
rect 9890 13800 10120 13895
rect 10240 13800 10470 13895
rect 10590 13800 10820 13895
rect 10940 13800 11170 13895
rect 11290 13800 11520 13895
rect 11640 13800 11870 13895
rect 11990 13800 12220 13895
rect 12340 13800 12570 13895
rect 12690 13800 12920 13895
rect 13040 13800 13270 13895
rect 13390 13800 13620 13895
rect 13740 13800 13970 13895
rect 14090 13800 14320 13895
rect 14440 13800 14670 13895
rect 230 13680 280 13800
rect 12080 13680 12130 13800
rect -1260 13595 -1030 13680
rect -910 13595 -680 13680
rect -560 13595 -330 13680
rect -210 13595 20 13680
rect 140 13595 370 13680
rect 490 13595 720 13680
rect 840 13595 1070 13680
rect 1190 13595 1420 13680
rect 1540 13595 1770 13680
rect -1260 13545 1770 13595
rect -1260 13450 -1030 13545
rect -910 13450 -680 13545
rect -560 13450 -330 13545
rect -210 13450 20 13545
rect 140 13450 370 13545
rect 490 13450 720 13545
rect 840 13450 1070 13545
rect 1190 13450 1420 13545
rect 1540 13450 1770 13545
rect 9540 13595 9770 13680
rect 9890 13595 10120 13680
rect 10240 13595 10470 13680
rect 10590 13595 10820 13680
rect 10940 13595 11170 13680
rect 11290 13595 11520 13680
rect 11640 13595 11870 13680
rect 11990 13595 12220 13680
rect 12340 13595 12570 13680
rect 12690 13595 12920 13680
rect 13040 13595 13270 13680
rect 13390 13595 13620 13680
rect 13740 13595 13970 13680
rect 14090 13595 14320 13680
rect 14440 13595 14670 13680
rect 9540 13545 14670 13595
rect 9540 13450 9770 13545
rect 9890 13450 10120 13545
rect 10240 13450 10470 13545
rect 10590 13450 10820 13545
rect 10940 13450 11170 13545
rect 11290 13450 11520 13545
rect 11640 13450 11870 13545
rect 11990 13450 12220 13545
rect 12340 13450 12570 13545
rect 12690 13450 12920 13545
rect 13040 13450 13270 13545
rect 13390 13450 13620 13545
rect 13740 13450 13970 13545
rect 14090 13450 14320 13545
rect 14440 13450 14670 13545
rect 230 13330 280 13450
rect 12080 13330 12130 13450
rect -1260 13245 -1030 13330
rect -910 13245 -680 13330
rect -560 13245 -330 13330
rect -210 13245 20 13330
rect 140 13245 370 13330
rect 490 13245 720 13330
rect 840 13245 1070 13330
rect 1190 13245 1420 13330
rect 1540 13245 1770 13330
rect -1260 13195 1770 13245
rect -1260 13100 -1030 13195
rect -910 13100 -680 13195
rect -560 13100 -330 13195
rect -210 13100 20 13195
rect 140 13100 370 13195
rect 490 13100 720 13195
rect 840 13100 1070 13195
rect 1190 13100 1420 13195
rect 1540 13100 1770 13195
rect 9540 13245 9770 13330
rect 9890 13245 10120 13330
rect 10240 13245 10470 13330
rect 10590 13245 10820 13330
rect 10940 13245 11170 13330
rect 11290 13245 11520 13330
rect 11640 13245 11870 13330
rect 11990 13245 12220 13330
rect 12340 13245 12570 13330
rect 12690 13245 12920 13330
rect 13040 13245 13270 13330
rect 13390 13245 13620 13330
rect 13740 13245 13970 13330
rect 14090 13245 14320 13330
rect 14440 13245 14670 13330
rect 9540 13195 14670 13245
rect 9540 13100 9770 13195
rect 9890 13100 10120 13195
rect 10240 13100 10470 13195
rect 10590 13100 10820 13195
rect 10940 13100 11170 13195
rect 11290 13100 11520 13195
rect 11640 13100 11870 13195
rect 11990 13100 12220 13195
rect 12340 13100 12570 13195
rect 12690 13100 12920 13195
rect 13040 13100 13270 13195
rect 13390 13100 13620 13195
rect 13740 13100 13970 13195
rect 14090 13100 14320 13195
rect 14440 13100 14670 13195
rect 230 12980 280 13100
rect 12080 12980 12130 13100
rect -1260 12895 -1030 12980
rect -910 12895 -680 12980
rect -560 12895 -330 12980
rect -210 12895 20 12980
rect 140 12895 370 12980
rect 490 12895 720 12980
rect 840 12895 1070 12980
rect 1190 12895 1420 12980
rect 1540 12895 1770 12980
rect -1260 12845 1770 12895
rect -1260 12750 -1030 12845
rect -910 12750 -680 12845
rect -560 12750 -330 12845
rect -210 12750 20 12845
rect 140 12750 370 12845
rect 490 12750 720 12845
rect 840 12750 1070 12845
rect 1190 12750 1420 12845
rect 1540 12750 1770 12845
rect 9540 12895 9770 12980
rect 9890 12895 10120 12980
rect 10240 12895 10470 12980
rect 10590 12895 10820 12980
rect 10940 12895 11170 12980
rect 11290 12895 11520 12980
rect 11640 12895 11870 12980
rect 11990 12895 12220 12980
rect 12340 12895 12570 12980
rect 12690 12895 12920 12980
rect 13040 12895 13270 12980
rect 13390 12895 13620 12980
rect 13740 12895 13970 12980
rect 14090 12895 14320 12980
rect 14440 12895 14670 12980
rect 9540 12845 14670 12895
rect 9540 12750 9770 12845
rect 9890 12750 10120 12845
rect 10240 12750 10470 12845
rect 10590 12750 10820 12845
rect 10940 12750 11170 12845
rect 11290 12750 11520 12845
rect 11640 12750 11870 12845
rect 11990 12750 12220 12845
rect 12340 12750 12570 12845
rect 12690 12750 12920 12845
rect 13040 12750 13270 12845
rect 13390 12750 13620 12845
rect 13740 12750 13970 12845
rect 14090 12750 14320 12845
rect 14440 12750 14670 12845
rect 230 12630 280 12750
rect 12080 12630 12130 12750
rect -1260 12545 -1030 12630
rect -910 12545 -680 12630
rect -560 12545 -330 12630
rect -210 12545 20 12630
rect 140 12545 370 12630
rect 490 12545 720 12630
rect 840 12545 1070 12630
rect 1190 12545 1420 12630
rect 1540 12545 1770 12630
rect -1260 12495 1770 12545
rect -1260 12400 -1030 12495
rect -910 12400 -680 12495
rect -560 12400 -330 12495
rect -210 12400 20 12495
rect 140 12400 370 12495
rect 490 12400 720 12495
rect 840 12400 1070 12495
rect 1190 12400 1420 12495
rect 1540 12400 1770 12495
rect 9540 12545 9770 12630
rect 9890 12545 10120 12630
rect 10240 12545 10470 12630
rect 10590 12545 10820 12630
rect 10940 12545 11170 12630
rect 11290 12545 11520 12630
rect 11640 12545 11870 12630
rect 11990 12545 12220 12630
rect 12340 12545 12570 12630
rect 12690 12545 12920 12630
rect 13040 12545 13270 12630
rect 13390 12545 13620 12630
rect 13740 12545 13970 12630
rect 14090 12545 14320 12630
rect 14440 12545 14670 12630
rect 9540 12495 14670 12545
rect 9540 12400 9770 12495
rect 9890 12400 10120 12495
rect 10240 12400 10470 12495
rect 10590 12400 10820 12495
rect 10940 12400 11170 12495
rect 11290 12400 11520 12495
rect 11640 12400 11870 12495
rect 11990 12400 12220 12495
rect 12340 12400 12570 12495
rect 12690 12400 12920 12495
rect 13040 12400 13270 12495
rect 13390 12400 13620 12495
rect 13740 12400 13970 12495
rect 14090 12400 14320 12495
rect 14440 12400 14670 12495
rect 230 12280 280 12400
rect 12080 12280 12130 12400
rect -1260 12195 -1030 12280
rect -910 12195 -680 12280
rect -560 12195 -330 12280
rect -210 12195 20 12280
rect 140 12195 370 12280
rect 490 12195 720 12280
rect 840 12195 1070 12280
rect 1190 12195 1420 12280
rect 1540 12195 1770 12280
rect -1260 12145 1770 12195
rect -1260 12050 -1030 12145
rect -910 12050 -680 12145
rect -560 12050 -330 12145
rect -210 12050 20 12145
rect 140 12050 370 12145
rect 490 12050 720 12145
rect 840 12050 1070 12145
rect 1190 12050 1420 12145
rect 1540 12050 1770 12145
rect 9540 12195 9770 12280
rect 9890 12195 10120 12280
rect 10240 12195 10470 12280
rect 10590 12195 10820 12280
rect 10940 12195 11170 12280
rect 11290 12195 11520 12280
rect 11640 12195 11870 12280
rect 11990 12195 12220 12280
rect 12340 12195 12570 12280
rect 12690 12195 12920 12280
rect 13040 12195 13270 12280
rect 13390 12195 13620 12280
rect 13740 12195 13970 12280
rect 14090 12195 14320 12280
rect 14440 12195 14670 12280
rect 9540 12145 14670 12195
rect 9540 12050 9770 12145
rect 9890 12050 10120 12145
rect 10240 12050 10470 12145
rect 10590 12050 10820 12145
rect 10940 12050 11170 12145
rect 11290 12050 11520 12145
rect 11640 12050 11870 12145
rect 11990 12050 12220 12145
rect 12340 12050 12570 12145
rect 12690 12050 12920 12145
rect 13040 12050 13270 12145
rect 13390 12050 13620 12145
rect 13740 12050 13970 12145
rect 14090 12050 14320 12145
rect 14440 12050 14670 12145
rect 230 11930 280 12050
rect 12080 11930 12130 12050
rect -1260 11845 -1030 11930
rect -910 11845 -680 11930
rect -560 11845 -330 11930
rect -210 11845 20 11930
rect 140 11845 370 11930
rect 490 11845 720 11930
rect 840 11845 1070 11930
rect 1190 11845 1420 11930
rect 1540 11845 1770 11930
rect -1260 11795 1770 11845
rect -1260 11700 -1030 11795
rect -910 11700 -680 11795
rect -560 11700 -330 11795
rect -210 11700 20 11795
rect 140 11700 370 11795
rect 490 11700 720 11795
rect 840 11700 1070 11795
rect 1190 11700 1420 11795
rect 1540 11700 1770 11795
rect 9540 11845 9770 11930
rect 9890 11845 10120 11930
rect 10240 11845 10470 11930
rect 10590 11845 10820 11930
rect 10940 11845 11170 11930
rect 11290 11845 11520 11930
rect 11640 11845 11870 11930
rect 11990 11845 12220 11930
rect 12340 11845 12570 11930
rect 12690 11845 12920 11930
rect 13040 11845 13270 11930
rect 13390 11845 13620 11930
rect 13740 11845 13970 11930
rect 14090 11845 14320 11930
rect 14440 11845 14670 11930
rect 9540 11795 14670 11845
rect 9540 11700 9770 11795
rect 9890 11700 10120 11795
rect 10240 11700 10470 11795
rect 10590 11700 10820 11795
rect 10940 11700 11170 11795
rect 11290 11700 11520 11795
rect 11640 11700 11870 11795
rect 11990 11700 12220 11795
rect 12340 11700 12570 11795
rect 12690 11700 12920 11795
rect 13040 11700 13270 11795
rect 13390 11700 13620 11795
rect 13740 11700 13970 11795
rect 14090 11700 14320 11795
rect 14440 11700 14670 11795
rect 230 11580 280 11700
rect 12080 11580 12130 11700
rect -1260 11495 -1030 11580
rect -910 11495 -680 11580
rect -560 11495 -330 11580
rect -210 11495 20 11580
rect 140 11495 370 11580
rect 490 11495 720 11580
rect 840 11495 1070 11580
rect 1190 11495 1420 11580
rect 1540 11495 1770 11580
rect -1260 11445 1770 11495
rect -1260 11350 -1030 11445
rect -910 11350 -680 11445
rect -560 11350 -330 11445
rect -210 11350 20 11445
rect 140 11350 370 11445
rect 490 11350 720 11445
rect 840 11350 1070 11445
rect 1190 11350 1420 11445
rect 1540 11350 1770 11445
rect 9540 11495 9770 11580
rect 9890 11495 10120 11580
rect 10240 11495 10470 11580
rect 10590 11495 10820 11580
rect 10940 11495 11170 11580
rect 11290 11495 11520 11580
rect 11640 11495 11870 11580
rect 11990 11495 12220 11580
rect 12340 11495 12570 11580
rect 12690 11495 12920 11580
rect 13040 11495 13270 11580
rect 13390 11495 13620 11580
rect 13740 11495 13970 11580
rect 14090 11495 14320 11580
rect 14440 11495 14670 11580
rect 9540 11445 14670 11495
rect 9540 11350 9770 11445
rect 9890 11350 10120 11445
rect 10240 11350 10470 11445
rect 10590 11350 10820 11445
rect 10940 11350 11170 11445
rect 11290 11350 11520 11445
rect 11640 11350 11870 11445
rect 11990 11350 12220 11445
rect 12340 11350 12570 11445
rect 12690 11350 12920 11445
rect 13040 11350 13270 11445
rect 13390 11350 13620 11445
rect 13740 11350 13970 11445
rect 14090 11350 14320 11445
rect 14440 11350 14670 11445
rect 230 11230 280 11350
rect 12080 11230 12130 11350
rect -1260 11145 -1030 11230
rect -910 11145 -680 11230
rect -560 11145 -330 11230
rect -210 11145 20 11230
rect 140 11145 370 11230
rect 490 11145 720 11230
rect 840 11145 1070 11230
rect 1190 11145 1420 11230
rect 1540 11145 1770 11230
rect -1260 11095 1770 11145
rect -1260 11000 -1030 11095
rect -910 11000 -680 11095
rect -560 11000 -330 11095
rect -210 11000 20 11095
rect 140 11000 370 11095
rect 490 11000 720 11095
rect 840 11000 1070 11095
rect 1190 11000 1420 11095
rect 1540 11000 1770 11095
rect 9540 11145 9770 11230
rect 9890 11145 10120 11230
rect 10240 11145 10470 11230
rect 10590 11145 10820 11230
rect 10940 11145 11170 11230
rect 11290 11145 11520 11230
rect 11640 11145 11870 11230
rect 11990 11145 12220 11230
rect 12340 11145 12570 11230
rect 12690 11145 12920 11230
rect 13040 11145 13270 11230
rect 13390 11145 13620 11230
rect 13740 11145 13970 11230
rect 14090 11145 14320 11230
rect 14440 11145 14670 11230
rect 9540 11095 14670 11145
rect 9540 11000 9770 11095
rect 9890 11000 10120 11095
rect 10240 11000 10470 11095
rect 10590 11000 10820 11095
rect 10940 11000 11170 11095
rect 11290 11000 11520 11095
rect 11640 11000 11870 11095
rect 11990 11000 12220 11095
rect 12340 11000 12570 11095
rect 12690 11000 12920 11095
rect 13040 11000 13270 11095
rect 13390 11000 13620 11095
rect 13740 11000 13970 11095
rect 14090 11000 14320 11095
rect 14440 11000 14670 11095
rect 230 10880 280 11000
rect 12080 10880 12130 11000
rect -1260 10795 -1030 10880
rect -910 10795 -680 10880
rect -560 10795 -330 10880
rect -210 10795 20 10880
rect 140 10795 370 10880
rect 490 10795 720 10880
rect 840 10795 1070 10880
rect 1190 10795 1420 10880
rect 1540 10795 1770 10880
rect -1260 10745 1770 10795
rect -1260 10650 -1030 10745
rect -910 10650 -680 10745
rect -560 10650 -330 10745
rect -210 10650 20 10745
rect 140 10650 370 10745
rect 490 10650 720 10745
rect 840 10650 1070 10745
rect 1190 10650 1420 10745
rect 1540 10650 1770 10745
rect 9540 10795 9770 10880
rect 9890 10795 10120 10880
rect 10240 10795 10470 10880
rect 10590 10795 10820 10880
rect 10940 10795 11170 10880
rect 11290 10795 11520 10880
rect 11640 10795 11870 10880
rect 11990 10795 12220 10880
rect 12340 10795 12570 10880
rect 12690 10795 12920 10880
rect 13040 10795 13270 10880
rect 13390 10795 13620 10880
rect 13740 10795 13970 10880
rect 14090 10795 14320 10880
rect 14440 10795 14670 10880
rect 9540 10745 14670 10795
rect 9540 10650 9770 10745
rect 9890 10650 10120 10745
rect 10240 10650 10470 10745
rect 10590 10650 10820 10745
rect 10940 10650 11170 10745
rect 11290 10650 11520 10745
rect 11640 10650 11870 10745
rect 11990 10650 12220 10745
rect 12340 10650 12570 10745
rect 12690 10650 12920 10745
rect 13040 10650 13270 10745
rect 13390 10650 13620 10745
rect 13740 10650 13970 10745
rect 14090 10650 14320 10745
rect 14440 10650 14670 10745
rect 230 10530 280 10650
rect 12080 10530 12130 10650
rect -1260 10445 -1030 10530
rect -910 10445 -680 10530
rect -560 10445 -330 10530
rect -210 10445 20 10530
rect 140 10445 370 10530
rect 490 10445 720 10530
rect 840 10445 1070 10530
rect 1190 10445 1420 10530
rect 1540 10445 1770 10530
rect -1260 10395 1770 10445
rect -1260 10300 -1030 10395
rect -910 10300 -680 10395
rect -560 10300 -330 10395
rect -210 10300 20 10395
rect 140 10300 370 10395
rect 490 10300 720 10395
rect 840 10300 1070 10395
rect 1190 10300 1420 10395
rect 1540 10300 1770 10395
rect 9540 10445 9770 10530
rect 9890 10445 10120 10530
rect 10240 10445 10470 10530
rect 10590 10445 10820 10530
rect 10940 10445 11170 10530
rect 11290 10445 11520 10530
rect 11640 10445 11870 10530
rect 11990 10445 12220 10530
rect 12340 10445 12570 10530
rect 12690 10445 12920 10530
rect 13040 10445 13270 10530
rect 13390 10445 13620 10530
rect 13740 10445 13970 10530
rect 14090 10445 14320 10530
rect 14440 10445 14670 10530
rect 9540 10395 14670 10445
rect 9540 10300 9770 10395
rect 9890 10300 10120 10395
rect 10240 10300 10470 10395
rect 10590 10300 10820 10395
rect 10940 10300 11170 10395
rect 11290 10300 11520 10395
rect 11640 10300 11870 10395
rect 11990 10300 12220 10395
rect 12340 10300 12570 10395
rect 12690 10300 12920 10395
rect 13040 10300 13270 10395
rect 13390 10300 13620 10395
rect 13740 10300 13970 10395
rect 14090 10300 14320 10395
rect 14440 10300 14670 10395
rect 230 10180 280 10300
rect 12080 10180 12130 10300
rect -4840 9615 -1640 10155
rect -1260 10095 -1030 10180
rect -910 10095 -680 10180
rect -560 10095 -330 10180
rect -210 10095 20 10180
rect 140 10095 370 10180
rect 490 10095 720 10180
rect 840 10095 1070 10180
rect 1190 10095 1420 10180
rect 1540 10095 1770 10180
rect -1260 10090 1770 10095
rect 9540 10095 9770 10180
rect 9890 10095 10120 10180
rect 10240 10095 10470 10180
rect 10590 10095 10820 10180
rect 10940 10095 11170 10180
rect 11290 10095 11520 10180
rect 11640 10095 11870 10180
rect 11990 10095 12220 10180
rect 12340 10095 12570 10180
rect 12690 10095 12920 10180
rect 13040 10095 13270 10180
rect 13390 10095 13620 10180
rect 13740 10095 13970 10180
rect 14090 10095 14320 10180
rect 14440 10095 14670 10180
rect -1260 10085 2095 10090
rect -1260 10055 2060 10085
rect 2090 10055 2095 10085
rect -1260 10050 2095 10055
rect -1260 10045 1770 10050
rect -1260 9950 -1030 10045
rect -910 9950 -680 10045
rect -560 9950 -330 10045
rect -210 9950 20 10045
rect 140 9950 370 10045
rect 490 9950 720 10045
rect 840 9950 1070 10045
rect 1190 9950 1420 10045
rect 1540 9950 1770 10045
rect 9540 10045 14670 10095
rect 9540 9950 9770 10045
rect 9890 9950 10120 10045
rect 10240 9950 10470 10045
rect 10590 9950 10820 10045
rect 10940 9950 11170 10045
rect 11290 9950 11520 10045
rect 11640 9950 11870 10045
rect 11990 9950 12220 10045
rect 12340 9950 12570 10045
rect 12690 9950 12920 10045
rect 13040 9950 13270 10045
rect 13390 9950 13620 10045
rect 13740 9950 13970 10045
rect 14090 9950 14320 10045
rect 14440 9950 14670 10045
rect 12080 9830 12130 9950
rect 9540 9745 9770 9830
rect 9890 9745 10120 9830
rect 10240 9745 10470 9830
rect 10590 9745 10820 9830
rect 10940 9745 11170 9830
rect 11290 9745 11520 9830
rect 11640 9745 11870 9830
rect 11990 9745 12220 9830
rect 12340 9745 12570 9830
rect 12690 9745 12920 9830
rect 13040 9745 13270 9830
rect 13390 9745 13620 9830
rect 13740 9745 13970 9830
rect 14090 9745 14320 9830
rect 14440 9745 14670 9830
rect 9540 9695 14670 9745
rect -4840 9565 -4805 9615
rect -4755 9565 -4710 9615
rect -4660 9565 -4615 9615
rect -4565 9565 -4515 9615
rect -4465 9565 -4415 9615
rect -4365 9565 -4315 9615
rect -4265 9565 -4220 9615
rect -4170 9565 -4125 9615
rect -4075 9565 -4005 9615
rect -3955 9565 -3910 9615
rect -3860 9565 -3815 9615
rect -3765 9565 -3715 9615
rect -3665 9565 -3615 9615
rect -3565 9565 -3515 9615
rect -3465 9565 -3420 9615
rect -3370 9565 -3325 9615
rect -3275 9565 -3205 9615
rect -3155 9565 -3110 9615
rect -3060 9565 -3015 9615
rect -2965 9565 -2915 9615
rect -2865 9565 -2815 9615
rect -2765 9565 -2715 9615
rect -2665 9565 -2620 9615
rect -2570 9565 -2525 9615
rect -2475 9565 -2405 9615
rect -2355 9565 -2310 9615
rect -2260 9565 -2215 9615
rect -2165 9565 -2115 9615
rect -2065 9565 -2015 9615
rect -1965 9565 -1915 9615
rect -1865 9565 -1820 9615
rect -1770 9565 -1725 9615
rect -1675 9565 -1640 9615
rect -4840 9525 -1640 9565
rect -4840 9475 -4805 9525
rect -4755 9475 -4710 9525
rect -4660 9475 -4615 9525
rect -4565 9475 -4515 9525
rect -4465 9475 -4415 9525
rect -4365 9475 -4315 9525
rect -4265 9475 -4220 9525
rect -4170 9475 -4125 9525
rect -4075 9475 -4005 9525
rect -3955 9475 -3910 9525
rect -3860 9475 -3815 9525
rect -3765 9475 -3715 9525
rect -3665 9475 -3615 9525
rect -3565 9475 -3515 9525
rect -3465 9475 -3420 9525
rect -3370 9475 -3325 9525
rect -3275 9475 -3205 9525
rect -3155 9475 -3110 9525
rect -3060 9475 -3015 9525
rect -2965 9475 -2915 9525
rect -2865 9475 -2815 9525
rect -2765 9475 -2715 9525
rect -2665 9475 -2620 9525
rect -2570 9475 -2525 9525
rect -2475 9475 -2405 9525
rect -2355 9475 -2310 9525
rect -2260 9475 -2215 9525
rect -2165 9475 -2115 9525
rect -2065 9475 -2015 9525
rect -1965 9475 -1915 9525
rect -1865 9475 -1820 9525
rect -1770 9475 -1725 9525
rect -1675 9475 -1640 9525
rect -4840 9425 -1640 9475
rect -4840 9375 -4805 9425
rect -4755 9375 -4710 9425
rect -4660 9375 -4615 9425
rect -4565 9375 -4515 9425
rect -4465 9375 -4415 9425
rect -4365 9375 -4315 9425
rect -4265 9375 -4220 9425
rect -4170 9375 -4125 9425
rect -4075 9375 -4005 9425
rect -3955 9375 -3910 9425
rect -3860 9375 -3815 9425
rect -3765 9375 -3715 9425
rect -3665 9375 -3615 9425
rect -3565 9375 -3515 9425
rect -3465 9375 -3420 9425
rect -3370 9375 -3325 9425
rect -3275 9375 -3205 9425
rect -3155 9375 -3110 9425
rect -3060 9375 -3015 9425
rect -2965 9375 -2915 9425
rect -2865 9375 -2815 9425
rect -2765 9375 -2715 9425
rect -2665 9375 -2620 9425
rect -2570 9375 -2525 9425
rect -2475 9375 -2405 9425
rect -2355 9375 -2310 9425
rect -2260 9375 -2215 9425
rect -2165 9375 -2115 9425
rect -2065 9375 -2015 9425
rect -1965 9375 -1915 9425
rect -1865 9375 -1820 9425
rect -1770 9375 -1725 9425
rect -1675 9375 -1640 9425
rect -4840 9335 -1640 9375
rect -4840 9285 -4805 9335
rect -4755 9285 -4710 9335
rect -4660 9285 -4615 9335
rect -4565 9285 -4515 9335
rect -4465 9285 -4415 9335
rect -4365 9285 -4315 9335
rect -4265 9285 -4220 9335
rect -4170 9285 -4125 9335
rect -4075 9285 -4005 9335
rect -3955 9285 -3910 9335
rect -3860 9285 -3815 9335
rect -3765 9285 -3715 9335
rect -3665 9285 -3615 9335
rect -3565 9285 -3515 9335
rect -3465 9285 -3420 9335
rect -3370 9285 -3325 9335
rect -3275 9285 -3205 9335
rect -3155 9285 -3110 9335
rect -3060 9285 -3015 9335
rect -2965 9285 -2915 9335
rect -2865 9285 -2815 9335
rect -2765 9285 -2715 9335
rect -2665 9285 -2620 9335
rect -2570 9285 -2525 9335
rect -2475 9285 -2405 9335
rect -2355 9285 -2310 9335
rect -2260 9285 -2215 9335
rect -2165 9285 -2115 9335
rect -2065 9285 -2015 9335
rect -1965 9285 -1915 9335
rect -1865 9285 -1820 9335
rect -1770 9285 -1725 9335
rect -1675 9285 -1640 9335
rect -4840 9215 -1640 9285
rect -4840 9165 -4805 9215
rect -4755 9165 -4710 9215
rect -4660 9165 -4615 9215
rect -4565 9165 -4515 9215
rect -4465 9165 -4415 9215
rect -4365 9165 -4315 9215
rect -4265 9165 -4220 9215
rect -4170 9165 -4125 9215
rect -4075 9165 -4005 9215
rect -3955 9165 -3910 9215
rect -3860 9165 -3815 9215
rect -3765 9165 -3715 9215
rect -3665 9165 -3615 9215
rect -3565 9165 -3515 9215
rect -3465 9165 -3420 9215
rect -3370 9165 -3325 9215
rect -3275 9165 -3205 9215
rect -3155 9165 -3110 9215
rect -3060 9165 -3015 9215
rect -2965 9165 -2915 9215
rect -2865 9165 -2815 9215
rect -2765 9165 -2715 9215
rect -2665 9165 -2620 9215
rect -2570 9165 -2525 9215
rect -2475 9165 -2405 9215
rect -2355 9165 -2310 9215
rect -2260 9165 -2215 9215
rect -2165 9165 -2115 9215
rect -2065 9165 -2015 9215
rect -1965 9165 -1915 9215
rect -1865 9165 -1820 9215
rect -1770 9165 -1725 9215
rect -1675 9165 -1640 9215
rect -4840 9125 -1640 9165
rect -4840 9075 -4805 9125
rect -4755 9075 -4710 9125
rect -4660 9075 -4615 9125
rect -4565 9075 -4515 9125
rect -4465 9075 -4415 9125
rect -4365 9075 -4315 9125
rect -4265 9075 -4220 9125
rect -4170 9075 -4125 9125
rect -4075 9075 -4005 9125
rect -3955 9075 -3910 9125
rect -3860 9075 -3815 9125
rect -3765 9075 -3715 9125
rect -3665 9075 -3615 9125
rect -3565 9075 -3515 9125
rect -3465 9075 -3420 9125
rect -3370 9075 -3325 9125
rect -3275 9075 -3205 9125
rect -3155 9075 -3110 9125
rect -3060 9075 -3015 9125
rect -2965 9075 -2915 9125
rect -2865 9075 -2815 9125
rect -2765 9075 -2715 9125
rect -2665 9075 -2620 9125
rect -2570 9075 -2525 9125
rect -2475 9075 -2405 9125
rect -2355 9075 -2310 9125
rect -2260 9075 -2215 9125
rect -2165 9075 -2115 9125
rect -2065 9075 -2015 9125
rect -1965 9075 -1915 9125
rect -1865 9075 -1820 9125
rect -1770 9075 -1725 9125
rect -1675 9075 -1640 9125
rect -4840 9025 -1640 9075
rect -4840 8975 -4805 9025
rect -4755 8975 -4710 9025
rect -4660 8975 -4615 9025
rect -4565 8975 -4515 9025
rect -4465 8975 -4415 9025
rect -4365 8975 -4315 9025
rect -4265 8975 -4220 9025
rect -4170 8975 -4125 9025
rect -4075 8975 -4005 9025
rect -3955 8975 -3910 9025
rect -3860 8975 -3815 9025
rect -3765 8975 -3715 9025
rect -3665 8975 -3615 9025
rect -3565 8975 -3515 9025
rect -3465 8975 -3420 9025
rect -3370 8975 -3325 9025
rect -3275 8975 -3205 9025
rect -3155 8975 -3110 9025
rect -3060 8975 -3015 9025
rect -2965 8975 -2915 9025
rect -2865 8975 -2815 9025
rect -2765 8975 -2715 9025
rect -2665 8975 -2620 9025
rect -2570 8975 -2525 9025
rect -2475 8975 -2405 9025
rect -2355 8975 -2310 9025
rect -2260 8975 -2215 9025
rect -2165 8975 -2115 9025
rect -2065 8975 -2015 9025
rect -1965 8975 -1915 9025
rect -1865 8975 -1820 9025
rect -1770 8975 -1725 9025
rect -1675 8975 -1640 9025
rect -4840 8935 -1640 8975
rect -4840 8885 -4805 8935
rect -4755 8885 -4710 8935
rect -4660 8885 -4615 8935
rect -4565 8885 -4515 8935
rect -4465 8885 -4415 8935
rect -4365 8885 -4315 8935
rect -4265 8885 -4220 8935
rect -4170 8885 -4125 8935
rect -4075 8885 -4005 8935
rect -3955 8885 -3910 8935
rect -3860 8885 -3815 8935
rect -3765 8885 -3715 8935
rect -3665 8885 -3615 8935
rect -3565 8885 -3515 8935
rect -3465 8885 -3420 8935
rect -3370 8885 -3325 8935
rect -3275 8885 -3205 8935
rect -3155 8885 -3110 8935
rect -3060 8885 -3015 8935
rect -2965 8885 -2915 8935
rect -2865 8885 -2815 8935
rect -2765 8885 -2715 8935
rect -2665 8885 -2620 8935
rect -2570 8885 -2525 8935
rect -2475 8885 -2405 8935
rect -2355 8885 -2310 8935
rect -2260 8885 -2215 8935
rect -2165 8885 -2115 8935
rect -2065 8885 -2015 8935
rect -1965 8885 -1915 8935
rect -1865 8885 -1820 8935
rect -1770 8885 -1725 8935
rect -1675 8885 -1640 8935
rect -4840 8815 -1640 8885
rect -4840 8765 -4805 8815
rect -4755 8765 -4710 8815
rect -4660 8765 -4615 8815
rect -4565 8765 -4515 8815
rect -4465 8765 -4415 8815
rect -4365 8765 -4315 8815
rect -4265 8765 -4220 8815
rect -4170 8765 -4125 8815
rect -4075 8765 -4005 8815
rect -3955 8765 -3910 8815
rect -3860 8765 -3815 8815
rect -3765 8765 -3715 8815
rect -3665 8765 -3615 8815
rect -3565 8765 -3515 8815
rect -3465 8765 -3420 8815
rect -3370 8765 -3325 8815
rect -3275 8765 -3205 8815
rect -3155 8765 -3110 8815
rect -3060 8765 -3015 8815
rect -2965 8765 -2915 8815
rect -2865 8765 -2815 8815
rect -2765 8765 -2715 8815
rect -2665 8765 -2620 8815
rect -2570 8765 -2525 8815
rect -2475 8765 -2405 8815
rect -2355 8765 -2310 8815
rect -2260 8765 -2215 8815
rect -2165 8765 -2115 8815
rect -2065 8765 -2015 8815
rect -1965 8765 -1915 8815
rect -1865 8765 -1820 8815
rect -1770 8765 -1725 8815
rect -1675 8765 -1640 8815
rect -4840 8725 -1640 8765
rect -4840 8675 -4805 8725
rect -4755 8675 -4710 8725
rect -4660 8675 -4615 8725
rect -4565 8675 -4515 8725
rect -4465 8675 -4415 8725
rect -4365 8675 -4315 8725
rect -4265 8675 -4220 8725
rect -4170 8675 -4125 8725
rect -4075 8675 -4005 8725
rect -3955 8675 -3910 8725
rect -3860 8675 -3815 8725
rect -3765 8675 -3715 8725
rect -3665 8675 -3615 8725
rect -3565 8675 -3515 8725
rect -3465 8675 -3420 8725
rect -3370 8675 -3325 8725
rect -3275 8675 -3205 8725
rect -3155 8675 -3110 8725
rect -3060 8675 -3015 8725
rect -2965 8675 -2915 8725
rect -2865 8675 -2815 8725
rect -2765 8675 -2715 8725
rect -2665 8675 -2620 8725
rect -2570 8675 -2525 8725
rect -2475 8675 -2405 8725
rect -2355 8675 -2310 8725
rect -2260 8675 -2215 8725
rect -2165 8675 -2115 8725
rect -2065 8675 -2015 8725
rect -1965 8675 -1915 8725
rect -1865 8675 -1820 8725
rect -1770 8675 -1725 8725
rect -1675 8675 -1640 8725
rect -4840 8625 -1640 8675
rect -4840 8575 -4805 8625
rect -4755 8575 -4710 8625
rect -4660 8575 -4615 8625
rect -4565 8575 -4515 8625
rect -4465 8575 -4415 8625
rect -4365 8575 -4315 8625
rect -4265 8575 -4220 8625
rect -4170 8575 -4125 8625
rect -4075 8575 -4005 8625
rect -3955 8575 -3910 8625
rect -3860 8575 -3815 8625
rect -3765 8575 -3715 8625
rect -3665 8575 -3615 8625
rect -3565 8575 -3515 8625
rect -3465 8575 -3420 8625
rect -3370 8575 -3325 8625
rect -3275 8575 -3205 8625
rect -3155 8575 -3110 8625
rect -3060 8575 -3015 8625
rect -2965 8575 -2915 8625
rect -2865 8575 -2815 8625
rect -2765 8575 -2715 8625
rect -2665 8575 -2620 8625
rect -2570 8575 -2525 8625
rect -2475 8575 -2405 8625
rect -2355 8575 -2310 8625
rect -2260 8575 -2215 8625
rect -2165 8575 -2115 8625
rect -2065 8575 -2015 8625
rect -1965 8575 -1915 8625
rect -1865 8575 -1820 8625
rect -1770 8575 -1725 8625
rect -1675 8575 -1640 8625
rect -4840 8535 -1640 8575
rect -4840 8485 -4805 8535
rect -4755 8485 -4710 8535
rect -4660 8485 -4615 8535
rect -4565 8485 -4515 8535
rect -4465 8485 -4415 8535
rect -4365 8485 -4315 8535
rect -4265 8485 -4220 8535
rect -4170 8485 -4125 8535
rect -4075 8485 -4005 8535
rect -3955 8485 -3910 8535
rect -3860 8485 -3815 8535
rect -3765 8485 -3715 8535
rect -3665 8485 -3615 8535
rect -3565 8485 -3515 8535
rect -3465 8485 -3420 8535
rect -3370 8485 -3325 8535
rect -3275 8485 -3205 8535
rect -3155 8485 -3110 8535
rect -3060 8485 -3015 8535
rect -2965 8485 -2915 8535
rect -2865 8485 -2815 8535
rect -2765 8485 -2715 8535
rect -2665 8485 -2620 8535
rect -2570 8485 -2525 8535
rect -2475 8485 -2405 8535
rect -2355 8485 -2310 8535
rect -2260 8485 -2215 8535
rect -2165 8485 -2115 8535
rect -2065 8485 -2015 8535
rect -1965 8485 -1915 8535
rect -1865 8485 -1820 8535
rect -1770 8485 -1725 8535
rect -1675 8485 -1640 8535
rect -4840 8415 -1640 8485
rect -4840 8365 -4805 8415
rect -4755 8365 -4710 8415
rect -4660 8365 -4615 8415
rect -4565 8365 -4515 8415
rect -4465 8365 -4415 8415
rect -4365 8365 -4315 8415
rect -4265 8365 -4220 8415
rect -4170 8365 -4125 8415
rect -4075 8365 -4005 8415
rect -3955 8365 -3910 8415
rect -3860 8365 -3815 8415
rect -3765 8365 -3715 8415
rect -3665 8365 -3615 8415
rect -3565 8365 -3515 8415
rect -3465 8365 -3420 8415
rect -3370 8365 -3325 8415
rect -3275 8365 -3205 8415
rect -3155 8365 -3110 8415
rect -3060 8365 -3015 8415
rect -2965 8365 -2915 8415
rect -2865 8365 -2815 8415
rect -2765 8365 -2715 8415
rect -2665 8365 -2620 8415
rect -2570 8365 -2525 8415
rect -2475 8365 -2405 8415
rect -2355 8365 -2310 8415
rect -2260 8365 -2215 8415
rect -2165 8365 -2115 8415
rect -2065 8365 -2015 8415
rect -1965 8365 -1915 8415
rect -1865 8365 -1820 8415
rect -1770 8365 -1725 8415
rect -1675 8365 -1640 8415
rect -4840 8325 -1640 8365
rect -4840 8275 -4805 8325
rect -4755 8275 -4710 8325
rect -4660 8275 -4615 8325
rect -4565 8275 -4515 8325
rect -4465 8275 -4415 8325
rect -4365 8275 -4315 8325
rect -4265 8275 -4220 8325
rect -4170 8275 -4125 8325
rect -4075 8275 -4005 8325
rect -3955 8275 -3910 8325
rect -3860 8275 -3815 8325
rect -3765 8275 -3715 8325
rect -3665 8275 -3615 8325
rect -3565 8275 -3515 8325
rect -3465 8275 -3420 8325
rect -3370 8275 -3325 8325
rect -3275 8275 -3205 8325
rect -3155 8275 -3110 8325
rect -3060 8275 -3015 8325
rect -2965 8275 -2915 8325
rect -2865 8275 -2815 8325
rect -2765 8275 -2715 8325
rect -2665 8275 -2620 8325
rect -2570 8275 -2525 8325
rect -2475 8275 -2405 8325
rect -2355 8275 -2310 8325
rect -2260 8275 -2215 8325
rect -2165 8275 -2115 8325
rect -2065 8275 -2015 8325
rect -1965 8275 -1915 8325
rect -1865 8275 -1820 8325
rect -1770 8275 -1725 8325
rect -1675 8275 -1640 8325
rect -4840 8225 -1640 8275
rect -4840 8175 -4805 8225
rect -4755 8175 -4710 8225
rect -4660 8175 -4615 8225
rect -4565 8175 -4515 8225
rect -4465 8175 -4415 8225
rect -4365 8175 -4315 8225
rect -4265 8175 -4220 8225
rect -4170 8175 -4125 8225
rect -4075 8175 -4005 8225
rect -3955 8175 -3910 8225
rect -3860 8175 -3815 8225
rect -3765 8175 -3715 8225
rect -3665 8175 -3615 8225
rect -3565 8175 -3515 8225
rect -3465 8175 -3420 8225
rect -3370 8175 -3325 8225
rect -3275 8175 -3205 8225
rect -3155 8175 -3110 8225
rect -3060 8175 -3015 8225
rect -2965 8175 -2915 8225
rect -2865 8175 -2815 8225
rect -2765 8175 -2715 8225
rect -2665 8175 -2620 8225
rect -2570 8175 -2525 8225
rect -2475 8175 -2405 8225
rect -2355 8175 -2310 8225
rect -2260 8175 -2215 8225
rect -2165 8175 -2115 8225
rect -2065 8175 -2015 8225
rect -1965 8175 -1915 8225
rect -1865 8175 -1820 8225
rect -1770 8175 -1725 8225
rect -1675 8175 -1640 8225
rect -4840 8135 -1640 8175
rect -4840 8085 -4805 8135
rect -4755 8085 -4710 8135
rect -4660 8085 -4615 8135
rect -4565 8085 -4515 8135
rect -4465 8085 -4415 8135
rect -4365 8085 -4315 8135
rect -4265 8085 -4220 8135
rect -4170 8085 -4125 8135
rect -4075 8085 -4005 8135
rect -3955 8085 -3910 8135
rect -3860 8085 -3815 8135
rect -3765 8085 -3715 8135
rect -3665 8085 -3615 8135
rect -3565 8085 -3515 8135
rect -3465 8085 -3420 8135
rect -3370 8085 -3325 8135
rect -3275 8085 -3205 8135
rect -3155 8085 -3110 8135
rect -3060 8085 -3015 8135
rect -2965 8085 -2915 8135
rect -2865 8085 -2815 8135
rect -2765 8085 -2715 8135
rect -2665 8085 -2620 8135
rect -2570 8085 -2525 8135
rect -2475 8085 -2405 8135
rect -2355 8085 -2310 8135
rect -2260 8085 -2215 8135
rect -2165 8085 -2115 8135
rect -2065 8085 -2015 8135
rect -1965 8085 -1915 8135
rect -1865 8085 -1820 8135
rect -1770 8085 -1725 8135
rect -1675 8085 -1640 8135
rect -4840 8015 -1640 8085
rect -4840 7965 -4805 8015
rect -4755 7965 -4710 8015
rect -4660 7965 -4615 8015
rect -4565 7965 -4515 8015
rect -4465 7965 -4415 8015
rect -4365 7965 -4315 8015
rect -4265 7965 -4220 8015
rect -4170 7965 -4125 8015
rect -4075 7965 -4005 8015
rect -3955 7965 -3910 8015
rect -3860 7965 -3815 8015
rect -3765 7965 -3715 8015
rect -3665 7965 -3615 8015
rect -3565 7965 -3515 8015
rect -3465 7965 -3420 8015
rect -3370 7965 -3325 8015
rect -3275 7965 -3205 8015
rect -3155 7965 -3110 8015
rect -3060 7965 -3015 8015
rect -2965 7965 -2915 8015
rect -2865 7965 -2815 8015
rect -2765 7965 -2715 8015
rect -2665 7965 -2620 8015
rect -2570 7965 -2525 8015
rect -2475 7965 -2405 8015
rect -2355 7965 -2310 8015
rect -2260 7965 -2215 8015
rect -2165 7965 -2115 8015
rect -2065 7965 -2015 8015
rect -1965 7965 -1915 8015
rect -1865 7965 -1820 8015
rect -1770 7965 -1725 8015
rect -1675 7965 -1640 8015
rect -4840 7925 -1640 7965
rect -4840 7875 -4805 7925
rect -4755 7875 -4710 7925
rect -4660 7875 -4615 7925
rect -4565 7875 -4515 7925
rect -4465 7875 -4415 7925
rect -4365 7875 -4315 7925
rect -4265 7875 -4220 7925
rect -4170 7875 -4125 7925
rect -4075 7875 -4005 7925
rect -3955 7875 -3910 7925
rect -3860 7875 -3815 7925
rect -3765 7875 -3715 7925
rect -3665 7875 -3615 7925
rect -3565 7875 -3515 7925
rect -3465 7875 -3420 7925
rect -3370 7875 -3325 7925
rect -3275 7875 -3205 7925
rect -3155 7875 -3110 7925
rect -3060 7875 -3015 7925
rect -2965 7875 -2915 7925
rect -2865 7875 -2815 7925
rect -2765 7875 -2715 7925
rect -2665 7875 -2620 7925
rect -2570 7875 -2525 7925
rect -2475 7875 -2405 7925
rect -2355 7875 -2310 7925
rect -2260 7875 -2215 7925
rect -2165 7875 -2115 7925
rect -2065 7875 -2015 7925
rect -1965 7875 -1915 7925
rect -1865 7875 -1820 7925
rect -1770 7875 -1725 7925
rect -1675 7875 -1640 7925
rect -4840 7825 -1640 7875
rect -4840 7775 -4805 7825
rect -4755 7775 -4710 7825
rect -4660 7775 -4615 7825
rect -4565 7775 -4515 7825
rect -4465 7775 -4415 7825
rect -4365 7775 -4315 7825
rect -4265 7775 -4220 7825
rect -4170 7775 -4125 7825
rect -4075 7775 -4005 7825
rect -3955 7775 -3910 7825
rect -3860 7775 -3815 7825
rect -3765 7775 -3715 7825
rect -3665 7775 -3615 7825
rect -3565 7775 -3515 7825
rect -3465 7775 -3420 7825
rect -3370 7775 -3325 7825
rect -3275 7775 -3205 7825
rect -3155 7775 -3110 7825
rect -3060 7775 -3015 7825
rect -2965 7775 -2915 7825
rect -2865 7775 -2815 7825
rect -2765 7775 -2715 7825
rect -2665 7775 -2620 7825
rect -2570 7775 -2525 7825
rect -2475 7775 -2405 7825
rect -2355 7775 -2310 7825
rect -2260 7775 -2215 7825
rect -2165 7775 -2115 7825
rect -2065 7775 -2015 7825
rect -1965 7775 -1915 7825
rect -1865 7775 -1820 7825
rect -1770 7775 -1725 7825
rect -1675 7775 -1640 7825
rect -4840 7735 -1640 7775
rect -4840 7685 -4805 7735
rect -4755 7685 -4710 7735
rect -4660 7685 -4615 7735
rect -4565 7685 -4515 7735
rect -4465 7685 -4415 7735
rect -4365 7685 -4315 7735
rect -4265 7685 -4220 7735
rect -4170 7685 -4125 7735
rect -4075 7685 -4005 7735
rect -3955 7685 -3910 7735
rect -3860 7685 -3815 7735
rect -3765 7685 -3715 7735
rect -3665 7685 -3615 7735
rect -3565 7685 -3515 7735
rect -3465 7685 -3420 7735
rect -3370 7685 -3325 7735
rect -3275 7685 -3205 7735
rect -3155 7685 -3110 7735
rect -3060 7685 -3015 7735
rect -2965 7685 -2915 7735
rect -2865 7685 -2815 7735
rect -2765 7685 -2715 7735
rect -2665 7685 -2620 7735
rect -2570 7685 -2525 7735
rect -2475 7685 -2405 7735
rect -2355 7685 -2310 7735
rect -2260 7685 -2215 7735
rect -2165 7685 -2115 7735
rect -2065 7685 -2015 7735
rect -1965 7685 -1915 7735
rect -1865 7685 -1820 7735
rect -1770 7685 -1725 7735
rect -1675 7685 -1640 7735
rect -4840 7615 -1640 7685
rect -4840 7565 -4805 7615
rect -4755 7565 -4710 7615
rect -4660 7565 -4615 7615
rect -4565 7565 -4515 7615
rect -4465 7565 -4415 7615
rect -4365 7565 -4315 7615
rect -4265 7565 -4220 7615
rect -4170 7565 -4125 7615
rect -4075 7565 -4005 7615
rect -3955 7565 -3910 7615
rect -3860 7565 -3815 7615
rect -3765 7565 -3715 7615
rect -3665 7565 -3615 7615
rect -3565 7565 -3515 7615
rect -3465 7565 -3420 7615
rect -3370 7565 -3325 7615
rect -3275 7565 -3205 7615
rect -3155 7565 -3110 7615
rect -3060 7565 -3015 7615
rect -2965 7565 -2915 7615
rect -2865 7565 -2815 7615
rect -2765 7565 -2715 7615
rect -2665 7565 -2620 7615
rect -2570 7565 -2525 7615
rect -2475 7565 -2405 7615
rect -2355 7565 -2310 7615
rect -2260 7565 -2215 7615
rect -2165 7565 -2115 7615
rect -2065 7565 -2015 7615
rect -1965 7565 -1915 7615
rect -1865 7565 -1820 7615
rect -1770 7565 -1725 7615
rect -1675 7565 -1640 7615
rect -4840 7525 -1640 7565
rect -4840 7475 -4805 7525
rect -4755 7475 -4710 7525
rect -4660 7475 -4615 7525
rect -4565 7475 -4515 7525
rect -4465 7475 -4415 7525
rect -4365 7475 -4315 7525
rect -4265 7475 -4220 7525
rect -4170 7475 -4125 7525
rect -4075 7475 -4005 7525
rect -3955 7475 -3910 7525
rect -3860 7475 -3815 7525
rect -3765 7475 -3715 7525
rect -3665 7475 -3615 7525
rect -3565 7475 -3515 7525
rect -3465 7475 -3420 7525
rect -3370 7475 -3325 7525
rect -3275 7475 -3205 7525
rect -3155 7475 -3110 7525
rect -3060 7475 -3015 7525
rect -2965 7475 -2915 7525
rect -2865 7475 -2815 7525
rect -2765 7475 -2715 7525
rect -2665 7475 -2620 7525
rect -2570 7475 -2525 7525
rect -2475 7475 -2405 7525
rect -2355 7475 -2310 7525
rect -2260 7475 -2215 7525
rect -2165 7475 -2115 7525
rect -2065 7475 -2015 7525
rect -1965 7475 -1915 7525
rect -1865 7475 -1820 7525
rect -1770 7475 -1725 7525
rect -1675 7475 -1640 7525
rect -4840 7425 -1640 7475
rect -4840 7375 -4805 7425
rect -4755 7375 -4710 7425
rect -4660 7375 -4615 7425
rect -4565 7375 -4515 7425
rect -4465 7375 -4415 7425
rect -4365 7375 -4315 7425
rect -4265 7375 -4220 7425
rect -4170 7375 -4125 7425
rect -4075 7375 -4005 7425
rect -3955 7375 -3910 7425
rect -3860 7375 -3815 7425
rect -3765 7375 -3715 7425
rect -3665 7375 -3615 7425
rect -3565 7375 -3515 7425
rect -3465 7375 -3420 7425
rect -3370 7375 -3325 7425
rect -3275 7375 -3205 7425
rect -3155 7375 -3110 7425
rect -3060 7375 -3015 7425
rect -2965 7375 -2915 7425
rect -2865 7375 -2815 7425
rect -2765 7375 -2715 7425
rect -2665 7375 -2620 7425
rect -2570 7375 -2525 7425
rect -2475 7375 -2405 7425
rect -2355 7375 -2310 7425
rect -2260 7375 -2215 7425
rect -2165 7375 -2115 7425
rect -2065 7375 -2015 7425
rect -1965 7375 -1915 7425
rect -1865 7375 -1820 7425
rect -1770 7375 -1725 7425
rect -1675 7375 -1640 7425
rect -4840 7335 -1640 7375
rect -4840 7285 -4805 7335
rect -4755 7285 -4710 7335
rect -4660 7285 -4615 7335
rect -4565 7285 -4515 7335
rect -4465 7285 -4415 7335
rect -4365 7285 -4315 7335
rect -4265 7285 -4220 7335
rect -4170 7285 -4125 7335
rect -4075 7285 -4005 7335
rect -3955 7285 -3910 7335
rect -3860 7285 -3815 7335
rect -3765 7285 -3715 7335
rect -3665 7285 -3615 7335
rect -3565 7285 -3515 7335
rect -3465 7285 -3420 7335
rect -3370 7285 -3325 7335
rect -3275 7285 -3205 7335
rect -3155 7285 -3110 7335
rect -3060 7285 -3015 7335
rect -2965 7285 -2915 7335
rect -2865 7285 -2815 7335
rect -2765 7285 -2715 7335
rect -2665 7285 -2620 7335
rect -2570 7285 -2525 7335
rect -2475 7285 -2405 7335
rect -2355 7285 -2310 7335
rect -2260 7285 -2215 7335
rect -2165 7285 -2115 7335
rect -2065 7285 -2015 7335
rect -1965 7285 -1915 7335
rect -1865 7285 -1820 7335
rect -1770 7285 -1725 7335
rect -1675 7285 -1640 7335
rect -4840 7215 -1640 7285
rect -4840 7165 -4805 7215
rect -4755 7165 -4710 7215
rect -4660 7165 -4615 7215
rect -4565 7165 -4515 7215
rect -4465 7165 -4415 7215
rect -4365 7165 -4315 7215
rect -4265 7165 -4220 7215
rect -4170 7165 -4125 7215
rect -4075 7165 -4005 7215
rect -3955 7165 -3910 7215
rect -3860 7165 -3815 7215
rect -3765 7165 -3715 7215
rect -3665 7165 -3615 7215
rect -3565 7165 -3515 7215
rect -3465 7165 -3420 7215
rect -3370 7165 -3325 7215
rect -3275 7165 -3205 7215
rect -3155 7165 -3110 7215
rect -3060 7165 -3015 7215
rect -2965 7165 -2915 7215
rect -2865 7165 -2815 7215
rect -2765 7165 -2715 7215
rect -2665 7165 -2620 7215
rect -2570 7165 -2525 7215
rect -2475 7165 -2405 7215
rect -2355 7165 -2310 7215
rect -2260 7165 -2215 7215
rect -2165 7165 -2115 7215
rect -2065 7165 -2015 7215
rect -1965 7165 -1915 7215
rect -1865 7165 -1820 7215
rect -1770 7165 -1725 7215
rect -1675 7165 -1640 7215
rect -4840 7125 -1640 7165
rect -4840 7075 -4805 7125
rect -4755 7075 -4710 7125
rect -4660 7075 -4615 7125
rect -4565 7075 -4515 7125
rect -4465 7075 -4415 7125
rect -4365 7075 -4315 7125
rect -4265 7075 -4220 7125
rect -4170 7075 -4125 7125
rect -4075 7075 -4005 7125
rect -3955 7075 -3910 7125
rect -3860 7075 -3815 7125
rect -3765 7075 -3715 7125
rect -3665 7075 -3615 7125
rect -3565 7075 -3515 7125
rect -3465 7075 -3420 7125
rect -3370 7075 -3325 7125
rect -3275 7075 -3205 7125
rect -3155 7075 -3110 7125
rect -3060 7075 -3015 7125
rect -2965 7075 -2915 7125
rect -2865 7075 -2815 7125
rect -2765 7075 -2715 7125
rect -2665 7075 -2620 7125
rect -2570 7075 -2525 7125
rect -2475 7075 -2405 7125
rect -2355 7075 -2310 7125
rect -2260 7075 -2215 7125
rect -2165 7075 -2115 7125
rect -2065 7075 -2015 7125
rect -1965 7075 -1915 7125
rect -1865 7075 -1820 7125
rect -1770 7075 -1725 7125
rect -1675 7075 -1640 7125
rect -4840 7025 -1640 7075
rect -4840 6975 -4805 7025
rect -4755 6975 -4710 7025
rect -4660 6975 -4615 7025
rect -4565 6975 -4515 7025
rect -4465 6975 -4415 7025
rect -4365 6975 -4315 7025
rect -4265 6975 -4220 7025
rect -4170 6975 -4125 7025
rect -4075 6975 -4005 7025
rect -3955 6975 -3910 7025
rect -3860 6975 -3815 7025
rect -3765 6975 -3715 7025
rect -3665 6975 -3615 7025
rect -3565 6975 -3515 7025
rect -3465 6975 -3420 7025
rect -3370 6975 -3325 7025
rect -3275 6975 -3205 7025
rect -3155 6975 -3110 7025
rect -3060 6975 -3015 7025
rect -2965 6975 -2915 7025
rect -2865 6975 -2815 7025
rect -2765 6975 -2715 7025
rect -2665 6975 -2620 7025
rect -2570 6975 -2525 7025
rect -2475 6975 -2405 7025
rect -2355 6975 -2310 7025
rect -2260 6975 -2215 7025
rect -2165 6975 -2115 7025
rect -2065 6975 -2015 7025
rect -1965 6975 -1915 7025
rect -1865 6975 -1820 7025
rect -1770 6975 -1725 7025
rect -1675 6975 -1640 7025
rect -4840 6935 -1640 6975
rect -4840 6885 -4805 6935
rect -4755 6885 -4710 6935
rect -4660 6885 -4615 6935
rect -4565 6885 -4515 6935
rect -4465 6885 -4415 6935
rect -4365 6885 -4315 6935
rect -4265 6885 -4220 6935
rect -4170 6885 -4125 6935
rect -4075 6885 -4005 6935
rect -3955 6885 -3910 6935
rect -3860 6885 -3815 6935
rect -3765 6885 -3715 6935
rect -3665 6885 -3615 6935
rect -3565 6885 -3515 6935
rect -3465 6885 -3420 6935
rect -3370 6885 -3325 6935
rect -3275 6885 -3205 6935
rect -3155 6885 -3110 6935
rect -3060 6885 -3015 6935
rect -2965 6885 -2915 6935
rect -2865 6885 -2815 6935
rect -2765 6885 -2715 6935
rect -2665 6885 -2620 6935
rect -2570 6885 -2525 6935
rect -2475 6885 -2405 6935
rect -2355 6885 -2310 6935
rect -2260 6885 -2215 6935
rect -2165 6885 -2115 6935
rect -2065 6885 -2015 6935
rect -1965 6885 -1915 6935
rect -1865 6885 -1820 6935
rect -1770 6885 -1725 6935
rect -1675 6885 -1640 6935
rect -4840 6815 -1640 6885
rect -4840 6765 -4805 6815
rect -4755 6765 -4710 6815
rect -4660 6765 -4615 6815
rect -4565 6765 -4515 6815
rect -4465 6765 -4415 6815
rect -4365 6765 -4315 6815
rect -4265 6765 -4220 6815
rect -4170 6765 -4125 6815
rect -4075 6765 -4005 6815
rect -3955 6765 -3910 6815
rect -3860 6765 -3815 6815
rect -3765 6765 -3715 6815
rect -3665 6765 -3615 6815
rect -3565 6765 -3515 6815
rect -3465 6765 -3420 6815
rect -3370 6765 -3325 6815
rect -3275 6765 -3205 6815
rect -3155 6765 -3110 6815
rect -3060 6765 -3015 6815
rect -2965 6765 -2915 6815
rect -2865 6765 -2815 6815
rect -2765 6765 -2715 6815
rect -2665 6765 -2620 6815
rect -2570 6765 -2525 6815
rect -2475 6765 -2405 6815
rect -2355 6765 -2310 6815
rect -2260 6765 -2215 6815
rect -2165 6765 -2115 6815
rect -2065 6765 -2015 6815
rect -1965 6765 -1915 6815
rect -1865 6765 -1820 6815
rect -1770 6765 -1725 6815
rect -1675 6765 -1640 6815
rect -4840 6725 -1640 6765
rect -4840 6675 -4805 6725
rect -4755 6675 -4710 6725
rect -4660 6675 -4615 6725
rect -4565 6675 -4515 6725
rect -4465 6675 -4415 6725
rect -4365 6675 -4315 6725
rect -4265 6675 -4220 6725
rect -4170 6675 -4125 6725
rect -4075 6675 -4005 6725
rect -3955 6675 -3910 6725
rect -3860 6675 -3815 6725
rect -3765 6675 -3715 6725
rect -3665 6675 -3615 6725
rect -3565 6675 -3515 6725
rect -3465 6675 -3420 6725
rect -3370 6675 -3325 6725
rect -3275 6675 -3205 6725
rect -3155 6675 -3110 6725
rect -3060 6675 -3015 6725
rect -2965 6675 -2915 6725
rect -2865 6675 -2815 6725
rect -2765 6675 -2715 6725
rect -2665 6675 -2620 6725
rect -2570 6675 -2525 6725
rect -2475 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6675 -1640 6725
rect -4840 6625 -1640 6675
rect -4840 6575 -4805 6625
rect -4755 6575 -4710 6625
rect -4660 6575 -4615 6625
rect -4565 6575 -4515 6625
rect -4465 6575 -4415 6625
rect -4365 6575 -4315 6625
rect -4265 6575 -4220 6625
rect -4170 6575 -4125 6625
rect -4075 6575 -4005 6625
rect -3955 6575 -3910 6625
rect -3860 6575 -3815 6625
rect -3765 6575 -3715 6625
rect -3665 6575 -3615 6625
rect -3565 6575 -3515 6625
rect -3465 6575 -3420 6625
rect -3370 6575 -3325 6625
rect -3275 6575 -3205 6625
rect -3155 6575 -3110 6625
rect -3060 6575 -3015 6625
rect -2965 6575 -2915 6625
rect -2865 6575 -2815 6625
rect -2765 6575 -2715 6625
rect -2665 6575 -2620 6625
rect -2570 6575 -2525 6625
rect -2475 6575 -2405 6625
rect -2355 6575 -2310 6625
rect -2260 6575 -2215 6625
rect -2165 6575 -2115 6625
rect -2065 6575 -2015 6625
rect -1965 6575 -1915 6625
rect -1865 6575 -1820 6625
rect -1770 6575 -1725 6625
rect -1675 6575 -1640 6625
rect -4840 6535 -1640 6575
rect -4840 6485 -4805 6535
rect -4755 6485 -4710 6535
rect -4660 6485 -4615 6535
rect -4565 6485 -4515 6535
rect -4465 6485 -4415 6535
rect -4365 6485 -4315 6535
rect -4265 6485 -4220 6535
rect -4170 6485 -4125 6535
rect -4075 6485 -4005 6535
rect -3955 6485 -3910 6535
rect -3860 6485 -3815 6535
rect -3765 6485 -3715 6535
rect -3665 6485 -3615 6535
rect -3565 6485 -3515 6535
rect -3465 6485 -3420 6535
rect -3370 6485 -3325 6535
rect -3275 6485 -3205 6535
rect -3155 6485 -3110 6535
rect -3060 6485 -3015 6535
rect -2965 6485 -2915 6535
rect -2865 6485 -2815 6535
rect -2765 6485 -2715 6535
rect -2665 6485 -2620 6535
rect -2570 6485 -2525 6535
rect -2475 6485 -2405 6535
rect -2355 6485 -2310 6535
rect -2260 6485 -2215 6535
rect -2165 6485 -2115 6535
rect -2065 6485 -2015 6535
rect -1965 6485 -1915 6535
rect -1865 6485 -1820 6535
rect -1770 6485 -1725 6535
rect -1675 6485 -1640 6535
rect -4840 6450 -1640 6485
rect -90 9640 -30 9650
rect -90 9600 -80 9640
rect -40 9600 -30 9640
rect -90 9575 -30 9600
rect -90 9535 -80 9575
rect -40 9535 -30 9575
rect -90 9505 -30 9535
rect -90 9465 -80 9505
rect -40 9465 -30 9505
rect -90 9435 -30 9465
rect -90 9395 -80 9435
rect -40 9395 -30 9435
rect -90 9365 -30 9395
rect -90 9325 -80 9365
rect -40 9325 -30 9365
rect -90 9300 -30 9325
rect -90 9260 -80 9300
rect -40 9260 -30 9300
rect -90 9240 -30 9260
rect -90 9200 -80 9240
rect -40 9200 -30 9240
rect -90 9175 -30 9200
rect -90 9135 -80 9175
rect -40 9135 -30 9175
rect -90 9105 -30 9135
rect -90 9065 -80 9105
rect -40 9065 -30 9105
rect -90 9035 -30 9065
rect -90 8995 -80 9035
rect -40 8995 -30 9035
rect -90 8965 -30 8995
rect -90 8925 -80 8965
rect -40 8925 -30 8965
rect -90 8900 -30 8925
rect -90 8860 -80 8900
rect -40 8860 -30 8900
rect -90 8840 -30 8860
rect -90 8800 -80 8840
rect -40 8800 -30 8840
rect -90 8775 -30 8800
rect -90 8735 -80 8775
rect -40 8735 -30 8775
rect -90 8705 -30 8735
rect -90 8665 -80 8705
rect -40 8665 -30 8705
rect -90 8635 -30 8665
rect -90 8595 -80 8635
rect -40 8595 -30 8635
rect -90 8565 -30 8595
rect -90 8525 -80 8565
rect -40 8525 -30 8565
rect -90 8500 -30 8525
rect -90 8460 -80 8500
rect -40 8460 -30 8500
rect -90 8440 -30 8460
rect -90 8400 -80 8440
rect -40 8400 -30 8440
rect -90 8375 -30 8400
rect -90 8335 -80 8375
rect -40 8335 -30 8375
rect -90 8305 -30 8335
rect -90 8265 -80 8305
rect -40 8265 -30 8305
rect -90 8235 -30 8265
rect -90 8195 -80 8235
rect -40 8195 -30 8235
rect -90 8165 -30 8195
rect -90 8125 -80 8165
rect -40 8125 -30 8165
rect -90 8100 -30 8125
rect -90 8060 -80 8100
rect -40 8060 -30 8100
rect -90 8040 -30 8060
rect -90 8000 -80 8040
rect -40 8000 -30 8040
rect -90 7975 -30 8000
rect -90 7935 -80 7975
rect -40 7935 -30 7975
rect -90 7905 -30 7935
rect -90 7865 -80 7905
rect -40 7865 -30 7905
rect -90 7835 -30 7865
rect -90 7795 -80 7835
rect -40 7795 -30 7835
rect -90 7765 -30 7795
rect -90 7725 -80 7765
rect -40 7725 -30 7765
rect -90 7700 -30 7725
rect -90 7660 -80 7700
rect -40 7660 -30 7700
rect -90 7640 -30 7660
rect -90 7600 -80 7640
rect -40 7600 -30 7640
rect -90 7575 -30 7600
rect -90 7535 -80 7575
rect -40 7535 -30 7575
rect -90 7505 -30 7535
rect -90 7465 -80 7505
rect -40 7465 -30 7505
rect -90 7435 -30 7465
rect -90 7395 -80 7435
rect -40 7395 -30 7435
rect -90 7365 -30 7395
rect -90 7325 -80 7365
rect -40 7325 -30 7365
rect -90 7300 -30 7325
rect -90 7260 -80 7300
rect -40 7260 -30 7300
rect -90 7240 -30 7260
rect -90 7200 -80 7240
rect -40 7200 -30 7240
rect -90 7175 -30 7200
rect -90 7135 -80 7175
rect -40 7135 -30 7175
rect -90 7105 -30 7135
rect -90 7065 -80 7105
rect -40 7065 -30 7105
rect -90 7035 -30 7065
rect -90 6995 -80 7035
rect -40 6995 -30 7035
rect -90 6965 -30 6995
rect -90 6925 -80 6965
rect -40 6925 -30 6965
rect -90 6900 -30 6925
rect -90 6860 -80 6900
rect -40 6860 -30 6900
rect -90 6840 -30 6860
rect -90 6800 -80 6840
rect -40 6800 -30 6840
rect -90 6775 -30 6800
rect -90 6735 -80 6775
rect -40 6735 -30 6775
rect -90 6705 -30 6735
rect -90 6665 -80 6705
rect -40 6665 -30 6705
rect -90 6635 -30 6665
rect -90 6595 -80 6635
rect -40 6595 -30 6635
rect -90 6565 -30 6595
rect -90 6525 -80 6565
rect -40 6525 -30 6565
rect -90 6500 -30 6525
rect -90 6460 -80 6500
rect -40 6460 -30 6500
rect -90 6450 -30 6460
rect 260 9640 320 9650
rect 260 9600 270 9640
rect 310 9600 320 9640
rect 260 9575 320 9600
rect 260 9535 270 9575
rect 310 9535 320 9575
rect 260 9505 320 9535
rect 260 9465 270 9505
rect 310 9465 320 9505
rect 260 9435 320 9465
rect 260 9395 270 9435
rect 310 9395 320 9435
rect 260 9365 320 9395
rect 260 9325 270 9365
rect 310 9325 320 9365
rect 260 9300 320 9325
rect 260 9260 270 9300
rect 310 9260 320 9300
rect 260 9240 320 9260
rect 260 9200 270 9240
rect 310 9200 320 9240
rect 260 9175 320 9200
rect 260 9135 270 9175
rect 310 9135 320 9175
rect 260 9105 320 9135
rect 260 9065 270 9105
rect 310 9065 320 9105
rect 260 9035 320 9065
rect 260 8995 270 9035
rect 310 8995 320 9035
rect 260 8965 320 8995
rect 260 8925 270 8965
rect 310 8925 320 8965
rect 260 8900 320 8925
rect 260 8860 270 8900
rect 310 8860 320 8900
rect 260 8840 320 8860
rect 260 8800 270 8840
rect 310 8800 320 8840
rect 260 8775 320 8800
rect 260 8735 270 8775
rect 310 8735 320 8775
rect 260 8705 320 8735
rect 260 8665 270 8705
rect 310 8665 320 8705
rect 260 8635 320 8665
rect 260 8595 270 8635
rect 310 8595 320 8635
rect 260 8565 320 8595
rect 260 8525 270 8565
rect 310 8525 320 8565
rect 260 8500 320 8525
rect 260 8460 270 8500
rect 310 8460 320 8500
rect 260 8440 320 8460
rect 260 8400 270 8440
rect 310 8400 320 8440
rect 260 8375 320 8400
rect 260 8335 270 8375
rect 310 8335 320 8375
rect 260 8305 320 8335
rect 260 8265 270 8305
rect 310 8265 320 8305
rect 260 8235 320 8265
rect 260 8195 270 8235
rect 310 8195 320 8235
rect 260 8165 320 8195
rect 260 8125 270 8165
rect 310 8125 320 8165
rect 260 8100 320 8125
rect 260 8060 270 8100
rect 310 8060 320 8100
rect 260 8040 320 8060
rect 260 8000 270 8040
rect 310 8000 320 8040
rect 260 7975 320 8000
rect 260 7935 270 7975
rect 310 7935 320 7975
rect 260 7905 320 7935
rect 260 7865 270 7905
rect 310 7865 320 7905
rect 260 7835 320 7865
rect 260 7795 270 7835
rect 310 7795 320 7835
rect 260 7765 320 7795
rect 260 7725 270 7765
rect 310 7725 320 7765
rect 260 7700 320 7725
rect 260 7660 270 7700
rect 310 7660 320 7700
rect 260 7640 320 7660
rect 260 7600 270 7640
rect 310 7600 320 7640
rect 260 7575 320 7600
rect 260 7535 270 7575
rect 310 7535 320 7575
rect 260 7505 320 7535
rect 260 7465 270 7505
rect 310 7465 320 7505
rect 260 7435 320 7465
rect 260 7395 270 7435
rect 310 7395 320 7435
rect 260 7365 320 7395
rect 260 7325 270 7365
rect 310 7325 320 7365
rect 260 7300 320 7325
rect 260 7260 270 7300
rect 310 7260 320 7300
rect 260 7240 320 7260
rect 260 7200 270 7240
rect 310 7200 320 7240
rect 260 7175 320 7200
rect 260 7135 270 7175
rect 310 7135 320 7175
rect 260 7105 320 7135
rect 260 7065 270 7105
rect 310 7065 320 7105
rect 260 7035 320 7065
rect 260 6995 270 7035
rect 310 6995 320 7035
rect 260 6965 320 6995
rect 260 6925 270 6965
rect 310 6925 320 6965
rect 260 6900 320 6925
rect 260 6860 270 6900
rect 310 6860 320 6900
rect 260 6840 320 6860
rect 260 6800 270 6840
rect 310 6800 320 6840
rect 260 6775 320 6800
rect 260 6735 270 6775
rect 310 6735 320 6775
rect 260 6705 320 6735
rect 260 6665 270 6705
rect 310 6665 320 6705
rect 260 6635 320 6665
rect 260 6595 270 6635
rect 310 6595 320 6635
rect 260 6565 320 6595
rect 260 6525 270 6565
rect 310 6525 320 6565
rect 260 6500 320 6525
rect 260 6460 270 6500
rect 310 6460 320 6500
rect 260 6450 320 6460
rect 610 9640 670 9650
rect 610 9600 620 9640
rect 660 9600 670 9640
rect 610 9575 670 9600
rect 610 9535 620 9575
rect 660 9535 670 9575
rect 610 9505 670 9535
rect 610 9465 620 9505
rect 660 9465 670 9505
rect 610 9435 670 9465
rect 610 9395 620 9435
rect 660 9395 670 9435
rect 610 9365 670 9395
rect 610 9325 620 9365
rect 660 9325 670 9365
rect 610 9300 670 9325
rect 610 9260 620 9300
rect 660 9260 670 9300
rect 610 9240 670 9260
rect 610 9200 620 9240
rect 660 9200 670 9240
rect 610 9175 670 9200
rect 610 9135 620 9175
rect 660 9135 670 9175
rect 610 9105 670 9135
rect 610 9065 620 9105
rect 660 9065 670 9105
rect 610 9035 670 9065
rect 610 8995 620 9035
rect 660 8995 670 9035
rect 610 8965 670 8995
rect 610 8925 620 8965
rect 660 8925 670 8965
rect 610 8900 670 8925
rect 610 8860 620 8900
rect 660 8860 670 8900
rect 610 8840 670 8860
rect 610 8800 620 8840
rect 660 8800 670 8840
rect 610 8775 670 8800
rect 610 8735 620 8775
rect 660 8735 670 8775
rect 610 8705 670 8735
rect 610 8665 620 8705
rect 660 8665 670 8705
rect 610 8635 670 8665
rect 610 8595 620 8635
rect 660 8595 670 8635
rect 610 8565 670 8595
rect 610 8525 620 8565
rect 660 8525 670 8565
rect 610 8500 670 8525
rect 610 8460 620 8500
rect 660 8460 670 8500
rect 610 8440 670 8460
rect 610 8400 620 8440
rect 660 8400 670 8440
rect 610 8375 670 8400
rect 610 8335 620 8375
rect 660 8335 670 8375
rect 610 8305 670 8335
rect 610 8265 620 8305
rect 660 8265 670 8305
rect 610 8235 670 8265
rect 610 8195 620 8235
rect 660 8195 670 8235
rect 610 8165 670 8195
rect 610 8125 620 8165
rect 660 8125 670 8165
rect 610 8100 670 8125
rect 610 8060 620 8100
rect 660 8060 670 8100
rect 610 8040 670 8060
rect 610 8000 620 8040
rect 660 8000 670 8040
rect 610 7975 670 8000
rect 610 7935 620 7975
rect 660 7935 670 7975
rect 610 7905 670 7935
rect 610 7865 620 7905
rect 660 7865 670 7905
rect 610 7835 670 7865
rect 610 7795 620 7835
rect 660 7795 670 7835
rect 610 7765 670 7795
rect 610 7725 620 7765
rect 660 7725 670 7765
rect 610 7700 670 7725
rect 610 7660 620 7700
rect 660 7660 670 7700
rect 610 7640 670 7660
rect 610 7600 620 7640
rect 660 7600 670 7640
rect 610 7575 670 7600
rect 610 7535 620 7575
rect 660 7535 670 7575
rect 610 7505 670 7535
rect 610 7465 620 7505
rect 660 7465 670 7505
rect 610 7435 670 7465
rect 610 7395 620 7435
rect 660 7395 670 7435
rect 610 7365 670 7395
rect 610 7325 620 7365
rect 660 7325 670 7365
rect 610 7300 670 7325
rect 610 7260 620 7300
rect 660 7260 670 7300
rect 610 7240 670 7260
rect 610 7200 620 7240
rect 660 7200 670 7240
rect 610 7175 670 7200
rect 610 7135 620 7175
rect 660 7135 670 7175
rect 610 7105 670 7135
rect 610 7065 620 7105
rect 660 7065 670 7105
rect 610 7035 670 7065
rect 610 6995 620 7035
rect 660 6995 670 7035
rect 610 6965 670 6995
rect 610 6925 620 6965
rect 660 6925 670 6965
rect 610 6900 670 6925
rect 610 6860 620 6900
rect 660 6860 670 6900
rect 610 6840 670 6860
rect 610 6800 620 6840
rect 660 6800 670 6840
rect 610 6775 670 6800
rect 610 6735 620 6775
rect 660 6735 670 6775
rect 610 6705 670 6735
rect 610 6665 620 6705
rect 660 6665 670 6705
rect 610 6635 670 6665
rect 610 6595 620 6635
rect 660 6595 670 6635
rect 610 6565 670 6595
rect 610 6525 620 6565
rect 660 6525 670 6565
rect 610 6500 670 6525
rect 610 6460 620 6500
rect 660 6460 670 6500
rect 610 6450 670 6460
rect 1310 9640 1370 9650
rect 1310 9600 1320 9640
rect 1360 9600 1370 9640
rect 1310 9575 1370 9600
rect 1310 9535 1320 9575
rect 1360 9535 1370 9575
rect 1310 9505 1370 9535
rect 1310 9465 1320 9505
rect 1360 9465 1370 9505
rect 1310 9435 1370 9465
rect 1310 9395 1320 9435
rect 1360 9395 1370 9435
rect 1310 9365 1370 9395
rect 1310 9325 1320 9365
rect 1360 9325 1370 9365
rect 1310 9300 1370 9325
rect 1310 9260 1320 9300
rect 1360 9260 1370 9300
rect 1310 9240 1370 9260
rect 1310 9200 1320 9240
rect 1360 9200 1370 9240
rect 1310 9175 1370 9200
rect 1310 9135 1320 9175
rect 1360 9135 1370 9175
rect 1310 9105 1370 9135
rect 1310 9065 1320 9105
rect 1360 9065 1370 9105
rect 1310 9035 1370 9065
rect 1310 8995 1320 9035
rect 1360 8995 1370 9035
rect 1310 8965 1370 8995
rect 1310 8925 1320 8965
rect 1360 8925 1370 8965
rect 1310 8900 1370 8925
rect 1310 8860 1320 8900
rect 1360 8860 1370 8900
rect 1310 8840 1370 8860
rect 1310 8800 1320 8840
rect 1360 8800 1370 8840
rect 1310 8775 1370 8800
rect 1310 8735 1320 8775
rect 1360 8735 1370 8775
rect 1310 8705 1370 8735
rect 1310 8665 1320 8705
rect 1360 8665 1370 8705
rect 1310 8635 1370 8665
rect 1310 8595 1320 8635
rect 1360 8595 1370 8635
rect 1310 8565 1370 8595
rect 1310 8525 1320 8565
rect 1360 8525 1370 8565
rect 1310 8500 1370 8525
rect 1310 8460 1320 8500
rect 1360 8460 1370 8500
rect 1310 8440 1370 8460
rect 1310 8400 1320 8440
rect 1360 8400 1370 8440
rect 1310 8375 1370 8400
rect 1310 8335 1320 8375
rect 1360 8335 1370 8375
rect 1310 8305 1370 8335
rect 1310 8265 1320 8305
rect 1360 8265 1370 8305
rect 1310 8235 1370 8265
rect 1310 8195 1320 8235
rect 1360 8195 1370 8235
rect 1310 8165 1370 8195
rect 1310 8125 1320 8165
rect 1360 8125 1370 8165
rect 1310 8100 1370 8125
rect 1310 8060 1320 8100
rect 1360 8060 1370 8100
rect 1310 8040 1370 8060
rect 1310 8000 1320 8040
rect 1360 8000 1370 8040
rect 1310 7975 1370 8000
rect 1310 7935 1320 7975
rect 1360 7935 1370 7975
rect 1310 7905 1370 7935
rect 1310 7865 1320 7905
rect 1360 7865 1370 7905
rect 1310 7835 1370 7865
rect 1310 7795 1320 7835
rect 1360 7795 1370 7835
rect 1310 7765 1370 7795
rect 1310 7725 1320 7765
rect 1360 7725 1370 7765
rect 1310 7700 1370 7725
rect 1310 7660 1320 7700
rect 1360 7660 1370 7700
rect 1310 7640 1370 7660
rect 1310 7600 1320 7640
rect 1360 7600 1370 7640
rect 1310 7575 1370 7600
rect 1310 7535 1320 7575
rect 1360 7535 1370 7575
rect 1310 7505 1370 7535
rect 1310 7465 1320 7505
rect 1360 7465 1370 7505
rect 1310 7435 1370 7465
rect 1310 7395 1320 7435
rect 1360 7395 1370 7435
rect 1310 7365 1370 7395
rect 1310 7325 1320 7365
rect 1360 7325 1370 7365
rect 1310 7300 1370 7325
rect 1310 7260 1320 7300
rect 1360 7260 1370 7300
rect 1310 7240 1370 7260
rect 1310 7200 1320 7240
rect 1360 7200 1370 7240
rect 1310 7175 1370 7200
rect 1310 7135 1320 7175
rect 1360 7135 1370 7175
rect 1310 7105 1370 7135
rect 1310 7065 1320 7105
rect 1360 7065 1370 7105
rect 1310 7035 1370 7065
rect 1310 6995 1320 7035
rect 1360 6995 1370 7035
rect 1310 6965 1370 6995
rect 1310 6925 1320 6965
rect 1360 6925 1370 6965
rect 1310 6900 1370 6925
rect 1310 6860 1320 6900
rect 1360 6860 1370 6900
rect 1310 6840 1370 6860
rect 1310 6800 1320 6840
rect 1360 6800 1370 6840
rect 1310 6775 1370 6800
rect 1310 6735 1320 6775
rect 1360 6735 1370 6775
rect 1310 6705 1370 6735
rect 1310 6665 1320 6705
rect 1360 6665 1370 6705
rect 1310 6635 1370 6665
rect 1310 6595 1320 6635
rect 1360 6595 1370 6635
rect 1310 6565 1370 6595
rect 1310 6525 1320 6565
rect 1360 6525 1370 6565
rect 1310 6500 1370 6525
rect 1310 6460 1320 6500
rect 1360 6460 1370 6500
rect 1310 6450 1370 6460
rect 1660 9640 1720 9650
rect 1660 9600 1670 9640
rect 1710 9600 1720 9640
rect 1660 9575 1720 9600
rect 1660 9535 1670 9575
rect 1710 9535 1720 9575
rect 1660 9505 1720 9535
rect 1660 9465 1670 9505
rect 1710 9465 1720 9505
rect 1660 9435 1720 9465
rect 1660 9395 1670 9435
rect 1710 9395 1720 9435
rect 1660 9365 1720 9395
rect 1660 9325 1670 9365
rect 1710 9325 1720 9365
rect 1660 9300 1720 9325
rect 1660 9260 1670 9300
rect 1710 9260 1720 9300
rect 1660 9240 1720 9260
rect 1660 9200 1670 9240
rect 1710 9200 1720 9240
rect 1660 9175 1720 9200
rect 1660 9135 1670 9175
rect 1710 9135 1720 9175
rect 1660 9105 1720 9135
rect 1660 9065 1670 9105
rect 1710 9065 1720 9105
rect 1660 9035 1720 9065
rect 1660 8995 1670 9035
rect 1710 8995 1720 9035
rect 1660 8965 1720 8995
rect 1660 8925 1670 8965
rect 1710 8925 1720 8965
rect 1660 8900 1720 8925
rect 1660 8860 1670 8900
rect 1710 8860 1720 8900
rect 1660 8840 1720 8860
rect 1660 8800 1670 8840
rect 1710 8800 1720 8840
rect 1660 8775 1720 8800
rect 1660 8735 1670 8775
rect 1710 8735 1720 8775
rect 1660 8705 1720 8735
rect 1660 8665 1670 8705
rect 1710 8665 1720 8705
rect 1660 8635 1720 8665
rect 1660 8595 1670 8635
rect 1710 8595 1720 8635
rect 1660 8565 1720 8595
rect 1660 8525 1670 8565
rect 1710 8525 1720 8565
rect 1660 8500 1720 8525
rect 1660 8460 1670 8500
rect 1710 8460 1720 8500
rect 1660 8440 1720 8460
rect 1660 8400 1670 8440
rect 1710 8400 1720 8440
rect 1660 8375 1720 8400
rect 1660 8335 1670 8375
rect 1710 8335 1720 8375
rect 1660 8305 1720 8335
rect 1660 8265 1670 8305
rect 1710 8265 1720 8305
rect 1660 8235 1720 8265
rect 1660 8195 1670 8235
rect 1710 8195 1720 8235
rect 1660 8165 1720 8195
rect 1660 8125 1670 8165
rect 1710 8125 1720 8165
rect 1660 8100 1720 8125
rect 1660 8060 1670 8100
rect 1710 8060 1720 8100
rect 1660 8040 1720 8060
rect 1660 8000 1670 8040
rect 1710 8000 1720 8040
rect 1660 7975 1720 8000
rect 1660 7935 1670 7975
rect 1710 7935 1720 7975
rect 1660 7905 1720 7935
rect 1660 7865 1670 7905
rect 1710 7865 1720 7905
rect 1660 7835 1720 7865
rect 1660 7795 1670 7835
rect 1710 7795 1720 7835
rect 1660 7765 1720 7795
rect 1660 7725 1670 7765
rect 1710 7725 1720 7765
rect 1660 7700 1720 7725
rect 1660 7660 1670 7700
rect 1710 7660 1720 7700
rect 1660 7640 1720 7660
rect 1660 7600 1670 7640
rect 1710 7600 1720 7640
rect 1660 7575 1720 7600
rect 1660 7535 1670 7575
rect 1710 7535 1720 7575
rect 1660 7505 1720 7535
rect 1660 7465 1670 7505
rect 1710 7465 1720 7505
rect 1660 7435 1720 7465
rect 1660 7395 1670 7435
rect 1710 7395 1720 7435
rect 1660 7365 1720 7395
rect 1660 7325 1670 7365
rect 1710 7325 1720 7365
rect 1660 7300 1720 7325
rect 1660 7260 1670 7300
rect 1710 7260 1720 7300
rect 1660 7240 1720 7260
rect 1660 7200 1670 7240
rect 1710 7200 1720 7240
rect 1660 7175 1720 7200
rect 1660 7135 1670 7175
rect 1710 7135 1720 7175
rect 1660 7105 1720 7135
rect 1660 7065 1670 7105
rect 1710 7065 1720 7105
rect 1660 7035 1720 7065
rect 1660 6995 1670 7035
rect 1710 6995 1720 7035
rect 1660 6965 1720 6995
rect 1660 6925 1670 6965
rect 1710 6925 1720 6965
rect 1660 6900 1720 6925
rect 1660 6860 1670 6900
rect 1710 6860 1720 6900
rect 1660 6840 1720 6860
rect 1660 6800 1670 6840
rect 1710 6800 1720 6840
rect 1660 6775 1720 6800
rect 1660 6735 1670 6775
rect 1710 6735 1720 6775
rect 1660 6705 1720 6735
rect 1660 6665 1670 6705
rect 1710 6665 1720 6705
rect 1660 6635 1720 6665
rect 1660 6595 1670 6635
rect 1710 6595 1720 6635
rect 1660 6565 1720 6595
rect 1660 6525 1670 6565
rect 1710 6525 1720 6565
rect 1660 6500 1720 6525
rect 1660 6460 1670 6500
rect 1710 6460 1720 6500
rect 1660 6450 1720 6460
rect 2375 9640 2435 9650
rect 2375 9600 2385 9640
rect 2425 9600 2435 9640
rect 2375 9575 2435 9600
rect 2375 9535 2385 9575
rect 2425 9535 2435 9575
rect 2375 9505 2435 9535
rect 2375 9465 2385 9505
rect 2425 9465 2435 9505
rect 2375 9435 2435 9465
rect 2375 9395 2385 9435
rect 2425 9395 2435 9435
rect 2375 9365 2435 9395
rect 2375 9325 2385 9365
rect 2425 9325 2435 9365
rect 2375 9300 2435 9325
rect 2375 9260 2385 9300
rect 2425 9260 2435 9300
rect 2375 9240 2435 9260
rect 2375 9200 2385 9240
rect 2425 9200 2435 9240
rect 2375 9175 2435 9200
rect 2375 9135 2385 9175
rect 2425 9135 2435 9175
rect 2375 9105 2435 9135
rect 2375 9065 2385 9105
rect 2425 9065 2435 9105
rect 2375 9035 2435 9065
rect 2375 8995 2385 9035
rect 2425 8995 2435 9035
rect 2375 8965 2435 8995
rect 2375 8925 2385 8965
rect 2425 8925 2435 8965
rect 2375 8900 2435 8925
rect 2375 8860 2385 8900
rect 2425 8860 2435 8900
rect 2375 8840 2435 8860
rect 2375 8800 2385 8840
rect 2425 8800 2435 8840
rect 2375 8775 2435 8800
rect 2375 8735 2385 8775
rect 2425 8735 2435 8775
rect 2375 8705 2435 8735
rect 2375 8665 2385 8705
rect 2425 8665 2435 8705
rect 2375 8635 2435 8665
rect 2375 8595 2385 8635
rect 2425 8595 2435 8635
rect 2375 8565 2435 8595
rect 2375 8525 2385 8565
rect 2425 8525 2435 8565
rect 2375 8500 2435 8525
rect 2375 8460 2385 8500
rect 2425 8460 2435 8500
rect 2375 8440 2435 8460
rect 2375 8400 2385 8440
rect 2425 8400 2435 8440
rect 2375 8375 2435 8400
rect 2375 8335 2385 8375
rect 2425 8335 2435 8375
rect 2375 8305 2435 8335
rect 2375 8265 2385 8305
rect 2425 8265 2435 8305
rect 2375 8235 2435 8265
rect 2375 8195 2385 8235
rect 2425 8195 2435 8235
rect 2375 8165 2435 8195
rect 2375 8125 2385 8165
rect 2425 8125 2435 8165
rect 2375 8100 2435 8125
rect 2375 8060 2385 8100
rect 2425 8060 2435 8100
rect 2375 8040 2435 8060
rect 2375 8000 2385 8040
rect 2425 8000 2435 8040
rect 2375 7975 2435 8000
rect 2375 7935 2385 7975
rect 2425 7935 2435 7975
rect 2375 7905 2435 7935
rect 2375 7865 2385 7905
rect 2425 7865 2435 7905
rect 2375 7835 2435 7865
rect 2375 7795 2385 7835
rect 2425 7795 2435 7835
rect 2375 7765 2435 7795
rect 2375 7725 2385 7765
rect 2425 7725 2435 7765
rect 2375 7700 2435 7725
rect 2375 7660 2385 7700
rect 2425 7660 2435 7700
rect 2375 7640 2435 7660
rect 2375 7600 2385 7640
rect 2425 7600 2435 7640
rect 2375 7575 2435 7600
rect 2375 7535 2385 7575
rect 2425 7535 2435 7575
rect 2375 7505 2435 7535
rect 2375 7465 2385 7505
rect 2425 7465 2435 7505
rect 2375 7435 2435 7465
rect 2375 7395 2385 7435
rect 2425 7395 2435 7435
rect 2375 7365 2435 7395
rect 2375 7325 2385 7365
rect 2425 7325 2435 7365
rect 2375 7300 2435 7325
rect 2375 7260 2385 7300
rect 2425 7260 2435 7300
rect 2375 7240 2435 7260
rect 2375 7200 2385 7240
rect 2425 7200 2435 7240
rect 2375 7175 2435 7200
rect 2375 7135 2385 7175
rect 2425 7135 2435 7175
rect 2375 7105 2435 7135
rect 2375 7065 2385 7105
rect 2425 7065 2435 7105
rect 2375 7035 2435 7065
rect 2375 6995 2385 7035
rect 2425 6995 2435 7035
rect 2375 6965 2435 6995
rect 2375 6925 2385 6965
rect 2425 6925 2435 6965
rect 2375 6900 2435 6925
rect 2375 6860 2385 6900
rect 2425 6860 2435 6900
rect 2375 6840 2435 6860
rect 2375 6800 2385 6840
rect 2425 6800 2435 6840
rect 2375 6775 2435 6800
rect 2375 6735 2385 6775
rect 2425 6735 2435 6775
rect 2375 6705 2435 6735
rect 2375 6665 2385 6705
rect 2425 6665 2435 6705
rect 2375 6635 2435 6665
rect 2375 6595 2385 6635
rect 2425 6595 2435 6635
rect 2375 6565 2435 6595
rect 2375 6525 2385 6565
rect 2425 6525 2435 6565
rect 2375 6500 2435 6525
rect 2375 6460 2385 6500
rect 2425 6460 2435 6500
rect 2375 6450 2435 6460
rect 3225 9640 3285 9650
rect 3225 9600 3235 9640
rect 3275 9600 3285 9640
rect 3225 9575 3285 9600
rect 3225 9535 3235 9575
rect 3275 9535 3285 9575
rect 3225 9505 3285 9535
rect 3225 9465 3235 9505
rect 3275 9465 3285 9505
rect 3225 9435 3285 9465
rect 3225 9395 3235 9435
rect 3275 9395 3285 9435
rect 3225 9365 3285 9395
rect 3225 9325 3235 9365
rect 3275 9325 3285 9365
rect 3225 9300 3285 9325
rect 3225 9260 3235 9300
rect 3275 9260 3285 9300
rect 3225 9240 3285 9260
rect 3225 9200 3235 9240
rect 3275 9200 3285 9240
rect 3225 9175 3285 9200
rect 3225 9135 3235 9175
rect 3275 9135 3285 9175
rect 3225 9105 3285 9135
rect 3225 9065 3235 9105
rect 3275 9065 3285 9105
rect 3225 9035 3285 9065
rect 3225 8995 3235 9035
rect 3275 8995 3285 9035
rect 3225 8965 3285 8995
rect 3225 8925 3235 8965
rect 3275 8925 3285 8965
rect 3225 8900 3285 8925
rect 3225 8860 3235 8900
rect 3275 8860 3285 8900
rect 3225 8840 3285 8860
rect 3225 8800 3235 8840
rect 3275 8800 3285 8840
rect 3225 8775 3285 8800
rect 3225 8735 3235 8775
rect 3275 8735 3285 8775
rect 3225 8705 3285 8735
rect 3225 8665 3235 8705
rect 3275 8665 3285 8705
rect 3225 8635 3285 8665
rect 3225 8595 3235 8635
rect 3275 8595 3285 8635
rect 3225 8565 3285 8595
rect 3225 8525 3235 8565
rect 3275 8525 3285 8565
rect 3225 8500 3285 8525
rect 3225 8460 3235 8500
rect 3275 8460 3285 8500
rect 3225 8440 3285 8460
rect 3225 8400 3235 8440
rect 3275 8400 3285 8440
rect 3225 8375 3285 8400
rect 3225 8335 3235 8375
rect 3275 8335 3285 8375
rect 3225 8305 3285 8335
rect 3225 8265 3235 8305
rect 3275 8265 3285 8305
rect 3225 8235 3285 8265
rect 3225 8195 3235 8235
rect 3275 8195 3285 8235
rect 3225 8165 3285 8195
rect 3225 8125 3235 8165
rect 3275 8125 3285 8165
rect 3225 8100 3285 8125
rect 3225 8060 3235 8100
rect 3275 8060 3285 8100
rect 3225 8040 3285 8060
rect 3225 8000 3235 8040
rect 3275 8000 3285 8040
rect 3225 7975 3285 8000
rect 3225 7935 3235 7975
rect 3275 7935 3285 7975
rect 3225 7905 3285 7935
rect 3225 7865 3235 7905
rect 3275 7865 3285 7905
rect 3225 7835 3285 7865
rect 3225 7795 3235 7835
rect 3275 7795 3285 7835
rect 3225 7765 3285 7795
rect 3225 7725 3235 7765
rect 3275 7725 3285 7765
rect 3225 7700 3285 7725
rect 3225 7660 3235 7700
rect 3275 7660 3285 7700
rect 3225 7640 3285 7660
rect 3225 7600 3235 7640
rect 3275 7600 3285 7640
rect 3225 7575 3285 7600
rect 3225 7535 3235 7575
rect 3275 7535 3285 7575
rect 3225 7505 3285 7535
rect 3225 7465 3235 7505
rect 3275 7465 3285 7505
rect 3225 7435 3285 7465
rect 3225 7395 3235 7435
rect 3275 7395 3285 7435
rect 3225 7365 3285 7395
rect 3225 7325 3235 7365
rect 3275 7325 3285 7365
rect 3225 7300 3285 7325
rect 3225 7260 3235 7300
rect 3275 7260 3285 7300
rect 3225 7240 3285 7260
rect 3225 7200 3235 7240
rect 3275 7200 3285 7240
rect 3225 7175 3285 7200
rect 3225 7135 3235 7175
rect 3275 7135 3285 7175
rect 3225 7105 3285 7135
rect 3225 7065 3235 7105
rect 3275 7065 3285 7105
rect 3225 7035 3285 7065
rect 3225 6995 3235 7035
rect 3275 6995 3285 7035
rect 3225 6965 3285 6995
rect 3225 6925 3235 6965
rect 3275 6925 3285 6965
rect 3225 6900 3285 6925
rect 3225 6860 3235 6900
rect 3275 6860 3285 6900
rect 3225 6840 3285 6860
rect 3225 6800 3235 6840
rect 3275 6800 3285 6840
rect 3225 6775 3285 6800
rect 3225 6735 3235 6775
rect 3275 6735 3285 6775
rect 3225 6705 3285 6735
rect 3225 6665 3235 6705
rect 3275 6665 3285 6705
rect 3225 6635 3285 6665
rect 3225 6595 3235 6635
rect 3275 6595 3285 6635
rect 3225 6565 3285 6595
rect 3225 6525 3235 6565
rect 3275 6525 3285 6565
rect 3225 6500 3285 6525
rect 3225 6460 3235 6500
rect 3275 6460 3285 6500
rect 3225 6450 3285 6460
rect 5635 9640 5695 9650
rect 5635 9600 5645 9640
rect 5685 9600 5695 9640
rect 5635 9575 5695 9600
rect 5635 9535 5645 9575
rect 5685 9535 5695 9575
rect 5635 9505 5695 9535
rect 5635 9465 5645 9505
rect 5685 9465 5695 9505
rect 5635 9435 5695 9465
rect 5635 9395 5645 9435
rect 5685 9395 5695 9435
rect 5635 9365 5695 9395
rect 5635 9325 5645 9365
rect 5685 9325 5695 9365
rect 5635 9300 5695 9325
rect 5635 9260 5645 9300
rect 5685 9260 5695 9300
rect 5635 9240 5695 9260
rect 5635 9200 5645 9240
rect 5685 9200 5695 9240
rect 5635 9175 5695 9200
rect 5635 9135 5645 9175
rect 5685 9135 5695 9175
rect 5635 9105 5695 9135
rect 5635 9065 5645 9105
rect 5685 9065 5695 9105
rect 5635 9035 5695 9065
rect 5635 8995 5645 9035
rect 5685 8995 5695 9035
rect 5635 8965 5695 8995
rect 5635 8925 5645 8965
rect 5685 8925 5695 8965
rect 5635 8900 5695 8925
rect 5635 8860 5645 8900
rect 5685 8860 5695 8900
rect 5635 8840 5695 8860
rect 5635 8800 5645 8840
rect 5685 8800 5695 8840
rect 5635 8775 5695 8800
rect 5635 8735 5645 8775
rect 5685 8735 5695 8775
rect 5635 8705 5695 8735
rect 5635 8665 5645 8705
rect 5685 8665 5695 8705
rect 5635 8635 5695 8665
rect 5635 8595 5645 8635
rect 5685 8595 5695 8635
rect 5635 8565 5695 8595
rect 5635 8525 5645 8565
rect 5685 8525 5695 8565
rect 5635 8500 5695 8525
rect 5635 8460 5645 8500
rect 5685 8460 5695 8500
rect 5635 8440 5695 8460
rect 5635 8400 5645 8440
rect 5685 8400 5695 8440
rect 5635 8375 5695 8400
rect 5635 8335 5645 8375
rect 5685 8335 5695 8375
rect 5635 8305 5695 8335
rect 5635 8265 5645 8305
rect 5685 8265 5695 8305
rect 5635 8235 5695 8265
rect 5635 8195 5645 8235
rect 5685 8195 5695 8235
rect 5635 8165 5695 8195
rect 5635 8125 5645 8165
rect 5685 8125 5695 8165
rect 5635 8100 5695 8125
rect 5635 8060 5645 8100
rect 5685 8060 5695 8100
rect 5635 8040 5695 8060
rect 5635 8000 5645 8040
rect 5685 8000 5695 8040
rect 5635 7975 5695 8000
rect 5635 7935 5645 7975
rect 5685 7935 5695 7975
rect 5635 7905 5695 7935
rect 5635 7865 5645 7905
rect 5685 7865 5695 7905
rect 5635 7835 5695 7865
rect 5635 7795 5645 7835
rect 5685 7795 5695 7835
rect 5635 7765 5695 7795
rect 5635 7725 5645 7765
rect 5685 7725 5695 7765
rect 5635 7700 5695 7725
rect 5635 7660 5645 7700
rect 5685 7660 5695 7700
rect 5635 7640 5695 7660
rect 5635 7600 5645 7640
rect 5685 7600 5695 7640
rect 5635 7575 5695 7600
rect 5635 7535 5645 7575
rect 5685 7535 5695 7575
rect 5635 7505 5695 7535
rect 5635 7465 5645 7505
rect 5685 7465 5695 7505
rect 5635 7435 5695 7465
rect 5635 7395 5645 7435
rect 5685 7395 5695 7435
rect 5635 7365 5695 7395
rect 5635 7325 5645 7365
rect 5685 7325 5695 7365
rect 5635 7300 5695 7325
rect 5635 7260 5645 7300
rect 5685 7260 5695 7300
rect 5635 7240 5695 7260
rect 5635 7200 5645 7240
rect 5685 7200 5695 7240
rect 5635 7175 5695 7200
rect 5635 7135 5645 7175
rect 5685 7135 5695 7175
rect 5635 7105 5695 7135
rect 5635 7065 5645 7105
rect 5685 7065 5695 7105
rect 5635 7035 5695 7065
rect 5635 6995 5645 7035
rect 5685 6995 5695 7035
rect 5635 6965 5695 6995
rect 5635 6925 5645 6965
rect 5685 6925 5695 6965
rect 5635 6900 5695 6925
rect 5635 6860 5645 6900
rect 5685 6860 5695 6900
rect 5635 6840 5695 6860
rect 5635 6800 5645 6840
rect 5685 6800 5695 6840
rect 5635 6775 5695 6800
rect 5635 6735 5645 6775
rect 5685 6735 5695 6775
rect 5635 6705 5695 6735
rect 5635 6665 5645 6705
rect 5685 6665 5695 6705
rect 5635 6635 5695 6665
rect 5635 6595 5645 6635
rect 5685 6595 5695 6635
rect 5635 6565 5695 6595
rect 5635 6525 5645 6565
rect 5685 6525 5695 6565
rect 5635 6500 5695 6525
rect 5635 6460 5645 6500
rect 5685 6460 5695 6500
rect 5635 6450 5695 6460
rect 6290 9640 6350 9650
rect 6290 9600 6300 9640
rect 6340 9600 6350 9640
rect 6290 9575 6350 9600
rect 6290 9535 6300 9575
rect 6340 9535 6350 9575
rect 6290 9505 6350 9535
rect 6290 9465 6300 9505
rect 6340 9465 6350 9505
rect 6290 9435 6350 9465
rect 6290 9395 6300 9435
rect 6340 9395 6350 9435
rect 6290 9365 6350 9395
rect 6290 9325 6300 9365
rect 6340 9325 6350 9365
rect 6290 9300 6350 9325
rect 6290 9260 6300 9300
rect 6340 9260 6350 9300
rect 6290 9240 6350 9260
rect 6290 9200 6300 9240
rect 6340 9200 6350 9240
rect 6290 9175 6350 9200
rect 6290 9135 6300 9175
rect 6340 9135 6350 9175
rect 6290 9105 6350 9135
rect 6290 9065 6300 9105
rect 6340 9065 6350 9105
rect 6290 9035 6350 9065
rect 6290 8995 6300 9035
rect 6340 8995 6350 9035
rect 6290 8965 6350 8995
rect 6290 8925 6300 8965
rect 6340 8925 6350 8965
rect 6290 8900 6350 8925
rect 6290 8860 6300 8900
rect 6340 8860 6350 8900
rect 6290 8840 6350 8860
rect 6290 8800 6300 8840
rect 6340 8800 6350 8840
rect 6290 8775 6350 8800
rect 6290 8735 6300 8775
rect 6340 8735 6350 8775
rect 6290 8705 6350 8735
rect 6290 8665 6300 8705
rect 6340 8665 6350 8705
rect 6290 8635 6350 8665
rect 6290 8595 6300 8635
rect 6340 8595 6350 8635
rect 6290 8565 6350 8595
rect 6290 8525 6300 8565
rect 6340 8525 6350 8565
rect 6290 8500 6350 8525
rect 6290 8460 6300 8500
rect 6340 8460 6350 8500
rect 6290 8440 6350 8460
rect 6290 8400 6300 8440
rect 6340 8400 6350 8440
rect 6290 8375 6350 8400
rect 6290 8335 6300 8375
rect 6340 8335 6350 8375
rect 6290 8305 6350 8335
rect 6290 8265 6300 8305
rect 6340 8265 6350 8305
rect 6290 8235 6350 8265
rect 6290 8195 6300 8235
rect 6340 8195 6350 8235
rect 6290 8165 6350 8195
rect 6290 8125 6300 8165
rect 6340 8125 6350 8165
rect 6290 8100 6350 8125
rect 6290 8060 6300 8100
rect 6340 8060 6350 8100
rect 6290 8040 6350 8060
rect 6290 8000 6300 8040
rect 6340 8000 6350 8040
rect 6290 7975 6350 8000
rect 6290 7935 6300 7975
rect 6340 7935 6350 7975
rect 6290 7905 6350 7935
rect 6290 7865 6300 7905
rect 6340 7865 6350 7905
rect 6290 7835 6350 7865
rect 6290 7795 6300 7835
rect 6340 7795 6350 7835
rect 6290 7765 6350 7795
rect 6290 7725 6300 7765
rect 6340 7725 6350 7765
rect 6290 7700 6350 7725
rect 6290 7660 6300 7700
rect 6340 7660 6350 7700
rect 6290 7640 6350 7660
rect 6290 7600 6300 7640
rect 6340 7600 6350 7640
rect 6290 7575 6350 7600
rect 6290 7535 6300 7575
rect 6340 7535 6350 7575
rect 6290 7505 6350 7535
rect 6290 7465 6300 7505
rect 6340 7465 6350 7505
rect 6290 7435 6350 7465
rect 6290 7395 6300 7435
rect 6340 7395 6350 7435
rect 6290 7365 6350 7395
rect 6290 7325 6300 7365
rect 6340 7325 6350 7365
rect 6290 7300 6350 7325
rect 6290 7260 6300 7300
rect 6340 7260 6350 7300
rect 6290 7240 6350 7260
rect 6290 7200 6300 7240
rect 6340 7200 6350 7240
rect 6290 7175 6350 7200
rect 6290 7135 6300 7175
rect 6340 7135 6350 7175
rect 6290 7105 6350 7135
rect 6290 7065 6300 7105
rect 6340 7065 6350 7105
rect 6290 7035 6350 7065
rect 6290 6995 6300 7035
rect 6340 6995 6350 7035
rect 6290 6965 6350 6995
rect 6290 6925 6300 6965
rect 6340 6925 6350 6965
rect 6290 6900 6350 6925
rect 6290 6860 6300 6900
rect 6340 6860 6350 6900
rect 6290 6840 6350 6860
rect 6290 6800 6300 6840
rect 6340 6800 6350 6840
rect 6290 6775 6350 6800
rect 6290 6735 6300 6775
rect 6340 6735 6350 6775
rect 6290 6705 6350 6735
rect 6290 6665 6300 6705
rect 6340 6665 6350 6705
rect 6290 6635 6350 6665
rect 6290 6595 6300 6635
rect 6340 6595 6350 6635
rect 6290 6565 6350 6595
rect 6290 6525 6300 6565
rect 6340 6525 6350 6565
rect 6290 6500 6350 6525
rect 6290 6460 6300 6500
rect 6340 6460 6350 6500
rect 6290 6450 6350 6460
rect 6580 9640 6640 9650
rect 6580 9600 6590 9640
rect 6630 9600 6640 9640
rect 6580 9575 6640 9600
rect 6580 9535 6590 9575
rect 6630 9535 6640 9575
rect 6580 9505 6640 9535
rect 6580 9465 6590 9505
rect 6630 9465 6640 9505
rect 6580 9435 6640 9465
rect 6580 9395 6590 9435
rect 6630 9395 6640 9435
rect 6580 9365 6640 9395
rect 6580 9325 6590 9365
rect 6630 9325 6640 9365
rect 6580 9300 6640 9325
rect 6580 9260 6590 9300
rect 6630 9260 6640 9300
rect 6580 9240 6640 9260
rect 6580 9200 6590 9240
rect 6630 9200 6640 9240
rect 6580 9175 6640 9200
rect 6580 9135 6590 9175
rect 6630 9135 6640 9175
rect 6580 9105 6640 9135
rect 6580 9065 6590 9105
rect 6630 9065 6640 9105
rect 6580 9035 6640 9065
rect 6580 8995 6590 9035
rect 6630 8995 6640 9035
rect 6580 8965 6640 8995
rect 6580 8925 6590 8965
rect 6630 8925 6640 8965
rect 6580 8900 6640 8925
rect 6580 8860 6590 8900
rect 6630 8860 6640 8900
rect 6580 8840 6640 8860
rect 6580 8800 6590 8840
rect 6630 8800 6640 8840
rect 6580 8775 6640 8800
rect 6580 8735 6590 8775
rect 6630 8735 6640 8775
rect 6580 8705 6640 8735
rect 6580 8665 6590 8705
rect 6630 8665 6640 8705
rect 6580 8635 6640 8665
rect 6580 8595 6590 8635
rect 6630 8595 6640 8635
rect 6580 8565 6640 8595
rect 6580 8525 6590 8565
rect 6630 8525 6640 8565
rect 6580 8500 6640 8525
rect 6580 8460 6590 8500
rect 6630 8460 6640 8500
rect 6580 8440 6640 8460
rect 6580 8400 6590 8440
rect 6630 8400 6640 8440
rect 6580 8375 6640 8400
rect 6580 8335 6590 8375
rect 6630 8335 6640 8375
rect 6580 8305 6640 8335
rect 6580 8265 6590 8305
rect 6630 8265 6640 8305
rect 6580 8235 6640 8265
rect 6580 8195 6590 8235
rect 6630 8195 6640 8235
rect 6580 8165 6640 8195
rect 6580 8125 6590 8165
rect 6630 8125 6640 8165
rect 6580 8100 6640 8125
rect 6580 8060 6590 8100
rect 6630 8060 6640 8100
rect 6580 8040 6640 8060
rect 6580 8000 6590 8040
rect 6630 8000 6640 8040
rect 6580 7975 6640 8000
rect 6580 7935 6590 7975
rect 6630 7935 6640 7975
rect 6580 7905 6640 7935
rect 6580 7865 6590 7905
rect 6630 7865 6640 7905
rect 6580 7835 6640 7865
rect 6580 7795 6590 7835
rect 6630 7795 6640 7835
rect 6580 7765 6640 7795
rect 6580 7725 6590 7765
rect 6630 7725 6640 7765
rect 6580 7700 6640 7725
rect 6580 7660 6590 7700
rect 6630 7660 6640 7700
rect 6580 7640 6640 7660
rect 6580 7600 6590 7640
rect 6630 7600 6640 7640
rect 6580 7575 6640 7600
rect 6580 7535 6590 7575
rect 6630 7535 6640 7575
rect 6580 7505 6640 7535
rect 6580 7465 6590 7505
rect 6630 7465 6640 7505
rect 6580 7435 6640 7465
rect 6580 7395 6590 7435
rect 6630 7395 6640 7435
rect 6580 7365 6640 7395
rect 6580 7325 6590 7365
rect 6630 7325 6640 7365
rect 6580 7300 6640 7325
rect 6580 7260 6590 7300
rect 6630 7260 6640 7300
rect 6580 7240 6640 7260
rect 6580 7200 6590 7240
rect 6630 7200 6640 7240
rect 6580 7175 6640 7200
rect 6580 7135 6590 7175
rect 6630 7135 6640 7175
rect 6580 7105 6640 7135
rect 6580 7065 6590 7105
rect 6630 7065 6640 7105
rect 6580 7035 6640 7065
rect 6580 6995 6590 7035
rect 6630 6995 6640 7035
rect 6580 6965 6640 6995
rect 6580 6925 6590 6965
rect 6630 6925 6640 6965
rect 6580 6900 6640 6925
rect 6580 6860 6590 6900
rect 6630 6860 6640 6900
rect 6580 6840 6640 6860
rect 6580 6800 6590 6840
rect 6630 6800 6640 6840
rect 6580 6775 6640 6800
rect 6580 6735 6590 6775
rect 6630 6735 6640 6775
rect 6580 6705 6640 6735
rect 6580 6665 6590 6705
rect 6630 6665 6640 6705
rect 6580 6635 6640 6665
rect 6580 6595 6590 6635
rect 6630 6595 6640 6635
rect 6580 6565 6640 6595
rect 6580 6525 6590 6565
rect 6630 6525 6640 6565
rect 6580 6500 6640 6525
rect 6580 6460 6590 6500
rect 6630 6460 6640 6500
rect 6580 6450 6640 6460
rect 7260 9640 7320 9650
rect 7260 9600 7270 9640
rect 7310 9600 7320 9640
rect 7260 9575 7320 9600
rect 7260 9535 7270 9575
rect 7310 9535 7320 9575
rect 7260 9505 7320 9535
rect 7260 9465 7270 9505
rect 7310 9465 7320 9505
rect 7260 9435 7320 9465
rect 7260 9395 7270 9435
rect 7310 9395 7320 9435
rect 7260 9365 7320 9395
rect 7260 9325 7270 9365
rect 7310 9325 7320 9365
rect 7260 9300 7320 9325
rect 7260 9260 7270 9300
rect 7310 9260 7320 9300
rect 7260 9240 7320 9260
rect 7260 9200 7270 9240
rect 7310 9200 7320 9240
rect 7260 9175 7320 9200
rect 7260 9135 7270 9175
rect 7310 9135 7320 9175
rect 7260 9105 7320 9135
rect 7260 9065 7270 9105
rect 7310 9065 7320 9105
rect 7260 9035 7320 9065
rect 7260 8995 7270 9035
rect 7310 8995 7320 9035
rect 7260 8965 7320 8995
rect 7260 8925 7270 8965
rect 7310 8925 7320 8965
rect 7260 8900 7320 8925
rect 7260 8860 7270 8900
rect 7310 8860 7320 8900
rect 7260 8840 7320 8860
rect 7260 8800 7270 8840
rect 7310 8800 7320 8840
rect 7260 8775 7320 8800
rect 7260 8735 7270 8775
rect 7310 8735 7320 8775
rect 7260 8705 7320 8735
rect 7260 8665 7270 8705
rect 7310 8665 7320 8705
rect 7260 8635 7320 8665
rect 7260 8595 7270 8635
rect 7310 8595 7320 8635
rect 7260 8565 7320 8595
rect 7260 8525 7270 8565
rect 7310 8525 7320 8565
rect 7260 8500 7320 8525
rect 7260 8460 7270 8500
rect 7310 8460 7320 8500
rect 7260 8440 7320 8460
rect 7260 8400 7270 8440
rect 7310 8400 7320 8440
rect 7260 8375 7320 8400
rect 7260 8335 7270 8375
rect 7310 8335 7320 8375
rect 7260 8305 7320 8335
rect 7260 8265 7270 8305
rect 7310 8265 7320 8305
rect 7260 8235 7320 8265
rect 7260 8195 7270 8235
rect 7310 8195 7320 8235
rect 7260 8165 7320 8195
rect 7260 8125 7270 8165
rect 7310 8125 7320 8165
rect 7260 8100 7320 8125
rect 7260 8060 7270 8100
rect 7310 8060 7320 8100
rect 7260 8040 7320 8060
rect 7260 8000 7270 8040
rect 7310 8000 7320 8040
rect 7260 7975 7320 8000
rect 7260 7935 7270 7975
rect 7310 7935 7320 7975
rect 7260 7905 7320 7935
rect 7260 7865 7270 7905
rect 7310 7865 7320 7905
rect 7260 7835 7320 7865
rect 7260 7795 7270 7835
rect 7310 7795 7320 7835
rect 7260 7765 7320 7795
rect 7260 7725 7270 7765
rect 7310 7725 7320 7765
rect 7260 7700 7320 7725
rect 7260 7660 7270 7700
rect 7310 7660 7320 7700
rect 7260 7640 7320 7660
rect 7260 7600 7270 7640
rect 7310 7600 7320 7640
rect 7260 7575 7320 7600
rect 7260 7535 7270 7575
rect 7310 7535 7320 7575
rect 7260 7505 7320 7535
rect 7260 7465 7270 7505
rect 7310 7465 7320 7505
rect 7260 7435 7320 7465
rect 7260 7395 7270 7435
rect 7310 7395 7320 7435
rect 7260 7365 7320 7395
rect 7260 7325 7270 7365
rect 7310 7325 7320 7365
rect 7260 7300 7320 7325
rect 7260 7260 7270 7300
rect 7310 7260 7320 7300
rect 7260 7240 7320 7260
rect 7260 7200 7270 7240
rect 7310 7200 7320 7240
rect 7260 7175 7320 7200
rect 7260 7135 7270 7175
rect 7310 7135 7320 7175
rect 7260 7105 7320 7135
rect 7260 7065 7270 7105
rect 7310 7065 7320 7105
rect 7260 7035 7320 7065
rect 7260 6995 7270 7035
rect 7310 6995 7320 7035
rect 7260 6965 7320 6995
rect 7260 6925 7270 6965
rect 7310 6925 7320 6965
rect 7260 6900 7320 6925
rect 7260 6860 7270 6900
rect 7310 6860 7320 6900
rect 7260 6840 7320 6860
rect 7260 6800 7270 6840
rect 7310 6800 7320 6840
rect 7260 6775 7320 6800
rect 7260 6735 7270 6775
rect 7310 6735 7320 6775
rect 7260 6705 7320 6735
rect 7260 6665 7270 6705
rect 7310 6665 7320 6705
rect 7260 6635 7320 6665
rect 7260 6595 7270 6635
rect 7310 6595 7320 6635
rect 7260 6565 7320 6595
rect 7260 6525 7270 6565
rect 7310 6525 7320 6565
rect 7260 6500 7320 6525
rect 7260 6460 7270 6500
rect 7310 6460 7320 6500
rect 7260 6450 7320 6460
rect 7610 9640 7670 9650
rect 7610 9600 7620 9640
rect 7660 9600 7670 9640
rect 7610 9575 7670 9600
rect 7610 9535 7620 9575
rect 7660 9535 7670 9575
rect 7610 9505 7670 9535
rect 7610 9465 7620 9505
rect 7660 9465 7670 9505
rect 7610 9435 7670 9465
rect 7610 9395 7620 9435
rect 7660 9395 7670 9435
rect 7610 9365 7670 9395
rect 7610 9325 7620 9365
rect 7660 9325 7670 9365
rect 7610 9300 7670 9325
rect 7610 9260 7620 9300
rect 7660 9260 7670 9300
rect 7610 9240 7670 9260
rect 7610 9200 7620 9240
rect 7660 9200 7670 9240
rect 7610 9175 7670 9200
rect 7610 9135 7620 9175
rect 7660 9135 7670 9175
rect 7610 9105 7670 9135
rect 7610 9065 7620 9105
rect 7660 9065 7670 9105
rect 7610 9035 7670 9065
rect 7610 8995 7620 9035
rect 7660 8995 7670 9035
rect 7610 8965 7670 8995
rect 7610 8925 7620 8965
rect 7660 8925 7670 8965
rect 7610 8900 7670 8925
rect 7610 8860 7620 8900
rect 7660 8860 7670 8900
rect 7610 8840 7670 8860
rect 7610 8800 7620 8840
rect 7660 8800 7670 8840
rect 7610 8775 7670 8800
rect 7610 8735 7620 8775
rect 7660 8735 7670 8775
rect 7610 8705 7670 8735
rect 7610 8665 7620 8705
rect 7660 8665 7670 8705
rect 7610 8635 7670 8665
rect 7610 8595 7620 8635
rect 7660 8595 7670 8635
rect 7610 8565 7670 8595
rect 7610 8525 7620 8565
rect 7660 8525 7670 8565
rect 7610 8500 7670 8525
rect 7610 8460 7620 8500
rect 7660 8460 7670 8500
rect 7610 8440 7670 8460
rect 7610 8400 7620 8440
rect 7660 8400 7670 8440
rect 7610 8375 7670 8400
rect 7610 8335 7620 8375
rect 7660 8335 7670 8375
rect 7610 8305 7670 8335
rect 7610 8265 7620 8305
rect 7660 8265 7670 8305
rect 7610 8235 7670 8265
rect 7610 8195 7620 8235
rect 7660 8195 7670 8235
rect 7610 8165 7670 8195
rect 7610 8125 7620 8165
rect 7660 8125 7670 8165
rect 7610 8100 7670 8125
rect 7610 8060 7620 8100
rect 7660 8060 7670 8100
rect 7610 8040 7670 8060
rect 7610 8000 7620 8040
rect 7660 8000 7670 8040
rect 7610 7975 7670 8000
rect 7610 7935 7620 7975
rect 7660 7935 7670 7975
rect 7610 7905 7670 7935
rect 7610 7865 7620 7905
rect 7660 7865 7670 7905
rect 7610 7835 7670 7865
rect 7610 7795 7620 7835
rect 7660 7795 7670 7835
rect 7610 7765 7670 7795
rect 7610 7725 7620 7765
rect 7660 7725 7670 7765
rect 7610 7700 7670 7725
rect 7610 7660 7620 7700
rect 7660 7660 7670 7700
rect 7610 7640 7670 7660
rect 7610 7600 7620 7640
rect 7660 7600 7670 7640
rect 7610 7575 7670 7600
rect 7610 7535 7620 7575
rect 7660 7535 7670 7575
rect 7610 7505 7670 7535
rect 7610 7465 7620 7505
rect 7660 7465 7670 7505
rect 7610 7435 7670 7465
rect 7610 7395 7620 7435
rect 7660 7395 7670 7435
rect 7610 7365 7670 7395
rect 7610 7325 7620 7365
rect 7660 7325 7670 7365
rect 7610 7300 7670 7325
rect 7610 7260 7620 7300
rect 7660 7260 7670 7300
rect 7610 7240 7670 7260
rect 7610 7200 7620 7240
rect 7660 7200 7670 7240
rect 7610 7175 7670 7200
rect 7610 7135 7620 7175
rect 7660 7135 7670 7175
rect 7610 7105 7670 7135
rect 7610 7065 7620 7105
rect 7660 7065 7670 7105
rect 7610 7035 7670 7065
rect 7610 6995 7620 7035
rect 7660 6995 7670 7035
rect 7610 6965 7670 6995
rect 7610 6925 7620 6965
rect 7660 6925 7670 6965
rect 7610 6900 7670 6925
rect 7610 6860 7620 6900
rect 7660 6860 7670 6900
rect 7610 6840 7670 6860
rect 7610 6800 7620 6840
rect 7660 6800 7670 6840
rect 7610 6775 7670 6800
rect 7610 6735 7620 6775
rect 7660 6735 7670 6775
rect 7610 6705 7670 6735
rect 7610 6665 7620 6705
rect 7660 6665 7670 6705
rect 7610 6635 7670 6665
rect 7610 6595 7620 6635
rect 7660 6595 7670 6635
rect 7610 6565 7670 6595
rect 7610 6525 7620 6565
rect 7660 6525 7670 6565
rect 7610 6500 7670 6525
rect 7610 6460 7620 6500
rect 7660 6460 7670 6500
rect 7610 6450 7670 6460
rect 8310 9640 8370 9650
rect 8310 9600 8320 9640
rect 8360 9600 8370 9640
rect 8310 9575 8370 9600
rect 8310 9535 8320 9575
rect 8360 9535 8370 9575
rect 8310 9505 8370 9535
rect 8310 9465 8320 9505
rect 8360 9465 8370 9505
rect 8310 9435 8370 9465
rect 8310 9395 8320 9435
rect 8360 9395 8370 9435
rect 8310 9365 8370 9395
rect 8310 9325 8320 9365
rect 8360 9325 8370 9365
rect 8310 9300 8370 9325
rect 8310 9260 8320 9300
rect 8360 9260 8370 9300
rect 8310 9240 8370 9260
rect 8310 9200 8320 9240
rect 8360 9200 8370 9240
rect 8310 9175 8370 9200
rect 8310 9135 8320 9175
rect 8360 9135 8370 9175
rect 8310 9105 8370 9135
rect 8310 9065 8320 9105
rect 8360 9065 8370 9105
rect 8310 9035 8370 9065
rect 8310 8995 8320 9035
rect 8360 8995 8370 9035
rect 8310 8965 8370 8995
rect 8310 8925 8320 8965
rect 8360 8925 8370 8965
rect 8310 8900 8370 8925
rect 8310 8860 8320 8900
rect 8360 8860 8370 8900
rect 8310 8840 8370 8860
rect 8310 8800 8320 8840
rect 8360 8800 8370 8840
rect 8310 8775 8370 8800
rect 8310 8735 8320 8775
rect 8360 8735 8370 8775
rect 8310 8705 8370 8735
rect 8310 8665 8320 8705
rect 8360 8665 8370 8705
rect 8310 8635 8370 8665
rect 8310 8595 8320 8635
rect 8360 8595 8370 8635
rect 8310 8565 8370 8595
rect 8310 8525 8320 8565
rect 8360 8525 8370 8565
rect 8310 8500 8370 8525
rect 8310 8460 8320 8500
rect 8360 8460 8370 8500
rect 8310 8440 8370 8460
rect 8310 8400 8320 8440
rect 8360 8400 8370 8440
rect 8310 8375 8370 8400
rect 8310 8335 8320 8375
rect 8360 8335 8370 8375
rect 8310 8305 8370 8335
rect 8310 8265 8320 8305
rect 8360 8265 8370 8305
rect 8310 8235 8370 8265
rect 8310 8195 8320 8235
rect 8360 8195 8370 8235
rect 8310 8165 8370 8195
rect 8310 8125 8320 8165
rect 8360 8125 8370 8165
rect 8310 8100 8370 8125
rect 8310 8060 8320 8100
rect 8360 8060 8370 8100
rect 8310 8040 8370 8060
rect 8310 8000 8320 8040
rect 8360 8000 8370 8040
rect 8310 7975 8370 8000
rect 8310 7935 8320 7975
rect 8360 7935 8370 7975
rect 8310 7905 8370 7935
rect 8310 7865 8320 7905
rect 8360 7865 8370 7905
rect 8310 7835 8370 7865
rect 8310 7795 8320 7835
rect 8360 7795 8370 7835
rect 8310 7765 8370 7795
rect 8310 7725 8320 7765
rect 8360 7725 8370 7765
rect 8310 7700 8370 7725
rect 8310 7660 8320 7700
rect 8360 7660 8370 7700
rect 8310 7640 8370 7660
rect 8310 7600 8320 7640
rect 8360 7600 8370 7640
rect 8310 7575 8370 7600
rect 8310 7535 8320 7575
rect 8360 7535 8370 7575
rect 8310 7505 8370 7535
rect 8310 7465 8320 7505
rect 8360 7465 8370 7505
rect 8310 7435 8370 7465
rect 8310 7395 8320 7435
rect 8360 7395 8370 7435
rect 8310 7365 8370 7395
rect 8310 7325 8320 7365
rect 8360 7325 8370 7365
rect 8310 7300 8370 7325
rect 8310 7260 8320 7300
rect 8360 7260 8370 7300
rect 8310 7240 8370 7260
rect 8310 7200 8320 7240
rect 8360 7200 8370 7240
rect 8310 7175 8370 7200
rect 8310 7135 8320 7175
rect 8360 7135 8370 7175
rect 8310 7105 8370 7135
rect 8310 7065 8320 7105
rect 8360 7065 8370 7105
rect 8310 7035 8370 7065
rect 8310 6995 8320 7035
rect 8360 6995 8370 7035
rect 8310 6965 8370 6995
rect 8310 6925 8320 6965
rect 8360 6925 8370 6965
rect 8310 6900 8370 6925
rect 8310 6860 8320 6900
rect 8360 6860 8370 6900
rect 8310 6840 8370 6860
rect 8310 6800 8320 6840
rect 8360 6800 8370 6840
rect 8310 6775 8370 6800
rect 8310 6735 8320 6775
rect 8360 6735 8370 6775
rect 8310 6705 8370 6735
rect 8310 6665 8320 6705
rect 8360 6665 8370 6705
rect 8310 6635 8370 6665
rect 8310 6595 8320 6635
rect 8360 6595 8370 6635
rect 8310 6565 8370 6595
rect 8310 6525 8320 6565
rect 8360 6525 8370 6565
rect 8310 6500 8370 6525
rect 8310 6460 8320 6500
rect 8360 6460 8370 6500
rect 8310 6450 8370 6460
rect 8660 9640 8720 9650
rect 8660 9600 8670 9640
rect 8710 9600 8720 9640
rect 8660 9575 8720 9600
rect 8660 9535 8670 9575
rect 8710 9535 8720 9575
rect 8660 9505 8720 9535
rect 8660 9465 8670 9505
rect 8710 9465 8720 9505
rect 8660 9435 8720 9465
rect 8660 9395 8670 9435
rect 8710 9395 8720 9435
rect 8660 9365 8720 9395
rect 8660 9325 8670 9365
rect 8710 9325 8720 9365
rect 8660 9300 8720 9325
rect 8660 9260 8670 9300
rect 8710 9260 8720 9300
rect 8660 9240 8720 9260
rect 8660 9200 8670 9240
rect 8710 9200 8720 9240
rect 8660 9175 8720 9200
rect 8660 9135 8670 9175
rect 8710 9135 8720 9175
rect 8660 9105 8720 9135
rect 8660 9065 8670 9105
rect 8710 9065 8720 9105
rect 8660 9035 8720 9065
rect 8660 8995 8670 9035
rect 8710 8995 8720 9035
rect 8660 8965 8720 8995
rect 8660 8925 8670 8965
rect 8710 8925 8720 8965
rect 8660 8900 8720 8925
rect 8660 8860 8670 8900
rect 8710 8860 8720 8900
rect 8660 8840 8720 8860
rect 8660 8800 8670 8840
rect 8710 8800 8720 8840
rect 8660 8775 8720 8800
rect 8660 8735 8670 8775
rect 8710 8735 8720 8775
rect 8660 8705 8720 8735
rect 8660 8665 8670 8705
rect 8710 8665 8720 8705
rect 8660 8635 8720 8665
rect 8660 8595 8670 8635
rect 8710 8595 8720 8635
rect 8660 8565 8720 8595
rect 8660 8525 8670 8565
rect 8710 8525 8720 8565
rect 8660 8500 8720 8525
rect 8660 8460 8670 8500
rect 8710 8460 8720 8500
rect 8660 8440 8720 8460
rect 8660 8400 8670 8440
rect 8710 8400 8720 8440
rect 8660 8375 8720 8400
rect 8660 8335 8670 8375
rect 8710 8335 8720 8375
rect 8660 8305 8720 8335
rect 8660 8265 8670 8305
rect 8710 8265 8720 8305
rect 8660 8235 8720 8265
rect 8660 8195 8670 8235
rect 8710 8195 8720 8235
rect 8660 8165 8720 8195
rect 8660 8125 8670 8165
rect 8710 8125 8720 8165
rect 8660 8100 8720 8125
rect 8660 8060 8670 8100
rect 8710 8060 8720 8100
rect 8660 8040 8720 8060
rect 8660 8000 8670 8040
rect 8710 8000 8720 8040
rect 8660 7975 8720 8000
rect 8660 7935 8670 7975
rect 8710 7935 8720 7975
rect 8660 7905 8720 7935
rect 8660 7865 8670 7905
rect 8710 7865 8720 7905
rect 8660 7835 8720 7865
rect 8660 7795 8670 7835
rect 8710 7795 8720 7835
rect 8660 7765 8720 7795
rect 8660 7725 8670 7765
rect 8710 7725 8720 7765
rect 8660 7700 8720 7725
rect 8660 7660 8670 7700
rect 8710 7660 8720 7700
rect 8660 7640 8720 7660
rect 8660 7600 8670 7640
rect 8710 7600 8720 7640
rect 8660 7575 8720 7600
rect 8660 7535 8670 7575
rect 8710 7535 8720 7575
rect 8660 7505 8720 7535
rect 8660 7465 8670 7505
rect 8710 7465 8720 7505
rect 8660 7435 8720 7465
rect 8660 7395 8670 7435
rect 8710 7395 8720 7435
rect 8660 7365 8720 7395
rect 8660 7325 8670 7365
rect 8710 7325 8720 7365
rect 8660 7300 8720 7325
rect 8660 7260 8670 7300
rect 8710 7260 8720 7300
rect 8660 7240 8720 7260
rect 8660 7200 8670 7240
rect 8710 7200 8720 7240
rect 8660 7175 8720 7200
rect 8660 7135 8670 7175
rect 8710 7135 8720 7175
rect 8660 7105 8720 7135
rect 8660 7065 8670 7105
rect 8710 7065 8720 7105
rect 8660 7035 8720 7065
rect 8660 6995 8670 7035
rect 8710 6995 8720 7035
rect 8660 6965 8720 6995
rect 8660 6925 8670 6965
rect 8710 6925 8720 6965
rect 8660 6900 8720 6925
rect 8660 6860 8670 6900
rect 8710 6860 8720 6900
rect 8660 6840 8720 6860
rect 8660 6800 8670 6840
rect 8710 6800 8720 6840
rect 8660 6775 8720 6800
rect 8660 6735 8670 6775
rect 8710 6735 8720 6775
rect 8660 6705 8720 6735
rect 8660 6665 8670 6705
rect 8710 6665 8720 6705
rect 8660 6635 8720 6665
rect 8660 6595 8670 6635
rect 8710 6595 8720 6635
rect 8660 6565 8720 6595
rect 8660 6525 8670 6565
rect 8710 6525 8720 6565
rect 8660 6500 8720 6525
rect 8660 6460 8670 6500
rect 8710 6460 8720 6500
rect 8660 6450 8720 6460
rect 9010 9640 9070 9650
rect 9010 9600 9020 9640
rect 9060 9600 9070 9640
rect 9540 9600 9770 9695
rect 9890 9600 10120 9695
rect 10240 9600 10470 9695
rect 10590 9600 10820 9695
rect 10940 9600 11170 9695
rect 11290 9600 11520 9695
rect 11640 9600 11870 9695
rect 11990 9600 12220 9695
rect 12340 9600 12570 9695
rect 12690 9600 12920 9695
rect 13040 9600 13270 9695
rect 13390 9600 13620 9695
rect 13740 9600 13970 9695
rect 14090 9600 14320 9695
rect 14440 9600 14670 9695
rect 14790 9615 17990 17395
rect 9010 9575 9070 9600
rect 9010 9535 9020 9575
rect 9060 9535 9070 9575
rect 9010 9505 9070 9535
rect 9010 9465 9020 9505
rect 9060 9465 9070 9505
rect 12080 9480 12130 9600
rect 14790 9565 14825 9615
rect 14875 9565 14920 9615
rect 14970 9565 15015 9615
rect 15065 9565 15115 9615
rect 15165 9565 15215 9615
rect 15265 9565 15315 9615
rect 15365 9565 15410 9615
rect 15460 9565 15505 9615
rect 15555 9565 15625 9615
rect 15675 9565 15720 9615
rect 15770 9565 15815 9615
rect 15865 9565 15915 9615
rect 15965 9565 16015 9615
rect 16065 9565 16115 9615
rect 16165 9565 16210 9615
rect 16260 9565 16305 9615
rect 16355 9565 16425 9615
rect 16475 9565 16520 9615
rect 16570 9565 16615 9615
rect 16665 9565 16715 9615
rect 16765 9565 16815 9615
rect 16865 9565 16915 9615
rect 16965 9565 17010 9615
rect 17060 9565 17105 9615
rect 17155 9565 17225 9615
rect 17275 9565 17320 9615
rect 17370 9565 17415 9615
rect 17465 9565 17515 9615
rect 17565 9565 17615 9615
rect 17665 9565 17715 9615
rect 17765 9565 17810 9615
rect 17860 9565 17905 9615
rect 17955 9565 17990 9615
rect 14790 9525 17990 9565
rect 9010 9435 9070 9465
rect 9010 9395 9020 9435
rect 9060 9395 9070 9435
rect 9010 9365 9070 9395
rect 9010 9325 9020 9365
rect 9060 9325 9070 9365
rect 9010 9300 9070 9325
rect 9010 9260 9020 9300
rect 9060 9260 9070 9300
rect 9010 9240 9070 9260
rect 9540 9395 9770 9480
rect 9890 9395 10120 9480
rect 10240 9395 10470 9480
rect 10590 9395 10820 9480
rect 10940 9395 11170 9480
rect 11290 9395 11520 9480
rect 11640 9395 11870 9480
rect 11990 9395 12220 9480
rect 12340 9395 12570 9480
rect 12690 9395 12920 9480
rect 13040 9395 13270 9480
rect 13390 9395 13620 9480
rect 13740 9395 13970 9480
rect 14090 9395 14320 9480
rect 14440 9395 14670 9480
rect 9540 9345 14670 9395
rect 9540 9250 9770 9345
rect 9890 9250 10120 9345
rect 10240 9250 10470 9345
rect 10590 9250 10820 9345
rect 10940 9250 11170 9345
rect 11290 9250 11520 9345
rect 11640 9250 11870 9345
rect 11990 9250 12220 9345
rect 12340 9250 12570 9345
rect 12690 9250 12920 9345
rect 13040 9250 13270 9345
rect 13390 9250 13620 9345
rect 13740 9250 13970 9345
rect 14090 9250 14320 9345
rect 14440 9250 14670 9345
rect 14790 9475 14825 9525
rect 14875 9475 14920 9525
rect 14970 9475 15015 9525
rect 15065 9475 15115 9525
rect 15165 9475 15215 9525
rect 15265 9475 15315 9525
rect 15365 9475 15410 9525
rect 15460 9475 15505 9525
rect 15555 9475 15625 9525
rect 15675 9475 15720 9525
rect 15770 9475 15815 9525
rect 15865 9475 15915 9525
rect 15965 9475 16015 9525
rect 16065 9475 16115 9525
rect 16165 9475 16210 9525
rect 16260 9475 16305 9525
rect 16355 9475 16425 9525
rect 16475 9475 16520 9525
rect 16570 9475 16615 9525
rect 16665 9475 16715 9525
rect 16765 9475 16815 9525
rect 16865 9475 16915 9525
rect 16965 9475 17010 9525
rect 17060 9475 17105 9525
rect 17155 9475 17225 9525
rect 17275 9475 17320 9525
rect 17370 9475 17415 9525
rect 17465 9475 17515 9525
rect 17565 9475 17615 9525
rect 17665 9475 17715 9525
rect 17765 9475 17810 9525
rect 17860 9475 17905 9525
rect 17955 9475 17990 9525
rect 14790 9425 17990 9475
rect 14790 9375 14825 9425
rect 14875 9375 14920 9425
rect 14970 9375 15015 9425
rect 15065 9375 15115 9425
rect 15165 9375 15215 9425
rect 15265 9375 15315 9425
rect 15365 9375 15410 9425
rect 15460 9375 15505 9425
rect 15555 9375 15625 9425
rect 15675 9375 15720 9425
rect 15770 9375 15815 9425
rect 15865 9375 15915 9425
rect 15965 9375 16015 9425
rect 16065 9375 16115 9425
rect 16165 9375 16210 9425
rect 16260 9375 16305 9425
rect 16355 9375 16425 9425
rect 16475 9375 16520 9425
rect 16570 9375 16615 9425
rect 16665 9375 16715 9425
rect 16765 9375 16815 9425
rect 16865 9375 16915 9425
rect 16965 9375 17010 9425
rect 17060 9375 17105 9425
rect 17155 9375 17225 9425
rect 17275 9375 17320 9425
rect 17370 9375 17415 9425
rect 17465 9375 17515 9425
rect 17565 9375 17615 9425
rect 17665 9375 17715 9425
rect 17765 9375 17810 9425
rect 17860 9375 17905 9425
rect 17955 9375 17990 9425
rect 14790 9335 17990 9375
rect 14790 9285 14825 9335
rect 14875 9285 14920 9335
rect 14970 9285 15015 9335
rect 15065 9285 15115 9335
rect 15165 9285 15215 9335
rect 15265 9285 15315 9335
rect 15365 9285 15410 9335
rect 15460 9285 15505 9335
rect 15555 9285 15625 9335
rect 15675 9285 15720 9335
rect 15770 9285 15815 9335
rect 15865 9285 15915 9335
rect 15965 9285 16015 9335
rect 16065 9285 16115 9335
rect 16165 9285 16210 9335
rect 16260 9285 16305 9335
rect 16355 9285 16425 9335
rect 16475 9285 16520 9335
rect 16570 9285 16615 9335
rect 16665 9285 16715 9335
rect 16765 9285 16815 9335
rect 16865 9285 16915 9335
rect 16965 9285 17010 9335
rect 17060 9285 17105 9335
rect 17155 9285 17225 9335
rect 17275 9285 17320 9335
rect 17370 9285 17415 9335
rect 17465 9285 17515 9335
rect 17565 9285 17615 9335
rect 17665 9285 17715 9335
rect 17765 9285 17810 9335
rect 17860 9285 17905 9335
rect 17955 9285 17990 9335
rect 9010 9200 9020 9240
rect 9060 9200 9070 9240
rect 9010 9175 9070 9200
rect 9010 9135 9020 9175
rect 9060 9135 9070 9175
rect 9010 9105 9070 9135
rect 12080 9130 12130 9250
rect 14790 9215 17990 9285
rect 14790 9165 14825 9215
rect 14875 9165 14920 9215
rect 14970 9165 15015 9215
rect 15065 9165 15115 9215
rect 15165 9165 15215 9215
rect 15265 9165 15315 9215
rect 15365 9165 15410 9215
rect 15460 9165 15505 9215
rect 15555 9165 15625 9215
rect 15675 9165 15720 9215
rect 15770 9165 15815 9215
rect 15865 9165 15915 9215
rect 15965 9165 16015 9215
rect 16065 9165 16115 9215
rect 16165 9165 16210 9215
rect 16260 9165 16305 9215
rect 16355 9165 16425 9215
rect 16475 9165 16520 9215
rect 16570 9165 16615 9215
rect 16665 9165 16715 9215
rect 16765 9165 16815 9215
rect 16865 9165 16915 9215
rect 16965 9165 17010 9215
rect 17060 9165 17105 9215
rect 17155 9165 17225 9215
rect 17275 9165 17320 9215
rect 17370 9165 17415 9215
rect 17465 9165 17515 9215
rect 17565 9165 17615 9215
rect 17665 9165 17715 9215
rect 17765 9165 17810 9215
rect 17860 9165 17905 9215
rect 17955 9165 17990 9215
rect 9010 9065 9020 9105
rect 9060 9065 9070 9105
rect 9010 9035 9070 9065
rect 9010 8995 9020 9035
rect 9060 8995 9070 9035
rect 9010 8965 9070 8995
rect 9010 8925 9020 8965
rect 9060 8925 9070 8965
rect 9010 8900 9070 8925
rect 9540 9045 9770 9130
rect 9890 9045 10120 9130
rect 10240 9045 10470 9130
rect 10590 9045 10820 9130
rect 10940 9045 11170 9130
rect 11290 9045 11520 9130
rect 11640 9045 11870 9130
rect 11990 9045 12220 9130
rect 12340 9045 12570 9130
rect 12690 9045 12920 9130
rect 13040 9045 13270 9130
rect 13390 9045 13620 9130
rect 13740 9045 13970 9130
rect 14090 9045 14320 9130
rect 14440 9045 14670 9130
rect 9540 8995 14670 9045
rect 9540 8900 9770 8995
rect 9890 8900 10120 8995
rect 10240 8900 10470 8995
rect 10590 8900 10820 8995
rect 10940 8900 11170 8995
rect 11290 8900 11520 8995
rect 11640 8900 11870 8995
rect 11990 8900 12220 8995
rect 12340 8900 12570 8995
rect 12690 8900 12920 8995
rect 13040 8900 13270 8995
rect 13390 8900 13620 8995
rect 13740 8900 13970 8995
rect 14090 8900 14320 8995
rect 14440 8900 14670 8995
rect 14790 9125 17990 9165
rect 14790 9075 14825 9125
rect 14875 9075 14920 9125
rect 14970 9075 15015 9125
rect 15065 9075 15115 9125
rect 15165 9075 15215 9125
rect 15265 9075 15315 9125
rect 15365 9075 15410 9125
rect 15460 9075 15505 9125
rect 15555 9075 15625 9125
rect 15675 9075 15720 9125
rect 15770 9075 15815 9125
rect 15865 9075 15915 9125
rect 15965 9075 16015 9125
rect 16065 9075 16115 9125
rect 16165 9075 16210 9125
rect 16260 9075 16305 9125
rect 16355 9075 16425 9125
rect 16475 9075 16520 9125
rect 16570 9075 16615 9125
rect 16665 9075 16715 9125
rect 16765 9075 16815 9125
rect 16865 9075 16915 9125
rect 16965 9075 17010 9125
rect 17060 9075 17105 9125
rect 17155 9075 17225 9125
rect 17275 9075 17320 9125
rect 17370 9075 17415 9125
rect 17465 9075 17515 9125
rect 17565 9075 17615 9125
rect 17665 9075 17715 9125
rect 17765 9075 17810 9125
rect 17860 9075 17905 9125
rect 17955 9075 17990 9125
rect 14790 9025 17990 9075
rect 14790 8975 14825 9025
rect 14875 8975 14920 9025
rect 14970 8975 15015 9025
rect 15065 8975 15115 9025
rect 15165 8975 15215 9025
rect 15265 8975 15315 9025
rect 15365 8975 15410 9025
rect 15460 8975 15505 9025
rect 15555 8975 15625 9025
rect 15675 8975 15720 9025
rect 15770 8975 15815 9025
rect 15865 8975 15915 9025
rect 15965 8975 16015 9025
rect 16065 8975 16115 9025
rect 16165 8975 16210 9025
rect 16260 8975 16305 9025
rect 16355 8975 16425 9025
rect 16475 8975 16520 9025
rect 16570 8975 16615 9025
rect 16665 8975 16715 9025
rect 16765 8975 16815 9025
rect 16865 8975 16915 9025
rect 16965 8975 17010 9025
rect 17060 8975 17105 9025
rect 17155 8975 17225 9025
rect 17275 8975 17320 9025
rect 17370 8975 17415 9025
rect 17465 8975 17515 9025
rect 17565 8975 17615 9025
rect 17665 8975 17715 9025
rect 17765 8975 17810 9025
rect 17860 8975 17905 9025
rect 17955 8975 17990 9025
rect 14790 8935 17990 8975
rect 9010 8860 9020 8900
rect 9060 8860 9070 8900
rect 9010 8840 9070 8860
rect 9010 8800 9020 8840
rect 9060 8800 9070 8840
rect 9010 8775 9070 8800
rect 12080 8780 12130 8900
rect 14790 8885 14825 8935
rect 14875 8885 14920 8935
rect 14970 8885 15015 8935
rect 15065 8885 15115 8935
rect 15165 8885 15215 8935
rect 15265 8885 15315 8935
rect 15365 8885 15410 8935
rect 15460 8885 15505 8935
rect 15555 8885 15625 8935
rect 15675 8885 15720 8935
rect 15770 8885 15815 8935
rect 15865 8885 15915 8935
rect 15965 8885 16015 8935
rect 16065 8885 16115 8935
rect 16165 8885 16210 8935
rect 16260 8885 16305 8935
rect 16355 8885 16425 8935
rect 16475 8885 16520 8935
rect 16570 8885 16615 8935
rect 16665 8885 16715 8935
rect 16765 8885 16815 8935
rect 16865 8885 16915 8935
rect 16965 8885 17010 8935
rect 17060 8885 17105 8935
rect 17155 8885 17225 8935
rect 17275 8885 17320 8935
rect 17370 8885 17415 8935
rect 17465 8885 17515 8935
rect 17565 8885 17615 8935
rect 17665 8885 17715 8935
rect 17765 8885 17810 8935
rect 17860 8885 17905 8935
rect 17955 8885 17990 8935
rect 14790 8815 17990 8885
rect 9010 8735 9020 8775
rect 9060 8735 9070 8775
rect 9010 8705 9070 8735
rect 9010 8665 9020 8705
rect 9060 8665 9070 8705
rect 9010 8635 9070 8665
rect 9010 8595 9020 8635
rect 9060 8595 9070 8635
rect 9010 8565 9070 8595
rect 9010 8525 9020 8565
rect 9060 8525 9070 8565
rect 9540 8695 9770 8780
rect 9890 8695 10120 8780
rect 10240 8695 10470 8780
rect 10590 8695 10820 8780
rect 10940 8695 11170 8780
rect 11290 8695 11520 8780
rect 11640 8695 11870 8780
rect 11990 8695 12220 8780
rect 12340 8695 12570 8780
rect 12690 8695 12920 8780
rect 13040 8695 13270 8780
rect 13390 8695 13620 8780
rect 13740 8695 13970 8780
rect 14090 8695 14320 8780
rect 14440 8695 14670 8780
rect 9540 8645 14670 8695
rect 9540 8550 9770 8645
rect 9890 8550 10120 8645
rect 10240 8550 10470 8645
rect 10590 8550 10820 8645
rect 10940 8550 11170 8645
rect 11290 8550 11520 8645
rect 11640 8550 11870 8645
rect 11990 8550 12220 8645
rect 12340 8550 12570 8645
rect 12690 8550 12920 8645
rect 13040 8550 13270 8645
rect 13390 8550 13620 8645
rect 13740 8550 13970 8645
rect 14090 8550 14320 8645
rect 14440 8550 14670 8645
rect 14790 8765 14825 8815
rect 14875 8765 14920 8815
rect 14970 8765 15015 8815
rect 15065 8765 15115 8815
rect 15165 8765 15215 8815
rect 15265 8765 15315 8815
rect 15365 8765 15410 8815
rect 15460 8765 15505 8815
rect 15555 8765 15625 8815
rect 15675 8765 15720 8815
rect 15770 8765 15815 8815
rect 15865 8765 15915 8815
rect 15965 8765 16015 8815
rect 16065 8765 16115 8815
rect 16165 8765 16210 8815
rect 16260 8765 16305 8815
rect 16355 8765 16425 8815
rect 16475 8765 16520 8815
rect 16570 8765 16615 8815
rect 16665 8765 16715 8815
rect 16765 8765 16815 8815
rect 16865 8765 16915 8815
rect 16965 8765 17010 8815
rect 17060 8765 17105 8815
rect 17155 8765 17225 8815
rect 17275 8765 17320 8815
rect 17370 8765 17415 8815
rect 17465 8765 17515 8815
rect 17565 8765 17615 8815
rect 17665 8765 17715 8815
rect 17765 8765 17810 8815
rect 17860 8765 17905 8815
rect 17955 8765 17990 8815
rect 14790 8725 17990 8765
rect 14790 8675 14825 8725
rect 14875 8675 14920 8725
rect 14970 8675 15015 8725
rect 15065 8675 15115 8725
rect 15165 8675 15215 8725
rect 15265 8675 15315 8725
rect 15365 8675 15410 8725
rect 15460 8675 15505 8725
rect 15555 8675 15625 8725
rect 15675 8675 15720 8725
rect 15770 8675 15815 8725
rect 15865 8675 15915 8725
rect 15965 8675 16015 8725
rect 16065 8675 16115 8725
rect 16165 8675 16210 8725
rect 16260 8675 16305 8725
rect 16355 8675 16425 8725
rect 16475 8675 16520 8725
rect 16570 8675 16615 8725
rect 16665 8675 16715 8725
rect 16765 8675 16815 8725
rect 16865 8675 16915 8725
rect 16965 8675 17010 8725
rect 17060 8675 17105 8725
rect 17155 8675 17225 8725
rect 17275 8675 17320 8725
rect 17370 8675 17415 8725
rect 17465 8675 17515 8725
rect 17565 8675 17615 8725
rect 17665 8675 17715 8725
rect 17765 8675 17810 8725
rect 17860 8675 17905 8725
rect 17955 8675 17990 8725
rect 14790 8625 17990 8675
rect 14790 8575 14825 8625
rect 14875 8575 14920 8625
rect 14970 8575 15015 8625
rect 15065 8575 15115 8625
rect 15165 8575 15215 8625
rect 15265 8575 15315 8625
rect 15365 8575 15410 8625
rect 15460 8575 15505 8625
rect 15555 8575 15625 8625
rect 15675 8575 15720 8625
rect 15770 8575 15815 8625
rect 15865 8575 15915 8625
rect 15965 8575 16015 8625
rect 16065 8575 16115 8625
rect 16165 8575 16210 8625
rect 16260 8575 16305 8625
rect 16355 8575 16425 8625
rect 16475 8575 16520 8625
rect 16570 8575 16615 8625
rect 16665 8575 16715 8625
rect 16765 8575 16815 8625
rect 16865 8575 16915 8625
rect 16965 8575 17010 8625
rect 17060 8575 17105 8625
rect 17155 8575 17225 8625
rect 17275 8575 17320 8625
rect 17370 8575 17415 8625
rect 17465 8575 17515 8625
rect 17565 8575 17615 8625
rect 17665 8575 17715 8625
rect 17765 8575 17810 8625
rect 17860 8575 17905 8625
rect 17955 8575 17990 8625
rect 9010 8500 9070 8525
rect 9010 8460 9020 8500
rect 9060 8460 9070 8500
rect 9010 8440 9070 8460
rect 9010 8400 9020 8440
rect 9060 8400 9070 8440
rect 12080 8430 12130 8550
rect 14790 8535 17990 8575
rect 14790 8485 14825 8535
rect 14875 8485 14920 8535
rect 14970 8485 15015 8535
rect 15065 8485 15115 8535
rect 15165 8485 15215 8535
rect 15265 8485 15315 8535
rect 15365 8485 15410 8535
rect 15460 8485 15505 8535
rect 15555 8485 15625 8535
rect 15675 8485 15720 8535
rect 15770 8485 15815 8535
rect 15865 8485 15915 8535
rect 15965 8485 16015 8535
rect 16065 8485 16115 8535
rect 16165 8485 16210 8535
rect 16260 8485 16305 8535
rect 16355 8485 16425 8535
rect 16475 8485 16520 8535
rect 16570 8485 16615 8535
rect 16665 8485 16715 8535
rect 16765 8485 16815 8535
rect 16865 8485 16915 8535
rect 16965 8485 17010 8535
rect 17060 8485 17105 8535
rect 17155 8485 17225 8535
rect 17275 8485 17320 8535
rect 17370 8485 17415 8535
rect 17465 8485 17515 8535
rect 17565 8485 17615 8535
rect 17665 8485 17715 8535
rect 17765 8485 17810 8535
rect 17860 8485 17905 8535
rect 17955 8485 17990 8535
rect 9010 8375 9070 8400
rect 9010 8335 9020 8375
rect 9060 8335 9070 8375
rect 9010 8305 9070 8335
rect 9010 8265 9020 8305
rect 9060 8265 9070 8305
rect 9010 8235 9070 8265
rect 9010 8195 9020 8235
rect 9060 8195 9070 8235
rect 9540 8345 9770 8430
rect 9890 8345 10120 8430
rect 10240 8345 10470 8430
rect 10590 8345 10820 8430
rect 10940 8345 11170 8430
rect 11290 8345 11520 8430
rect 11640 8345 11870 8430
rect 11990 8345 12220 8430
rect 12340 8345 12570 8430
rect 12690 8345 12920 8430
rect 13040 8345 13270 8430
rect 13390 8345 13620 8430
rect 13740 8345 13970 8430
rect 14090 8345 14320 8430
rect 14440 8345 14670 8430
rect 9540 8295 14670 8345
rect 9540 8200 9770 8295
rect 9890 8200 10120 8295
rect 10240 8200 10470 8295
rect 10590 8200 10820 8295
rect 10940 8200 11170 8295
rect 11290 8200 11520 8295
rect 11640 8200 11870 8295
rect 11990 8200 12220 8295
rect 12340 8200 12570 8295
rect 12690 8200 12920 8295
rect 13040 8200 13270 8295
rect 13390 8200 13620 8295
rect 13740 8200 13970 8295
rect 14090 8200 14320 8295
rect 14440 8200 14670 8295
rect 14790 8415 17990 8485
rect 14790 8365 14825 8415
rect 14875 8365 14920 8415
rect 14970 8365 15015 8415
rect 15065 8365 15115 8415
rect 15165 8365 15215 8415
rect 15265 8365 15315 8415
rect 15365 8365 15410 8415
rect 15460 8365 15505 8415
rect 15555 8365 15625 8415
rect 15675 8365 15720 8415
rect 15770 8365 15815 8415
rect 15865 8365 15915 8415
rect 15965 8365 16015 8415
rect 16065 8365 16115 8415
rect 16165 8365 16210 8415
rect 16260 8365 16305 8415
rect 16355 8365 16425 8415
rect 16475 8365 16520 8415
rect 16570 8365 16615 8415
rect 16665 8365 16715 8415
rect 16765 8365 16815 8415
rect 16865 8365 16915 8415
rect 16965 8365 17010 8415
rect 17060 8365 17105 8415
rect 17155 8365 17225 8415
rect 17275 8365 17320 8415
rect 17370 8365 17415 8415
rect 17465 8365 17515 8415
rect 17565 8365 17615 8415
rect 17665 8365 17715 8415
rect 17765 8365 17810 8415
rect 17860 8365 17905 8415
rect 17955 8365 17990 8415
rect 14790 8325 17990 8365
rect 14790 8275 14825 8325
rect 14875 8275 14920 8325
rect 14970 8275 15015 8325
rect 15065 8275 15115 8325
rect 15165 8275 15215 8325
rect 15265 8275 15315 8325
rect 15365 8275 15410 8325
rect 15460 8275 15505 8325
rect 15555 8275 15625 8325
rect 15675 8275 15720 8325
rect 15770 8275 15815 8325
rect 15865 8275 15915 8325
rect 15965 8275 16015 8325
rect 16065 8275 16115 8325
rect 16165 8275 16210 8325
rect 16260 8275 16305 8325
rect 16355 8275 16425 8325
rect 16475 8275 16520 8325
rect 16570 8275 16615 8325
rect 16665 8275 16715 8325
rect 16765 8275 16815 8325
rect 16865 8275 16915 8325
rect 16965 8275 17010 8325
rect 17060 8275 17105 8325
rect 17155 8275 17225 8325
rect 17275 8275 17320 8325
rect 17370 8275 17415 8325
rect 17465 8275 17515 8325
rect 17565 8275 17615 8325
rect 17665 8275 17715 8325
rect 17765 8275 17810 8325
rect 17860 8275 17905 8325
rect 17955 8275 17990 8325
rect 14790 8225 17990 8275
rect 9010 8165 9070 8195
rect 9010 8125 9020 8165
rect 9060 8125 9070 8165
rect 9010 8100 9070 8125
rect 9010 8060 9020 8100
rect 9060 8060 9070 8100
rect 12080 8080 12130 8200
rect 14790 8175 14825 8225
rect 14875 8175 14920 8225
rect 14970 8175 15015 8225
rect 15065 8175 15115 8225
rect 15165 8175 15215 8225
rect 15265 8175 15315 8225
rect 15365 8175 15410 8225
rect 15460 8175 15505 8225
rect 15555 8175 15625 8225
rect 15675 8175 15720 8225
rect 15770 8175 15815 8225
rect 15865 8175 15915 8225
rect 15965 8175 16015 8225
rect 16065 8175 16115 8225
rect 16165 8175 16210 8225
rect 16260 8175 16305 8225
rect 16355 8175 16425 8225
rect 16475 8175 16520 8225
rect 16570 8175 16615 8225
rect 16665 8175 16715 8225
rect 16765 8175 16815 8225
rect 16865 8175 16915 8225
rect 16965 8175 17010 8225
rect 17060 8175 17105 8225
rect 17155 8175 17225 8225
rect 17275 8175 17320 8225
rect 17370 8175 17415 8225
rect 17465 8175 17515 8225
rect 17565 8175 17615 8225
rect 17665 8175 17715 8225
rect 17765 8175 17810 8225
rect 17860 8175 17905 8225
rect 17955 8175 17990 8225
rect 14790 8135 17990 8175
rect 14790 8085 14825 8135
rect 14875 8085 14920 8135
rect 14970 8085 15015 8135
rect 15065 8085 15115 8135
rect 15165 8085 15215 8135
rect 15265 8085 15315 8135
rect 15365 8085 15410 8135
rect 15460 8085 15505 8135
rect 15555 8085 15625 8135
rect 15675 8085 15720 8135
rect 15770 8085 15815 8135
rect 15865 8085 15915 8135
rect 15965 8085 16015 8135
rect 16065 8085 16115 8135
rect 16165 8085 16210 8135
rect 16260 8085 16305 8135
rect 16355 8085 16425 8135
rect 16475 8085 16520 8135
rect 16570 8085 16615 8135
rect 16665 8085 16715 8135
rect 16765 8085 16815 8135
rect 16865 8085 16915 8135
rect 16965 8085 17010 8135
rect 17060 8085 17105 8135
rect 17155 8085 17225 8135
rect 17275 8085 17320 8135
rect 17370 8085 17415 8135
rect 17465 8085 17515 8135
rect 17565 8085 17615 8135
rect 17665 8085 17715 8135
rect 17765 8085 17810 8135
rect 17860 8085 17905 8135
rect 17955 8085 17990 8135
rect 9010 8040 9070 8060
rect 9010 8000 9020 8040
rect 9060 8000 9070 8040
rect 9010 7975 9070 8000
rect 9010 7935 9020 7975
rect 9060 7935 9070 7975
rect 9010 7905 9070 7935
rect 9010 7865 9020 7905
rect 9060 7865 9070 7905
rect 9010 7835 9070 7865
rect 9540 7995 9770 8080
rect 9890 7995 10120 8080
rect 10240 7995 10470 8080
rect 10590 7995 10820 8080
rect 10940 7995 11170 8080
rect 11290 7995 11520 8080
rect 11640 7995 11870 8080
rect 11990 7995 12220 8080
rect 12340 7995 12570 8080
rect 12690 7995 12920 8080
rect 13040 7995 13270 8080
rect 13390 7995 13620 8080
rect 13740 7995 13970 8080
rect 14090 7995 14320 8080
rect 14440 7995 14670 8080
rect 9540 7945 14670 7995
rect 9540 7850 9770 7945
rect 9890 7850 10120 7945
rect 10240 7850 10470 7945
rect 10590 7850 10820 7945
rect 10940 7850 11170 7945
rect 11290 7850 11520 7945
rect 11640 7850 11870 7945
rect 11990 7850 12220 7945
rect 12340 7850 12570 7945
rect 12690 7850 12920 7945
rect 13040 7850 13270 7945
rect 13390 7850 13620 7945
rect 13740 7850 13970 7945
rect 14090 7850 14320 7945
rect 14440 7850 14670 7945
rect 14790 8015 17990 8085
rect 14790 7965 14825 8015
rect 14875 7965 14920 8015
rect 14970 7965 15015 8015
rect 15065 7965 15115 8015
rect 15165 7965 15215 8015
rect 15265 7965 15315 8015
rect 15365 7965 15410 8015
rect 15460 7965 15505 8015
rect 15555 7965 15625 8015
rect 15675 7965 15720 8015
rect 15770 7965 15815 8015
rect 15865 7965 15915 8015
rect 15965 7965 16015 8015
rect 16065 7965 16115 8015
rect 16165 7965 16210 8015
rect 16260 7965 16305 8015
rect 16355 7965 16425 8015
rect 16475 7965 16520 8015
rect 16570 7965 16615 8015
rect 16665 7965 16715 8015
rect 16765 7965 16815 8015
rect 16865 7965 16915 8015
rect 16965 7965 17010 8015
rect 17060 7965 17105 8015
rect 17155 7965 17225 8015
rect 17275 7965 17320 8015
rect 17370 7965 17415 8015
rect 17465 7965 17515 8015
rect 17565 7965 17615 8015
rect 17665 7965 17715 8015
rect 17765 7965 17810 8015
rect 17860 7965 17905 8015
rect 17955 7965 17990 8015
rect 14790 7925 17990 7965
rect 14790 7875 14825 7925
rect 14875 7875 14920 7925
rect 14970 7875 15015 7925
rect 15065 7875 15115 7925
rect 15165 7875 15215 7925
rect 15265 7875 15315 7925
rect 15365 7875 15410 7925
rect 15460 7875 15505 7925
rect 15555 7875 15625 7925
rect 15675 7875 15720 7925
rect 15770 7875 15815 7925
rect 15865 7875 15915 7925
rect 15965 7875 16015 7925
rect 16065 7875 16115 7925
rect 16165 7875 16210 7925
rect 16260 7875 16305 7925
rect 16355 7875 16425 7925
rect 16475 7875 16520 7925
rect 16570 7875 16615 7925
rect 16665 7875 16715 7925
rect 16765 7875 16815 7925
rect 16865 7875 16915 7925
rect 16965 7875 17010 7925
rect 17060 7875 17105 7925
rect 17155 7875 17225 7925
rect 17275 7875 17320 7925
rect 17370 7875 17415 7925
rect 17465 7875 17515 7925
rect 17565 7875 17615 7925
rect 17665 7875 17715 7925
rect 17765 7875 17810 7925
rect 17860 7875 17905 7925
rect 17955 7875 17990 7925
rect 9010 7795 9020 7835
rect 9060 7795 9070 7835
rect 9010 7765 9070 7795
rect 9010 7725 9020 7765
rect 9060 7725 9070 7765
rect 12080 7730 12130 7850
rect 14790 7825 17990 7875
rect 14790 7775 14825 7825
rect 14875 7775 14920 7825
rect 14970 7775 15015 7825
rect 15065 7775 15115 7825
rect 15165 7775 15215 7825
rect 15265 7775 15315 7825
rect 15365 7775 15410 7825
rect 15460 7775 15505 7825
rect 15555 7775 15625 7825
rect 15675 7775 15720 7825
rect 15770 7775 15815 7825
rect 15865 7775 15915 7825
rect 15965 7775 16015 7825
rect 16065 7775 16115 7825
rect 16165 7775 16210 7825
rect 16260 7775 16305 7825
rect 16355 7775 16425 7825
rect 16475 7775 16520 7825
rect 16570 7775 16615 7825
rect 16665 7775 16715 7825
rect 16765 7775 16815 7825
rect 16865 7775 16915 7825
rect 16965 7775 17010 7825
rect 17060 7775 17105 7825
rect 17155 7775 17225 7825
rect 17275 7775 17320 7825
rect 17370 7775 17415 7825
rect 17465 7775 17515 7825
rect 17565 7775 17615 7825
rect 17665 7775 17715 7825
rect 17765 7775 17810 7825
rect 17860 7775 17905 7825
rect 17955 7775 17990 7825
rect 14790 7735 17990 7775
rect 9010 7700 9070 7725
rect 9010 7660 9020 7700
rect 9060 7660 9070 7700
rect 9010 7640 9070 7660
rect 9010 7600 9020 7640
rect 9060 7600 9070 7640
rect 9010 7575 9070 7600
rect 9010 7535 9020 7575
rect 9060 7535 9070 7575
rect 9010 7505 9070 7535
rect 9010 7465 9020 7505
rect 9060 7465 9070 7505
rect 9540 7645 9770 7730
rect 9890 7645 10120 7730
rect 10240 7645 10470 7730
rect 10590 7645 10820 7730
rect 10940 7645 11170 7730
rect 11290 7645 11520 7730
rect 11640 7645 11870 7730
rect 11990 7645 12220 7730
rect 12340 7645 12570 7730
rect 12690 7645 12920 7730
rect 13040 7645 13270 7730
rect 13390 7645 13620 7730
rect 13740 7645 13970 7730
rect 14090 7645 14320 7730
rect 14440 7645 14670 7730
rect 9540 7595 14670 7645
rect 9540 7500 9770 7595
rect 9890 7500 10120 7595
rect 10240 7500 10470 7595
rect 10590 7500 10820 7595
rect 10940 7500 11170 7595
rect 11290 7500 11520 7595
rect 11640 7500 11870 7595
rect 11990 7500 12220 7595
rect 12340 7500 12570 7595
rect 12690 7500 12920 7595
rect 13040 7500 13270 7595
rect 13390 7500 13620 7595
rect 13740 7500 13970 7595
rect 14090 7500 14320 7595
rect 14440 7500 14670 7595
rect 14790 7685 14825 7735
rect 14875 7685 14920 7735
rect 14970 7685 15015 7735
rect 15065 7685 15115 7735
rect 15165 7685 15215 7735
rect 15265 7685 15315 7735
rect 15365 7685 15410 7735
rect 15460 7685 15505 7735
rect 15555 7685 15625 7735
rect 15675 7685 15720 7735
rect 15770 7685 15815 7735
rect 15865 7685 15915 7735
rect 15965 7685 16015 7735
rect 16065 7685 16115 7735
rect 16165 7685 16210 7735
rect 16260 7685 16305 7735
rect 16355 7685 16425 7735
rect 16475 7685 16520 7735
rect 16570 7685 16615 7735
rect 16665 7685 16715 7735
rect 16765 7685 16815 7735
rect 16865 7685 16915 7735
rect 16965 7685 17010 7735
rect 17060 7685 17105 7735
rect 17155 7685 17225 7735
rect 17275 7685 17320 7735
rect 17370 7685 17415 7735
rect 17465 7685 17515 7735
rect 17565 7685 17615 7735
rect 17665 7685 17715 7735
rect 17765 7685 17810 7735
rect 17860 7685 17905 7735
rect 17955 7685 17990 7735
rect 14790 7615 17990 7685
rect 14790 7565 14825 7615
rect 14875 7565 14920 7615
rect 14970 7565 15015 7615
rect 15065 7565 15115 7615
rect 15165 7565 15215 7615
rect 15265 7565 15315 7615
rect 15365 7565 15410 7615
rect 15460 7565 15505 7615
rect 15555 7565 15625 7615
rect 15675 7565 15720 7615
rect 15770 7565 15815 7615
rect 15865 7565 15915 7615
rect 15965 7565 16015 7615
rect 16065 7565 16115 7615
rect 16165 7565 16210 7615
rect 16260 7565 16305 7615
rect 16355 7565 16425 7615
rect 16475 7565 16520 7615
rect 16570 7565 16615 7615
rect 16665 7565 16715 7615
rect 16765 7565 16815 7615
rect 16865 7565 16915 7615
rect 16965 7565 17010 7615
rect 17060 7565 17105 7615
rect 17155 7565 17225 7615
rect 17275 7565 17320 7615
rect 17370 7565 17415 7615
rect 17465 7565 17515 7615
rect 17565 7565 17615 7615
rect 17665 7565 17715 7615
rect 17765 7565 17810 7615
rect 17860 7565 17905 7615
rect 17955 7565 17990 7615
rect 14790 7525 17990 7565
rect 9010 7435 9070 7465
rect 9010 7395 9020 7435
rect 9060 7395 9070 7435
rect 9010 7365 9070 7395
rect 12080 7380 12130 7500
rect 14790 7475 14825 7525
rect 14875 7475 14920 7525
rect 14970 7475 15015 7525
rect 15065 7475 15115 7525
rect 15165 7475 15215 7525
rect 15265 7475 15315 7525
rect 15365 7475 15410 7525
rect 15460 7475 15505 7525
rect 15555 7475 15625 7525
rect 15675 7475 15720 7525
rect 15770 7475 15815 7525
rect 15865 7475 15915 7525
rect 15965 7475 16015 7525
rect 16065 7475 16115 7525
rect 16165 7475 16210 7525
rect 16260 7475 16305 7525
rect 16355 7475 16425 7525
rect 16475 7475 16520 7525
rect 16570 7475 16615 7525
rect 16665 7475 16715 7525
rect 16765 7475 16815 7525
rect 16865 7475 16915 7525
rect 16965 7475 17010 7525
rect 17060 7475 17105 7525
rect 17155 7475 17225 7525
rect 17275 7475 17320 7525
rect 17370 7475 17415 7525
rect 17465 7475 17515 7525
rect 17565 7475 17615 7525
rect 17665 7475 17715 7525
rect 17765 7475 17810 7525
rect 17860 7475 17905 7525
rect 17955 7475 17990 7525
rect 14790 7425 17990 7475
rect 9010 7325 9020 7365
rect 9060 7325 9070 7365
rect 9010 7300 9070 7325
rect 9010 7260 9020 7300
rect 9060 7260 9070 7300
rect 9010 7240 9070 7260
rect 9010 7200 9020 7240
rect 9060 7200 9070 7240
rect 9010 7175 9070 7200
rect 9010 7135 9020 7175
rect 9060 7135 9070 7175
rect 9540 7295 9770 7380
rect 9890 7295 10120 7380
rect 10240 7295 10470 7380
rect 10590 7295 10820 7380
rect 10940 7295 11170 7380
rect 11290 7295 11520 7380
rect 11640 7295 11870 7380
rect 11990 7295 12220 7380
rect 12340 7295 12570 7380
rect 12690 7295 12920 7380
rect 13040 7295 13270 7380
rect 13390 7295 13620 7380
rect 13740 7295 13970 7380
rect 14090 7295 14320 7380
rect 14440 7295 14670 7380
rect 9540 7245 14670 7295
rect 9540 7150 9770 7245
rect 9890 7150 10120 7245
rect 10240 7150 10470 7245
rect 10590 7150 10820 7245
rect 10940 7150 11170 7245
rect 11290 7150 11520 7245
rect 11640 7150 11870 7245
rect 11990 7150 12220 7245
rect 12340 7150 12570 7245
rect 12690 7150 12920 7245
rect 13040 7150 13270 7245
rect 13390 7150 13620 7245
rect 13740 7150 13970 7245
rect 14090 7150 14320 7245
rect 14440 7150 14670 7245
rect 14790 7375 14825 7425
rect 14875 7375 14920 7425
rect 14970 7375 15015 7425
rect 15065 7375 15115 7425
rect 15165 7375 15215 7425
rect 15265 7375 15315 7425
rect 15365 7375 15410 7425
rect 15460 7375 15505 7425
rect 15555 7375 15625 7425
rect 15675 7375 15720 7425
rect 15770 7375 15815 7425
rect 15865 7375 15915 7425
rect 15965 7375 16015 7425
rect 16065 7375 16115 7425
rect 16165 7375 16210 7425
rect 16260 7375 16305 7425
rect 16355 7375 16425 7425
rect 16475 7375 16520 7425
rect 16570 7375 16615 7425
rect 16665 7375 16715 7425
rect 16765 7375 16815 7425
rect 16865 7375 16915 7425
rect 16965 7375 17010 7425
rect 17060 7375 17105 7425
rect 17155 7375 17225 7425
rect 17275 7375 17320 7425
rect 17370 7375 17415 7425
rect 17465 7375 17515 7425
rect 17565 7375 17615 7425
rect 17665 7375 17715 7425
rect 17765 7375 17810 7425
rect 17860 7375 17905 7425
rect 17955 7375 17990 7425
rect 14790 7335 17990 7375
rect 14790 7285 14825 7335
rect 14875 7285 14920 7335
rect 14970 7285 15015 7335
rect 15065 7285 15115 7335
rect 15165 7285 15215 7335
rect 15265 7285 15315 7335
rect 15365 7285 15410 7335
rect 15460 7285 15505 7335
rect 15555 7285 15625 7335
rect 15675 7285 15720 7335
rect 15770 7285 15815 7335
rect 15865 7285 15915 7335
rect 15965 7285 16015 7335
rect 16065 7285 16115 7335
rect 16165 7285 16210 7335
rect 16260 7285 16305 7335
rect 16355 7285 16425 7335
rect 16475 7285 16520 7335
rect 16570 7285 16615 7335
rect 16665 7285 16715 7335
rect 16765 7285 16815 7335
rect 16865 7285 16915 7335
rect 16965 7285 17010 7335
rect 17060 7285 17105 7335
rect 17155 7285 17225 7335
rect 17275 7285 17320 7335
rect 17370 7285 17415 7335
rect 17465 7285 17515 7335
rect 17565 7285 17615 7335
rect 17665 7285 17715 7335
rect 17765 7285 17810 7335
rect 17860 7285 17905 7335
rect 17955 7285 17990 7335
rect 14790 7215 17990 7285
rect 14790 7165 14825 7215
rect 14875 7165 14920 7215
rect 14970 7165 15015 7215
rect 15065 7165 15115 7215
rect 15165 7165 15215 7215
rect 15265 7165 15315 7215
rect 15365 7165 15410 7215
rect 15460 7165 15505 7215
rect 15555 7165 15625 7215
rect 15675 7165 15720 7215
rect 15770 7165 15815 7215
rect 15865 7165 15915 7215
rect 15965 7165 16015 7215
rect 16065 7165 16115 7215
rect 16165 7165 16210 7215
rect 16260 7165 16305 7215
rect 16355 7165 16425 7215
rect 16475 7165 16520 7215
rect 16570 7165 16615 7215
rect 16665 7165 16715 7215
rect 16765 7165 16815 7215
rect 16865 7165 16915 7215
rect 16965 7165 17010 7215
rect 17060 7165 17105 7215
rect 17155 7165 17225 7215
rect 17275 7165 17320 7215
rect 17370 7165 17415 7215
rect 17465 7165 17515 7215
rect 17565 7165 17615 7215
rect 17665 7165 17715 7215
rect 17765 7165 17810 7215
rect 17860 7165 17905 7215
rect 17955 7165 17990 7215
rect 9010 7105 9070 7135
rect 9010 7065 9020 7105
rect 9060 7065 9070 7105
rect 9010 7035 9070 7065
rect 9010 6995 9020 7035
rect 9060 6995 9070 7035
rect 12080 7030 12130 7150
rect 14790 7125 17990 7165
rect 14790 7075 14825 7125
rect 14875 7075 14920 7125
rect 14970 7075 15015 7125
rect 15065 7075 15115 7125
rect 15165 7075 15215 7125
rect 15265 7075 15315 7125
rect 15365 7075 15410 7125
rect 15460 7075 15505 7125
rect 15555 7075 15625 7125
rect 15675 7075 15720 7125
rect 15770 7075 15815 7125
rect 15865 7075 15915 7125
rect 15965 7075 16015 7125
rect 16065 7075 16115 7125
rect 16165 7075 16210 7125
rect 16260 7075 16305 7125
rect 16355 7075 16425 7125
rect 16475 7075 16520 7125
rect 16570 7075 16615 7125
rect 16665 7075 16715 7125
rect 16765 7075 16815 7125
rect 16865 7075 16915 7125
rect 16965 7075 17010 7125
rect 17060 7075 17105 7125
rect 17155 7075 17225 7125
rect 17275 7075 17320 7125
rect 17370 7075 17415 7125
rect 17465 7075 17515 7125
rect 17565 7075 17615 7125
rect 17665 7075 17715 7125
rect 17765 7075 17810 7125
rect 17860 7075 17905 7125
rect 17955 7075 17990 7125
rect 9010 6965 9070 6995
rect 9010 6925 9020 6965
rect 9060 6925 9070 6965
rect 9010 6900 9070 6925
rect 9010 6860 9020 6900
rect 9060 6860 9070 6900
rect 9010 6840 9070 6860
rect 9010 6800 9020 6840
rect 9060 6800 9070 6840
rect 9540 6945 9770 7030
rect 9890 6945 10120 7030
rect 10240 6945 10470 7030
rect 10590 6945 10820 7030
rect 10940 6945 11170 7030
rect 11290 6945 11520 7030
rect 11640 6945 11870 7030
rect 11990 6945 12220 7030
rect 12340 6945 12570 7030
rect 12690 6945 12920 7030
rect 13040 6945 13270 7030
rect 13390 6945 13620 7030
rect 13740 6945 13970 7030
rect 14090 6945 14320 7030
rect 14440 6945 14670 7030
rect 9540 6895 14670 6945
rect 9540 6800 9770 6895
rect 9890 6800 10120 6895
rect 10240 6800 10470 6895
rect 10590 6800 10820 6895
rect 10940 6800 11170 6895
rect 11290 6800 11520 6895
rect 11640 6800 11870 6895
rect 11990 6800 12220 6895
rect 12340 6800 12570 6895
rect 12690 6800 12920 6895
rect 13040 6800 13270 6895
rect 13390 6800 13620 6895
rect 13740 6800 13970 6895
rect 14090 6800 14320 6895
rect 14440 6800 14670 6895
rect 14790 7025 17990 7075
rect 14790 6975 14825 7025
rect 14875 6975 14920 7025
rect 14970 6975 15015 7025
rect 15065 6975 15115 7025
rect 15165 6975 15215 7025
rect 15265 6975 15315 7025
rect 15365 6975 15410 7025
rect 15460 6975 15505 7025
rect 15555 6975 15625 7025
rect 15675 6975 15720 7025
rect 15770 6975 15815 7025
rect 15865 6975 15915 7025
rect 15965 6975 16015 7025
rect 16065 6975 16115 7025
rect 16165 6975 16210 7025
rect 16260 6975 16305 7025
rect 16355 6975 16425 7025
rect 16475 6975 16520 7025
rect 16570 6975 16615 7025
rect 16665 6975 16715 7025
rect 16765 6975 16815 7025
rect 16865 6975 16915 7025
rect 16965 6975 17010 7025
rect 17060 6975 17105 7025
rect 17155 6975 17225 7025
rect 17275 6975 17320 7025
rect 17370 6975 17415 7025
rect 17465 6975 17515 7025
rect 17565 6975 17615 7025
rect 17665 6975 17715 7025
rect 17765 6975 17810 7025
rect 17860 6975 17905 7025
rect 17955 6975 17990 7025
rect 14790 6935 17990 6975
rect 14790 6885 14825 6935
rect 14875 6885 14920 6935
rect 14970 6885 15015 6935
rect 15065 6885 15115 6935
rect 15165 6885 15215 6935
rect 15265 6885 15315 6935
rect 15365 6885 15410 6935
rect 15460 6885 15505 6935
rect 15555 6885 15625 6935
rect 15675 6885 15720 6935
rect 15770 6885 15815 6935
rect 15865 6885 15915 6935
rect 15965 6885 16015 6935
rect 16065 6885 16115 6935
rect 16165 6885 16210 6935
rect 16260 6885 16305 6935
rect 16355 6885 16425 6935
rect 16475 6885 16520 6935
rect 16570 6885 16615 6935
rect 16665 6885 16715 6935
rect 16765 6885 16815 6935
rect 16865 6885 16915 6935
rect 16965 6885 17010 6935
rect 17060 6885 17105 6935
rect 17155 6885 17225 6935
rect 17275 6885 17320 6935
rect 17370 6885 17415 6935
rect 17465 6885 17515 6935
rect 17565 6885 17615 6935
rect 17665 6885 17715 6935
rect 17765 6885 17810 6935
rect 17860 6885 17905 6935
rect 17955 6885 17990 6935
rect 14790 6815 17990 6885
rect 9010 6775 9070 6800
rect 9010 6735 9020 6775
rect 9060 6735 9070 6775
rect 9010 6705 9070 6735
rect 9010 6665 9020 6705
rect 9060 6665 9070 6705
rect 12080 6680 12130 6800
rect 14790 6765 14825 6815
rect 14875 6765 14920 6815
rect 14970 6765 15015 6815
rect 15065 6765 15115 6815
rect 15165 6765 15215 6815
rect 15265 6765 15315 6815
rect 15365 6765 15410 6815
rect 15460 6765 15505 6815
rect 15555 6765 15625 6815
rect 15675 6765 15720 6815
rect 15770 6765 15815 6815
rect 15865 6765 15915 6815
rect 15965 6765 16015 6815
rect 16065 6765 16115 6815
rect 16165 6765 16210 6815
rect 16260 6765 16305 6815
rect 16355 6765 16425 6815
rect 16475 6765 16520 6815
rect 16570 6765 16615 6815
rect 16665 6765 16715 6815
rect 16765 6765 16815 6815
rect 16865 6765 16915 6815
rect 16965 6765 17010 6815
rect 17060 6765 17105 6815
rect 17155 6765 17225 6815
rect 17275 6765 17320 6815
rect 17370 6765 17415 6815
rect 17465 6765 17515 6815
rect 17565 6765 17615 6815
rect 17665 6765 17715 6815
rect 17765 6765 17810 6815
rect 17860 6765 17905 6815
rect 17955 6765 17990 6815
rect 14790 6725 17990 6765
rect 9010 6635 9070 6665
rect 9010 6595 9020 6635
rect 9060 6595 9070 6635
rect 9010 6565 9070 6595
rect 9010 6525 9020 6565
rect 9060 6525 9070 6565
rect 9010 6500 9070 6525
rect 9010 6460 9020 6500
rect 9060 6460 9070 6500
rect 9010 6450 9070 6460
rect 9540 6595 9770 6680
rect 9890 6595 10120 6680
rect 10240 6595 10470 6680
rect 10590 6595 10820 6680
rect 10940 6595 11170 6680
rect 11290 6595 11520 6680
rect 11640 6595 11870 6680
rect 11990 6595 12220 6680
rect 12340 6595 12570 6680
rect 12690 6595 12920 6680
rect 13040 6595 13270 6680
rect 13390 6595 13620 6680
rect 13740 6595 13970 6680
rect 14090 6595 14320 6680
rect 14440 6595 14670 6680
rect 9540 6545 14670 6595
rect 9540 6450 9770 6545
rect 9890 6450 10120 6545
rect 10240 6450 10470 6545
rect 10590 6450 10820 6545
rect 10940 6450 11170 6545
rect 11290 6450 11520 6545
rect 11640 6450 11870 6545
rect 11990 6450 12220 6545
rect 12340 6450 12570 6545
rect 12690 6450 12920 6545
rect 13040 6450 13270 6545
rect 13390 6450 13620 6545
rect 13740 6450 13970 6545
rect 14090 6450 14320 6545
rect 14440 6450 14670 6545
rect 14790 6675 14825 6725
rect 14875 6675 14920 6725
rect 14970 6675 15015 6725
rect 15065 6675 15115 6725
rect 15165 6675 15215 6725
rect 15265 6675 15315 6725
rect 15365 6675 15410 6725
rect 15460 6675 15505 6725
rect 15555 6675 15625 6725
rect 15675 6675 15720 6725
rect 15770 6675 15815 6725
rect 15865 6675 15915 6725
rect 15965 6675 16015 6725
rect 16065 6675 16115 6725
rect 16165 6675 16210 6725
rect 16260 6675 16305 6725
rect 16355 6675 16425 6725
rect 16475 6675 16520 6725
rect 16570 6675 16615 6725
rect 16665 6675 16715 6725
rect 16765 6675 16815 6725
rect 16865 6675 16915 6725
rect 16965 6675 17010 6725
rect 17060 6675 17105 6725
rect 17155 6675 17225 6725
rect 17275 6675 17320 6725
rect 17370 6675 17415 6725
rect 17465 6675 17515 6725
rect 17565 6675 17615 6725
rect 17665 6675 17715 6725
rect 17765 6675 17810 6725
rect 17860 6675 17905 6725
rect 17955 6675 17990 6725
rect 14790 6625 17990 6675
rect 14790 6575 14825 6625
rect 14875 6575 14920 6625
rect 14970 6575 15015 6625
rect 15065 6575 15115 6625
rect 15165 6575 15215 6625
rect 15265 6575 15315 6625
rect 15365 6575 15410 6625
rect 15460 6575 15505 6625
rect 15555 6575 15625 6625
rect 15675 6575 15720 6625
rect 15770 6575 15815 6625
rect 15865 6575 15915 6625
rect 15965 6575 16015 6625
rect 16065 6575 16115 6625
rect 16165 6575 16210 6625
rect 16260 6575 16305 6625
rect 16355 6575 16425 6625
rect 16475 6575 16520 6625
rect 16570 6575 16615 6625
rect 16665 6575 16715 6625
rect 16765 6575 16815 6625
rect 16865 6575 16915 6625
rect 16965 6575 17010 6625
rect 17060 6575 17105 6625
rect 17155 6575 17225 6625
rect 17275 6575 17320 6625
rect 17370 6575 17415 6625
rect 17465 6575 17515 6625
rect 17565 6575 17615 6625
rect 17665 6575 17715 6625
rect 17765 6575 17810 6625
rect 17860 6575 17905 6625
rect 17955 6575 17990 6625
rect 14790 6535 17990 6575
rect 14790 6485 14825 6535
rect 14875 6485 14920 6535
rect 14970 6485 15015 6535
rect 15065 6485 15115 6535
rect 15165 6485 15215 6535
rect 15265 6485 15315 6535
rect 15365 6485 15410 6535
rect 15460 6485 15505 6535
rect 15555 6485 15625 6535
rect 15675 6485 15720 6535
rect 15770 6485 15815 6535
rect 15865 6485 15915 6535
rect 15965 6485 16015 6535
rect 16065 6485 16115 6535
rect 16165 6485 16210 6535
rect 16260 6485 16305 6535
rect 16355 6485 16425 6535
rect 16475 6485 16520 6535
rect 16570 6485 16615 6535
rect 16665 6485 16715 6535
rect 16765 6485 16815 6535
rect 16865 6485 16915 6535
rect 16965 6485 17010 6535
rect 17060 6485 17105 6535
rect 17155 6485 17225 6535
rect 17275 6485 17320 6535
rect 17370 6485 17415 6535
rect 17465 6485 17515 6535
rect 17565 6485 17615 6535
rect 17665 6485 17715 6535
rect 17765 6485 17810 6535
rect 17860 6485 17905 6535
rect 17955 6485 17990 6535
rect 1500 1370 1510 1380
rect -90 -1300 -30 -1290
rect -90 -1340 -80 -1300
rect -40 -1340 -30 -1300
rect -90 -1365 -30 -1340
rect -90 -1405 -80 -1365
rect -40 -1405 -30 -1365
rect -90 -1435 -30 -1405
rect -90 -1475 -80 -1435
rect -40 -1475 -30 -1435
rect -90 -1505 -30 -1475
rect -90 -1545 -80 -1505
rect -40 -1545 -30 -1505
rect -90 -1575 -30 -1545
rect -90 -1615 -80 -1575
rect -40 -1615 -30 -1575
rect -90 -1640 -30 -1615
rect -90 -1680 -80 -1640
rect -40 -1680 -30 -1640
rect -90 -1700 -30 -1680
rect -90 -1740 -80 -1700
rect -40 -1740 -30 -1700
rect -90 -1765 -30 -1740
rect -90 -1805 -80 -1765
rect -40 -1805 -30 -1765
rect -90 -1835 -30 -1805
rect -90 -1875 -80 -1835
rect -40 -1875 -30 -1835
rect -90 -1905 -30 -1875
rect -90 -1945 -80 -1905
rect -40 -1945 -30 -1905
rect -90 -1975 -30 -1945
rect -90 -2015 -80 -1975
rect -40 -2015 -30 -1975
rect -90 -2040 -30 -2015
rect -90 -2080 -80 -2040
rect -40 -2080 -30 -2040
rect -90 -2100 -30 -2080
rect -90 -2140 -80 -2100
rect -40 -2140 -30 -2100
rect -90 -2165 -30 -2140
rect -90 -2205 -80 -2165
rect -40 -2205 -30 -2165
rect -90 -2235 -30 -2205
rect -90 -2275 -80 -2235
rect -40 -2275 -30 -2235
rect -90 -2305 -30 -2275
rect -90 -2345 -80 -2305
rect -40 -2345 -30 -2305
rect -90 -2375 -30 -2345
rect -90 -2415 -80 -2375
rect -40 -2415 -30 -2375
rect -90 -2440 -30 -2415
rect -90 -2480 -80 -2440
rect -40 -2480 -30 -2440
rect -90 -2500 -30 -2480
rect -90 -2540 -80 -2500
rect -40 -2540 -30 -2500
rect -90 -2565 -30 -2540
rect -90 -2605 -80 -2565
rect -40 -2605 -30 -2565
rect -90 -2635 -30 -2605
rect -90 -2675 -80 -2635
rect -40 -2675 -30 -2635
rect -90 -2705 -30 -2675
rect -90 -2745 -80 -2705
rect -40 -2745 -30 -2705
rect -90 -2775 -30 -2745
rect -90 -2815 -80 -2775
rect -40 -2815 -30 -2775
rect -90 -2840 -30 -2815
rect -90 -2880 -80 -2840
rect -40 -2880 -30 -2840
rect -90 -2900 -30 -2880
rect -90 -2940 -80 -2900
rect -40 -2940 -30 -2900
rect -90 -2965 -30 -2940
rect -90 -3005 -80 -2965
rect -40 -3005 -30 -2965
rect -90 -3035 -30 -3005
rect -90 -3075 -80 -3035
rect -40 -3075 -30 -3035
rect -90 -3105 -30 -3075
rect -90 -3145 -80 -3105
rect -40 -3145 -30 -3105
rect -90 -3175 -30 -3145
rect -90 -3215 -80 -3175
rect -40 -3215 -30 -3175
rect -90 -3240 -30 -3215
rect -90 -3280 -80 -3240
rect -40 -3280 -30 -3240
rect -90 -3300 -30 -3280
rect -90 -3340 -80 -3300
rect -40 -3340 -30 -3300
rect -90 -3365 -30 -3340
rect -90 -3405 -80 -3365
rect -40 -3405 -30 -3365
rect -90 -3435 -30 -3405
rect -90 -3475 -80 -3435
rect -40 -3475 -30 -3435
rect -90 -3505 -30 -3475
rect -90 -3545 -80 -3505
rect -40 -3545 -30 -3505
rect -90 -3575 -30 -3545
rect -90 -3615 -80 -3575
rect -40 -3615 -30 -3575
rect -90 -3640 -30 -3615
rect -90 -3680 -80 -3640
rect -40 -3680 -30 -3640
rect -90 -3700 -30 -3680
rect -90 -3740 -80 -3700
rect -40 -3740 -30 -3700
rect -90 -3765 -30 -3740
rect -90 -3805 -80 -3765
rect -40 -3805 -30 -3765
rect -90 -3835 -30 -3805
rect -90 -3875 -80 -3835
rect -40 -3875 -30 -3835
rect -90 -3905 -30 -3875
rect -90 -3945 -80 -3905
rect -40 -3945 -30 -3905
rect -90 -3975 -30 -3945
rect -90 -4015 -80 -3975
rect -40 -4015 -30 -3975
rect -90 -4040 -30 -4015
rect -90 -4080 -80 -4040
rect -40 -4080 -30 -4040
rect -90 -4100 -30 -4080
rect -90 -4140 -80 -4100
rect -40 -4140 -30 -4100
rect -90 -4165 -30 -4140
rect -90 -4205 -80 -4165
rect -40 -4205 -30 -4165
rect -90 -4235 -30 -4205
rect -90 -4275 -80 -4235
rect -40 -4275 -30 -4235
rect -90 -4305 -30 -4275
rect -90 -4345 -80 -4305
rect -40 -4345 -30 -4305
rect -90 -4375 -30 -4345
rect -90 -4415 -80 -4375
rect -40 -4415 -30 -4375
rect -90 -4440 -30 -4415
rect -90 -4480 -80 -4440
rect -40 -4480 -30 -4440
rect -90 -4490 -30 -4480
rect 260 -1300 320 -1290
rect 260 -1340 270 -1300
rect 310 -1340 320 -1300
rect 260 -1365 320 -1340
rect 260 -1405 270 -1365
rect 310 -1405 320 -1365
rect 260 -1435 320 -1405
rect 260 -1475 270 -1435
rect 310 -1475 320 -1435
rect 260 -1505 320 -1475
rect 260 -1545 270 -1505
rect 310 -1545 320 -1505
rect 260 -1575 320 -1545
rect 260 -1615 270 -1575
rect 310 -1615 320 -1575
rect 260 -1640 320 -1615
rect 260 -1680 270 -1640
rect 310 -1680 320 -1640
rect 260 -1700 320 -1680
rect 260 -1740 270 -1700
rect 310 -1740 320 -1700
rect 260 -1765 320 -1740
rect 260 -1805 270 -1765
rect 310 -1805 320 -1765
rect 260 -1835 320 -1805
rect 260 -1875 270 -1835
rect 310 -1875 320 -1835
rect 260 -1905 320 -1875
rect 260 -1945 270 -1905
rect 310 -1945 320 -1905
rect 260 -1975 320 -1945
rect 260 -2015 270 -1975
rect 310 -2015 320 -1975
rect 260 -2040 320 -2015
rect 260 -2080 270 -2040
rect 310 -2080 320 -2040
rect 260 -2100 320 -2080
rect 260 -2140 270 -2100
rect 310 -2140 320 -2100
rect 260 -2165 320 -2140
rect 260 -2205 270 -2165
rect 310 -2205 320 -2165
rect 260 -2235 320 -2205
rect 260 -2275 270 -2235
rect 310 -2275 320 -2235
rect 260 -2305 320 -2275
rect 260 -2345 270 -2305
rect 310 -2345 320 -2305
rect 260 -2375 320 -2345
rect 260 -2415 270 -2375
rect 310 -2415 320 -2375
rect 260 -2440 320 -2415
rect 260 -2480 270 -2440
rect 310 -2480 320 -2440
rect 260 -2500 320 -2480
rect 260 -2540 270 -2500
rect 310 -2540 320 -2500
rect 260 -2565 320 -2540
rect 260 -2605 270 -2565
rect 310 -2605 320 -2565
rect 260 -2635 320 -2605
rect 260 -2675 270 -2635
rect 310 -2675 320 -2635
rect 260 -2705 320 -2675
rect 260 -2745 270 -2705
rect 310 -2745 320 -2705
rect 260 -2775 320 -2745
rect 260 -2815 270 -2775
rect 310 -2815 320 -2775
rect 260 -2840 320 -2815
rect 260 -2880 270 -2840
rect 310 -2880 320 -2840
rect 260 -2900 320 -2880
rect 260 -2940 270 -2900
rect 310 -2940 320 -2900
rect 260 -2965 320 -2940
rect 260 -3005 270 -2965
rect 310 -3005 320 -2965
rect 260 -3035 320 -3005
rect 260 -3075 270 -3035
rect 310 -3075 320 -3035
rect 260 -3105 320 -3075
rect 260 -3145 270 -3105
rect 310 -3145 320 -3105
rect 260 -3175 320 -3145
rect 260 -3215 270 -3175
rect 310 -3215 320 -3175
rect 260 -3240 320 -3215
rect 260 -3280 270 -3240
rect 310 -3280 320 -3240
rect 260 -3300 320 -3280
rect 260 -3340 270 -3300
rect 310 -3340 320 -3300
rect 260 -3365 320 -3340
rect 260 -3405 270 -3365
rect 310 -3405 320 -3365
rect 260 -3435 320 -3405
rect 260 -3475 270 -3435
rect 310 -3475 320 -3435
rect 260 -3505 320 -3475
rect 260 -3545 270 -3505
rect 310 -3545 320 -3505
rect 260 -3575 320 -3545
rect 260 -3615 270 -3575
rect 310 -3615 320 -3575
rect 260 -3640 320 -3615
rect 260 -3680 270 -3640
rect 310 -3680 320 -3640
rect 260 -3700 320 -3680
rect 260 -3740 270 -3700
rect 310 -3740 320 -3700
rect 260 -3765 320 -3740
rect 260 -3805 270 -3765
rect 310 -3805 320 -3765
rect 260 -3835 320 -3805
rect 260 -3875 270 -3835
rect 310 -3875 320 -3835
rect 260 -3905 320 -3875
rect 260 -3945 270 -3905
rect 310 -3945 320 -3905
rect 260 -3975 320 -3945
rect 260 -4015 270 -3975
rect 310 -4015 320 -3975
rect 260 -4040 320 -4015
rect 260 -4080 270 -4040
rect 310 -4080 320 -4040
rect 260 -4100 320 -4080
rect 260 -4140 270 -4100
rect 310 -4140 320 -4100
rect 260 -4165 320 -4140
rect 260 -4205 270 -4165
rect 310 -4205 320 -4165
rect 260 -4235 320 -4205
rect 260 -4275 270 -4235
rect 310 -4275 320 -4235
rect 260 -4305 320 -4275
rect 260 -4345 270 -4305
rect 310 -4345 320 -4305
rect 260 -4375 320 -4345
rect 260 -4415 270 -4375
rect 310 -4415 320 -4375
rect 260 -4440 320 -4415
rect 260 -4480 270 -4440
rect 310 -4480 320 -4440
rect 260 -4490 320 -4480
rect 610 -1300 670 -1290
rect 610 -1340 620 -1300
rect 660 -1340 670 -1300
rect 610 -1365 670 -1340
rect 610 -1405 620 -1365
rect 660 -1405 670 -1365
rect 610 -1435 670 -1405
rect 610 -1475 620 -1435
rect 660 -1475 670 -1435
rect 610 -1505 670 -1475
rect 610 -1545 620 -1505
rect 660 -1545 670 -1505
rect 610 -1575 670 -1545
rect 610 -1615 620 -1575
rect 660 -1615 670 -1575
rect 610 -1640 670 -1615
rect 610 -1680 620 -1640
rect 660 -1680 670 -1640
rect 610 -1700 670 -1680
rect 610 -1740 620 -1700
rect 660 -1740 670 -1700
rect 610 -1765 670 -1740
rect 610 -1805 620 -1765
rect 660 -1805 670 -1765
rect 610 -1835 670 -1805
rect 610 -1875 620 -1835
rect 660 -1875 670 -1835
rect 610 -1905 670 -1875
rect 610 -1945 620 -1905
rect 660 -1945 670 -1905
rect 610 -1975 670 -1945
rect 610 -2015 620 -1975
rect 660 -2015 670 -1975
rect 610 -2040 670 -2015
rect 610 -2080 620 -2040
rect 660 -2080 670 -2040
rect 610 -2100 670 -2080
rect 610 -2140 620 -2100
rect 660 -2140 670 -2100
rect 610 -2165 670 -2140
rect 610 -2205 620 -2165
rect 660 -2205 670 -2165
rect 610 -2235 670 -2205
rect 610 -2275 620 -2235
rect 660 -2275 670 -2235
rect 610 -2305 670 -2275
rect 610 -2345 620 -2305
rect 660 -2345 670 -2305
rect 610 -2375 670 -2345
rect 610 -2415 620 -2375
rect 660 -2415 670 -2375
rect 610 -2440 670 -2415
rect 610 -2480 620 -2440
rect 660 -2480 670 -2440
rect 610 -2500 670 -2480
rect 610 -2540 620 -2500
rect 660 -2540 670 -2500
rect 610 -2565 670 -2540
rect 610 -2605 620 -2565
rect 660 -2605 670 -2565
rect 610 -2635 670 -2605
rect 610 -2675 620 -2635
rect 660 -2675 670 -2635
rect 610 -2705 670 -2675
rect 610 -2745 620 -2705
rect 660 -2745 670 -2705
rect 610 -2775 670 -2745
rect 610 -2815 620 -2775
rect 660 -2815 670 -2775
rect 610 -2840 670 -2815
rect 610 -2880 620 -2840
rect 660 -2880 670 -2840
rect 610 -2900 670 -2880
rect 610 -2940 620 -2900
rect 660 -2940 670 -2900
rect 610 -2965 670 -2940
rect 610 -3005 620 -2965
rect 660 -3005 670 -2965
rect 610 -3035 670 -3005
rect 610 -3075 620 -3035
rect 660 -3075 670 -3035
rect 610 -3105 670 -3075
rect 610 -3145 620 -3105
rect 660 -3145 670 -3105
rect 610 -3175 670 -3145
rect 610 -3215 620 -3175
rect 660 -3215 670 -3175
rect 610 -3240 670 -3215
rect 610 -3280 620 -3240
rect 660 -3280 670 -3240
rect 610 -3300 670 -3280
rect 610 -3340 620 -3300
rect 660 -3340 670 -3300
rect 610 -3365 670 -3340
rect 610 -3405 620 -3365
rect 660 -3405 670 -3365
rect 610 -3435 670 -3405
rect 610 -3475 620 -3435
rect 660 -3475 670 -3435
rect 610 -3505 670 -3475
rect 610 -3545 620 -3505
rect 660 -3545 670 -3505
rect 610 -3575 670 -3545
rect 610 -3615 620 -3575
rect 660 -3615 670 -3575
rect 610 -3640 670 -3615
rect 610 -3680 620 -3640
rect 660 -3680 670 -3640
rect 610 -3700 670 -3680
rect 610 -3740 620 -3700
rect 660 -3740 670 -3700
rect 610 -3765 670 -3740
rect 610 -3805 620 -3765
rect 660 -3805 670 -3765
rect 610 -3835 670 -3805
rect 610 -3875 620 -3835
rect 660 -3875 670 -3835
rect 610 -3905 670 -3875
rect 610 -3945 620 -3905
rect 660 -3945 670 -3905
rect 610 -3975 670 -3945
rect 610 -4015 620 -3975
rect 660 -4015 670 -3975
rect 610 -4040 670 -4015
rect 610 -4080 620 -4040
rect 660 -4080 670 -4040
rect 610 -4100 670 -4080
rect 610 -4140 620 -4100
rect 660 -4140 670 -4100
rect 610 -4165 670 -4140
rect 610 -4205 620 -4165
rect 660 -4205 670 -4165
rect 610 -4235 670 -4205
rect 610 -4275 620 -4235
rect 660 -4275 670 -4235
rect 610 -4305 670 -4275
rect 610 -4345 620 -4305
rect 660 -4345 670 -4305
rect 610 -4375 670 -4345
rect 610 -4415 620 -4375
rect 660 -4415 670 -4375
rect 610 -4440 670 -4415
rect 610 -4480 620 -4440
rect 660 -4480 670 -4440
rect 610 -4490 670 -4480
rect 960 -1300 1020 -1290
rect 960 -1340 970 -1300
rect 1010 -1340 1020 -1300
rect 960 -1365 1020 -1340
rect 960 -1405 970 -1365
rect 1010 -1405 1020 -1365
rect 960 -1435 1020 -1405
rect 960 -1475 970 -1435
rect 1010 -1475 1020 -1435
rect 960 -1505 1020 -1475
rect 960 -1545 970 -1505
rect 1010 -1545 1020 -1505
rect 960 -1575 1020 -1545
rect 960 -1615 970 -1575
rect 1010 -1615 1020 -1575
rect 960 -1640 1020 -1615
rect 960 -1680 970 -1640
rect 1010 -1680 1020 -1640
rect 960 -1700 1020 -1680
rect 960 -1740 970 -1700
rect 1010 -1740 1020 -1700
rect 960 -1765 1020 -1740
rect 960 -1805 970 -1765
rect 1010 -1805 1020 -1765
rect 960 -1835 1020 -1805
rect 960 -1875 970 -1835
rect 1010 -1875 1020 -1835
rect 960 -1905 1020 -1875
rect 960 -1945 970 -1905
rect 1010 -1945 1020 -1905
rect 960 -1975 1020 -1945
rect 960 -2015 970 -1975
rect 1010 -2015 1020 -1975
rect 960 -2040 1020 -2015
rect 960 -2080 970 -2040
rect 1010 -2080 1020 -2040
rect 960 -2100 1020 -2080
rect 960 -2140 970 -2100
rect 1010 -2140 1020 -2100
rect 960 -2165 1020 -2140
rect 960 -2205 970 -2165
rect 1010 -2205 1020 -2165
rect 960 -2235 1020 -2205
rect 960 -2275 970 -2235
rect 1010 -2275 1020 -2235
rect 960 -2305 1020 -2275
rect 960 -2345 970 -2305
rect 1010 -2345 1020 -2305
rect 960 -2375 1020 -2345
rect 960 -2415 970 -2375
rect 1010 -2415 1020 -2375
rect 960 -2440 1020 -2415
rect 960 -2480 970 -2440
rect 1010 -2480 1020 -2440
rect 960 -2500 1020 -2480
rect 960 -2540 970 -2500
rect 1010 -2540 1020 -2500
rect 960 -2565 1020 -2540
rect 960 -2605 970 -2565
rect 1010 -2605 1020 -2565
rect 960 -2635 1020 -2605
rect 960 -2675 970 -2635
rect 1010 -2675 1020 -2635
rect 960 -2705 1020 -2675
rect 960 -2745 970 -2705
rect 1010 -2745 1020 -2705
rect 960 -2775 1020 -2745
rect 960 -2815 970 -2775
rect 1010 -2815 1020 -2775
rect 960 -2840 1020 -2815
rect 960 -2880 970 -2840
rect 1010 -2880 1020 -2840
rect 960 -2900 1020 -2880
rect 960 -2940 970 -2900
rect 1010 -2940 1020 -2900
rect 960 -2965 1020 -2940
rect 960 -3005 970 -2965
rect 1010 -3005 1020 -2965
rect 960 -3035 1020 -3005
rect 960 -3075 970 -3035
rect 1010 -3075 1020 -3035
rect 960 -3105 1020 -3075
rect 960 -3145 970 -3105
rect 1010 -3145 1020 -3105
rect 960 -3175 1020 -3145
rect 960 -3215 970 -3175
rect 1010 -3215 1020 -3175
rect 960 -3240 1020 -3215
rect 960 -3280 970 -3240
rect 1010 -3280 1020 -3240
rect 960 -3300 1020 -3280
rect 960 -3340 970 -3300
rect 1010 -3340 1020 -3300
rect 960 -3365 1020 -3340
rect 960 -3405 970 -3365
rect 1010 -3405 1020 -3365
rect 960 -3435 1020 -3405
rect 960 -3475 970 -3435
rect 1010 -3475 1020 -3435
rect 960 -3505 1020 -3475
rect 960 -3545 970 -3505
rect 1010 -3545 1020 -3505
rect 960 -3575 1020 -3545
rect 960 -3615 970 -3575
rect 1010 -3615 1020 -3575
rect 960 -3640 1020 -3615
rect 960 -3680 970 -3640
rect 1010 -3680 1020 -3640
rect 960 -3700 1020 -3680
rect 960 -3740 970 -3700
rect 1010 -3740 1020 -3700
rect 960 -3765 1020 -3740
rect 960 -3805 970 -3765
rect 1010 -3805 1020 -3765
rect 960 -3835 1020 -3805
rect 960 -3875 970 -3835
rect 1010 -3875 1020 -3835
rect 960 -3905 1020 -3875
rect 960 -3945 970 -3905
rect 1010 -3945 1020 -3905
rect 960 -3975 1020 -3945
rect 960 -4015 970 -3975
rect 1010 -4015 1020 -3975
rect 960 -4040 1020 -4015
rect 960 -4080 970 -4040
rect 1010 -4080 1020 -4040
rect 960 -4100 1020 -4080
rect 960 -4140 970 -4100
rect 1010 -4140 1020 -4100
rect 960 -4165 1020 -4140
rect 960 -4205 970 -4165
rect 1010 -4205 1020 -4165
rect 960 -4235 1020 -4205
rect 960 -4275 970 -4235
rect 1010 -4275 1020 -4235
rect 960 -4305 1020 -4275
rect 960 -4345 970 -4305
rect 1010 -4345 1020 -4305
rect 960 -4375 1020 -4345
rect 960 -4415 970 -4375
rect 1010 -4415 1020 -4375
rect 960 -4440 1020 -4415
rect 960 -4480 970 -4440
rect 1010 -4480 1020 -4440
rect 960 -4490 1020 -4480
rect 1310 -1300 1370 -1290
rect 1310 -1340 1320 -1300
rect 1360 -1340 1370 -1300
rect 1310 -1365 1370 -1340
rect 1310 -1405 1320 -1365
rect 1360 -1405 1370 -1365
rect 1310 -1435 1370 -1405
rect 1310 -1475 1320 -1435
rect 1360 -1475 1370 -1435
rect 1310 -1505 1370 -1475
rect 1310 -1545 1320 -1505
rect 1360 -1545 1370 -1505
rect 1310 -1575 1370 -1545
rect 1310 -1615 1320 -1575
rect 1360 -1615 1370 -1575
rect 1310 -1640 1370 -1615
rect 1310 -1680 1320 -1640
rect 1360 -1680 1370 -1640
rect 1310 -1700 1370 -1680
rect 1310 -1740 1320 -1700
rect 1360 -1740 1370 -1700
rect 1310 -1765 1370 -1740
rect 1310 -1805 1320 -1765
rect 1360 -1805 1370 -1765
rect 1310 -1835 1370 -1805
rect 1310 -1875 1320 -1835
rect 1360 -1875 1370 -1835
rect 1310 -1905 1370 -1875
rect 1310 -1945 1320 -1905
rect 1360 -1945 1370 -1905
rect 1310 -1975 1370 -1945
rect 1310 -2015 1320 -1975
rect 1360 -2015 1370 -1975
rect 1310 -2040 1370 -2015
rect 1310 -2080 1320 -2040
rect 1360 -2080 1370 -2040
rect 1310 -2100 1370 -2080
rect 1310 -2140 1320 -2100
rect 1360 -2140 1370 -2100
rect 1310 -2165 1370 -2140
rect 1310 -2205 1320 -2165
rect 1360 -2205 1370 -2165
rect 1310 -2235 1370 -2205
rect 1310 -2275 1320 -2235
rect 1360 -2275 1370 -2235
rect 1310 -2305 1370 -2275
rect 1310 -2345 1320 -2305
rect 1360 -2345 1370 -2305
rect 1310 -2375 1370 -2345
rect 1310 -2415 1320 -2375
rect 1360 -2415 1370 -2375
rect 1310 -2440 1370 -2415
rect 1310 -2480 1320 -2440
rect 1360 -2480 1370 -2440
rect 1310 -2500 1370 -2480
rect 1310 -2540 1320 -2500
rect 1360 -2540 1370 -2500
rect 1310 -2565 1370 -2540
rect 1310 -2605 1320 -2565
rect 1360 -2605 1370 -2565
rect 1310 -2635 1370 -2605
rect 1310 -2675 1320 -2635
rect 1360 -2675 1370 -2635
rect 1310 -2705 1370 -2675
rect 1310 -2745 1320 -2705
rect 1360 -2745 1370 -2705
rect 1310 -2775 1370 -2745
rect 1310 -2815 1320 -2775
rect 1360 -2815 1370 -2775
rect 1310 -2840 1370 -2815
rect 1310 -2880 1320 -2840
rect 1360 -2880 1370 -2840
rect 1310 -2900 1370 -2880
rect 1310 -2940 1320 -2900
rect 1360 -2940 1370 -2900
rect 1310 -2965 1370 -2940
rect 1310 -3005 1320 -2965
rect 1360 -3005 1370 -2965
rect 1310 -3035 1370 -3005
rect 1310 -3075 1320 -3035
rect 1360 -3075 1370 -3035
rect 1310 -3105 1370 -3075
rect 1310 -3145 1320 -3105
rect 1360 -3145 1370 -3105
rect 1310 -3175 1370 -3145
rect 1310 -3215 1320 -3175
rect 1360 -3215 1370 -3175
rect 1310 -3240 1370 -3215
rect 1310 -3280 1320 -3240
rect 1360 -3280 1370 -3240
rect 1310 -3300 1370 -3280
rect 1310 -3340 1320 -3300
rect 1360 -3340 1370 -3300
rect 1310 -3365 1370 -3340
rect 1310 -3405 1320 -3365
rect 1360 -3405 1370 -3365
rect 1310 -3435 1370 -3405
rect 1310 -3475 1320 -3435
rect 1360 -3475 1370 -3435
rect 1310 -3505 1370 -3475
rect 1310 -3545 1320 -3505
rect 1360 -3545 1370 -3505
rect 1310 -3575 1370 -3545
rect 1310 -3615 1320 -3575
rect 1360 -3615 1370 -3575
rect 1310 -3640 1370 -3615
rect 1310 -3680 1320 -3640
rect 1360 -3680 1370 -3640
rect 1310 -3700 1370 -3680
rect 1310 -3740 1320 -3700
rect 1360 -3740 1370 -3700
rect 1310 -3765 1370 -3740
rect 1310 -3805 1320 -3765
rect 1360 -3805 1370 -3765
rect 1310 -3835 1370 -3805
rect 1310 -3875 1320 -3835
rect 1360 -3875 1370 -3835
rect 1310 -3905 1370 -3875
rect 1310 -3945 1320 -3905
rect 1360 -3945 1370 -3905
rect 1310 -3975 1370 -3945
rect 1310 -4015 1320 -3975
rect 1360 -4015 1370 -3975
rect 1310 -4040 1370 -4015
rect 1310 -4080 1320 -4040
rect 1360 -4080 1370 -4040
rect 1310 -4100 1370 -4080
rect 1310 -4140 1320 -4100
rect 1360 -4140 1370 -4100
rect 1310 -4165 1370 -4140
rect 1310 -4205 1320 -4165
rect 1360 -4205 1370 -4165
rect 1310 -4235 1370 -4205
rect 1310 -4275 1320 -4235
rect 1360 -4275 1370 -4235
rect 1310 -4305 1370 -4275
rect 1310 -4345 1320 -4305
rect 1360 -4345 1370 -4305
rect 1310 -4375 1370 -4345
rect 1310 -4415 1320 -4375
rect 1360 -4415 1370 -4375
rect 1310 -4440 1370 -4415
rect 1310 -4480 1320 -4440
rect 1360 -4480 1370 -4440
rect 1310 -4490 1370 -4480
rect 1660 -1300 1720 -1290
rect 1660 -1340 1670 -1300
rect 1710 -1340 1720 -1300
rect 1660 -1365 1720 -1340
rect 1660 -1405 1670 -1365
rect 1710 -1405 1720 -1365
rect 1660 -1435 1720 -1405
rect 1660 -1475 1670 -1435
rect 1710 -1475 1720 -1435
rect 1660 -1505 1720 -1475
rect 1660 -1545 1670 -1505
rect 1710 -1545 1720 -1505
rect 1660 -1575 1720 -1545
rect 1660 -1615 1670 -1575
rect 1710 -1615 1720 -1575
rect 1660 -1640 1720 -1615
rect 1660 -1680 1670 -1640
rect 1710 -1680 1720 -1640
rect 1660 -1700 1720 -1680
rect 1660 -1740 1670 -1700
rect 1710 -1740 1720 -1700
rect 1660 -1765 1720 -1740
rect 1660 -1805 1670 -1765
rect 1710 -1805 1720 -1765
rect 1660 -1835 1720 -1805
rect 1660 -1875 1670 -1835
rect 1710 -1875 1720 -1835
rect 1660 -1905 1720 -1875
rect 1660 -1945 1670 -1905
rect 1710 -1945 1720 -1905
rect 1660 -1975 1720 -1945
rect 1660 -2015 1670 -1975
rect 1710 -2015 1720 -1975
rect 1660 -2040 1720 -2015
rect 1660 -2080 1670 -2040
rect 1710 -2080 1720 -2040
rect 1660 -2100 1720 -2080
rect 1660 -2140 1670 -2100
rect 1710 -2140 1720 -2100
rect 1660 -2165 1720 -2140
rect 1660 -2205 1670 -2165
rect 1710 -2205 1720 -2165
rect 1660 -2235 1720 -2205
rect 1660 -2275 1670 -2235
rect 1710 -2275 1720 -2235
rect 1660 -2305 1720 -2275
rect 1660 -2345 1670 -2305
rect 1710 -2345 1720 -2305
rect 1660 -2375 1720 -2345
rect 1660 -2415 1670 -2375
rect 1710 -2415 1720 -2375
rect 1660 -2440 1720 -2415
rect 1660 -2480 1670 -2440
rect 1710 -2480 1720 -2440
rect 1660 -2500 1720 -2480
rect 1660 -2540 1670 -2500
rect 1710 -2540 1720 -2500
rect 1660 -2565 1720 -2540
rect 1660 -2605 1670 -2565
rect 1710 -2605 1720 -2565
rect 1660 -2635 1720 -2605
rect 1660 -2675 1670 -2635
rect 1710 -2675 1720 -2635
rect 1660 -2705 1720 -2675
rect 1660 -2745 1670 -2705
rect 1710 -2745 1720 -2705
rect 1660 -2775 1720 -2745
rect 1660 -2815 1670 -2775
rect 1710 -2815 1720 -2775
rect 1660 -2840 1720 -2815
rect 1660 -2880 1670 -2840
rect 1710 -2880 1720 -2840
rect 1660 -2900 1720 -2880
rect 1660 -2940 1670 -2900
rect 1710 -2940 1720 -2900
rect 1660 -2965 1720 -2940
rect 1660 -3005 1670 -2965
rect 1710 -3005 1720 -2965
rect 1660 -3035 1720 -3005
rect 1660 -3075 1670 -3035
rect 1710 -3075 1720 -3035
rect 1660 -3105 1720 -3075
rect 1660 -3145 1670 -3105
rect 1710 -3145 1720 -3105
rect 1660 -3175 1720 -3145
rect 1660 -3215 1670 -3175
rect 1710 -3215 1720 -3175
rect 1660 -3240 1720 -3215
rect 1660 -3280 1670 -3240
rect 1710 -3280 1720 -3240
rect 1660 -3300 1720 -3280
rect 1660 -3340 1670 -3300
rect 1710 -3340 1720 -3300
rect 1660 -3365 1720 -3340
rect 1660 -3405 1670 -3365
rect 1710 -3405 1720 -3365
rect 1660 -3435 1720 -3405
rect 1660 -3475 1670 -3435
rect 1710 -3475 1720 -3435
rect 1660 -3505 1720 -3475
rect 1660 -3545 1670 -3505
rect 1710 -3545 1720 -3505
rect 1660 -3575 1720 -3545
rect 1660 -3615 1670 -3575
rect 1710 -3615 1720 -3575
rect 1660 -3640 1720 -3615
rect 1660 -3680 1670 -3640
rect 1710 -3680 1720 -3640
rect 1660 -3700 1720 -3680
rect 1660 -3740 1670 -3700
rect 1710 -3740 1720 -3700
rect 1660 -3765 1720 -3740
rect 1660 -3805 1670 -3765
rect 1710 -3805 1720 -3765
rect 1660 -3835 1720 -3805
rect 1660 -3875 1670 -3835
rect 1710 -3875 1720 -3835
rect 1660 -3905 1720 -3875
rect 1660 -3945 1670 -3905
rect 1710 -3945 1720 -3905
rect 1660 -3975 1720 -3945
rect 1660 -4015 1670 -3975
rect 1710 -4015 1720 -3975
rect 1660 -4040 1720 -4015
rect 1660 -4080 1670 -4040
rect 1710 -4080 1720 -4040
rect 1660 -4100 1720 -4080
rect 1660 -4140 1670 -4100
rect 1710 -4140 1720 -4100
rect 1660 -4165 1720 -4140
rect 1660 -4205 1670 -4165
rect 1710 -4205 1720 -4165
rect 1660 -4235 1720 -4205
rect 1660 -4275 1670 -4235
rect 1710 -4275 1720 -4235
rect 1660 -4305 1720 -4275
rect 1660 -4345 1670 -4305
rect 1710 -4345 1720 -4305
rect 1660 -4375 1720 -4345
rect 1660 -4415 1670 -4375
rect 1710 -4415 1720 -4375
rect 1660 -4440 1720 -4415
rect 1660 -4480 1670 -4440
rect 1710 -4480 1720 -4440
rect 1660 -4490 1720 -4480
rect 2010 -1300 2070 -1290
rect 2010 -1340 2020 -1300
rect 2060 -1340 2070 -1300
rect 2010 -1365 2070 -1340
rect 2010 -1405 2020 -1365
rect 2060 -1405 2070 -1365
rect 2010 -1435 2070 -1405
rect 2010 -1475 2020 -1435
rect 2060 -1475 2070 -1435
rect 2010 -1505 2070 -1475
rect 2010 -1545 2020 -1505
rect 2060 -1545 2070 -1505
rect 2010 -1575 2070 -1545
rect 2010 -1615 2020 -1575
rect 2060 -1615 2070 -1575
rect 2010 -1640 2070 -1615
rect 2010 -1680 2020 -1640
rect 2060 -1680 2070 -1640
rect 2010 -1700 2070 -1680
rect 2010 -1740 2020 -1700
rect 2060 -1740 2070 -1700
rect 2010 -1765 2070 -1740
rect 2010 -1805 2020 -1765
rect 2060 -1805 2070 -1765
rect 2010 -1835 2070 -1805
rect 2010 -1875 2020 -1835
rect 2060 -1875 2070 -1835
rect 2010 -1905 2070 -1875
rect 2010 -1945 2020 -1905
rect 2060 -1945 2070 -1905
rect 2010 -1975 2070 -1945
rect 2010 -2015 2020 -1975
rect 2060 -2015 2070 -1975
rect 2010 -2040 2070 -2015
rect 2010 -2080 2020 -2040
rect 2060 -2080 2070 -2040
rect 2010 -2100 2070 -2080
rect 2010 -2140 2020 -2100
rect 2060 -2140 2070 -2100
rect 2010 -2165 2070 -2140
rect 2010 -2205 2020 -2165
rect 2060 -2205 2070 -2165
rect 2010 -2235 2070 -2205
rect 2010 -2275 2020 -2235
rect 2060 -2275 2070 -2235
rect 2010 -2305 2070 -2275
rect 2010 -2345 2020 -2305
rect 2060 -2345 2070 -2305
rect 2010 -2375 2070 -2345
rect 2010 -2415 2020 -2375
rect 2060 -2415 2070 -2375
rect 2010 -2440 2070 -2415
rect 2010 -2480 2020 -2440
rect 2060 -2480 2070 -2440
rect 2010 -2500 2070 -2480
rect 2010 -2540 2020 -2500
rect 2060 -2540 2070 -2500
rect 2010 -2565 2070 -2540
rect 2010 -2605 2020 -2565
rect 2060 -2605 2070 -2565
rect 2010 -2635 2070 -2605
rect 2010 -2675 2020 -2635
rect 2060 -2675 2070 -2635
rect 2010 -2705 2070 -2675
rect 2010 -2745 2020 -2705
rect 2060 -2745 2070 -2705
rect 2010 -2775 2070 -2745
rect 2010 -2815 2020 -2775
rect 2060 -2815 2070 -2775
rect 2010 -2840 2070 -2815
rect 2010 -2880 2020 -2840
rect 2060 -2880 2070 -2840
rect 2010 -2900 2070 -2880
rect 2010 -2940 2020 -2900
rect 2060 -2940 2070 -2900
rect 2010 -2965 2070 -2940
rect 2010 -3005 2020 -2965
rect 2060 -3005 2070 -2965
rect 2010 -3035 2070 -3005
rect 2010 -3075 2020 -3035
rect 2060 -3075 2070 -3035
rect 2010 -3105 2070 -3075
rect 2010 -3145 2020 -3105
rect 2060 -3145 2070 -3105
rect 2010 -3175 2070 -3145
rect 2010 -3215 2020 -3175
rect 2060 -3215 2070 -3175
rect 2010 -3240 2070 -3215
rect 2010 -3280 2020 -3240
rect 2060 -3280 2070 -3240
rect 2010 -3300 2070 -3280
rect 2010 -3340 2020 -3300
rect 2060 -3340 2070 -3300
rect 2010 -3365 2070 -3340
rect 2010 -3405 2020 -3365
rect 2060 -3405 2070 -3365
rect 2010 -3435 2070 -3405
rect 2010 -3475 2020 -3435
rect 2060 -3475 2070 -3435
rect 2010 -3505 2070 -3475
rect 2010 -3545 2020 -3505
rect 2060 -3545 2070 -3505
rect 2010 -3575 2070 -3545
rect 2010 -3615 2020 -3575
rect 2060 -3615 2070 -3575
rect 2010 -3640 2070 -3615
rect 2010 -3680 2020 -3640
rect 2060 -3680 2070 -3640
rect 2010 -3700 2070 -3680
rect 2010 -3740 2020 -3700
rect 2060 -3740 2070 -3700
rect 2010 -3765 2070 -3740
rect 2010 -3805 2020 -3765
rect 2060 -3805 2070 -3765
rect 2010 -3835 2070 -3805
rect 2010 -3875 2020 -3835
rect 2060 -3875 2070 -3835
rect 2010 -3905 2070 -3875
rect 2010 -3945 2020 -3905
rect 2060 -3945 2070 -3905
rect 2010 -3975 2070 -3945
rect 2010 -4015 2020 -3975
rect 2060 -4015 2070 -3975
rect 2010 -4040 2070 -4015
rect 2010 -4080 2020 -4040
rect 2060 -4080 2070 -4040
rect 2010 -4100 2070 -4080
rect 2010 -4140 2020 -4100
rect 2060 -4140 2070 -4100
rect 2010 -4165 2070 -4140
rect 2010 -4205 2020 -4165
rect 2060 -4205 2070 -4165
rect 2010 -4235 2070 -4205
rect 2010 -4275 2020 -4235
rect 2060 -4275 2070 -4235
rect 2010 -4305 2070 -4275
rect 2010 -4345 2020 -4305
rect 2060 -4345 2070 -4305
rect 2010 -4375 2070 -4345
rect 2010 -4415 2020 -4375
rect 2060 -4415 2070 -4375
rect 2010 -4440 2070 -4415
rect 2010 -4480 2020 -4440
rect 2060 -4480 2070 -4440
rect 2010 -4490 2070 -4480
rect 2360 -1300 2420 -1290
rect 2360 -1340 2370 -1300
rect 2410 -1340 2420 -1300
rect 2360 -1365 2420 -1340
rect 2360 -1405 2370 -1365
rect 2410 -1405 2420 -1365
rect 2360 -1435 2420 -1405
rect 2360 -1475 2370 -1435
rect 2410 -1475 2420 -1435
rect 2360 -1505 2420 -1475
rect 2360 -1545 2370 -1505
rect 2410 -1545 2420 -1505
rect 2360 -1575 2420 -1545
rect 2360 -1615 2370 -1575
rect 2410 -1615 2420 -1575
rect 2360 -1640 2420 -1615
rect 2360 -1680 2370 -1640
rect 2410 -1680 2420 -1640
rect 2360 -1700 2420 -1680
rect 2360 -1740 2370 -1700
rect 2410 -1740 2420 -1700
rect 2360 -1765 2420 -1740
rect 2360 -1805 2370 -1765
rect 2410 -1805 2420 -1765
rect 2360 -1835 2420 -1805
rect 2360 -1875 2370 -1835
rect 2410 -1875 2420 -1835
rect 2360 -1905 2420 -1875
rect 2360 -1945 2370 -1905
rect 2410 -1945 2420 -1905
rect 2360 -1975 2420 -1945
rect 2360 -2015 2370 -1975
rect 2410 -2015 2420 -1975
rect 2360 -2040 2420 -2015
rect 2360 -2080 2370 -2040
rect 2410 -2080 2420 -2040
rect 2360 -2100 2420 -2080
rect 2360 -2140 2370 -2100
rect 2410 -2140 2420 -2100
rect 2360 -2165 2420 -2140
rect 2360 -2205 2370 -2165
rect 2410 -2205 2420 -2165
rect 2360 -2235 2420 -2205
rect 2360 -2275 2370 -2235
rect 2410 -2275 2420 -2235
rect 2360 -2305 2420 -2275
rect 2360 -2345 2370 -2305
rect 2410 -2345 2420 -2305
rect 2360 -2375 2420 -2345
rect 2360 -2415 2370 -2375
rect 2410 -2415 2420 -2375
rect 2360 -2440 2420 -2415
rect 2360 -2480 2370 -2440
rect 2410 -2480 2420 -2440
rect 2360 -2500 2420 -2480
rect 2360 -2540 2370 -2500
rect 2410 -2540 2420 -2500
rect 2360 -2565 2420 -2540
rect 2360 -2605 2370 -2565
rect 2410 -2605 2420 -2565
rect 2360 -2635 2420 -2605
rect 2360 -2675 2370 -2635
rect 2410 -2675 2420 -2635
rect 2360 -2705 2420 -2675
rect 2360 -2745 2370 -2705
rect 2410 -2745 2420 -2705
rect 2360 -2775 2420 -2745
rect 2360 -2815 2370 -2775
rect 2410 -2815 2420 -2775
rect 2360 -2840 2420 -2815
rect 2360 -2880 2370 -2840
rect 2410 -2880 2420 -2840
rect 2360 -2900 2420 -2880
rect 2360 -2940 2370 -2900
rect 2410 -2940 2420 -2900
rect 2360 -2965 2420 -2940
rect 2360 -3005 2370 -2965
rect 2410 -3005 2420 -2965
rect 2360 -3035 2420 -3005
rect 2360 -3075 2370 -3035
rect 2410 -3075 2420 -3035
rect 2360 -3105 2420 -3075
rect 2360 -3145 2370 -3105
rect 2410 -3145 2420 -3105
rect 2360 -3175 2420 -3145
rect 2360 -3215 2370 -3175
rect 2410 -3215 2420 -3175
rect 2360 -3240 2420 -3215
rect 2360 -3280 2370 -3240
rect 2410 -3280 2420 -3240
rect 2360 -3300 2420 -3280
rect 2360 -3340 2370 -3300
rect 2410 -3340 2420 -3300
rect 2360 -3365 2420 -3340
rect 2360 -3405 2370 -3365
rect 2410 -3405 2420 -3365
rect 2360 -3435 2420 -3405
rect 2360 -3475 2370 -3435
rect 2410 -3475 2420 -3435
rect 2360 -3505 2420 -3475
rect 2360 -3545 2370 -3505
rect 2410 -3545 2420 -3505
rect 2360 -3575 2420 -3545
rect 2360 -3615 2370 -3575
rect 2410 -3615 2420 -3575
rect 2360 -3640 2420 -3615
rect 2360 -3680 2370 -3640
rect 2410 -3680 2420 -3640
rect 2360 -3700 2420 -3680
rect 2360 -3740 2370 -3700
rect 2410 -3740 2420 -3700
rect 2360 -3765 2420 -3740
rect 2360 -3805 2370 -3765
rect 2410 -3805 2420 -3765
rect 2360 -3835 2420 -3805
rect 2360 -3875 2370 -3835
rect 2410 -3875 2420 -3835
rect 2360 -3905 2420 -3875
rect 2360 -3945 2370 -3905
rect 2410 -3945 2420 -3905
rect 2360 -3975 2420 -3945
rect 2360 -4015 2370 -3975
rect 2410 -4015 2420 -3975
rect 2360 -4040 2420 -4015
rect 2360 -4080 2370 -4040
rect 2410 -4080 2420 -4040
rect 2360 -4100 2420 -4080
rect 2360 -4140 2370 -4100
rect 2410 -4140 2420 -4100
rect 2360 -4165 2420 -4140
rect 2360 -4205 2370 -4165
rect 2410 -4205 2420 -4165
rect 2360 -4235 2420 -4205
rect 2360 -4275 2370 -4235
rect 2410 -4275 2420 -4235
rect 2360 -4305 2420 -4275
rect 2360 -4345 2370 -4305
rect 2410 -4345 2420 -4305
rect 2360 -4375 2420 -4345
rect 2360 -4415 2370 -4375
rect 2410 -4415 2420 -4375
rect 2360 -4440 2420 -4415
rect 2360 -4480 2370 -4440
rect 2410 -4480 2420 -4440
rect 2360 -4490 2420 -4480
rect 2710 -1300 2770 -1290
rect 2710 -1340 2720 -1300
rect 2760 -1340 2770 -1300
rect 2710 -1365 2770 -1340
rect 2710 -1405 2720 -1365
rect 2760 -1405 2770 -1365
rect 2710 -1435 2770 -1405
rect 2710 -1475 2720 -1435
rect 2760 -1475 2770 -1435
rect 2710 -1505 2770 -1475
rect 2710 -1545 2720 -1505
rect 2760 -1545 2770 -1505
rect 2710 -1575 2770 -1545
rect 2710 -1615 2720 -1575
rect 2760 -1615 2770 -1575
rect 2710 -1640 2770 -1615
rect 2710 -1680 2720 -1640
rect 2760 -1680 2770 -1640
rect 2710 -1700 2770 -1680
rect 2710 -1740 2720 -1700
rect 2760 -1740 2770 -1700
rect 2710 -1765 2770 -1740
rect 2710 -1805 2720 -1765
rect 2760 -1805 2770 -1765
rect 2710 -1835 2770 -1805
rect 2710 -1875 2720 -1835
rect 2760 -1875 2770 -1835
rect 2710 -1905 2770 -1875
rect 2710 -1945 2720 -1905
rect 2760 -1945 2770 -1905
rect 2710 -1975 2770 -1945
rect 2710 -2015 2720 -1975
rect 2760 -2015 2770 -1975
rect 2710 -2040 2770 -2015
rect 2710 -2080 2720 -2040
rect 2760 -2080 2770 -2040
rect 2710 -2100 2770 -2080
rect 2710 -2140 2720 -2100
rect 2760 -2140 2770 -2100
rect 2710 -2165 2770 -2140
rect 2710 -2205 2720 -2165
rect 2760 -2205 2770 -2165
rect 2710 -2235 2770 -2205
rect 2710 -2275 2720 -2235
rect 2760 -2275 2770 -2235
rect 2710 -2305 2770 -2275
rect 2710 -2345 2720 -2305
rect 2760 -2345 2770 -2305
rect 2710 -2375 2770 -2345
rect 2710 -2415 2720 -2375
rect 2760 -2415 2770 -2375
rect 2710 -2440 2770 -2415
rect 2710 -2480 2720 -2440
rect 2760 -2480 2770 -2440
rect 2710 -2500 2770 -2480
rect 2710 -2540 2720 -2500
rect 2760 -2540 2770 -2500
rect 2710 -2565 2770 -2540
rect 2710 -2605 2720 -2565
rect 2760 -2605 2770 -2565
rect 2710 -2635 2770 -2605
rect 2710 -2675 2720 -2635
rect 2760 -2675 2770 -2635
rect 2710 -2705 2770 -2675
rect 2710 -2745 2720 -2705
rect 2760 -2745 2770 -2705
rect 2710 -2775 2770 -2745
rect 2710 -2815 2720 -2775
rect 2760 -2815 2770 -2775
rect 2710 -2840 2770 -2815
rect 2710 -2880 2720 -2840
rect 2760 -2880 2770 -2840
rect 2710 -2900 2770 -2880
rect 2710 -2940 2720 -2900
rect 2760 -2940 2770 -2900
rect 2710 -2965 2770 -2940
rect 2710 -3005 2720 -2965
rect 2760 -3005 2770 -2965
rect 2710 -3035 2770 -3005
rect 2710 -3075 2720 -3035
rect 2760 -3075 2770 -3035
rect 2710 -3105 2770 -3075
rect 2710 -3145 2720 -3105
rect 2760 -3145 2770 -3105
rect 2710 -3175 2770 -3145
rect 2710 -3215 2720 -3175
rect 2760 -3215 2770 -3175
rect 2710 -3240 2770 -3215
rect 2710 -3280 2720 -3240
rect 2760 -3280 2770 -3240
rect 2710 -3300 2770 -3280
rect 2710 -3340 2720 -3300
rect 2760 -3340 2770 -3300
rect 2710 -3365 2770 -3340
rect 2710 -3405 2720 -3365
rect 2760 -3405 2770 -3365
rect 2710 -3435 2770 -3405
rect 2710 -3475 2720 -3435
rect 2760 -3475 2770 -3435
rect 2710 -3505 2770 -3475
rect 2710 -3545 2720 -3505
rect 2760 -3545 2770 -3505
rect 2710 -3575 2770 -3545
rect 2710 -3615 2720 -3575
rect 2760 -3615 2770 -3575
rect 2710 -3640 2770 -3615
rect 2710 -3680 2720 -3640
rect 2760 -3680 2770 -3640
rect 2710 -3700 2770 -3680
rect 2710 -3740 2720 -3700
rect 2760 -3740 2770 -3700
rect 2710 -3765 2770 -3740
rect 2710 -3805 2720 -3765
rect 2760 -3805 2770 -3765
rect 2710 -3835 2770 -3805
rect 2710 -3875 2720 -3835
rect 2760 -3875 2770 -3835
rect 2710 -3905 2770 -3875
rect 2710 -3945 2720 -3905
rect 2760 -3945 2770 -3905
rect 2710 -3975 2770 -3945
rect 2710 -4015 2720 -3975
rect 2760 -4015 2770 -3975
rect 2710 -4040 2770 -4015
rect 2710 -4080 2720 -4040
rect 2760 -4080 2770 -4040
rect 2710 -4100 2770 -4080
rect 2710 -4140 2720 -4100
rect 2760 -4140 2770 -4100
rect 2710 -4165 2770 -4140
rect 2710 -4205 2720 -4165
rect 2760 -4205 2770 -4165
rect 2710 -4235 2770 -4205
rect 2710 -4275 2720 -4235
rect 2760 -4275 2770 -4235
rect 2710 -4305 2770 -4275
rect 2710 -4345 2720 -4305
rect 2760 -4345 2770 -4305
rect 2710 -4375 2770 -4345
rect 2710 -4415 2720 -4375
rect 2760 -4415 2770 -4375
rect 2710 -4440 2770 -4415
rect 2710 -4480 2720 -4440
rect 2760 -4480 2770 -4440
rect 2710 -4490 2770 -4480
rect 3060 -1300 3120 -1290
rect 3060 -1340 3070 -1300
rect 3110 -1340 3120 -1300
rect 3060 -1365 3120 -1340
rect 3060 -1405 3070 -1365
rect 3110 -1405 3120 -1365
rect 3060 -1435 3120 -1405
rect 3060 -1475 3070 -1435
rect 3110 -1475 3120 -1435
rect 3060 -1505 3120 -1475
rect 3060 -1545 3070 -1505
rect 3110 -1545 3120 -1505
rect 3060 -1575 3120 -1545
rect 3060 -1615 3070 -1575
rect 3110 -1615 3120 -1575
rect 3060 -1640 3120 -1615
rect 3060 -1680 3070 -1640
rect 3110 -1680 3120 -1640
rect 3060 -1700 3120 -1680
rect 3060 -1740 3070 -1700
rect 3110 -1740 3120 -1700
rect 3060 -1765 3120 -1740
rect 3060 -1805 3070 -1765
rect 3110 -1805 3120 -1765
rect 3060 -1835 3120 -1805
rect 3060 -1875 3070 -1835
rect 3110 -1875 3120 -1835
rect 3060 -1905 3120 -1875
rect 3060 -1945 3070 -1905
rect 3110 -1945 3120 -1905
rect 3060 -1975 3120 -1945
rect 3060 -2015 3070 -1975
rect 3110 -2015 3120 -1975
rect 3060 -2040 3120 -2015
rect 3060 -2080 3070 -2040
rect 3110 -2080 3120 -2040
rect 3060 -2100 3120 -2080
rect 3060 -2140 3070 -2100
rect 3110 -2140 3120 -2100
rect 3060 -2165 3120 -2140
rect 3060 -2205 3070 -2165
rect 3110 -2205 3120 -2165
rect 3060 -2235 3120 -2205
rect 3060 -2275 3070 -2235
rect 3110 -2275 3120 -2235
rect 3060 -2305 3120 -2275
rect 3060 -2345 3070 -2305
rect 3110 -2345 3120 -2305
rect 3060 -2375 3120 -2345
rect 3060 -2415 3070 -2375
rect 3110 -2415 3120 -2375
rect 3060 -2440 3120 -2415
rect 3060 -2480 3070 -2440
rect 3110 -2480 3120 -2440
rect 3060 -2500 3120 -2480
rect 3060 -2540 3070 -2500
rect 3110 -2540 3120 -2500
rect 3060 -2565 3120 -2540
rect 3060 -2605 3070 -2565
rect 3110 -2605 3120 -2565
rect 3060 -2635 3120 -2605
rect 3060 -2675 3070 -2635
rect 3110 -2675 3120 -2635
rect 3060 -2705 3120 -2675
rect 3060 -2745 3070 -2705
rect 3110 -2745 3120 -2705
rect 3060 -2775 3120 -2745
rect 3060 -2815 3070 -2775
rect 3110 -2815 3120 -2775
rect 3060 -2840 3120 -2815
rect 3060 -2880 3070 -2840
rect 3110 -2880 3120 -2840
rect 3060 -2900 3120 -2880
rect 3060 -2940 3070 -2900
rect 3110 -2940 3120 -2900
rect 3060 -2965 3120 -2940
rect 3060 -3005 3070 -2965
rect 3110 -3005 3120 -2965
rect 3060 -3035 3120 -3005
rect 3060 -3075 3070 -3035
rect 3110 -3075 3120 -3035
rect 3060 -3105 3120 -3075
rect 3060 -3145 3070 -3105
rect 3110 -3145 3120 -3105
rect 3060 -3175 3120 -3145
rect 3060 -3215 3070 -3175
rect 3110 -3215 3120 -3175
rect 3060 -3240 3120 -3215
rect 3060 -3280 3070 -3240
rect 3110 -3280 3120 -3240
rect 3060 -3300 3120 -3280
rect 3060 -3340 3070 -3300
rect 3110 -3340 3120 -3300
rect 3060 -3365 3120 -3340
rect 3060 -3405 3070 -3365
rect 3110 -3405 3120 -3365
rect 3060 -3435 3120 -3405
rect 3060 -3475 3070 -3435
rect 3110 -3475 3120 -3435
rect 3060 -3505 3120 -3475
rect 3060 -3545 3070 -3505
rect 3110 -3545 3120 -3505
rect 3060 -3575 3120 -3545
rect 3060 -3615 3070 -3575
rect 3110 -3615 3120 -3575
rect 3060 -3640 3120 -3615
rect 3060 -3680 3070 -3640
rect 3110 -3680 3120 -3640
rect 3060 -3700 3120 -3680
rect 3060 -3740 3070 -3700
rect 3110 -3740 3120 -3700
rect 3060 -3765 3120 -3740
rect 3060 -3805 3070 -3765
rect 3110 -3805 3120 -3765
rect 3060 -3835 3120 -3805
rect 3060 -3875 3070 -3835
rect 3110 -3875 3120 -3835
rect 3060 -3905 3120 -3875
rect 3060 -3945 3070 -3905
rect 3110 -3945 3120 -3905
rect 3060 -3975 3120 -3945
rect 3060 -4015 3070 -3975
rect 3110 -4015 3120 -3975
rect 3060 -4040 3120 -4015
rect 3060 -4080 3070 -4040
rect 3110 -4080 3120 -4040
rect 3060 -4100 3120 -4080
rect 3060 -4140 3070 -4100
rect 3110 -4140 3120 -4100
rect 3060 -4165 3120 -4140
rect 3060 -4205 3070 -4165
rect 3110 -4205 3120 -4165
rect 3060 -4235 3120 -4205
rect 3060 -4275 3070 -4235
rect 3110 -4275 3120 -4235
rect 3060 -4305 3120 -4275
rect 3060 -4345 3070 -4305
rect 3110 -4345 3120 -4305
rect 3060 -4375 3120 -4345
rect 3060 -4415 3070 -4375
rect 3110 -4415 3120 -4375
rect 3060 -4440 3120 -4415
rect 3060 -4480 3070 -4440
rect 3110 -4480 3120 -4440
rect 3060 -4490 3120 -4480
rect 3410 -1300 3470 -1290
rect 3410 -1340 3420 -1300
rect 3460 -1340 3470 -1300
rect 3410 -1365 3470 -1340
rect 3410 -1405 3420 -1365
rect 3460 -1405 3470 -1365
rect 3410 -1435 3470 -1405
rect 3410 -1475 3420 -1435
rect 3460 -1475 3470 -1435
rect 3410 -1505 3470 -1475
rect 3410 -1545 3420 -1505
rect 3460 -1545 3470 -1505
rect 3410 -1575 3470 -1545
rect 3410 -1615 3420 -1575
rect 3460 -1615 3470 -1575
rect 3410 -1640 3470 -1615
rect 3410 -1680 3420 -1640
rect 3460 -1680 3470 -1640
rect 3410 -1700 3470 -1680
rect 3410 -1740 3420 -1700
rect 3460 -1740 3470 -1700
rect 3410 -1765 3470 -1740
rect 3410 -1805 3420 -1765
rect 3460 -1805 3470 -1765
rect 3410 -1835 3470 -1805
rect 3410 -1875 3420 -1835
rect 3460 -1875 3470 -1835
rect 3410 -1905 3470 -1875
rect 3410 -1945 3420 -1905
rect 3460 -1945 3470 -1905
rect 3410 -1975 3470 -1945
rect 3410 -2015 3420 -1975
rect 3460 -2015 3470 -1975
rect 3410 -2040 3470 -2015
rect 3410 -2080 3420 -2040
rect 3460 -2080 3470 -2040
rect 3410 -2100 3470 -2080
rect 3410 -2140 3420 -2100
rect 3460 -2140 3470 -2100
rect 3410 -2165 3470 -2140
rect 3410 -2205 3420 -2165
rect 3460 -2205 3470 -2165
rect 3410 -2235 3470 -2205
rect 3410 -2275 3420 -2235
rect 3460 -2275 3470 -2235
rect 3410 -2305 3470 -2275
rect 3410 -2345 3420 -2305
rect 3460 -2345 3470 -2305
rect 3410 -2375 3470 -2345
rect 3410 -2415 3420 -2375
rect 3460 -2415 3470 -2375
rect 3410 -2440 3470 -2415
rect 3410 -2480 3420 -2440
rect 3460 -2480 3470 -2440
rect 3410 -2500 3470 -2480
rect 3410 -2540 3420 -2500
rect 3460 -2540 3470 -2500
rect 3410 -2565 3470 -2540
rect 3410 -2605 3420 -2565
rect 3460 -2605 3470 -2565
rect 3410 -2635 3470 -2605
rect 3410 -2675 3420 -2635
rect 3460 -2675 3470 -2635
rect 3410 -2705 3470 -2675
rect 3410 -2745 3420 -2705
rect 3460 -2745 3470 -2705
rect 3410 -2775 3470 -2745
rect 3410 -2815 3420 -2775
rect 3460 -2815 3470 -2775
rect 3410 -2840 3470 -2815
rect 3410 -2880 3420 -2840
rect 3460 -2880 3470 -2840
rect 3410 -2900 3470 -2880
rect 3410 -2940 3420 -2900
rect 3460 -2940 3470 -2900
rect 3410 -2965 3470 -2940
rect 3410 -3005 3420 -2965
rect 3460 -3005 3470 -2965
rect 3410 -3035 3470 -3005
rect 3410 -3075 3420 -3035
rect 3460 -3075 3470 -3035
rect 3410 -3105 3470 -3075
rect 3410 -3145 3420 -3105
rect 3460 -3145 3470 -3105
rect 3410 -3175 3470 -3145
rect 3410 -3215 3420 -3175
rect 3460 -3215 3470 -3175
rect 3410 -3240 3470 -3215
rect 3410 -3280 3420 -3240
rect 3460 -3280 3470 -3240
rect 3410 -3300 3470 -3280
rect 3410 -3340 3420 -3300
rect 3460 -3340 3470 -3300
rect 3410 -3365 3470 -3340
rect 3410 -3405 3420 -3365
rect 3460 -3405 3470 -3365
rect 3410 -3435 3470 -3405
rect 3410 -3475 3420 -3435
rect 3460 -3475 3470 -3435
rect 3410 -3505 3470 -3475
rect 3410 -3545 3420 -3505
rect 3460 -3545 3470 -3505
rect 3410 -3575 3470 -3545
rect 3410 -3615 3420 -3575
rect 3460 -3615 3470 -3575
rect 3410 -3640 3470 -3615
rect 3410 -3680 3420 -3640
rect 3460 -3680 3470 -3640
rect 3410 -3700 3470 -3680
rect 3410 -3740 3420 -3700
rect 3460 -3740 3470 -3700
rect 3410 -3765 3470 -3740
rect 3410 -3805 3420 -3765
rect 3460 -3805 3470 -3765
rect 3410 -3835 3470 -3805
rect 3410 -3875 3420 -3835
rect 3460 -3875 3470 -3835
rect 3410 -3905 3470 -3875
rect 3410 -3945 3420 -3905
rect 3460 -3945 3470 -3905
rect 3410 -3975 3470 -3945
rect 3410 -4015 3420 -3975
rect 3460 -4015 3470 -3975
rect 3410 -4040 3470 -4015
rect 3410 -4080 3420 -4040
rect 3460 -4080 3470 -4040
rect 3410 -4100 3470 -4080
rect 3410 -4140 3420 -4100
rect 3460 -4140 3470 -4100
rect 3410 -4165 3470 -4140
rect 3410 -4205 3420 -4165
rect 3460 -4205 3470 -4165
rect 3410 -4235 3470 -4205
rect 3410 -4275 3420 -4235
rect 3460 -4275 3470 -4235
rect 3410 -4305 3470 -4275
rect 3410 -4345 3420 -4305
rect 3460 -4345 3470 -4305
rect 3410 -4375 3470 -4345
rect 3410 -4415 3420 -4375
rect 3460 -4415 3470 -4375
rect 3410 -4440 3470 -4415
rect 3410 -4480 3420 -4440
rect 3460 -4480 3470 -4440
rect 3410 -4490 3470 -4480
rect 3760 -1300 3820 -1290
rect 3760 -1340 3770 -1300
rect 3810 -1340 3820 -1300
rect 3760 -1365 3820 -1340
rect 3760 -1405 3770 -1365
rect 3810 -1405 3820 -1365
rect 3760 -1435 3820 -1405
rect 3760 -1475 3770 -1435
rect 3810 -1475 3820 -1435
rect 3760 -1505 3820 -1475
rect 3760 -1545 3770 -1505
rect 3810 -1545 3820 -1505
rect 3760 -1575 3820 -1545
rect 3760 -1615 3770 -1575
rect 3810 -1615 3820 -1575
rect 3760 -1640 3820 -1615
rect 3760 -1680 3770 -1640
rect 3810 -1680 3820 -1640
rect 3760 -1700 3820 -1680
rect 3760 -1740 3770 -1700
rect 3810 -1740 3820 -1700
rect 3760 -1765 3820 -1740
rect 3760 -1805 3770 -1765
rect 3810 -1805 3820 -1765
rect 3760 -1835 3820 -1805
rect 3760 -1875 3770 -1835
rect 3810 -1875 3820 -1835
rect 3760 -1905 3820 -1875
rect 3760 -1945 3770 -1905
rect 3810 -1945 3820 -1905
rect 3760 -1975 3820 -1945
rect 3760 -2015 3770 -1975
rect 3810 -2015 3820 -1975
rect 3760 -2040 3820 -2015
rect 3760 -2080 3770 -2040
rect 3810 -2080 3820 -2040
rect 3760 -2100 3820 -2080
rect 3760 -2140 3770 -2100
rect 3810 -2140 3820 -2100
rect 3760 -2165 3820 -2140
rect 3760 -2205 3770 -2165
rect 3810 -2205 3820 -2165
rect 3760 -2235 3820 -2205
rect 3760 -2275 3770 -2235
rect 3810 -2275 3820 -2235
rect 3760 -2305 3820 -2275
rect 3760 -2345 3770 -2305
rect 3810 -2345 3820 -2305
rect 3760 -2375 3820 -2345
rect 3760 -2415 3770 -2375
rect 3810 -2415 3820 -2375
rect 3760 -2440 3820 -2415
rect 3760 -2480 3770 -2440
rect 3810 -2480 3820 -2440
rect 3760 -2500 3820 -2480
rect 3760 -2540 3770 -2500
rect 3810 -2540 3820 -2500
rect 3760 -2565 3820 -2540
rect 3760 -2605 3770 -2565
rect 3810 -2605 3820 -2565
rect 3760 -2635 3820 -2605
rect 3760 -2675 3770 -2635
rect 3810 -2675 3820 -2635
rect 3760 -2705 3820 -2675
rect 3760 -2745 3770 -2705
rect 3810 -2745 3820 -2705
rect 3760 -2775 3820 -2745
rect 3760 -2815 3770 -2775
rect 3810 -2815 3820 -2775
rect 3760 -2840 3820 -2815
rect 3760 -2880 3770 -2840
rect 3810 -2880 3820 -2840
rect 3760 -2900 3820 -2880
rect 3760 -2940 3770 -2900
rect 3810 -2940 3820 -2900
rect 3760 -2965 3820 -2940
rect 3760 -3005 3770 -2965
rect 3810 -3005 3820 -2965
rect 3760 -3035 3820 -3005
rect 3760 -3075 3770 -3035
rect 3810 -3075 3820 -3035
rect 3760 -3105 3820 -3075
rect 3760 -3145 3770 -3105
rect 3810 -3145 3820 -3105
rect 3760 -3175 3820 -3145
rect 3760 -3215 3770 -3175
rect 3810 -3215 3820 -3175
rect 3760 -3240 3820 -3215
rect 3760 -3280 3770 -3240
rect 3810 -3280 3820 -3240
rect 3760 -3300 3820 -3280
rect 3760 -3340 3770 -3300
rect 3810 -3340 3820 -3300
rect 3760 -3365 3820 -3340
rect 3760 -3405 3770 -3365
rect 3810 -3405 3820 -3365
rect 3760 -3435 3820 -3405
rect 3760 -3475 3770 -3435
rect 3810 -3475 3820 -3435
rect 3760 -3505 3820 -3475
rect 3760 -3545 3770 -3505
rect 3810 -3545 3820 -3505
rect 3760 -3575 3820 -3545
rect 3760 -3615 3770 -3575
rect 3810 -3615 3820 -3575
rect 3760 -3640 3820 -3615
rect 3760 -3680 3770 -3640
rect 3810 -3680 3820 -3640
rect 3760 -3700 3820 -3680
rect 3760 -3740 3770 -3700
rect 3810 -3740 3820 -3700
rect 3760 -3765 3820 -3740
rect 3760 -3805 3770 -3765
rect 3810 -3805 3820 -3765
rect 3760 -3835 3820 -3805
rect 3760 -3875 3770 -3835
rect 3810 -3875 3820 -3835
rect 3760 -3905 3820 -3875
rect 3760 -3945 3770 -3905
rect 3810 -3945 3820 -3905
rect 3760 -3975 3820 -3945
rect 3760 -4015 3770 -3975
rect 3810 -4015 3820 -3975
rect 3760 -4040 3820 -4015
rect 3760 -4080 3770 -4040
rect 3810 -4080 3820 -4040
rect 3760 -4100 3820 -4080
rect 3760 -4140 3770 -4100
rect 3810 -4140 3820 -4100
rect 3760 -4165 3820 -4140
rect 3760 -4205 3770 -4165
rect 3810 -4205 3820 -4165
rect 3760 -4235 3820 -4205
rect 3760 -4275 3770 -4235
rect 3810 -4275 3820 -4235
rect 3760 -4305 3820 -4275
rect 3760 -4345 3770 -4305
rect 3810 -4345 3820 -4305
rect 3760 -4375 3820 -4345
rect 3760 -4415 3770 -4375
rect 3810 -4415 3820 -4375
rect 3760 -4440 3820 -4415
rect 3760 -4480 3770 -4440
rect 3810 -4480 3820 -4440
rect 3760 -4490 3820 -4480
rect 4110 -1300 4170 -1290
rect 4110 -1340 4120 -1300
rect 4160 -1340 4170 -1300
rect 4110 -1365 4170 -1340
rect 4110 -1405 4120 -1365
rect 4160 -1405 4170 -1365
rect 4110 -1435 4170 -1405
rect 4110 -1475 4120 -1435
rect 4160 -1475 4170 -1435
rect 4110 -1505 4170 -1475
rect 4110 -1545 4120 -1505
rect 4160 -1545 4170 -1505
rect 4110 -1575 4170 -1545
rect 4110 -1615 4120 -1575
rect 4160 -1615 4170 -1575
rect 4110 -1640 4170 -1615
rect 4110 -1680 4120 -1640
rect 4160 -1680 4170 -1640
rect 4110 -1700 4170 -1680
rect 4110 -1740 4120 -1700
rect 4160 -1740 4170 -1700
rect 4110 -1765 4170 -1740
rect 4110 -1805 4120 -1765
rect 4160 -1805 4170 -1765
rect 4110 -1835 4170 -1805
rect 4110 -1875 4120 -1835
rect 4160 -1875 4170 -1835
rect 4110 -1905 4170 -1875
rect 4110 -1945 4120 -1905
rect 4160 -1945 4170 -1905
rect 4110 -1975 4170 -1945
rect 4110 -2015 4120 -1975
rect 4160 -2015 4170 -1975
rect 4110 -2040 4170 -2015
rect 4110 -2080 4120 -2040
rect 4160 -2080 4170 -2040
rect 4110 -2100 4170 -2080
rect 4110 -2140 4120 -2100
rect 4160 -2140 4170 -2100
rect 4110 -2165 4170 -2140
rect 4110 -2205 4120 -2165
rect 4160 -2205 4170 -2165
rect 4110 -2235 4170 -2205
rect 4110 -2275 4120 -2235
rect 4160 -2275 4170 -2235
rect 4110 -2305 4170 -2275
rect 4110 -2345 4120 -2305
rect 4160 -2345 4170 -2305
rect 4110 -2375 4170 -2345
rect 4110 -2415 4120 -2375
rect 4160 -2415 4170 -2375
rect 4110 -2440 4170 -2415
rect 4110 -2480 4120 -2440
rect 4160 -2480 4170 -2440
rect 4110 -2500 4170 -2480
rect 4110 -2540 4120 -2500
rect 4160 -2540 4170 -2500
rect 4110 -2565 4170 -2540
rect 4110 -2605 4120 -2565
rect 4160 -2605 4170 -2565
rect 4110 -2635 4170 -2605
rect 4110 -2675 4120 -2635
rect 4160 -2675 4170 -2635
rect 4110 -2705 4170 -2675
rect 4110 -2745 4120 -2705
rect 4160 -2745 4170 -2705
rect 4110 -2775 4170 -2745
rect 4110 -2815 4120 -2775
rect 4160 -2815 4170 -2775
rect 4110 -2840 4170 -2815
rect 4110 -2880 4120 -2840
rect 4160 -2880 4170 -2840
rect 4110 -2900 4170 -2880
rect 4110 -2940 4120 -2900
rect 4160 -2940 4170 -2900
rect 4110 -2965 4170 -2940
rect 4110 -3005 4120 -2965
rect 4160 -3005 4170 -2965
rect 4110 -3035 4170 -3005
rect 4110 -3075 4120 -3035
rect 4160 -3075 4170 -3035
rect 4110 -3105 4170 -3075
rect 4110 -3145 4120 -3105
rect 4160 -3145 4170 -3105
rect 4110 -3175 4170 -3145
rect 4110 -3215 4120 -3175
rect 4160 -3215 4170 -3175
rect 4110 -3240 4170 -3215
rect 4110 -3280 4120 -3240
rect 4160 -3280 4170 -3240
rect 4110 -3300 4170 -3280
rect 4110 -3340 4120 -3300
rect 4160 -3340 4170 -3300
rect 4110 -3365 4170 -3340
rect 4110 -3405 4120 -3365
rect 4160 -3405 4170 -3365
rect 4110 -3435 4170 -3405
rect 4110 -3475 4120 -3435
rect 4160 -3475 4170 -3435
rect 4110 -3505 4170 -3475
rect 4110 -3545 4120 -3505
rect 4160 -3545 4170 -3505
rect 4110 -3575 4170 -3545
rect 4110 -3615 4120 -3575
rect 4160 -3615 4170 -3575
rect 4110 -3640 4170 -3615
rect 4110 -3680 4120 -3640
rect 4160 -3680 4170 -3640
rect 4110 -3700 4170 -3680
rect 4110 -3740 4120 -3700
rect 4160 -3740 4170 -3700
rect 4110 -3765 4170 -3740
rect 4110 -3805 4120 -3765
rect 4160 -3805 4170 -3765
rect 4110 -3835 4170 -3805
rect 4110 -3875 4120 -3835
rect 4160 -3875 4170 -3835
rect 4110 -3905 4170 -3875
rect 4110 -3945 4120 -3905
rect 4160 -3945 4170 -3905
rect 4110 -3975 4170 -3945
rect 4110 -4015 4120 -3975
rect 4160 -4015 4170 -3975
rect 4110 -4040 4170 -4015
rect 4110 -4080 4120 -4040
rect 4160 -4080 4170 -4040
rect 4110 -4100 4170 -4080
rect 4110 -4140 4120 -4100
rect 4160 -4140 4170 -4100
rect 4110 -4165 4170 -4140
rect 4110 -4205 4120 -4165
rect 4160 -4205 4170 -4165
rect 4110 -4235 4170 -4205
rect 4110 -4275 4120 -4235
rect 4160 -4275 4170 -4235
rect 4110 -4305 4170 -4275
rect 4110 -4345 4120 -4305
rect 4160 -4345 4170 -4305
rect 4110 -4375 4170 -4345
rect 4110 -4415 4120 -4375
rect 4160 -4415 4170 -4375
rect 4110 -4440 4170 -4415
rect 4110 -4480 4120 -4440
rect 4160 -4480 4170 -4440
rect 4110 -4490 4170 -4480
rect 4460 -1300 4520 -1290
rect 4460 -1340 4470 -1300
rect 4510 -1340 4520 -1300
rect 4460 -1365 4520 -1340
rect 4460 -1405 4470 -1365
rect 4510 -1405 4520 -1365
rect 4460 -1435 4520 -1405
rect 4460 -1475 4470 -1435
rect 4510 -1475 4520 -1435
rect 4460 -1505 4520 -1475
rect 4460 -1545 4470 -1505
rect 4510 -1545 4520 -1505
rect 4460 -1575 4520 -1545
rect 4460 -1615 4470 -1575
rect 4510 -1615 4520 -1575
rect 4460 -1640 4520 -1615
rect 4460 -1680 4470 -1640
rect 4510 -1680 4520 -1640
rect 4460 -1700 4520 -1680
rect 4460 -1740 4470 -1700
rect 4510 -1740 4520 -1700
rect 4460 -1765 4520 -1740
rect 4460 -1805 4470 -1765
rect 4510 -1805 4520 -1765
rect 4460 -1835 4520 -1805
rect 4460 -1875 4470 -1835
rect 4510 -1875 4520 -1835
rect 4460 -1905 4520 -1875
rect 4460 -1945 4470 -1905
rect 4510 -1945 4520 -1905
rect 4460 -1975 4520 -1945
rect 4460 -2015 4470 -1975
rect 4510 -2015 4520 -1975
rect 4460 -2040 4520 -2015
rect 4460 -2080 4470 -2040
rect 4510 -2080 4520 -2040
rect 4460 -2100 4520 -2080
rect 4460 -2140 4470 -2100
rect 4510 -2140 4520 -2100
rect 4460 -2165 4520 -2140
rect 4460 -2205 4470 -2165
rect 4510 -2205 4520 -2165
rect 4460 -2235 4520 -2205
rect 4460 -2275 4470 -2235
rect 4510 -2275 4520 -2235
rect 4460 -2305 4520 -2275
rect 4460 -2345 4470 -2305
rect 4510 -2345 4520 -2305
rect 4460 -2375 4520 -2345
rect 4460 -2415 4470 -2375
rect 4510 -2415 4520 -2375
rect 4460 -2440 4520 -2415
rect 4460 -2480 4470 -2440
rect 4510 -2480 4520 -2440
rect 4460 -2500 4520 -2480
rect 4460 -2540 4470 -2500
rect 4510 -2540 4520 -2500
rect 4460 -2565 4520 -2540
rect 4460 -2605 4470 -2565
rect 4510 -2605 4520 -2565
rect 4460 -2635 4520 -2605
rect 4460 -2675 4470 -2635
rect 4510 -2675 4520 -2635
rect 4460 -2705 4520 -2675
rect 4460 -2745 4470 -2705
rect 4510 -2745 4520 -2705
rect 4460 -2775 4520 -2745
rect 4460 -2815 4470 -2775
rect 4510 -2815 4520 -2775
rect 4460 -2840 4520 -2815
rect 4460 -2880 4470 -2840
rect 4510 -2880 4520 -2840
rect 4460 -2900 4520 -2880
rect 4460 -2940 4470 -2900
rect 4510 -2940 4520 -2900
rect 4460 -2965 4520 -2940
rect 4460 -3005 4470 -2965
rect 4510 -3005 4520 -2965
rect 4460 -3035 4520 -3005
rect 4460 -3075 4470 -3035
rect 4510 -3075 4520 -3035
rect 4460 -3105 4520 -3075
rect 4460 -3145 4470 -3105
rect 4510 -3145 4520 -3105
rect 4460 -3175 4520 -3145
rect 4460 -3215 4470 -3175
rect 4510 -3215 4520 -3175
rect 4460 -3240 4520 -3215
rect 4460 -3280 4470 -3240
rect 4510 -3280 4520 -3240
rect 4460 -3300 4520 -3280
rect 4460 -3340 4470 -3300
rect 4510 -3340 4520 -3300
rect 4460 -3365 4520 -3340
rect 4460 -3405 4470 -3365
rect 4510 -3405 4520 -3365
rect 4460 -3435 4520 -3405
rect 4460 -3475 4470 -3435
rect 4510 -3475 4520 -3435
rect 4460 -3505 4520 -3475
rect 4460 -3545 4470 -3505
rect 4510 -3545 4520 -3505
rect 4460 -3575 4520 -3545
rect 4460 -3615 4470 -3575
rect 4510 -3615 4520 -3575
rect 4460 -3640 4520 -3615
rect 4460 -3680 4470 -3640
rect 4510 -3680 4520 -3640
rect 4460 -3700 4520 -3680
rect 4460 -3740 4470 -3700
rect 4510 -3740 4520 -3700
rect 4460 -3765 4520 -3740
rect 4460 -3805 4470 -3765
rect 4510 -3805 4520 -3765
rect 4460 -3835 4520 -3805
rect 4460 -3875 4470 -3835
rect 4510 -3875 4520 -3835
rect 4460 -3905 4520 -3875
rect 4460 -3945 4470 -3905
rect 4510 -3945 4520 -3905
rect 4460 -3975 4520 -3945
rect 4460 -4015 4470 -3975
rect 4510 -4015 4520 -3975
rect 4460 -4040 4520 -4015
rect 4460 -4080 4470 -4040
rect 4510 -4080 4520 -4040
rect 4460 -4100 4520 -4080
rect 4460 -4140 4470 -4100
rect 4510 -4140 4520 -4100
rect 4460 -4165 4520 -4140
rect 4460 -4205 4470 -4165
rect 4510 -4205 4520 -4165
rect 4460 -4235 4520 -4205
rect 4460 -4275 4470 -4235
rect 4510 -4275 4520 -4235
rect 4460 -4305 4520 -4275
rect 4460 -4345 4470 -4305
rect 4510 -4345 4520 -4305
rect 4460 -4375 4520 -4345
rect 4460 -4415 4470 -4375
rect 4510 -4415 4520 -4375
rect 4460 -4440 4520 -4415
rect 4460 -4480 4470 -4440
rect 4510 -4480 4520 -4440
rect 4460 -4490 4520 -4480
rect 4810 -1300 4870 -1290
rect 4810 -1340 4820 -1300
rect 4860 -1340 4870 -1300
rect 4810 -1365 4870 -1340
rect 4810 -1405 4820 -1365
rect 4860 -1405 4870 -1365
rect 4810 -1435 4870 -1405
rect 4810 -1475 4820 -1435
rect 4860 -1475 4870 -1435
rect 4810 -1505 4870 -1475
rect 4810 -1545 4820 -1505
rect 4860 -1545 4870 -1505
rect 4810 -1575 4870 -1545
rect 4810 -1615 4820 -1575
rect 4860 -1615 4870 -1575
rect 4810 -1640 4870 -1615
rect 4810 -1680 4820 -1640
rect 4860 -1680 4870 -1640
rect 4810 -1700 4870 -1680
rect 4810 -1740 4820 -1700
rect 4860 -1740 4870 -1700
rect 4810 -1765 4870 -1740
rect 4810 -1805 4820 -1765
rect 4860 -1805 4870 -1765
rect 4810 -1835 4870 -1805
rect 4810 -1875 4820 -1835
rect 4860 -1875 4870 -1835
rect 4810 -1905 4870 -1875
rect 4810 -1945 4820 -1905
rect 4860 -1945 4870 -1905
rect 4810 -1975 4870 -1945
rect 4810 -2015 4820 -1975
rect 4860 -2015 4870 -1975
rect 4810 -2040 4870 -2015
rect 4810 -2080 4820 -2040
rect 4860 -2080 4870 -2040
rect 4810 -2100 4870 -2080
rect 4810 -2140 4820 -2100
rect 4860 -2140 4870 -2100
rect 4810 -2165 4870 -2140
rect 4810 -2205 4820 -2165
rect 4860 -2205 4870 -2165
rect 4810 -2235 4870 -2205
rect 4810 -2275 4820 -2235
rect 4860 -2275 4870 -2235
rect 4810 -2305 4870 -2275
rect 4810 -2345 4820 -2305
rect 4860 -2345 4870 -2305
rect 4810 -2375 4870 -2345
rect 4810 -2415 4820 -2375
rect 4860 -2415 4870 -2375
rect 4810 -2440 4870 -2415
rect 4810 -2480 4820 -2440
rect 4860 -2480 4870 -2440
rect 4810 -2500 4870 -2480
rect 4810 -2540 4820 -2500
rect 4860 -2540 4870 -2500
rect 4810 -2565 4870 -2540
rect 4810 -2605 4820 -2565
rect 4860 -2605 4870 -2565
rect 4810 -2635 4870 -2605
rect 4810 -2675 4820 -2635
rect 4860 -2675 4870 -2635
rect 4810 -2705 4870 -2675
rect 4810 -2745 4820 -2705
rect 4860 -2745 4870 -2705
rect 4810 -2775 4870 -2745
rect 4810 -2815 4820 -2775
rect 4860 -2815 4870 -2775
rect 4810 -2840 4870 -2815
rect 4810 -2880 4820 -2840
rect 4860 -2880 4870 -2840
rect 4810 -2900 4870 -2880
rect 4810 -2940 4820 -2900
rect 4860 -2940 4870 -2900
rect 4810 -2965 4870 -2940
rect 4810 -3005 4820 -2965
rect 4860 -3005 4870 -2965
rect 4810 -3035 4870 -3005
rect 4810 -3075 4820 -3035
rect 4860 -3075 4870 -3035
rect 4810 -3105 4870 -3075
rect 4810 -3145 4820 -3105
rect 4860 -3145 4870 -3105
rect 4810 -3175 4870 -3145
rect 4810 -3215 4820 -3175
rect 4860 -3215 4870 -3175
rect 4810 -3240 4870 -3215
rect 4810 -3280 4820 -3240
rect 4860 -3280 4870 -3240
rect 4810 -3300 4870 -3280
rect 4810 -3340 4820 -3300
rect 4860 -3340 4870 -3300
rect 4810 -3365 4870 -3340
rect 4810 -3405 4820 -3365
rect 4860 -3405 4870 -3365
rect 4810 -3435 4870 -3405
rect 4810 -3475 4820 -3435
rect 4860 -3475 4870 -3435
rect 4810 -3505 4870 -3475
rect 4810 -3545 4820 -3505
rect 4860 -3545 4870 -3505
rect 4810 -3575 4870 -3545
rect 4810 -3615 4820 -3575
rect 4860 -3615 4870 -3575
rect 4810 -3640 4870 -3615
rect 4810 -3680 4820 -3640
rect 4860 -3680 4870 -3640
rect 4810 -3700 4870 -3680
rect 4810 -3740 4820 -3700
rect 4860 -3740 4870 -3700
rect 4810 -3765 4870 -3740
rect 4810 -3805 4820 -3765
rect 4860 -3805 4870 -3765
rect 4810 -3835 4870 -3805
rect 4810 -3875 4820 -3835
rect 4860 -3875 4870 -3835
rect 4810 -3905 4870 -3875
rect 4810 -3945 4820 -3905
rect 4860 -3945 4870 -3905
rect 4810 -3975 4870 -3945
rect 4810 -4015 4820 -3975
rect 4860 -4015 4870 -3975
rect 4810 -4040 4870 -4015
rect 4810 -4080 4820 -4040
rect 4860 -4080 4870 -4040
rect 4810 -4100 4870 -4080
rect 4810 -4140 4820 -4100
rect 4860 -4140 4870 -4100
rect 4810 -4165 4870 -4140
rect 4810 -4205 4820 -4165
rect 4860 -4205 4870 -4165
rect 4810 -4235 4870 -4205
rect 4810 -4275 4820 -4235
rect 4860 -4275 4870 -4235
rect 4810 -4305 4870 -4275
rect 4810 -4345 4820 -4305
rect 4860 -4345 4870 -4305
rect 4810 -4375 4870 -4345
rect 4810 -4415 4820 -4375
rect 4860 -4415 4870 -4375
rect 4810 -4440 4870 -4415
rect 4810 -4480 4820 -4440
rect 4860 -4480 4870 -4440
rect 4810 -4490 4870 -4480
rect 5160 -1300 5220 -1290
rect 5160 -1340 5170 -1300
rect 5210 -1340 5220 -1300
rect 5160 -1365 5220 -1340
rect 5160 -1405 5170 -1365
rect 5210 -1405 5220 -1365
rect 5160 -1435 5220 -1405
rect 5160 -1475 5170 -1435
rect 5210 -1475 5220 -1435
rect 5160 -1505 5220 -1475
rect 5160 -1545 5170 -1505
rect 5210 -1545 5220 -1505
rect 5160 -1575 5220 -1545
rect 5160 -1615 5170 -1575
rect 5210 -1615 5220 -1575
rect 5160 -1640 5220 -1615
rect 5160 -1680 5170 -1640
rect 5210 -1680 5220 -1640
rect 5160 -1700 5220 -1680
rect 5160 -1740 5170 -1700
rect 5210 -1740 5220 -1700
rect 5160 -1765 5220 -1740
rect 5160 -1805 5170 -1765
rect 5210 -1805 5220 -1765
rect 5160 -1835 5220 -1805
rect 5160 -1875 5170 -1835
rect 5210 -1875 5220 -1835
rect 5160 -1905 5220 -1875
rect 5160 -1945 5170 -1905
rect 5210 -1945 5220 -1905
rect 5160 -1975 5220 -1945
rect 5160 -2015 5170 -1975
rect 5210 -2015 5220 -1975
rect 5160 -2040 5220 -2015
rect 5160 -2080 5170 -2040
rect 5210 -2080 5220 -2040
rect 5160 -2100 5220 -2080
rect 5160 -2140 5170 -2100
rect 5210 -2140 5220 -2100
rect 5160 -2165 5220 -2140
rect 5160 -2205 5170 -2165
rect 5210 -2205 5220 -2165
rect 5160 -2235 5220 -2205
rect 5160 -2275 5170 -2235
rect 5210 -2275 5220 -2235
rect 5160 -2305 5220 -2275
rect 5160 -2345 5170 -2305
rect 5210 -2345 5220 -2305
rect 5160 -2375 5220 -2345
rect 5160 -2415 5170 -2375
rect 5210 -2415 5220 -2375
rect 5160 -2440 5220 -2415
rect 5160 -2480 5170 -2440
rect 5210 -2480 5220 -2440
rect 5160 -2500 5220 -2480
rect 5160 -2540 5170 -2500
rect 5210 -2540 5220 -2500
rect 5160 -2565 5220 -2540
rect 5160 -2605 5170 -2565
rect 5210 -2605 5220 -2565
rect 5160 -2635 5220 -2605
rect 5160 -2675 5170 -2635
rect 5210 -2675 5220 -2635
rect 5160 -2705 5220 -2675
rect 5160 -2745 5170 -2705
rect 5210 -2745 5220 -2705
rect 5160 -2775 5220 -2745
rect 5160 -2815 5170 -2775
rect 5210 -2815 5220 -2775
rect 5160 -2840 5220 -2815
rect 5160 -2880 5170 -2840
rect 5210 -2880 5220 -2840
rect 5160 -2900 5220 -2880
rect 5160 -2940 5170 -2900
rect 5210 -2940 5220 -2900
rect 5160 -2965 5220 -2940
rect 5160 -3005 5170 -2965
rect 5210 -3005 5220 -2965
rect 5160 -3035 5220 -3005
rect 5160 -3075 5170 -3035
rect 5210 -3075 5220 -3035
rect 5160 -3105 5220 -3075
rect 5160 -3145 5170 -3105
rect 5210 -3145 5220 -3105
rect 5160 -3175 5220 -3145
rect 5160 -3215 5170 -3175
rect 5210 -3215 5220 -3175
rect 5160 -3240 5220 -3215
rect 5160 -3280 5170 -3240
rect 5210 -3280 5220 -3240
rect 5160 -3300 5220 -3280
rect 5160 -3340 5170 -3300
rect 5210 -3340 5220 -3300
rect 5160 -3365 5220 -3340
rect 5160 -3405 5170 -3365
rect 5210 -3405 5220 -3365
rect 5160 -3435 5220 -3405
rect 5160 -3475 5170 -3435
rect 5210 -3475 5220 -3435
rect 5160 -3505 5220 -3475
rect 5160 -3545 5170 -3505
rect 5210 -3545 5220 -3505
rect 5160 -3575 5220 -3545
rect 5160 -3615 5170 -3575
rect 5210 -3615 5220 -3575
rect 5160 -3640 5220 -3615
rect 5160 -3680 5170 -3640
rect 5210 -3680 5220 -3640
rect 5160 -3700 5220 -3680
rect 5160 -3740 5170 -3700
rect 5210 -3740 5220 -3700
rect 5160 -3765 5220 -3740
rect 5160 -3805 5170 -3765
rect 5210 -3805 5220 -3765
rect 5160 -3835 5220 -3805
rect 5160 -3875 5170 -3835
rect 5210 -3875 5220 -3835
rect 5160 -3905 5220 -3875
rect 5160 -3945 5170 -3905
rect 5210 -3945 5220 -3905
rect 5160 -3975 5220 -3945
rect 5160 -4015 5170 -3975
rect 5210 -4015 5220 -3975
rect 5160 -4040 5220 -4015
rect 5160 -4080 5170 -4040
rect 5210 -4080 5220 -4040
rect 5160 -4100 5220 -4080
rect 5160 -4140 5170 -4100
rect 5210 -4140 5220 -4100
rect 5160 -4165 5220 -4140
rect 5160 -4205 5170 -4165
rect 5210 -4205 5220 -4165
rect 5160 -4235 5220 -4205
rect 5160 -4275 5170 -4235
rect 5210 -4275 5220 -4235
rect 5160 -4305 5220 -4275
rect 5160 -4345 5170 -4305
rect 5210 -4345 5220 -4305
rect 5160 -4375 5220 -4345
rect 5160 -4415 5170 -4375
rect 5210 -4415 5220 -4375
rect 5160 -4440 5220 -4415
rect 5160 -4480 5170 -4440
rect 5210 -4480 5220 -4440
rect 5160 -4490 5220 -4480
rect 5510 -1300 5570 -1290
rect 5510 -1340 5520 -1300
rect 5560 -1340 5570 -1300
rect 5510 -1365 5570 -1340
rect 5510 -1405 5520 -1365
rect 5560 -1405 5570 -1365
rect 5510 -1435 5570 -1405
rect 5510 -1475 5520 -1435
rect 5560 -1475 5570 -1435
rect 5510 -1505 5570 -1475
rect 5510 -1545 5520 -1505
rect 5560 -1545 5570 -1505
rect 5510 -1575 5570 -1545
rect 5510 -1615 5520 -1575
rect 5560 -1615 5570 -1575
rect 5510 -1640 5570 -1615
rect 5510 -1680 5520 -1640
rect 5560 -1680 5570 -1640
rect 5510 -1700 5570 -1680
rect 5510 -1740 5520 -1700
rect 5560 -1740 5570 -1700
rect 5510 -1765 5570 -1740
rect 5510 -1805 5520 -1765
rect 5560 -1805 5570 -1765
rect 5510 -1835 5570 -1805
rect 5510 -1875 5520 -1835
rect 5560 -1875 5570 -1835
rect 5510 -1905 5570 -1875
rect 5510 -1945 5520 -1905
rect 5560 -1945 5570 -1905
rect 5510 -1975 5570 -1945
rect 5510 -2015 5520 -1975
rect 5560 -2015 5570 -1975
rect 5510 -2040 5570 -2015
rect 5510 -2080 5520 -2040
rect 5560 -2080 5570 -2040
rect 5510 -2100 5570 -2080
rect 5510 -2140 5520 -2100
rect 5560 -2140 5570 -2100
rect 5510 -2165 5570 -2140
rect 5510 -2205 5520 -2165
rect 5560 -2205 5570 -2165
rect 5510 -2235 5570 -2205
rect 5510 -2275 5520 -2235
rect 5560 -2275 5570 -2235
rect 5510 -2305 5570 -2275
rect 5510 -2345 5520 -2305
rect 5560 -2345 5570 -2305
rect 5510 -2375 5570 -2345
rect 5510 -2415 5520 -2375
rect 5560 -2415 5570 -2375
rect 5510 -2440 5570 -2415
rect 5510 -2480 5520 -2440
rect 5560 -2480 5570 -2440
rect 5510 -2500 5570 -2480
rect 5510 -2540 5520 -2500
rect 5560 -2540 5570 -2500
rect 5510 -2565 5570 -2540
rect 5510 -2605 5520 -2565
rect 5560 -2605 5570 -2565
rect 5510 -2635 5570 -2605
rect 5510 -2675 5520 -2635
rect 5560 -2675 5570 -2635
rect 5510 -2705 5570 -2675
rect 5510 -2745 5520 -2705
rect 5560 -2745 5570 -2705
rect 5510 -2775 5570 -2745
rect 5510 -2815 5520 -2775
rect 5560 -2815 5570 -2775
rect 5510 -2840 5570 -2815
rect 5510 -2880 5520 -2840
rect 5560 -2880 5570 -2840
rect 5510 -2900 5570 -2880
rect 5510 -2940 5520 -2900
rect 5560 -2940 5570 -2900
rect 5510 -2965 5570 -2940
rect 5510 -3005 5520 -2965
rect 5560 -3005 5570 -2965
rect 5510 -3035 5570 -3005
rect 5510 -3075 5520 -3035
rect 5560 -3075 5570 -3035
rect 5510 -3105 5570 -3075
rect 5510 -3145 5520 -3105
rect 5560 -3145 5570 -3105
rect 5510 -3175 5570 -3145
rect 5510 -3215 5520 -3175
rect 5560 -3215 5570 -3175
rect 5510 -3240 5570 -3215
rect 5510 -3280 5520 -3240
rect 5560 -3280 5570 -3240
rect 5510 -3300 5570 -3280
rect 5510 -3340 5520 -3300
rect 5560 -3340 5570 -3300
rect 5510 -3365 5570 -3340
rect 5510 -3405 5520 -3365
rect 5560 -3405 5570 -3365
rect 5510 -3435 5570 -3405
rect 5510 -3475 5520 -3435
rect 5560 -3475 5570 -3435
rect 5510 -3505 5570 -3475
rect 5510 -3545 5520 -3505
rect 5560 -3545 5570 -3505
rect 5510 -3575 5570 -3545
rect 5510 -3615 5520 -3575
rect 5560 -3615 5570 -3575
rect 5510 -3640 5570 -3615
rect 5510 -3680 5520 -3640
rect 5560 -3680 5570 -3640
rect 5510 -3700 5570 -3680
rect 5510 -3740 5520 -3700
rect 5560 -3740 5570 -3700
rect 5510 -3765 5570 -3740
rect 5510 -3805 5520 -3765
rect 5560 -3805 5570 -3765
rect 5510 -3835 5570 -3805
rect 5510 -3875 5520 -3835
rect 5560 -3875 5570 -3835
rect 5510 -3905 5570 -3875
rect 5510 -3945 5520 -3905
rect 5560 -3945 5570 -3905
rect 5510 -3975 5570 -3945
rect 5510 -4015 5520 -3975
rect 5560 -4015 5570 -3975
rect 5510 -4040 5570 -4015
rect 5510 -4080 5520 -4040
rect 5560 -4080 5570 -4040
rect 5510 -4100 5570 -4080
rect 5510 -4140 5520 -4100
rect 5560 -4140 5570 -4100
rect 5510 -4165 5570 -4140
rect 5510 -4205 5520 -4165
rect 5560 -4205 5570 -4165
rect 5510 -4235 5570 -4205
rect 5510 -4275 5520 -4235
rect 5560 -4275 5570 -4235
rect 5510 -4305 5570 -4275
rect 5510 -4345 5520 -4305
rect 5560 -4345 5570 -4305
rect 5510 -4375 5570 -4345
rect 5510 -4415 5520 -4375
rect 5560 -4415 5570 -4375
rect 5510 -4440 5570 -4415
rect 5510 -4480 5520 -4440
rect 5560 -4480 5570 -4440
rect 5510 -4490 5570 -4480
rect 5860 -1300 5920 -1290
rect 5860 -1340 5870 -1300
rect 5910 -1340 5920 -1300
rect 5860 -1365 5920 -1340
rect 5860 -1405 5870 -1365
rect 5910 -1405 5920 -1365
rect 5860 -1435 5920 -1405
rect 5860 -1475 5870 -1435
rect 5910 -1475 5920 -1435
rect 5860 -1505 5920 -1475
rect 5860 -1545 5870 -1505
rect 5910 -1545 5920 -1505
rect 5860 -1575 5920 -1545
rect 5860 -1615 5870 -1575
rect 5910 -1615 5920 -1575
rect 5860 -1640 5920 -1615
rect 5860 -1680 5870 -1640
rect 5910 -1680 5920 -1640
rect 5860 -1700 5920 -1680
rect 5860 -1740 5870 -1700
rect 5910 -1740 5920 -1700
rect 5860 -1765 5920 -1740
rect 5860 -1805 5870 -1765
rect 5910 -1805 5920 -1765
rect 5860 -1835 5920 -1805
rect 5860 -1875 5870 -1835
rect 5910 -1875 5920 -1835
rect 5860 -1905 5920 -1875
rect 5860 -1945 5870 -1905
rect 5910 -1945 5920 -1905
rect 5860 -1975 5920 -1945
rect 5860 -2015 5870 -1975
rect 5910 -2015 5920 -1975
rect 5860 -2040 5920 -2015
rect 5860 -2080 5870 -2040
rect 5910 -2080 5920 -2040
rect 5860 -2100 5920 -2080
rect 5860 -2140 5870 -2100
rect 5910 -2140 5920 -2100
rect 5860 -2165 5920 -2140
rect 5860 -2205 5870 -2165
rect 5910 -2205 5920 -2165
rect 5860 -2235 5920 -2205
rect 5860 -2275 5870 -2235
rect 5910 -2275 5920 -2235
rect 5860 -2305 5920 -2275
rect 5860 -2345 5870 -2305
rect 5910 -2345 5920 -2305
rect 5860 -2375 5920 -2345
rect 5860 -2415 5870 -2375
rect 5910 -2415 5920 -2375
rect 5860 -2440 5920 -2415
rect 5860 -2480 5870 -2440
rect 5910 -2480 5920 -2440
rect 5860 -2500 5920 -2480
rect 5860 -2540 5870 -2500
rect 5910 -2540 5920 -2500
rect 5860 -2565 5920 -2540
rect 5860 -2605 5870 -2565
rect 5910 -2605 5920 -2565
rect 5860 -2635 5920 -2605
rect 5860 -2675 5870 -2635
rect 5910 -2675 5920 -2635
rect 5860 -2705 5920 -2675
rect 5860 -2745 5870 -2705
rect 5910 -2745 5920 -2705
rect 5860 -2775 5920 -2745
rect 5860 -2815 5870 -2775
rect 5910 -2815 5920 -2775
rect 5860 -2840 5920 -2815
rect 5860 -2880 5870 -2840
rect 5910 -2880 5920 -2840
rect 5860 -2900 5920 -2880
rect 5860 -2940 5870 -2900
rect 5910 -2940 5920 -2900
rect 5860 -2965 5920 -2940
rect 5860 -3005 5870 -2965
rect 5910 -3005 5920 -2965
rect 5860 -3035 5920 -3005
rect 5860 -3075 5870 -3035
rect 5910 -3075 5920 -3035
rect 5860 -3105 5920 -3075
rect 5860 -3145 5870 -3105
rect 5910 -3145 5920 -3105
rect 5860 -3175 5920 -3145
rect 5860 -3215 5870 -3175
rect 5910 -3215 5920 -3175
rect 5860 -3240 5920 -3215
rect 5860 -3280 5870 -3240
rect 5910 -3280 5920 -3240
rect 5860 -3300 5920 -3280
rect 5860 -3340 5870 -3300
rect 5910 -3340 5920 -3300
rect 5860 -3365 5920 -3340
rect 5860 -3405 5870 -3365
rect 5910 -3405 5920 -3365
rect 5860 -3435 5920 -3405
rect 5860 -3475 5870 -3435
rect 5910 -3475 5920 -3435
rect 5860 -3505 5920 -3475
rect 5860 -3545 5870 -3505
rect 5910 -3545 5920 -3505
rect 5860 -3575 5920 -3545
rect 5860 -3615 5870 -3575
rect 5910 -3615 5920 -3575
rect 5860 -3640 5920 -3615
rect 5860 -3680 5870 -3640
rect 5910 -3680 5920 -3640
rect 5860 -3700 5920 -3680
rect 5860 -3740 5870 -3700
rect 5910 -3740 5920 -3700
rect 5860 -3765 5920 -3740
rect 5860 -3805 5870 -3765
rect 5910 -3805 5920 -3765
rect 5860 -3835 5920 -3805
rect 5860 -3875 5870 -3835
rect 5910 -3875 5920 -3835
rect 5860 -3905 5920 -3875
rect 5860 -3945 5870 -3905
rect 5910 -3945 5920 -3905
rect 5860 -3975 5920 -3945
rect 5860 -4015 5870 -3975
rect 5910 -4015 5920 -3975
rect 5860 -4040 5920 -4015
rect 5860 -4080 5870 -4040
rect 5910 -4080 5920 -4040
rect 5860 -4100 5920 -4080
rect 5860 -4140 5870 -4100
rect 5910 -4140 5920 -4100
rect 5860 -4165 5920 -4140
rect 5860 -4205 5870 -4165
rect 5910 -4205 5920 -4165
rect 5860 -4235 5920 -4205
rect 5860 -4275 5870 -4235
rect 5910 -4275 5920 -4235
rect 5860 -4305 5920 -4275
rect 5860 -4345 5870 -4305
rect 5910 -4345 5920 -4305
rect 5860 -4375 5920 -4345
rect 5860 -4415 5870 -4375
rect 5910 -4415 5920 -4375
rect 5860 -4440 5920 -4415
rect 5860 -4480 5870 -4440
rect 5910 -4480 5920 -4440
rect 5860 -4490 5920 -4480
rect 6210 -1300 6270 -1290
rect 6210 -1340 6220 -1300
rect 6260 -1340 6270 -1300
rect 6210 -1365 6270 -1340
rect 6210 -1405 6220 -1365
rect 6260 -1405 6270 -1365
rect 6210 -1435 6270 -1405
rect 6210 -1475 6220 -1435
rect 6260 -1475 6270 -1435
rect 6210 -1505 6270 -1475
rect 6210 -1545 6220 -1505
rect 6260 -1545 6270 -1505
rect 6210 -1575 6270 -1545
rect 6210 -1615 6220 -1575
rect 6260 -1615 6270 -1575
rect 6210 -1640 6270 -1615
rect 6210 -1680 6220 -1640
rect 6260 -1680 6270 -1640
rect 6210 -1700 6270 -1680
rect 6210 -1740 6220 -1700
rect 6260 -1740 6270 -1700
rect 6210 -1765 6270 -1740
rect 6210 -1805 6220 -1765
rect 6260 -1805 6270 -1765
rect 6210 -1835 6270 -1805
rect 6210 -1875 6220 -1835
rect 6260 -1875 6270 -1835
rect 6210 -1905 6270 -1875
rect 6210 -1945 6220 -1905
rect 6260 -1945 6270 -1905
rect 6210 -1975 6270 -1945
rect 6210 -2015 6220 -1975
rect 6260 -2015 6270 -1975
rect 6210 -2040 6270 -2015
rect 6210 -2080 6220 -2040
rect 6260 -2080 6270 -2040
rect 6210 -2100 6270 -2080
rect 6210 -2140 6220 -2100
rect 6260 -2140 6270 -2100
rect 6210 -2165 6270 -2140
rect 6210 -2205 6220 -2165
rect 6260 -2205 6270 -2165
rect 6210 -2235 6270 -2205
rect 6210 -2275 6220 -2235
rect 6260 -2275 6270 -2235
rect 6210 -2305 6270 -2275
rect 6210 -2345 6220 -2305
rect 6260 -2345 6270 -2305
rect 6210 -2375 6270 -2345
rect 6210 -2415 6220 -2375
rect 6260 -2415 6270 -2375
rect 6210 -2440 6270 -2415
rect 6210 -2480 6220 -2440
rect 6260 -2480 6270 -2440
rect 6210 -2500 6270 -2480
rect 6210 -2540 6220 -2500
rect 6260 -2540 6270 -2500
rect 6210 -2565 6270 -2540
rect 6210 -2605 6220 -2565
rect 6260 -2605 6270 -2565
rect 6210 -2635 6270 -2605
rect 6210 -2675 6220 -2635
rect 6260 -2675 6270 -2635
rect 6210 -2705 6270 -2675
rect 6210 -2745 6220 -2705
rect 6260 -2745 6270 -2705
rect 6210 -2775 6270 -2745
rect 6210 -2815 6220 -2775
rect 6260 -2815 6270 -2775
rect 6210 -2840 6270 -2815
rect 6210 -2880 6220 -2840
rect 6260 -2880 6270 -2840
rect 6210 -2900 6270 -2880
rect 6210 -2940 6220 -2900
rect 6260 -2940 6270 -2900
rect 6210 -2965 6270 -2940
rect 6210 -3005 6220 -2965
rect 6260 -3005 6270 -2965
rect 6210 -3035 6270 -3005
rect 6210 -3075 6220 -3035
rect 6260 -3075 6270 -3035
rect 6210 -3105 6270 -3075
rect 6210 -3145 6220 -3105
rect 6260 -3145 6270 -3105
rect 6210 -3175 6270 -3145
rect 6210 -3215 6220 -3175
rect 6260 -3215 6270 -3175
rect 6210 -3240 6270 -3215
rect 6210 -3280 6220 -3240
rect 6260 -3280 6270 -3240
rect 6210 -3300 6270 -3280
rect 6210 -3340 6220 -3300
rect 6260 -3340 6270 -3300
rect 6210 -3365 6270 -3340
rect 6210 -3405 6220 -3365
rect 6260 -3405 6270 -3365
rect 6210 -3435 6270 -3405
rect 6210 -3475 6220 -3435
rect 6260 -3475 6270 -3435
rect 6210 -3505 6270 -3475
rect 6210 -3545 6220 -3505
rect 6260 -3545 6270 -3505
rect 6210 -3575 6270 -3545
rect 6210 -3615 6220 -3575
rect 6260 -3615 6270 -3575
rect 6210 -3640 6270 -3615
rect 6210 -3680 6220 -3640
rect 6260 -3680 6270 -3640
rect 6210 -3700 6270 -3680
rect 6210 -3740 6220 -3700
rect 6260 -3740 6270 -3700
rect 6210 -3765 6270 -3740
rect 6210 -3805 6220 -3765
rect 6260 -3805 6270 -3765
rect 6210 -3835 6270 -3805
rect 6210 -3875 6220 -3835
rect 6260 -3875 6270 -3835
rect 6210 -3905 6270 -3875
rect 6210 -3945 6220 -3905
rect 6260 -3945 6270 -3905
rect 6210 -3975 6270 -3945
rect 6210 -4015 6220 -3975
rect 6260 -4015 6270 -3975
rect 6210 -4040 6270 -4015
rect 6210 -4080 6220 -4040
rect 6260 -4080 6270 -4040
rect 6210 -4100 6270 -4080
rect 6210 -4140 6220 -4100
rect 6260 -4140 6270 -4100
rect 6210 -4165 6270 -4140
rect 6210 -4205 6220 -4165
rect 6260 -4205 6270 -4165
rect 6210 -4235 6270 -4205
rect 6210 -4275 6220 -4235
rect 6260 -4275 6270 -4235
rect 6210 -4305 6270 -4275
rect 6210 -4345 6220 -4305
rect 6260 -4345 6270 -4305
rect 6210 -4375 6270 -4345
rect 6210 -4415 6220 -4375
rect 6260 -4415 6270 -4375
rect 6210 -4440 6270 -4415
rect 6210 -4480 6220 -4440
rect 6260 -4480 6270 -4440
rect 6210 -4490 6270 -4480
rect 6560 -1300 6620 -1290
rect 6560 -1340 6570 -1300
rect 6610 -1340 6620 -1300
rect 6560 -1365 6620 -1340
rect 6560 -1405 6570 -1365
rect 6610 -1405 6620 -1365
rect 6560 -1435 6620 -1405
rect 6560 -1475 6570 -1435
rect 6610 -1475 6620 -1435
rect 6560 -1505 6620 -1475
rect 6560 -1545 6570 -1505
rect 6610 -1545 6620 -1505
rect 6560 -1575 6620 -1545
rect 6560 -1615 6570 -1575
rect 6610 -1615 6620 -1575
rect 6560 -1640 6620 -1615
rect 6560 -1680 6570 -1640
rect 6610 -1680 6620 -1640
rect 6560 -1700 6620 -1680
rect 6560 -1740 6570 -1700
rect 6610 -1740 6620 -1700
rect 6560 -1765 6620 -1740
rect 6560 -1805 6570 -1765
rect 6610 -1805 6620 -1765
rect 6560 -1835 6620 -1805
rect 6560 -1875 6570 -1835
rect 6610 -1875 6620 -1835
rect 6560 -1905 6620 -1875
rect 6560 -1945 6570 -1905
rect 6610 -1945 6620 -1905
rect 6560 -1975 6620 -1945
rect 6560 -2015 6570 -1975
rect 6610 -2015 6620 -1975
rect 6560 -2040 6620 -2015
rect 6560 -2080 6570 -2040
rect 6610 -2080 6620 -2040
rect 6560 -2100 6620 -2080
rect 6560 -2140 6570 -2100
rect 6610 -2140 6620 -2100
rect 6560 -2165 6620 -2140
rect 6560 -2205 6570 -2165
rect 6610 -2205 6620 -2165
rect 6560 -2235 6620 -2205
rect 6560 -2275 6570 -2235
rect 6610 -2275 6620 -2235
rect 6560 -2305 6620 -2275
rect 6560 -2345 6570 -2305
rect 6610 -2345 6620 -2305
rect 6560 -2375 6620 -2345
rect 6560 -2415 6570 -2375
rect 6610 -2415 6620 -2375
rect 6560 -2440 6620 -2415
rect 6560 -2480 6570 -2440
rect 6610 -2480 6620 -2440
rect 6560 -2500 6620 -2480
rect 6560 -2540 6570 -2500
rect 6610 -2540 6620 -2500
rect 6560 -2565 6620 -2540
rect 6560 -2605 6570 -2565
rect 6610 -2605 6620 -2565
rect 6560 -2635 6620 -2605
rect 6560 -2675 6570 -2635
rect 6610 -2675 6620 -2635
rect 6560 -2705 6620 -2675
rect 6560 -2745 6570 -2705
rect 6610 -2745 6620 -2705
rect 6560 -2775 6620 -2745
rect 6560 -2815 6570 -2775
rect 6610 -2815 6620 -2775
rect 6560 -2840 6620 -2815
rect 6560 -2880 6570 -2840
rect 6610 -2880 6620 -2840
rect 6560 -2900 6620 -2880
rect 6560 -2940 6570 -2900
rect 6610 -2940 6620 -2900
rect 6560 -2965 6620 -2940
rect 6560 -3005 6570 -2965
rect 6610 -3005 6620 -2965
rect 6560 -3035 6620 -3005
rect 6560 -3075 6570 -3035
rect 6610 -3075 6620 -3035
rect 6560 -3105 6620 -3075
rect 6560 -3145 6570 -3105
rect 6610 -3145 6620 -3105
rect 6560 -3175 6620 -3145
rect 6560 -3215 6570 -3175
rect 6610 -3215 6620 -3175
rect 6560 -3240 6620 -3215
rect 6560 -3280 6570 -3240
rect 6610 -3280 6620 -3240
rect 6560 -3300 6620 -3280
rect 6560 -3340 6570 -3300
rect 6610 -3340 6620 -3300
rect 6560 -3365 6620 -3340
rect 6560 -3405 6570 -3365
rect 6610 -3405 6620 -3365
rect 6560 -3435 6620 -3405
rect 6560 -3475 6570 -3435
rect 6610 -3475 6620 -3435
rect 6560 -3505 6620 -3475
rect 6560 -3545 6570 -3505
rect 6610 -3545 6620 -3505
rect 6560 -3575 6620 -3545
rect 6560 -3615 6570 -3575
rect 6610 -3615 6620 -3575
rect 6560 -3640 6620 -3615
rect 6560 -3680 6570 -3640
rect 6610 -3680 6620 -3640
rect 6560 -3700 6620 -3680
rect 6560 -3740 6570 -3700
rect 6610 -3740 6620 -3700
rect 6560 -3765 6620 -3740
rect 6560 -3805 6570 -3765
rect 6610 -3805 6620 -3765
rect 6560 -3835 6620 -3805
rect 6560 -3875 6570 -3835
rect 6610 -3875 6620 -3835
rect 6560 -3905 6620 -3875
rect 6560 -3945 6570 -3905
rect 6610 -3945 6620 -3905
rect 6560 -3975 6620 -3945
rect 6560 -4015 6570 -3975
rect 6610 -4015 6620 -3975
rect 6560 -4040 6620 -4015
rect 6560 -4080 6570 -4040
rect 6610 -4080 6620 -4040
rect 6560 -4100 6620 -4080
rect 6560 -4140 6570 -4100
rect 6610 -4140 6620 -4100
rect 6560 -4165 6620 -4140
rect 6560 -4205 6570 -4165
rect 6610 -4205 6620 -4165
rect 6560 -4235 6620 -4205
rect 6560 -4275 6570 -4235
rect 6610 -4275 6620 -4235
rect 6560 -4305 6620 -4275
rect 6560 -4345 6570 -4305
rect 6610 -4345 6620 -4305
rect 6560 -4375 6620 -4345
rect 6560 -4415 6570 -4375
rect 6610 -4415 6620 -4375
rect 6560 -4440 6620 -4415
rect 6560 -4480 6570 -4440
rect 6610 -4480 6620 -4440
rect 6560 -4490 6620 -4480
rect 6910 -1300 6970 -1290
rect 6910 -1340 6920 -1300
rect 6960 -1340 6970 -1300
rect 6910 -1365 6970 -1340
rect 6910 -1405 6920 -1365
rect 6960 -1405 6970 -1365
rect 6910 -1435 6970 -1405
rect 6910 -1475 6920 -1435
rect 6960 -1475 6970 -1435
rect 6910 -1505 6970 -1475
rect 6910 -1545 6920 -1505
rect 6960 -1545 6970 -1505
rect 6910 -1575 6970 -1545
rect 6910 -1615 6920 -1575
rect 6960 -1615 6970 -1575
rect 6910 -1640 6970 -1615
rect 6910 -1680 6920 -1640
rect 6960 -1680 6970 -1640
rect 6910 -1700 6970 -1680
rect 6910 -1740 6920 -1700
rect 6960 -1740 6970 -1700
rect 6910 -1765 6970 -1740
rect 6910 -1805 6920 -1765
rect 6960 -1805 6970 -1765
rect 6910 -1835 6970 -1805
rect 6910 -1875 6920 -1835
rect 6960 -1875 6970 -1835
rect 6910 -1905 6970 -1875
rect 6910 -1945 6920 -1905
rect 6960 -1945 6970 -1905
rect 6910 -1975 6970 -1945
rect 6910 -2015 6920 -1975
rect 6960 -2015 6970 -1975
rect 6910 -2040 6970 -2015
rect 6910 -2080 6920 -2040
rect 6960 -2080 6970 -2040
rect 6910 -2100 6970 -2080
rect 6910 -2140 6920 -2100
rect 6960 -2140 6970 -2100
rect 6910 -2165 6970 -2140
rect 6910 -2205 6920 -2165
rect 6960 -2205 6970 -2165
rect 6910 -2235 6970 -2205
rect 6910 -2275 6920 -2235
rect 6960 -2275 6970 -2235
rect 6910 -2305 6970 -2275
rect 6910 -2345 6920 -2305
rect 6960 -2345 6970 -2305
rect 6910 -2375 6970 -2345
rect 6910 -2415 6920 -2375
rect 6960 -2415 6970 -2375
rect 6910 -2440 6970 -2415
rect 6910 -2480 6920 -2440
rect 6960 -2480 6970 -2440
rect 6910 -2500 6970 -2480
rect 6910 -2540 6920 -2500
rect 6960 -2540 6970 -2500
rect 6910 -2565 6970 -2540
rect 6910 -2605 6920 -2565
rect 6960 -2605 6970 -2565
rect 6910 -2635 6970 -2605
rect 6910 -2675 6920 -2635
rect 6960 -2675 6970 -2635
rect 6910 -2705 6970 -2675
rect 6910 -2745 6920 -2705
rect 6960 -2745 6970 -2705
rect 6910 -2775 6970 -2745
rect 6910 -2815 6920 -2775
rect 6960 -2815 6970 -2775
rect 6910 -2840 6970 -2815
rect 6910 -2880 6920 -2840
rect 6960 -2880 6970 -2840
rect 6910 -2900 6970 -2880
rect 6910 -2940 6920 -2900
rect 6960 -2940 6970 -2900
rect 6910 -2965 6970 -2940
rect 6910 -3005 6920 -2965
rect 6960 -3005 6970 -2965
rect 6910 -3035 6970 -3005
rect 6910 -3075 6920 -3035
rect 6960 -3075 6970 -3035
rect 6910 -3105 6970 -3075
rect 6910 -3145 6920 -3105
rect 6960 -3145 6970 -3105
rect 6910 -3175 6970 -3145
rect 6910 -3215 6920 -3175
rect 6960 -3215 6970 -3175
rect 6910 -3240 6970 -3215
rect 6910 -3280 6920 -3240
rect 6960 -3280 6970 -3240
rect 6910 -3300 6970 -3280
rect 6910 -3340 6920 -3300
rect 6960 -3340 6970 -3300
rect 6910 -3365 6970 -3340
rect 6910 -3405 6920 -3365
rect 6960 -3405 6970 -3365
rect 6910 -3435 6970 -3405
rect 6910 -3475 6920 -3435
rect 6960 -3475 6970 -3435
rect 6910 -3505 6970 -3475
rect 6910 -3545 6920 -3505
rect 6960 -3545 6970 -3505
rect 6910 -3575 6970 -3545
rect 6910 -3615 6920 -3575
rect 6960 -3615 6970 -3575
rect 6910 -3640 6970 -3615
rect 6910 -3680 6920 -3640
rect 6960 -3680 6970 -3640
rect 6910 -3700 6970 -3680
rect 6910 -3740 6920 -3700
rect 6960 -3740 6970 -3700
rect 6910 -3765 6970 -3740
rect 6910 -3805 6920 -3765
rect 6960 -3805 6970 -3765
rect 6910 -3835 6970 -3805
rect 6910 -3875 6920 -3835
rect 6960 -3875 6970 -3835
rect 6910 -3905 6970 -3875
rect 6910 -3945 6920 -3905
rect 6960 -3945 6970 -3905
rect 6910 -3975 6970 -3945
rect 6910 -4015 6920 -3975
rect 6960 -4015 6970 -3975
rect 6910 -4040 6970 -4015
rect 6910 -4080 6920 -4040
rect 6960 -4080 6970 -4040
rect 6910 -4100 6970 -4080
rect 6910 -4140 6920 -4100
rect 6960 -4140 6970 -4100
rect 6910 -4165 6970 -4140
rect 6910 -4205 6920 -4165
rect 6960 -4205 6970 -4165
rect 6910 -4235 6970 -4205
rect 6910 -4275 6920 -4235
rect 6960 -4275 6970 -4235
rect 6910 -4305 6970 -4275
rect 6910 -4345 6920 -4305
rect 6960 -4345 6970 -4305
rect 6910 -4375 6970 -4345
rect 6910 -4415 6920 -4375
rect 6960 -4415 6970 -4375
rect 6910 -4440 6970 -4415
rect 6910 -4480 6920 -4440
rect 6960 -4480 6970 -4440
rect 6910 -4490 6970 -4480
rect 7260 -1300 7320 -1290
rect 7260 -1340 7270 -1300
rect 7310 -1340 7320 -1300
rect 7260 -1365 7320 -1340
rect 7260 -1405 7270 -1365
rect 7310 -1405 7320 -1365
rect 7260 -1435 7320 -1405
rect 7260 -1475 7270 -1435
rect 7310 -1475 7320 -1435
rect 7260 -1505 7320 -1475
rect 7260 -1545 7270 -1505
rect 7310 -1545 7320 -1505
rect 7260 -1575 7320 -1545
rect 7260 -1615 7270 -1575
rect 7310 -1615 7320 -1575
rect 7260 -1640 7320 -1615
rect 7260 -1680 7270 -1640
rect 7310 -1680 7320 -1640
rect 7260 -1700 7320 -1680
rect 7260 -1740 7270 -1700
rect 7310 -1740 7320 -1700
rect 7260 -1765 7320 -1740
rect 7260 -1805 7270 -1765
rect 7310 -1805 7320 -1765
rect 7260 -1835 7320 -1805
rect 7260 -1875 7270 -1835
rect 7310 -1875 7320 -1835
rect 7260 -1905 7320 -1875
rect 7260 -1945 7270 -1905
rect 7310 -1945 7320 -1905
rect 7260 -1975 7320 -1945
rect 7260 -2015 7270 -1975
rect 7310 -2015 7320 -1975
rect 7260 -2040 7320 -2015
rect 7260 -2080 7270 -2040
rect 7310 -2080 7320 -2040
rect 7260 -2100 7320 -2080
rect 7260 -2140 7270 -2100
rect 7310 -2140 7320 -2100
rect 7260 -2165 7320 -2140
rect 7260 -2205 7270 -2165
rect 7310 -2205 7320 -2165
rect 7260 -2235 7320 -2205
rect 7260 -2275 7270 -2235
rect 7310 -2275 7320 -2235
rect 7260 -2305 7320 -2275
rect 7260 -2345 7270 -2305
rect 7310 -2345 7320 -2305
rect 7260 -2375 7320 -2345
rect 7260 -2415 7270 -2375
rect 7310 -2415 7320 -2375
rect 7260 -2440 7320 -2415
rect 7260 -2480 7270 -2440
rect 7310 -2480 7320 -2440
rect 7260 -2500 7320 -2480
rect 7260 -2540 7270 -2500
rect 7310 -2540 7320 -2500
rect 7260 -2565 7320 -2540
rect 7260 -2605 7270 -2565
rect 7310 -2605 7320 -2565
rect 7260 -2635 7320 -2605
rect 7260 -2675 7270 -2635
rect 7310 -2675 7320 -2635
rect 7260 -2705 7320 -2675
rect 7260 -2745 7270 -2705
rect 7310 -2745 7320 -2705
rect 7260 -2775 7320 -2745
rect 7260 -2815 7270 -2775
rect 7310 -2815 7320 -2775
rect 7260 -2840 7320 -2815
rect 7260 -2880 7270 -2840
rect 7310 -2880 7320 -2840
rect 7260 -2900 7320 -2880
rect 7260 -2940 7270 -2900
rect 7310 -2940 7320 -2900
rect 7260 -2965 7320 -2940
rect 7260 -3005 7270 -2965
rect 7310 -3005 7320 -2965
rect 7260 -3035 7320 -3005
rect 7260 -3075 7270 -3035
rect 7310 -3075 7320 -3035
rect 7260 -3105 7320 -3075
rect 7260 -3145 7270 -3105
rect 7310 -3145 7320 -3105
rect 7260 -3175 7320 -3145
rect 7260 -3215 7270 -3175
rect 7310 -3215 7320 -3175
rect 7260 -3240 7320 -3215
rect 7260 -3280 7270 -3240
rect 7310 -3280 7320 -3240
rect 7260 -3300 7320 -3280
rect 7260 -3340 7270 -3300
rect 7310 -3340 7320 -3300
rect 7260 -3365 7320 -3340
rect 7260 -3405 7270 -3365
rect 7310 -3405 7320 -3365
rect 7260 -3435 7320 -3405
rect 7260 -3475 7270 -3435
rect 7310 -3475 7320 -3435
rect 7260 -3505 7320 -3475
rect 7260 -3545 7270 -3505
rect 7310 -3545 7320 -3505
rect 7260 -3575 7320 -3545
rect 7260 -3615 7270 -3575
rect 7310 -3615 7320 -3575
rect 7260 -3640 7320 -3615
rect 7260 -3680 7270 -3640
rect 7310 -3680 7320 -3640
rect 7260 -3700 7320 -3680
rect 7260 -3740 7270 -3700
rect 7310 -3740 7320 -3700
rect 7260 -3765 7320 -3740
rect 7260 -3805 7270 -3765
rect 7310 -3805 7320 -3765
rect 7260 -3835 7320 -3805
rect 7260 -3875 7270 -3835
rect 7310 -3875 7320 -3835
rect 7260 -3905 7320 -3875
rect 7260 -3945 7270 -3905
rect 7310 -3945 7320 -3905
rect 7260 -3975 7320 -3945
rect 7260 -4015 7270 -3975
rect 7310 -4015 7320 -3975
rect 7260 -4040 7320 -4015
rect 7260 -4080 7270 -4040
rect 7310 -4080 7320 -4040
rect 7260 -4100 7320 -4080
rect 7260 -4140 7270 -4100
rect 7310 -4140 7320 -4100
rect 7260 -4165 7320 -4140
rect 7260 -4205 7270 -4165
rect 7310 -4205 7320 -4165
rect 7260 -4235 7320 -4205
rect 7260 -4275 7270 -4235
rect 7310 -4275 7320 -4235
rect 7260 -4305 7320 -4275
rect 7260 -4345 7270 -4305
rect 7310 -4345 7320 -4305
rect 7260 -4375 7320 -4345
rect 7260 -4415 7270 -4375
rect 7310 -4415 7320 -4375
rect 7260 -4440 7320 -4415
rect 7260 -4480 7270 -4440
rect 7310 -4480 7320 -4440
rect 7260 -4490 7320 -4480
rect 7610 -1300 7670 -1290
rect 7610 -1340 7620 -1300
rect 7660 -1340 7670 -1300
rect 7610 -1365 7670 -1340
rect 7610 -1405 7620 -1365
rect 7660 -1405 7670 -1365
rect 7610 -1435 7670 -1405
rect 7610 -1475 7620 -1435
rect 7660 -1475 7670 -1435
rect 7610 -1505 7670 -1475
rect 7610 -1545 7620 -1505
rect 7660 -1545 7670 -1505
rect 7610 -1575 7670 -1545
rect 7610 -1615 7620 -1575
rect 7660 -1615 7670 -1575
rect 7610 -1640 7670 -1615
rect 7610 -1680 7620 -1640
rect 7660 -1680 7670 -1640
rect 7610 -1700 7670 -1680
rect 7610 -1740 7620 -1700
rect 7660 -1740 7670 -1700
rect 7610 -1765 7670 -1740
rect 7610 -1805 7620 -1765
rect 7660 -1805 7670 -1765
rect 7610 -1835 7670 -1805
rect 7610 -1875 7620 -1835
rect 7660 -1875 7670 -1835
rect 7610 -1905 7670 -1875
rect 7610 -1945 7620 -1905
rect 7660 -1945 7670 -1905
rect 7610 -1975 7670 -1945
rect 7610 -2015 7620 -1975
rect 7660 -2015 7670 -1975
rect 7610 -2040 7670 -2015
rect 7610 -2080 7620 -2040
rect 7660 -2080 7670 -2040
rect 7610 -2100 7670 -2080
rect 7610 -2140 7620 -2100
rect 7660 -2140 7670 -2100
rect 7610 -2165 7670 -2140
rect 7610 -2205 7620 -2165
rect 7660 -2205 7670 -2165
rect 7610 -2235 7670 -2205
rect 7610 -2275 7620 -2235
rect 7660 -2275 7670 -2235
rect 7610 -2305 7670 -2275
rect 7610 -2345 7620 -2305
rect 7660 -2345 7670 -2305
rect 7610 -2375 7670 -2345
rect 7610 -2415 7620 -2375
rect 7660 -2415 7670 -2375
rect 7610 -2440 7670 -2415
rect 7610 -2480 7620 -2440
rect 7660 -2480 7670 -2440
rect 7610 -2500 7670 -2480
rect 7610 -2540 7620 -2500
rect 7660 -2540 7670 -2500
rect 7610 -2565 7670 -2540
rect 7610 -2605 7620 -2565
rect 7660 -2605 7670 -2565
rect 7610 -2635 7670 -2605
rect 7610 -2675 7620 -2635
rect 7660 -2675 7670 -2635
rect 7610 -2705 7670 -2675
rect 7610 -2745 7620 -2705
rect 7660 -2745 7670 -2705
rect 7610 -2775 7670 -2745
rect 7610 -2815 7620 -2775
rect 7660 -2815 7670 -2775
rect 7610 -2840 7670 -2815
rect 7610 -2880 7620 -2840
rect 7660 -2880 7670 -2840
rect 7610 -2900 7670 -2880
rect 7610 -2940 7620 -2900
rect 7660 -2940 7670 -2900
rect 7610 -2965 7670 -2940
rect 7610 -3005 7620 -2965
rect 7660 -3005 7670 -2965
rect 7610 -3035 7670 -3005
rect 7610 -3075 7620 -3035
rect 7660 -3075 7670 -3035
rect 7610 -3105 7670 -3075
rect 7610 -3145 7620 -3105
rect 7660 -3145 7670 -3105
rect 7610 -3175 7670 -3145
rect 7610 -3215 7620 -3175
rect 7660 -3215 7670 -3175
rect 7610 -3240 7670 -3215
rect 7610 -3280 7620 -3240
rect 7660 -3280 7670 -3240
rect 7610 -3300 7670 -3280
rect 7610 -3340 7620 -3300
rect 7660 -3340 7670 -3300
rect 7610 -3365 7670 -3340
rect 7610 -3405 7620 -3365
rect 7660 -3405 7670 -3365
rect 7610 -3435 7670 -3405
rect 7610 -3475 7620 -3435
rect 7660 -3475 7670 -3435
rect 7610 -3505 7670 -3475
rect 7610 -3545 7620 -3505
rect 7660 -3545 7670 -3505
rect 7610 -3575 7670 -3545
rect 7610 -3615 7620 -3575
rect 7660 -3615 7670 -3575
rect 7610 -3640 7670 -3615
rect 7610 -3680 7620 -3640
rect 7660 -3680 7670 -3640
rect 7610 -3700 7670 -3680
rect 7610 -3740 7620 -3700
rect 7660 -3740 7670 -3700
rect 7610 -3765 7670 -3740
rect 7610 -3805 7620 -3765
rect 7660 -3805 7670 -3765
rect 7610 -3835 7670 -3805
rect 7610 -3875 7620 -3835
rect 7660 -3875 7670 -3835
rect 7610 -3905 7670 -3875
rect 7610 -3945 7620 -3905
rect 7660 -3945 7670 -3905
rect 7610 -3975 7670 -3945
rect 7610 -4015 7620 -3975
rect 7660 -4015 7670 -3975
rect 7610 -4040 7670 -4015
rect 7610 -4080 7620 -4040
rect 7660 -4080 7670 -4040
rect 7610 -4100 7670 -4080
rect 7610 -4140 7620 -4100
rect 7660 -4140 7670 -4100
rect 7610 -4165 7670 -4140
rect 7610 -4205 7620 -4165
rect 7660 -4205 7670 -4165
rect 7610 -4235 7670 -4205
rect 7610 -4275 7620 -4235
rect 7660 -4275 7670 -4235
rect 7610 -4305 7670 -4275
rect 7610 -4345 7620 -4305
rect 7660 -4345 7670 -4305
rect 7610 -4375 7670 -4345
rect 7610 -4415 7620 -4375
rect 7660 -4415 7670 -4375
rect 7610 -4440 7670 -4415
rect 7610 -4480 7620 -4440
rect 7660 -4480 7670 -4440
rect 7610 -4490 7670 -4480
rect 7960 -1300 8020 -1290
rect 7960 -1340 7970 -1300
rect 8010 -1340 8020 -1300
rect 7960 -1365 8020 -1340
rect 7960 -1405 7970 -1365
rect 8010 -1405 8020 -1365
rect 7960 -1435 8020 -1405
rect 7960 -1475 7970 -1435
rect 8010 -1475 8020 -1435
rect 7960 -1505 8020 -1475
rect 7960 -1545 7970 -1505
rect 8010 -1545 8020 -1505
rect 7960 -1575 8020 -1545
rect 7960 -1615 7970 -1575
rect 8010 -1615 8020 -1575
rect 7960 -1640 8020 -1615
rect 7960 -1680 7970 -1640
rect 8010 -1680 8020 -1640
rect 7960 -1700 8020 -1680
rect 7960 -1740 7970 -1700
rect 8010 -1740 8020 -1700
rect 7960 -1765 8020 -1740
rect 7960 -1805 7970 -1765
rect 8010 -1805 8020 -1765
rect 7960 -1835 8020 -1805
rect 7960 -1875 7970 -1835
rect 8010 -1875 8020 -1835
rect 7960 -1905 8020 -1875
rect 7960 -1945 7970 -1905
rect 8010 -1945 8020 -1905
rect 7960 -1975 8020 -1945
rect 7960 -2015 7970 -1975
rect 8010 -2015 8020 -1975
rect 7960 -2040 8020 -2015
rect 7960 -2080 7970 -2040
rect 8010 -2080 8020 -2040
rect 7960 -2100 8020 -2080
rect 7960 -2140 7970 -2100
rect 8010 -2140 8020 -2100
rect 7960 -2165 8020 -2140
rect 7960 -2205 7970 -2165
rect 8010 -2205 8020 -2165
rect 7960 -2235 8020 -2205
rect 7960 -2275 7970 -2235
rect 8010 -2275 8020 -2235
rect 7960 -2305 8020 -2275
rect 7960 -2345 7970 -2305
rect 8010 -2345 8020 -2305
rect 7960 -2375 8020 -2345
rect 7960 -2415 7970 -2375
rect 8010 -2415 8020 -2375
rect 7960 -2440 8020 -2415
rect 7960 -2480 7970 -2440
rect 8010 -2480 8020 -2440
rect 7960 -2500 8020 -2480
rect 7960 -2540 7970 -2500
rect 8010 -2540 8020 -2500
rect 7960 -2565 8020 -2540
rect 7960 -2605 7970 -2565
rect 8010 -2605 8020 -2565
rect 7960 -2635 8020 -2605
rect 7960 -2675 7970 -2635
rect 8010 -2675 8020 -2635
rect 7960 -2705 8020 -2675
rect 7960 -2745 7970 -2705
rect 8010 -2745 8020 -2705
rect 7960 -2775 8020 -2745
rect 7960 -2815 7970 -2775
rect 8010 -2815 8020 -2775
rect 7960 -2840 8020 -2815
rect 7960 -2880 7970 -2840
rect 8010 -2880 8020 -2840
rect 7960 -2900 8020 -2880
rect 7960 -2940 7970 -2900
rect 8010 -2940 8020 -2900
rect 7960 -2965 8020 -2940
rect 7960 -3005 7970 -2965
rect 8010 -3005 8020 -2965
rect 7960 -3035 8020 -3005
rect 7960 -3075 7970 -3035
rect 8010 -3075 8020 -3035
rect 7960 -3105 8020 -3075
rect 7960 -3145 7970 -3105
rect 8010 -3145 8020 -3105
rect 7960 -3175 8020 -3145
rect 7960 -3215 7970 -3175
rect 8010 -3215 8020 -3175
rect 7960 -3240 8020 -3215
rect 7960 -3280 7970 -3240
rect 8010 -3280 8020 -3240
rect 7960 -3300 8020 -3280
rect 7960 -3340 7970 -3300
rect 8010 -3340 8020 -3300
rect 7960 -3365 8020 -3340
rect 7960 -3405 7970 -3365
rect 8010 -3405 8020 -3365
rect 7960 -3435 8020 -3405
rect 7960 -3475 7970 -3435
rect 8010 -3475 8020 -3435
rect 7960 -3505 8020 -3475
rect 7960 -3545 7970 -3505
rect 8010 -3545 8020 -3505
rect 7960 -3575 8020 -3545
rect 7960 -3615 7970 -3575
rect 8010 -3615 8020 -3575
rect 7960 -3640 8020 -3615
rect 7960 -3680 7970 -3640
rect 8010 -3680 8020 -3640
rect 7960 -3700 8020 -3680
rect 7960 -3740 7970 -3700
rect 8010 -3740 8020 -3700
rect 7960 -3765 8020 -3740
rect 7960 -3805 7970 -3765
rect 8010 -3805 8020 -3765
rect 7960 -3835 8020 -3805
rect 7960 -3875 7970 -3835
rect 8010 -3875 8020 -3835
rect 7960 -3905 8020 -3875
rect 7960 -3945 7970 -3905
rect 8010 -3945 8020 -3905
rect 7960 -3975 8020 -3945
rect 7960 -4015 7970 -3975
rect 8010 -4015 8020 -3975
rect 7960 -4040 8020 -4015
rect 7960 -4080 7970 -4040
rect 8010 -4080 8020 -4040
rect 7960 -4100 8020 -4080
rect 7960 -4140 7970 -4100
rect 8010 -4140 8020 -4100
rect 7960 -4165 8020 -4140
rect 7960 -4205 7970 -4165
rect 8010 -4205 8020 -4165
rect 7960 -4235 8020 -4205
rect 7960 -4275 7970 -4235
rect 8010 -4275 8020 -4235
rect 7960 -4305 8020 -4275
rect 7960 -4345 7970 -4305
rect 8010 -4345 8020 -4305
rect 7960 -4375 8020 -4345
rect 7960 -4415 7970 -4375
rect 8010 -4415 8020 -4375
rect 7960 -4440 8020 -4415
rect 7960 -4480 7970 -4440
rect 8010 -4480 8020 -4440
rect 7960 -4490 8020 -4480
rect 8310 -1300 8370 -1290
rect 8310 -1340 8320 -1300
rect 8360 -1340 8370 -1300
rect 8310 -1365 8370 -1340
rect 8310 -1405 8320 -1365
rect 8360 -1405 8370 -1365
rect 8310 -1435 8370 -1405
rect 8310 -1475 8320 -1435
rect 8360 -1475 8370 -1435
rect 8310 -1505 8370 -1475
rect 8310 -1545 8320 -1505
rect 8360 -1545 8370 -1505
rect 8310 -1575 8370 -1545
rect 8310 -1615 8320 -1575
rect 8360 -1615 8370 -1575
rect 8310 -1640 8370 -1615
rect 8310 -1680 8320 -1640
rect 8360 -1680 8370 -1640
rect 8310 -1700 8370 -1680
rect 8310 -1740 8320 -1700
rect 8360 -1740 8370 -1700
rect 8310 -1765 8370 -1740
rect 8310 -1805 8320 -1765
rect 8360 -1805 8370 -1765
rect 8310 -1835 8370 -1805
rect 8310 -1875 8320 -1835
rect 8360 -1875 8370 -1835
rect 8310 -1905 8370 -1875
rect 8310 -1945 8320 -1905
rect 8360 -1945 8370 -1905
rect 8310 -1975 8370 -1945
rect 8310 -2015 8320 -1975
rect 8360 -2015 8370 -1975
rect 8310 -2040 8370 -2015
rect 8310 -2080 8320 -2040
rect 8360 -2080 8370 -2040
rect 8310 -2100 8370 -2080
rect 8310 -2140 8320 -2100
rect 8360 -2140 8370 -2100
rect 8310 -2165 8370 -2140
rect 8310 -2205 8320 -2165
rect 8360 -2205 8370 -2165
rect 8310 -2235 8370 -2205
rect 8310 -2275 8320 -2235
rect 8360 -2275 8370 -2235
rect 8310 -2305 8370 -2275
rect 8310 -2345 8320 -2305
rect 8360 -2345 8370 -2305
rect 8310 -2375 8370 -2345
rect 8310 -2415 8320 -2375
rect 8360 -2415 8370 -2375
rect 8310 -2440 8370 -2415
rect 8310 -2480 8320 -2440
rect 8360 -2480 8370 -2440
rect 8310 -2500 8370 -2480
rect 8310 -2540 8320 -2500
rect 8360 -2540 8370 -2500
rect 8310 -2565 8370 -2540
rect 8310 -2605 8320 -2565
rect 8360 -2605 8370 -2565
rect 8310 -2635 8370 -2605
rect 8310 -2675 8320 -2635
rect 8360 -2675 8370 -2635
rect 8310 -2705 8370 -2675
rect 8310 -2745 8320 -2705
rect 8360 -2745 8370 -2705
rect 8310 -2775 8370 -2745
rect 8310 -2815 8320 -2775
rect 8360 -2815 8370 -2775
rect 8310 -2840 8370 -2815
rect 8310 -2880 8320 -2840
rect 8360 -2880 8370 -2840
rect 8310 -2900 8370 -2880
rect 8310 -2940 8320 -2900
rect 8360 -2940 8370 -2900
rect 8310 -2965 8370 -2940
rect 8310 -3005 8320 -2965
rect 8360 -3005 8370 -2965
rect 8310 -3035 8370 -3005
rect 8310 -3075 8320 -3035
rect 8360 -3075 8370 -3035
rect 8310 -3105 8370 -3075
rect 8310 -3145 8320 -3105
rect 8360 -3145 8370 -3105
rect 8310 -3175 8370 -3145
rect 8310 -3215 8320 -3175
rect 8360 -3215 8370 -3175
rect 8310 -3240 8370 -3215
rect 8310 -3280 8320 -3240
rect 8360 -3280 8370 -3240
rect 8310 -3300 8370 -3280
rect 8310 -3340 8320 -3300
rect 8360 -3340 8370 -3300
rect 8310 -3365 8370 -3340
rect 8310 -3405 8320 -3365
rect 8360 -3405 8370 -3365
rect 8310 -3435 8370 -3405
rect 8310 -3475 8320 -3435
rect 8360 -3475 8370 -3435
rect 8310 -3505 8370 -3475
rect 8310 -3545 8320 -3505
rect 8360 -3545 8370 -3505
rect 8310 -3575 8370 -3545
rect 8310 -3615 8320 -3575
rect 8360 -3615 8370 -3575
rect 8310 -3640 8370 -3615
rect 8310 -3680 8320 -3640
rect 8360 -3680 8370 -3640
rect 8310 -3700 8370 -3680
rect 8310 -3740 8320 -3700
rect 8360 -3740 8370 -3700
rect 8310 -3765 8370 -3740
rect 8310 -3805 8320 -3765
rect 8360 -3805 8370 -3765
rect 8310 -3835 8370 -3805
rect 8310 -3875 8320 -3835
rect 8360 -3875 8370 -3835
rect 8310 -3905 8370 -3875
rect 8310 -3945 8320 -3905
rect 8360 -3945 8370 -3905
rect 8310 -3975 8370 -3945
rect 8310 -4015 8320 -3975
rect 8360 -4015 8370 -3975
rect 8310 -4040 8370 -4015
rect 8310 -4080 8320 -4040
rect 8360 -4080 8370 -4040
rect 8310 -4100 8370 -4080
rect 8310 -4140 8320 -4100
rect 8360 -4140 8370 -4100
rect 8310 -4165 8370 -4140
rect 8310 -4205 8320 -4165
rect 8360 -4205 8370 -4165
rect 8310 -4235 8370 -4205
rect 8310 -4275 8320 -4235
rect 8360 -4275 8370 -4235
rect 8310 -4305 8370 -4275
rect 8310 -4345 8320 -4305
rect 8360 -4345 8370 -4305
rect 8310 -4375 8370 -4345
rect 8310 -4415 8320 -4375
rect 8360 -4415 8370 -4375
rect 8310 -4440 8370 -4415
rect 8310 -4480 8320 -4440
rect 8360 -4480 8370 -4440
rect 8310 -4490 8370 -4480
rect 8660 -1300 8720 -1290
rect 8660 -1340 8670 -1300
rect 8710 -1340 8720 -1300
rect 8660 -1365 8720 -1340
rect 8660 -1405 8670 -1365
rect 8710 -1405 8720 -1365
rect 8660 -1435 8720 -1405
rect 8660 -1475 8670 -1435
rect 8710 -1475 8720 -1435
rect 8660 -1505 8720 -1475
rect 8660 -1545 8670 -1505
rect 8710 -1545 8720 -1505
rect 8660 -1575 8720 -1545
rect 8660 -1615 8670 -1575
rect 8710 -1615 8720 -1575
rect 8660 -1640 8720 -1615
rect 8660 -1680 8670 -1640
rect 8710 -1680 8720 -1640
rect 8660 -1700 8720 -1680
rect 8660 -1740 8670 -1700
rect 8710 -1740 8720 -1700
rect 8660 -1765 8720 -1740
rect 8660 -1805 8670 -1765
rect 8710 -1805 8720 -1765
rect 8660 -1835 8720 -1805
rect 8660 -1875 8670 -1835
rect 8710 -1875 8720 -1835
rect 8660 -1905 8720 -1875
rect 8660 -1945 8670 -1905
rect 8710 -1945 8720 -1905
rect 8660 -1975 8720 -1945
rect 8660 -2015 8670 -1975
rect 8710 -2015 8720 -1975
rect 8660 -2040 8720 -2015
rect 8660 -2080 8670 -2040
rect 8710 -2080 8720 -2040
rect 8660 -2100 8720 -2080
rect 8660 -2140 8670 -2100
rect 8710 -2140 8720 -2100
rect 8660 -2165 8720 -2140
rect 8660 -2205 8670 -2165
rect 8710 -2205 8720 -2165
rect 8660 -2235 8720 -2205
rect 8660 -2275 8670 -2235
rect 8710 -2275 8720 -2235
rect 8660 -2305 8720 -2275
rect 8660 -2345 8670 -2305
rect 8710 -2345 8720 -2305
rect 8660 -2375 8720 -2345
rect 8660 -2415 8670 -2375
rect 8710 -2415 8720 -2375
rect 8660 -2440 8720 -2415
rect 8660 -2480 8670 -2440
rect 8710 -2480 8720 -2440
rect 8660 -2500 8720 -2480
rect 8660 -2540 8670 -2500
rect 8710 -2540 8720 -2500
rect 8660 -2565 8720 -2540
rect 8660 -2605 8670 -2565
rect 8710 -2605 8720 -2565
rect 8660 -2635 8720 -2605
rect 8660 -2675 8670 -2635
rect 8710 -2675 8720 -2635
rect 8660 -2705 8720 -2675
rect 8660 -2745 8670 -2705
rect 8710 -2745 8720 -2705
rect 8660 -2775 8720 -2745
rect 8660 -2815 8670 -2775
rect 8710 -2815 8720 -2775
rect 8660 -2840 8720 -2815
rect 8660 -2880 8670 -2840
rect 8710 -2880 8720 -2840
rect 8660 -2900 8720 -2880
rect 8660 -2940 8670 -2900
rect 8710 -2940 8720 -2900
rect 8660 -2965 8720 -2940
rect 8660 -3005 8670 -2965
rect 8710 -3005 8720 -2965
rect 8660 -3035 8720 -3005
rect 8660 -3075 8670 -3035
rect 8710 -3075 8720 -3035
rect 8660 -3105 8720 -3075
rect 8660 -3145 8670 -3105
rect 8710 -3145 8720 -3105
rect 8660 -3175 8720 -3145
rect 8660 -3215 8670 -3175
rect 8710 -3215 8720 -3175
rect 8660 -3240 8720 -3215
rect 8660 -3280 8670 -3240
rect 8710 -3280 8720 -3240
rect 8660 -3300 8720 -3280
rect 8660 -3340 8670 -3300
rect 8710 -3340 8720 -3300
rect 8660 -3365 8720 -3340
rect 8660 -3405 8670 -3365
rect 8710 -3405 8720 -3365
rect 8660 -3435 8720 -3405
rect 8660 -3475 8670 -3435
rect 8710 -3475 8720 -3435
rect 8660 -3505 8720 -3475
rect 8660 -3545 8670 -3505
rect 8710 -3545 8720 -3505
rect 8660 -3575 8720 -3545
rect 8660 -3615 8670 -3575
rect 8710 -3615 8720 -3575
rect 8660 -3640 8720 -3615
rect 8660 -3680 8670 -3640
rect 8710 -3680 8720 -3640
rect 8660 -3700 8720 -3680
rect 8660 -3740 8670 -3700
rect 8710 -3740 8720 -3700
rect 8660 -3765 8720 -3740
rect 8660 -3805 8670 -3765
rect 8710 -3805 8720 -3765
rect 8660 -3835 8720 -3805
rect 8660 -3875 8670 -3835
rect 8710 -3875 8720 -3835
rect 8660 -3905 8720 -3875
rect 8660 -3945 8670 -3905
rect 8710 -3945 8720 -3905
rect 8660 -3975 8720 -3945
rect 8660 -4015 8670 -3975
rect 8710 -4015 8720 -3975
rect 8660 -4040 8720 -4015
rect 8660 -4080 8670 -4040
rect 8710 -4080 8720 -4040
rect 8660 -4100 8720 -4080
rect 8660 -4140 8670 -4100
rect 8710 -4140 8720 -4100
rect 8660 -4165 8720 -4140
rect 8660 -4205 8670 -4165
rect 8710 -4205 8720 -4165
rect 8660 -4235 8720 -4205
rect 8660 -4275 8670 -4235
rect 8710 -4275 8720 -4235
rect 8660 -4305 8720 -4275
rect 8660 -4345 8670 -4305
rect 8710 -4345 8720 -4305
rect 8660 -4375 8720 -4345
rect 8660 -4415 8670 -4375
rect 8710 -4415 8720 -4375
rect 8660 -4440 8720 -4415
rect 8660 -4480 8670 -4440
rect 8710 -4480 8720 -4440
rect 8660 -4490 8720 -4480
rect 14790 -1325 17990 6485
rect 14790 -1375 14825 -1325
rect 14875 -1375 14920 -1325
rect 14970 -1375 15015 -1325
rect 15065 -1375 15115 -1325
rect 15165 -1375 15215 -1325
rect 15265 -1375 15315 -1325
rect 15365 -1375 15410 -1325
rect 15460 -1375 15505 -1325
rect 15555 -1375 15625 -1325
rect 15675 -1375 15720 -1325
rect 15770 -1375 15815 -1325
rect 15865 -1375 15915 -1325
rect 15965 -1375 16015 -1325
rect 16065 -1375 16115 -1325
rect 16165 -1375 16210 -1325
rect 16260 -1375 16305 -1325
rect 16355 -1375 16425 -1325
rect 16475 -1375 16520 -1325
rect 16570 -1375 16615 -1325
rect 16665 -1375 16715 -1325
rect 16765 -1375 16815 -1325
rect 16865 -1375 16915 -1325
rect 16965 -1375 17010 -1325
rect 17060 -1375 17105 -1325
rect 17155 -1375 17225 -1325
rect 17275 -1375 17320 -1325
rect 17370 -1375 17415 -1325
rect 17465 -1375 17515 -1325
rect 17565 -1375 17615 -1325
rect 17665 -1375 17715 -1325
rect 17765 -1375 17810 -1325
rect 17860 -1375 17905 -1325
rect 17955 -1375 17990 -1325
rect 14790 -1415 17990 -1375
rect 14790 -1465 14825 -1415
rect 14875 -1465 14920 -1415
rect 14970 -1465 15015 -1415
rect 15065 -1465 15115 -1415
rect 15165 -1465 15215 -1415
rect 15265 -1465 15315 -1415
rect 15365 -1465 15410 -1415
rect 15460 -1465 15505 -1415
rect 15555 -1465 15625 -1415
rect 15675 -1465 15720 -1415
rect 15770 -1465 15815 -1415
rect 15865 -1465 15915 -1415
rect 15965 -1465 16015 -1415
rect 16065 -1465 16115 -1415
rect 16165 -1465 16210 -1415
rect 16260 -1465 16305 -1415
rect 16355 -1465 16425 -1415
rect 16475 -1465 16520 -1415
rect 16570 -1465 16615 -1415
rect 16665 -1465 16715 -1415
rect 16765 -1465 16815 -1415
rect 16865 -1465 16915 -1415
rect 16965 -1465 17010 -1415
rect 17060 -1465 17105 -1415
rect 17155 -1465 17225 -1415
rect 17275 -1465 17320 -1415
rect 17370 -1465 17415 -1415
rect 17465 -1465 17515 -1415
rect 17565 -1465 17615 -1415
rect 17665 -1465 17715 -1415
rect 17765 -1465 17810 -1415
rect 17860 -1465 17905 -1415
rect 17955 -1465 17990 -1415
rect 14790 -1515 17990 -1465
rect 14790 -1565 14825 -1515
rect 14875 -1565 14920 -1515
rect 14970 -1565 15015 -1515
rect 15065 -1565 15115 -1515
rect 15165 -1565 15215 -1515
rect 15265 -1565 15315 -1515
rect 15365 -1565 15410 -1515
rect 15460 -1565 15505 -1515
rect 15555 -1565 15625 -1515
rect 15675 -1565 15720 -1515
rect 15770 -1565 15815 -1515
rect 15865 -1565 15915 -1515
rect 15965 -1565 16015 -1515
rect 16065 -1565 16115 -1515
rect 16165 -1565 16210 -1515
rect 16260 -1565 16305 -1515
rect 16355 -1565 16425 -1515
rect 16475 -1565 16520 -1515
rect 16570 -1565 16615 -1515
rect 16665 -1565 16715 -1515
rect 16765 -1565 16815 -1515
rect 16865 -1565 16915 -1515
rect 16965 -1565 17010 -1515
rect 17060 -1565 17105 -1515
rect 17155 -1565 17225 -1515
rect 17275 -1565 17320 -1515
rect 17370 -1565 17415 -1515
rect 17465 -1565 17515 -1515
rect 17565 -1565 17615 -1515
rect 17665 -1565 17715 -1515
rect 17765 -1565 17810 -1515
rect 17860 -1565 17905 -1515
rect 17955 -1565 17990 -1515
rect 14790 -1605 17990 -1565
rect 14790 -1655 14825 -1605
rect 14875 -1655 14920 -1605
rect 14970 -1655 15015 -1605
rect 15065 -1655 15115 -1605
rect 15165 -1655 15215 -1605
rect 15265 -1655 15315 -1605
rect 15365 -1655 15410 -1605
rect 15460 -1655 15505 -1605
rect 15555 -1655 15625 -1605
rect 15675 -1655 15720 -1605
rect 15770 -1655 15815 -1605
rect 15865 -1655 15915 -1605
rect 15965 -1655 16015 -1605
rect 16065 -1655 16115 -1605
rect 16165 -1655 16210 -1605
rect 16260 -1655 16305 -1605
rect 16355 -1655 16425 -1605
rect 16475 -1655 16520 -1605
rect 16570 -1655 16615 -1605
rect 16665 -1655 16715 -1605
rect 16765 -1655 16815 -1605
rect 16865 -1655 16915 -1605
rect 16965 -1655 17010 -1605
rect 17060 -1655 17105 -1605
rect 17155 -1655 17225 -1605
rect 17275 -1655 17320 -1605
rect 17370 -1655 17415 -1605
rect 17465 -1655 17515 -1605
rect 17565 -1655 17615 -1605
rect 17665 -1655 17715 -1605
rect 17765 -1655 17810 -1605
rect 17860 -1655 17905 -1605
rect 17955 -1655 17990 -1605
rect 14790 -1725 17990 -1655
rect 14790 -1775 14825 -1725
rect 14875 -1775 14920 -1725
rect 14970 -1775 15015 -1725
rect 15065 -1775 15115 -1725
rect 15165 -1775 15215 -1725
rect 15265 -1775 15315 -1725
rect 15365 -1775 15410 -1725
rect 15460 -1775 15505 -1725
rect 15555 -1775 15625 -1725
rect 15675 -1775 15720 -1725
rect 15770 -1775 15815 -1725
rect 15865 -1775 15915 -1725
rect 15965 -1775 16015 -1725
rect 16065 -1775 16115 -1725
rect 16165 -1775 16210 -1725
rect 16260 -1775 16305 -1725
rect 16355 -1775 16425 -1725
rect 16475 -1775 16520 -1725
rect 16570 -1775 16615 -1725
rect 16665 -1775 16715 -1725
rect 16765 -1775 16815 -1725
rect 16865 -1775 16915 -1725
rect 16965 -1775 17010 -1725
rect 17060 -1775 17105 -1725
rect 17155 -1775 17225 -1725
rect 17275 -1775 17320 -1725
rect 17370 -1775 17415 -1725
rect 17465 -1775 17515 -1725
rect 17565 -1775 17615 -1725
rect 17665 -1775 17715 -1725
rect 17765 -1775 17810 -1725
rect 17860 -1775 17905 -1725
rect 17955 -1775 17990 -1725
rect 14790 -1815 17990 -1775
rect 14790 -1865 14825 -1815
rect 14875 -1865 14920 -1815
rect 14970 -1865 15015 -1815
rect 15065 -1865 15115 -1815
rect 15165 -1865 15215 -1815
rect 15265 -1865 15315 -1815
rect 15365 -1865 15410 -1815
rect 15460 -1865 15505 -1815
rect 15555 -1865 15625 -1815
rect 15675 -1865 15720 -1815
rect 15770 -1865 15815 -1815
rect 15865 -1865 15915 -1815
rect 15965 -1865 16015 -1815
rect 16065 -1865 16115 -1815
rect 16165 -1865 16210 -1815
rect 16260 -1865 16305 -1815
rect 16355 -1865 16425 -1815
rect 16475 -1865 16520 -1815
rect 16570 -1865 16615 -1815
rect 16665 -1865 16715 -1815
rect 16765 -1865 16815 -1815
rect 16865 -1865 16915 -1815
rect 16965 -1865 17010 -1815
rect 17060 -1865 17105 -1815
rect 17155 -1865 17225 -1815
rect 17275 -1865 17320 -1815
rect 17370 -1865 17415 -1815
rect 17465 -1865 17515 -1815
rect 17565 -1865 17615 -1815
rect 17665 -1865 17715 -1815
rect 17765 -1865 17810 -1815
rect 17860 -1865 17905 -1815
rect 17955 -1865 17990 -1815
rect 14790 -1915 17990 -1865
rect 14790 -1965 14825 -1915
rect 14875 -1965 14920 -1915
rect 14970 -1965 15015 -1915
rect 15065 -1965 15115 -1915
rect 15165 -1965 15215 -1915
rect 15265 -1965 15315 -1915
rect 15365 -1965 15410 -1915
rect 15460 -1965 15505 -1915
rect 15555 -1965 15625 -1915
rect 15675 -1965 15720 -1915
rect 15770 -1965 15815 -1915
rect 15865 -1965 15915 -1915
rect 15965 -1965 16015 -1915
rect 16065 -1965 16115 -1915
rect 16165 -1965 16210 -1915
rect 16260 -1965 16305 -1915
rect 16355 -1965 16425 -1915
rect 16475 -1965 16520 -1915
rect 16570 -1965 16615 -1915
rect 16665 -1965 16715 -1915
rect 16765 -1965 16815 -1915
rect 16865 -1965 16915 -1915
rect 16965 -1965 17010 -1915
rect 17060 -1965 17105 -1915
rect 17155 -1965 17225 -1915
rect 17275 -1965 17320 -1915
rect 17370 -1965 17415 -1915
rect 17465 -1965 17515 -1915
rect 17565 -1965 17615 -1915
rect 17665 -1965 17715 -1915
rect 17765 -1965 17810 -1915
rect 17860 -1965 17905 -1915
rect 17955 -1965 17990 -1915
rect 14790 -2005 17990 -1965
rect 14790 -2055 14825 -2005
rect 14875 -2055 14920 -2005
rect 14970 -2055 15015 -2005
rect 15065 -2055 15115 -2005
rect 15165 -2055 15215 -2005
rect 15265 -2055 15315 -2005
rect 15365 -2055 15410 -2005
rect 15460 -2055 15505 -2005
rect 15555 -2055 15625 -2005
rect 15675 -2055 15720 -2005
rect 15770 -2055 15815 -2005
rect 15865 -2055 15915 -2005
rect 15965 -2055 16015 -2005
rect 16065 -2055 16115 -2005
rect 16165 -2055 16210 -2005
rect 16260 -2055 16305 -2005
rect 16355 -2055 16425 -2005
rect 16475 -2055 16520 -2005
rect 16570 -2055 16615 -2005
rect 16665 -2055 16715 -2005
rect 16765 -2055 16815 -2005
rect 16865 -2055 16915 -2005
rect 16965 -2055 17010 -2005
rect 17060 -2055 17105 -2005
rect 17155 -2055 17225 -2005
rect 17275 -2055 17320 -2005
rect 17370 -2055 17415 -2005
rect 17465 -2055 17515 -2005
rect 17565 -2055 17615 -2005
rect 17665 -2055 17715 -2005
rect 17765 -2055 17810 -2005
rect 17860 -2055 17905 -2005
rect 17955 -2055 17990 -2005
rect 14790 -2125 17990 -2055
rect 14790 -2175 14825 -2125
rect 14875 -2175 14920 -2125
rect 14970 -2175 15015 -2125
rect 15065 -2175 15115 -2125
rect 15165 -2175 15215 -2125
rect 15265 -2175 15315 -2125
rect 15365 -2175 15410 -2125
rect 15460 -2175 15505 -2125
rect 15555 -2175 15625 -2125
rect 15675 -2175 15720 -2125
rect 15770 -2175 15815 -2125
rect 15865 -2175 15915 -2125
rect 15965 -2175 16015 -2125
rect 16065 -2175 16115 -2125
rect 16165 -2175 16210 -2125
rect 16260 -2175 16305 -2125
rect 16355 -2175 16425 -2125
rect 16475 -2175 16520 -2125
rect 16570 -2175 16615 -2125
rect 16665 -2175 16715 -2125
rect 16765 -2175 16815 -2125
rect 16865 -2175 16915 -2125
rect 16965 -2175 17010 -2125
rect 17060 -2175 17105 -2125
rect 17155 -2175 17225 -2125
rect 17275 -2175 17320 -2125
rect 17370 -2175 17415 -2125
rect 17465 -2175 17515 -2125
rect 17565 -2175 17615 -2125
rect 17665 -2175 17715 -2125
rect 17765 -2175 17810 -2125
rect 17860 -2175 17905 -2125
rect 17955 -2175 17990 -2125
rect 14790 -2215 17990 -2175
rect 14790 -2265 14825 -2215
rect 14875 -2265 14920 -2215
rect 14970 -2265 15015 -2215
rect 15065 -2265 15115 -2215
rect 15165 -2265 15215 -2215
rect 15265 -2265 15315 -2215
rect 15365 -2265 15410 -2215
rect 15460 -2265 15505 -2215
rect 15555 -2265 15625 -2215
rect 15675 -2265 15720 -2215
rect 15770 -2265 15815 -2215
rect 15865 -2265 15915 -2215
rect 15965 -2265 16015 -2215
rect 16065 -2265 16115 -2215
rect 16165 -2265 16210 -2215
rect 16260 -2265 16305 -2215
rect 16355 -2265 16425 -2215
rect 16475 -2265 16520 -2215
rect 16570 -2265 16615 -2215
rect 16665 -2265 16715 -2215
rect 16765 -2265 16815 -2215
rect 16865 -2265 16915 -2215
rect 16965 -2265 17010 -2215
rect 17060 -2265 17105 -2215
rect 17155 -2265 17225 -2215
rect 17275 -2265 17320 -2215
rect 17370 -2265 17415 -2215
rect 17465 -2265 17515 -2215
rect 17565 -2265 17615 -2215
rect 17665 -2265 17715 -2215
rect 17765 -2265 17810 -2215
rect 17860 -2265 17905 -2215
rect 17955 -2265 17990 -2215
rect 14790 -2315 17990 -2265
rect 14790 -2365 14825 -2315
rect 14875 -2365 14920 -2315
rect 14970 -2365 15015 -2315
rect 15065 -2365 15115 -2315
rect 15165 -2365 15215 -2315
rect 15265 -2365 15315 -2315
rect 15365 -2365 15410 -2315
rect 15460 -2365 15505 -2315
rect 15555 -2365 15625 -2315
rect 15675 -2365 15720 -2315
rect 15770 -2365 15815 -2315
rect 15865 -2365 15915 -2315
rect 15965 -2365 16015 -2315
rect 16065 -2365 16115 -2315
rect 16165 -2365 16210 -2315
rect 16260 -2365 16305 -2315
rect 16355 -2365 16425 -2315
rect 16475 -2365 16520 -2315
rect 16570 -2365 16615 -2315
rect 16665 -2365 16715 -2315
rect 16765 -2365 16815 -2315
rect 16865 -2365 16915 -2315
rect 16965 -2365 17010 -2315
rect 17060 -2365 17105 -2315
rect 17155 -2365 17225 -2315
rect 17275 -2365 17320 -2315
rect 17370 -2365 17415 -2315
rect 17465 -2365 17515 -2315
rect 17565 -2365 17615 -2315
rect 17665 -2365 17715 -2315
rect 17765 -2365 17810 -2315
rect 17860 -2365 17905 -2315
rect 17955 -2365 17990 -2315
rect 14790 -2405 17990 -2365
rect 14790 -2455 14825 -2405
rect 14875 -2455 14920 -2405
rect 14970 -2455 15015 -2405
rect 15065 -2455 15115 -2405
rect 15165 -2455 15215 -2405
rect 15265 -2455 15315 -2405
rect 15365 -2455 15410 -2405
rect 15460 -2455 15505 -2405
rect 15555 -2455 15625 -2405
rect 15675 -2455 15720 -2405
rect 15770 -2455 15815 -2405
rect 15865 -2455 15915 -2405
rect 15965 -2455 16015 -2405
rect 16065 -2455 16115 -2405
rect 16165 -2455 16210 -2405
rect 16260 -2455 16305 -2405
rect 16355 -2455 16425 -2405
rect 16475 -2455 16520 -2405
rect 16570 -2455 16615 -2405
rect 16665 -2455 16715 -2405
rect 16765 -2455 16815 -2405
rect 16865 -2455 16915 -2405
rect 16965 -2455 17010 -2405
rect 17060 -2455 17105 -2405
rect 17155 -2455 17225 -2405
rect 17275 -2455 17320 -2405
rect 17370 -2455 17415 -2405
rect 17465 -2455 17515 -2405
rect 17565 -2455 17615 -2405
rect 17665 -2455 17715 -2405
rect 17765 -2455 17810 -2405
rect 17860 -2455 17905 -2405
rect 17955 -2455 17990 -2405
rect 14790 -2525 17990 -2455
rect 14790 -2575 14825 -2525
rect 14875 -2575 14920 -2525
rect 14970 -2575 15015 -2525
rect 15065 -2575 15115 -2525
rect 15165 -2575 15215 -2525
rect 15265 -2575 15315 -2525
rect 15365 -2575 15410 -2525
rect 15460 -2575 15505 -2525
rect 15555 -2575 15625 -2525
rect 15675 -2575 15720 -2525
rect 15770 -2575 15815 -2525
rect 15865 -2575 15915 -2525
rect 15965 -2575 16015 -2525
rect 16065 -2575 16115 -2525
rect 16165 -2575 16210 -2525
rect 16260 -2575 16305 -2525
rect 16355 -2575 16425 -2525
rect 16475 -2575 16520 -2525
rect 16570 -2575 16615 -2525
rect 16665 -2575 16715 -2525
rect 16765 -2575 16815 -2525
rect 16865 -2575 16915 -2525
rect 16965 -2575 17010 -2525
rect 17060 -2575 17105 -2525
rect 17155 -2575 17225 -2525
rect 17275 -2575 17320 -2525
rect 17370 -2575 17415 -2525
rect 17465 -2575 17515 -2525
rect 17565 -2575 17615 -2525
rect 17665 -2575 17715 -2525
rect 17765 -2575 17810 -2525
rect 17860 -2575 17905 -2525
rect 17955 -2575 17990 -2525
rect 14790 -2615 17990 -2575
rect 14790 -2665 14825 -2615
rect 14875 -2665 14920 -2615
rect 14970 -2665 15015 -2615
rect 15065 -2665 15115 -2615
rect 15165 -2665 15215 -2615
rect 15265 -2665 15315 -2615
rect 15365 -2665 15410 -2615
rect 15460 -2665 15505 -2615
rect 15555 -2665 15625 -2615
rect 15675 -2665 15720 -2615
rect 15770 -2665 15815 -2615
rect 15865 -2665 15915 -2615
rect 15965 -2665 16015 -2615
rect 16065 -2665 16115 -2615
rect 16165 -2665 16210 -2615
rect 16260 -2665 16305 -2615
rect 16355 -2665 16425 -2615
rect 16475 -2665 16520 -2615
rect 16570 -2665 16615 -2615
rect 16665 -2665 16715 -2615
rect 16765 -2665 16815 -2615
rect 16865 -2665 16915 -2615
rect 16965 -2665 17010 -2615
rect 17060 -2665 17105 -2615
rect 17155 -2665 17225 -2615
rect 17275 -2665 17320 -2615
rect 17370 -2665 17415 -2615
rect 17465 -2665 17515 -2615
rect 17565 -2665 17615 -2615
rect 17665 -2665 17715 -2615
rect 17765 -2665 17810 -2615
rect 17860 -2665 17905 -2615
rect 17955 -2665 17990 -2615
rect 14790 -2715 17990 -2665
rect 14790 -2765 14825 -2715
rect 14875 -2765 14920 -2715
rect 14970 -2765 15015 -2715
rect 15065 -2765 15115 -2715
rect 15165 -2765 15215 -2715
rect 15265 -2765 15315 -2715
rect 15365 -2765 15410 -2715
rect 15460 -2765 15505 -2715
rect 15555 -2765 15625 -2715
rect 15675 -2765 15720 -2715
rect 15770 -2765 15815 -2715
rect 15865 -2765 15915 -2715
rect 15965 -2765 16015 -2715
rect 16065 -2765 16115 -2715
rect 16165 -2765 16210 -2715
rect 16260 -2765 16305 -2715
rect 16355 -2765 16425 -2715
rect 16475 -2765 16520 -2715
rect 16570 -2765 16615 -2715
rect 16665 -2765 16715 -2715
rect 16765 -2765 16815 -2715
rect 16865 -2765 16915 -2715
rect 16965 -2765 17010 -2715
rect 17060 -2765 17105 -2715
rect 17155 -2765 17225 -2715
rect 17275 -2765 17320 -2715
rect 17370 -2765 17415 -2715
rect 17465 -2765 17515 -2715
rect 17565 -2765 17615 -2715
rect 17665 -2765 17715 -2715
rect 17765 -2765 17810 -2715
rect 17860 -2765 17905 -2715
rect 17955 -2765 17990 -2715
rect 14790 -2805 17990 -2765
rect 14790 -2855 14825 -2805
rect 14875 -2855 14920 -2805
rect 14970 -2855 15015 -2805
rect 15065 -2855 15115 -2805
rect 15165 -2855 15215 -2805
rect 15265 -2855 15315 -2805
rect 15365 -2855 15410 -2805
rect 15460 -2855 15505 -2805
rect 15555 -2855 15625 -2805
rect 15675 -2855 15720 -2805
rect 15770 -2855 15815 -2805
rect 15865 -2855 15915 -2805
rect 15965 -2855 16015 -2805
rect 16065 -2855 16115 -2805
rect 16165 -2855 16210 -2805
rect 16260 -2855 16305 -2805
rect 16355 -2855 16425 -2805
rect 16475 -2855 16520 -2805
rect 16570 -2855 16615 -2805
rect 16665 -2855 16715 -2805
rect 16765 -2855 16815 -2805
rect 16865 -2855 16915 -2805
rect 16965 -2855 17010 -2805
rect 17060 -2855 17105 -2805
rect 17155 -2855 17225 -2805
rect 17275 -2855 17320 -2805
rect 17370 -2855 17415 -2805
rect 17465 -2855 17515 -2805
rect 17565 -2855 17615 -2805
rect 17665 -2855 17715 -2805
rect 17765 -2855 17810 -2805
rect 17860 -2855 17905 -2805
rect 17955 -2855 17990 -2805
rect 14790 -2925 17990 -2855
rect 14790 -2975 14825 -2925
rect 14875 -2975 14920 -2925
rect 14970 -2975 15015 -2925
rect 15065 -2975 15115 -2925
rect 15165 -2975 15215 -2925
rect 15265 -2975 15315 -2925
rect 15365 -2975 15410 -2925
rect 15460 -2975 15505 -2925
rect 15555 -2975 15625 -2925
rect 15675 -2975 15720 -2925
rect 15770 -2975 15815 -2925
rect 15865 -2975 15915 -2925
rect 15965 -2975 16015 -2925
rect 16065 -2975 16115 -2925
rect 16165 -2975 16210 -2925
rect 16260 -2975 16305 -2925
rect 16355 -2975 16425 -2925
rect 16475 -2975 16520 -2925
rect 16570 -2975 16615 -2925
rect 16665 -2975 16715 -2925
rect 16765 -2975 16815 -2925
rect 16865 -2975 16915 -2925
rect 16965 -2975 17010 -2925
rect 17060 -2975 17105 -2925
rect 17155 -2975 17225 -2925
rect 17275 -2975 17320 -2925
rect 17370 -2975 17415 -2925
rect 17465 -2975 17515 -2925
rect 17565 -2975 17615 -2925
rect 17665 -2975 17715 -2925
rect 17765 -2975 17810 -2925
rect 17860 -2975 17905 -2925
rect 17955 -2975 17990 -2925
rect 14790 -3015 17990 -2975
rect 14790 -3065 14825 -3015
rect 14875 -3065 14920 -3015
rect 14970 -3065 15015 -3015
rect 15065 -3065 15115 -3015
rect 15165 -3065 15215 -3015
rect 15265 -3065 15315 -3015
rect 15365 -3065 15410 -3015
rect 15460 -3065 15505 -3015
rect 15555 -3065 15625 -3015
rect 15675 -3065 15720 -3015
rect 15770 -3065 15815 -3015
rect 15865 -3065 15915 -3015
rect 15965 -3065 16015 -3015
rect 16065 -3065 16115 -3015
rect 16165 -3065 16210 -3015
rect 16260 -3065 16305 -3015
rect 16355 -3065 16425 -3015
rect 16475 -3065 16520 -3015
rect 16570 -3065 16615 -3015
rect 16665 -3065 16715 -3015
rect 16765 -3065 16815 -3015
rect 16865 -3065 16915 -3015
rect 16965 -3065 17010 -3015
rect 17060 -3065 17105 -3015
rect 17155 -3065 17225 -3015
rect 17275 -3065 17320 -3015
rect 17370 -3065 17415 -3015
rect 17465 -3065 17515 -3015
rect 17565 -3065 17615 -3015
rect 17665 -3065 17715 -3015
rect 17765 -3065 17810 -3015
rect 17860 -3065 17905 -3015
rect 17955 -3065 17990 -3015
rect 14790 -3115 17990 -3065
rect 14790 -3165 14825 -3115
rect 14875 -3165 14920 -3115
rect 14970 -3165 15015 -3115
rect 15065 -3165 15115 -3115
rect 15165 -3165 15215 -3115
rect 15265 -3165 15315 -3115
rect 15365 -3165 15410 -3115
rect 15460 -3165 15505 -3115
rect 15555 -3165 15625 -3115
rect 15675 -3165 15720 -3115
rect 15770 -3165 15815 -3115
rect 15865 -3165 15915 -3115
rect 15965 -3165 16015 -3115
rect 16065 -3165 16115 -3115
rect 16165 -3165 16210 -3115
rect 16260 -3165 16305 -3115
rect 16355 -3165 16425 -3115
rect 16475 -3165 16520 -3115
rect 16570 -3165 16615 -3115
rect 16665 -3165 16715 -3115
rect 16765 -3165 16815 -3115
rect 16865 -3165 16915 -3115
rect 16965 -3165 17010 -3115
rect 17060 -3165 17105 -3115
rect 17155 -3165 17225 -3115
rect 17275 -3165 17320 -3115
rect 17370 -3165 17415 -3115
rect 17465 -3165 17515 -3115
rect 17565 -3165 17615 -3115
rect 17665 -3165 17715 -3115
rect 17765 -3165 17810 -3115
rect 17860 -3165 17905 -3115
rect 17955 -3165 17990 -3115
rect 14790 -3205 17990 -3165
rect 14790 -3255 14825 -3205
rect 14875 -3255 14920 -3205
rect 14970 -3255 15015 -3205
rect 15065 -3255 15115 -3205
rect 15165 -3255 15215 -3205
rect 15265 -3255 15315 -3205
rect 15365 -3255 15410 -3205
rect 15460 -3255 15505 -3205
rect 15555 -3255 15625 -3205
rect 15675 -3255 15720 -3205
rect 15770 -3255 15815 -3205
rect 15865 -3255 15915 -3205
rect 15965 -3255 16015 -3205
rect 16065 -3255 16115 -3205
rect 16165 -3255 16210 -3205
rect 16260 -3255 16305 -3205
rect 16355 -3255 16425 -3205
rect 16475 -3255 16520 -3205
rect 16570 -3255 16615 -3205
rect 16665 -3255 16715 -3205
rect 16765 -3255 16815 -3205
rect 16865 -3255 16915 -3205
rect 16965 -3255 17010 -3205
rect 17060 -3255 17105 -3205
rect 17155 -3255 17225 -3205
rect 17275 -3255 17320 -3205
rect 17370 -3255 17415 -3205
rect 17465 -3255 17515 -3205
rect 17565 -3255 17615 -3205
rect 17665 -3255 17715 -3205
rect 17765 -3255 17810 -3205
rect 17860 -3255 17905 -3205
rect 17955 -3255 17990 -3205
rect 14790 -3325 17990 -3255
rect 14790 -3375 14825 -3325
rect 14875 -3375 14920 -3325
rect 14970 -3375 15015 -3325
rect 15065 -3375 15115 -3325
rect 15165 -3375 15215 -3325
rect 15265 -3375 15315 -3325
rect 15365 -3375 15410 -3325
rect 15460 -3375 15505 -3325
rect 15555 -3375 15625 -3325
rect 15675 -3375 15720 -3325
rect 15770 -3375 15815 -3325
rect 15865 -3375 15915 -3325
rect 15965 -3375 16015 -3325
rect 16065 -3375 16115 -3325
rect 16165 -3375 16210 -3325
rect 16260 -3375 16305 -3325
rect 16355 -3375 16425 -3325
rect 16475 -3375 16520 -3325
rect 16570 -3375 16615 -3325
rect 16665 -3375 16715 -3325
rect 16765 -3375 16815 -3325
rect 16865 -3375 16915 -3325
rect 16965 -3375 17010 -3325
rect 17060 -3375 17105 -3325
rect 17155 -3375 17225 -3325
rect 17275 -3375 17320 -3325
rect 17370 -3375 17415 -3325
rect 17465 -3375 17515 -3325
rect 17565 -3375 17615 -3325
rect 17665 -3375 17715 -3325
rect 17765 -3375 17810 -3325
rect 17860 -3375 17905 -3325
rect 17955 -3375 17990 -3325
rect 14790 -3415 17990 -3375
rect 14790 -3465 14825 -3415
rect 14875 -3465 14920 -3415
rect 14970 -3465 15015 -3415
rect 15065 -3465 15115 -3415
rect 15165 -3465 15215 -3415
rect 15265 -3465 15315 -3415
rect 15365 -3465 15410 -3415
rect 15460 -3465 15505 -3415
rect 15555 -3465 15625 -3415
rect 15675 -3465 15720 -3415
rect 15770 -3465 15815 -3415
rect 15865 -3465 15915 -3415
rect 15965 -3465 16015 -3415
rect 16065 -3465 16115 -3415
rect 16165 -3465 16210 -3415
rect 16260 -3465 16305 -3415
rect 16355 -3465 16425 -3415
rect 16475 -3465 16520 -3415
rect 16570 -3465 16615 -3415
rect 16665 -3465 16715 -3415
rect 16765 -3465 16815 -3415
rect 16865 -3465 16915 -3415
rect 16965 -3465 17010 -3415
rect 17060 -3465 17105 -3415
rect 17155 -3465 17225 -3415
rect 17275 -3465 17320 -3415
rect 17370 -3465 17415 -3415
rect 17465 -3465 17515 -3415
rect 17565 -3465 17615 -3415
rect 17665 -3465 17715 -3415
rect 17765 -3465 17810 -3415
rect 17860 -3465 17905 -3415
rect 17955 -3465 17990 -3415
rect 14790 -3515 17990 -3465
rect 14790 -3565 14825 -3515
rect 14875 -3565 14920 -3515
rect 14970 -3565 15015 -3515
rect 15065 -3565 15115 -3515
rect 15165 -3565 15215 -3515
rect 15265 -3565 15315 -3515
rect 15365 -3565 15410 -3515
rect 15460 -3565 15505 -3515
rect 15555 -3565 15625 -3515
rect 15675 -3565 15720 -3515
rect 15770 -3565 15815 -3515
rect 15865 -3565 15915 -3515
rect 15965 -3565 16015 -3515
rect 16065 -3565 16115 -3515
rect 16165 -3565 16210 -3515
rect 16260 -3565 16305 -3515
rect 16355 -3565 16425 -3515
rect 16475 -3565 16520 -3515
rect 16570 -3565 16615 -3515
rect 16665 -3565 16715 -3515
rect 16765 -3565 16815 -3515
rect 16865 -3565 16915 -3515
rect 16965 -3565 17010 -3515
rect 17060 -3565 17105 -3515
rect 17155 -3565 17225 -3515
rect 17275 -3565 17320 -3515
rect 17370 -3565 17415 -3515
rect 17465 -3565 17515 -3515
rect 17565 -3565 17615 -3515
rect 17665 -3565 17715 -3515
rect 17765 -3565 17810 -3515
rect 17860 -3565 17905 -3515
rect 17955 -3565 17990 -3515
rect 14790 -3605 17990 -3565
rect 14790 -3655 14825 -3605
rect 14875 -3655 14920 -3605
rect 14970 -3655 15015 -3605
rect 15065 -3655 15115 -3605
rect 15165 -3655 15215 -3605
rect 15265 -3655 15315 -3605
rect 15365 -3655 15410 -3605
rect 15460 -3655 15505 -3605
rect 15555 -3655 15625 -3605
rect 15675 -3655 15720 -3605
rect 15770 -3655 15815 -3605
rect 15865 -3655 15915 -3605
rect 15965 -3655 16015 -3605
rect 16065 -3655 16115 -3605
rect 16165 -3655 16210 -3605
rect 16260 -3655 16305 -3605
rect 16355 -3655 16425 -3605
rect 16475 -3655 16520 -3605
rect 16570 -3655 16615 -3605
rect 16665 -3655 16715 -3605
rect 16765 -3655 16815 -3605
rect 16865 -3655 16915 -3605
rect 16965 -3655 17010 -3605
rect 17060 -3655 17105 -3605
rect 17155 -3655 17225 -3605
rect 17275 -3655 17320 -3605
rect 17370 -3655 17415 -3605
rect 17465 -3655 17515 -3605
rect 17565 -3655 17615 -3605
rect 17665 -3655 17715 -3605
rect 17765 -3655 17810 -3605
rect 17860 -3655 17905 -3605
rect 17955 -3655 17990 -3605
rect 14790 -3725 17990 -3655
rect 14790 -3775 14825 -3725
rect 14875 -3775 14920 -3725
rect 14970 -3775 15015 -3725
rect 15065 -3775 15115 -3725
rect 15165 -3775 15215 -3725
rect 15265 -3775 15315 -3725
rect 15365 -3775 15410 -3725
rect 15460 -3775 15505 -3725
rect 15555 -3775 15625 -3725
rect 15675 -3775 15720 -3725
rect 15770 -3775 15815 -3725
rect 15865 -3775 15915 -3725
rect 15965 -3775 16015 -3725
rect 16065 -3775 16115 -3725
rect 16165 -3775 16210 -3725
rect 16260 -3775 16305 -3725
rect 16355 -3775 16425 -3725
rect 16475 -3775 16520 -3725
rect 16570 -3775 16615 -3725
rect 16665 -3775 16715 -3725
rect 16765 -3775 16815 -3725
rect 16865 -3775 16915 -3725
rect 16965 -3775 17010 -3725
rect 17060 -3775 17105 -3725
rect 17155 -3775 17225 -3725
rect 17275 -3775 17320 -3725
rect 17370 -3775 17415 -3725
rect 17465 -3775 17515 -3725
rect 17565 -3775 17615 -3725
rect 17665 -3775 17715 -3725
rect 17765 -3775 17810 -3725
rect 17860 -3775 17905 -3725
rect 17955 -3775 17990 -3725
rect 14790 -3815 17990 -3775
rect 14790 -3865 14825 -3815
rect 14875 -3865 14920 -3815
rect 14970 -3865 15015 -3815
rect 15065 -3865 15115 -3815
rect 15165 -3865 15215 -3815
rect 15265 -3865 15315 -3815
rect 15365 -3865 15410 -3815
rect 15460 -3865 15505 -3815
rect 15555 -3865 15625 -3815
rect 15675 -3865 15720 -3815
rect 15770 -3865 15815 -3815
rect 15865 -3865 15915 -3815
rect 15965 -3865 16015 -3815
rect 16065 -3865 16115 -3815
rect 16165 -3865 16210 -3815
rect 16260 -3865 16305 -3815
rect 16355 -3865 16425 -3815
rect 16475 -3865 16520 -3815
rect 16570 -3865 16615 -3815
rect 16665 -3865 16715 -3815
rect 16765 -3865 16815 -3815
rect 16865 -3865 16915 -3815
rect 16965 -3865 17010 -3815
rect 17060 -3865 17105 -3815
rect 17155 -3865 17225 -3815
rect 17275 -3865 17320 -3815
rect 17370 -3865 17415 -3815
rect 17465 -3865 17515 -3815
rect 17565 -3865 17615 -3815
rect 17665 -3865 17715 -3815
rect 17765 -3865 17810 -3815
rect 17860 -3865 17905 -3815
rect 17955 -3865 17990 -3815
rect 14790 -3915 17990 -3865
rect 14790 -3965 14825 -3915
rect 14875 -3965 14920 -3915
rect 14970 -3965 15015 -3915
rect 15065 -3965 15115 -3915
rect 15165 -3965 15215 -3915
rect 15265 -3965 15315 -3915
rect 15365 -3965 15410 -3915
rect 15460 -3965 15505 -3915
rect 15555 -3965 15625 -3915
rect 15675 -3965 15720 -3915
rect 15770 -3965 15815 -3915
rect 15865 -3965 15915 -3915
rect 15965 -3965 16015 -3915
rect 16065 -3965 16115 -3915
rect 16165 -3965 16210 -3915
rect 16260 -3965 16305 -3915
rect 16355 -3965 16425 -3915
rect 16475 -3965 16520 -3915
rect 16570 -3965 16615 -3915
rect 16665 -3965 16715 -3915
rect 16765 -3965 16815 -3915
rect 16865 -3965 16915 -3915
rect 16965 -3965 17010 -3915
rect 17060 -3965 17105 -3915
rect 17155 -3965 17225 -3915
rect 17275 -3965 17320 -3915
rect 17370 -3965 17415 -3915
rect 17465 -3965 17515 -3915
rect 17565 -3965 17615 -3915
rect 17665 -3965 17715 -3915
rect 17765 -3965 17810 -3915
rect 17860 -3965 17905 -3915
rect 17955 -3965 17990 -3915
rect 14790 -4005 17990 -3965
rect 14790 -4055 14825 -4005
rect 14875 -4055 14920 -4005
rect 14970 -4055 15015 -4005
rect 15065 -4055 15115 -4005
rect 15165 -4055 15215 -4005
rect 15265 -4055 15315 -4005
rect 15365 -4055 15410 -4005
rect 15460 -4055 15505 -4005
rect 15555 -4055 15625 -4005
rect 15675 -4055 15720 -4005
rect 15770 -4055 15815 -4005
rect 15865 -4055 15915 -4005
rect 15965 -4055 16015 -4005
rect 16065 -4055 16115 -4005
rect 16165 -4055 16210 -4005
rect 16260 -4055 16305 -4005
rect 16355 -4055 16425 -4005
rect 16475 -4055 16520 -4005
rect 16570 -4055 16615 -4005
rect 16665 -4055 16715 -4005
rect 16765 -4055 16815 -4005
rect 16865 -4055 16915 -4005
rect 16965 -4055 17010 -4005
rect 17060 -4055 17105 -4005
rect 17155 -4055 17225 -4005
rect 17275 -4055 17320 -4005
rect 17370 -4055 17415 -4005
rect 17465 -4055 17515 -4005
rect 17565 -4055 17615 -4005
rect 17665 -4055 17715 -4005
rect 17765 -4055 17810 -4005
rect 17860 -4055 17905 -4005
rect 17955 -4055 17990 -4005
rect 14790 -4125 17990 -4055
rect 14790 -4175 14825 -4125
rect 14875 -4175 14920 -4125
rect 14970 -4175 15015 -4125
rect 15065 -4175 15115 -4125
rect 15165 -4175 15215 -4125
rect 15265 -4175 15315 -4125
rect 15365 -4175 15410 -4125
rect 15460 -4175 15505 -4125
rect 15555 -4175 15625 -4125
rect 15675 -4175 15720 -4125
rect 15770 -4175 15815 -4125
rect 15865 -4175 15915 -4125
rect 15965 -4175 16015 -4125
rect 16065 -4175 16115 -4125
rect 16165 -4175 16210 -4125
rect 16260 -4175 16305 -4125
rect 16355 -4175 16425 -4125
rect 16475 -4175 16520 -4125
rect 16570 -4175 16615 -4125
rect 16665 -4175 16715 -4125
rect 16765 -4175 16815 -4125
rect 16865 -4175 16915 -4125
rect 16965 -4175 17010 -4125
rect 17060 -4175 17105 -4125
rect 17155 -4175 17225 -4125
rect 17275 -4175 17320 -4125
rect 17370 -4175 17415 -4125
rect 17465 -4175 17515 -4125
rect 17565 -4175 17615 -4125
rect 17665 -4175 17715 -4125
rect 17765 -4175 17810 -4125
rect 17860 -4175 17905 -4125
rect 17955 -4175 17990 -4125
rect 14790 -4215 17990 -4175
rect 14790 -4265 14825 -4215
rect 14875 -4265 14920 -4215
rect 14970 -4265 15015 -4215
rect 15065 -4265 15115 -4215
rect 15165 -4265 15215 -4215
rect 15265 -4265 15315 -4215
rect 15365 -4265 15410 -4215
rect 15460 -4265 15505 -4215
rect 15555 -4265 15625 -4215
rect 15675 -4265 15720 -4215
rect 15770 -4265 15815 -4215
rect 15865 -4265 15915 -4215
rect 15965 -4265 16015 -4215
rect 16065 -4265 16115 -4215
rect 16165 -4265 16210 -4215
rect 16260 -4265 16305 -4215
rect 16355 -4265 16425 -4215
rect 16475 -4265 16520 -4215
rect 16570 -4265 16615 -4215
rect 16665 -4265 16715 -4215
rect 16765 -4265 16815 -4215
rect 16865 -4265 16915 -4215
rect 16965 -4265 17010 -4215
rect 17060 -4265 17105 -4215
rect 17155 -4265 17225 -4215
rect 17275 -4265 17320 -4215
rect 17370 -4265 17415 -4215
rect 17465 -4265 17515 -4215
rect 17565 -4265 17615 -4215
rect 17665 -4265 17715 -4215
rect 17765 -4265 17810 -4215
rect 17860 -4265 17905 -4215
rect 17955 -4265 17990 -4215
rect 14790 -4315 17990 -4265
rect 14790 -4365 14825 -4315
rect 14875 -4365 14920 -4315
rect 14970 -4365 15015 -4315
rect 15065 -4365 15115 -4315
rect 15165 -4365 15215 -4315
rect 15265 -4365 15315 -4315
rect 15365 -4365 15410 -4315
rect 15460 -4365 15505 -4315
rect 15555 -4365 15625 -4315
rect 15675 -4365 15720 -4315
rect 15770 -4365 15815 -4315
rect 15865 -4365 15915 -4315
rect 15965 -4365 16015 -4315
rect 16065 -4365 16115 -4315
rect 16165 -4365 16210 -4315
rect 16260 -4365 16305 -4315
rect 16355 -4365 16425 -4315
rect 16475 -4365 16520 -4315
rect 16570 -4365 16615 -4315
rect 16665 -4365 16715 -4315
rect 16765 -4365 16815 -4315
rect 16865 -4365 16915 -4315
rect 16965 -4365 17010 -4315
rect 17060 -4365 17105 -4315
rect 17155 -4365 17225 -4315
rect 17275 -4365 17320 -4315
rect 17370 -4365 17415 -4315
rect 17465 -4365 17515 -4315
rect 17565 -4365 17615 -4315
rect 17665 -4365 17715 -4315
rect 17765 -4365 17810 -4315
rect 17860 -4365 17905 -4315
rect 17955 -4365 17990 -4315
rect 14790 -4405 17990 -4365
rect 14790 -4455 14825 -4405
rect 14875 -4455 14920 -4405
rect 14970 -4455 15015 -4405
rect 15065 -4455 15115 -4405
rect 15165 -4455 15215 -4405
rect 15265 -4455 15315 -4405
rect 15365 -4455 15410 -4405
rect 15460 -4455 15505 -4405
rect 15555 -4455 15625 -4405
rect 15675 -4455 15720 -4405
rect 15770 -4455 15815 -4405
rect 15865 -4455 15915 -4405
rect 15965 -4455 16015 -4405
rect 16065 -4455 16115 -4405
rect 16165 -4455 16210 -4405
rect 16260 -4455 16305 -4405
rect 16355 -4455 16425 -4405
rect 16475 -4455 16520 -4405
rect 16570 -4455 16615 -4405
rect 16665 -4455 16715 -4405
rect 16765 -4455 16815 -4405
rect 16865 -4455 16915 -4405
rect 16965 -4455 17010 -4405
rect 17060 -4455 17105 -4405
rect 17155 -4455 17225 -4405
rect 17275 -4455 17320 -4405
rect 17370 -4455 17415 -4405
rect 17465 -4455 17515 -4405
rect 17565 -4455 17615 -4405
rect 17665 -4455 17715 -4405
rect 17765 -4455 17810 -4405
rect 17860 -4455 17905 -4405
rect 17955 -4455 17990 -4405
rect 14790 -4490 17990 -4455
<< via3 >>
rect 2330 20910 2370 20915
rect 2330 20880 2335 20910
rect 2335 20880 2365 20910
rect 2365 20880 2370 20910
rect 2330 20875 2370 20880
rect 2330 20845 2370 20850
rect 2330 20815 2335 20845
rect 2335 20815 2365 20845
rect 2365 20815 2370 20845
rect 2330 20810 2370 20815
rect 2330 20775 2370 20780
rect 2330 20745 2335 20775
rect 2335 20745 2365 20775
rect 2365 20745 2370 20775
rect 2330 20740 2370 20745
rect 2330 20705 2370 20710
rect 2330 20675 2335 20705
rect 2335 20675 2365 20705
rect 2365 20675 2370 20705
rect 2330 20670 2370 20675
rect 2330 20635 2370 20640
rect 2330 20605 2335 20635
rect 2335 20605 2365 20635
rect 2365 20605 2370 20635
rect 2330 20600 2370 20605
rect 2330 20570 2370 20575
rect 2330 20540 2335 20570
rect 2335 20540 2365 20570
rect 2365 20540 2370 20570
rect 2330 20535 2370 20540
rect 2330 20510 2370 20515
rect 2330 20480 2335 20510
rect 2335 20480 2365 20510
rect 2365 20480 2370 20510
rect 2330 20475 2370 20480
rect 2330 20445 2370 20450
rect 2330 20415 2335 20445
rect 2335 20415 2365 20445
rect 2365 20415 2370 20445
rect 2330 20410 2370 20415
rect 2330 20375 2370 20380
rect 2330 20345 2335 20375
rect 2335 20345 2365 20375
rect 2365 20345 2370 20375
rect 2330 20340 2370 20345
rect 2330 20305 2370 20310
rect 2330 20275 2335 20305
rect 2335 20275 2365 20305
rect 2365 20275 2370 20305
rect 2330 20270 2370 20275
rect 2330 20235 2370 20240
rect 2330 20205 2335 20235
rect 2335 20205 2365 20235
rect 2365 20205 2370 20235
rect 2330 20200 2370 20205
rect 2330 20170 2370 20175
rect 2330 20140 2335 20170
rect 2335 20140 2365 20170
rect 2365 20140 2370 20170
rect 2330 20135 2370 20140
rect 2330 20110 2370 20115
rect 2330 20080 2335 20110
rect 2335 20080 2365 20110
rect 2365 20080 2370 20110
rect 2330 20075 2370 20080
rect 2330 20045 2370 20050
rect 2330 20015 2335 20045
rect 2335 20015 2365 20045
rect 2365 20015 2370 20045
rect 2330 20010 2370 20015
rect 2330 19975 2370 19980
rect 2330 19945 2335 19975
rect 2335 19945 2365 19975
rect 2365 19945 2370 19975
rect 2330 19940 2370 19945
rect 2330 19905 2370 19910
rect 2330 19875 2335 19905
rect 2335 19875 2365 19905
rect 2365 19875 2370 19905
rect 2330 19870 2370 19875
rect 2330 19835 2370 19840
rect 2330 19805 2335 19835
rect 2335 19805 2365 19835
rect 2365 19805 2370 19835
rect 2330 19800 2370 19805
rect 2330 19770 2370 19775
rect 2330 19740 2335 19770
rect 2335 19740 2365 19770
rect 2365 19740 2370 19770
rect 2330 19735 2370 19740
rect 2330 19710 2370 19715
rect 2330 19680 2335 19710
rect 2335 19680 2365 19710
rect 2365 19680 2370 19710
rect 2330 19675 2370 19680
rect 2330 19645 2370 19650
rect 2330 19615 2335 19645
rect 2335 19615 2365 19645
rect 2365 19615 2370 19645
rect 2330 19610 2370 19615
rect 2330 19575 2370 19580
rect 2330 19545 2335 19575
rect 2335 19545 2365 19575
rect 2365 19545 2370 19575
rect 2330 19540 2370 19545
rect 2330 19505 2370 19510
rect 2330 19475 2335 19505
rect 2335 19475 2365 19505
rect 2365 19475 2370 19505
rect 2330 19470 2370 19475
rect 2330 19435 2370 19440
rect 2330 19405 2335 19435
rect 2335 19405 2365 19435
rect 2365 19405 2370 19435
rect 2330 19400 2370 19405
rect 2330 19370 2370 19375
rect 2330 19340 2335 19370
rect 2335 19340 2365 19370
rect 2365 19340 2370 19370
rect 2330 19335 2370 19340
rect 2330 19310 2370 19315
rect 2330 19280 2335 19310
rect 2335 19280 2365 19310
rect 2365 19280 2370 19310
rect 2330 19275 2370 19280
rect 2330 19245 2370 19250
rect 2330 19215 2335 19245
rect 2335 19215 2365 19245
rect 2365 19215 2370 19245
rect 2330 19210 2370 19215
rect 2330 19175 2370 19180
rect 2330 19145 2335 19175
rect 2335 19145 2365 19175
rect 2365 19145 2370 19175
rect 2330 19140 2370 19145
rect 2330 19105 2370 19110
rect 2330 19075 2335 19105
rect 2335 19075 2365 19105
rect 2365 19075 2370 19105
rect 2330 19070 2370 19075
rect 2330 19035 2370 19040
rect 2330 19005 2335 19035
rect 2335 19005 2365 19035
rect 2365 19005 2370 19035
rect 2330 19000 2370 19005
rect 2330 18970 2370 18975
rect 2330 18940 2335 18970
rect 2335 18940 2365 18970
rect 2365 18940 2370 18970
rect 2330 18935 2370 18940
rect 2330 18910 2370 18915
rect 2330 18880 2335 18910
rect 2335 18880 2365 18910
rect 2365 18880 2370 18910
rect 2330 18875 2370 18880
rect 2330 18845 2370 18850
rect 2330 18815 2335 18845
rect 2335 18815 2365 18845
rect 2365 18815 2370 18845
rect 2330 18810 2370 18815
rect 2330 18775 2370 18780
rect 2330 18745 2335 18775
rect 2335 18745 2365 18775
rect 2365 18745 2370 18775
rect 2330 18740 2370 18745
rect 2330 18705 2370 18710
rect 2330 18675 2335 18705
rect 2335 18675 2365 18705
rect 2365 18675 2370 18705
rect 2330 18670 2370 18675
rect 2330 18635 2370 18640
rect 2330 18605 2335 18635
rect 2335 18605 2365 18635
rect 2365 18605 2370 18635
rect 2330 18600 2370 18605
rect 2330 18570 2370 18575
rect 2330 18540 2335 18570
rect 2335 18540 2365 18570
rect 2365 18540 2370 18570
rect 2330 18535 2370 18540
rect 2330 18510 2370 18515
rect 2330 18480 2335 18510
rect 2335 18480 2365 18510
rect 2365 18480 2370 18510
rect 2330 18475 2370 18480
rect 2330 18445 2370 18450
rect 2330 18415 2335 18445
rect 2335 18415 2365 18445
rect 2365 18415 2370 18445
rect 2330 18410 2370 18415
rect 2330 18375 2370 18380
rect 2330 18345 2335 18375
rect 2335 18345 2365 18375
rect 2365 18345 2370 18375
rect 2330 18340 2370 18345
rect 2330 18305 2370 18310
rect 2330 18275 2335 18305
rect 2335 18275 2365 18305
rect 2365 18275 2370 18305
rect 2330 18270 2370 18275
rect 2330 18235 2370 18240
rect 2330 18205 2335 18235
rect 2335 18205 2365 18235
rect 2365 18205 2370 18235
rect 2330 18200 2370 18205
rect 2330 18170 2370 18175
rect 2330 18140 2335 18170
rect 2335 18140 2365 18170
rect 2365 18140 2370 18170
rect 2330 18135 2370 18140
rect 2330 18110 2370 18115
rect 2330 18080 2335 18110
rect 2335 18080 2365 18110
rect 2365 18080 2370 18110
rect 2330 18075 2370 18080
rect 2330 18045 2370 18050
rect 2330 18015 2335 18045
rect 2335 18015 2365 18045
rect 2365 18015 2370 18045
rect 2330 18010 2370 18015
rect 2330 17975 2370 17980
rect 2330 17945 2335 17975
rect 2335 17945 2365 17975
rect 2365 17945 2370 17975
rect 2330 17940 2370 17945
rect 2330 17905 2370 17910
rect 2330 17875 2335 17905
rect 2335 17875 2365 17905
rect 2365 17875 2370 17905
rect 2330 17870 2370 17875
rect 2330 17835 2370 17840
rect 2330 17805 2335 17835
rect 2335 17805 2365 17835
rect 2365 17805 2370 17835
rect 2330 17800 2370 17805
rect 2330 17770 2370 17775
rect 2330 17740 2335 17770
rect 2335 17740 2365 17770
rect 2365 17740 2370 17770
rect 2330 17735 2370 17740
rect 6700 20910 6740 20915
rect 6700 20880 6705 20910
rect 6705 20880 6735 20910
rect 6735 20880 6740 20910
rect 6700 20875 6740 20880
rect 6700 20845 6740 20850
rect 6700 20815 6705 20845
rect 6705 20815 6735 20845
rect 6735 20815 6740 20845
rect 6700 20810 6740 20815
rect 6700 20775 6740 20780
rect 6700 20745 6705 20775
rect 6705 20745 6735 20775
rect 6735 20745 6740 20775
rect 6700 20740 6740 20745
rect 6700 20705 6740 20710
rect 6700 20675 6705 20705
rect 6705 20675 6735 20705
rect 6735 20675 6740 20705
rect 6700 20670 6740 20675
rect 6700 20635 6740 20640
rect 6700 20605 6705 20635
rect 6705 20605 6735 20635
rect 6735 20605 6740 20635
rect 6700 20600 6740 20605
rect 6700 20570 6740 20575
rect 6700 20540 6705 20570
rect 6705 20540 6735 20570
rect 6735 20540 6740 20570
rect 6700 20535 6740 20540
rect 6700 20510 6740 20515
rect 6700 20480 6705 20510
rect 6705 20480 6735 20510
rect 6735 20480 6740 20510
rect 6700 20475 6740 20480
rect 6700 20445 6740 20450
rect 6700 20415 6705 20445
rect 6705 20415 6735 20445
rect 6735 20415 6740 20445
rect 6700 20410 6740 20415
rect 6700 20375 6740 20380
rect 6700 20345 6705 20375
rect 6705 20345 6735 20375
rect 6735 20345 6740 20375
rect 6700 20340 6740 20345
rect 6700 20305 6740 20310
rect 6700 20275 6705 20305
rect 6705 20275 6735 20305
rect 6735 20275 6740 20305
rect 6700 20270 6740 20275
rect 6700 20235 6740 20240
rect 6700 20205 6705 20235
rect 6705 20205 6735 20235
rect 6735 20205 6740 20235
rect 6700 20200 6740 20205
rect 6700 20170 6740 20175
rect 6700 20140 6705 20170
rect 6705 20140 6735 20170
rect 6735 20140 6740 20170
rect 6700 20135 6740 20140
rect 6700 20110 6740 20115
rect 6700 20080 6705 20110
rect 6705 20080 6735 20110
rect 6735 20080 6740 20110
rect 6700 20075 6740 20080
rect 6700 20045 6740 20050
rect 6700 20015 6705 20045
rect 6705 20015 6735 20045
rect 6735 20015 6740 20045
rect 6700 20010 6740 20015
rect 6700 19975 6740 19980
rect 6700 19945 6705 19975
rect 6705 19945 6735 19975
rect 6735 19945 6740 19975
rect 6700 19940 6740 19945
rect 6700 19905 6740 19910
rect 6700 19875 6705 19905
rect 6705 19875 6735 19905
rect 6735 19875 6740 19905
rect 6700 19870 6740 19875
rect 6700 19835 6740 19840
rect 6700 19805 6705 19835
rect 6705 19805 6735 19835
rect 6735 19805 6740 19835
rect 6700 19800 6740 19805
rect 6700 19770 6740 19775
rect 6700 19740 6705 19770
rect 6705 19740 6735 19770
rect 6735 19740 6740 19770
rect 6700 19735 6740 19740
rect 6700 19710 6740 19715
rect 6700 19680 6705 19710
rect 6705 19680 6735 19710
rect 6735 19680 6740 19710
rect 6700 19675 6740 19680
rect 6700 19645 6740 19650
rect 6700 19615 6705 19645
rect 6705 19615 6735 19645
rect 6735 19615 6740 19645
rect 6700 19610 6740 19615
rect 6700 19575 6740 19580
rect 6700 19545 6705 19575
rect 6705 19545 6735 19575
rect 6735 19545 6740 19575
rect 6700 19540 6740 19545
rect 6700 19505 6740 19510
rect 6700 19475 6705 19505
rect 6705 19475 6735 19505
rect 6735 19475 6740 19505
rect 6700 19470 6740 19475
rect 6700 19435 6740 19440
rect 6700 19405 6705 19435
rect 6705 19405 6735 19435
rect 6735 19405 6740 19435
rect 6700 19400 6740 19405
rect 6700 19370 6740 19375
rect 6700 19340 6705 19370
rect 6705 19340 6735 19370
rect 6735 19340 6740 19370
rect 6700 19335 6740 19340
rect 6700 19310 6740 19315
rect 6700 19280 6705 19310
rect 6705 19280 6735 19310
rect 6735 19280 6740 19310
rect 6700 19275 6740 19280
rect 6700 19245 6740 19250
rect 6700 19215 6705 19245
rect 6705 19215 6735 19245
rect 6735 19215 6740 19245
rect 6700 19210 6740 19215
rect 6700 19175 6740 19180
rect 6700 19145 6705 19175
rect 6705 19145 6735 19175
rect 6735 19145 6740 19175
rect 6700 19140 6740 19145
rect 6700 19105 6740 19110
rect 6700 19075 6705 19105
rect 6705 19075 6735 19105
rect 6735 19075 6740 19105
rect 6700 19070 6740 19075
rect 6700 19035 6740 19040
rect 6700 19005 6705 19035
rect 6705 19005 6735 19035
rect 6735 19005 6740 19035
rect 6700 19000 6740 19005
rect 6700 18970 6740 18975
rect 6700 18940 6705 18970
rect 6705 18940 6735 18970
rect 6735 18940 6740 18970
rect 6700 18935 6740 18940
rect 6700 18910 6740 18915
rect 6700 18880 6705 18910
rect 6705 18880 6735 18910
rect 6735 18880 6740 18910
rect 6700 18875 6740 18880
rect 6700 18845 6740 18850
rect 6700 18815 6705 18845
rect 6705 18815 6735 18845
rect 6735 18815 6740 18845
rect 6700 18810 6740 18815
rect 6700 18775 6740 18780
rect 6700 18745 6705 18775
rect 6705 18745 6735 18775
rect 6735 18745 6740 18775
rect 6700 18740 6740 18745
rect 6700 18705 6740 18710
rect 6700 18675 6705 18705
rect 6705 18675 6735 18705
rect 6735 18675 6740 18705
rect 6700 18670 6740 18675
rect 6700 18635 6740 18640
rect 6700 18605 6705 18635
rect 6705 18605 6735 18635
rect 6735 18605 6740 18635
rect 6700 18600 6740 18605
rect 6700 18570 6740 18575
rect 6700 18540 6705 18570
rect 6705 18540 6735 18570
rect 6735 18540 6740 18570
rect 6700 18535 6740 18540
rect 6700 18510 6740 18515
rect 6700 18480 6705 18510
rect 6705 18480 6735 18510
rect 6735 18480 6740 18510
rect 6700 18475 6740 18480
rect 6700 18445 6740 18450
rect 6700 18415 6705 18445
rect 6705 18415 6735 18445
rect 6735 18415 6740 18445
rect 6700 18410 6740 18415
rect 6700 18375 6740 18380
rect 6700 18345 6705 18375
rect 6705 18345 6735 18375
rect 6735 18345 6740 18375
rect 6700 18340 6740 18345
rect 6700 18305 6740 18310
rect 6700 18275 6705 18305
rect 6705 18275 6735 18305
rect 6735 18275 6740 18305
rect 6700 18270 6740 18275
rect 6700 18235 6740 18240
rect 6700 18205 6705 18235
rect 6705 18205 6735 18235
rect 6735 18205 6740 18235
rect 6700 18200 6740 18205
rect 6700 18170 6740 18175
rect 6700 18140 6705 18170
rect 6705 18140 6735 18170
rect 6735 18140 6740 18170
rect 6700 18135 6740 18140
rect 6700 18110 6740 18115
rect 6700 18080 6705 18110
rect 6705 18080 6735 18110
rect 6735 18080 6740 18110
rect 6700 18075 6740 18080
rect 6700 18045 6740 18050
rect 6700 18015 6705 18045
rect 6705 18015 6735 18045
rect 6735 18015 6740 18045
rect 6700 18010 6740 18015
rect 6700 17975 6740 17980
rect 6700 17945 6705 17975
rect 6705 17945 6735 17975
rect 6735 17945 6740 17975
rect 6700 17940 6740 17945
rect 6700 17905 6740 17910
rect 6700 17875 6705 17905
rect 6705 17875 6735 17905
rect 6735 17875 6740 17905
rect 6700 17870 6740 17875
rect 6700 17835 6740 17840
rect 6700 17805 6705 17835
rect 6705 17805 6735 17835
rect 6735 17805 6740 17835
rect 6700 17800 6740 17805
rect 6700 17770 6740 17775
rect 6700 17740 6705 17770
rect 6705 17740 6735 17770
rect 6735 17740 6740 17770
rect 6700 17735 6740 17740
rect 14825 20840 14875 20890
rect 14920 20840 14970 20890
rect 15015 20840 15065 20890
rect 15115 20840 15165 20890
rect 15215 20840 15265 20890
rect 15315 20840 15365 20890
rect 15410 20840 15460 20890
rect 15505 20840 15555 20890
rect 15625 20840 15675 20890
rect 15720 20840 15770 20890
rect 15815 20840 15865 20890
rect 15915 20840 15965 20890
rect 16015 20840 16065 20890
rect 16115 20840 16165 20890
rect 16210 20840 16260 20890
rect 16305 20840 16355 20890
rect 16425 20840 16475 20890
rect 16520 20840 16570 20890
rect 16615 20840 16665 20890
rect 16715 20840 16765 20890
rect 16815 20840 16865 20890
rect 16915 20840 16965 20890
rect 17010 20840 17060 20890
rect 17105 20840 17155 20890
rect 17225 20840 17275 20890
rect 17320 20840 17370 20890
rect 17415 20840 17465 20890
rect 17515 20840 17565 20890
rect 17615 20840 17665 20890
rect 17715 20840 17765 20890
rect 17810 20840 17860 20890
rect 17905 20840 17955 20890
rect 14825 20750 14875 20800
rect 14920 20750 14970 20800
rect 15015 20750 15065 20800
rect 15115 20750 15165 20800
rect 15215 20750 15265 20800
rect 15315 20750 15365 20800
rect 15410 20750 15460 20800
rect 15505 20750 15555 20800
rect 15625 20750 15675 20800
rect 15720 20750 15770 20800
rect 15815 20750 15865 20800
rect 15915 20750 15965 20800
rect 16015 20750 16065 20800
rect 16115 20750 16165 20800
rect 16210 20750 16260 20800
rect 16305 20750 16355 20800
rect 16425 20750 16475 20800
rect 16520 20750 16570 20800
rect 16615 20750 16665 20800
rect 16715 20750 16765 20800
rect 16815 20750 16865 20800
rect 16915 20750 16965 20800
rect 17010 20750 17060 20800
rect 17105 20750 17155 20800
rect 17225 20750 17275 20800
rect 17320 20750 17370 20800
rect 17415 20750 17465 20800
rect 17515 20750 17565 20800
rect 17615 20750 17665 20800
rect 17715 20750 17765 20800
rect 17810 20750 17860 20800
rect 17905 20750 17955 20800
rect 14825 20650 14875 20700
rect 14920 20650 14970 20700
rect 15015 20650 15065 20700
rect 15115 20650 15165 20700
rect 15215 20650 15265 20700
rect 15315 20650 15365 20700
rect 15410 20650 15460 20700
rect 15505 20650 15555 20700
rect 15625 20650 15675 20700
rect 15720 20650 15770 20700
rect 15815 20650 15865 20700
rect 15915 20650 15965 20700
rect 16015 20650 16065 20700
rect 16115 20650 16165 20700
rect 16210 20650 16260 20700
rect 16305 20650 16355 20700
rect 16425 20650 16475 20700
rect 16520 20650 16570 20700
rect 16615 20650 16665 20700
rect 16715 20650 16765 20700
rect 16815 20650 16865 20700
rect 16915 20650 16965 20700
rect 17010 20650 17060 20700
rect 17105 20650 17155 20700
rect 17225 20650 17275 20700
rect 17320 20650 17370 20700
rect 17415 20650 17465 20700
rect 17515 20650 17565 20700
rect 17615 20650 17665 20700
rect 17715 20650 17765 20700
rect 17810 20650 17860 20700
rect 17905 20650 17955 20700
rect 14825 20560 14875 20610
rect 14920 20560 14970 20610
rect 15015 20560 15065 20610
rect 15115 20560 15165 20610
rect 15215 20560 15265 20610
rect 15315 20560 15365 20610
rect 15410 20560 15460 20610
rect 15505 20560 15555 20610
rect 15625 20560 15675 20610
rect 15720 20560 15770 20610
rect 15815 20560 15865 20610
rect 15915 20560 15965 20610
rect 16015 20560 16065 20610
rect 16115 20560 16165 20610
rect 16210 20560 16260 20610
rect 16305 20560 16355 20610
rect 16425 20560 16475 20610
rect 16520 20560 16570 20610
rect 16615 20560 16665 20610
rect 16715 20560 16765 20610
rect 16815 20560 16865 20610
rect 16915 20560 16965 20610
rect 17010 20560 17060 20610
rect 17105 20560 17155 20610
rect 17225 20560 17275 20610
rect 17320 20560 17370 20610
rect 17415 20560 17465 20610
rect 17515 20560 17565 20610
rect 17615 20560 17665 20610
rect 17715 20560 17765 20610
rect 17810 20560 17860 20610
rect 17905 20560 17955 20610
rect 14825 20440 14875 20490
rect 14920 20440 14970 20490
rect 15015 20440 15065 20490
rect 15115 20440 15165 20490
rect 15215 20440 15265 20490
rect 15315 20440 15365 20490
rect 15410 20440 15460 20490
rect 15505 20440 15555 20490
rect 15625 20440 15675 20490
rect 15720 20440 15770 20490
rect 15815 20440 15865 20490
rect 15915 20440 15965 20490
rect 16015 20440 16065 20490
rect 16115 20440 16165 20490
rect 16210 20440 16260 20490
rect 16305 20440 16355 20490
rect 16425 20440 16475 20490
rect 16520 20440 16570 20490
rect 16615 20440 16665 20490
rect 16715 20440 16765 20490
rect 16815 20440 16865 20490
rect 16915 20440 16965 20490
rect 17010 20440 17060 20490
rect 17105 20440 17155 20490
rect 17225 20440 17275 20490
rect 17320 20440 17370 20490
rect 17415 20440 17465 20490
rect 17515 20440 17565 20490
rect 17615 20440 17665 20490
rect 17715 20440 17765 20490
rect 17810 20440 17860 20490
rect 17905 20440 17955 20490
rect 14825 20350 14875 20400
rect 14920 20350 14970 20400
rect 15015 20350 15065 20400
rect 15115 20350 15165 20400
rect 15215 20350 15265 20400
rect 15315 20350 15365 20400
rect 15410 20350 15460 20400
rect 15505 20350 15555 20400
rect 15625 20350 15675 20400
rect 15720 20350 15770 20400
rect 15815 20350 15865 20400
rect 15915 20350 15965 20400
rect 16015 20350 16065 20400
rect 16115 20350 16165 20400
rect 16210 20350 16260 20400
rect 16305 20350 16355 20400
rect 16425 20350 16475 20400
rect 16520 20350 16570 20400
rect 16615 20350 16665 20400
rect 16715 20350 16765 20400
rect 16815 20350 16865 20400
rect 16915 20350 16965 20400
rect 17010 20350 17060 20400
rect 17105 20350 17155 20400
rect 17225 20350 17275 20400
rect 17320 20350 17370 20400
rect 17415 20350 17465 20400
rect 17515 20350 17565 20400
rect 17615 20350 17665 20400
rect 17715 20350 17765 20400
rect 17810 20350 17860 20400
rect 17905 20350 17955 20400
rect 14825 20250 14875 20300
rect 14920 20250 14970 20300
rect 15015 20250 15065 20300
rect 15115 20250 15165 20300
rect 15215 20250 15265 20300
rect 15315 20250 15365 20300
rect 15410 20250 15460 20300
rect 15505 20250 15555 20300
rect 15625 20250 15675 20300
rect 15720 20250 15770 20300
rect 15815 20250 15865 20300
rect 15915 20250 15965 20300
rect 16015 20250 16065 20300
rect 16115 20250 16165 20300
rect 16210 20250 16260 20300
rect 16305 20250 16355 20300
rect 16425 20250 16475 20300
rect 16520 20250 16570 20300
rect 16615 20250 16665 20300
rect 16715 20250 16765 20300
rect 16815 20250 16865 20300
rect 16915 20250 16965 20300
rect 17010 20250 17060 20300
rect 17105 20250 17155 20300
rect 17225 20250 17275 20300
rect 17320 20250 17370 20300
rect 17415 20250 17465 20300
rect 17515 20250 17565 20300
rect 17615 20250 17665 20300
rect 17715 20250 17765 20300
rect 17810 20250 17860 20300
rect 17905 20250 17955 20300
rect 14825 20160 14875 20210
rect 14920 20160 14970 20210
rect 15015 20160 15065 20210
rect 15115 20160 15165 20210
rect 15215 20160 15265 20210
rect 15315 20160 15365 20210
rect 15410 20160 15460 20210
rect 15505 20160 15555 20210
rect 15625 20160 15675 20210
rect 15720 20160 15770 20210
rect 15815 20160 15865 20210
rect 15915 20160 15965 20210
rect 16015 20160 16065 20210
rect 16115 20160 16165 20210
rect 16210 20160 16260 20210
rect 16305 20160 16355 20210
rect 16425 20160 16475 20210
rect 16520 20160 16570 20210
rect 16615 20160 16665 20210
rect 16715 20160 16765 20210
rect 16815 20160 16865 20210
rect 16915 20160 16965 20210
rect 17010 20160 17060 20210
rect 17105 20160 17155 20210
rect 17225 20160 17275 20210
rect 17320 20160 17370 20210
rect 17415 20160 17465 20210
rect 17515 20160 17565 20210
rect 17615 20160 17665 20210
rect 17715 20160 17765 20210
rect 17810 20160 17860 20210
rect 17905 20160 17955 20210
rect 14825 20040 14875 20090
rect 14920 20040 14970 20090
rect 15015 20040 15065 20090
rect 15115 20040 15165 20090
rect 15215 20040 15265 20090
rect 15315 20040 15365 20090
rect 15410 20040 15460 20090
rect 15505 20040 15555 20090
rect 15625 20040 15675 20090
rect 15720 20040 15770 20090
rect 15815 20040 15865 20090
rect 15915 20040 15965 20090
rect 16015 20040 16065 20090
rect 16115 20040 16165 20090
rect 16210 20040 16260 20090
rect 16305 20040 16355 20090
rect 16425 20040 16475 20090
rect 16520 20040 16570 20090
rect 16615 20040 16665 20090
rect 16715 20040 16765 20090
rect 16815 20040 16865 20090
rect 16915 20040 16965 20090
rect 17010 20040 17060 20090
rect 17105 20040 17155 20090
rect 17225 20040 17275 20090
rect 17320 20040 17370 20090
rect 17415 20040 17465 20090
rect 17515 20040 17565 20090
rect 17615 20040 17665 20090
rect 17715 20040 17765 20090
rect 17810 20040 17860 20090
rect 17905 20040 17955 20090
rect 14825 19950 14875 20000
rect 14920 19950 14970 20000
rect 15015 19950 15065 20000
rect 15115 19950 15165 20000
rect 15215 19950 15265 20000
rect 15315 19950 15365 20000
rect 15410 19950 15460 20000
rect 15505 19950 15555 20000
rect 15625 19950 15675 20000
rect 15720 19950 15770 20000
rect 15815 19950 15865 20000
rect 15915 19950 15965 20000
rect 16015 19950 16065 20000
rect 16115 19950 16165 20000
rect 16210 19950 16260 20000
rect 16305 19950 16355 20000
rect 16425 19950 16475 20000
rect 16520 19950 16570 20000
rect 16615 19950 16665 20000
rect 16715 19950 16765 20000
rect 16815 19950 16865 20000
rect 16915 19950 16965 20000
rect 17010 19950 17060 20000
rect 17105 19950 17155 20000
rect 17225 19950 17275 20000
rect 17320 19950 17370 20000
rect 17415 19950 17465 20000
rect 17515 19950 17565 20000
rect 17615 19950 17665 20000
rect 17715 19950 17765 20000
rect 17810 19950 17860 20000
rect 17905 19950 17955 20000
rect 14825 19850 14875 19900
rect 14920 19850 14970 19900
rect 15015 19850 15065 19900
rect 15115 19850 15165 19900
rect 15215 19850 15265 19900
rect 15315 19850 15365 19900
rect 15410 19850 15460 19900
rect 15505 19850 15555 19900
rect 15625 19850 15675 19900
rect 15720 19850 15770 19900
rect 15815 19850 15865 19900
rect 15915 19850 15965 19900
rect 16015 19850 16065 19900
rect 16115 19850 16165 19900
rect 16210 19850 16260 19900
rect 16305 19850 16355 19900
rect 16425 19850 16475 19900
rect 16520 19850 16570 19900
rect 16615 19850 16665 19900
rect 16715 19850 16765 19900
rect 16815 19850 16865 19900
rect 16915 19850 16965 19900
rect 17010 19850 17060 19900
rect 17105 19850 17155 19900
rect 17225 19850 17275 19900
rect 17320 19850 17370 19900
rect 17415 19850 17465 19900
rect 17515 19850 17565 19900
rect 17615 19850 17665 19900
rect 17715 19850 17765 19900
rect 17810 19850 17860 19900
rect 17905 19850 17955 19900
rect 14825 19760 14875 19810
rect 14920 19760 14970 19810
rect 15015 19760 15065 19810
rect 15115 19760 15165 19810
rect 15215 19760 15265 19810
rect 15315 19760 15365 19810
rect 15410 19760 15460 19810
rect 15505 19760 15555 19810
rect 15625 19760 15675 19810
rect 15720 19760 15770 19810
rect 15815 19760 15865 19810
rect 15915 19760 15965 19810
rect 16015 19760 16065 19810
rect 16115 19760 16165 19810
rect 16210 19760 16260 19810
rect 16305 19760 16355 19810
rect 16425 19760 16475 19810
rect 16520 19760 16570 19810
rect 16615 19760 16665 19810
rect 16715 19760 16765 19810
rect 16815 19760 16865 19810
rect 16915 19760 16965 19810
rect 17010 19760 17060 19810
rect 17105 19760 17155 19810
rect 17225 19760 17275 19810
rect 17320 19760 17370 19810
rect 17415 19760 17465 19810
rect 17515 19760 17565 19810
rect 17615 19760 17665 19810
rect 17715 19760 17765 19810
rect 17810 19760 17860 19810
rect 17905 19760 17955 19810
rect 14825 19640 14875 19690
rect 14920 19640 14970 19690
rect 15015 19640 15065 19690
rect 15115 19640 15165 19690
rect 15215 19640 15265 19690
rect 15315 19640 15365 19690
rect 15410 19640 15460 19690
rect 15505 19640 15555 19690
rect 15625 19640 15675 19690
rect 15720 19640 15770 19690
rect 15815 19640 15865 19690
rect 15915 19640 15965 19690
rect 16015 19640 16065 19690
rect 16115 19640 16165 19690
rect 16210 19640 16260 19690
rect 16305 19640 16355 19690
rect 16425 19640 16475 19690
rect 16520 19640 16570 19690
rect 16615 19640 16665 19690
rect 16715 19640 16765 19690
rect 16815 19640 16865 19690
rect 16915 19640 16965 19690
rect 17010 19640 17060 19690
rect 17105 19640 17155 19690
rect 17225 19640 17275 19690
rect 17320 19640 17370 19690
rect 17415 19640 17465 19690
rect 17515 19640 17565 19690
rect 17615 19640 17665 19690
rect 17715 19640 17765 19690
rect 17810 19640 17860 19690
rect 17905 19640 17955 19690
rect 14825 19550 14875 19600
rect 14920 19550 14970 19600
rect 15015 19550 15065 19600
rect 15115 19550 15165 19600
rect 15215 19550 15265 19600
rect 15315 19550 15365 19600
rect 15410 19550 15460 19600
rect 15505 19550 15555 19600
rect 15625 19550 15675 19600
rect 15720 19550 15770 19600
rect 15815 19550 15865 19600
rect 15915 19550 15965 19600
rect 16015 19550 16065 19600
rect 16115 19550 16165 19600
rect 16210 19550 16260 19600
rect 16305 19550 16355 19600
rect 16425 19550 16475 19600
rect 16520 19550 16570 19600
rect 16615 19550 16665 19600
rect 16715 19550 16765 19600
rect 16815 19550 16865 19600
rect 16915 19550 16965 19600
rect 17010 19550 17060 19600
rect 17105 19550 17155 19600
rect 17225 19550 17275 19600
rect 17320 19550 17370 19600
rect 17415 19550 17465 19600
rect 17515 19550 17565 19600
rect 17615 19550 17665 19600
rect 17715 19550 17765 19600
rect 17810 19550 17860 19600
rect 17905 19550 17955 19600
rect 14825 19450 14875 19500
rect 14920 19450 14970 19500
rect 15015 19450 15065 19500
rect 15115 19450 15165 19500
rect 15215 19450 15265 19500
rect 15315 19450 15365 19500
rect 15410 19450 15460 19500
rect 15505 19450 15555 19500
rect 15625 19450 15675 19500
rect 15720 19450 15770 19500
rect 15815 19450 15865 19500
rect 15915 19450 15965 19500
rect 16015 19450 16065 19500
rect 16115 19450 16165 19500
rect 16210 19450 16260 19500
rect 16305 19450 16355 19500
rect 16425 19450 16475 19500
rect 16520 19450 16570 19500
rect 16615 19450 16665 19500
rect 16715 19450 16765 19500
rect 16815 19450 16865 19500
rect 16915 19450 16965 19500
rect 17010 19450 17060 19500
rect 17105 19450 17155 19500
rect 17225 19450 17275 19500
rect 17320 19450 17370 19500
rect 17415 19450 17465 19500
rect 17515 19450 17565 19500
rect 17615 19450 17665 19500
rect 17715 19450 17765 19500
rect 17810 19450 17860 19500
rect 17905 19450 17955 19500
rect 14825 19360 14875 19410
rect 14920 19360 14970 19410
rect 15015 19360 15065 19410
rect 15115 19360 15165 19410
rect 15215 19360 15265 19410
rect 15315 19360 15365 19410
rect 15410 19360 15460 19410
rect 15505 19360 15555 19410
rect 15625 19360 15675 19410
rect 15720 19360 15770 19410
rect 15815 19360 15865 19410
rect 15915 19360 15965 19410
rect 16015 19360 16065 19410
rect 16115 19360 16165 19410
rect 16210 19360 16260 19410
rect 16305 19360 16355 19410
rect 16425 19360 16475 19410
rect 16520 19360 16570 19410
rect 16615 19360 16665 19410
rect 16715 19360 16765 19410
rect 16815 19360 16865 19410
rect 16915 19360 16965 19410
rect 17010 19360 17060 19410
rect 17105 19360 17155 19410
rect 17225 19360 17275 19410
rect 17320 19360 17370 19410
rect 17415 19360 17465 19410
rect 17515 19360 17565 19410
rect 17615 19360 17665 19410
rect 17715 19360 17765 19410
rect 17810 19360 17860 19410
rect 17905 19360 17955 19410
rect 14825 19240 14875 19290
rect 14920 19240 14970 19290
rect 15015 19240 15065 19290
rect 15115 19240 15165 19290
rect 15215 19240 15265 19290
rect 15315 19240 15365 19290
rect 15410 19240 15460 19290
rect 15505 19240 15555 19290
rect 15625 19240 15675 19290
rect 15720 19240 15770 19290
rect 15815 19240 15865 19290
rect 15915 19240 15965 19290
rect 16015 19240 16065 19290
rect 16115 19240 16165 19290
rect 16210 19240 16260 19290
rect 16305 19240 16355 19290
rect 16425 19240 16475 19290
rect 16520 19240 16570 19290
rect 16615 19240 16665 19290
rect 16715 19240 16765 19290
rect 16815 19240 16865 19290
rect 16915 19240 16965 19290
rect 17010 19240 17060 19290
rect 17105 19240 17155 19290
rect 17225 19240 17275 19290
rect 17320 19240 17370 19290
rect 17415 19240 17465 19290
rect 17515 19240 17565 19290
rect 17615 19240 17665 19290
rect 17715 19240 17765 19290
rect 17810 19240 17860 19290
rect 17905 19240 17955 19290
rect 14825 19150 14875 19200
rect 14920 19150 14970 19200
rect 15015 19150 15065 19200
rect 15115 19150 15165 19200
rect 15215 19150 15265 19200
rect 15315 19150 15365 19200
rect 15410 19150 15460 19200
rect 15505 19150 15555 19200
rect 15625 19150 15675 19200
rect 15720 19150 15770 19200
rect 15815 19150 15865 19200
rect 15915 19150 15965 19200
rect 16015 19150 16065 19200
rect 16115 19150 16165 19200
rect 16210 19150 16260 19200
rect 16305 19150 16355 19200
rect 16425 19150 16475 19200
rect 16520 19150 16570 19200
rect 16615 19150 16665 19200
rect 16715 19150 16765 19200
rect 16815 19150 16865 19200
rect 16915 19150 16965 19200
rect 17010 19150 17060 19200
rect 17105 19150 17155 19200
rect 17225 19150 17275 19200
rect 17320 19150 17370 19200
rect 17415 19150 17465 19200
rect 17515 19150 17565 19200
rect 17615 19150 17665 19200
rect 17715 19150 17765 19200
rect 17810 19150 17860 19200
rect 17905 19150 17955 19200
rect 14825 19050 14875 19100
rect 14920 19050 14970 19100
rect 15015 19050 15065 19100
rect 15115 19050 15165 19100
rect 15215 19050 15265 19100
rect 15315 19050 15365 19100
rect 15410 19050 15460 19100
rect 15505 19050 15555 19100
rect 15625 19050 15675 19100
rect 15720 19050 15770 19100
rect 15815 19050 15865 19100
rect 15915 19050 15965 19100
rect 16015 19050 16065 19100
rect 16115 19050 16165 19100
rect 16210 19050 16260 19100
rect 16305 19050 16355 19100
rect 16425 19050 16475 19100
rect 16520 19050 16570 19100
rect 16615 19050 16665 19100
rect 16715 19050 16765 19100
rect 16815 19050 16865 19100
rect 16915 19050 16965 19100
rect 17010 19050 17060 19100
rect 17105 19050 17155 19100
rect 17225 19050 17275 19100
rect 17320 19050 17370 19100
rect 17415 19050 17465 19100
rect 17515 19050 17565 19100
rect 17615 19050 17665 19100
rect 17715 19050 17765 19100
rect 17810 19050 17860 19100
rect 17905 19050 17955 19100
rect 14825 18960 14875 19010
rect 14920 18960 14970 19010
rect 15015 18960 15065 19010
rect 15115 18960 15165 19010
rect 15215 18960 15265 19010
rect 15315 18960 15365 19010
rect 15410 18960 15460 19010
rect 15505 18960 15555 19010
rect 15625 18960 15675 19010
rect 15720 18960 15770 19010
rect 15815 18960 15865 19010
rect 15915 18960 15965 19010
rect 16015 18960 16065 19010
rect 16115 18960 16165 19010
rect 16210 18960 16260 19010
rect 16305 18960 16355 19010
rect 16425 18960 16475 19010
rect 16520 18960 16570 19010
rect 16615 18960 16665 19010
rect 16715 18960 16765 19010
rect 16815 18960 16865 19010
rect 16915 18960 16965 19010
rect 17010 18960 17060 19010
rect 17105 18960 17155 19010
rect 17225 18960 17275 19010
rect 17320 18960 17370 19010
rect 17415 18960 17465 19010
rect 17515 18960 17565 19010
rect 17615 18960 17665 19010
rect 17715 18960 17765 19010
rect 17810 18960 17860 19010
rect 17905 18960 17955 19010
rect 14825 18840 14875 18890
rect 14920 18840 14970 18890
rect 15015 18840 15065 18890
rect 15115 18840 15165 18890
rect 15215 18840 15265 18890
rect 15315 18840 15365 18890
rect 15410 18840 15460 18890
rect 15505 18840 15555 18890
rect 15625 18840 15675 18890
rect 15720 18840 15770 18890
rect 15815 18840 15865 18890
rect 15915 18840 15965 18890
rect 16015 18840 16065 18890
rect 16115 18840 16165 18890
rect 16210 18840 16260 18890
rect 16305 18840 16355 18890
rect 16425 18840 16475 18890
rect 16520 18840 16570 18890
rect 16615 18840 16665 18890
rect 16715 18840 16765 18890
rect 16815 18840 16865 18890
rect 16915 18840 16965 18890
rect 17010 18840 17060 18890
rect 17105 18840 17155 18890
rect 17225 18840 17275 18890
rect 17320 18840 17370 18890
rect 17415 18840 17465 18890
rect 17515 18840 17565 18890
rect 17615 18840 17665 18890
rect 17715 18840 17765 18890
rect 17810 18840 17860 18890
rect 17905 18840 17955 18890
rect 14825 18750 14875 18800
rect 14920 18750 14970 18800
rect 15015 18750 15065 18800
rect 15115 18750 15165 18800
rect 15215 18750 15265 18800
rect 15315 18750 15365 18800
rect 15410 18750 15460 18800
rect 15505 18750 15555 18800
rect 15625 18750 15675 18800
rect 15720 18750 15770 18800
rect 15815 18750 15865 18800
rect 15915 18750 15965 18800
rect 16015 18750 16065 18800
rect 16115 18750 16165 18800
rect 16210 18750 16260 18800
rect 16305 18750 16355 18800
rect 16425 18750 16475 18800
rect 16520 18750 16570 18800
rect 16615 18750 16665 18800
rect 16715 18750 16765 18800
rect 16815 18750 16865 18800
rect 16915 18750 16965 18800
rect 17010 18750 17060 18800
rect 17105 18750 17155 18800
rect 17225 18750 17275 18800
rect 17320 18750 17370 18800
rect 17415 18750 17465 18800
rect 17515 18750 17565 18800
rect 17615 18750 17665 18800
rect 17715 18750 17765 18800
rect 17810 18750 17860 18800
rect 17905 18750 17955 18800
rect 14825 18650 14875 18700
rect 14920 18650 14970 18700
rect 15015 18650 15065 18700
rect 15115 18650 15165 18700
rect 15215 18650 15265 18700
rect 15315 18650 15365 18700
rect 15410 18650 15460 18700
rect 15505 18650 15555 18700
rect 15625 18650 15675 18700
rect 15720 18650 15770 18700
rect 15815 18650 15865 18700
rect 15915 18650 15965 18700
rect 16015 18650 16065 18700
rect 16115 18650 16165 18700
rect 16210 18650 16260 18700
rect 16305 18650 16355 18700
rect 16425 18650 16475 18700
rect 16520 18650 16570 18700
rect 16615 18650 16665 18700
rect 16715 18650 16765 18700
rect 16815 18650 16865 18700
rect 16915 18650 16965 18700
rect 17010 18650 17060 18700
rect 17105 18650 17155 18700
rect 17225 18650 17275 18700
rect 17320 18650 17370 18700
rect 17415 18650 17465 18700
rect 17515 18650 17565 18700
rect 17615 18650 17665 18700
rect 17715 18650 17765 18700
rect 17810 18650 17860 18700
rect 17905 18650 17955 18700
rect 14825 18560 14875 18610
rect 14920 18560 14970 18610
rect 15015 18560 15065 18610
rect 15115 18560 15165 18610
rect 15215 18560 15265 18610
rect 15315 18560 15365 18610
rect 15410 18560 15460 18610
rect 15505 18560 15555 18610
rect 15625 18560 15675 18610
rect 15720 18560 15770 18610
rect 15815 18560 15865 18610
rect 15915 18560 15965 18610
rect 16015 18560 16065 18610
rect 16115 18560 16165 18610
rect 16210 18560 16260 18610
rect 16305 18560 16355 18610
rect 16425 18560 16475 18610
rect 16520 18560 16570 18610
rect 16615 18560 16665 18610
rect 16715 18560 16765 18610
rect 16815 18560 16865 18610
rect 16915 18560 16965 18610
rect 17010 18560 17060 18610
rect 17105 18560 17155 18610
rect 17225 18560 17275 18610
rect 17320 18560 17370 18610
rect 17415 18560 17465 18610
rect 17515 18560 17565 18610
rect 17615 18560 17665 18610
rect 17715 18560 17765 18610
rect 17810 18560 17860 18610
rect 17905 18560 17955 18610
rect 14825 18440 14875 18490
rect 14920 18440 14970 18490
rect 15015 18440 15065 18490
rect 15115 18440 15165 18490
rect 15215 18440 15265 18490
rect 15315 18440 15365 18490
rect 15410 18440 15460 18490
rect 15505 18440 15555 18490
rect 15625 18440 15675 18490
rect 15720 18440 15770 18490
rect 15815 18440 15865 18490
rect 15915 18440 15965 18490
rect 16015 18440 16065 18490
rect 16115 18440 16165 18490
rect 16210 18440 16260 18490
rect 16305 18440 16355 18490
rect 16425 18440 16475 18490
rect 16520 18440 16570 18490
rect 16615 18440 16665 18490
rect 16715 18440 16765 18490
rect 16815 18440 16865 18490
rect 16915 18440 16965 18490
rect 17010 18440 17060 18490
rect 17105 18440 17155 18490
rect 17225 18440 17275 18490
rect 17320 18440 17370 18490
rect 17415 18440 17465 18490
rect 17515 18440 17565 18490
rect 17615 18440 17665 18490
rect 17715 18440 17765 18490
rect 17810 18440 17860 18490
rect 17905 18440 17955 18490
rect 14825 18350 14875 18400
rect 14920 18350 14970 18400
rect 15015 18350 15065 18400
rect 15115 18350 15165 18400
rect 15215 18350 15265 18400
rect 15315 18350 15365 18400
rect 15410 18350 15460 18400
rect 15505 18350 15555 18400
rect 15625 18350 15675 18400
rect 15720 18350 15770 18400
rect 15815 18350 15865 18400
rect 15915 18350 15965 18400
rect 16015 18350 16065 18400
rect 16115 18350 16165 18400
rect 16210 18350 16260 18400
rect 16305 18350 16355 18400
rect 16425 18350 16475 18400
rect 16520 18350 16570 18400
rect 16615 18350 16665 18400
rect 16715 18350 16765 18400
rect 16815 18350 16865 18400
rect 16915 18350 16965 18400
rect 17010 18350 17060 18400
rect 17105 18350 17155 18400
rect 17225 18350 17275 18400
rect 17320 18350 17370 18400
rect 17415 18350 17465 18400
rect 17515 18350 17565 18400
rect 17615 18350 17665 18400
rect 17715 18350 17765 18400
rect 17810 18350 17860 18400
rect 17905 18350 17955 18400
rect 14825 18250 14875 18300
rect 14920 18250 14970 18300
rect 15015 18250 15065 18300
rect 15115 18250 15165 18300
rect 15215 18250 15265 18300
rect 15315 18250 15365 18300
rect 15410 18250 15460 18300
rect 15505 18250 15555 18300
rect 15625 18250 15675 18300
rect 15720 18250 15770 18300
rect 15815 18250 15865 18300
rect 15915 18250 15965 18300
rect 16015 18250 16065 18300
rect 16115 18250 16165 18300
rect 16210 18250 16260 18300
rect 16305 18250 16355 18300
rect 16425 18250 16475 18300
rect 16520 18250 16570 18300
rect 16615 18250 16665 18300
rect 16715 18250 16765 18300
rect 16815 18250 16865 18300
rect 16915 18250 16965 18300
rect 17010 18250 17060 18300
rect 17105 18250 17155 18300
rect 17225 18250 17275 18300
rect 17320 18250 17370 18300
rect 17415 18250 17465 18300
rect 17515 18250 17565 18300
rect 17615 18250 17665 18300
rect 17715 18250 17765 18300
rect 17810 18250 17860 18300
rect 17905 18250 17955 18300
rect 14825 18160 14875 18210
rect 14920 18160 14970 18210
rect 15015 18160 15065 18210
rect 15115 18160 15165 18210
rect 15215 18160 15265 18210
rect 15315 18160 15365 18210
rect 15410 18160 15460 18210
rect 15505 18160 15555 18210
rect 15625 18160 15675 18210
rect 15720 18160 15770 18210
rect 15815 18160 15865 18210
rect 15915 18160 15965 18210
rect 16015 18160 16065 18210
rect 16115 18160 16165 18210
rect 16210 18160 16260 18210
rect 16305 18160 16355 18210
rect 16425 18160 16475 18210
rect 16520 18160 16570 18210
rect 16615 18160 16665 18210
rect 16715 18160 16765 18210
rect 16815 18160 16865 18210
rect 16915 18160 16965 18210
rect 17010 18160 17060 18210
rect 17105 18160 17155 18210
rect 17225 18160 17275 18210
rect 17320 18160 17370 18210
rect 17415 18160 17465 18210
rect 17515 18160 17565 18210
rect 17615 18160 17665 18210
rect 17715 18160 17765 18210
rect 17810 18160 17860 18210
rect 17905 18160 17955 18210
rect 14825 18040 14875 18090
rect 14920 18040 14970 18090
rect 15015 18040 15065 18090
rect 15115 18040 15165 18090
rect 15215 18040 15265 18090
rect 15315 18040 15365 18090
rect 15410 18040 15460 18090
rect 15505 18040 15555 18090
rect 15625 18040 15675 18090
rect 15720 18040 15770 18090
rect 15815 18040 15865 18090
rect 15915 18040 15965 18090
rect 16015 18040 16065 18090
rect 16115 18040 16165 18090
rect 16210 18040 16260 18090
rect 16305 18040 16355 18090
rect 16425 18040 16475 18090
rect 16520 18040 16570 18090
rect 16615 18040 16665 18090
rect 16715 18040 16765 18090
rect 16815 18040 16865 18090
rect 16915 18040 16965 18090
rect 17010 18040 17060 18090
rect 17105 18040 17155 18090
rect 17225 18040 17275 18090
rect 17320 18040 17370 18090
rect 17415 18040 17465 18090
rect 17515 18040 17565 18090
rect 17615 18040 17665 18090
rect 17715 18040 17765 18090
rect 17810 18040 17860 18090
rect 17905 18040 17955 18090
rect 14825 17950 14875 18000
rect 14920 17950 14970 18000
rect 15015 17950 15065 18000
rect 15115 17950 15165 18000
rect 15215 17950 15265 18000
rect 15315 17950 15365 18000
rect 15410 17950 15460 18000
rect 15505 17950 15555 18000
rect 15625 17950 15675 18000
rect 15720 17950 15770 18000
rect 15815 17950 15865 18000
rect 15915 17950 15965 18000
rect 16015 17950 16065 18000
rect 16115 17950 16165 18000
rect 16210 17950 16260 18000
rect 16305 17950 16355 18000
rect 16425 17950 16475 18000
rect 16520 17950 16570 18000
rect 16615 17950 16665 18000
rect 16715 17950 16765 18000
rect 16815 17950 16865 18000
rect 16915 17950 16965 18000
rect 17010 17950 17060 18000
rect 17105 17950 17155 18000
rect 17225 17950 17275 18000
rect 17320 17950 17370 18000
rect 17415 17950 17465 18000
rect 17515 17950 17565 18000
rect 17615 17950 17665 18000
rect 17715 17950 17765 18000
rect 17810 17950 17860 18000
rect 17905 17950 17955 18000
rect 14825 17850 14875 17900
rect 14920 17850 14970 17900
rect 15015 17850 15065 17900
rect 15115 17850 15165 17900
rect 15215 17850 15265 17900
rect 15315 17850 15365 17900
rect 15410 17850 15460 17900
rect 15505 17850 15555 17900
rect 15625 17850 15675 17900
rect 15720 17850 15770 17900
rect 15815 17850 15865 17900
rect 15915 17850 15965 17900
rect 16015 17850 16065 17900
rect 16115 17850 16165 17900
rect 16210 17850 16260 17900
rect 16305 17850 16355 17900
rect 16425 17850 16475 17900
rect 16520 17850 16570 17900
rect 16615 17850 16665 17900
rect 16715 17850 16765 17900
rect 16815 17850 16865 17900
rect 16915 17850 16965 17900
rect 17010 17850 17060 17900
rect 17105 17850 17155 17900
rect 17225 17850 17275 17900
rect 17320 17850 17370 17900
rect 17415 17850 17465 17900
rect 17515 17850 17565 17900
rect 17615 17850 17665 17900
rect 17715 17850 17765 17900
rect 17810 17850 17860 17900
rect 17905 17850 17955 17900
rect 14825 17760 14875 17810
rect 14920 17760 14970 17810
rect 15015 17760 15065 17810
rect 15115 17760 15165 17810
rect 15215 17760 15265 17810
rect 15315 17760 15365 17810
rect 15410 17760 15460 17810
rect 15505 17760 15555 17810
rect 15625 17760 15675 17810
rect 15720 17760 15770 17810
rect 15815 17760 15865 17810
rect 15915 17760 15965 17810
rect 16015 17760 16065 17810
rect 16115 17760 16165 17810
rect 16210 17760 16260 17810
rect 16305 17760 16355 17810
rect 16425 17760 16475 17810
rect 16520 17760 16570 17810
rect 16615 17760 16665 17810
rect 16715 17760 16765 17810
rect 16815 17760 16865 17810
rect 16915 17760 16965 17810
rect 17010 17760 17060 17810
rect 17105 17760 17155 17810
rect 17225 17760 17275 17810
rect 17320 17760 17370 17810
rect 17415 17760 17465 17810
rect 17515 17760 17565 17810
rect 17615 17760 17665 17810
rect 17715 17760 17765 17810
rect 17810 17760 17860 17810
rect 17905 17760 17955 17810
rect -4805 9565 -4755 9615
rect -4710 9565 -4660 9615
rect -4615 9565 -4565 9615
rect -4515 9565 -4465 9615
rect -4415 9565 -4365 9615
rect -4315 9565 -4265 9615
rect -4220 9565 -4170 9615
rect -4125 9565 -4075 9615
rect -4005 9565 -3955 9615
rect -3910 9565 -3860 9615
rect -3815 9565 -3765 9615
rect -3715 9565 -3665 9615
rect -3615 9565 -3565 9615
rect -3515 9565 -3465 9615
rect -3420 9565 -3370 9615
rect -3325 9565 -3275 9615
rect -3205 9565 -3155 9615
rect -3110 9565 -3060 9615
rect -3015 9565 -2965 9615
rect -2915 9565 -2865 9615
rect -2815 9565 -2765 9615
rect -2715 9565 -2665 9615
rect -2620 9565 -2570 9615
rect -2525 9565 -2475 9615
rect -2405 9565 -2355 9615
rect -2310 9565 -2260 9615
rect -2215 9565 -2165 9615
rect -2115 9565 -2065 9615
rect -2015 9565 -1965 9615
rect -1915 9565 -1865 9615
rect -1820 9565 -1770 9615
rect -1725 9565 -1675 9615
rect -4805 9475 -4755 9525
rect -4710 9475 -4660 9525
rect -4615 9475 -4565 9525
rect -4515 9475 -4465 9525
rect -4415 9475 -4365 9525
rect -4315 9475 -4265 9525
rect -4220 9475 -4170 9525
rect -4125 9475 -4075 9525
rect -4005 9475 -3955 9525
rect -3910 9475 -3860 9525
rect -3815 9475 -3765 9525
rect -3715 9475 -3665 9525
rect -3615 9475 -3565 9525
rect -3515 9475 -3465 9525
rect -3420 9475 -3370 9525
rect -3325 9475 -3275 9525
rect -3205 9475 -3155 9525
rect -3110 9475 -3060 9525
rect -3015 9475 -2965 9525
rect -2915 9475 -2865 9525
rect -2815 9475 -2765 9525
rect -2715 9475 -2665 9525
rect -2620 9475 -2570 9525
rect -2525 9475 -2475 9525
rect -2405 9475 -2355 9525
rect -2310 9475 -2260 9525
rect -2215 9475 -2165 9525
rect -2115 9475 -2065 9525
rect -2015 9475 -1965 9525
rect -1915 9475 -1865 9525
rect -1820 9475 -1770 9525
rect -1725 9475 -1675 9525
rect -4805 9375 -4755 9425
rect -4710 9375 -4660 9425
rect -4615 9375 -4565 9425
rect -4515 9375 -4465 9425
rect -4415 9375 -4365 9425
rect -4315 9375 -4265 9425
rect -4220 9375 -4170 9425
rect -4125 9375 -4075 9425
rect -4005 9375 -3955 9425
rect -3910 9375 -3860 9425
rect -3815 9375 -3765 9425
rect -3715 9375 -3665 9425
rect -3615 9375 -3565 9425
rect -3515 9375 -3465 9425
rect -3420 9375 -3370 9425
rect -3325 9375 -3275 9425
rect -3205 9375 -3155 9425
rect -3110 9375 -3060 9425
rect -3015 9375 -2965 9425
rect -2915 9375 -2865 9425
rect -2815 9375 -2765 9425
rect -2715 9375 -2665 9425
rect -2620 9375 -2570 9425
rect -2525 9375 -2475 9425
rect -2405 9375 -2355 9425
rect -2310 9375 -2260 9425
rect -2215 9375 -2165 9425
rect -2115 9375 -2065 9425
rect -2015 9375 -1965 9425
rect -1915 9375 -1865 9425
rect -1820 9375 -1770 9425
rect -1725 9375 -1675 9425
rect -4805 9285 -4755 9335
rect -4710 9285 -4660 9335
rect -4615 9285 -4565 9335
rect -4515 9285 -4465 9335
rect -4415 9285 -4365 9335
rect -4315 9285 -4265 9335
rect -4220 9285 -4170 9335
rect -4125 9285 -4075 9335
rect -4005 9285 -3955 9335
rect -3910 9285 -3860 9335
rect -3815 9285 -3765 9335
rect -3715 9285 -3665 9335
rect -3615 9285 -3565 9335
rect -3515 9285 -3465 9335
rect -3420 9285 -3370 9335
rect -3325 9285 -3275 9335
rect -3205 9285 -3155 9335
rect -3110 9285 -3060 9335
rect -3015 9285 -2965 9335
rect -2915 9285 -2865 9335
rect -2815 9285 -2765 9335
rect -2715 9285 -2665 9335
rect -2620 9285 -2570 9335
rect -2525 9285 -2475 9335
rect -2405 9285 -2355 9335
rect -2310 9285 -2260 9335
rect -2215 9285 -2165 9335
rect -2115 9285 -2065 9335
rect -2015 9285 -1965 9335
rect -1915 9285 -1865 9335
rect -1820 9285 -1770 9335
rect -1725 9285 -1675 9335
rect -4805 9165 -4755 9215
rect -4710 9165 -4660 9215
rect -4615 9165 -4565 9215
rect -4515 9165 -4465 9215
rect -4415 9165 -4365 9215
rect -4315 9165 -4265 9215
rect -4220 9165 -4170 9215
rect -4125 9165 -4075 9215
rect -4005 9165 -3955 9215
rect -3910 9165 -3860 9215
rect -3815 9165 -3765 9215
rect -3715 9165 -3665 9215
rect -3615 9165 -3565 9215
rect -3515 9165 -3465 9215
rect -3420 9165 -3370 9215
rect -3325 9165 -3275 9215
rect -3205 9165 -3155 9215
rect -3110 9165 -3060 9215
rect -3015 9165 -2965 9215
rect -2915 9165 -2865 9215
rect -2815 9165 -2765 9215
rect -2715 9165 -2665 9215
rect -2620 9165 -2570 9215
rect -2525 9165 -2475 9215
rect -2405 9165 -2355 9215
rect -2310 9165 -2260 9215
rect -2215 9165 -2165 9215
rect -2115 9165 -2065 9215
rect -2015 9165 -1965 9215
rect -1915 9165 -1865 9215
rect -1820 9165 -1770 9215
rect -1725 9165 -1675 9215
rect -4805 9075 -4755 9125
rect -4710 9075 -4660 9125
rect -4615 9075 -4565 9125
rect -4515 9075 -4465 9125
rect -4415 9075 -4365 9125
rect -4315 9075 -4265 9125
rect -4220 9075 -4170 9125
rect -4125 9075 -4075 9125
rect -4005 9075 -3955 9125
rect -3910 9075 -3860 9125
rect -3815 9075 -3765 9125
rect -3715 9075 -3665 9125
rect -3615 9075 -3565 9125
rect -3515 9075 -3465 9125
rect -3420 9075 -3370 9125
rect -3325 9075 -3275 9125
rect -3205 9075 -3155 9125
rect -3110 9075 -3060 9125
rect -3015 9075 -2965 9125
rect -2915 9075 -2865 9125
rect -2815 9075 -2765 9125
rect -2715 9075 -2665 9125
rect -2620 9075 -2570 9125
rect -2525 9075 -2475 9125
rect -2405 9075 -2355 9125
rect -2310 9075 -2260 9125
rect -2215 9075 -2165 9125
rect -2115 9075 -2065 9125
rect -2015 9075 -1965 9125
rect -1915 9075 -1865 9125
rect -1820 9075 -1770 9125
rect -1725 9075 -1675 9125
rect -4805 8975 -4755 9025
rect -4710 8975 -4660 9025
rect -4615 8975 -4565 9025
rect -4515 8975 -4465 9025
rect -4415 8975 -4365 9025
rect -4315 8975 -4265 9025
rect -4220 8975 -4170 9025
rect -4125 8975 -4075 9025
rect -4005 8975 -3955 9025
rect -3910 8975 -3860 9025
rect -3815 8975 -3765 9025
rect -3715 8975 -3665 9025
rect -3615 8975 -3565 9025
rect -3515 8975 -3465 9025
rect -3420 8975 -3370 9025
rect -3325 8975 -3275 9025
rect -3205 8975 -3155 9025
rect -3110 8975 -3060 9025
rect -3015 8975 -2965 9025
rect -2915 8975 -2865 9025
rect -2815 8975 -2765 9025
rect -2715 8975 -2665 9025
rect -2620 8975 -2570 9025
rect -2525 8975 -2475 9025
rect -2405 8975 -2355 9025
rect -2310 8975 -2260 9025
rect -2215 8975 -2165 9025
rect -2115 8975 -2065 9025
rect -2015 8975 -1965 9025
rect -1915 8975 -1865 9025
rect -1820 8975 -1770 9025
rect -1725 8975 -1675 9025
rect -4805 8885 -4755 8935
rect -4710 8885 -4660 8935
rect -4615 8885 -4565 8935
rect -4515 8885 -4465 8935
rect -4415 8885 -4365 8935
rect -4315 8885 -4265 8935
rect -4220 8885 -4170 8935
rect -4125 8885 -4075 8935
rect -4005 8885 -3955 8935
rect -3910 8885 -3860 8935
rect -3815 8885 -3765 8935
rect -3715 8885 -3665 8935
rect -3615 8885 -3565 8935
rect -3515 8885 -3465 8935
rect -3420 8885 -3370 8935
rect -3325 8885 -3275 8935
rect -3205 8885 -3155 8935
rect -3110 8885 -3060 8935
rect -3015 8885 -2965 8935
rect -2915 8885 -2865 8935
rect -2815 8885 -2765 8935
rect -2715 8885 -2665 8935
rect -2620 8885 -2570 8935
rect -2525 8885 -2475 8935
rect -2405 8885 -2355 8935
rect -2310 8885 -2260 8935
rect -2215 8885 -2165 8935
rect -2115 8885 -2065 8935
rect -2015 8885 -1965 8935
rect -1915 8885 -1865 8935
rect -1820 8885 -1770 8935
rect -1725 8885 -1675 8935
rect -4805 8765 -4755 8815
rect -4710 8765 -4660 8815
rect -4615 8765 -4565 8815
rect -4515 8765 -4465 8815
rect -4415 8765 -4365 8815
rect -4315 8765 -4265 8815
rect -4220 8765 -4170 8815
rect -4125 8765 -4075 8815
rect -4005 8765 -3955 8815
rect -3910 8765 -3860 8815
rect -3815 8765 -3765 8815
rect -3715 8765 -3665 8815
rect -3615 8765 -3565 8815
rect -3515 8765 -3465 8815
rect -3420 8765 -3370 8815
rect -3325 8765 -3275 8815
rect -3205 8765 -3155 8815
rect -3110 8765 -3060 8815
rect -3015 8765 -2965 8815
rect -2915 8765 -2865 8815
rect -2815 8765 -2765 8815
rect -2715 8765 -2665 8815
rect -2620 8765 -2570 8815
rect -2525 8765 -2475 8815
rect -2405 8765 -2355 8815
rect -2310 8765 -2260 8815
rect -2215 8765 -2165 8815
rect -2115 8765 -2065 8815
rect -2015 8765 -1965 8815
rect -1915 8765 -1865 8815
rect -1820 8765 -1770 8815
rect -1725 8765 -1675 8815
rect -4805 8675 -4755 8725
rect -4710 8675 -4660 8725
rect -4615 8675 -4565 8725
rect -4515 8675 -4465 8725
rect -4415 8675 -4365 8725
rect -4315 8675 -4265 8725
rect -4220 8675 -4170 8725
rect -4125 8675 -4075 8725
rect -4005 8675 -3955 8725
rect -3910 8675 -3860 8725
rect -3815 8675 -3765 8725
rect -3715 8675 -3665 8725
rect -3615 8675 -3565 8725
rect -3515 8675 -3465 8725
rect -3420 8675 -3370 8725
rect -3325 8675 -3275 8725
rect -3205 8675 -3155 8725
rect -3110 8675 -3060 8725
rect -3015 8675 -2965 8725
rect -2915 8675 -2865 8725
rect -2815 8675 -2765 8725
rect -2715 8675 -2665 8725
rect -2620 8675 -2570 8725
rect -2525 8675 -2475 8725
rect -2405 8675 -2355 8725
rect -2310 8675 -2260 8725
rect -2215 8675 -2165 8725
rect -2115 8675 -2065 8725
rect -2015 8675 -1965 8725
rect -1915 8675 -1865 8725
rect -1820 8675 -1770 8725
rect -1725 8675 -1675 8725
rect -4805 8575 -4755 8625
rect -4710 8575 -4660 8625
rect -4615 8575 -4565 8625
rect -4515 8575 -4465 8625
rect -4415 8575 -4365 8625
rect -4315 8575 -4265 8625
rect -4220 8575 -4170 8625
rect -4125 8575 -4075 8625
rect -4005 8575 -3955 8625
rect -3910 8575 -3860 8625
rect -3815 8575 -3765 8625
rect -3715 8575 -3665 8625
rect -3615 8575 -3565 8625
rect -3515 8575 -3465 8625
rect -3420 8575 -3370 8625
rect -3325 8575 -3275 8625
rect -3205 8575 -3155 8625
rect -3110 8575 -3060 8625
rect -3015 8575 -2965 8625
rect -2915 8575 -2865 8625
rect -2815 8575 -2765 8625
rect -2715 8575 -2665 8625
rect -2620 8575 -2570 8625
rect -2525 8575 -2475 8625
rect -2405 8575 -2355 8625
rect -2310 8575 -2260 8625
rect -2215 8575 -2165 8625
rect -2115 8575 -2065 8625
rect -2015 8575 -1965 8625
rect -1915 8575 -1865 8625
rect -1820 8575 -1770 8625
rect -1725 8575 -1675 8625
rect -4805 8485 -4755 8535
rect -4710 8485 -4660 8535
rect -4615 8485 -4565 8535
rect -4515 8485 -4465 8535
rect -4415 8485 -4365 8535
rect -4315 8485 -4265 8535
rect -4220 8485 -4170 8535
rect -4125 8485 -4075 8535
rect -4005 8485 -3955 8535
rect -3910 8485 -3860 8535
rect -3815 8485 -3765 8535
rect -3715 8485 -3665 8535
rect -3615 8485 -3565 8535
rect -3515 8485 -3465 8535
rect -3420 8485 -3370 8535
rect -3325 8485 -3275 8535
rect -3205 8485 -3155 8535
rect -3110 8485 -3060 8535
rect -3015 8485 -2965 8535
rect -2915 8485 -2865 8535
rect -2815 8485 -2765 8535
rect -2715 8485 -2665 8535
rect -2620 8485 -2570 8535
rect -2525 8485 -2475 8535
rect -2405 8485 -2355 8535
rect -2310 8485 -2260 8535
rect -2215 8485 -2165 8535
rect -2115 8485 -2065 8535
rect -2015 8485 -1965 8535
rect -1915 8485 -1865 8535
rect -1820 8485 -1770 8535
rect -1725 8485 -1675 8535
rect -4805 8365 -4755 8415
rect -4710 8365 -4660 8415
rect -4615 8365 -4565 8415
rect -4515 8365 -4465 8415
rect -4415 8365 -4365 8415
rect -4315 8365 -4265 8415
rect -4220 8365 -4170 8415
rect -4125 8365 -4075 8415
rect -4005 8365 -3955 8415
rect -3910 8365 -3860 8415
rect -3815 8365 -3765 8415
rect -3715 8365 -3665 8415
rect -3615 8365 -3565 8415
rect -3515 8365 -3465 8415
rect -3420 8365 -3370 8415
rect -3325 8365 -3275 8415
rect -3205 8365 -3155 8415
rect -3110 8365 -3060 8415
rect -3015 8365 -2965 8415
rect -2915 8365 -2865 8415
rect -2815 8365 -2765 8415
rect -2715 8365 -2665 8415
rect -2620 8365 -2570 8415
rect -2525 8365 -2475 8415
rect -2405 8365 -2355 8415
rect -2310 8365 -2260 8415
rect -2215 8365 -2165 8415
rect -2115 8365 -2065 8415
rect -2015 8365 -1965 8415
rect -1915 8365 -1865 8415
rect -1820 8365 -1770 8415
rect -1725 8365 -1675 8415
rect -4805 8275 -4755 8325
rect -4710 8275 -4660 8325
rect -4615 8275 -4565 8325
rect -4515 8275 -4465 8325
rect -4415 8275 -4365 8325
rect -4315 8275 -4265 8325
rect -4220 8275 -4170 8325
rect -4125 8275 -4075 8325
rect -4005 8275 -3955 8325
rect -3910 8275 -3860 8325
rect -3815 8275 -3765 8325
rect -3715 8275 -3665 8325
rect -3615 8275 -3565 8325
rect -3515 8275 -3465 8325
rect -3420 8275 -3370 8325
rect -3325 8275 -3275 8325
rect -3205 8275 -3155 8325
rect -3110 8275 -3060 8325
rect -3015 8275 -2965 8325
rect -2915 8275 -2865 8325
rect -2815 8275 -2765 8325
rect -2715 8275 -2665 8325
rect -2620 8275 -2570 8325
rect -2525 8275 -2475 8325
rect -2405 8275 -2355 8325
rect -2310 8275 -2260 8325
rect -2215 8275 -2165 8325
rect -2115 8275 -2065 8325
rect -2015 8275 -1965 8325
rect -1915 8275 -1865 8325
rect -1820 8275 -1770 8325
rect -1725 8275 -1675 8325
rect -4805 8175 -4755 8225
rect -4710 8175 -4660 8225
rect -4615 8175 -4565 8225
rect -4515 8175 -4465 8225
rect -4415 8175 -4365 8225
rect -4315 8175 -4265 8225
rect -4220 8175 -4170 8225
rect -4125 8175 -4075 8225
rect -4005 8175 -3955 8225
rect -3910 8175 -3860 8225
rect -3815 8175 -3765 8225
rect -3715 8175 -3665 8225
rect -3615 8175 -3565 8225
rect -3515 8175 -3465 8225
rect -3420 8175 -3370 8225
rect -3325 8175 -3275 8225
rect -3205 8175 -3155 8225
rect -3110 8175 -3060 8225
rect -3015 8175 -2965 8225
rect -2915 8175 -2865 8225
rect -2815 8175 -2765 8225
rect -2715 8175 -2665 8225
rect -2620 8175 -2570 8225
rect -2525 8175 -2475 8225
rect -2405 8175 -2355 8225
rect -2310 8175 -2260 8225
rect -2215 8175 -2165 8225
rect -2115 8175 -2065 8225
rect -2015 8175 -1965 8225
rect -1915 8175 -1865 8225
rect -1820 8175 -1770 8225
rect -1725 8175 -1675 8225
rect -4805 8085 -4755 8135
rect -4710 8085 -4660 8135
rect -4615 8085 -4565 8135
rect -4515 8085 -4465 8135
rect -4415 8085 -4365 8135
rect -4315 8085 -4265 8135
rect -4220 8085 -4170 8135
rect -4125 8085 -4075 8135
rect -4005 8085 -3955 8135
rect -3910 8085 -3860 8135
rect -3815 8085 -3765 8135
rect -3715 8085 -3665 8135
rect -3615 8085 -3565 8135
rect -3515 8085 -3465 8135
rect -3420 8085 -3370 8135
rect -3325 8085 -3275 8135
rect -3205 8085 -3155 8135
rect -3110 8085 -3060 8135
rect -3015 8085 -2965 8135
rect -2915 8085 -2865 8135
rect -2815 8085 -2765 8135
rect -2715 8085 -2665 8135
rect -2620 8085 -2570 8135
rect -2525 8085 -2475 8135
rect -2405 8085 -2355 8135
rect -2310 8085 -2260 8135
rect -2215 8085 -2165 8135
rect -2115 8085 -2065 8135
rect -2015 8085 -1965 8135
rect -1915 8085 -1865 8135
rect -1820 8085 -1770 8135
rect -1725 8085 -1675 8135
rect -4805 7965 -4755 8015
rect -4710 7965 -4660 8015
rect -4615 7965 -4565 8015
rect -4515 7965 -4465 8015
rect -4415 7965 -4365 8015
rect -4315 7965 -4265 8015
rect -4220 7965 -4170 8015
rect -4125 7965 -4075 8015
rect -4005 7965 -3955 8015
rect -3910 7965 -3860 8015
rect -3815 7965 -3765 8015
rect -3715 7965 -3665 8015
rect -3615 7965 -3565 8015
rect -3515 7965 -3465 8015
rect -3420 7965 -3370 8015
rect -3325 7965 -3275 8015
rect -3205 7965 -3155 8015
rect -3110 7965 -3060 8015
rect -3015 7965 -2965 8015
rect -2915 7965 -2865 8015
rect -2815 7965 -2765 8015
rect -2715 7965 -2665 8015
rect -2620 7965 -2570 8015
rect -2525 7965 -2475 8015
rect -2405 7965 -2355 8015
rect -2310 7965 -2260 8015
rect -2215 7965 -2165 8015
rect -2115 7965 -2065 8015
rect -2015 7965 -1965 8015
rect -1915 7965 -1865 8015
rect -1820 7965 -1770 8015
rect -1725 7965 -1675 8015
rect -4805 7875 -4755 7925
rect -4710 7875 -4660 7925
rect -4615 7875 -4565 7925
rect -4515 7875 -4465 7925
rect -4415 7875 -4365 7925
rect -4315 7875 -4265 7925
rect -4220 7875 -4170 7925
rect -4125 7875 -4075 7925
rect -4005 7875 -3955 7925
rect -3910 7875 -3860 7925
rect -3815 7875 -3765 7925
rect -3715 7875 -3665 7925
rect -3615 7875 -3565 7925
rect -3515 7875 -3465 7925
rect -3420 7875 -3370 7925
rect -3325 7875 -3275 7925
rect -3205 7875 -3155 7925
rect -3110 7875 -3060 7925
rect -3015 7875 -2965 7925
rect -2915 7875 -2865 7925
rect -2815 7875 -2765 7925
rect -2715 7875 -2665 7925
rect -2620 7875 -2570 7925
rect -2525 7875 -2475 7925
rect -2405 7875 -2355 7925
rect -2310 7875 -2260 7925
rect -2215 7875 -2165 7925
rect -2115 7875 -2065 7925
rect -2015 7875 -1965 7925
rect -1915 7875 -1865 7925
rect -1820 7875 -1770 7925
rect -1725 7875 -1675 7925
rect -4805 7775 -4755 7825
rect -4710 7775 -4660 7825
rect -4615 7775 -4565 7825
rect -4515 7775 -4465 7825
rect -4415 7775 -4365 7825
rect -4315 7775 -4265 7825
rect -4220 7775 -4170 7825
rect -4125 7775 -4075 7825
rect -4005 7775 -3955 7825
rect -3910 7775 -3860 7825
rect -3815 7775 -3765 7825
rect -3715 7775 -3665 7825
rect -3615 7775 -3565 7825
rect -3515 7775 -3465 7825
rect -3420 7775 -3370 7825
rect -3325 7775 -3275 7825
rect -3205 7775 -3155 7825
rect -3110 7775 -3060 7825
rect -3015 7775 -2965 7825
rect -2915 7775 -2865 7825
rect -2815 7775 -2765 7825
rect -2715 7775 -2665 7825
rect -2620 7775 -2570 7825
rect -2525 7775 -2475 7825
rect -2405 7775 -2355 7825
rect -2310 7775 -2260 7825
rect -2215 7775 -2165 7825
rect -2115 7775 -2065 7825
rect -2015 7775 -1965 7825
rect -1915 7775 -1865 7825
rect -1820 7775 -1770 7825
rect -1725 7775 -1675 7825
rect -4805 7685 -4755 7735
rect -4710 7685 -4660 7735
rect -4615 7685 -4565 7735
rect -4515 7685 -4465 7735
rect -4415 7685 -4365 7735
rect -4315 7685 -4265 7735
rect -4220 7685 -4170 7735
rect -4125 7685 -4075 7735
rect -4005 7685 -3955 7735
rect -3910 7685 -3860 7735
rect -3815 7685 -3765 7735
rect -3715 7685 -3665 7735
rect -3615 7685 -3565 7735
rect -3515 7685 -3465 7735
rect -3420 7685 -3370 7735
rect -3325 7685 -3275 7735
rect -3205 7685 -3155 7735
rect -3110 7685 -3060 7735
rect -3015 7685 -2965 7735
rect -2915 7685 -2865 7735
rect -2815 7685 -2765 7735
rect -2715 7685 -2665 7735
rect -2620 7685 -2570 7735
rect -2525 7685 -2475 7735
rect -2405 7685 -2355 7735
rect -2310 7685 -2260 7735
rect -2215 7685 -2165 7735
rect -2115 7685 -2065 7735
rect -2015 7685 -1965 7735
rect -1915 7685 -1865 7735
rect -1820 7685 -1770 7735
rect -1725 7685 -1675 7735
rect -4805 7565 -4755 7615
rect -4710 7565 -4660 7615
rect -4615 7565 -4565 7615
rect -4515 7565 -4465 7615
rect -4415 7565 -4365 7615
rect -4315 7565 -4265 7615
rect -4220 7565 -4170 7615
rect -4125 7565 -4075 7615
rect -4005 7565 -3955 7615
rect -3910 7565 -3860 7615
rect -3815 7565 -3765 7615
rect -3715 7565 -3665 7615
rect -3615 7565 -3565 7615
rect -3515 7565 -3465 7615
rect -3420 7565 -3370 7615
rect -3325 7565 -3275 7615
rect -3205 7565 -3155 7615
rect -3110 7565 -3060 7615
rect -3015 7565 -2965 7615
rect -2915 7565 -2865 7615
rect -2815 7565 -2765 7615
rect -2715 7565 -2665 7615
rect -2620 7565 -2570 7615
rect -2525 7565 -2475 7615
rect -2405 7565 -2355 7615
rect -2310 7565 -2260 7615
rect -2215 7565 -2165 7615
rect -2115 7565 -2065 7615
rect -2015 7565 -1965 7615
rect -1915 7565 -1865 7615
rect -1820 7565 -1770 7615
rect -1725 7565 -1675 7615
rect -4805 7475 -4755 7525
rect -4710 7475 -4660 7525
rect -4615 7475 -4565 7525
rect -4515 7475 -4465 7525
rect -4415 7475 -4365 7525
rect -4315 7475 -4265 7525
rect -4220 7475 -4170 7525
rect -4125 7475 -4075 7525
rect -4005 7475 -3955 7525
rect -3910 7475 -3860 7525
rect -3815 7475 -3765 7525
rect -3715 7475 -3665 7525
rect -3615 7475 -3565 7525
rect -3515 7475 -3465 7525
rect -3420 7475 -3370 7525
rect -3325 7475 -3275 7525
rect -3205 7475 -3155 7525
rect -3110 7475 -3060 7525
rect -3015 7475 -2965 7525
rect -2915 7475 -2865 7525
rect -2815 7475 -2765 7525
rect -2715 7475 -2665 7525
rect -2620 7475 -2570 7525
rect -2525 7475 -2475 7525
rect -2405 7475 -2355 7525
rect -2310 7475 -2260 7525
rect -2215 7475 -2165 7525
rect -2115 7475 -2065 7525
rect -2015 7475 -1965 7525
rect -1915 7475 -1865 7525
rect -1820 7475 -1770 7525
rect -1725 7475 -1675 7525
rect -4805 7375 -4755 7425
rect -4710 7375 -4660 7425
rect -4615 7375 -4565 7425
rect -4515 7375 -4465 7425
rect -4415 7375 -4365 7425
rect -4315 7375 -4265 7425
rect -4220 7375 -4170 7425
rect -4125 7375 -4075 7425
rect -4005 7375 -3955 7425
rect -3910 7375 -3860 7425
rect -3815 7375 -3765 7425
rect -3715 7375 -3665 7425
rect -3615 7375 -3565 7425
rect -3515 7375 -3465 7425
rect -3420 7375 -3370 7425
rect -3325 7375 -3275 7425
rect -3205 7375 -3155 7425
rect -3110 7375 -3060 7425
rect -3015 7375 -2965 7425
rect -2915 7375 -2865 7425
rect -2815 7375 -2765 7425
rect -2715 7375 -2665 7425
rect -2620 7375 -2570 7425
rect -2525 7375 -2475 7425
rect -2405 7375 -2355 7425
rect -2310 7375 -2260 7425
rect -2215 7375 -2165 7425
rect -2115 7375 -2065 7425
rect -2015 7375 -1965 7425
rect -1915 7375 -1865 7425
rect -1820 7375 -1770 7425
rect -1725 7375 -1675 7425
rect -4805 7285 -4755 7335
rect -4710 7285 -4660 7335
rect -4615 7285 -4565 7335
rect -4515 7285 -4465 7335
rect -4415 7285 -4365 7335
rect -4315 7285 -4265 7335
rect -4220 7285 -4170 7335
rect -4125 7285 -4075 7335
rect -4005 7285 -3955 7335
rect -3910 7285 -3860 7335
rect -3815 7285 -3765 7335
rect -3715 7285 -3665 7335
rect -3615 7285 -3565 7335
rect -3515 7285 -3465 7335
rect -3420 7285 -3370 7335
rect -3325 7285 -3275 7335
rect -3205 7285 -3155 7335
rect -3110 7285 -3060 7335
rect -3015 7285 -2965 7335
rect -2915 7285 -2865 7335
rect -2815 7285 -2765 7335
rect -2715 7285 -2665 7335
rect -2620 7285 -2570 7335
rect -2525 7285 -2475 7335
rect -2405 7285 -2355 7335
rect -2310 7285 -2260 7335
rect -2215 7285 -2165 7335
rect -2115 7285 -2065 7335
rect -2015 7285 -1965 7335
rect -1915 7285 -1865 7335
rect -1820 7285 -1770 7335
rect -1725 7285 -1675 7335
rect -4805 7165 -4755 7215
rect -4710 7165 -4660 7215
rect -4615 7165 -4565 7215
rect -4515 7165 -4465 7215
rect -4415 7165 -4365 7215
rect -4315 7165 -4265 7215
rect -4220 7165 -4170 7215
rect -4125 7165 -4075 7215
rect -4005 7165 -3955 7215
rect -3910 7165 -3860 7215
rect -3815 7165 -3765 7215
rect -3715 7165 -3665 7215
rect -3615 7165 -3565 7215
rect -3515 7165 -3465 7215
rect -3420 7165 -3370 7215
rect -3325 7165 -3275 7215
rect -3205 7165 -3155 7215
rect -3110 7165 -3060 7215
rect -3015 7165 -2965 7215
rect -2915 7165 -2865 7215
rect -2815 7165 -2765 7215
rect -2715 7165 -2665 7215
rect -2620 7165 -2570 7215
rect -2525 7165 -2475 7215
rect -2405 7165 -2355 7215
rect -2310 7165 -2260 7215
rect -2215 7165 -2165 7215
rect -2115 7165 -2065 7215
rect -2015 7165 -1965 7215
rect -1915 7165 -1865 7215
rect -1820 7165 -1770 7215
rect -1725 7165 -1675 7215
rect -4805 7075 -4755 7125
rect -4710 7075 -4660 7125
rect -4615 7075 -4565 7125
rect -4515 7075 -4465 7125
rect -4415 7075 -4365 7125
rect -4315 7075 -4265 7125
rect -4220 7075 -4170 7125
rect -4125 7075 -4075 7125
rect -4005 7075 -3955 7125
rect -3910 7075 -3860 7125
rect -3815 7075 -3765 7125
rect -3715 7075 -3665 7125
rect -3615 7075 -3565 7125
rect -3515 7075 -3465 7125
rect -3420 7075 -3370 7125
rect -3325 7075 -3275 7125
rect -3205 7075 -3155 7125
rect -3110 7075 -3060 7125
rect -3015 7075 -2965 7125
rect -2915 7075 -2865 7125
rect -2815 7075 -2765 7125
rect -2715 7075 -2665 7125
rect -2620 7075 -2570 7125
rect -2525 7075 -2475 7125
rect -2405 7075 -2355 7125
rect -2310 7075 -2260 7125
rect -2215 7075 -2165 7125
rect -2115 7075 -2065 7125
rect -2015 7075 -1965 7125
rect -1915 7075 -1865 7125
rect -1820 7075 -1770 7125
rect -1725 7075 -1675 7125
rect -4805 6975 -4755 7025
rect -4710 6975 -4660 7025
rect -4615 6975 -4565 7025
rect -4515 6975 -4465 7025
rect -4415 6975 -4365 7025
rect -4315 6975 -4265 7025
rect -4220 6975 -4170 7025
rect -4125 6975 -4075 7025
rect -4005 6975 -3955 7025
rect -3910 6975 -3860 7025
rect -3815 6975 -3765 7025
rect -3715 6975 -3665 7025
rect -3615 6975 -3565 7025
rect -3515 6975 -3465 7025
rect -3420 6975 -3370 7025
rect -3325 6975 -3275 7025
rect -3205 6975 -3155 7025
rect -3110 6975 -3060 7025
rect -3015 6975 -2965 7025
rect -2915 6975 -2865 7025
rect -2815 6975 -2765 7025
rect -2715 6975 -2665 7025
rect -2620 6975 -2570 7025
rect -2525 6975 -2475 7025
rect -2405 6975 -2355 7025
rect -2310 6975 -2260 7025
rect -2215 6975 -2165 7025
rect -2115 6975 -2065 7025
rect -2015 6975 -1965 7025
rect -1915 6975 -1865 7025
rect -1820 6975 -1770 7025
rect -1725 6975 -1675 7025
rect -4805 6885 -4755 6935
rect -4710 6885 -4660 6935
rect -4615 6885 -4565 6935
rect -4515 6885 -4465 6935
rect -4415 6885 -4365 6935
rect -4315 6885 -4265 6935
rect -4220 6885 -4170 6935
rect -4125 6885 -4075 6935
rect -4005 6885 -3955 6935
rect -3910 6885 -3860 6935
rect -3815 6885 -3765 6935
rect -3715 6885 -3665 6935
rect -3615 6885 -3565 6935
rect -3515 6885 -3465 6935
rect -3420 6885 -3370 6935
rect -3325 6885 -3275 6935
rect -3205 6885 -3155 6935
rect -3110 6885 -3060 6935
rect -3015 6885 -2965 6935
rect -2915 6885 -2865 6935
rect -2815 6885 -2765 6935
rect -2715 6885 -2665 6935
rect -2620 6885 -2570 6935
rect -2525 6885 -2475 6935
rect -2405 6885 -2355 6935
rect -2310 6885 -2260 6935
rect -2215 6885 -2165 6935
rect -2115 6885 -2065 6935
rect -2015 6885 -1965 6935
rect -1915 6885 -1865 6935
rect -1820 6885 -1770 6935
rect -1725 6885 -1675 6935
rect -4805 6765 -4755 6815
rect -4710 6765 -4660 6815
rect -4615 6765 -4565 6815
rect -4515 6765 -4465 6815
rect -4415 6765 -4365 6815
rect -4315 6765 -4265 6815
rect -4220 6765 -4170 6815
rect -4125 6765 -4075 6815
rect -4005 6765 -3955 6815
rect -3910 6765 -3860 6815
rect -3815 6765 -3765 6815
rect -3715 6765 -3665 6815
rect -3615 6765 -3565 6815
rect -3515 6765 -3465 6815
rect -3420 6765 -3370 6815
rect -3325 6765 -3275 6815
rect -3205 6765 -3155 6815
rect -3110 6765 -3060 6815
rect -3015 6765 -2965 6815
rect -2915 6765 -2865 6815
rect -2815 6765 -2765 6815
rect -2715 6765 -2665 6815
rect -2620 6765 -2570 6815
rect -2525 6765 -2475 6815
rect -2405 6765 -2355 6815
rect -2310 6765 -2260 6815
rect -2215 6765 -2165 6815
rect -2115 6765 -2065 6815
rect -2015 6765 -1965 6815
rect -1915 6765 -1865 6815
rect -1820 6765 -1770 6815
rect -1725 6765 -1675 6815
rect -4805 6675 -4755 6725
rect -4710 6675 -4660 6725
rect -4615 6675 -4565 6725
rect -4515 6675 -4465 6725
rect -4415 6675 -4365 6725
rect -4315 6675 -4265 6725
rect -4220 6675 -4170 6725
rect -4125 6675 -4075 6725
rect -4005 6675 -3955 6725
rect -3910 6675 -3860 6725
rect -3815 6675 -3765 6725
rect -3715 6675 -3665 6725
rect -3615 6675 -3565 6725
rect -3515 6675 -3465 6725
rect -3420 6675 -3370 6725
rect -3325 6675 -3275 6725
rect -3205 6675 -3155 6725
rect -3110 6675 -3060 6725
rect -3015 6675 -2965 6725
rect -2915 6675 -2865 6725
rect -2815 6675 -2765 6725
rect -2715 6675 -2665 6725
rect -2620 6675 -2570 6725
rect -2525 6675 -2475 6725
rect -2405 6675 -2355 6725
rect -2310 6675 -2260 6725
rect -2215 6675 -2165 6725
rect -2115 6675 -2065 6725
rect -2015 6675 -1965 6725
rect -1915 6675 -1865 6725
rect -1820 6675 -1770 6725
rect -1725 6675 -1675 6725
rect -4805 6575 -4755 6625
rect -4710 6575 -4660 6625
rect -4615 6575 -4565 6625
rect -4515 6575 -4465 6625
rect -4415 6575 -4365 6625
rect -4315 6575 -4265 6625
rect -4220 6575 -4170 6625
rect -4125 6575 -4075 6625
rect -4005 6575 -3955 6625
rect -3910 6575 -3860 6625
rect -3815 6575 -3765 6625
rect -3715 6575 -3665 6625
rect -3615 6575 -3565 6625
rect -3515 6575 -3465 6625
rect -3420 6575 -3370 6625
rect -3325 6575 -3275 6625
rect -3205 6575 -3155 6625
rect -3110 6575 -3060 6625
rect -3015 6575 -2965 6625
rect -2915 6575 -2865 6625
rect -2815 6575 -2765 6625
rect -2715 6575 -2665 6625
rect -2620 6575 -2570 6625
rect -2525 6575 -2475 6625
rect -2405 6575 -2355 6625
rect -2310 6575 -2260 6625
rect -2215 6575 -2165 6625
rect -2115 6575 -2065 6625
rect -2015 6575 -1965 6625
rect -1915 6575 -1865 6625
rect -1820 6575 -1770 6625
rect -1725 6575 -1675 6625
rect -4805 6485 -4755 6535
rect -4710 6485 -4660 6535
rect -4615 6485 -4565 6535
rect -4515 6485 -4465 6535
rect -4415 6485 -4365 6535
rect -4315 6485 -4265 6535
rect -4220 6485 -4170 6535
rect -4125 6485 -4075 6535
rect -4005 6485 -3955 6535
rect -3910 6485 -3860 6535
rect -3815 6485 -3765 6535
rect -3715 6485 -3665 6535
rect -3615 6485 -3565 6535
rect -3515 6485 -3465 6535
rect -3420 6485 -3370 6535
rect -3325 6485 -3275 6535
rect -3205 6485 -3155 6535
rect -3110 6485 -3060 6535
rect -3015 6485 -2965 6535
rect -2915 6485 -2865 6535
rect -2815 6485 -2765 6535
rect -2715 6485 -2665 6535
rect -2620 6485 -2570 6535
rect -2525 6485 -2475 6535
rect -2405 6485 -2355 6535
rect -2310 6485 -2260 6535
rect -2215 6485 -2165 6535
rect -2115 6485 -2065 6535
rect -2015 6485 -1965 6535
rect -1915 6485 -1865 6535
rect -1820 6485 -1770 6535
rect -1725 6485 -1675 6535
rect -80 9635 -40 9640
rect -80 9605 -75 9635
rect -75 9605 -45 9635
rect -45 9605 -40 9635
rect -80 9600 -40 9605
rect -80 9570 -40 9575
rect -80 9540 -75 9570
rect -75 9540 -45 9570
rect -45 9540 -40 9570
rect -80 9535 -40 9540
rect -80 9500 -40 9505
rect -80 9470 -75 9500
rect -75 9470 -45 9500
rect -45 9470 -40 9500
rect -80 9465 -40 9470
rect -80 9430 -40 9435
rect -80 9400 -75 9430
rect -75 9400 -45 9430
rect -45 9400 -40 9430
rect -80 9395 -40 9400
rect -80 9360 -40 9365
rect -80 9330 -75 9360
rect -75 9330 -45 9360
rect -45 9330 -40 9360
rect -80 9325 -40 9330
rect -80 9295 -40 9300
rect -80 9265 -75 9295
rect -75 9265 -45 9295
rect -45 9265 -40 9295
rect -80 9260 -40 9265
rect -80 9235 -40 9240
rect -80 9205 -75 9235
rect -75 9205 -45 9235
rect -45 9205 -40 9235
rect -80 9200 -40 9205
rect -80 9170 -40 9175
rect -80 9140 -75 9170
rect -75 9140 -45 9170
rect -45 9140 -40 9170
rect -80 9135 -40 9140
rect -80 9100 -40 9105
rect -80 9070 -75 9100
rect -75 9070 -45 9100
rect -45 9070 -40 9100
rect -80 9065 -40 9070
rect -80 9030 -40 9035
rect -80 9000 -75 9030
rect -75 9000 -45 9030
rect -45 9000 -40 9030
rect -80 8995 -40 9000
rect -80 8960 -40 8965
rect -80 8930 -75 8960
rect -75 8930 -45 8960
rect -45 8930 -40 8960
rect -80 8925 -40 8930
rect -80 8895 -40 8900
rect -80 8865 -75 8895
rect -75 8865 -45 8895
rect -45 8865 -40 8895
rect -80 8860 -40 8865
rect -80 8835 -40 8840
rect -80 8805 -75 8835
rect -75 8805 -45 8835
rect -45 8805 -40 8835
rect -80 8800 -40 8805
rect -80 8770 -40 8775
rect -80 8740 -75 8770
rect -75 8740 -45 8770
rect -45 8740 -40 8770
rect -80 8735 -40 8740
rect -80 8700 -40 8705
rect -80 8670 -75 8700
rect -75 8670 -45 8700
rect -45 8670 -40 8700
rect -80 8665 -40 8670
rect -80 8630 -40 8635
rect -80 8600 -75 8630
rect -75 8600 -45 8630
rect -45 8600 -40 8630
rect -80 8595 -40 8600
rect -80 8560 -40 8565
rect -80 8530 -75 8560
rect -75 8530 -45 8560
rect -45 8530 -40 8560
rect -80 8525 -40 8530
rect -80 8495 -40 8500
rect -80 8465 -75 8495
rect -75 8465 -45 8495
rect -45 8465 -40 8495
rect -80 8460 -40 8465
rect -80 8435 -40 8440
rect -80 8405 -75 8435
rect -75 8405 -45 8435
rect -45 8405 -40 8435
rect -80 8400 -40 8405
rect -80 8370 -40 8375
rect -80 8340 -75 8370
rect -75 8340 -45 8370
rect -45 8340 -40 8370
rect -80 8335 -40 8340
rect -80 8300 -40 8305
rect -80 8270 -75 8300
rect -75 8270 -45 8300
rect -45 8270 -40 8300
rect -80 8265 -40 8270
rect -80 8230 -40 8235
rect -80 8200 -75 8230
rect -75 8200 -45 8230
rect -45 8200 -40 8230
rect -80 8195 -40 8200
rect -80 8160 -40 8165
rect -80 8130 -75 8160
rect -75 8130 -45 8160
rect -45 8130 -40 8160
rect -80 8125 -40 8130
rect -80 8095 -40 8100
rect -80 8065 -75 8095
rect -75 8065 -45 8095
rect -45 8065 -40 8095
rect -80 8060 -40 8065
rect -80 8035 -40 8040
rect -80 8005 -75 8035
rect -75 8005 -45 8035
rect -45 8005 -40 8035
rect -80 8000 -40 8005
rect -80 7970 -40 7975
rect -80 7940 -75 7970
rect -75 7940 -45 7970
rect -45 7940 -40 7970
rect -80 7935 -40 7940
rect -80 7900 -40 7905
rect -80 7870 -75 7900
rect -75 7870 -45 7900
rect -45 7870 -40 7900
rect -80 7865 -40 7870
rect -80 7830 -40 7835
rect -80 7800 -75 7830
rect -75 7800 -45 7830
rect -45 7800 -40 7830
rect -80 7795 -40 7800
rect -80 7760 -40 7765
rect -80 7730 -75 7760
rect -75 7730 -45 7760
rect -45 7730 -40 7760
rect -80 7725 -40 7730
rect -80 7695 -40 7700
rect -80 7665 -75 7695
rect -75 7665 -45 7695
rect -45 7665 -40 7695
rect -80 7660 -40 7665
rect -80 7635 -40 7640
rect -80 7605 -75 7635
rect -75 7605 -45 7635
rect -45 7605 -40 7635
rect -80 7600 -40 7605
rect -80 7570 -40 7575
rect -80 7540 -75 7570
rect -75 7540 -45 7570
rect -45 7540 -40 7570
rect -80 7535 -40 7540
rect -80 7500 -40 7505
rect -80 7470 -75 7500
rect -75 7470 -45 7500
rect -45 7470 -40 7500
rect -80 7465 -40 7470
rect -80 7430 -40 7435
rect -80 7400 -75 7430
rect -75 7400 -45 7430
rect -45 7400 -40 7430
rect -80 7395 -40 7400
rect -80 7360 -40 7365
rect -80 7330 -75 7360
rect -75 7330 -45 7360
rect -45 7330 -40 7360
rect -80 7325 -40 7330
rect -80 7295 -40 7300
rect -80 7265 -75 7295
rect -75 7265 -45 7295
rect -45 7265 -40 7295
rect -80 7260 -40 7265
rect -80 7235 -40 7240
rect -80 7205 -75 7235
rect -75 7205 -45 7235
rect -45 7205 -40 7235
rect -80 7200 -40 7205
rect -80 7170 -40 7175
rect -80 7140 -75 7170
rect -75 7140 -45 7170
rect -45 7140 -40 7170
rect -80 7135 -40 7140
rect -80 7100 -40 7105
rect -80 7070 -75 7100
rect -75 7070 -45 7100
rect -45 7070 -40 7100
rect -80 7065 -40 7070
rect -80 7030 -40 7035
rect -80 7000 -75 7030
rect -75 7000 -45 7030
rect -45 7000 -40 7030
rect -80 6995 -40 7000
rect -80 6960 -40 6965
rect -80 6930 -75 6960
rect -75 6930 -45 6960
rect -45 6930 -40 6960
rect -80 6925 -40 6930
rect -80 6895 -40 6900
rect -80 6865 -75 6895
rect -75 6865 -45 6895
rect -45 6865 -40 6895
rect -80 6860 -40 6865
rect -80 6835 -40 6840
rect -80 6805 -75 6835
rect -75 6805 -45 6835
rect -45 6805 -40 6835
rect -80 6800 -40 6805
rect -80 6770 -40 6775
rect -80 6740 -75 6770
rect -75 6740 -45 6770
rect -45 6740 -40 6770
rect -80 6735 -40 6740
rect -80 6700 -40 6705
rect -80 6670 -75 6700
rect -75 6670 -45 6700
rect -45 6670 -40 6700
rect -80 6665 -40 6670
rect -80 6630 -40 6635
rect -80 6600 -75 6630
rect -75 6600 -45 6630
rect -45 6600 -40 6630
rect -80 6595 -40 6600
rect -80 6560 -40 6565
rect -80 6530 -75 6560
rect -75 6530 -45 6560
rect -45 6530 -40 6560
rect -80 6525 -40 6530
rect -80 6495 -40 6500
rect -80 6465 -75 6495
rect -75 6465 -45 6495
rect -45 6465 -40 6495
rect -80 6460 -40 6465
rect 270 9635 310 9640
rect 270 9605 275 9635
rect 275 9605 305 9635
rect 305 9605 310 9635
rect 270 9600 310 9605
rect 270 9570 310 9575
rect 270 9540 275 9570
rect 275 9540 305 9570
rect 305 9540 310 9570
rect 270 9535 310 9540
rect 270 9500 310 9505
rect 270 9470 275 9500
rect 275 9470 305 9500
rect 305 9470 310 9500
rect 270 9465 310 9470
rect 270 9430 310 9435
rect 270 9400 275 9430
rect 275 9400 305 9430
rect 305 9400 310 9430
rect 270 9395 310 9400
rect 270 9360 310 9365
rect 270 9330 275 9360
rect 275 9330 305 9360
rect 305 9330 310 9360
rect 270 9325 310 9330
rect 270 9295 310 9300
rect 270 9265 275 9295
rect 275 9265 305 9295
rect 305 9265 310 9295
rect 270 9260 310 9265
rect 270 9235 310 9240
rect 270 9205 275 9235
rect 275 9205 305 9235
rect 305 9205 310 9235
rect 270 9200 310 9205
rect 270 9170 310 9175
rect 270 9140 275 9170
rect 275 9140 305 9170
rect 305 9140 310 9170
rect 270 9135 310 9140
rect 270 9100 310 9105
rect 270 9070 275 9100
rect 275 9070 305 9100
rect 305 9070 310 9100
rect 270 9065 310 9070
rect 270 9030 310 9035
rect 270 9000 275 9030
rect 275 9000 305 9030
rect 305 9000 310 9030
rect 270 8995 310 9000
rect 270 8960 310 8965
rect 270 8930 275 8960
rect 275 8930 305 8960
rect 305 8930 310 8960
rect 270 8925 310 8930
rect 270 8895 310 8900
rect 270 8865 275 8895
rect 275 8865 305 8895
rect 305 8865 310 8895
rect 270 8860 310 8865
rect 270 8835 310 8840
rect 270 8805 275 8835
rect 275 8805 305 8835
rect 305 8805 310 8835
rect 270 8800 310 8805
rect 270 8770 310 8775
rect 270 8740 275 8770
rect 275 8740 305 8770
rect 305 8740 310 8770
rect 270 8735 310 8740
rect 270 8700 310 8705
rect 270 8670 275 8700
rect 275 8670 305 8700
rect 305 8670 310 8700
rect 270 8665 310 8670
rect 270 8630 310 8635
rect 270 8600 275 8630
rect 275 8600 305 8630
rect 305 8600 310 8630
rect 270 8595 310 8600
rect 270 8560 310 8565
rect 270 8530 275 8560
rect 275 8530 305 8560
rect 305 8530 310 8560
rect 270 8525 310 8530
rect 270 8495 310 8500
rect 270 8465 275 8495
rect 275 8465 305 8495
rect 305 8465 310 8495
rect 270 8460 310 8465
rect 270 8435 310 8440
rect 270 8405 275 8435
rect 275 8405 305 8435
rect 305 8405 310 8435
rect 270 8400 310 8405
rect 270 8370 310 8375
rect 270 8340 275 8370
rect 275 8340 305 8370
rect 305 8340 310 8370
rect 270 8335 310 8340
rect 270 8300 310 8305
rect 270 8270 275 8300
rect 275 8270 305 8300
rect 305 8270 310 8300
rect 270 8265 310 8270
rect 270 8230 310 8235
rect 270 8200 275 8230
rect 275 8200 305 8230
rect 305 8200 310 8230
rect 270 8195 310 8200
rect 270 8160 310 8165
rect 270 8130 275 8160
rect 275 8130 305 8160
rect 305 8130 310 8160
rect 270 8125 310 8130
rect 270 8095 310 8100
rect 270 8065 275 8095
rect 275 8065 305 8095
rect 305 8065 310 8095
rect 270 8060 310 8065
rect 270 8035 310 8040
rect 270 8005 275 8035
rect 275 8005 305 8035
rect 305 8005 310 8035
rect 270 8000 310 8005
rect 270 7970 310 7975
rect 270 7940 275 7970
rect 275 7940 305 7970
rect 305 7940 310 7970
rect 270 7935 310 7940
rect 270 7900 310 7905
rect 270 7870 275 7900
rect 275 7870 305 7900
rect 305 7870 310 7900
rect 270 7865 310 7870
rect 270 7830 310 7835
rect 270 7800 275 7830
rect 275 7800 305 7830
rect 305 7800 310 7830
rect 270 7795 310 7800
rect 270 7760 310 7765
rect 270 7730 275 7760
rect 275 7730 305 7760
rect 305 7730 310 7760
rect 270 7725 310 7730
rect 270 7695 310 7700
rect 270 7665 275 7695
rect 275 7665 305 7695
rect 305 7665 310 7695
rect 270 7660 310 7665
rect 270 7635 310 7640
rect 270 7605 275 7635
rect 275 7605 305 7635
rect 305 7605 310 7635
rect 270 7600 310 7605
rect 270 7570 310 7575
rect 270 7540 275 7570
rect 275 7540 305 7570
rect 305 7540 310 7570
rect 270 7535 310 7540
rect 270 7500 310 7505
rect 270 7470 275 7500
rect 275 7470 305 7500
rect 305 7470 310 7500
rect 270 7465 310 7470
rect 270 7430 310 7435
rect 270 7400 275 7430
rect 275 7400 305 7430
rect 305 7400 310 7430
rect 270 7395 310 7400
rect 270 7360 310 7365
rect 270 7330 275 7360
rect 275 7330 305 7360
rect 305 7330 310 7360
rect 270 7325 310 7330
rect 270 7295 310 7300
rect 270 7265 275 7295
rect 275 7265 305 7295
rect 305 7265 310 7295
rect 270 7260 310 7265
rect 270 7235 310 7240
rect 270 7205 275 7235
rect 275 7205 305 7235
rect 305 7205 310 7235
rect 270 7200 310 7205
rect 270 7170 310 7175
rect 270 7140 275 7170
rect 275 7140 305 7170
rect 305 7140 310 7170
rect 270 7135 310 7140
rect 270 7100 310 7105
rect 270 7070 275 7100
rect 275 7070 305 7100
rect 305 7070 310 7100
rect 270 7065 310 7070
rect 270 7030 310 7035
rect 270 7000 275 7030
rect 275 7000 305 7030
rect 305 7000 310 7030
rect 270 6995 310 7000
rect 270 6960 310 6965
rect 270 6930 275 6960
rect 275 6930 305 6960
rect 305 6930 310 6960
rect 270 6925 310 6930
rect 270 6895 310 6900
rect 270 6865 275 6895
rect 275 6865 305 6895
rect 305 6865 310 6895
rect 270 6860 310 6865
rect 270 6835 310 6840
rect 270 6805 275 6835
rect 275 6805 305 6835
rect 305 6805 310 6835
rect 270 6800 310 6805
rect 270 6770 310 6775
rect 270 6740 275 6770
rect 275 6740 305 6770
rect 305 6740 310 6770
rect 270 6735 310 6740
rect 270 6700 310 6705
rect 270 6670 275 6700
rect 275 6670 305 6700
rect 305 6670 310 6700
rect 270 6665 310 6670
rect 270 6630 310 6635
rect 270 6600 275 6630
rect 275 6600 305 6630
rect 305 6600 310 6630
rect 270 6595 310 6600
rect 270 6560 310 6565
rect 270 6530 275 6560
rect 275 6530 305 6560
rect 305 6530 310 6560
rect 270 6525 310 6530
rect 270 6495 310 6500
rect 270 6465 275 6495
rect 275 6465 305 6495
rect 305 6465 310 6495
rect 270 6460 310 6465
rect 620 9635 660 9640
rect 620 9605 625 9635
rect 625 9605 655 9635
rect 655 9605 660 9635
rect 620 9600 660 9605
rect 620 9570 660 9575
rect 620 9540 625 9570
rect 625 9540 655 9570
rect 655 9540 660 9570
rect 620 9535 660 9540
rect 620 9500 660 9505
rect 620 9470 625 9500
rect 625 9470 655 9500
rect 655 9470 660 9500
rect 620 9465 660 9470
rect 620 9430 660 9435
rect 620 9400 625 9430
rect 625 9400 655 9430
rect 655 9400 660 9430
rect 620 9395 660 9400
rect 620 9360 660 9365
rect 620 9330 625 9360
rect 625 9330 655 9360
rect 655 9330 660 9360
rect 620 9325 660 9330
rect 620 9295 660 9300
rect 620 9265 625 9295
rect 625 9265 655 9295
rect 655 9265 660 9295
rect 620 9260 660 9265
rect 620 9235 660 9240
rect 620 9205 625 9235
rect 625 9205 655 9235
rect 655 9205 660 9235
rect 620 9200 660 9205
rect 620 9170 660 9175
rect 620 9140 625 9170
rect 625 9140 655 9170
rect 655 9140 660 9170
rect 620 9135 660 9140
rect 620 9100 660 9105
rect 620 9070 625 9100
rect 625 9070 655 9100
rect 655 9070 660 9100
rect 620 9065 660 9070
rect 620 9030 660 9035
rect 620 9000 625 9030
rect 625 9000 655 9030
rect 655 9000 660 9030
rect 620 8995 660 9000
rect 620 8960 660 8965
rect 620 8930 625 8960
rect 625 8930 655 8960
rect 655 8930 660 8960
rect 620 8925 660 8930
rect 620 8895 660 8900
rect 620 8865 625 8895
rect 625 8865 655 8895
rect 655 8865 660 8895
rect 620 8860 660 8865
rect 620 8835 660 8840
rect 620 8805 625 8835
rect 625 8805 655 8835
rect 655 8805 660 8835
rect 620 8800 660 8805
rect 620 8770 660 8775
rect 620 8740 625 8770
rect 625 8740 655 8770
rect 655 8740 660 8770
rect 620 8735 660 8740
rect 620 8700 660 8705
rect 620 8670 625 8700
rect 625 8670 655 8700
rect 655 8670 660 8700
rect 620 8665 660 8670
rect 620 8630 660 8635
rect 620 8600 625 8630
rect 625 8600 655 8630
rect 655 8600 660 8630
rect 620 8595 660 8600
rect 620 8560 660 8565
rect 620 8530 625 8560
rect 625 8530 655 8560
rect 655 8530 660 8560
rect 620 8525 660 8530
rect 620 8495 660 8500
rect 620 8465 625 8495
rect 625 8465 655 8495
rect 655 8465 660 8495
rect 620 8460 660 8465
rect 620 8435 660 8440
rect 620 8405 625 8435
rect 625 8405 655 8435
rect 655 8405 660 8435
rect 620 8400 660 8405
rect 620 8370 660 8375
rect 620 8340 625 8370
rect 625 8340 655 8370
rect 655 8340 660 8370
rect 620 8335 660 8340
rect 620 8300 660 8305
rect 620 8270 625 8300
rect 625 8270 655 8300
rect 655 8270 660 8300
rect 620 8265 660 8270
rect 620 8230 660 8235
rect 620 8200 625 8230
rect 625 8200 655 8230
rect 655 8200 660 8230
rect 620 8195 660 8200
rect 620 8160 660 8165
rect 620 8130 625 8160
rect 625 8130 655 8160
rect 655 8130 660 8160
rect 620 8125 660 8130
rect 620 8095 660 8100
rect 620 8065 625 8095
rect 625 8065 655 8095
rect 655 8065 660 8095
rect 620 8060 660 8065
rect 620 8035 660 8040
rect 620 8005 625 8035
rect 625 8005 655 8035
rect 655 8005 660 8035
rect 620 8000 660 8005
rect 620 7970 660 7975
rect 620 7940 625 7970
rect 625 7940 655 7970
rect 655 7940 660 7970
rect 620 7935 660 7940
rect 620 7900 660 7905
rect 620 7870 625 7900
rect 625 7870 655 7900
rect 655 7870 660 7900
rect 620 7865 660 7870
rect 620 7830 660 7835
rect 620 7800 625 7830
rect 625 7800 655 7830
rect 655 7800 660 7830
rect 620 7795 660 7800
rect 620 7760 660 7765
rect 620 7730 625 7760
rect 625 7730 655 7760
rect 655 7730 660 7760
rect 620 7725 660 7730
rect 620 7695 660 7700
rect 620 7665 625 7695
rect 625 7665 655 7695
rect 655 7665 660 7695
rect 620 7660 660 7665
rect 620 7635 660 7640
rect 620 7605 625 7635
rect 625 7605 655 7635
rect 655 7605 660 7635
rect 620 7600 660 7605
rect 620 7570 660 7575
rect 620 7540 625 7570
rect 625 7540 655 7570
rect 655 7540 660 7570
rect 620 7535 660 7540
rect 620 7500 660 7505
rect 620 7470 625 7500
rect 625 7470 655 7500
rect 655 7470 660 7500
rect 620 7465 660 7470
rect 620 7430 660 7435
rect 620 7400 625 7430
rect 625 7400 655 7430
rect 655 7400 660 7430
rect 620 7395 660 7400
rect 620 7360 660 7365
rect 620 7330 625 7360
rect 625 7330 655 7360
rect 655 7330 660 7360
rect 620 7325 660 7330
rect 620 7295 660 7300
rect 620 7265 625 7295
rect 625 7265 655 7295
rect 655 7265 660 7295
rect 620 7260 660 7265
rect 620 7235 660 7240
rect 620 7205 625 7235
rect 625 7205 655 7235
rect 655 7205 660 7235
rect 620 7200 660 7205
rect 620 7170 660 7175
rect 620 7140 625 7170
rect 625 7140 655 7170
rect 655 7140 660 7170
rect 620 7135 660 7140
rect 620 7100 660 7105
rect 620 7070 625 7100
rect 625 7070 655 7100
rect 655 7070 660 7100
rect 620 7065 660 7070
rect 620 7030 660 7035
rect 620 7000 625 7030
rect 625 7000 655 7030
rect 655 7000 660 7030
rect 620 6995 660 7000
rect 620 6960 660 6965
rect 620 6930 625 6960
rect 625 6930 655 6960
rect 655 6930 660 6960
rect 620 6925 660 6930
rect 620 6895 660 6900
rect 620 6865 625 6895
rect 625 6865 655 6895
rect 655 6865 660 6895
rect 620 6860 660 6865
rect 620 6835 660 6840
rect 620 6805 625 6835
rect 625 6805 655 6835
rect 655 6805 660 6835
rect 620 6800 660 6805
rect 620 6770 660 6775
rect 620 6740 625 6770
rect 625 6740 655 6770
rect 655 6740 660 6770
rect 620 6735 660 6740
rect 620 6700 660 6705
rect 620 6670 625 6700
rect 625 6670 655 6700
rect 655 6670 660 6700
rect 620 6665 660 6670
rect 620 6630 660 6635
rect 620 6600 625 6630
rect 625 6600 655 6630
rect 655 6600 660 6630
rect 620 6595 660 6600
rect 620 6560 660 6565
rect 620 6530 625 6560
rect 625 6530 655 6560
rect 655 6530 660 6560
rect 620 6525 660 6530
rect 620 6495 660 6500
rect 620 6465 625 6495
rect 625 6465 655 6495
rect 655 6465 660 6495
rect 620 6460 660 6465
rect 1320 9635 1360 9640
rect 1320 9605 1325 9635
rect 1325 9605 1355 9635
rect 1355 9605 1360 9635
rect 1320 9600 1360 9605
rect 1320 9570 1360 9575
rect 1320 9540 1325 9570
rect 1325 9540 1355 9570
rect 1355 9540 1360 9570
rect 1320 9535 1360 9540
rect 1320 9500 1360 9505
rect 1320 9470 1325 9500
rect 1325 9470 1355 9500
rect 1355 9470 1360 9500
rect 1320 9465 1360 9470
rect 1320 9430 1360 9435
rect 1320 9400 1325 9430
rect 1325 9400 1355 9430
rect 1355 9400 1360 9430
rect 1320 9395 1360 9400
rect 1320 9360 1360 9365
rect 1320 9330 1325 9360
rect 1325 9330 1355 9360
rect 1355 9330 1360 9360
rect 1320 9325 1360 9330
rect 1320 9295 1360 9300
rect 1320 9265 1325 9295
rect 1325 9265 1355 9295
rect 1355 9265 1360 9295
rect 1320 9260 1360 9265
rect 1320 9235 1360 9240
rect 1320 9205 1325 9235
rect 1325 9205 1355 9235
rect 1355 9205 1360 9235
rect 1320 9200 1360 9205
rect 1320 9170 1360 9175
rect 1320 9140 1325 9170
rect 1325 9140 1355 9170
rect 1355 9140 1360 9170
rect 1320 9135 1360 9140
rect 1320 9100 1360 9105
rect 1320 9070 1325 9100
rect 1325 9070 1355 9100
rect 1355 9070 1360 9100
rect 1320 9065 1360 9070
rect 1320 9030 1360 9035
rect 1320 9000 1325 9030
rect 1325 9000 1355 9030
rect 1355 9000 1360 9030
rect 1320 8995 1360 9000
rect 1320 8960 1360 8965
rect 1320 8930 1325 8960
rect 1325 8930 1355 8960
rect 1355 8930 1360 8960
rect 1320 8925 1360 8930
rect 1320 8895 1360 8900
rect 1320 8865 1325 8895
rect 1325 8865 1355 8895
rect 1355 8865 1360 8895
rect 1320 8860 1360 8865
rect 1320 8835 1360 8840
rect 1320 8805 1325 8835
rect 1325 8805 1355 8835
rect 1355 8805 1360 8835
rect 1320 8800 1360 8805
rect 1320 8770 1360 8775
rect 1320 8740 1325 8770
rect 1325 8740 1355 8770
rect 1355 8740 1360 8770
rect 1320 8735 1360 8740
rect 1320 8700 1360 8705
rect 1320 8670 1325 8700
rect 1325 8670 1355 8700
rect 1355 8670 1360 8700
rect 1320 8665 1360 8670
rect 1320 8630 1360 8635
rect 1320 8600 1325 8630
rect 1325 8600 1355 8630
rect 1355 8600 1360 8630
rect 1320 8595 1360 8600
rect 1320 8560 1360 8565
rect 1320 8530 1325 8560
rect 1325 8530 1355 8560
rect 1355 8530 1360 8560
rect 1320 8525 1360 8530
rect 1320 8495 1360 8500
rect 1320 8465 1325 8495
rect 1325 8465 1355 8495
rect 1355 8465 1360 8495
rect 1320 8460 1360 8465
rect 1320 8435 1360 8440
rect 1320 8405 1325 8435
rect 1325 8405 1355 8435
rect 1355 8405 1360 8435
rect 1320 8400 1360 8405
rect 1320 8370 1360 8375
rect 1320 8340 1325 8370
rect 1325 8340 1355 8370
rect 1355 8340 1360 8370
rect 1320 8335 1360 8340
rect 1320 8300 1360 8305
rect 1320 8270 1325 8300
rect 1325 8270 1355 8300
rect 1355 8270 1360 8300
rect 1320 8265 1360 8270
rect 1320 8230 1360 8235
rect 1320 8200 1325 8230
rect 1325 8200 1355 8230
rect 1355 8200 1360 8230
rect 1320 8195 1360 8200
rect 1320 8160 1360 8165
rect 1320 8130 1325 8160
rect 1325 8130 1355 8160
rect 1355 8130 1360 8160
rect 1320 8125 1360 8130
rect 1320 8095 1360 8100
rect 1320 8065 1325 8095
rect 1325 8065 1355 8095
rect 1355 8065 1360 8095
rect 1320 8060 1360 8065
rect 1320 8035 1360 8040
rect 1320 8005 1325 8035
rect 1325 8005 1355 8035
rect 1355 8005 1360 8035
rect 1320 8000 1360 8005
rect 1320 7970 1360 7975
rect 1320 7940 1325 7970
rect 1325 7940 1355 7970
rect 1355 7940 1360 7970
rect 1320 7935 1360 7940
rect 1320 7900 1360 7905
rect 1320 7870 1325 7900
rect 1325 7870 1355 7900
rect 1355 7870 1360 7900
rect 1320 7865 1360 7870
rect 1320 7830 1360 7835
rect 1320 7800 1325 7830
rect 1325 7800 1355 7830
rect 1355 7800 1360 7830
rect 1320 7795 1360 7800
rect 1320 7760 1360 7765
rect 1320 7730 1325 7760
rect 1325 7730 1355 7760
rect 1355 7730 1360 7760
rect 1320 7725 1360 7730
rect 1320 7695 1360 7700
rect 1320 7665 1325 7695
rect 1325 7665 1355 7695
rect 1355 7665 1360 7695
rect 1320 7660 1360 7665
rect 1320 7635 1360 7640
rect 1320 7605 1325 7635
rect 1325 7605 1355 7635
rect 1355 7605 1360 7635
rect 1320 7600 1360 7605
rect 1320 7570 1360 7575
rect 1320 7540 1325 7570
rect 1325 7540 1355 7570
rect 1355 7540 1360 7570
rect 1320 7535 1360 7540
rect 1320 7500 1360 7505
rect 1320 7470 1325 7500
rect 1325 7470 1355 7500
rect 1355 7470 1360 7500
rect 1320 7465 1360 7470
rect 1320 7430 1360 7435
rect 1320 7400 1325 7430
rect 1325 7400 1355 7430
rect 1355 7400 1360 7430
rect 1320 7395 1360 7400
rect 1320 7360 1360 7365
rect 1320 7330 1325 7360
rect 1325 7330 1355 7360
rect 1355 7330 1360 7360
rect 1320 7325 1360 7330
rect 1320 7295 1360 7300
rect 1320 7265 1325 7295
rect 1325 7265 1355 7295
rect 1355 7265 1360 7295
rect 1320 7260 1360 7265
rect 1320 7235 1360 7240
rect 1320 7205 1325 7235
rect 1325 7205 1355 7235
rect 1355 7205 1360 7235
rect 1320 7200 1360 7205
rect 1320 7170 1360 7175
rect 1320 7140 1325 7170
rect 1325 7140 1355 7170
rect 1355 7140 1360 7170
rect 1320 7135 1360 7140
rect 1320 7100 1360 7105
rect 1320 7070 1325 7100
rect 1325 7070 1355 7100
rect 1355 7070 1360 7100
rect 1320 7065 1360 7070
rect 1320 7030 1360 7035
rect 1320 7000 1325 7030
rect 1325 7000 1355 7030
rect 1355 7000 1360 7030
rect 1320 6995 1360 7000
rect 1320 6960 1360 6965
rect 1320 6930 1325 6960
rect 1325 6930 1355 6960
rect 1355 6930 1360 6960
rect 1320 6925 1360 6930
rect 1320 6895 1360 6900
rect 1320 6865 1325 6895
rect 1325 6865 1355 6895
rect 1355 6865 1360 6895
rect 1320 6860 1360 6865
rect 1320 6835 1360 6840
rect 1320 6805 1325 6835
rect 1325 6805 1355 6835
rect 1355 6805 1360 6835
rect 1320 6800 1360 6805
rect 1320 6770 1360 6775
rect 1320 6740 1325 6770
rect 1325 6740 1355 6770
rect 1355 6740 1360 6770
rect 1320 6735 1360 6740
rect 1320 6700 1360 6705
rect 1320 6670 1325 6700
rect 1325 6670 1355 6700
rect 1355 6670 1360 6700
rect 1320 6665 1360 6670
rect 1320 6630 1360 6635
rect 1320 6600 1325 6630
rect 1325 6600 1355 6630
rect 1355 6600 1360 6630
rect 1320 6595 1360 6600
rect 1320 6560 1360 6565
rect 1320 6530 1325 6560
rect 1325 6530 1355 6560
rect 1355 6530 1360 6560
rect 1320 6525 1360 6530
rect 1320 6495 1360 6500
rect 1320 6465 1325 6495
rect 1325 6465 1355 6495
rect 1355 6465 1360 6495
rect 1320 6460 1360 6465
rect 1670 9635 1710 9640
rect 1670 9605 1675 9635
rect 1675 9605 1705 9635
rect 1705 9605 1710 9635
rect 1670 9600 1710 9605
rect 1670 9570 1710 9575
rect 1670 9540 1675 9570
rect 1675 9540 1705 9570
rect 1705 9540 1710 9570
rect 1670 9535 1710 9540
rect 1670 9500 1710 9505
rect 1670 9470 1675 9500
rect 1675 9470 1705 9500
rect 1705 9470 1710 9500
rect 1670 9465 1710 9470
rect 1670 9430 1710 9435
rect 1670 9400 1675 9430
rect 1675 9400 1705 9430
rect 1705 9400 1710 9430
rect 1670 9395 1710 9400
rect 1670 9360 1710 9365
rect 1670 9330 1675 9360
rect 1675 9330 1705 9360
rect 1705 9330 1710 9360
rect 1670 9325 1710 9330
rect 1670 9295 1710 9300
rect 1670 9265 1675 9295
rect 1675 9265 1705 9295
rect 1705 9265 1710 9295
rect 1670 9260 1710 9265
rect 1670 9235 1710 9240
rect 1670 9205 1675 9235
rect 1675 9205 1705 9235
rect 1705 9205 1710 9235
rect 1670 9200 1710 9205
rect 1670 9170 1710 9175
rect 1670 9140 1675 9170
rect 1675 9140 1705 9170
rect 1705 9140 1710 9170
rect 1670 9135 1710 9140
rect 1670 9100 1710 9105
rect 1670 9070 1675 9100
rect 1675 9070 1705 9100
rect 1705 9070 1710 9100
rect 1670 9065 1710 9070
rect 1670 9030 1710 9035
rect 1670 9000 1675 9030
rect 1675 9000 1705 9030
rect 1705 9000 1710 9030
rect 1670 8995 1710 9000
rect 1670 8960 1710 8965
rect 1670 8930 1675 8960
rect 1675 8930 1705 8960
rect 1705 8930 1710 8960
rect 1670 8925 1710 8930
rect 1670 8895 1710 8900
rect 1670 8865 1675 8895
rect 1675 8865 1705 8895
rect 1705 8865 1710 8895
rect 1670 8860 1710 8865
rect 1670 8835 1710 8840
rect 1670 8805 1675 8835
rect 1675 8805 1705 8835
rect 1705 8805 1710 8835
rect 1670 8800 1710 8805
rect 1670 8770 1710 8775
rect 1670 8740 1675 8770
rect 1675 8740 1705 8770
rect 1705 8740 1710 8770
rect 1670 8735 1710 8740
rect 1670 8700 1710 8705
rect 1670 8670 1675 8700
rect 1675 8670 1705 8700
rect 1705 8670 1710 8700
rect 1670 8665 1710 8670
rect 1670 8630 1710 8635
rect 1670 8600 1675 8630
rect 1675 8600 1705 8630
rect 1705 8600 1710 8630
rect 1670 8595 1710 8600
rect 1670 8560 1710 8565
rect 1670 8530 1675 8560
rect 1675 8530 1705 8560
rect 1705 8530 1710 8560
rect 1670 8525 1710 8530
rect 1670 8495 1710 8500
rect 1670 8465 1675 8495
rect 1675 8465 1705 8495
rect 1705 8465 1710 8495
rect 1670 8460 1710 8465
rect 1670 8435 1710 8440
rect 1670 8405 1675 8435
rect 1675 8405 1705 8435
rect 1705 8405 1710 8435
rect 1670 8400 1710 8405
rect 1670 8370 1710 8375
rect 1670 8340 1675 8370
rect 1675 8340 1705 8370
rect 1705 8340 1710 8370
rect 1670 8335 1710 8340
rect 1670 8300 1710 8305
rect 1670 8270 1675 8300
rect 1675 8270 1705 8300
rect 1705 8270 1710 8300
rect 1670 8265 1710 8270
rect 1670 8230 1710 8235
rect 1670 8200 1675 8230
rect 1675 8200 1705 8230
rect 1705 8200 1710 8230
rect 1670 8195 1710 8200
rect 1670 8160 1710 8165
rect 1670 8130 1675 8160
rect 1675 8130 1705 8160
rect 1705 8130 1710 8160
rect 1670 8125 1710 8130
rect 1670 8095 1710 8100
rect 1670 8065 1675 8095
rect 1675 8065 1705 8095
rect 1705 8065 1710 8095
rect 1670 8060 1710 8065
rect 1670 8035 1710 8040
rect 1670 8005 1675 8035
rect 1675 8005 1705 8035
rect 1705 8005 1710 8035
rect 1670 8000 1710 8005
rect 1670 7970 1710 7975
rect 1670 7940 1675 7970
rect 1675 7940 1705 7970
rect 1705 7940 1710 7970
rect 1670 7935 1710 7940
rect 1670 7900 1710 7905
rect 1670 7870 1675 7900
rect 1675 7870 1705 7900
rect 1705 7870 1710 7900
rect 1670 7865 1710 7870
rect 1670 7830 1710 7835
rect 1670 7800 1675 7830
rect 1675 7800 1705 7830
rect 1705 7800 1710 7830
rect 1670 7795 1710 7800
rect 1670 7760 1710 7765
rect 1670 7730 1675 7760
rect 1675 7730 1705 7760
rect 1705 7730 1710 7760
rect 1670 7725 1710 7730
rect 1670 7695 1710 7700
rect 1670 7665 1675 7695
rect 1675 7665 1705 7695
rect 1705 7665 1710 7695
rect 1670 7660 1710 7665
rect 1670 7635 1710 7640
rect 1670 7605 1675 7635
rect 1675 7605 1705 7635
rect 1705 7605 1710 7635
rect 1670 7600 1710 7605
rect 1670 7570 1710 7575
rect 1670 7540 1675 7570
rect 1675 7540 1705 7570
rect 1705 7540 1710 7570
rect 1670 7535 1710 7540
rect 1670 7500 1710 7505
rect 1670 7470 1675 7500
rect 1675 7470 1705 7500
rect 1705 7470 1710 7500
rect 1670 7465 1710 7470
rect 1670 7430 1710 7435
rect 1670 7400 1675 7430
rect 1675 7400 1705 7430
rect 1705 7400 1710 7430
rect 1670 7395 1710 7400
rect 1670 7360 1710 7365
rect 1670 7330 1675 7360
rect 1675 7330 1705 7360
rect 1705 7330 1710 7360
rect 1670 7325 1710 7330
rect 1670 7295 1710 7300
rect 1670 7265 1675 7295
rect 1675 7265 1705 7295
rect 1705 7265 1710 7295
rect 1670 7260 1710 7265
rect 1670 7235 1710 7240
rect 1670 7205 1675 7235
rect 1675 7205 1705 7235
rect 1705 7205 1710 7235
rect 1670 7200 1710 7205
rect 1670 7170 1710 7175
rect 1670 7140 1675 7170
rect 1675 7140 1705 7170
rect 1705 7140 1710 7170
rect 1670 7135 1710 7140
rect 1670 7100 1710 7105
rect 1670 7070 1675 7100
rect 1675 7070 1705 7100
rect 1705 7070 1710 7100
rect 1670 7065 1710 7070
rect 1670 7030 1710 7035
rect 1670 7000 1675 7030
rect 1675 7000 1705 7030
rect 1705 7000 1710 7030
rect 1670 6995 1710 7000
rect 1670 6960 1710 6965
rect 1670 6930 1675 6960
rect 1675 6930 1705 6960
rect 1705 6930 1710 6960
rect 1670 6925 1710 6930
rect 1670 6895 1710 6900
rect 1670 6865 1675 6895
rect 1675 6865 1705 6895
rect 1705 6865 1710 6895
rect 1670 6860 1710 6865
rect 1670 6835 1710 6840
rect 1670 6805 1675 6835
rect 1675 6805 1705 6835
rect 1705 6805 1710 6835
rect 1670 6800 1710 6805
rect 1670 6770 1710 6775
rect 1670 6740 1675 6770
rect 1675 6740 1705 6770
rect 1705 6740 1710 6770
rect 1670 6735 1710 6740
rect 1670 6700 1710 6705
rect 1670 6670 1675 6700
rect 1675 6670 1705 6700
rect 1705 6670 1710 6700
rect 1670 6665 1710 6670
rect 1670 6630 1710 6635
rect 1670 6600 1675 6630
rect 1675 6600 1705 6630
rect 1705 6600 1710 6630
rect 1670 6595 1710 6600
rect 1670 6560 1710 6565
rect 1670 6530 1675 6560
rect 1675 6530 1705 6560
rect 1705 6530 1710 6560
rect 1670 6525 1710 6530
rect 1670 6495 1710 6500
rect 1670 6465 1675 6495
rect 1675 6465 1705 6495
rect 1705 6465 1710 6495
rect 1670 6460 1710 6465
rect 2385 9635 2425 9640
rect 2385 9605 2390 9635
rect 2390 9605 2420 9635
rect 2420 9605 2425 9635
rect 2385 9600 2425 9605
rect 2385 9570 2425 9575
rect 2385 9540 2390 9570
rect 2390 9540 2420 9570
rect 2420 9540 2425 9570
rect 2385 9535 2425 9540
rect 2385 9500 2425 9505
rect 2385 9470 2390 9500
rect 2390 9470 2420 9500
rect 2420 9470 2425 9500
rect 2385 9465 2425 9470
rect 2385 9430 2425 9435
rect 2385 9400 2390 9430
rect 2390 9400 2420 9430
rect 2420 9400 2425 9430
rect 2385 9395 2425 9400
rect 2385 9360 2425 9365
rect 2385 9330 2390 9360
rect 2390 9330 2420 9360
rect 2420 9330 2425 9360
rect 2385 9325 2425 9330
rect 2385 9295 2425 9300
rect 2385 9265 2390 9295
rect 2390 9265 2420 9295
rect 2420 9265 2425 9295
rect 2385 9260 2425 9265
rect 2385 9235 2425 9240
rect 2385 9205 2390 9235
rect 2390 9205 2420 9235
rect 2420 9205 2425 9235
rect 2385 9200 2425 9205
rect 2385 9170 2425 9175
rect 2385 9140 2390 9170
rect 2390 9140 2420 9170
rect 2420 9140 2425 9170
rect 2385 9135 2425 9140
rect 2385 9100 2425 9105
rect 2385 9070 2390 9100
rect 2390 9070 2420 9100
rect 2420 9070 2425 9100
rect 2385 9065 2425 9070
rect 2385 9030 2425 9035
rect 2385 9000 2390 9030
rect 2390 9000 2420 9030
rect 2420 9000 2425 9030
rect 2385 8995 2425 9000
rect 2385 8960 2425 8965
rect 2385 8930 2390 8960
rect 2390 8930 2420 8960
rect 2420 8930 2425 8960
rect 2385 8925 2425 8930
rect 2385 8895 2425 8900
rect 2385 8865 2390 8895
rect 2390 8865 2420 8895
rect 2420 8865 2425 8895
rect 2385 8860 2425 8865
rect 2385 8835 2425 8840
rect 2385 8805 2390 8835
rect 2390 8805 2420 8835
rect 2420 8805 2425 8835
rect 2385 8800 2425 8805
rect 2385 8770 2425 8775
rect 2385 8740 2390 8770
rect 2390 8740 2420 8770
rect 2420 8740 2425 8770
rect 2385 8735 2425 8740
rect 2385 8700 2425 8705
rect 2385 8670 2390 8700
rect 2390 8670 2420 8700
rect 2420 8670 2425 8700
rect 2385 8665 2425 8670
rect 2385 8630 2425 8635
rect 2385 8600 2390 8630
rect 2390 8600 2420 8630
rect 2420 8600 2425 8630
rect 2385 8595 2425 8600
rect 2385 8560 2425 8565
rect 2385 8530 2390 8560
rect 2390 8530 2420 8560
rect 2420 8530 2425 8560
rect 2385 8525 2425 8530
rect 2385 8495 2425 8500
rect 2385 8465 2390 8495
rect 2390 8465 2420 8495
rect 2420 8465 2425 8495
rect 2385 8460 2425 8465
rect 2385 8435 2425 8440
rect 2385 8405 2390 8435
rect 2390 8405 2420 8435
rect 2420 8405 2425 8435
rect 2385 8400 2425 8405
rect 2385 8370 2425 8375
rect 2385 8340 2390 8370
rect 2390 8340 2420 8370
rect 2420 8340 2425 8370
rect 2385 8335 2425 8340
rect 2385 8300 2425 8305
rect 2385 8270 2390 8300
rect 2390 8270 2420 8300
rect 2420 8270 2425 8300
rect 2385 8265 2425 8270
rect 2385 8230 2425 8235
rect 2385 8200 2390 8230
rect 2390 8200 2420 8230
rect 2420 8200 2425 8230
rect 2385 8195 2425 8200
rect 2385 8160 2425 8165
rect 2385 8130 2390 8160
rect 2390 8130 2420 8160
rect 2420 8130 2425 8160
rect 2385 8125 2425 8130
rect 2385 8095 2425 8100
rect 2385 8065 2390 8095
rect 2390 8065 2420 8095
rect 2420 8065 2425 8095
rect 2385 8060 2425 8065
rect 2385 8035 2425 8040
rect 2385 8005 2390 8035
rect 2390 8005 2420 8035
rect 2420 8005 2425 8035
rect 2385 8000 2425 8005
rect 2385 7970 2425 7975
rect 2385 7940 2390 7970
rect 2390 7940 2420 7970
rect 2420 7940 2425 7970
rect 2385 7935 2425 7940
rect 2385 7900 2425 7905
rect 2385 7870 2390 7900
rect 2390 7870 2420 7900
rect 2420 7870 2425 7900
rect 2385 7865 2425 7870
rect 2385 7830 2425 7835
rect 2385 7800 2390 7830
rect 2390 7800 2420 7830
rect 2420 7800 2425 7830
rect 2385 7795 2425 7800
rect 2385 7760 2425 7765
rect 2385 7730 2390 7760
rect 2390 7730 2420 7760
rect 2420 7730 2425 7760
rect 2385 7725 2425 7730
rect 2385 7695 2425 7700
rect 2385 7665 2390 7695
rect 2390 7665 2420 7695
rect 2420 7665 2425 7695
rect 2385 7660 2425 7665
rect 2385 7635 2425 7640
rect 2385 7605 2390 7635
rect 2390 7605 2420 7635
rect 2420 7605 2425 7635
rect 2385 7600 2425 7605
rect 2385 7570 2425 7575
rect 2385 7540 2390 7570
rect 2390 7540 2420 7570
rect 2420 7540 2425 7570
rect 2385 7535 2425 7540
rect 2385 7500 2425 7505
rect 2385 7470 2390 7500
rect 2390 7470 2420 7500
rect 2420 7470 2425 7500
rect 2385 7465 2425 7470
rect 2385 7430 2425 7435
rect 2385 7400 2390 7430
rect 2390 7400 2420 7430
rect 2420 7400 2425 7430
rect 2385 7395 2425 7400
rect 2385 7360 2425 7365
rect 2385 7330 2390 7360
rect 2390 7330 2420 7360
rect 2420 7330 2425 7360
rect 2385 7325 2425 7330
rect 2385 7295 2425 7300
rect 2385 7265 2390 7295
rect 2390 7265 2420 7295
rect 2420 7265 2425 7295
rect 2385 7260 2425 7265
rect 2385 7235 2425 7240
rect 2385 7205 2390 7235
rect 2390 7205 2420 7235
rect 2420 7205 2425 7235
rect 2385 7200 2425 7205
rect 2385 7170 2425 7175
rect 2385 7140 2390 7170
rect 2390 7140 2420 7170
rect 2420 7140 2425 7170
rect 2385 7135 2425 7140
rect 2385 7100 2425 7105
rect 2385 7070 2390 7100
rect 2390 7070 2420 7100
rect 2420 7070 2425 7100
rect 2385 7065 2425 7070
rect 2385 7030 2425 7035
rect 2385 7000 2390 7030
rect 2390 7000 2420 7030
rect 2420 7000 2425 7030
rect 2385 6995 2425 7000
rect 2385 6960 2425 6965
rect 2385 6930 2390 6960
rect 2390 6930 2420 6960
rect 2420 6930 2425 6960
rect 2385 6925 2425 6930
rect 2385 6895 2425 6900
rect 2385 6865 2390 6895
rect 2390 6865 2420 6895
rect 2420 6865 2425 6895
rect 2385 6860 2425 6865
rect 2385 6835 2425 6840
rect 2385 6805 2390 6835
rect 2390 6805 2420 6835
rect 2420 6805 2425 6835
rect 2385 6800 2425 6805
rect 2385 6770 2425 6775
rect 2385 6740 2390 6770
rect 2390 6740 2420 6770
rect 2420 6740 2425 6770
rect 2385 6735 2425 6740
rect 2385 6700 2425 6705
rect 2385 6670 2390 6700
rect 2390 6670 2420 6700
rect 2420 6670 2425 6700
rect 2385 6665 2425 6670
rect 2385 6630 2425 6635
rect 2385 6600 2390 6630
rect 2390 6600 2420 6630
rect 2420 6600 2425 6630
rect 2385 6595 2425 6600
rect 2385 6560 2425 6565
rect 2385 6530 2390 6560
rect 2390 6530 2420 6560
rect 2420 6530 2425 6560
rect 2385 6525 2425 6530
rect 2385 6495 2425 6500
rect 2385 6465 2390 6495
rect 2390 6465 2420 6495
rect 2420 6465 2425 6495
rect 2385 6460 2425 6465
rect 3235 9635 3275 9640
rect 3235 9605 3240 9635
rect 3240 9605 3270 9635
rect 3270 9605 3275 9635
rect 3235 9600 3275 9605
rect 3235 9570 3275 9575
rect 3235 9540 3240 9570
rect 3240 9540 3270 9570
rect 3270 9540 3275 9570
rect 3235 9535 3275 9540
rect 3235 9500 3275 9505
rect 3235 9470 3240 9500
rect 3240 9470 3270 9500
rect 3270 9470 3275 9500
rect 3235 9465 3275 9470
rect 3235 9430 3275 9435
rect 3235 9400 3240 9430
rect 3240 9400 3270 9430
rect 3270 9400 3275 9430
rect 3235 9395 3275 9400
rect 3235 9360 3275 9365
rect 3235 9330 3240 9360
rect 3240 9330 3270 9360
rect 3270 9330 3275 9360
rect 3235 9325 3275 9330
rect 3235 9295 3275 9300
rect 3235 9265 3240 9295
rect 3240 9265 3270 9295
rect 3270 9265 3275 9295
rect 3235 9260 3275 9265
rect 3235 9235 3275 9240
rect 3235 9205 3240 9235
rect 3240 9205 3270 9235
rect 3270 9205 3275 9235
rect 3235 9200 3275 9205
rect 3235 9170 3275 9175
rect 3235 9140 3240 9170
rect 3240 9140 3270 9170
rect 3270 9140 3275 9170
rect 3235 9135 3275 9140
rect 3235 9100 3275 9105
rect 3235 9070 3240 9100
rect 3240 9070 3270 9100
rect 3270 9070 3275 9100
rect 3235 9065 3275 9070
rect 3235 9030 3275 9035
rect 3235 9000 3240 9030
rect 3240 9000 3270 9030
rect 3270 9000 3275 9030
rect 3235 8995 3275 9000
rect 3235 8960 3275 8965
rect 3235 8930 3240 8960
rect 3240 8930 3270 8960
rect 3270 8930 3275 8960
rect 3235 8925 3275 8930
rect 3235 8895 3275 8900
rect 3235 8865 3240 8895
rect 3240 8865 3270 8895
rect 3270 8865 3275 8895
rect 3235 8860 3275 8865
rect 3235 8835 3275 8840
rect 3235 8805 3240 8835
rect 3240 8805 3270 8835
rect 3270 8805 3275 8835
rect 3235 8800 3275 8805
rect 3235 8770 3275 8775
rect 3235 8740 3240 8770
rect 3240 8740 3270 8770
rect 3270 8740 3275 8770
rect 3235 8735 3275 8740
rect 3235 8700 3275 8705
rect 3235 8670 3240 8700
rect 3240 8670 3270 8700
rect 3270 8670 3275 8700
rect 3235 8665 3275 8670
rect 3235 8630 3275 8635
rect 3235 8600 3240 8630
rect 3240 8600 3270 8630
rect 3270 8600 3275 8630
rect 3235 8595 3275 8600
rect 3235 8560 3275 8565
rect 3235 8530 3240 8560
rect 3240 8530 3270 8560
rect 3270 8530 3275 8560
rect 3235 8525 3275 8530
rect 3235 8495 3275 8500
rect 3235 8465 3240 8495
rect 3240 8465 3270 8495
rect 3270 8465 3275 8495
rect 3235 8460 3275 8465
rect 3235 8435 3275 8440
rect 3235 8405 3240 8435
rect 3240 8405 3270 8435
rect 3270 8405 3275 8435
rect 3235 8400 3275 8405
rect 3235 8370 3275 8375
rect 3235 8340 3240 8370
rect 3240 8340 3270 8370
rect 3270 8340 3275 8370
rect 3235 8335 3275 8340
rect 3235 8300 3275 8305
rect 3235 8270 3240 8300
rect 3240 8270 3270 8300
rect 3270 8270 3275 8300
rect 3235 8265 3275 8270
rect 3235 8230 3275 8235
rect 3235 8200 3240 8230
rect 3240 8200 3270 8230
rect 3270 8200 3275 8230
rect 3235 8195 3275 8200
rect 3235 8160 3275 8165
rect 3235 8130 3240 8160
rect 3240 8130 3270 8160
rect 3270 8130 3275 8160
rect 3235 8125 3275 8130
rect 3235 8095 3275 8100
rect 3235 8065 3240 8095
rect 3240 8065 3270 8095
rect 3270 8065 3275 8095
rect 3235 8060 3275 8065
rect 3235 8035 3275 8040
rect 3235 8005 3240 8035
rect 3240 8005 3270 8035
rect 3270 8005 3275 8035
rect 3235 8000 3275 8005
rect 3235 7970 3275 7975
rect 3235 7940 3240 7970
rect 3240 7940 3270 7970
rect 3270 7940 3275 7970
rect 3235 7935 3275 7940
rect 3235 7900 3275 7905
rect 3235 7870 3240 7900
rect 3240 7870 3270 7900
rect 3270 7870 3275 7900
rect 3235 7865 3275 7870
rect 3235 7830 3275 7835
rect 3235 7800 3240 7830
rect 3240 7800 3270 7830
rect 3270 7800 3275 7830
rect 3235 7795 3275 7800
rect 3235 7760 3275 7765
rect 3235 7730 3240 7760
rect 3240 7730 3270 7760
rect 3270 7730 3275 7760
rect 3235 7725 3275 7730
rect 3235 7695 3275 7700
rect 3235 7665 3240 7695
rect 3240 7665 3270 7695
rect 3270 7665 3275 7695
rect 3235 7660 3275 7665
rect 3235 7635 3275 7640
rect 3235 7605 3240 7635
rect 3240 7605 3270 7635
rect 3270 7605 3275 7635
rect 3235 7600 3275 7605
rect 3235 7570 3275 7575
rect 3235 7540 3240 7570
rect 3240 7540 3270 7570
rect 3270 7540 3275 7570
rect 3235 7535 3275 7540
rect 3235 7500 3275 7505
rect 3235 7470 3240 7500
rect 3240 7470 3270 7500
rect 3270 7470 3275 7500
rect 3235 7465 3275 7470
rect 3235 7430 3275 7435
rect 3235 7400 3240 7430
rect 3240 7400 3270 7430
rect 3270 7400 3275 7430
rect 3235 7395 3275 7400
rect 3235 7360 3275 7365
rect 3235 7330 3240 7360
rect 3240 7330 3270 7360
rect 3270 7330 3275 7360
rect 3235 7325 3275 7330
rect 3235 7295 3275 7300
rect 3235 7265 3240 7295
rect 3240 7265 3270 7295
rect 3270 7265 3275 7295
rect 3235 7260 3275 7265
rect 3235 7235 3275 7240
rect 3235 7205 3240 7235
rect 3240 7205 3270 7235
rect 3270 7205 3275 7235
rect 3235 7200 3275 7205
rect 3235 7170 3275 7175
rect 3235 7140 3240 7170
rect 3240 7140 3270 7170
rect 3270 7140 3275 7170
rect 3235 7135 3275 7140
rect 3235 7100 3275 7105
rect 3235 7070 3240 7100
rect 3240 7070 3270 7100
rect 3270 7070 3275 7100
rect 3235 7065 3275 7070
rect 3235 7030 3275 7035
rect 3235 7000 3240 7030
rect 3240 7000 3270 7030
rect 3270 7000 3275 7030
rect 3235 6995 3275 7000
rect 3235 6960 3275 6965
rect 3235 6930 3240 6960
rect 3240 6930 3270 6960
rect 3270 6930 3275 6960
rect 3235 6925 3275 6930
rect 3235 6895 3275 6900
rect 3235 6865 3240 6895
rect 3240 6865 3270 6895
rect 3270 6865 3275 6895
rect 3235 6860 3275 6865
rect 3235 6835 3275 6840
rect 3235 6805 3240 6835
rect 3240 6805 3270 6835
rect 3270 6805 3275 6835
rect 3235 6800 3275 6805
rect 3235 6770 3275 6775
rect 3235 6740 3240 6770
rect 3240 6740 3270 6770
rect 3270 6740 3275 6770
rect 3235 6735 3275 6740
rect 3235 6700 3275 6705
rect 3235 6670 3240 6700
rect 3240 6670 3270 6700
rect 3270 6670 3275 6700
rect 3235 6665 3275 6670
rect 3235 6630 3275 6635
rect 3235 6600 3240 6630
rect 3240 6600 3270 6630
rect 3270 6600 3275 6630
rect 3235 6595 3275 6600
rect 3235 6560 3275 6565
rect 3235 6530 3240 6560
rect 3240 6530 3270 6560
rect 3270 6530 3275 6560
rect 3235 6525 3275 6530
rect 3235 6495 3275 6500
rect 3235 6465 3240 6495
rect 3240 6465 3270 6495
rect 3270 6465 3275 6495
rect 3235 6460 3275 6465
rect 5645 9635 5685 9640
rect 5645 9605 5650 9635
rect 5650 9605 5680 9635
rect 5680 9605 5685 9635
rect 5645 9600 5685 9605
rect 5645 9570 5685 9575
rect 5645 9540 5650 9570
rect 5650 9540 5680 9570
rect 5680 9540 5685 9570
rect 5645 9535 5685 9540
rect 5645 9500 5685 9505
rect 5645 9470 5650 9500
rect 5650 9470 5680 9500
rect 5680 9470 5685 9500
rect 5645 9465 5685 9470
rect 5645 9430 5685 9435
rect 5645 9400 5650 9430
rect 5650 9400 5680 9430
rect 5680 9400 5685 9430
rect 5645 9395 5685 9400
rect 5645 9360 5685 9365
rect 5645 9330 5650 9360
rect 5650 9330 5680 9360
rect 5680 9330 5685 9360
rect 5645 9325 5685 9330
rect 5645 9295 5685 9300
rect 5645 9265 5650 9295
rect 5650 9265 5680 9295
rect 5680 9265 5685 9295
rect 5645 9260 5685 9265
rect 5645 9235 5685 9240
rect 5645 9205 5650 9235
rect 5650 9205 5680 9235
rect 5680 9205 5685 9235
rect 5645 9200 5685 9205
rect 5645 9170 5685 9175
rect 5645 9140 5650 9170
rect 5650 9140 5680 9170
rect 5680 9140 5685 9170
rect 5645 9135 5685 9140
rect 5645 9100 5685 9105
rect 5645 9070 5650 9100
rect 5650 9070 5680 9100
rect 5680 9070 5685 9100
rect 5645 9065 5685 9070
rect 5645 9030 5685 9035
rect 5645 9000 5650 9030
rect 5650 9000 5680 9030
rect 5680 9000 5685 9030
rect 5645 8995 5685 9000
rect 5645 8960 5685 8965
rect 5645 8930 5650 8960
rect 5650 8930 5680 8960
rect 5680 8930 5685 8960
rect 5645 8925 5685 8930
rect 5645 8895 5685 8900
rect 5645 8865 5650 8895
rect 5650 8865 5680 8895
rect 5680 8865 5685 8895
rect 5645 8860 5685 8865
rect 5645 8835 5685 8840
rect 5645 8805 5650 8835
rect 5650 8805 5680 8835
rect 5680 8805 5685 8835
rect 5645 8800 5685 8805
rect 5645 8770 5685 8775
rect 5645 8740 5650 8770
rect 5650 8740 5680 8770
rect 5680 8740 5685 8770
rect 5645 8735 5685 8740
rect 5645 8700 5685 8705
rect 5645 8670 5650 8700
rect 5650 8670 5680 8700
rect 5680 8670 5685 8700
rect 5645 8665 5685 8670
rect 5645 8630 5685 8635
rect 5645 8600 5650 8630
rect 5650 8600 5680 8630
rect 5680 8600 5685 8630
rect 5645 8595 5685 8600
rect 5645 8560 5685 8565
rect 5645 8530 5650 8560
rect 5650 8530 5680 8560
rect 5680 8530 5685 8560
rect 5645 8525 5685 8530
rect 5645 8495 5685 8500
rect 5645 8465 5650 8495
rect 5650 8465 5680 8495
rect 5680 8465 5685 8495
rect 5645 8460 5685 8465
rect 5645 8435 5685 8440
rect 5645 8405 5650 8435
rect 5650 8405 5680 8435
rect 5680 8405 5685 8435
rect 5645 8400 5685 8405
rect 5645 8370 5685 8375
rect 5645 8340 5650 8370
rect 5650 8340 5680 8370
rect 5680 8340 5685 8370
rect 5645 8335 5685 8340
rect 5645 8300 5685 8305
rect 5645 8270 5650 8300
rect 5650 8270 5680 8300
rect 5680 8270 5685 8300
rect 5645 8265 5685 8270
rect 5645 8230 5685 8235
rect 5645 8200 5650 8230
rect 5650 8200 5680 8230
rect 5680 8200 5685 8230
rect 5645 8195 5685 8200
rect 5645 8160 5685 8165
rect 5645 8130 5650 8160
rect 5650 8130 5680 8160
rect 5680 8130 5685 8160
rect 5645 8125 5685 8130
rect 5645 8095 5685 8100
rect 5645 8065 5650 8095
rect 5650 8065 5680 8095
rect 5680 8065 5685 8095
rect 5645 8060 5685 8065
rect 5645 8035 5685 8040
rect 5645 8005 5650 8035
rect 5650 8005 5680 8035
rect 5680 8005 5685 8035
rect 5645 8000 5685 8005
rect 5645 7970 5685 7975
rect 5645 7940 5650 7970
rect 5650 7940 5680 7970
rect 5680 7940 5685 7970
rect 5645 7935 5685 7940
rect 5645 7900 5685 7905
rect 5645 7870 5650 7900
rect 5650 7870 5680 7900
rect 5680 7870 5685 7900
rect 5645 7865 5685 7870
rect 5645 7830 5685 7835
rect 5645 7800 5650 7830
rect 5650 7800 5680 7830
rect 5680 7800 5685 7830
rect 5645 7795 5685 7800
rect 5645 7760 5685 7765
rect 5645 7730 5650 7760
rect 5650 7730 5680 7760
rect 5680 7730 5685 7760
rect 5645 7725 5685 7730
rect 5645 7695 5685 7700
rect 5645 7665 5650 7695
rect 5650 7665 5680 7695
rect 5680 7665 5685 7695
rect 5645 7660 5685 7665
rect 5645 7635 5685 7640
rect 5645 7605 5650 7635
rect 5650 7605 5680 7635
rect 5680 7605 5685 7635
rect 5645 7600 5685 7605
rect 5645 7570 5685 7575
rect 5645 7540 5650 7570
rect 5650 7540 5680 7570
rect 5680 7540 5685 7570
rect 5645 7535 5685 7540
rect 5645 7500 5685 7505
rect 5645 7470 5650 7500
rect 5650 7470 5680 7500
rect 5680 7470 5685 7500
rect 5645 7465 5685 7470
rect 5645 7430 5685 7435
rect 5645 7400 5650 7430
rect 5650 7400 5680 7430
rect 5680 7400 5685 7430
rect 5645 7395 5685 7400
rect 5645 7360 5685 7365
rect 5645 7330 5650 7360
rect 5650 7330 5680 7360
rect 5680 7330 5685 7360
rect 5645 7325 5685 7330
rect 5645 7295 5685 7300
rect 5645 7265 5650 7295
rect 5650 7265 5680 7295
rect 5680 7265 5685 7295
rect 5645 7260 5685 7265
rect 5645 7235 5685 7240
rect 5645 7205 5650 7235
rect 5650 7205 5680 7235
rect 5680 7205 5685 7235
rect 5645 7200 5685 7205
rect 5645 7170 5685 7175
rect 5645 7140 5650 7170
rect 5650 7140 5680 7170
rect 5680 7140 5685 7170
rect 5645 7135 5685 7140
rect 5645 7100 5685 7105
rect 5645 7070 5650 7100
rect 5650 7070 5680 7100
rect 5680 7070 5685 7100
rect 5645 7065 5685 7070
rect 5645 7030 5685 7035
rect 5645 7000 5650 7030
rect 5650 7000 5680 7030
rect 5680 7000 5685 7030
rect 5645 6995 5685 7000
rect 5645 6960 5685 6965
rect 5645 6930 5650 6960
rect 5650 6930 5680 6960
rect 5680 6930 5685 6960
rect 5645 6925 5685 6930
rect 5645 6895 5685 6900
rect 5645 6865 5650 6895
rect 5650 6865 5680 6895
rect 5680 6865 5685 6895
rect 5645 6860 5685 6865
rect 5645 6835 5685 6840
rect 5645 6805 5650 6835
rect 5650 6805 5680 6835
rect 5680 6805 5685 6835
rect 5645 6800 5685 6805
rect 5645 6770 5685 6775
rect 5645 6740 5650 6770
rect 5650 6740 5680 6770
rect 5680 6740 5685 6770
rect 5645 6735 5685 6740
rect 5645 6700 5685 6705
rect 5645 6670 5650 6700
rect 5650 6670 5680 6700
rect 5680 6670 5685 6700
rect 5645 6665 5685 6670
rect 5645 6630 5685 6635
rect 5645 6600 5650 6630
rect 5650 6600 5680 6630
rect 5680 6600 5685 6630
rect 5645 6595 5685 6600
rect 5645 6560 5685 6565
rect 5645 6530 5650 6560
rect 5650 6530 5680 6560
rect 5680 6530 5685 6560
rect 5645 6525 5685 6530
rect 5645 6495 5685 6500
rect 5645 6465 5650 6495
rect 5650 6465 5680 6495
rect 5680 6465 5685 6495
rect 5645 6460 5685 6465
rect 6300 9635 6340 9640
rect 6300 9605 6305 9635
rect 6305 9605 6335 9635
rect 6335 9605 6340 9635
rect 6300 9600 6340 9605
rect 6300 9570 6340 9575
rect 6300 9540 6305 9570
rect 6305 9540 6335 9570
rect 6335 9540 6340 9570
rect 6300 9535 6340 9540
rect 6300 9500 6340 9505
rect 6300 9470 6305 9500
rect 6305 9470 6335 9500
rect 6335 9470 6340 9500
rect 6300 9465 6340 9470
rect 6300 9430 6340 9435
rect 6300 9400 6305 9430
rect 6305 9400 6335 9430
rect 6335 9400 6340 9430
rect 6300 9395 6340 9400
rect 6300 9360 6340 9365
rect 6300 9330 6305 9360
rect 6305 9330 6335 9360
rect 6335 9330 6340 9360
rect 6300 9325 6340 9330
rect 6300 9295 6340 9300
rect 6300 9265 6305 9295
rect 6305 9265 6335 9295
rect 6335 9265 6340 9295
rect 6300 9260 6340 9265
rect 6300 9235 6340 9240
rect 6300 9205 6305 9235
rect 6305 9205 6335 9235
rect 6335 9205 6340 9235
rect 6300 9200 6340 9205
rect 6300 9170 6340 9175
rect 6300 9140 6305 9170
rect 6305 9140 6335 9170
rect 6335 9140 6340 9170
rect 6300 9135 6340 9140
rect 6300 9100 6340 9105
rect 6300 9070 6305 9100
rect 6305 9070 6335 9100
rect 6335 9070 6340 9100
rect 6300 9065 6340 9070
rect 6300 9030 6340 9035
rect 6300 9000 6305 9030
rect 6305 9000 6335 9030
rect 6335 9000 6340 9030
rect 6300 8995 6340 9000
rect 6300 8960 6340 8965
rect 6300 8930 6305 8960
rect 6305 8930 6335 8960
rect 6335 8930 6340 8960
rect 6300 8925 6340 8930
rect 6300 8895 6340 8900
rect 6300 8865 6305 8895
rect 6305 8865 6335 8895
rect 6335 8865 6340 8895
rect 6300 8860 6340 8865
rect 6300 8835 6340 8840
rect 6300 8805 6305 8835
rect 6305 8805 6335 8835
rect 6335 8805 6340 8835
rect 6300 8800 6340 8805
rect 6300 8770 6340 8775
rect 6300 8740 6305 8770
rect 6305 8740 6335 8770
rect 6335 8740 6340 8770
rect 6300 8735 6340 8740
rect 6300 8700 6340 8705
rect 6300 8670 6305 8700
rect 6305 8670 6335 8700
rect 6335 8670 6340 8700
rect 6300 8665 6340 8670
rect 6300 8630 6340 8635
rect 6300 8600 6305 8630
rect 6305 8600 6335 8630
rect 6335 8600 6340 8630
rect 6300 8595 6340 8600
rect 6300 8560 6340 8565
rect 6300 8530 6305 8560
rect 6305 8530 6335 8560
rect 6335 8530 6340 8560
rect 6300 8525 6340 8530
rect 6300 8495 6340 8500
rect 6300 8465 6305 8495
rect 6305 8465 6335 8495
rect 6335 8465 6340 8495
rect 6300 8460 6340 8465
rect 6300 8435 6340 8440
rect 6300 8405 6305 8435
rect 6305 8405 6335 8435
rect 6335 8405 6340 8435
rect 6300 8400 6340 8405
rect 6300 8370 6340 8375
rect 6300 8340 6305 8370
rect 6305 8340 6335 8370
rect 6335 8340 6340 8370
rect 6300 8335 6340 8340
rect 6300 8300 6340 8305
rect 6300 8270 6305 8300
rect 6305 8270 6335 8300
rect 6335 8270 6340 8300
rect 6300 8265 6340 8270
rect 6300 8230 6340 8235
rect 6300 8200 6305 8230
rect 6305 8200 6335 8230
rect 6335 8200 6340 8230
rect 6300 8195 6340 8200
rect 6300 8160 6340 8165
rect 6300 8130 6305 8160
rect 6305 8130 6335 8160
rect 6335 8130 6340 8160
rect 6300 8125 6340 8130
rect 6300 8095 6340 8100
rect 6300 8065 6305 8095
rect 6305 8065 6335 8095
rect 6335 8065 6340 8095
rect 6300 8060 6340 8065
rect 6300 8035 6340 8040
rect 6300 8005 6305 8035
rect 6305 8005 6335 8035
rect 6335 8005 6340 8035
rect 6300 8000 6340 8005
rect 6300 7970 6340 7975
rect 6300 7940 6305 7970
rect 6305 7940 6335 7970
rect 6335 7940 6340 7970
rect 6300 7935 6340 7940
rect 6300 7900 6340 7905
rect 6300 7870 6305 7900
rect 6305 7870 6335 7900
rect 6335 7870 6340 7900
rect 6300 7865 6340 7870
rect 6300 7830 6340 7835
rect 6300 7800 6305 7830
rect 6305 7800 6335 7830
rect 6335 7800 6340 7830
rect 6300 7795 6340 7800
rect 6300 7760 6340 7765
rect 6300 7730 6305 7760
rect 6305 7730 6335 7760
rect 6335 7730 6340 7760
rect 6300 7725 6340 7730
rect 6300 7695 6340 7700
rect 6300 7665 6305 7695
rect 6305 7665 6335 7695
rect 6335 7665 6340 7695
rect 6300 7660 6340 7665
rect 6300 7635 6340 7640
rect 6300 7605 6305 7635
rect 6305 7605 6335 7635
rect 6335 7605 6340 7635
rect 6300 7600 6340 7605
rect 6300 7570 6340 7575
rect 6300 7540 6305 7570
rect 6305 7540 6335 7570
rect 6335 7540 6340 7570
rect 6300 7535 6340 7540
rect 6300 7500 6340 7505
rect 6300 7470 6305 7500
rect 6305 7470 6335 7500
rect 6335 7470 6340 7500
rect 6300 7465 6340 7470
rect 6300 7430 6340 7435
rect 6300 7400 6305 7430
rect 6305 7400 6335 7430
rect 6335 7400 6340 7430
rect 6300 7395 6340 7400
rect 6300 7360 6340 7365
rect 6300 7330 6305 7360
rect 6305 7330 6335 7360
rect 6335 7330 6340 7360
rect 6300 7325 6340 7330
rect 6300 7295 6340 7300
rect 6300 7265 6305 7295
rect 6305 7265 6335 7295
rect 6335 7265 6340 7295
rect 6300 7260 6340 7265
rect 6300 7235 6340 7240
rect 6300 7205 6305 7235
rect 6305 7205 6335 7235
rect 6335 7205 6340 7235
rect 6300 7200 6340 7205
rect 6300 7170 6340 7175
rect 6300 7140 6305 7170
rect 6305 7140 6335 7170
rect 6335 7140 6340 7170
rect 6300 7135 6340 7140
rect 6300 7100 6340 7105
rect 6300 7070 6305 7100
rect 6305 7070 6335 7100
rect 6335 7070 6340 7100
rect 6300 7065 6340 7070
rect 6300 7030 6340 7035
rect 6300 7000 6305 7030
rect 6305 7000 6335 7030
rect 6335 7000 6340 7030
rect 6300 6995 6340 7000
rect 6300 6960 6340 6965
rect 6300 6930 6305 6960
rect 6305 6930 6335 6960
rect 6335 6930 6340 6960
rect 6300 6925 6340 6930
rect 6300 6895 6340 6900
rect 6300 6865 6305 6895
rect 6305 6865 6335 6895
rect 6335 6865 6340 6895
rect 6300 6860 6340 6865
rect 6300 6835 6340 6840
rect 6300 6805 6305 6835
rect 6305 6805 6335 6835
rect 6335 6805 6340 6835
rect 6300 6800 6340 6805
rect 6300 6770 6340 6775
rect 6300 6740 6305 6770
rect 6305 6740 6335 6770
rect 6335 6740 6340 6770
rect 6300 6735 6340 6740
rect 6300 6700 6340 6705
rect 6300 6670 6305 6700
rect 6305 6670 6335 6700
rect 6335 6670 6340 6700
rect 6300 6665 6340 6670
rect 6300 6630 6340 6635
rect 6300 6600 6305 6630
rect 6305 6600 6335 6630
rect 6335 6600 6340 6630
rect 6300 6595 6340 6600
rect 6300 6560 6340 6565
rect 6300 6530 6305 6560
rect 6305 6530 6335 6560
rect 6335 6530 6340 6560
rect 6300 6525 6340 6530
rect 6300 6495 6340 6500
rect 6300 6465 6305 6495
rect 6305 6465 6335 6495
rect 6335 6465 6340 6495
rect 6300 6460 6340 6465
rect 6590 9635 6630 9640
rect 6590 9605 6595 9635
rect 6595 9605 6625 9635
rect 6625 9605 6630 9635
rect 6590 9600 6630 9605
rect 6590 9570 6630 9575
rect 6590 9540 6595 9570
rect 6595 9540 6625 9570
rect 6625 9540 6630 9570
rect 6590 9535 6630 9540
rect 6590 9500 6630 9505
rect 6590 9470 6595 9500
rect 6595 9470 6625 9500
rect 6625 9470 6630 9500
rect 6590 9465 6630 9470
rect 6590 9430 6630 9435
rect 6590 9400 6595 9430
rect 6595 9400 6625 9430
rect 6625 9400 6630 9430
rect 6590 9395 6630 9400
rect 6590 9360 6630 9365
rect 6590 9330 6595 9360
rect 6595 9330 6625 9360
rect 6625 9330 6630 9360
rect 6590 9325 6630 9330
rect 6590 9295 6630 9300
rect 6590 9265 6595 9295
rect 6595 9265 6625 9295
rect 6625 9265 6630 9295
rect 6590 9260 6630 9265
rect 6590 9235 6630 9240
rect 6590 9205 6595 9235
rect 6595 9205 6625 9235
rect 6625 9205 6630 9235
rect 6590 9200 6630 9205
rect 6590 9170 6630 9175
rect 6590 9140 6595 9170
rect 6595 9140 6625 9170
rect 6625 9140 6630 9170
rect 6590 9135 6630 9140
rect 6590 9100 6630 9105
rect 6590 9070 6595 9100
rect 6595 9070 6625 9100
rect 6625 9070 6630 9100
rect 6590 9065 6630 9070
rect 6590 9030 6630 9035
rect 6590 9000 6595 9030
rect 6595 9000 6625 9030
rect 6625 9000 6630 9030
rect 6590 8995 6630 9000
rect 6590 8960 6630 8965
rect 6590 8930 6595 8960
rect 6595 8930 6625 8960
rect 6625 8930 6630 8960
rect 6590 8925 6630 8930
rect 6590 8895 6630 8900
rect 6590 8865 6595 8895
rect 6595 8865 6625 8895
rect 6625 8865 6630 8895
rect 6590 8860 6630 8865
rect 6590 8835 6630 8840
rect 6590 8805 6595 8835
rect 6595 8805 6625 8835
rect 6625 8805 6630 8835
rect 6590 8800 6630 8805
rect 6590 8770 6630 8775
rect 6590 8740 6595 8770
rect 6595 8740 6625 8770
rect 6625 8740 6630 8770
rect 6590 8735 6630 8740
rect 6590 8700 6630 8705
rect 6590 8670 6595 8700
rect 6595 8670 6625 8700
rect 6625 8670 6630 8700
rect 6590 8665 6630 8670
rect 6590 8630 6630 8635
rect 6590 8600 6595 8630
rect 6595 8600 6625 8630
rect 6625 8600 6630 8630
rect 6590 8595 6630 8600
rect 6590 8560 6630 8565
rect 6590 8530 6595 8560
rect 6595 8530 6625 8560
rect 6625 8530 6630 8560
rect 6590 8525 6630 8530
rect 6590 8495 6630 8500
rect 6590 8465 6595 8495
rect 6595 8465 6625 8495
rect 6625 8465 6630 8495
rect 6590 8460 6630 8465
rect 6590 8435 6630 8440
rect 6590 8405 6595 8435
rect 6595 8405 6625 8435
rect 6625 8405 6630 8435
rect 6590 8400 6630 8405
rect 6590 8370 6630 8375
rect 6590 8340 6595 8370
rect 6595 8340 6625 8370
rect 6625 8340 6630 8370
rect 6590 8335 6630 8340
rect 6590 8300 6630 8305
rect 6590 8270 6595 8300
rect 6595 8270 6625 8300
rect 6625 8270 6630 8300
rect 6590 8265 6630 8270
rect 6590 8230 6630 8235
rect 6590 8200 6595 8230
rect 6595 8200 6625 8230
rect 6625 8200 6630 8230
rect 6590 8195 6630 8200
rect 6590 8160 6630 8165
rect 6590 8130 6595 8160
rect 6595 8130 6625 8160
rect 6625 8130 6630 8160
rect 6590 8125 6630 8130
rect 6590 8095 6630 8100
rect 6590 8065 6595 8095
rect 6595 8065 6625 8095
rect 6625 8065 6630 8095
rect 6590 8060 6630 8065
rect 6590 8035 6630 8040
rect 6590 8005 6595 8035
rect 6595 8005 6625 8035
rect 6625 8005 6630 8035
rect 6590 8000 6630 8005
rect 6590 7970 6630 7975
rect 6590 7940 6595 7970
rect 6595 7940 6625 7970
rect 6625 7940 6630 7970
rect 6590 7935 6630 7940
rect 6590 7900 6630 7905
rect 6590 7870 6595 7900
rect 6595 7870 6625 7900
rect 6625 7870 6630 7900
rect 6590 7865 6630 7870
rect 6590 7830 6630 7835
rect 6590 7800 6595 7830
rect 6595 7800 6625 7830
rect 6625 7800 6630 7830
rect 6590 7795 6630 7800
rect 6590 7760 6630 7765
rect 6590 7730 6595 7760
rect 6595 7730 6625 7760
rect 6625 7730 6630 7760
rect 6590 7725 6630 7730
rect 6590 7695 6630 7700
rect 6590 7665 6595 7695
rect 6595 7665 6625 7695
rect 6625 7665 6630 7695
rect 6590 7660 6630 7665
rect 6590 7635 6630 7640
rect 6590 7605 6595 7635
rect 6595 7605 6625 7635
rect 6625 7605 6630 7635
rect 6590 7600 6630 7605
rect 6590 7570 6630 7575
rect 6590 7540 6595 7570
rect 6595 7540 6625 7570
rect 6625 7540 6630 7570
rect 6590 7535 6630 7540
rect 6590 7500 6630 7505
rect 6590 7470 6595 7500
rect 6595 7470 6625 7500
rect 6625 7470 6630 7500
rect 6590 7465 6630 7470
rect 6590 7430 6630 7435
rect 6590 7400 6595 7430
rect 6595 7400 6625 7430
rect 6625 7400 6630 7430
rect 6590 7395 6630 7400
rect 6590 7360 6630 7365
rect 6590 7330 6595 7360
rect 6595 7330 6625 7360
rect 6625 7330 6630 7360
rect 6590 7325 6630 7330
rect 6590 7295 6630 7300
rect 6590 7265 6595 7295
rect 6595 7265 6625 7295
rect 6625 7265 6630 7295
rect 6590 7260 6630 7265
rect 6590 7235 6630 7240
rect 6590 7205 6595 7235
rect 6595 7205 6625 7235
rect 6625 7205 6630 7235
rect 6590 7200 6630 7205
rect 6590 7170 6630 7175
rect 6590 7140 6595 7170
rect 6595 7140 6625 7170
rect 6625 7140 6630 7170
rect 6590 7135 6630 7140
rect 6590 7100 6630 7105
rect 6590 7070 6595 7100
rect 6595 7070 6625 7100
rect 6625 7070 6630 7100
rect 6590 7065 6630 7070
rect 6590 7030 6630 7035
rect 6590 7000 6595 7030
rect 6595 7000 6625 7030
rect 6625 7000 6630 7030
rect 6590 6995 6630 7000
rect 6590 6960 6630 6965
rect 6590 6930 6595 6960
rect 6595 6930 6625 6960
rect 6625 6930 6630 6960
rect 6590 6925 6630 6930
rect 6590 6895 6630 6900
rect 6590 6865 6595 6895
rect 6595 6865 6625 6895
rect 6625 6865 6630 6895
rect 6590 6860 6630 6865
rect 6590 6835 6630 6840
rect 6590 6805 6595 6835
rect 6595 6805 6625 6835
rect 6625 6805 6630 6835
rect 6590 6800 6630 6805
rect 6590 6770 6630 6775
rect 6590 6740 6595 6770
rect 6595 6740 6625 6770
rect 6625 6740 6630 6770
rect 6590 6735 6630 6740
rect 6590 6700 6630 6705
rect 6590 6670 6595 6700
rect 6595 6670 6625 6700
rect 6625 6670 6630 6700
rect 6590 6665 6630 6670
rect 6590 6630 6630 6635
rect 6590 6600 6595 6630
rect 6595 6600 6625 6630
rect 6625 6600 6630 6630
rect 6590 6595 6630 6600
rect 6590 6560 6630 6565
rect 6590 6530 6595 6560
rect 6595 6530 6625 6560
rect 6625 6530 6630 6560
rect 6590 6525 6630 6530
rect 6590 6495 6630 6500
rect 6590 6465 6595 6495
rect 6595 6465 6625 6495
rect 6625 6465 6630 6495
rect 6590 6460 6630 6465
rect 7270 9635 7310 9640
rect 7270 9605 7275 9635
rect 7275 9605 7305 9635
rect 7305 9605 7310 9635
rect 7270 9600 7310 9605
rect 7270 9570 7310 9575
rect 7270 9540 7275 9570
rect 7275 9540 7305 9570
rect 7305 9540 7310 9570
rect 7270 9535 7310 9540
rect 7270 9500 7310 9505
rect 7270 9470 7275 9500
rect 7275 9470 7305 9500
rect 7305 9470 7310 9500
rect 7270 9465 7310 9470
rect 7270 9430 7310 9435
rect 7270 9400 7275 9430
rect 7275 9400 7305 9430
rect 7305 9400 7310 9430
rect 7270 9395 7310 9400
rect 7270 9360 7310 9365
rect 7270 9330 7275 9360
rect 7275 9330 7305 9360
rect 7305 9330 7310 9360
rect 7270 9325 7310 9330
rect 7270 9295 7310 9300
rect 7270 9265 7275 9295
rect 7275 9265 7305 9295
rect 7305 9265 7310 9295
rect 7270 9260 7310 9265
rect 7270 9235 7310 9240
rect 7270 9205 7275 9235
rect 7275 9205 7305 9235
rect 7305 9205 7310 9235
rect 7270 9200 7310 9205
rect 7270 9170 7310 9175
rect 7270 9140 7275 9170
rect 7275 9140 7305 9170
rect 7305 9140 7310 9170
rect 7270 9135 7310 9140
rect 7270 9100 7310 9105
rect 7270 9070 7275 9100
rect 7275 9070 7305 9100
rect 7305 9070 7310 9100
rect 7270 9065 7310 9070
rect 7270 9030 7310 9035
rect 7270 9000 7275 9030
rect 7275 9000 7305 9030
rect 7305 9000 7310 9030
rect 7270 8995 7310 9000
rect 7270 8960 7310 8965
rect 7270 8930 7275 8960
rect 7275 8930 7305 8960
rect 7305 8930 7310 8960
rect 7270 8925 7310 8930
rect 7270 8895 7310 8900
rect 7270 8865 7275 8895
rect 7275 8865 7305 8895
rect 7305 8865 7310 8895
rect 7270 8860 7310 8865
rect 7270 8835 7310 8840
rect 7270 8805 7275 8835
rect 7275 8805 7305 8835
rect 7305 8805 7310 8835
rect 7270 8800 7310 8805
rect 7270 8770 7310 8775
rect 7270 8740 7275 8770
rect 7275 8740 7305 8770
rect 7305 8740 7310 8770
rect 7270 8735 7310 8740
rect 7270 8700 7310 8705
rect 7270 8670 7275 8700
rect 7275 8670 7305 8700
rect 7305 8670 7310 8700
rect 7270 8665 7310 8670
rect 7270 8630 7310 8635
rect 7270 8600 7275 8630
rect 7275 8600 7305 8630
rect 7305 8600 7310 8630
rect 7270 8595 7310 8600
rect 7270 8560 7310 8565
rect 7270 8530 7275 8560
rect 7275 8530 7305 8560
rect 7305 8530 7310 8560
rect 7270 8525 7310 8530
rect 7270 8495 7310 8500
rect 7270 8465 7275 8495
rect 7275 8465 7305 8495
rect 7305 8465 7310 8495
rect 7270 8460 7310 8465
rect 7270 8435 7310 8440
rect 7270 8405 7275 8435
rect 7275 8405 7305 8435
rect 7305 8405 7310 8435
rect 7270 8400 7310 8405
rect 7270 8370 7310 8375
rect 7270 8340 7275 8370
rect 7275 8340 7305 8370
rect 7305 8340 7310 8370
rect 7270 8335 7310 8340
rect 7270 8300 7310 8305
rect 7270 8270 7275 8300
rect 7275 8270 7305 8300
rect 7305 8270 7310 8300
rect 7270 8265 7310 8270
rect 7270 8230 7310 8235
rect 7270 8200 7275 8230
rect 7275 8200 7305 8230
rect 7305 8200 7310 8230
rect 7270 8195 7310 8200
rect 7270 8160 7310 8165
rect 7270 8130 7275 8160
rect 7275 8130 7305 8160
rect 7305 8130 7310 8160
rect 7270 8125 7310 8130
rect 7270 8095 7310 8100
rect 7270 8065 7275 8095
rect 7275 8065 7305 8095
rect 7305 8065 7310 8095
rect 7270 8060 7310 8065
rect 7270 8035 7310 8040
rect 7270 8005 7275 8035
rect 7275 8005 7305 8035
rect 7305 8005 7310 8035
rect 7270 8000 7310 8005
rect 7270 7970 7310 7975
rect 7270 7940 7275 7970
rect 7275 7940 7305 7970
rect 7305 7940 7310 7970
rect 7270 7935 7310 7940
rect 7270 7900 7310 7905
rect 7270 7870 7275 7900
rect 7275 7870 7305 7900
rect 7305 7870 7310 7900
rect 7270 7865 7310 7870
rect 7270 7830 7310 7835
rect 7270 7800 7275 7830
rect 7275 7800 7305 7830
rect 7305 7800 7310 7830
rect 7270 7795 7310 7800
rect 7270 7760 7310 7765
rect 7270 7730 7275 7760
rect 7275 7730 7305 7760
rect 7305 7730 7310 7760
rect 7270 7725 7310 7730
rect 7270 7695 7310 7700
rect 7270 7665 7275 7695
rect 7275 7665 7305 7695
rect 7305 7665 7310 7695
rect 7270 7660 7310 7665
rect 7270 7635 7310 7640
rect 7270 7605 7275 7635
rect 7275 7605 7305 7635
rect 7305 7605 7310 7635
rect 7270 7600 7310 7605
rect 7270 7570 7310 7575
rect 7270 7540 7275 7570
rect 7275 7540 7305 7570
rect 7305 7540 7310 7570
rect 7270 7535 7310 7540
rect 7270 7500 7310 7505
rect 7270 7470 7275 7500
rect 7275 7470 7305 7500
rect 7305 7470 7310 7500
rect 7270 7465 7310 7470
rect 7270 7430 7310 7435
rect 7270 7400 7275 7430
rect 7275 7400 7305 7430
rect 7305 7400 7310 7430
rect 7270 7395 7310 7400
rect 7270 7360 7310 7365
rect 7270 7330 7275 7360
rect 7275 7330 7305 7360
rect 7305 7330 7310 7360
rect 7270 7325 7310 7330
rect 7270 7295 7310 7300
rect 7270 7265 7275 7295
rect 7275 7265 7305 7295
rect 7305 7265 7310 7295
rect 7270 7260 7310 7265
rect 7270 7235 7310 7240
rect 7270 7205 7275 7235
rect 7275 7205 7305 7235
rect 7305 7205 7310 7235
rect 7270 7200 7310 7205
rect 7270 7170 7310 7175
rect 7270 7140 7275 7170
rect 7275 7140 7305 7170
rect 7305 7140 7310 7170
rect 7270 7135 7310 7140
rect 7270 7100 7310 7105
rect 7270 7070 7275 7100
rect 7275 7070 7305 7100
rect 7305 7070 7310 7100
rect 7270 7065 7310 7070
rect 7270 7030 7310 7035
rect 7270 7000 7275 7030
rect 7275 7000 7305 7030
rect 7305 7000 7310 7030
rect 7270 6995 7310 7000
rect 7270 6960 7310 6965
rect 7270 6930 7275 6960
rect 7275 6930 7305 6960
rect 7305 6930 7310 6960
rect 7270 6925 7310 6930
rect 7270 6895 7310 6900
rect 7270 6865 7275 6895
rect 7275 6865 7305 6895
rect 7305 6865 7310 6895
rect 7270 6860 7310 6865
rect 7270 6835 7310 6840
rect 7270 6805 7275 6835
rect 7275 6805 7305 6835
rect 7305 6805 7310 6835
rect 7270 6800 7310 6805
rect 7270 6770 7310 6775
rect 7270 6740 7275 6770
rect 7275 6740 7305 6770
rect 7305 6740 7310 6770
rect 7270 6735 7310 6740
rect 7270 6700 7310 6705
rect 7270 6670 7275 6700
rect 7275 6670 7305 6700
rect 7305 6670 7310 6700
rect 7270 6665 7310 6670
rect 7270 6630 7310 6635
rect 7270 6600 7275 6630
rect 7275 6600 7305 6630
rect 7305 6600 7310 6630
rect 7270 6595 7310 6600
rect 7270 6560 7310 6565
rect 7270 6530 7275 6560
rect 7275 6530 7305 6560
rect 7305 6530 7310 6560
rect 7270 6525 7310 6530
rect 7270 6495 7310 6500
rect 7270 6465 7275 6495
rect 7275 6465 7305 6495
rect 7305 6465 7310 6495
rect 7270 6460 7310 6465
rect 7620 9635 7660 9640
rect 7620 9605 7625 9635
rect 7625 9605 7655 9635
rect 7655 9605 7660 9635
rect 7620 9600 7660 9605
rect 7620 9570 7660 9575
rect 7620 9540 7625 9570
rect 7625 9540 7655 9570
rect 7655 9540 7660 9570
rect 7620 9535 7660 9540
rect 7620 9500 7660 9505
rect 7620 9470 7625 9500
rect 7625 9470 7655 9500
rect 7655 9470 7660 9500
rect 7620 9465 7660 9470
rect 7620 9430 7660 9435
rect 7620 9400 7625 9430
rect 7625 9400 7655 9430
rect 7655 9400 7660 9430
rect 7620 9395 7660 9400
rect 7620 9360 7660 9365
rect 7620 9330 7625 9360
rect 7625 9330 7655 9360
rect 7655 9330 7660 9360
rect 7620 9325 7660 9330
rect 7620 9295 7660 9300
rect 7620 9265 7625 9295
rect 7625 9265 7655 9295
rect 7655 9265 7660 9295
rect 7620 9260 7660 9265
rect 7620 9235 7660 9240
rect 7620 9205 7625 9235
rect 7625 9205 7655 9235
rect 7655 9205 7660 9235
rect 7620 9200 7660 9205
rect 7620 9170 7660 9175
rect 7620 9140 7625 9170
rect 7625 9140 7655 9170
rect 7655 9140 7660 9170
rect 7620 9135 7660 9140
rect 7620 9100 7660 9105
rect 7620 9070 7625 9100
rect 7625 9070 7655 9100
rect 7655 9070 7660 9100
rect 7620 9065 7660 9070
rect 7620 9030 7660 9035
rect 7620 9000 7625 9030
rect 7625 9000 7655 9030
rect 7655 9000 7660 9030
rect 7620 8995 7660 9000
rect 7620 8960 7660 8965
rect 7620 8930 7625 8960
rect 7625 8930 7655 8960
rect 7655 8930 7660 8960
rect 7620 8925 7660 8930
rect 7620 8895 7660 8900
rect 7620 8865 7625 8895
rect 7625 8865 7655 8895
rect 7655 8865 7660 8895
rect 7620 8860 7660 8865
rect 7620 8835 7660 8840
rect 7620 8805 7625 8835
rect 7625 8805 7655 8835
rect 7655 8805 7660 8835
rect 7620 8800 7660 8805
rect 7620 8770 7660 8775
rect 7620 8740 7625 8770
rect 7625 8740 7655 8770
rect 7655 8740 7660 8770
rect 7620 8735 7660 8740
rect 7620 8700 7660 8705
rect 7620 8670 7625 8700
rect 7625 8670 7655 8700
rect 7655 8670 7660 8700
rect 7620 8665 7660 8670
rect 7620 8630 7660 8635
rect 7620 8600 7625 8630
rect 7625 8600 7655 8630
rect 7655 8600 7660 8630
rect 7620 8595 7660 8600
rect 7620 8560 7660 8565
rect 7620 8530 7625 8560
rect 7625 8530 7655 8560
rect 7655 8530 7660 8560
rect 7620 8525 7660 8530
rect 7620 8495 7660 8500
rect 7620 8465 7625 8495
rect 7625 8465 7655 8495
rect 7655 8465 7660 8495
rect 7620 8460 7660 8465
rect 7620 8435 7660 8440
rect 7620 8405 7625 8435
rect 7625 8405 7655 8435
rect 7655 8405 7660 8435
rect 7620 8400 7660 8405
rect 7620 8370 7660 8375
rect 7620 8340 7625 8370
rect 7625 8340 7655 8370
rect 7655 8340 7660 8370
rect 7620 8335 7660 8340
rect 7620 8300 7660 8305
rect 7620 8270 7625 8300
rect 7625 8270 7655 8300
rect 7655 8270 7660 8300
rect 7620 8265 7660 8270
rect 7620 8230 7660 8235
rect 7620 8200 7625 8230
rect 7625 8200 7655 8230
rect 7655 8200 7660 8230
rect 7620 8195 7660 8200
rect 7620 8160 7660 8165
rect 7620 8130 7625 8160
rect 7625 8130 7655 8160
rect 7655 8130 7660 8160
rect 7620 8125 7660 8130
rect 7620 8095 7660 8100
rect 7620 8065 7625 8095
rect 7625 8065 7655 8095
rect 7655 8065 7660 8095
rect 7620 8060 7660 8065
rect 7620 8035 7660 8040
rect 7620 8005 7625 8035
rect 7625 8005 7655 8035
rect 7655 8005 7660 8035
rect 7620 8000 7660 8005
rect 7620 7970 7660 7975
rect 7620 7940 7625 7970
rect 7625 7940 7655 7970
rect 7655 7940 7660 7970
rect 7620 7935 7660 7940
rect 7620 7900 7660 7905
rect 7620 7870 7625 7900
rect 7625 7870 7655 7900
rect 7655 7870 7660 7900
rect 7620 7865 7660 7870
rect 7620 7830 7660 7835
rect 7620 7800 7625 7830
rect 7625 7800 7655 7830
rect 7655 7800 7660 7830
rect 7620 7795 7660 7800
rect 7620 7760 7660 7765
rect 7620 7730 7625 7760
rect 7625 7730 7655 7760
rect 7655 7730 7660 7760
rect 7620 7725 7660 7730
rect 7620 7695 7660 7700
rect 7620 7665 7625 7695
rect 7625 7665 7655 7695
rect 7655 7665 7660 7695
rect 7620 7660 7660 7665
rect 7620 7635 7660 7640
rect 7620 7605 7625 7635
rect 7625 7605 7655 7635
rect 7655 7605 7660 7635
rect 7620 7600 7660 7605
rect 7620 7570 7660 7575
rect 7620 7540 7625 7570
rect 7625 7540 7655 7570
rect 7655 7540 7660 7570
rect 7620 7535 7660 7540
rect 7620 7500 7660 7505
rect 7620 7470 7625 7500
rect 7625 7470 7655 7500
rect 7655 7470 7660 7500
rect 7620 7465 7660 7470
rect 7620 7430 7660 7435
rect 7620 7400 7625 7430
rect 7625 7400 7655 7430
rect 7655 7400 7660 7430
rect 7620 7395 7660 7400
rect 7620 7360 7660 7365
rect 7620 7330 7625 7360
rect 7625 7330 7655 7360
rect 7655 7330 7660 7360
rect 7620 7325 7660 7330
rect 7620 7295 7660 7300
rect 7620 7265 7625 7295
rect 7625 7265 7655 7295
rect 7655 7265 7660 7295
rect 7620 7260 7660 7265
rect 7620 7235 7660 7240
rect 7620 7205 7625 7235
rect 7625 7205 7655 7235
rect 7655 7205 7660 7235
rect 7620 7200 7660 7205
rect 7620 7170 7660 7175
rect 7620 7140 7625 7170
rect 7625 7140 7655 7170
rect 7655 7140 7660 7170
rect 7620 7135 7660 7140
rect 7620 7100 7660 7105
rect 7620 7070 7625 7100
rect 7625 7070 7655 7100
rect 7655 7070 7660 7100
rect 7620 7065 7660 7070
rect 7620 7030 7660 7035
rect 7620 7000 7625 7030
rect 7625 7000 7655 7030
rect 7655 7000 7660 7030
rect 7620 6995 7660 7000
rect 7620 6960 7660 6965
rect 7620 6930 7625 6960
rect 7625 6930 7655 6960
rect 7655 6930 7660 6960
rect 7620 6925 7660 6930
rect 7620 6895 7660 6900
rect 7620 6865 7625 6895
rect 7625 6865 7655 6895
rect 7655 6865 7660 6895
rect 7620 6860 7660 6865
rect 7620 6835 7660 6840
rect 7620 6805 7625 6835
rect 7625 6805 7655 6835
rect 7655 6805 7660 6835
rect 7620 6800 7660 6805
rect 7620 6770 7660 6775
rect 7620 6740 7625 6770
rect 7625 6740 7655 6770
rect 7655 6740 7660 6770
rect 7620 6735 7660 6740
rect 7620 6700 7660 6705
rect 7620 6670 7625 6700
rect 7625 6670 7655 6700
rect 7655 6670 7660 6700
rect 7620 6665 7660 6670
rect 7620 6630 7660 6635
rect 7620 6600 7625 6630
rect 7625 6600 7655 6630
rect 7655 6600 7660 6630
rect 7620 6595 7660 6600
rect 7620 6560 7660 6565
rect 7620 6530 7625 6560
rect 7625 6530 7655 6560
rect 7655 6530 7660 6560
rect 7620 6525 7660 6530
rect 7620 6495 7660 6500
rect 7620 6465 7625 6495
rect 7625 6465 7655 6495
rect 7655 6465 7660 6495
rect 7620 6460 7660 6465
rect 8320 9635 8360 9640
rect 8320 9605 8325 9635
rect 8325 9605 8355 9635
rect 8355 9605 8360 9635
rect 8320 9600 8360 9605
rect 8320 9570 8360 9575
rect 8320 9540 8325 9570
rect 8325 9540 8355 9570
rect 8355 9540 8360 9570
rect 8320 9535 8360 9540
rect 8320 9500 8360 9505
rect 8320 9470 8325 9500
rect 8325 9470 8355 9500
rect 8355 9470 8360 9500
rect 8320 9465 8360 9470
rect 8320 9430 8360 9435
rect 8320 9400 8325 9430
rect 8325 9400 8355 9430
rect 8355 9400 8360 9430
rect 8320 9395 8360 9400
rect 8320 9360 8360 9365
rect 8320 9330 8325 9360
rect 8325 9330 8355 9360
rect 8355 9330 8360 9360
rect 8320 9325 8360 9330
rect 8320 9295 8360 9300
rect 8320 9265 8325 9295
rect 8325 9265 8355 9295
rect 8355 9265 8360 9295
rect 8320 9260 8360 9265
rect 8320 9235 8360 9240
rect 8320 9205 8325 9235
rect 8325 9205 8355 9235
rect 8355 9205 8360 9235
rect 8320 9200 8360 9205
rect 8320 9170 8360 9175
rect 8320 9140 8325 9170
rect 8325 9140 8355 9170
rect 8355 9140 8360 9170
rect 8320 9135 8360 9140
rect 8320 9100 8360 9105
rect 8320 9070 8325 9100
rect 8325 9070 8355 9100
rect 8355 9070 8360 9100
rect 8320 9065 8360 9070
rect 8320 9030 8360 9035
rect 8320 9000 8325 9030
rect 8325 9000 8355 9030
rect 8355 9000 8360 9030
rect 8320 8995 8360 9000
rect 8320 8960 8360 8965
rect 8320 8930 8325 8960
rect 8325 8930 8355 8960
rect 8355 8930 8360 8960
rect 8320 8925 8360 8930
rect 8320 8895 8360 8900
rect 8320 8865 8325 8895
rect 8325 8865 8355 8895
rect 8355 8865 8360 8895
rect 8320 8860 8360 8865
rect 8320 8835 8360 8840
rect 8320 8805 8325 8835
rect 8325 8805 8355 8835
rect 8355 8805 8360 8835
rect 8320 8800 8360 8805
rect 8320 8770 8360 8775
rect 8320 8740 8325 8770
rect 8325 8740 8355 8770
rect 8355 8740 8360 8770
rect 8320 8735 8360 8740
rect 8320 8700 8360 8705
rect 8320 8670 8325 8700
rect 8325 8670 8355 8700
rect 8355 8670 8360 8700
rect 8320 8665 8360 8670
rect 8320 8630 8360 8635
rect 8320 8600 8325 8630
rect 8325 8600 8355 8630
rect 8355 8600 8360 8630
rect 8320 8595 8360 8600
rect 8320 8560 8360 8565
rect 8320 8530 8325 8560
rect 8325 8530 8355 8560
rect 8355 8530 8360 8560
rect 8320 8525 8360 8530
rect 8320 8495 8360 8500
rect 8320 8465 8325 8495
rect 8325 8465 8355 8495
rect 8355 8465 8360 8495
rect 8320 8460 8360 8465
rect 8320 8435 8360 8440
rect 8320 8405 8325 8435
rect 8325 8405 8355 8435
rect 8355 8405 8360 8435
rect 8320 8400 8360 8405
rect 8320 8370 8360 8375
rect 8320 8340 8325 8370
rect 8325 8340 8355 8370
rect 8355 8340 8360 8370
rect 8320 8335 8360 8340
rect 8320 8300 8360 8305
rect 8320 8270 8325 8300
rect 8325 8270 8355 8300
rect 8355 8270 8360 8300
rect 8320 8265 8360 8270
rect 8320 8230 8360 8235
rect 8320 8200 8325 8230
rect 8325 8200 8355 8230
rect 8355 8200 8360 8230
rect 8320 8195 8360 8200
rect 8320 8160 8360 8165
rect 8320 8130 8325 8160
rect 8325 8130 8355 8160
rect 8355 8130 8360 8160
rect 8320 8125 8360 8130
rect 8320 8095 8360 8100
rect 8320 8065 8325 8095
rect 8325 8065 8355 8095
rect 8355 8065 8360 8095
rect 8320 8060 8360 8065
rect 8320 8035 8360 8040
rect 8320 8005 8325 8035
rect 8325 8005 8355 8035
rect 8355 8005 8360 8035
rect 8320 8000 8360 8005
rect 8320 7970 8360 7975
rect 8320 7940 8325 7970
rect 8325 7940 8355 7970
rect 8355 7940 8360 7970
rect 8320 7935 8360 7940
rect 8320 7900 8360 7905
rect 8320 7870 8325 7900
rect 8325 7870 8355 7900
rect 8355 7870 8360 7900
rect 8320 7865 8360 7870
rect 8320 7830 8360 7835
rect 8320 7800 8325 7830
rect 8325 7800 8355 7830
rect 8355 7800 8360 7830
rect 8320 7795 8360 7800
rect 8320 7760 8360 7765
rect 8320 7730 8325 7760
rect 8325 7730 8355 7760
rect 8355 7730 8360 7760
rect 8320 7725 8360 7730
rect 8320 7695 8360 7700
rect 8320 7665 8325 7695
rect 8325 7665 8355 7695
rect 8355 7665 8360 7695
rect 8320 7660 8360 7665
rect 8320 7635 8360 7640
rect 8320 7605 8325 7635
rect 8325 7605 8355 7635
rect 8355 7605 8360 7635
rect 8320 7600 8360 7605
rect 8320 7570 8360 7575
rect 8320 7540 8325 7570
rect 8325 7540 8355 7570
rect 8355 7540 8360 7570
rect 8320 7535 8360 7540
rect 8320 7500 8360 7505
rect 8320 7470 8325 7500
rect 8325 7470 8355 7500
rect 8355 7470 8360 7500
rect 8320 7465 8360 7470
rect 8320 7430 8360 7435
rect 8320 7400 8325 7430
rect 8325 7400 8355 7430
rect 8355 7400 8360 7430
rect 8320 7395 8360 7400
rect 8320 7360 8360 7365
rect 8320 7330 8325 7360
rect 8325 7330 8355 7360
rect 8355 7330 8360 7360
rect 8320 7325 8360 7330
rect 8320 7295 8360 7300
rect 8320 7265 8325 7295
rect 8325 7265 8355 7295
rect 8355 7265 8360 7295
rect 8320 7260 8360 7265
rect 8320 7235 8360 7240
rect 8320 7205 8325 7235
rect 8325 7205 8355 7235
rect 8355 7205 8360 7235
rect 8320 7200 8360 7205
rect 8320 7170 8360 7175
rect 8320 7140 8325 7170
rect 8325 7140 8355 7170
rect 8355 7140 8360 7170
rect 8320 7135 8360 7140
rect 8320 7100 8360 7105
rect 8320 7070 8325 7100
rect 8325 7070 8355 7100
rect 8355 7070 8360 7100
rect 8320 7065 8360 7070
rect 8320 7030 8360 7035
rect 8320 7000 8325 7030
rect 8325 7000 8355 7030
rect 8355 7000 8360 7030
rect 8320 6995 8360 7000
rect 8320 6960 8360 6965
rect 8320 6930 8325 6960
rect 8325 6930 8355 6960
rect 8355 6930 8360 6960
rect 8320 6925 8360 6930
rect 8320 6895 8360 6900
rect 8320 6865 8325 6895
rect 8325 6865 8355 6895
rect 8355 6865 8360 6895
rect 8320 6860 8360 6865
rect 8320 6835 8360 6840
rect 8320 6805 8325 6835
rect 8325 6805 8355 6835
rect 8355 6805 8360 6835
rect 8320 6800 8360 6805
rect 8320 6770 8360 6775
rect 8320 6740 8325 6770
rect 8325 6740 8355 6770
rect 8355 6740 8360 6770
rect 8320 6735 8360 6740
rect 8320 6700 8360 6705
rect 8320 6670 8325 6700
rect 8325 6670 8355 6700
rect 8355 6670 8360 6700
rect 8320 6665 8360 6670
rect 8320 6630 8360 6635
rect 8320 6600 8325 6630
rect 8325 6600 8355 6630
rect 8355 6600 8360 6630
rect 8320 6595 8360 6600
rect 8320 6560 8360 6565
rect 8320 6530 8325 6560
rect 8325 6530 8355 6560
rect 8355 6530 8360 6560
rect 8320 6525 8360 6530
rect 8320 6495 8360 6500
rect 8320 6465 8325 6495
rect 8325 6465 8355 6495
rect 8355 6465 8360 6495
rect 8320 6460 8360 6465
rect 8670 9635 8710 9640
rect 8670 9605 8675 9635
rect 8675 9605 8705 9635
rect 8705 9605 8710 9635
rect 8670 9600 8710 9605
rect 8670 9570 8710 9575
rect 8670 9540 8675 9570
rect 8675 9540 8705 9570
rect 8705 9540 8710 9570
rect 8670 9535 8710 9540
rect 8670 9500 8710 9505
rect 8670 9470 8675 9500
rect 8675 9470 8705 9500
rect 8705 9470 8710 9500
rect 8670 9465 8710 9470
rect 8670 9430 8710 9435
rect 8670 9400 8675 9430
rect 8675 9400 8705 9430
rect 8705 9400 8710 9430
rect 8670 9395 8710 9400
rect 8670 9360 8710 9365
rect 8670 9330 8675 9360
rect 8675 9330 8705 9360
rect 8705 9330 8710 9360
rect 8670 9325 8710 9330
rect 8670 9295 8710 9300
rect 8670 9265 8675 9295
rect 8675 9265 8705 9295
rect 8705 9265 8710 9295
rect 8670 9260 8710 9265
rect 8670 9235 8710 9240
rect 8670 9205 8675 9235
rect 8675 9205 8705 9235
rect 8705 9205 8710 9235
rect 8670 9200 8710 9205
rect 8670 9170 8710 9175
rect 8670 9140 8675 9170
rect 8675 9140 8705 9170
rect 8705 9140 8710 9170
rect 8670 9135 8710 9140
rect 8670 9100 8710 9105
rect 8670 9070 8675 9100
rect 8675 9070 8705 9100
rect 8705 9070 8710 9100
rect 8670 9065 8710 9070
rect 8670 9030 8710 9035
rect 8670 9000 8675 9030
rect 8675 9000 8705 9030
rect 8705 9000 8710 9030
rect 8670 8995 8710 9000
rect 8670 8960 8710 8965
rect 8670 8930 8675 8960
rect 8675 8930 8705 8960
rect 8705 8930 8710 8960
rect 8670 8925 8710 8930
rect 8670 8895 8710 8900
rect 8670 8865 8675 8895
rect 8675 8865 8705 8895
rect 8705 8865 8710 8895
rect 8670 8860 8710 8865
rect 8670 8835 8710 8840
rect 8670 8805 8675 8835
rect 8675 8805 8705 8835
rect 8705 8805 8710 8835
rect 8670 8800 8710 8805
rect 8670 8770 8710 8775
rect 8670 8740 8675 8770
rect 8675 8740 8705 8770
rect 8705 8740 8710 8770
rect 8670 8735 8710 8740
rect 8670 8700 8710 8705
rect 8670 8670 8675 8700
rect 8675 8670 8705 8700
rect 8705 8670 8710 8700
rect 8670 8665 8710 8670
rect 8670 8630 8710 8635
rect 8670 8600 8675 8630
rect 8675 8600 8705 8630
rect 8705 8600 8710 8630
rect 8670 8595 8710 8600
rect 8670 8560 8710 8565
rect 8670 8530 8675 8560
rect 8675 8530 8705 8560
rect 8705 8530 8710 8560
rect 8670 8525 8710 8530
rect 8670 8495 8710 8500
rect 8670 8465 8675 8495
rect 8675 8465 8705 8495
rect 8705 8465 8710 8495
rect 8670 8460 8710 8465
rect 8670 8435 8710 8440
rect 8670 8405 8675 8435
rect 8675 8405 8705 8435
rect 8705 8405 8710 8435
rect 8670 8400 8710 8405
rect 8670 8370 8710 8375
rect 8670 8340 8675 8370
rect 8675 8340 8705 8370
rect 8705 8340 8710 8370
rect 8670 8335 8710 8340
rect 8670 8300 8710 8305
rect 8670 8270 8675 8300
rect 8675 8270 8705 8300
rect 8705 8270 8710 8300
rect 8670 8265 8710 8270
rect 8670 8230 8710 8235
rect 8670 8200 8675 8230
rect 8675 8200 8705 8230
rect 8705 8200 8710 8230
rect 8670 8195 8710 8200
rect 8670 8160 8710 8165
rect 8670 8130 8675 8160
rect 8675 8130 8705 8160
rect 8705 8130 8710 8160
rect 8670 8125 8710 8130
rect 8670 8095 8710 8100
rect 8670 8065 8675 8095
rect 8675 8065 8705 8095
rect 8705 8065 8710 8095
rect 8670 8060 8710 8065
rect 8670 8035 8710 8040
rect 8670 8005 8675 8035
rect 8675 8005 8705 8035
rect 8705 8005 8710 8035
rect 8670 8000 8710 8005
rect 8670 7970 8710 7975
rect 8670 7940 8675 7970
rect 8675 7940 8705 7970
rect 8705 7940 8710 7970
rect 8670 7935 8710 7940
rect 8670 7900 8710 7905
rect 8670 7870 8675 7900
rect 8675 7870 8705 7900
rect 8705 7870 8710 7900
rect 8670 7865 8710 7870
rect 8670 7830 8710 7835
rect 8670 7800 8675 7830
rect 8675 7800 8705 7830
rect 8705 7800 8710 7830
rect 8670 7795 8710 7800
rect 8670 7760 8710 7765
rect 8670 7730 8675 7760
rect 8675 7730 8705 7760
rect 8705 7730 8710 7760
rect 8670 7725 8710 7730
rect 8670 7695 8710 7700
rect 8670 7665 8675 7695
rect 8675 7665 8705 7695
rect 8705 7665 8710 7695
rect 8670 7660 8710 7665
rect 8670 7635 8710 7640
rect 8670 7605 8675 7635
rect 8675 7605 8705 7635
rect 8705 7605 8710 7635
rect 8670 7600 8710 7605
rect 8670 7570 8710 7575
rect 8670 7540 8675 7570
rect 8675 7540 8705 7570
rect 8705 7540 8710 7570
rect 8670 7535 8710 7540
rect 8670 7500 8710 7505
rect 8670 7470 8675 7500
rect 8675 7470 8705 7500
rect 8705 7470 8710 7500
rect 8670 7465 8710 7470
rect 8670 7430 8710 7435
rect 8670 7400 8675 7430
rect 8675 7400 8705 7430
rect 8705 7400 8710 7430
rect 8670 7395 8710 7400
rect 8670 7360 8710 7365
rect 8670 7330 8675 7360
rect 8675 7330 8705 7360
rect 8705 7330 8710 7360
rect 8670 7325 8710 7330
rect 8670 7295 8710 7300
rect 8670 7265 8675 7295
rect 8675 7265 8705 7295
rect 8705 7265 8710 7295
rect 8670 7260 8710 7265
rect 8670 7235 8710 7240
rect 8670 7205 8675 7235
rect 8675 7205 8705 7235
rect 8705 7205 8710 7235
rect 8670 7200 8710 7205
rect 8670 7170 8710 7175
rect 8670 7140 8675 7170
rect 8675 7140 8705 7170
rect 8705 7140 8710 7170
rect 8670 7135 8710 7140
rect 8670 7100 8710 7105
rect 8670 7070 8675 7100
rect 8675 7070 8705 7100
rect 8705 7070 8710 7100
rect 8670 7065 8710 7070
rect 8670 7030 8710 7035
rect 8670 7000 8675 7030
rect 8675 7000 8705 7030
rect 8705 7000 8710 7030
rect 8670 6995 8710 7000
rect 8670 6960 8710 6965
rect 8670 6930 8675 6960
rect 8675 6930 8705 6960
rect 8705 6930 8710 6960
rect 8670 6925 8710 6930
rect 8670 6895 8710 6900
rect 8670 6865 8675 6895
rect 8675 6865 8705 6895
rect 8705 6865 8710 6895
rect 8670 6860 8710 6865
rect 8670 6835 8710 6840
rect 8670 6805 8675 6835
rect 8675 6805 8705 6835
rect 8705 6805 8710 6835
rect 8670 6800 8710 6805
rect 8670 6770 8710 6775
rect 8670 6740 8675 6770
rect 8675 6740 8705 6770
rect 8705 6740 8710 6770
rect 8670 6735 8710 6740
rect 8670 6700 8710 6705
rect 8670 6670 8675 6700
rect 8675 6670 8705 6700
rect 8705 6670 8710 6700
rect 8670 6665 8710 6670
rect 8670 6630 8710 6635
rect 8670 6600 8675 6630
rect 8675 6600 8705 6630
rect 8705 6600 8710 6630
rect 8670 6595 8710 6600
rect 8670 6560 8710 6565
rect 8670 6530 8675 6560
rect 8675 6530 8705 6560
rect 8705 6530 8710 6560
rect 8670 6525 8710 6530
rect 8670 6495 8710 6500
rect 8670 6465 8675 6495
rect 8675 6465 8705 6495
rect 8705 6465 8710 6495
rect 8670 6460 8710 6465
rect 9020 9635 9060 9640
rect 9020 9605 9025 9635
rect 9025 9605 9055 9635
rect 9055 9605 9060 9635
rect 9020 9600 9060 9605
rect 9020 9570 9060 9575
rect 9020 9540 9025 9570
rect 9025 9540 9055 9570
rect 9055 9540 9060 9570
rect 9020 9535 9060 9540
rect 9020 9500 9060 9505
rect 9020 9470 9025 9500
rect 9025 9470 9055 9500
rect 9055 9470 9060 9500
rect 9020 9465 9060 9470
rect 14825 9565 14875 9615
rect 14920 9565 14970 9615
rect 15015 9565 15065 9615
rect 15115 9565 15165 9615
rect 15215 9565 15265 9615
rect 15315 9565 15365 9615
rect 15410 9565 15460 9615
rect 15505 9565 15555 9615
rect 15625 9565 15675 9615
rect 15720 9565 15770 9615
rect 15815 9565 15865 9615
rect 15915 9565 15965 9615
rect 16015 9565 16065 9615
rect 16115 9565 16165 9615
rect 16210 9565 16260 9615
rect 16305 9565 16355 9615
rect 16425 9565 16475 9615
rect 16520 9565 16570 9615
rect 16615 9565 16665 9615
rect 16715 9565 16765 9615
rect 16815 9565 16865 9615
rect 16915 9565 16965 9615
rect 17010 9565 17060 9615
rect 17105 9565 17155 9615
rect 17225 9565 17275 9615
rect 17320 9565 17370 9615
rect 17415 9565 17465 9615
rect 17515 9565 17565 9615
rect 17615 9565 17665 9615
rect 17715 9565 17765 9615
rect 17810 9565 17860 9615
rect 17905 9565 17955 9615
rect 9020 9430 9060 9435
rect 9020 9400 9025 9430
rect 9025 9400 9055 9430
rect 9055 9400 9060 9430
rect 9020 9395 9060 9400
rect 9020 9360 9060 9365
rect 9020 9330 9025 9360
rect 9025 9330 9055 9360
rect 9055 9330 9060 9360
rect 9020 9325 9060 9330
rect 9020 9295 9060 9300
rect 9020 9265 9025 9295
rect 9025 9265 9055 9295
rect 9055 9265 9060 9295
rect 9020 9260 9060 9265
rect 14825 9475 14875 9525
rect 14920 9475 14970 9525
rect 15015 9475 15065 9525
rect 15115 9475 15165 9525
rect 15215 9475 15265 9525
rect 15315 9475 15365 9525
rect 15410 9475 15460 9525
rect 15505 9475 15555 9525
rect 15625 9475 15675 9525
rect 15720 9475 15770 9525
rect 15815 9475 15865 9525
rect 15915 9475 15965 9525
rect 16015 9475 16065 9525
rect 16115 9475 16165 9525
rect 16210 9475 16260 9525
rect 16305 9475 16355 9525
rect 16425 9475 16475 9525
rect 16520 9475 16570 9525
rect 16615 9475 16665 9525
rect 16715 9475 16765 9525
rect 16815 9475 16865 9525
rect 16915 9475 16965 9525
rect 17010 9475 17060 9525
rect 17105 9475 17155 9525
rect 17225 9475 17275 9525
rect 17320 9475 17370 9525
rect 17415 9475 17465 9525
rect 17515 9475 17565 9525
rect 17615 9475 17665 9525
rect 17715 9475 17765 9525
rect 17810 9475 17860 9525
rect 17905 9475 17955 9525
rect 14825 9375 14875 9425
rect 14920 9375 14970 9425
rect 15015 9375 15065 9425
rect 15115 9375 15165 9425
rect 15215 9375 15265 9425
rect 15315 9375 15365 9425
rect 15410 9375 15460 9425
rect 15505 9375 15555 9425
rect 15625 9375 15675 9425
rect 15720 9375 15770 9425
rect 15815 9375 15865 9425
rect 15915 9375 15965 9425
rect 16015 9375 16065 9425
rect 16115 9375 16165 9425
rect 16210 9375 16260 9425
rect 16305 9375 16355 9425
rect 16425 9375 16475 9425
rect 16520 9375 16570 9425
rect 16615 9375 16665 9425
rect 16715 9375 16765 9425
rect 16815 9375 16865 9425
rect 16915 9375 16965 9425
rect 17010 9375 17060 9425
rect 17105 9375 17155 9425
rect 17225 9375 17275 9425
rect 17320 9375 17370 9425
rect 17415 9375 17465 9425
rect 17515 9375 17565 9425
rect 17615 9375 17665 9425
rect 17715 9375 17765 9425
rect 17810 9375 17860 9425
rect 17905 9375 17955 9425
rect 14825 9285 14875 9335
rect 14920 9285 14970 9335
rect 15015 9285 15065 9335
rect 15115 9285 15165 9335
rect 15215 9285 15265 9335
rect 15315 9285 15365 9335
rect 15410 9285 15460 9335
rect 15505 9285 15555 9335
rect 15625 9285 15675 9335
rect 15720 9285 15770 9335
rect 15815 9285 15865 9335
rect 15915 9285 15965 9335
rect 16015 9285 16065 9335
rect 16115 9285 16165 9335
rect 16210 9285 16260 9335
rect 16305 9285 16355 9335
rect 16425 9285 16475 9335
rect 16520 9285 16570 9335
rect 16615 9285 16665 9335
rect 16715 9285 16765 9335
rect 16815 9285 16865 9335
rect 16915 9285 16965 9335
rect 17010 9285 17060 9335
rect 17105 9285 17155 9335
rect 17225 9285 17275 9335
rect 17320 9285 17370 9335
rect 17415 9285 17465 9335
rect 17515 9285 17565 9335
rect 17615 9285 17665 9335
rect 17715 9285 17765 9335
rect 17810 9285 17860 9335
rect 17905 9285 17955 9335
rect 9020 9235 9060 9240
rect 9020 9205 9025 9235
rect 9025 9205 9055 9235
rect 9055 9205 9060 9235
rect 9020 9200 9060 9205
rect 9020 9170 9060 9175
rect 9020 9140 9025 9170
rect 9025 9140 9055 9170
rect 9055 9140 9060 9170
rect 9020 9135 9060 9140
rect 14825 9165 14875 9215
rect 14920 9165 14970 9215
rect 15015 9165 15065 9215
rect 15115 9165 15165 9215
rect 15215 9165 15265 9215
rect 15315 9165 15365 9215
rect 15410 9165 15460 9215
rect 15505 9165 15555 9215
rect 15625 9165 15675 9215
rect 15720 9165 15770 9215
rect 15815 9165 15865 9215
rect 15915 9165 15965 9215
rect 16015 9165 16065 9215
rect 16115 9165 16165 9215
rect 16210 9165 16260 9215
rect 16305 9165 16355 9215
rect 16425 9165 16475 9215
rect 16520 9165 16570 9215
rect 16615 9165 16665 9215
rect 16715 9165 16765 9215
rect 16815 9165 16865 9215
rect 16915 9165 16965 9215
rect 17010 9165 17060 9215
rect 17105 9165 17155 9215
rect 17225 9165 17275 9215
rect 17320 9165 17370 9215
rect 17415 9165 17465 9215
rect 17515 9165 17565 9215
rect 17615 9165 17665 9215
rect 17715 9165 17765 9215
rect 17810 9165 17860 9215
rect 17905 9165 17955 9215
rect 9020 9100 9060 9105
rect 9020 9070 9025 9100
rect 9025 9070 9055 9100
rect 9055 9070 9060 9100
rect 9020 9065 9060 9070
rect 9020 9030 9060 9035
rect 9020 9000 9025 9030
rect 9025 9000 9055 9030
rect 9055 9000 9060 9030
rect 9020 8995 9060 9000
rect 9020 8960 9060 8965
rect 9020 8930 9025 8960
rect 9025 8930 9055 8960
rect 9055 8930 9060 8960
rect 9020 8925 9060 8930
rect 14825 9075 14875 9125
rect 14920 9075 14970 9125
rect 15015 9075 15065 9125
rect 15115 9075 15165 9125
rect 15215 9075 15265 9125
rect 15315 9075 15365 9125
rect 15410 9075 15460 9125
rect 15505 9075 15555 9125
rect 15625 9075 15675 9125
rect 15720 9075 15770 9125
rect 15815 9075 15865 9125
rect 15915 9075 15965 9125
rect 16015 9075 16065 9125
rect 16115 9075 16165 9125
rect 16210 9075 16260 9125
rect 16305 9075 16355 9125
rect 16425 9075 16475 9125
rect 16520 9075 16570 9125
rect 16615 9075 16665 9125
rect 16715 9075 16765 9125
rect 16815 9075 16865 9125
rect 16915 9075 16965 9125
rect 17010 9075 17060 9125
rect 17105 9075 17155 9125
rect 17225 9075 17275 9125
rect 17320 9075 17370 9125
rect 17415 9075 17465 9125
rect 17515 9075 17565 9125
rect 17615 9075 17665 9125
rect 17715 9075 17765 9125
rect 17810 9075 17860 9125
rect 17905 9075 17955 9125
rect 14825 8975 14875 9025
rect 14920 8975 14970 9025
rect 15015 8975 15065 9025
rect 15115 8975 15165 9025
rect 15215 8975 15265 9025
rect 15315 8975 15365 9025
rect 15410 8975 15460 9025
rect 15505 8975 15555 9025
rect 15625 8975 15675 9025
rect 15720 8975 15770 9025
rect 15815 8975 15865 9025
rect 15915 8975 15965 9025
rect 16015 8975 16065 9025
rect 16115 8975 16165 9025
rect 16210 8975 16260 9025
rect 16305 8975 16355 9025
rect 16425 8975 16475 9025
rect 16520 8975 16570 9025
rect 16615 8975 16665 9025
rect 16715 8975 16765 9025
rect 16815 8975 16865 9025
rect 16915 8975 16965 9025
rect 17010 8975 17060 9025
rect 17105 8975 17155 9025
rect 17225 8975 17275 9025
rect 17320 8975 17370 9025
rect 17415 8975 17465 9025
rect 17515 8975 17565 9025
rect 17615 8975 17665 9025
rect 17715 8975 17765 9025
rect 17810 8975 17860 9025
rect 17905 8975 17955 9025
rect 9020 8895 9060 8900
rect 9020 8865 9025 8895
rect 9025 8865 9055 8895
rect 9055 8865 9060 8895
rect 9020 8860 9060 8865
rect 9020 8835 9060 8840
rect 9020 8805 9025 8835
rect 9025 8805 9055 8835
rect 9055 8805 9060 8835
rect 9020 8800 9060 8805
rect 14825 8885 14875 8935
rect 14920 8885 14970 8935
rect 15015 8885 15065 8935
rect 15115 8885 15165 8935
rect 15215 8885 15265 8935
rect 15315 8885 15365 8935
rect 15410 8885 15460 8935
rect 15505 8885 15555 8935
rect 15625 8885 15675 8935
rect 15720 8885 15770 8935
rect 15815 8885 15865 8935
rect 15915 8885 15965 8935
rect 16015 8885 16065 8935
rect 16115 8885 16165 8935
rect 16210 8885 16260 8935
rect 16305 8885 16355 8935
rect 16425 8885 16475 8935
rect 16520 8885 16570 8935
rect 16615 8885 16665 8935
rect 16715 8885 16765 8935
rect 16815 8885 16865 8935
rect 16915 8885 16965 8935
rect 17010 8885 17060 8935
rect 17105 8885 17155 8935
rect 17225 8885 17275 8935
rect 17320 8885 17370 8935
rect 17415 8885 17465 8935
rect 17515 8885 17565 8935
rect 17615 8885 17665 8935
rect 17715 8885 17765 8935
rect 17810 8885 17860 8935
rect 17905 8885 17955 8935
rect 9020 8770 9060 8775
rect 9020 8740 9025 8770
rect 9025 8740 9055 8770
rect 9055 8740 9060 8770
rect 9020 8735 9060 8740
rect 9020 8700 9060 8705
rect 9020 8670 9025 8700
rect 9025 8670 9055 8700
rect 9055 8670 9060 8700
rect 9020 8665 9060 8670
rect 9020 8630 9060 8635
rect 9020 8600 9025 8630
rect 9025 8600 9055 8630
rect 9055 8600 9060 8630
rect 9020 8595 9060 8600
rect 9020 8560 9060 8565
rect 9020 8530 9025 8560
rect 9025 8530 9055 8560
rect 9055 8530 9060 8560
rect 9020 8525 9060 8530
rect 14825 8765 14875 8815
rect 14920 8765 14970 8815
rect 15015 8765 15065 8815
rect 15115 8765 15165 8815
rect 15215 8765 15265 8815
rect 15315 8765 15365 8815
rect 15410 8765 15460 8815
rect 15505 8765 15555 8815
rect 15625 8765 15675 8815
rect 15720 8765 15770 8815
rect 15815 8765 15865 8815
rect 15915 8765 15965 8815
rect 16015 8765 16065 8815
rect 16115 8765 16165 8815
rect 16210 8765 16260 8815
rect 16305 8765 16355 8815
rect 16425 8765 16475 8815
rect 16520 8765 16570 8815
rect 16615 8765 16665 8815
rect 16715 8765 16765 8815
rect 16815 8765 16865 8815
rect 16915 8765 16965 8815
rect 17010 8765 17060 8815
rect 17105 8765 17155 8815
rect 17225 8765 17275 8815
rect 17320 8765 17370 8815
rect 17415 8765 17465 8815
rect 17515 8765 17565 8815
rect 17615 8765 17665 8815
rect 17715 8765 17765 8815
rect 17810 8765 17860 8815
rect 17905 8765 17955 8815
rect 14825 8675 14875 8725
rect 14920 8675 14970 8725
rect 15015 8675 15065 8725
rect 15115 8675 15165 8725
rect 15215 8675 15265 8725
rect 15315 8675 15365 8725
rect 15410 8675 15460 8725
rect 15505 8675 15555 8725
rect 15625 8675 15675 8725
rect 15720 8675 15770 8725
rect 15815 8675 15865 8725
rect 15915 8675 15965 8725
rect 16015 8675 16065 8725
rect 16115 8675 16165 8725
rect 16210 8675 16260 8725
rect 16305 8675 16355 8725
rect 16425 8675 16475 8725
rect 16520 8675 16570 8725
rect 16615 8675 16665 8725
rect 16715 8675 16765 8725
rect 16815 8675 16865 8725
rect 16915 8675 16965 8725
rect 17010 8675 17060 8725
rect 17105 8675 17155 8725
rect 17225 8675 17275 8725
rect 17320 8675 17370 8725
rect 17415 8675 17465 8725
rect 17515 8675 17565 8725
rect 17615 8675 17665 8725
rect 17715 8675 17765 8725
rect 17810 8675 17860 8725
rect 17905 8675 17955 8725
rect 14825 8575 14875 8625
rect 14920 8575 14970 8625
rect 15015 8575 15065 8625
rect 15115 8575 15165 8625
rect 15215 8575 15265 8625
rect 15315 8575 15365 8625
rect 15410 8575 15460 8625
rect 15505 8575 15555 8625
rect 15625 8575 15675 8625
rect 15720 8575 15770 8625
rect 15815 8575 15865 8625
rect 15915 8575 15965 8625
rect 16015 8575 16065 8625
rect 16115 8575 16165 8625
rect 16210 8575 16260 8625
rect 16305 8575 16355 8625
rect 16425 8575 16475 8625
rect 16520 8575 16570 8625
rect 16615 8575 16665 8625
rect 16715 8575 16765 8625
rect 16815 8575 16865 8625
rect 16915 8575 16965 8625
rect 17010 8575 17060 8625
rect 17105 8575 17155 8625
rect 17225 8575 17275 8625
rect 17320 8575 17370 8625
rect 17415 8575 17465 8625
rect 17515 8575 17565 8625
rect 17615 8575 17665 8625
rect 17715 8575 17765 8625
rect 17810 8575 17860 8625
rect 17905 8575 17955 8625
rect 9020 8495 9060 8500
rect 9020 8465 9025 8495
rect 9025 8465 9055 8495
rect 9055 8465 9060 8495
rect 9020 8460 9060 8465
rect 9020 8435 9060 8440
rect 9020 8405 9025 8435
rect 9025 8405 9055 8435
rect 9055 8405 9060 8435
rect 9020 8400 9060 8405
rect 14825 8485 14875 8535
rect 14920 8485 14970 8535
rect 15015 8485 15065 8535
rect 15115 8485 15165 8535
rect 15215 8485 15265 8535
rect 15315 8485 15365 8535
rect 15410 8485 15460 8535
rect 15505 8485 15555 8535
rect 15625 8485 15675 8535
rect 15720 8485 15770 8535
rect 15815 8485 15865 8535
rect 15915 8485 15965 8535
rect 16015 8485 16065 8535
rect 16115 8485 16165 8535
rect 16210 8485 16260 8535
rect 16305 8485 16355 8535
rect 16425 8485 16475 8535
rect 16520 8485 16570 8535
rect 16615 8485 16665 8535
rect 16715 8485 16765 8535
rect 16815 8485 16865 8535
rect 16915 8485 16965 8535
rect 17010 8485 17060 8535
rect 17105 8485 17155 8535
rect 17225 8485 17275 8535
rect 17320 8485 17370 8535
rect 17415 8485 17465 8535
rect 17515 8485 17565 8535
rect 17615 8485 17665 8535
rect 17715 8485 17765 8535
rect 17810 8485 17860 8535
rect 17905 8485 17955 8535
rect 9020 8370 9060 8375
rect 9020 8340 9025 8370
rect 9025 8340 9055 8370
rect 9055 8340 9060 8370
rect 9020 8335 9060 8340
rect 9020 8300 9060 8305
rect 9020 8270 9025 8300
rect 9025 8270 9055 8300
rect 9055 8270 9060 8300
rect 9020 8265 9060 8270
rect 9020 8230 9060 8235
rect 9020 8200 9025 8230
rect 9025 8200 9055 8230
rect 9055 8200 9060 8230
rect 9020 8195 9060 8200
rect 14825 8365 14875 8415
rect 14920 8365 14970 8415
rect 15015 8365 15065 8415
rect 15115 8365 15165 8415
rect 15215 8365 15265 8415
rect 15315 8365 15365 8415
rect 15410 8365 15460 8415
rect 15505 8365 15555 8415
rect 15625 8365 15675 8415
rect 15720 8365 15770 8415
rect 15815 8365 15865 8415
rect 15915 8365 15965 8415
rect 16015 8365 16065 8415
rect 16115 8365 16165 8415
rect 16210 8365 16260 8415
rect 16305 8365 16355 8415
rect 16425 8365 16475 8415
rect 16520 8365 16570 8415
rect 16615 8365 16665 8415
rect 16715 8365 16765 8415
rect 16815 8365 16865 8415
rect 16915 8365 16965 8415
rect 17010 8365 17060 8415
rect 17105 8365 17155 8415
rect 17225 8365 17275 8415
rect 17320 8365 17370 8415
rect 17415 8365 17465 8415
rect 17515 8365 17565 8415
rect 17615 8365 17665 8415
rect 17715 8365 17765 8415
rect 17810 8365 17860 8415
rect 17905 8365 17955 8415
rect 14825 8275 14875 8325
rect 14920 8275 14970 8325
rect 15015 8275 15065 8325
rect 15115 8275 15165 8325
rect 15215 8275 15265 8325
rect 15315 8275 15365 8325
rect 15410 8275 15460 8325
rect 15505 8275 15555 8325
rect 15625 8275 15675 8325
rect 15720 8275 15770 8325
rect 15815 8275 15865 8325
rect 15915 8275 15965 8325
rect 16015 8275 16065 8325
rect 16115 8275 16165 8325
rect 16210 8275 16260 8325
rect 16305 8275 16355 8325
rect 16425 8275 16475 8325
rect 16520 8275 16570 8325
rect 16615 8275 16665 8325
rect 16715 8275 16765 8325
rect 16815 8275 16865 8325
rect 16915 8275 16965 8325
rect 17010 8275 17060 8325
rect 17105 8275 17155 8325
rect 17225 8275 17275 8325
rect 17320 8275 17370 8325
rect 17415 8275 17465 8325
rect 17515 8275 17565 8325
rect 17615 8275 17665 8325
rect 17715 8275 17765 8325
rect 17810 8275 17860 8325
rect 17905 8275 17955 8325
rect 9020 8160 9060 8165
rect 9020 8130 9025 8160
rect 9025 8130 9055 8160
rect 9055 8130 9060 8160
rect 9020 8125 9060 8130
rect 9020 8095 9060 8100
rect 9020 8065 9025 8095
rect 9025 8065 9055 8095
rect 9055 8065 9060 8095
rect 9020 8060 9060 8065
rect 14825 8175 14875 8225
rect 14920 8175 14970 8225
rect 15015 8175 15065 8225
rect 15115 8175 15165 8225
rect 15215 8175 15265 8225
rect 15315 8175 15365 8225
rect 15410 8175 15460 8225
rect 15505 8175 15555 8225
rect 15625 8175 15675 8225
rect 15720 8175 15770 8225
rect 15815 8175 15865 8225
rect 15915 8175 15965 8225
rect 16015 8175 16065 8225
rect 16115 8175 16165 8225
rect 16210 8175 16260 8225
rect 16305 8175 16355 8225
rect 16425 8175 16475 8225
rect 16520 8175 16570 8225
rect 16615 8175 16665 8225
rect 16715 8175 16765 8225
rect 16815 8175 16865 8225
rect 16915 8175 16965 8225
rect 17010 8175 17060 8225
rect 17105 8175 17155 8225
rect 17225 8175 17275 8225
rect 17320 8175 17370 8225
rect 17415 8175 17465 8225
rect 17515 8175 17565 8225
rect 17615 8175 17665 8225
rect 17715 8175 17765 8225
rect 17810 8175 17860 8225
rect 17905 8175 17955 8225
rect 14825 8085 14875 8135
rect 14920 8085 14970 8135
rect 15015 8085 15065 8135
rect 15115 8085 15165 8135
rect 15215 8085 15265 8135
rect 15315 8085 15365 8135
rect 15410 8085 15460 8135
rect 15505 8085 15555 8135
rect 15625 8085 15675 8135
rect 15720 8085 15770 8135
rect 15815 8085 15865 8135
rect 15915 8085 15965 8135
rect 16015 8085 16065 8135
rect 16115 8085 16165 8135
rect 16210 8085 16260 8135
rect 16305 8085 16355 8135
rect 16425 8085 16475 8135
rect 16520 8085 16570 8135
rect 16615 8085 16665 8135
rect 16715 8085 16765 8135
rect 16815 8085 16865 8135
rect 16915 8085 16965 8135
rect 17010 8085 17060 8135
rect 17105 8085 17155 8135
rect 17225 8085 17275 8135
rect 17320 8085 17370 8135
rect 17415 8085 17465 8135
rect 17515 8085 17565 8135
rect 17615 8085 17665 8135
rect 17715 8085 17765 8135
rect 17810 8085 17860 8135
rect 17905 8085 17955 8135
rect 9020 8035 9060 8040
rect 9020 8005 9025 8035
rect 9025 8005 9055 8035
rect 9055 8005 9060 8035
rect 9020 8000 9060 8005
rect 9020 7970 9060 7975
rect 9020 7940 9025 7970
rect 9025 7940 9055 7970
rect 9055 7940 9060 7970
rect 9020 7935 9060 7940
rect 9020 7900 9060 7905
rect 9020 7870 9025 7900
rect 9025 7870 9055 7900
rect 9055 7870 9060 7900
rect 9020 7865 9060 7870
rect 14825 7965 14875 8015
rect 14920 7965 14970 8015
rect 15015 7965 15065 8015
rect 15115 7965 15165 8015
rect 15215 7965 15265 8015
rect 15315 7965 15365 8015
rect 15410 7965 15460 8015
rect 15505 7965 15555 8015
rect 15625 7965 15675 8015
rect 15720 7965 15770 8015
rect 15815 7965 15865 8015
rect 15915 7965 15965 8015
rect 16015 7965 16065 8015
rect 16115 7965 16165 8015
rect 16210 7965 16260 8015
rect 16305 7965 16355 8015
rect 16425 7965 16475 8015
rect 16520 7965 16570 8015
rect 16615 7965 16665 8015
rect 16715 7965 16765 8015
rect 16815 7965 16865 8015
rect 16915 7965 16965 8015
rect 17010 7965 17060 8015
rect 17105 7965 17155 8015
rect 17225 7965 17275 8015
rect 17320 7965 17370 8015
rect 17415 7965 17465 8015
rect 17515 7965 17565 8015
rect 17615 7965 17665 8015
rect 17715 7965 17765 8015
rect 17810 7965 17860 8015
rect 17905 7965 17955 8015
rect 14825 7875 14875 7925
rect 14920 7875 14970 7925
rect 15015 7875 15065 7925
rect 15115 7875 15165 7925
rect 15215 7875 15265 7925
rect 15315 7875 15365 7925
rect 15410 7875 15460 7925
rect 15505 7875 15555 7925
rect 15625 7875 15675 7925
rect 15720 7875 15770 7925
rect 15815 7875 15865 7925
rect 15915 7875 15965 7925
rect 16015 7875 16065 7925
rect 16115 7875 16165 7925
rect 16210 7875 16260 7925
rect 16305 7875 16355 7925
rect 16425 7875 16475 7925
rect 16520 7875 16570 7925
rect 16615 7875 16665 7925
rect 16715 7875 16765 7925
rect 16815 7875 16865 7925
rect 16915 7875 16965 7925
rect 17010 7875 17060 7925
rect 17105 7875 17155 7925
rect 17225 7875 17275 7925
rect 17320 7875 17370 7925
rect 17415 7875 17465 7925
rect 17515 7875 17565 7925
rect 17615 7875 17665 7925
rect 17715 7875 17765 7925
rect 17810 7875 17860 7925
rect 17905 7875 17955 7925
rect 9020 7830 9060 7835
rect 9020 7800 9025 7830
rect 9025 7800 9055 7830
rect 9055 7800 9060 7830
rect 9020 7795 9060 7800
rect 9020 7760 9060 7765
rect 9020 7730 9025 7760
rect 9025 7730 9055 7760
rect 9055 7730 9060 7760
rect 9020 7725 9060 7730
rect 14825 7775 14875 7825
rect 14920 7775 14970 7825
rect 15015 7775 15065 7825
rect 15115 7775 15165 7825
rect 15215 7775 15265 7825
rect 15315 7775 15365 7825
rect 15410 7775 15460 7825
rect 15505 7775 15555 7825
rect 15625 7775 15675 7825
rect 15720 7775 15770 7825
rect 15815 7775 15865 7825
rect 15915 7775 15965 7825
rect 16015 7775 16065 7825
rect 16115 7775 16165 7825
rect 16210 7775 16260 7825
rect 16305 7775 16355 7825
rect 16425 7775 16475 7825
rect 16520 7775 16570 7825
rect 16615 7775 16665 7825
rect 16715 7775 16765 7825
rect 16815 7775 16865 7825
rect 16915 7775 16965 7825
rect 17010 7775 17060 7825
rect 17105 7775 17155 7825
rect 17225 7775 17275 7825
rect 17320 7775 17370 7825
rect 17415 7775 17465 7825
rect 17515 7775 17565 7825
rect 17615 7775 17665 7825
rect 17715 7775 17765 7825
rect 17810 7775 17860 7825
rect 17905 7775 17955 7825
rect 9020 7695 9060 7700
rect 9020 7665 9025 7695
rect 9025 7665 9055 7695
rect 9055 7665 9060 7695
rect 9020 7660 9060 7665
rect 9020 7635 9060 7640
rect 9020 7605 9025 7635
rect 9025 7605 9055 7635
rect 9055 7605 9060 7635
rect 9020 7600 9060 7605
rect 9020 7570 9060 7575
rect 9020 7540 9025 7570
rect 9025 7540 9055 7570
rect 9055 7540 9060 7570
rect 9020 7535 9060 7540
rect 9020 7500 9060 7505
rect 9020 7470 9025 7500
rect 9025 7470 9055 7500
rect 9055 7470 9060 7500
rect 9020 7465 9060 7470
rect 14825 7685 14875 7735
rect 14920 7685 14970 7735
rect 15015 7685 15065 7735
rect 15115 7685 15165 7735
rect 15215 7685 15265 7735
rect 15315 7685 15365 7735
rect 15410 7685 15460 7735
rect 15505 7685 15555 7735
rect 15625 7685 15675 7735
rect 15720 7685 15770 7735
rect 15815 7685 15865 7735
rect 15915 7685 15965 7735
rect 16015 7685 16065 7735
rect 16115 7685 16165 7735
rect 16210 7685 16260 7735
rect 16305 7685 16355 7735
rect 16425 7685 16475 7735
rect 16520 7685 16570 7735
rect 16615 7685 16665 7735
rect 16715 7685 16765 7735
rect 16815 7685 16865 7735
rect 16915 7685 16965 7735
rect 17010 7685 17060 7735
rect 17105 7685 17155 7735
rect 17225 7685 17275 7735
rect 17320 7685 17370 7735
rect 17415 7685 17465 7735
rect 17515 7685 17565 7735
rect 17615 7685 17665 7735
rect 17715 7685 17765 7735
rect 17810 7685 17860 7735
rect 17905 7685 17955 7735
rect 14825 7565 14875 7615
rect 14920 7565 14970 7615
rect 15015 7565 15065 7615
rect 15115 7565 15165 7615
rect 15215 7565 15265 7615
rect 15315 7565 15365 7615
rect 15410 7565 15460 7615
rect 15505 7565 15555 7615
rect 15625 7565 15675 7615
rect 15720 7565 15770 7615
rect 15815 7565 15865 7615
rect 15915 7565 15965 7615
rect 16015 7565 16065 7615
rect 16115 7565 16165 7615
rect 16210 7565 16260 7615
rect 16305 7565 16355 7615
rect 16425 7565 16475 7615
rect 16520 7565 16570 7615
rect 16615 7565 16665 7615
rect 16715 7565 16765 7615
rect 16815 7565 16865 7615
rect 16915 7565 16965 7615
rect 17010 7565 17060 7615
rect 17105 7565 17155 7615
rect 17225 7565 17275 7615
rect 17320 7565 17370 7615
rect 17415 7565 17465 7615
rect 17515 7565 17565 7615
rect 17615 7565 17665 7615
rect 17715 7565 17765 7615
rect 17810 7565 17860 7615
rect 17905 7565 17955 7615
rect 9020 7430 9060 7435
rect 9020 7400 9025 7430
rect 9025 7400 9055 7430
rect 9055 7400 9060 7430
rect 9020 7395 9060 7400
rect 14825 7475 14875 7525
rect 14920 7475 14970 7525
rect 15015 7475 15065 7525
rect 15115 7475 15165 7525
rect 15215 7475 15265 7525
rect 15315 7475 15365 7525
rect 15410 7475 15460 7525
rect 15505 7475 15555 7525
rect 15625 7475 15675 7525
rect 15720 7475 15770 7525
rect 15815 7475 15865 7525
rect 15915 7475 15965 7525
rect 16015 7475 16065 7525
rect 16115 7475 16165 7525
rect 16210 7475 16260 7525
rect 16305 7475 16355 7525
rect 16425 7475 16475 7525
rect 16520 7475 16570 7525
rect 16615 7475 16665 7525
rect 16715 7475 16765 7525
rect 16815 7475 16865 7525
rect 16915 7475 16965 7525
rect 17010 7475 17060 7525
rect 17105 7475 17155 7525
rect 17225 7475 17275 7525
rect 17320 7475 17370 7525
rect 17415 7475 17465 7525
rect 17515 7475 17565 7525
rect 17615 7475 17665 7525
rect 17715 7475 17765 7525
rect 17810 7475 17860 7525
rect 17905 7475 17955 7525
rect 9020 7360 9060 7365
rect 9020 7330 9025 7360
rect 9025 7330 9055 7360
rect 9055 7330 9060 7360
rect 9020 7325 9060 7330
rect 9020 7295 9060 7300
rect 9020 7265 9025 7295
rect 9025 7265 9055 7295
rect 9055 7265 9060 7295
rect 9020 7260 9060 7265
rect 9020 7235 9060 7240
rect 9020 7205 9025 7235
rect 9025 7205 9055 7235
rect 9055 7205 9060 7235
rect 9020 7200 9060 7205
rect 9020 7170 9060 7175
rect 9020 7140 9025 7170
rect 9025 7140 9055 7170
rect 9055 7140 9060 7170
rect 9020 7135 9060 7140
rect 14825 7375 14875 7425
rect 14920 7375 14970 7425
rect 15015 7375 15065 7425
rect 15115 7375 15165 7425
rect 15215 7375 15265 7425
rect 15315 7375 15365 7425
rect 15410 7375 15460 7425
rect 15505 7375 15555 7425
rect 15625 7375 15675 7425
rect 15720 7375 15770 7425
rect 15815 7375 15865 7425
rect 15915 7375 15965 7425
rect 16015 7375 16065 7425
rect 16115 7375 16165 7425
rect 16210 7375 16260 7425
rect 16305 7375 16355 7425
rect 16425 7375 16475 7425
rect 16520 7375 16570 7425
rect 16615 7375 16665 7425
rect 16715 7375 16765 7425
rect 16815 7375 16865 7425
rect 16915 7375 16965 7425
rect 17010 7375 17060 7425
rect 17105 7375 17155 7425
rect 17225 7375 17275 7425
rect 17320 7375 17370 7425
rect 17415 7375 17465 7425
rect 17515 7375 17565 7425
rect 17615 7375 17665 7425
rect 17715 7375 17765 7425
rect 17810 7375 17860 7425
rect 17905 7375 17955 7425
rect 14825 7285 14875 7335
rect 14920 7285 14970 7335
rect 15015 7285 15065 7335
rect 15115 7285 15165 7335
rect 15215 7285 15265 7335
rect 15315 7285 15365 7335
rect 15410 7285 15460 7335
rect 15505 7285 15555 7335
rect 15625 7285 15675 7335
rect 15720 7285 15770 7335
rect 15815 7285 15865 7335
rect 15915 7285 15965 7335
rect 16015 7285 16065 7335
rect 16115 7285 16165 7335
rect 16210 7285 16260 7335
rect 16305 7285 16355 7335
rect 16425 7285 16475 7335
rect 16520 7285 16570 7335
rect 16615 7285 16665 7335
rect 16715 7285 16765 7335
rect 16815 7285 16865 7335
rect 16915 7285 16965 7335
rect 17010 7285 17060 7335
rect 17105 7285 17155 7335
rect 17225 7285 17275 7335
rect 17320 7285 17370 7335
rect 17415 7285 17465 7335
rect 17515 7285 17565 7335
rect 17615 7285 17665 7335
rect 17715 7285 17765 7335
rect 17810 7285 17860 7335
rect 17905 7285 17955 7335
rect 14825 7165 14875 7215
rect 14920 7165 14970 7215
rect 15015 7165 15065 7215
rect 15115 7165 15165 7215
rect 15215 7165 15265 7215
rect 15315 7165 15365 7215
rect 15410 7165 15460 7215
rect 15505 7165 15555 7215
rect 15625 7165 15675 7215
rect 15720 7165 15770 7215
rect 15815 7165 15865 7215
rect 15915 7165 15965 7215
rect 16015 7165 16065 7215
rect 16115 7165 16165 7215
rect 16210 7165 16260 7215
rect 16305 7165 16355 7215
rect 16425 7165 16475 7215
rect 16520 7165 16570 7215
rect 16615 7165 16665 7215
rect 16715 7165 16765 7215
rect 16815 7165 16865 7215
rect 16915 7165 16965 7215
rect 17010 7165 17060 7215
rect 17105 7165 17155 7215
rect 17225 7165 17275 7215
rect 17320 7165 17370 7215
rect 17415 7165 17465 7215
rect 17515 7165 17565 7215
rect 17615 7165 17665 7215
rect 17715 7165 17765 7215
rect 17810 7165 17860 7215
rect 17905 7165 17955 7215
rect 9020 7100 9060 7105
rect 9020 7070 9025 7100
rect 9025 7070 9055 7100
rect 9055 7070 9060 7100
rect 9020 7065 9060 7070
rect 9020 7030 9060 7035
rect 9020 7000 9025 7030
rect 9025 7000 9055 7030
rect 9055 7000 9060 7030
rect 9020 6995 9060 7000
rect 14825 7075 14875 7125
rect 14920 7075 14970 7125
rect 15015 7075 15065 7125
rect 15115 7075 15165 7125
rect 15215 7075 15265 7125
rect 15315 7075 15365 7125
rect 15410 7075 15460 7125
rect 15505 7075 15555 7125
rect 15625 7075 15675 7125
rect 15720 7075 15770 7125
rect 15815 7075 15865 7125
rect 15915 7075 15965 7125
rect 16015 7075 16065 7125
rect 16115 7075 16165 7125
rect 16210 7075 16260 7125
rect 16305 7075 16355 7125
rect 16425 7075 16475 7125
rect 16520 7075 16570 7125
rect 16615 7075 16665 7125
rect 16715 7075 16765 7125
rect 16815 7075 16865 7125
rect 16915 7075 16965 7125
rect 17010 7075 17060 7125
rect 17105 7075 17155 7125
rect 17225 7075 17275 7125
rect 17320 7075 17370 7125
rect 17415 7075 17465 7125
rect 17515 7075 17565 7125
rect 17615 7075 17665 7125
rect 17715 7075 17765 7125
rect 17810 7075 17860 7125
rect 17905 7075 17955 7125
rect 9020 6960 9060 6965
rect 9020 6930 9025 6960
rect 9025 6930 9055 6960
rect 9055 6930 9060 6960
rect 9020 6925 9060 6930
rect 9020 6895 9060 6900
rect 9020 6865 9025 6895
rect 9025 6865 9055 6895
rect 9055 6865 9060 6895
rect 9020 6860 9060 6865
rect 9020 6835 9060 6840
rect 9020 6805 9025 6835
rect 9025 6805 9055 6835
rect 9055 6805 9060 6835
rect 9020 6800 9060 6805
rect 14825 6975 14875 7025
rect 14920 6975 14970 7025
rect 15015 6975 15065 7025
rect 15115 6975 15165 7025
rect 15215 6975 15265 7025
rect 15315 6975 15365 7025
rect 15410 6975 15460 7025
rect 15505 6975 15555 7025
rect 15625 6975 15675 7025
rect 15720 6975 15770 7025
rect 15815 6975 15865 7025
rect 15915 6975 15965 7025
rect 16015 6975 16065 7025
rect 16115 6975 16165 7025
rect 16210 6975 16260 7025
rect 16305 6975 16355 7025
rect 16425 6975 16475 7025
rect 16520 6975 16570 7025
rect 16615 6975 16665 7025
rect 16715 6975 16765 7025
rect 16815 6975 16865 7025
rect 16915 6975 16965 7025
rect 17010 6975 17060 7025
rect 17105 6975 17155 7025
rect 17225 6975 17275 7025
rect 17320 6975 17370 7025
rect 17415 6975 17465 7025
rect 17515 6975 17565 7025
rect 17615 6975 17665 7025
rect 17715 6975 17765 7025
rect 17810 6975 17860 7025
rect 17905 6975 17955 7025
rect 14825 6885 14875 6935
rect 14920 6885 14970 6935
rect 15015 6885 15065 6935
rect 15115 6885 15165 6935
rect 15215 6885 15265 6935
rect 15315 6885 15365 6935
rect 15410 6885 15460 6935
rect 15505 6885 15555 6935
rect 15625 6885 15675 6935
rect 15720 6885 15770 6935
rect 15815 6885 15865 6935
rect 15915 6885 15965 6935
rect 16015 6885 16065 6935
rect 16115 6885 16165 6935
rect 16210 6885 16260 6935
rect 16305 6885 16355 6935
rect 16425 6885 16475 6935
rect 16520 6885 16570 6935
rect 16615 6885 16665 6935
rect 16715 6885 16765 6935
rect 16815 6885 16865 6935
rect 16915 6885 16965 6935
rect 17010 6885 17060 6935
rect 17105 6885 17155 6935
rect 17225 6885 17275 6935
rect 17320 6885 17370 6935
rect 17415 6885 17465 6935
rect 17515 6885 17565 6935
rect 17615 6885 17665 6935
rect 17715 6885 17765 6935
rect 17810 6885 17860 6935
rect 17905 6885 17955 6935
rect 9020 6770 9060 6775
rect 9020 6740 9025 6770
rect 9025 6740 9055 6770
rect 9055 6740 9060 6770
rect 9020 6735 9060 6740
rect 9020 6700 9060 6705
rect 9020 6670 9025 6700
rect 9025 6670 9055 6700
rect 9055 6670 9060 6700
rect 9020 6665 9060 6670
rect 14825 6765 14875 6815
rect 14920 6765 14970 6815
rect 15015 6765 15065 6815
rect 15115 6765 15165 6815
rect 15215 6765 15265 6815
rect 15315 6765 15365 6815
rect 15410 6765 15460 6815
rect 15505 6765 15555 6815
rect 15625 6765 15675 6815
rect 15720 6765 15770 6815
rect 15815 6765 15865 6815
rect 15915 6765 15965 6815
rect 16015 6765 16065 6815
rect 16115 6765 16165 6815
rect 16210 6765 16260 6815
rect 16305 6765 16355 6815
rect 16425 6765 16475 6815
rect 16520 6765 16570 6815
rect 16615 6765 16665 6815
rect 16715 6765 16765 6815
rect 16815 6765 16865 6815
rect 16915 6765 16965 6815
rect 17010 6765 17060 6815
rect 17105 6765 17155 6815
rect 17225 6765 17275 6815
rect 17320 6765 17370 6815
rect 17415 6765 17465 6815
rect 17515 6765 17565 6815
rect 17615 6765 17665 6815
rect 17715 6765 17765 6815
rect 17810 6765 17860 6815
rect 17905 6765 17955 6815
rect 9020 6630 9060 6635
rect 9020 6600 9025 6630
rect 9025 6600 9055 6630
rect 9055 6600 9060 6630
rect 9020 6595 9060 6600
rect 9020 6560 9060 6565
rect 9020 6530 9025 6560
rect 9025 6530 9055 6560
rect 9055 6530 9060 6560
rect 9020 6525 9060 6530
rect 9020 6495 9060 6500
rect 9020 6465 9025 6495
rect 9025 6465 9055 6495
rect 9055 6465 9060 6495
rect 9020 6460 9060 6465
rect 14825 6675 14875 6725
rect 14920 6675 14970 6725
rect 15015 6675 15065 6725
rect 15115 6675 15165 6725
rect 15215 6675 15265 6725
rect 15315 6675 15365 6725
rect 15410 6675 15460 6725
rect 15505 6675 15555 6725
rect 15625 6675 15675 6725
rect 15720 6675 15770 6725
rect 15815 6675 15865 6725
rect 15915 6675 15965 6725
rect 16015 6675 16065 6725
rect 16115 6675 16165 6725
rect 16210 6675 16260 6725
rect 16305 6675 16355 6725
rect 16425 6675 16475 6725
rect 16520 6675 16570 6725
rect 16615 6675 16665 6725
rect 16715 6675 16765 6725
rect 16815 6675 16865 6725
rect 16915 6675 16965 6725
rect 17010 6675 17060 6725
rect 17105 6675 17155 6725
rect 17225 6675 17275 6725
rect 17320 6675 17370 6725
rect 17415 6675 17465 6725
rect 17515 6675 17565 6725
rect 17615 6675 17665 6725
rect 17715 6675 17765 6725
rect 17810 6675 17860 6725
rect 17905 6675 17955 6725
rect 14825 6575 14875 6625
rect 14920 6575 14970 6625
rect 15015 6575 15065 6625
rect 15115 6575 15165 6625
rect 15215 6575 15265 6625
rect 15315 6575 15365 6625
rect 15410 6575 15460 6625
rect 15505 6575 15555 6625
rect 15625 6575 15675 6625
rect 15720 6575 15770 6625
rect 15815 6575 15865 6625
rect 15915 6575 15965 6625
rect 16015 6575 16065 6625
rect 16115 6575 16165 6625
rect 16210 6575 16260 6625
rect 16305 6575 16355 6625
rect 16425 6575 16475 6625
rect 16520 6575 16570 6625
rect 16615 6575 16665 6625
rect 16715 6575 16765 6625
rect 16815 6575 16865 6625
rect 16915 6575 16965 6625
rect 17010 6575 17060 6625
rect 17105 6575 17155 6625
rect 17225 6575 17275 6625
rect 17320 6575 17370 6625
rect 17415 6575 17465 6625
rect 17515 6575 17565 6625
rect 17615 6575 17665 6625
rect 17715 6575 17765 6625
rect 17810 6575 17860 6625
rect 17905 6575 17955 6625
rect 14825 6485 14875 6535
rect 14920 6485 14970 6535
rect 15015 6485 15065 6535
rect 15115 6485 15165 6535
rect 15215 6485 15265 6535
rect 15315 6485 15365 6535
rect 15410 6485 15460 6535
rect 15505 6485 15555 6535
rect 15625 6485 15675 6535
rect 15720 6485 15770 6535
rect 15815 6485 15865 6535
rect 15915 6485 15965 6535
rect 16015 6485 16065 6535
rect 16115 6485 16165 6535
rect 16210 6485 16260 6535
rect 16305 6485 16355 6535
rect 16425 6485 16475 6535
rect 16520 6485 16570 6535
rect 16615 6485 16665 6535
rect 16715 6485 16765 6535
rect 16815 6485 16865 6535
rect 16915 6485 16965 6535
rect 17010 6485 17060 6535
rect 17105 6485 17155 6535
rect 17225 6485 17275 6535
rect 17320 6485 17370 6535
rect 17415 6485 17465 6535
rect 17515 6485 17565 6535
rect 17615 6485 17665 6535
rect 17715 6485 17765 6535
rect 17810 6485 17860 6535
rect 17905 6485 17955 6535
rect -80 -1305 -40 -1300
rect -80 -1335 -75 -1305
rect -75 -1335 -45 -1305
rect -45 -1335 -40 -1305
rect -80 -1340 -40 -1335
rect -80 -1370 -40 -1365
rect -80 -1400 -75 -1370
rect -75 -1400 -45 -1370
rect -45 -1400 -40 -1370
rect -80 -1405 -40 -1400
rect -80 -1440 -40 -1435
rect -80 -1470 -75 -1440
rect -75 -1470 -45 -1440
rect -45 -1470 -40 -1440
rect -80 -1475 -40 -1470
rect -80 -1510 -40 -1505
rect -80 -1540 -75 -1510
rect -75 -1540 -45 -1510
rect -45 -1540 -40 -1510
rect -80 -1545 -40 -1540
rect -80 -1580 -40 -1575
rect -80 -1610 -75 -1580
rect -75 -1610 -45 -1580
rect -45 -1610 -40 -1580
rect -80 -1615 -40 -1610
rect -80 -1645 -40 -1640
rect -80 -1675 -75 -1645
rect -75 -1675 -45 -1645
rect -45 -1675 -40 -1645
rect -80 -1680 -40 -1675
rect -80 -1705 -40 -1700
rect -80 -1735 -75 -1705
rect -75 -1735 -45 -1705
rect -45 -1735 -40 -1705
rect -80 -1740 -40 -1735
rect -80 -1770 -40 -1765
rect -80 -1800 -75 -1770
rect -75 -1800 -45 -1770
rect -45 -1800 -40 -1770
rect -80 -1805 -40 -1800
rect -80 -1840 -40 -1835
rect -80 -1870 -75 -1840
rect -75 -1870 -45 -1840
rect -45 -1870 -40 -1840
rect -80 -1875 -40 -1870
rect -80 -1910 -40 -1905
rect -80 -1940 -75 -1910
rect -75 -1940 -45 -1910
rect -45 -1940 -40 -1910
rect -80 -1945 -40 -1940
rect -80 -1980 -40 -1975
rect -80 -2010 -75 -1980
rect -75 -2010 -45 -1980
rect -45 -2010 -40 -1980
rect -80 -2015 -40 -2010
rect -80 -2045 -40 -2040
rect -80 -2075 -75 -2045
rect -75 -2075 -45 -2045
rect -45 -2075 -40 -2045
rect -80 -2080 -40 -2075
rect -80 -2105 -40 -2100
rect -80 -2135 -75 -2105
rect -75 -2135 -45 -2105
rect -45 -2135 -40 -2105
rect -80 -2140 -40 -2135
rect -80 -2170 -40 -2165
rect -80 -2200 -75 -2170
rect -75 -2200 -45 -2170
rect -45 -2200 -40 -2170
rect -80 -2205 -40 -2200
rect -80 -2240 -40 -2235
rect -80 -2270 -75 -2240
rect -75 -2270 -45 -2240
rect -45 -2270 -40 -2240
rect -80 -2275 -40 -2270
rect -80 -2310 -40 -2305
rect -80 -2340 -75 -2310
rect -75 -2340 -45 -2310
rect -45 -2340 -40 -2310
rect -80 -2345 -40 -2340
rect -80 -2380 -40 -2375
rect -80 -2410 -75 -2380
rect -75 -2410 -45 -2380
rect -45 -2410 -40 -2380
rect -80 -2415 -40 -2410
rect -80 -2445 -40 -2440
rect -80 -2475 -75 -2445
rect -75 -2475 -45 -2445
rect -45 -2475 -40 -2445
rect -80 -2480 -40 -2475
rect -80 -2505 -40 -2500
rect -80 -2535 -75 -2505
rect -75 -2535 -45 -2505
rect -45 -2535 -40 -2505
rect -80 -2540 -40 -2535
rect -80 -2570 -40 -2565
rect -80 -2600 -75 -2570
rect -75 -2600 -45 -2570
rect -45 -2600 -40 -2570
rect -80 -2605 -40 -2600
rect -80 -2640 -40 -2635
rect -80 -2670 -75 -2640
rect -75 -2670 -45 -2640
rect -45 -2670 -40 -2640
rect -80 -2675 -40 -2670
rect -80 -2710 -40 -2705
rect -80 -2740 -75 -2710
rect -75 -2740 -45 -2710
rect -45 -2740 -40 -2710
rect -80 -2745 -40 -2740
rect -80 -2780 -40 -2775
rect -80 -2810 -75 -2780
rect -75 -2810 -45 -2780
rect -45 -2810 -40 -2780
rect -80 -2815 -40 -2810
rect -80 -2845 -40 -2840
rect -80 -2875 -75 -2845
rect -75 -2875 -45 -2845
rect -45 -2875 -40 -2845
rect -80 -2880 -40 -2875
rect -80 -2905 -40 -2900
rect -80 -2935 -75 -2905
rect -75 -2935 -45 -2905
rect -45 -2935 -40 -2905
rect -80 -2940 -40 -2935
rect -80 -2970 -40 -2965
rect -80 -3000 -75 -2970
rect -75 -3000 -45 -2970
rect -45 -3000 -40 -2970
rect -80 -3005 -40 -3000
rect -80 -3040 -40 -3035
rect -80 -3070 -75 -3040
rect -75 -3070 -45 -3040
rect -45 -3070 -40 -3040
rect -80 -3075 -40 -3070
rect -80 -3110 -40 -3105
rect -80 -3140 -75 -3110
rect -75 -3140 -45 -3110
rect -45 -3140 -40 -3110
rect -80 -3145 -40 -3140
rect -80 -3180 -40 -3175
rect -80 -3210 -75 -3180
rect -75 -3210 -45 -3180
rect -45 -3210 -40 -3180
rect -80 -3215 -40 -3210
rect -80 -3245 -40 -3240
rect -80 -3275 -75 -3245
rect -75 -3275 -45 -3245
rect -45 -3275 -40 -3245
rect -80 -3280 -40 -3275
rect -80 -3305 -40 -3300
rect -80 -3335 -75 -3305
rect -75 -3335 -45 -3305
rect -45 -3335 -40 -3305
rect -80 -3340 -40 -3335
rect -80 -3370 -40 -3365
rect -80 -3400 -75 -3370
rect -75 -3400 -45 -3370
rect -45 -3400 -40 -3370
rect -80 -3405 -40 -3400
rect -80 -3440 -40 -3435
rect -80 -3470 -75 -3440
rect -75 -3470 -45 -3440
rect -45 -3470 -40 -3440
rect -80 -3475 -40 -3470
rect -80 -3510 -40 -3505
rect -80 -3540 -75 -3510
rect -75 -3540 -45 -3510
rect -45 -3540 -40 -3510
rect -80 -3545 -40 -3540
rect -80 -3580 -40 -3575
rect -80 -3610 -75 -3580
rect -75 -3610 -45 -3580
rect -45 -3610 -40 -3580
rect -80 -3615 -40 -3610
rect -80 -3645 -40 -3640
rect -80 -3675 -75 -3645
rect -75 -3675 -45 -3645
rect -45 -3675 -40 -3645
rect -80 -3680 -40 -3675
rect -80 -3705 -40 -3700
rect -80 -3735 -75 -3705
rect -75 -3735 -45 -3705
rect -45 -3735 -40 -3705
rect -80 -3740 -40 -3735
rect -80 -3770 -40 -3765
rect -80 -3800 -75 -3770
rect -75 -3800 -45 -3770
rect -45 -3800 -40 -3770
rect -80 -3805 -40 -3800
rect -80 -3840 -40 -3835
rect -80 -3870 -75 -3840
rect -75 -3870 -45 -3840
rect -45 -3870 -40 -3840
rect -80 -3875 -40 -3870
rect -80 -3910 -40 -3905
rect -80 -3940 -75 -3910
rect -75 -3940 -45 -3910
rect -45 -3940 -40 -3910
rect -80 -3945 -40 -3940
rect -80 -3980 -40 -3975
rect -80 -4010 -75 -3980
rect -75 -4010 -45 -3980
rect -45 -4010 -40 -3980
rect -80 -4015 -40 -4010
rect -80 -4045 -40 -4040
rect -80 -4075 -75 -4045
rect -75 -4075 -45 -4045
rect -45 -4075 -40 -4045
rect -80 -4080 -40 -4075
rect -80 -4105 -40 -4100
rect -80 -4135 -75 -4105
rect -75 -4135 -45 -4105
rect -45 -4135 -40 -4105
rect -80 -4140 -40 -4135
rect -80 -4170 -40 -4165
rect -80 -4200 -75 -4170
rect -75 -4200 -45 -4170
rect -45 -4200 -40 -4170
rect -80 -4205 -40 -4200
rect -80 -4240 -40 -4235
rect -80 -4270 -75 -4240
rect -75 -4270 -45 -4240
rect -45 -4270 -40 -4240
rect -80 -4275 -40 -4270
rect -80 -4310 -40 -4305
rect -80 -4340 -75 -4310
rect -75 -4340 -45 -4310
rect -45 -4340 -40 -4310
rect -80 -4345 -40 -4340
rect -80 -4380 -40 -4375
rect -80 -4410 -75 -4380
rect -75 -4410 -45 -4380
rect -45 -4410 -40 -4380
rect -80 -4415 -40 -4410
rect -80 -4445 -40 -4440
rect -80 -4475 -75 -4445
rect -75 -4475 -45 -4445
rect -45 -4475 -40 -4445
rect -80 -4480 -40 -4475
rect 270 -1305 310 -1300
rect 270 -1335 275 -1305
rect 275 -1335 305 -1305
rect 305 -1335 310 -1305
rect 270 -1340 310 -1335
rect 270 -1370 310 -1365
rect 270 -1400 275 -1370
rect 275 -1400 305 -1370
rect 305 -1400 310 -1370
rect 270 -1405 310 -1400
rect 270 -1440 310 -1435
rect 270 -1470 275 -1440
rect 275 -1470 305 -1440
rect 305 -1470 310 -1440
rect 270 -1475 310 -1470
rect 270 -1510 310 -1505
rect 270 -1540 275 -1510
rect 275 -1540 305 -1510
rect 305 -1540 310 -1510
rect 270 -1545 310 -1540
rect 270 -1580 310 -1575
rect 270 -1610 275 -1580
rect 275 -1610 305 -1580
rect 305 -1610 310 -1580
rect 270 -1615 310 -1610
rect 270 -1645 310 -1640
rect 270 -1675 275 -1645
rect 275 -1675 305 -1645
rect 305 -1675 310 -1645
rect 270 -1680 310 -1675
rect 270 -1705 310 -1700
rect 270 -1735 275 -1705
rect 275 -1735 305 -1705
rect 305 -1735 310 -1705
rect 270 -1740 310 -1735
rect 270 -1770 310 -1765
rect 270 -1800 275 -1770
rect 275 -1800 305 -1770
rect 305 -1800 310 -1770
rect 270 -1805 310 -1800
rect 270 -1840 310 -1835
rect 270 -1870 275 -1840
rect 275 -1870 305 -1840
rect 305 -1870 310 -1840
rect 270 -1875 310 -1870
rect 270 -1910 310 -1905
rect 270 -1940 275 -1910
rect 275 -1940 305 -1910
rect 305 -1940 310 -1910
rect 270 -1945 310 -1940
rect 270 -1980 310 -1975
rect 270 -2010 275 -1980
rect 275 -2010 305 -1980
rect 305 -2010 310 -1980
rect 270 -2015 310 -2010
rect 270 -2045 310 -2040
rect 270 -2075 275 -2045
rect 275 -2075 305 -2045
rect 305 -2075 310 -2045
rect 270 -2080 310 -2075
rect 270 -2105 310 -2100
rect 270 -2135 275 -2105
rect 275 -2135 305 -2105
rect 305 -2135 310 -2105
rect 270 -2140 310 -2135
rect 270 -2170 310 -2165
rect 270 -2200 275 -2170
rect 275 -2200 305 -2170
rect 305 -2200 310 -2170
rect 270 -2205 310 -2200
rect 270 -2240 310 -2235
rect 270 -2270 275 -2240
rect 275 -2270 305 -2240
rect 305 -2270 310 -2240
rect 270 -2275 310 -2270
rect 270 -2310 310 -2305
rect 270 -2340 275 -2310
rect 275 -2340 305 -2310
rect 305 -2340 310 -2310
rect 270 -2345 310 -2340
rect 270 -2380 310 -2375
rect 270 -2410 275 -2380
rect 275 -2410 305 -2380
rect 305 -2410 310 -2380
rect 270 -2415 310 -2410
rect 270 -2445 310 -2440
rect 270 -2475 275 -2445
rect 275 -2475 305 -2445
rect 305 -2475 310 -2445
rect 270 -2480 310 -2475
rect 270 -2505 310 -2500
rect 270 -2535 275 -2505
rect 275 -2535 305 -2505
rect 305 -2535 310 -2505
rect 270 -2540 310 -2535
rect 270 -2570 310 -2565
rect 270 -2600 275 -2570
rect 275 -2600 305 -2570
rect 305 -2600 310 -2570
rect 270 -2605 310 -2600
rect 270 -2640 310 -2635
rect 270 -2670 275 -2640
rect 275 -2670 305 -2640
rect 305 -2670 310 -2640
rect 270 -2675 310 -2670
rect 270 -2710 310 -2705
rect 270 -2740 275 -2710
rect 275 -2740 305 -2710
rect 305 -2740 310 -2710
rect 270 -2745 310 -2740
rect 270 -2780 310 -2775
rect 270 -2810 275 -2780
rect 275 -2810 305 -2780
rect 305 -2810 310 -2780
rect 270 -2815 310 -2810
rect 270 -2845 310 -2840
rect 270 -2875 275 -2845
rect 275 -2875 305 -2845
rect 305 -2875 310 -2845
rect 270 -2880 310 -2875
rect 270 -2905 310 -2900
rect 270 -2935 275 -2905
rect 275 -2935 305 -2905
rect 305 -2935 310 -2905
rect 270 -2940 310 -2935
rect 270 -2970 310 -2965
rect 270 -3000 275 -2970
rect 275 -3000 305 -2970
rect 305 -3000 310 -2970
rect 270 -3005 310 -3000
rect 270 -3040 310 -3035
rect 270 -3070 275 -3040
rect 275 -3070 305 -3040
rect 305 -3070 310 -3040
rect 270 -3075 310 -3070
rect 270 -3110 310 -3105
rect 270 -3140 275 -3110
rect 275 -3140 305 -3110
rect 305 -3140 310 -3110
rect 270 -3145 310 -3140
rect 270 -3180 310 -3175
rect 270 -3210 275 -3180
rect 275 -3210 305 -3180
rect 305 -3210 310 -3180
rect 270 -3215 310 -3210
rect 270 -3245 310 -3240
rect 270 -3275 275 -3245
rect 275 -3275 305 -3245
rect 305 -3275 310 -3245
rect 270 -3280 310 -3275
rect 270 -3305 310 -3300
rect 270 -3335 275 -3305
rect 275 -3335 305 -3305
rect 305 -3335 310 -3305
rect 270 -3340 310 -3335
rect 270 -3370 310 -3365
rect 270 -3400 275 -3370
rect 275 -3400 305 -3370
rect 305 -3400 310 -3370
rect 270 -3405 310 -3400
rect 270 -3440 310 -3435
rect 270 -3470 275 -3440
rect 275 -3470 305 -3440
rect 305 -3470 310 -3440
rect 270 -3475 310 -3470
rect 270 -3510 310 -3505
rect 270 -3540 275 -3510
rect 275 -3540 305 -3510
rect 305 -3540 310 -3510
rect 270 -3545 310 -3540
rect 270 -3580 310 -3575
rect 270 -3610 275 -3580
rect 275 -3610 305 -3580
rect 305 -3610 310 -3580
rect 270 -3615 310 -3610
rect 270 -3645 310 -3640
rect 270 -3675 275 -3645
rect 275 -3675 305 -3645
rect 305 -3675 310 -3645
rect 270 -3680 310 -3675
rect 270 -3705 310 -3700
rect 270 -3735 275 -3705
rect 275 -3735 305 -3705
rect 305 -3735 310 -3705
rect 270 -3740 310 -3735
rect 270 -3770 310 -3765
rect 270 -3800 275 -3770
rect 275 -3800 305 -3770
rect 305 -3800 310 -3770
rect 270 -3805 310 -3800
rect 270 -3840 310 -3835
rect 270 -3870 275 -3840
rect 275 -3870 305 -3840
rect 305 -3870 310 -3840
rect 270 -3875 310 -3870
rect 270 -3910 310 -3905
rect 270 -3940 275 -3910
rect 275 -3940 305 -3910
rect 305 -3940 310 -3910
rect 270 -3945 310 -3940
rect 270 -3980 310 -3975
rect 270 -4010 275 -3980
rect 275 -4010 305 -3980
rect 305 -4010 310 -3980
rect 270 -4015 310 -4010
rect 270 -4045 310 -4040
rect 270 -4075 275 -4045
rect 275 -4075 305 -4045
rect 305 -4075 310 -4045
rect 270 -4080 310 -4075
rect 270 -4105 310 -4100
rect 270 -4135 275 -4105
rect 275 -4135 305 -4105
rect 305 -4135 310 -4105
rect 270 -4140 310 -4135
rect 270 -4170 310 -4165
rect 270 -4200 275 -4170
rect 275 -4200 305 -4170
rect 305 -4200 310 -4170
rect 270 -4205 310 -4200
rect 270 -4240 310 -4235
rect 270 -4270 275 -4240
rect 275 -4270 305 -4240
rect 305 -4270 310 -4240
rect 270 -4275 310 -4270
rect 270 -4310 310 -4305
rect 270 -4340 275 -4310
rect 275 -4340 305 -4310
rect 305 -4340 310 -4310
rect 270 -4345 310 -4340
rect 270 -4380 310 -4375
rect 270 -4410 275 -4380
rect 275 -4410 305 -4380
rect 305 -4410 310 -4380
rect 270 -4415 310 -4410
rect 270 -4445 310 -4440
rect 270 -4475 275 -4445
rect 275 -4475 305 -4445
rect 305 -4475 310 -4445
rect 270 -4480 310 -4475
rect 620 -1305 660 -1300
rect 620 -1335 625 -1305
rect 625 -1335 655 -1305
rect 655 -1335 660 -1305
rect 620 -1340 660 -1335
rect 620 -1370 660 -1365
rect 620 -1400 625 -1370
rect 625 -1400 655 -1370
rect 655 -1400 660 -1370
rect 620 -1405 660 -1400
rect 620 -1440 660 -1435
rect 620 -1470 625 -1440
rect 625 -1470 655 -1440
rect 655 -1470 660 -1440
rect 620 -1475 660 -1470
rect 620 -1510 660 -1505
rect 620 -1540 625 -1510
rect 625 -1540 655 -1510
rect 655 -1540 660 -1510
rect 620 -1545 660 -1540
rect 620 -1580 660 -1575
rect 620 -1610 625 -1580
rect 625 -1610 655 -1580
rect 655 -1610 660 -1580
rect 620 -1615 660 -1610
rect 620 -1645 660 -1640
rect 620 -1675 625 -1645
rect 625 -1675 655 -1645
rect 655 -1675 660 -1645
rect 620 -1680 660 -1675
rect 620 -1705 660 -1700
rect 620 -1735 625 -1705
rect 625 -1735 655 -1705
rect 655 -1735 660 -1705
rect 620 -1740 660 -1735
rect 620 -1770 660 -1765
rect 620 -1800 625 -1770
rect 625 -1800 655 -1770
rect 655 -1800 660 -1770
rect 620 -1805 660 -1800
rect 620 -1840 660 -1835
rect 620 -1870 625 -1840
rect 625 -1870 655 -1840
rect 655 -1870 660 -1840
rect 620 -1875 660 -1870
rect 620 -1910 660 -1905
rect 620 -1940 625 -1910
rect 625 -1940 655 -1910
rect 655 -1940 660 -1910
rect 620 -1945 660 -1940
rect 620 -1980 660 -1975
rect 620 -2010 625 -1980
rect 625 -2010 655 -1980
rect 655 -2010 660 -1980
rect 620 -2015 660 -2010
rect 620 -2045 660 -2040
rect 620 -2075 625 -2045
rect 625 -2075 655 -2045
rect 655 -2075 660 -2045
rect 620 -2080 660 -2075
rect 620 -2105 660 -2100
rect 620 -2135 625 -2105
rect 625 -2135 655 -2105
rect 655 -2135 660 -2105
rect 620 -2140 660 -2135
rect 620 -2170 660 -2165
rect 620 -2200 625 -2170
rect 625 -2200 655 -2170
rect 655 -2200 660 -2170
rect 620 -2205 660 -2200
rect 620 -2240 660 -2235
rect 620 -2270 625 -2240
rect 625 -2270 655 -2240
rect 655 -2270 660 -2240
rect 620 -2275 660 -2270
rect 620 -2310 660 -2305
rect 620 -2340 625 -2310
rect 625 -2340 655 -2310
rect 655 -2340 660 -2310
rect 620 -2345 660 -2340
rect 620 -2380 660 -2375
rect 620 -2410 625 -2380
rect 625 -2410 655 -2380
rect 655 -2410 660 -2380
rect 620 -2415 660 -2410
rect 620 -2445 660 -2440
rect 620 -2475 625 -2445
rect 625 -2475 655 -2445
rect 655 -2475 660 -2445
rect 620 -2480 660 -2475
rect 620 -2505 660 -2500
rect 620 -2535 625 -2505
rect 625 -2535 655 -2505
rect 655 -2535 660 -2505
rect 620 -2540 660 -2535
rect 620 -2570 660 -2565
rect 620 -2600 625 -2570
rect 625 -2600 655 -2570
rect 655 -2600 660 -2570
rect 620 -2605 660 -2600
rect 620 -2640 660 -2635
rect 620 -2670 625 -2640
rect 625 -2670 655 -2640
rect 655 -2670 660 -2640
rect 620 -2675 660 -2670
rect 620 -2710 660 -2705
rect 620 -2740 625 -2710
rect 625 -2740 655 -2710
rect 655 -2740 660 -2710
rect 620 -2745 660 -2740
rect 620 -2780 660 -2775
rect 620 -2810 625 -2780
rect 625 -2810 655 -2780
rect 655 -2810 660 -2780
rect 620 -2815 660 -2810
rect 620 -2845 660 -2840
rect 620 -2875 625 -2845
rect 625 -2875 655 -2845
rect 655 -2875 660 -2845
rect 620 -2880 660 -2875
rect 620 -2905 660 -2900
rect 620 -2935 625 -2905
rect 625 -2935 655 -2905
rect 655 -2935 660 -2905
rect 620 -2940 660 -2935
rect 620 -2970 660 -2965
rect 620 -3000 625 -2970
rect 625 -3000 655 -2970
rect 655 -3000 660 -2970
rect 620 -3005 660 -3000
rect 620 -3040 660 -3035
rect 620 -3070 625 -3040
rect 625 -3070 655 -3040
rect 655 -3070 660 -3040
rect 620 -3075 660 -3070
rect 620 -3110 660 -3105
rect 620 -3140 625 -3110
rect 625 -3140 655 -3110
rect 655 -3140 660 -3110
rect 620 -3145 660 -3140
rect 620 -3180 660 -3175
rect 620 -3210 625 -3180
rect 625 -3210 655 -3180
rect 655 -3210 660 -3180
rect 620 -3215 660 -3210
rect 620 -3245 660 -3240
rect 620 -3275 625 -3245
rect 625 -3275 655 -3245
rect 655 -3275 660 -3245
rect 620 -3280 660 -3275
rect 620 -3305 660 -3300
rect 620 -3335 625 -3305
rect 625 -3335 655 -3305
rect 655 -3335 660 -3305
rect 620 -3340 660 -3335
rect 620 -3370 660 -3365
rect 620 -3400 625 -3370
rect 625 -3400 655 -3370
rect 655 -3400 660 -3370
rect 620 -3405 660 -3400
rect 620 -3440 660 -3435
rect 620 -3470 625 -3440
rect 625 -3470 655 -3440
rect 655 -3470 660 -3440
rect 620 -3475 660 -3470
rect 620 -3510 660 -3505
rect 620 -3540 625 -3510
rect 625 -3540 655 -3510
rect 655 -3540 660 -3510
rect 620 -3545 660 -3540
rect 620 -3580 660 -3575
rect 620 -3610 625 -3580
rect 625 -3610 655 -3580
rect 655 -3610 660 -3580
rect 620 -3615 660 -3610
rect 620 -3645 660 -3640
rect 620 -3675 625 -3645
rect 625 -3675 655 -3645
rect 655 -3675 660 -3645
rect 620 -3680 660 -3675
rect 620 -3705 660 -3700
rect 620 -3735 625 -3705
rect 625 -3735 655 -3705
rect 655 -3735 660 -3705
rect 620 -3740 660 -3735
rect 620 -3770 660 -3765
rect 620 -3800 625 -3770
rect 625 -3800 655 -3770
rect 655 -3800 660 -3770
rect 620 -3805 660 -3800
rect 620 -3840 660 -3835
rect 620 -3870 625 -3840
rect 625 -3870 655 -3840
rect 655 -3870 660 -3840
rect 620 -3875 660 -3870
rect 620 -3910 660 -3905
rect 620 -3940 625 -3910
rect 625 -3940 655 -3910
rect 655 -3940 660 -3910
rect 620 -3945 660 -3940
rect 620 -3980 660 -3975
rect 620 -4010 625 -3980
rect 625 -4010 655 -3980
rect 655 -4010 660 -3980
rect 620 -4015 660 -4010
rect 620 -4045 660 -4040
rect 620 -4075 625 -4045
rect 625 -4075 655 -4045
rect 655 -4075 660 -4045
rect 620 -4080 660 -4075
rect 620 -4105 660 -4100
rect 620 -4135 625 -4105
rect 625 -4135 655 -4105
rect 655 -4135 660 -4105
rect 620 -4140 660 -4135
rect 620 -4170 660 -4165
rect 620 -4200 625 -4170
rect 625 -4200 655 -4170
rect 655 -4200 660 -4170
rect 620 -4205 660 -4200
rect 620 -4240 660 -4235
rect 620 -4270 625 -4240
rect 625 -4270 655 -4240
rect 655 -4270 660 -4240
rect 620 -4275 660 -4270
rect 620 -4310 660 -4305
rect 620 -4340 625 -4310
rect 625 -4340 655 -4310
rect 655 -4340 660 -4310
rect 620 -4345 660 -4340
rect 620 -4380 660 -4375
rect 620 -4410 625 -4380
rect 625 -4410 655 -4380
rect 655 -4410 660 -4380
rect 620 -4415 660 -4410
rect 620 -4445 660 -4440
rect 620 -4475 625 -4445
rect 625 -4475 655 -4445
rect 655 -4475 660 -4445
rect 620 -4480 660 -4475
rect 970 -1305 1010 -1300
rect 970 -1335 975 -1305
rect 975 -1335 1005 -1305
rect 1005 -1335 1010 -1305
rect 970 -1340 1010 -1335
rect 970 -1370 1010 -1365
rect 970 -1400 975 -1370
rect 975 -1400 1005 -1370
rect 1005 -1400 1010 -1370
rect 970 -1405 1010 -1400
rect 970 -1440 1010 -1435
rect 970 -1470 975 -1440
rect 975 -1470 1005 -1440
rect 1005 -1470 1010 -1440
rect 970 -1475 1010 -1470
rect 970 -1510 1010 -1505
rect 970 -1540 975 -1510
rect 975 -1540 1005 -1510
rect 1005 -1540 1010 -1510
rect 970 -1545 1010 -1540
rect 970 -1580 1010 -1575
rect 970 -1610 975 -1580
rect 975 -1610 1005 -1580
rect 1005 -1610 1010 -1580
rect 970 -1615 1010 -1610
rect 970 -1645 1010 -1640
rect 970 -1675 975 -1645
rect 975 -1675 1005 -1645
rect 1005 -1675 1010 -1645
rect 970 -1680 1010 -1675
rect 970 -1705 1010 -1700
rect 970 -1735 975 -1705
rect 975 -1735 1005 -1705
rect 1005 -1735 1010 -1705
rect 970 -1740 1010 -1735
rect 970 -1770 1010 -1765
rect 970 -1800 975 -1770
rect 975 -1800 1005 -1770
rect 1005 -1800 1010 -1770
rect 970 -1805 1010 -1800
rect 970 -1840 1010 -1835
rect 970 -1870 975 -1840
rect 975 -1870 1005 -1840
rect 1005 -1870 1010 -1840
rect 970 -1875 1010 -1870
rect 970 -1910 1010 -1905
rect 970 -1940 975 -1910
rect 975 -1940 1005 -1910
rect 1005 -1940 1010 -1910
rect 970 -1945 1010 -1940
rect 970 -1980 1010 -1975
rect 970 -2010 975 -1980
rect 975 -2010 1005 -1980
rect 1005 -2010 1010 -1980
rect 970 -2015 1010 -2010
rect 970 -2045 1010 -2040
rect 970 -2075 975 -2045
rect 975 -2075 1005 -2045
rect 1005 -2075 1010 -2045
rect 970 -2080 1010 -2075
rect 970 -2105 1010 -2100
rect 970 -2135 975 -2105
rect 975 -2135 1005 -2105
rect 1005 -2135 1010 -2105
rect 970 -2140 1010 -2135
rect 970 -2170 1010 -2165
rect 970 -2200 975 -2170
rect 975 -2200 1005 -2170
rect 1005 -2200 1010 -2170
rect 970 -2205 1010 -2200
rect 970 -2240 1010 -2235
rect 970 -2270 975 -2240
rect 975 -2270 1005 -2240
rect 1005 -2270 1010 -2240
rect 970 -2275 1010 -2270
rect 970 -2310 1010 -2305
rect 970 -2340 975 -2310
rect 975 -2340 1005 -2310
rect 1005 -2340 1010 -2310
rect 970 -2345 1010 -2340
rect 970 -2380 1010 -2375
rect 970 -2410 975 -2380
rect 975 -2410 1005 -2380
rect 1005 -2410 1010 -2380
rect 970 -2415 1010 -2410
rect 970 -2445 1010 -2440
rect 970 -2475 975 -2445
rect 975 -2475 1005 -2445
rect 1005 -2475 1010 -2445
rect 970 -2480 1010 -2475
rect 970 -2505 1010 -2500
rect 970 -2535 975 -2505
rect 975 -2535 1005 -2505
rect 1005 -2535 1010 -2505
rect 970 -2540 1010 -2535
rect 970 -2570 1010 -2565
rect 970 -2600 975 -2570
rect 975 -2600 1005 -2570
rect 1005 -2600 1010 -2570
rect 970 -2605 1010 -2600
rect 970 -2640 1010 -2635
rect 970 -2670 975 -2640
rect 975 -2670 1005 -2640
rect 1005 -2670 1010 -2640
rect 970 -2675 1010 -2670
rect 970 -2710 1010 -2705
rect 970 -2740 975 -2710
rect 975 -2740 1005 -2710
rect 1005 -2740 1010 -2710
rect 970 -2745 1010 -2740
rect 970 -2780 1010 -2775
rect 970 -2810 975 -2780
rect 975 -2810 1005 -2780
rect 1005 -2810 1010 -2780
rect 970 -2815 1010 -2810
rect 970 -2845 1010 -2840
rect 970 -2875 975 -2845
rect 975 -2875 1005 -2845
rect 1005 -2875 1010 -2845
rect 970 -2880 1010 -2875
rect 970 -2905 1010 -2900
rect 970 -2935 975 -2905
rect 975 -2935 1005 -2905
rect 1005 -2935 1010 -2905
rect 970 -2940 1010 -2935
rect 970 -2970 1010 -2965
rect 970 -3000 975 -2970
rect 975 -3000 1005 -2970
rect 1005 -3000 1010 -2970
rect 970 -3005 1010 -3000
rect 970 -3040 1010 -3035
rect 970 -3070 975 -3040
rect 975 -3070 1005 -3040
rect 1005 -3070 1010 -3040
rect 970 -3075 1010 -3070
rect 970 -3110 1010 -3105
rect 970 -3140 975 -3110
rect 975 -3140 1005 -3110
rect 1005 -3140 1010 -3110
rect 970 -3145 1010 -3140
rect 970 -3180 1010 -3175
rect 970 -3210 975 -3180
rect 975 -3210 1005 -3180
rect 1005 -3210 1010 -3180
rect 970 -3215 1010 -3210
rect 970 -3245 1010 -3240
rect 970 -3275 975 -3245
rect 975 -3275 1005 -3245
rect 1005 -3275 1010 -3245
rect 970 -3280 1010 -3275
rect 970 -3305 1010 -3300
rect 970 -3335 975 -3305
rect 975 -3335 1005 -3305
rect 1005 -3335 1010 -3305
rect 970 -3340 1010 -3335
rect 970 -3370 1010 -3365
rect 970 -3400 975 -3370
rect 975 -3400 1005 -3370
rect 1005 -3400 1010 -3370
rect 970 -3405 1010 -3400
rect 970 -3440 1010 -3435
rect 970 -3470 975 -3440
rect 975 -3470 1005 -3440
rect 1005 -3470 1010 -3440
rect 970 -3475 1010 -3470
rect 970 -3510 1010 -3505
rect 970 -3540 975 -3510
rect 975 -3540 1005 -3510
rect 1005 -3540 1010 -3510
rect 970 -3545 1010 -3540
rect 970 -3580 1010 -3575
rect 970 -3610 975 -3580
rect 975 -3610 1005 -3580
rect 1005 -3610 1010 -3580
rect 970 -3615 1010 -3610
rect 970 -3645 1010 -3640
rect 970 -3675 975 -3645
rect 975 -3675 1005 -3645
rect 1005 -3675 1010 -3645
rect 970 -3680 1010 -3675
rect 970 -3705 1010 -3700
rect 970 -3735 975 -3705
rect 975 -3735 1005 -3705
rect 1005 -3735 1010 -3705
rect 970 -3740 1010 -3735
rect 970 -3770 1010 -3765
rect 970 -3800 975 -3770
rect 975 -3800 1005 -3770
rect 1005 -3800 1010 -3770
rect 970 -3805 1010 -3800
rect 970 -3840 1010 -3835
rect 970 -3870 975 -3840
rect 975 -3870 1005 -3840
rect 1005 -3870 1010 -3840
rect 970 -3875 1010 -3870
rect 970 -3910 1010 -3905
rect 970 -3940 975 -3910
rect 975 -3940 1005 -3910
rect 1005 -3940 1010 -3910
rect 970 -3945 1010 -3940
rect 970 -3980 1010 -3975
rect 970 -4010 975 -3980
rect 975 -4010 1005 -3980
rect 1005 -4010 1010 -3980
rect 970 -4015 1010 -4010
rect 970 -4045 1010 -4040
rect 970 -4075 975 -4045
rect 975 -4075 1005 -4045
rect 1005 -4075 1010 -4045
rect 970 -4080 1010 -4075
rect 970 -4105 1010 -4100
rect 970 -4135 975 -4105
rect 975 -4135 1005 -4105
rect 1005 -4135 1010 -4105
rect 970 -4140 1010 -4135
rect 970 -4170 1010 -4165
rect 970 -4200 975 -4170
rect 975 -4200 1005 -4170
rect 1005 -4200 1010 -4170
rect 970 -4205 1010 -4200
rect 970 -4240 1010 -4235
rect 970 -4270 975 -4240
rect 975 -4270 1005 -4240
rect 1005 -4270 1010 -4240
rect 970 -4275 1010 -4270
rect 970 -4310 1010 -4305
rect 970 -4340 975 -4310
rect 975 -4340 1005 -4310
rect 1005 -4340 1010 -4310
rect 970 -4345 1010 -4340
rect 970 -4380 1010 -4375
rect 970 -4410 975 -4380
rect 975 -4410 1005 -4380
rect 1005 -4410 1010 -4380
rect 970 -4415 1010 -4410
rect 970 -4445 1010 -4440
rect 970 -4475 975 -4445
rect 975 -4475 1005 -4445
rect 1005 -4475 1010 -4445
rect 970 -4480 1010 -4475
rect 1320 -1305 1360 -1300
rect 1320 -1335 1325 -1305
rect 1325 -1335 1355 -1305
rect 1355 -1335 1360 -1305
rect 1320 -1340 1360 -1335
rect 1320 -1370 1360 -1365
rect 1320 -1400 1325 -1370
rect 1325 -1400 1355 -1370
rect 1355 -1400 1360 -1370
rect 1320 -1405 1360 -1400
rect 1320 -1440 1360 -1435
rect 1320 -1470 1325 -1440
rect 1325 -1470 1355 -1440
rect 1355 -1470 1360 -1440
rect 1320 -1475 1360 -1470
rect 1320 -1510 1360 -1505
rect 1320 -1540 1325 -1510
rect 1325 -1540 1355 -1510
rect 1355 -1540 1360 -1510
rect 1320 -1545 1360 -1540
rect 1320 -1580 1360 -1575
rect 1320 -1610 1325 -1580
rect 1325 -1610 1355 -1580
rect 1355 -1610 1360 -1580
rect 1320 -1615 1360 -1610
rect 1320 -1645 1360 -1640
rect 1320 -1675 1325 -1645
rect 1325 -1675 1355 -1645
rect 1355 -1675 1360 -1645
rect 1320 -1680 1360 -1675
rect 1320 -1705 1360 -1700
rect 1320 -1735 1325 -1705
rect 1325 -1735 1355 -1705
rect 1355 -1735 1360 -1705
rect 1320 -1740 1360 -1735
rect 1320 -1770 1360 -1765
rect 1320 -1800 1325 -1770
rect 1325 -1800 1355 -1770
rect 1355 -1800 1360 -1770
rect 1320 -1805 1360 -1800
rect 1320 -1840 1360 -1835
rect 1320 -1870 1325 -1840
rect 1325 -1870 1355 -1840
rect 1355 -1870 1360 -1840
rect 1320 -1875 1360 -1870
rect 1320 -1910 1360 -1905
rect 1320 -1940 1325 -1910
rect 1325 -1940 1355 -1910
rect 1355 -1940 1360 -1910
rect 1320 -1945 1360 -1940
rect 1320 -1980 1360 -1975
rect 1320 -2010 1325 -1980
rect 1325 -2010 1355 -1980
rect 1355 -2010 1360 -1980
rect 1320 -2015 1360 -2010
rect 1320 -2045 1360 -2040
rect 1320 -2075 1325 -2045
rect 1325 -2075 1355 -2045
rect 1355 -2075 1360 -2045
rect 1320 -2080 1360 -2075
rect 1320 -2105 1360 -2100
rect 1320 -2135 1325 -2105
rect 1325 -2135 1355 -2105
rect 1355 -2135 1360 -2105
rect 1320 -2140 1360 -2135
rect 1320 -2170 1360 -2165
rect 1320 -2200 1325 -2170
rect 1325 -2200 1355 -2170
rect 1355 -2200 1360 -2170
rect 1320 -2205 1360 -2200
rect 1320 -2240 1360 -2235
rect 1320 -2270 1325 -2240
rect 1325 -2270 1355 -2240
rect 1355 -2270 1360 -2240
rect 1320 -2275 1360 -2270
rect 1320 -2310 1360 -2305
rect 1320 -2340 1325 -2310
rect 1325 -2340 1355 -2310
rect 1355 -2340 1360 -2310
rect 1320 -2345 1360 -2340
rect 1320 -2380 1360 -2375
rect 1320 -2410 1325 -2380
rect 1325 -2410 1355 -2380
rect 1355 -2410 1360 -2380
rect 1320 -2415 1360 -2410
rect 1320 -2445 1360 -2440
rect 1320 -2475 1325 -2445
rect 1325 -2475 1355 -2445
rect 1355 -2475 1360 -2445
rect 1320 -2480 1360 -2475
rect 1320 -2505 1360 -2500
rect 1320 -2535 1325 -2505
rect 1325 -2535 1355 -2505
rect 1355 -2535 1360 -2505
rect 1320 -2540 1360 -2535
rect 1320 -2570 1360 -2565
rect 1320 -2600 1325 -2570
rect 1325 -2600 1355 -2570
rect 1355 -2600 1360 -2570
rect 1320 -2605 1360 -2600
rect 1320 -2640 1360 -2635
rect 1320 -2670 1325 -2640
rect 1325 -2670 1355 -2640
rect 1355 -2670 1360 -2640
rect 1320 -2675 1360 -2670
rect 1320 -2710 1360 -2705
rect 1320 -2740 1325 -2710
rect 1325 -2740 1355 -2710
rect 1355 -2740 1360 -2710
rect 1320 -2745 1360 -2740
rect 1320 -2780 1360 -2775
rect 1320 -2810 1325 -2780
rect 1325 -2810 1355 -2780
rect 1355 -2810 1360 -2780
rect 1320 -2815 1360 -2810
rect 1320 -2845 1360 -2840
rect 1320 -2875 1325 -2845
rect 1325 -2875 1355 -2845
rect 1355 -2875 1360 -2845
rect 1320 -2880 1360 -2875
rect 1320 -2905 1360 -2900
rect 1320 -2935 1325 -2905
rect 1325 -2935 1355 -2905
rect 1355 -2935 1360 -2905
rect 1320 -2940 1360 -2935
rect 1320 -2970 1360 -2965
rect 1320 -3000 1325 -2970
rect 1325 -3000 1355 -2970
rect 1355 -3000 1360 -2970
rect 1320 -3005 1360 -3000
rect 1320 -3040 1360 -3035
rect 1320 -3070 1325 -3040
rect 1325 -3070 1355 -3040
rect 1355 -3070 1360 -3040
rect 1320 -3075 1360 -3070
rect 1320 -3110 1360 -3105
rect 1320 -3140 1325 -3110
rect 1325 -3140 1355 -3110
rect 1355 -3140 1360 -3110
rect 1320 -3145 1360 -3140
rect 1320 -3180 1360 -3175
rect 1320 -3210 1325 -3180
rect 1325 -3210 1355 -3180
rect 1355 -3210 1360 -3180
rect 1320 -3215 1360 -3210
rect 1320 -3245 1360 -3240
rect 1320 -3275 1325 -3245
rect 1325 -3275 1355 -3245
rect 1355 -3275 1360 -3245
rect 1320 -3280 1360 -3275
rect 1320 -3305 1360 -3300
rect 1320 -3335 1325 -3305
rect 1325 -3335 1355 -3305
rect 1355 -3335 1360 -3305
rect 1320 -3340 1360 -3335
rect 1320 -3370 1360 -3365
rect 1320 -3400 1325 -3370
rect 1325 -3400 1355 -3370
rect 1355 -3400 1360 -3370
rect 1320 -3405 1360 -3400
rect 1320 -3440 1360 -3435
rect 1320 -3470 1325 -3440
rect 1325 -3470 1355 -3440
rect 1355 -3470 1360 -3440
rect 1320 -3475 1360 -3470
rect 1320 -3510 1360 -3505
rect 1320 -3540 1325 -3510
rect 1325 -3540 1355 -3510
rect 1355 -3540 1360 -3510
rect 1320 -3545 1360 -3540
rect 1320 -3580 1360 -3575
rect 1320 -3610 1325 -3580
rect 1325 -3610 1355 -3580
rect 1355 -3610 1360 -3580
rect 1320 -3615 1360 -3610
rect 1320 -3645 1360 -3640
rect 1320 -3675 1325 -3645
rect 1325 -3675 1355 -3645
rect 1355 -3675 1360 -3645
rect 1320 -3680 1360 -3675
rect 1320 -3705 1360 -3700
rect 1320 -3735 1325 -3705
rect 1325 -3735 1355 -3705
rect 1355 -3735 1360 -3705
rect 1320 -3740 1360 -3735
rect 1320 -3770 1360 -3765
rect 1320 -3800 1325 -3770
rect 1325 -3800 1355 -3770
rect 1355 -3800 1360 -3770
rect 1320 -3805 1360 -3800
rect 1320 -3840 1360 -3835
rect 1320 -3870 1325 -3840
rect 1325 -3870 1355 -3840
rect 1355 -3870 1360 -3840
rect 1320 -3875 1360 -3870
rect 1320 -3910 1360 -3905
rect 1320 -3940 1325 -3910
rect 1325 -3940 1355 -3910
rect 1355 -3940 1360 -3910
rect 1320 -3945 1360 -3940
rect 1320 -3980 1360 -3975
rect 1320 -4010 1325 -3980
rect 1325 -4010 1355 -3980
rect 1355 -4010 1360 -3980
rect 1320 -4015 1360 -4010
rect 1320 -4045 1360 -4040
rect 1320 -4075 1325 -4045
rect 1325 -4075 1355 -4045
rect 1355 -4075 1360 -4045
rect 1320 -4080 1360 -4075
rect 1320 -4105 1360 -4100
rect 1320 -4135 1325 -4105
rect 1325 -4135 1355 -4105
rect 1355 -4135 1360 -4105
rect 1320 -4140 1360 -4135
rect 1320 -4170 1360 -4165
rect 1320 -4200 1325 -4170
rect 1325 -4200 1355 -4170
rect 1355 -4200 1360 -4170
rect 1320 -4205 1360 -4200
rect 1320 -4240 1360 -4235
rect 1320 -4270 1325 -4240
rect 1325 -4270 1355 -4240
rect 1355 -4270 1360 -4240
rect 1320 -4275 1360 -4270
rect 1320 -4310 1360 -4305
rect 1320 -4340 1325 -4310
rect 1325 -4340 1355 -4310
rect 1355 -4340 1360 -4310
rect 1320 -4345 1360 -4340
rect 1320 -4380 1360 -4375
rect 1320 -4410 1325 -4380
rect 1325 -4410 1355 -4380
rect 1355 -4410 1360 -4380
rect 1320 -4415 1360 -4410
rect 1320 -4445 1360 -4440
rect 1320 -4475 1325 -4445
rect 1325 -4475 1355 -4445
rect 1355 -4475 1360 -4445
rect 1320 -4480 1360 -4475
rect 1670 -1305 1710 -1300
rect 1670 -1335 1675 -1305
rect 1675 -1335 1705 -1305
rect 1705 -1335 1710 -1305
rect 1670 -1340 1710 -1335
rect 1670 -1370 1710 -1365
rect 1670 -1400 1675 -1370
rect 1675 -1400 1705 -1370
rect 1705 -1400 1710 -1370
rect 1670 -1405 1710 -1400
rect 1670 -1440 1710 -1435
rect 1670 -1470 1675 -1440
rect 1675 -1470 1705 -1440
rect 1705 -1470 1710 -1440
rect 1670 -1475 1710 -1470
rect 1670 -1510 1710 -1505
rect 1670 -1540 1675 -1510
rect 1675 -1540 1705 -1510
rect 1705 -1540 1710 -1510
rect 1670 -1545 1710 -1540
rect 1670 -1580 1710 -1575
rect 1670 -1610 1675 -1580
rect 1675 -1610 1705 -1580
rect 1705 -1610 1710 -1580
rect 1670 -1615 1710 -1610
rect 1670 -1645 1710 -1640
rect 1670 -1675 1675 -1645
rect 1675 -1675 1705 -1645
rect 1705 -1675 1710 -1645
rect 1670 -1680 1710 -1675
rect 1670 -1705 1710 -1700
rect 1670 -1735 1675 -1705
rect 1675 -1735 1705 -1705
rect 1705 -1735 1710 -1705
rect 1670 -1740 1710 -1735
rect 1670 -1770 1710 -1765
rect 1670 -1800 1675 -1770
rect 1675 -1800 1705 -1770
rect 1705 -1800 1710 -1770
rect 1670 -1805 1710 -1800
rect 1670 -1840 1710 -1835
rect 1670 -1870 1675 -1840
rect 1675 -1870 1705 -1840
rect 1705 -1870 1710 -1840
rect 1670 -1875 1710 -1870
rect 1670 -1910 1710 -1905
rect 1670 -1940 1675 -1910
rect 1675 -1940 1705 -1910
rect 1705 -1940 1710 -1910
rect 1670 -1945 1710 -1940
rect 1670 -1980 1710 -1975
rect 1670 -2010 1675 -1980
rect 1675 -2010 1705 -1980
rect 1705 -2010 1710 -1980
rect 1670 -2015 1710 -2010
rect 1670 -2045 1710 -2040
rect 1670 -2075 1675 -2045
rect 1675 -2075 1705 -2045
rect 1705 -2075 1710 -2045
rect 1670 -2080 1710 -2075
rect 1670 -2105 1710 -2100
rect 1670 -2135 1675 -2105
rect 1675 -2135 1705 -2105
rect 1705 -2135 1710 -2105
rect 1670 -2140 1710 -2135
rect 1670 -2170 1710 -2165
rect 1670 -2200 1675 -2170
rect 1675 -2200 1705 -2170
rect 1705 -2200 1710 -2170
rect 1670 -2205 1710 -2200
rect 1670 -2240 1710 -2235
rect 1670 -2270 1675 -2240
rect 1675 -2270 1705 -2240
rect 1705 -2270 1710 -2240
rect 1670 -2275 1710 -2270
rect 1670 -2310 1710 -2305
rect 1670 -2340 1675 -2310
rect 1675 -2340 1705 -2310
rect 1705 -2340 1710 -2310
rect 1670 -2345 1710 -2340
rect 1670 -2380 1710 -2375
rect 1670 -2410 1675 -2380
rect 1675 -2410 1705 -2380
rect 1705 -2410 1710 -2380
rect 1670 -2415 1710 -2410
rect 1670 -2445 1710 -2440
rect 1670 -2475 1675 -2445
rect 1675 -2475 1705 -2445
rect 1705 -2475 1710 -2445
rect 1670 -2480 1710 -2475
rect 1670 -2505 1710 -2500
rect 1670 -2535 1675 -2505
rect 1675 -2535 1705 -2505
rect 1705 -2535 1710 -2505
rect 1670 -2540 1710 -2535
rect 1670 -2570 1710 -2565
rect 1670 -2600 1675 -2570
rect 1675 -2600 1705 -2570
rect 1705 -2600 1710 -2570
rect 1670 -2605 1710 -2600
rect 1670 -2640 1710 -2635
rect 1670 -2670 1675 -2640
rect 1675 -2670 1705 -2640
rect 1705 -2670 1710 -2640
rect 1670 -2675 1710 -2670
rect 1670 -2710 1710 -2705
rect 1670 -2740 1675 -2710
rect 1675 -2740 1705 -2710
rect 1705 -2740 1710 -2710
rect 1670 -2745 1710 -2740
rect 1670 -2780 1710 -2775
rect 1670 -2810 1675 -2780
rect 1675 -2810 1705 -2780
rect 1705 -2810 1710 -2780
rect 1670 -2815 1710 -2810
rect 1670 -2845 1710 -2840
rect 1670 -2875 1675 -2845
rect 1675 -2875 1705 -2845
rect 1705 -2875 1710 -2845
rect 1670 -2880 1710 -2875
rect 1670 -2905 1710 -2900
rect 1670 -2935 1675 -2905
rect 1675 -2935 1705 -2905
rect 1705 -2935 1710 -2905
rect 1670 -2940 1710 -2935
rect 1670 -2970 1710 -2965
rect 1670 -3000 1675 -2970
rect 1675 -3000 1705 -2970
rect 1705 -3000 1710 -2970
rect 1670 -3005 1710 -3000
rect 1670 -3040 1710 -3035
rect 1670 -3070 1675 -3040
rect 1675 -3070 1705 -3040
rect 1705 -3070 1710 -3040
rect 1670 -3075 1710 -3070
rect 1670 -3110 1710 -3105
rect 1670 -3140 1675 -3110
rect 1675 -3140 1705 -3110
rect 1705 -3140 1710 -3110
rect 1670 -3145 1710 -3140
rect 1670 -3180 1710 -3175
rect 1670 -3210 1675 -3180
rect 1675 -3210 1705 -3180
rect 1705 -3210 1710 -3180
rect 1670 -3215 1710 -3210
rect 1670 -3245 1710 -3240
rect 1670 -3275 1675 -3245
rect 1675 -3275 1705 -3245
rect 1705 -3275 1710 -3245
rect 1670 -3280 1710 -3275
rect 1670 -3305 1710 -3300
rect 1670 -3335 1675 -3305
rect 1675 -3335 1705 -3305
rect 1705 -3335 1710 -3305
rect 1670 -3340 1710 -3335
rect 1670 -3370 1710 -3365
rect 1670 -3400 1675 -3370
rect 1675 -3400 1705 -3370
rect 1705 -3400 1710 -3370
rect 1670 -3405 1710 -3400
rect 1670 -3440 1710 -3435
rect 1670 -3470 1675 -3440
rect 1675 -3470 1705 -3440
rect 1705 -3470 1710 -3440
rect 1670 -3475 1710 -3470
rect 1670 -3510 1710 -3505
rect 1670 -3540 1675 -3510
rect 1675 -3540 1705 -3510
rect 1705 -3540 1710 -3510
rect 1670 -3545 1710 -3540
rect 1670 -3580 1710 -3575
rect 1670 -3610 1675 -3580
rect 1675 -3610 1705 -3580
rect 1705 -3610 1710 -3580
rect 1670 -3615 1710 -3610
rect 1670 -3645 1710 -3640
rect 1670 -3675 1675 -3645
rect 1675 -3675 1705 -3645
rect 1705 -3675 1710 -3645
rect 1670 -3680 1710 -3675
rect 1670 -3705 1710 -3700
rect 1670 -3735 1675 -3705
rect 1675 -3735 1705 -3705
rect 1705 -3735 1710 -3705
rect 1670 -3740 1710 -3735
rect 1670 -3770 1710 -3765
rect 1670 -3800 1675 -3770
rect 1675 -3800 1705 -3770
rect 1705 -3800 1710 -3770
rect 1670 -3805 1710 -3800
rect 1670 -3840 1710 -3835
rect 1670 -3870 1675 -3840
rect 1675 -3870 1705 -3840
rect 1705 -3870 1710 -3840
rect 1670 -3875 1710 -3870
rect 1670 -3910 1710 -3905
rect 1670 -3940 1675 -3910
rect 1675 -3940 1705 -3910
rect 1705 -3940 1710 -3910
rect 1670 -3945 1710 -3940
rect 1670 -3980 1710 -3975
rect 1670 -4010 1675 -3980
rect 1675 -4010 1705 -3980
rect 1705 -4010 1710 -3980
rect 1670 -4015 1710 -4010
rect 1670 -4045 1710 -4040
rect 1670 -4075 1675 -4045
rect 1675 -4075 1705 -4045
rect 1705 -4075 1710 -4045
rect 1670 -4080 1710 -4075
rect 1670 -4105 1710 -4100
rect 1670 -4135 1675 -4105
rect 1675 -4135 1705 -4105
rect 1705 -4135 1710 -4105
rect 1670 -4140 1710 -4135
rect 1670 -4170 1710 -4165
rect 1670 -4200 1675 -4170
rect 1675 -4200 1705 -4170
rect 1705 -4200 1710 -4170
rect 1670 -4205 1710 -4200
rect 1670 -4240 1710 -4235
rect 1670 -4270 1675 -4240
rect 1675 -4270 1705 -4240
rect 1705 -4270 1710 -4240
rect 1670 -4275 1710 -4270
rect 1670 -4310 1710 -4305
rect 1670 -4340 1675 -4310
rect 1675 -4340 1705 -4310
rect 1705 -4340 1710 -4310
rect 1670 -4345 1710 -4340
rect 1670 -4380 1710 -4375
rect 1670 -4410 1675 -4380
rect 1675 -4410 1705 -4380
rect 1705 -4410 1710 -4380
rect 1670 -4415 1710 -4410
rect 1670 -4445 1710 -4440
rect 1670 -4475 1675 -4445
rect 1675 -4475 1705 -4445
rect 1705 -4475 1710 -4445
rect 1670 -4480 1710 -4475
rect 2020 -1305 2060 -1300
rect 2020 -1335 2025 -1305
rect 2025 -1335 2055 -1305
rect 2055 -1335 2060 -1305
rect 2020 -1340 2060 -1335
rect 2020 -1370 2060 -1365
rect 2020 -1400 2025 -1370
rect 2025 -1400 2055 -1370
rect 2055 -1400 2060 -1370
rect 2020 -1405 2060 -1400
rect 2020 -1440 2060 -1435
rect 2020 -1470 2025 -1440
rect 2025 -1470 2055 -1440
rect 2055 -1470 2060 -1440
rect 2020 -1475 2060 -1470
rect 2020 -1510 2060 -1505
rect 2020 -1540 2025 -1510
rect 2025 -1540 2055 -1510
rect 2055 -1540 2060 -1510
rect 2020 -1545 2060 -1540
rect 2020 -1580 2060 -1575
rect 2020 -1610 2025 -1580
rect 2025 -1610 2055 -1580
rect 2055 -1610 2060 -1580
rect 2020 -1615 2060 -1610
rect 2020 -1645 2060 -1640
rect 2020 -1675 2025 -1645
rect 2025 -1675 2055 -1645
rect 2055 -1675 2060 -1645
rect 2020 -1680 2060 -1675
rect 2020 -1705 2060 -1700
rect 2020 -1735 2025 -1705
rect 2025 -1735 2055 -1705
rect 2055 -1735 2060 -1705
rect 2020 -1740 2060 -1735
rect 2020 -1770 2060 -1765
rect 2020 -1800 2025 -1770
rect 2025 -1800 2055 -1770
rect 2055 -1800 2060 -1770
rect 2020 -1805 2060 -1800
rect 2020 -1840 2060 -1835
rect 2020 -1870 2025 -1840
rect 2025 -1870 2055 -1840
rect 2055 -1870 2060 -1840
rect 2020 -1875 2060 -1870
rect 2020 -1910 2060 -1905
rect 2020 -1940 2025 -1910
rect 2025 -1940 2055 -1910
rect 2055 -1940 2060 -1910
rect 2020 -1945 2060 -1940
rect 2020 -1980 2060 -1975
rect 2020 -2010 2025 -1980
rect 2025 -2010 2055 -1980
rect 2055 -2010 2060 -1980
rect 2020 -2015 2060 -2010
rect 2020 -2045 2060 -2040
rect 2020 -2075 2025 -2045
rect 2025 -2075 2055 -2045
rect 2055 -2075 2060 -2045
rect 2020 -2080 2060 -2075
rect 2020 -2105 2060 -2100
rect 2020 -2135 2025 -2105
rect 2025 -2135 2055 -2105
rect 2055 -2135 2060 -2105
rect 2020 -2140 2060 -2135
rect 2020 -2170 2060 -2165
rect 2020 -2200 2025 -2170
rect 2025 -2200 2055 -2170
rect 2055 -2200 2060 -2170
rect 2020 -2205 2060 -2200
rect 2020 -2240 2060 -2235
rect 2020 -2270 2025 -2240
rect 2025 -2270 2055 -2240
rect 2055 -2270 2060 -2240
rect 2020 -2275 2060 -2270
rect 2020 -2310 2060 -2305
rect 2020 -2340 2025 -2310
rect 2025 -2340 2055 -2310
rect 2055 -2340 2060 -2310
rect 2020 -2345 2060 -2340
rect 2020 -2380 2060 -2375
rect 2020 -2410 2025 -2380
rect 2025 -2410 2055 -2380
rect 2055 -2410 2060 -2380
rect 2020 -2415 2060 -2410
rect 2020 -2445 2060 -2440
rect 2020 -2475 2025 -2445
rect 2025 -2475 2055 -2445
rect 2055 -2475 2060 -2445
rect 2020 -2480 2060 -2475
rect 2020 -2505 2060 -2500
rect 2020 -2535 2025 -2505
rect 2025 -2535 2055 -2505
rect 2055 -2535 2060 -2505
rect 2020 -2540 2060 -2535
rect 2020 -2570 2060 -2565
rect 2020 -2600 2025 -2570
rect 2025 -2600 2055 -2570
rect 2055 -2600 2060 -2570
rect 2020 -2605 2060 -2600
rect 2020 -2640 2060 -2635
rect 2020 -2670 2025 -2640
rect 2025 -2670 2055 -2640
rect 2055 -2670 2060 -2640
rect 2020 -2675 2060 -2670
rect 2020 -2710 2060 -2705
rect 2020 -2740 2025 -2710
rect 2025 -2740 2055 -2710
rect 2055 -2740 2060 -2710
rect 2020 -2745 2060 -2740
rect 2020 -2780 2060 -2775
rect 2020 -2810 2025 -2780
rect 2025 -2810 2055 -2780
rect 2055 -2810 2060 -2780
rect 2020 -2815 2060 -2810
rect 2020 -2845 2060 -2840
rect 2020 -2875 2025 -2845
rect 2025 -2875 2055 -2845
rect 2055 -2875 2060 -2845
rect 2020 -2880 2060 -2875
rect 2020 -2905 2060 -2900
rect 2020 -2935 2025 -2905
rect 2025 -2935 2055 -2905
rect 2055 -2935 2060 -2905
rect 2020 -2940 2060 -2935
rect 2020 -2970 2060 -2965
rect 2020 -3000 2025 -2970
rect 2025 -3000 2055 -2970
rect 2055 -3000 2060 -2970
rect 2020 -3005 2060 -3000
rect 2020 -3040 2060 -3035
rect 2020 -3070 2025 -3040
rect 2025 -3070 2055 -3040
rect 2055 -3070 2060 -3040
rect 2020 -3075 2060 -3070
rect 2020 -3110 2060 -3105
rect 2020 -3140 2025 -3110
rect 2025 -3140 2055 -3110
rect 2055 -3140 2060 -3110
rect 2020 -3145 2060 -3140
rect 2020 -3180 2060 -3175
rect 2020 -3210 2025 -3180
rect 2025 -3210 2055 -3180
rect 2055 -3210 2060 -3180
rect 2020 -3215 2060 -3210
rect 2020 -3245 2060 -3240
rect 2020 -3275 2025 -3245
rect 2025 -3275 2055 -3245
rect 2055 -3275 2060 -3245
rect 2020 -3280 2060 -3275
rect 2020 -3305 2060 -3300
rect 2020 -3335 2025 -3305
rect 2025 -3335 2055 -3305
rect 2055 -3335 2060 -3305
rect 2020 -3340 2060 -3335
rect 2020 -3370 2060 -3365
rect 2020 -3400 2025 -3370
rect 2025 -3400 2055 -3370
rect 2055 -3400 2060 -3370
rect 2020 -3405 2060 -3400
rect 2020 -3440 2060 -3435
rect 2020 -3470 2025 -3440
rect 2025 -3470 2055 -3440
rect 2055 -3470 2060 -3440
rect 2020 -3475 2060 -3470
rect 2020 -3510 2060 -3505
rect 2020 -3540 2025 -3510
rect 2025 -3540 2055 -3510
rect 2055 -3540 2060 -3510
rect 2020 -3545 2060 -3540
rect 2020 -3580 2060 -3575
rect 2020 -3610 2025 -3580
rect 2025 -3610 2055 -3580
rect 2055 -3610 2060 -3580
rect 2020 -3615 2060 -3610
rect 2020 -3645 2060 -3640
rect 2020 -3675 2025 -3645
rect 2025 -3675 2055 -3645
rect 2055 -3675 2060 -3645
rect 2020 -3680 2060 -3675
rect 2020 -3705 2060 -3700
rect 2020 -3735 2025 -3705
rect 2025 -3735 2055 -3705
rect 2055 -3735 2060 -3705
rect 2020 -3740 2060 -3735
rect 2020 -3770 2060 -3765
rect 2020 -3800 2025 -3770
rect 2025 -3800 2055 -3770
rect 2055 -3800 2060 -3770
rect 2020 -3805 2060 -3800
rect 2020 -3840 2060 -3835
rect 2020 -3870 2025 -3840
rect 2025 -3870 2055 -3840
rect 2055 -3870 2060 -3840
rect 2020 -3875 2060 -3870
rect 2020 -3910 2060 -3905
rect 2020 -3940 2025 -3910
rect 2025 -3940 2055 -3910
rect 2055 -3940 2060 -3910
rect 2020 -3945 2060 -3940
rect 2020 -3980 2060 -3975
rect 2020 -4010 2025 -3980
rect 2025 -4010 2055 -3980
rect 2055 -4010 2060 -3980
rect 2020 -4015 2060 -4010
rect 2020 -4045 2060 -4040
rect 2020 -4075 2025 -4045
rect 2025 -4075 2055 -4045
rect 2055 -4075 2060 -4045
rect 2020 -4080 2060 -4075
rect 2020 -4105 2060 -4100
rect 2020 -4135 2025 -4105
rect 2025 -4135 2055 -4105
rect 2055 -4135 2060 -4105
rect 2020 -4140 2060 -4135
rect 2020 -4170 2060 -4165
rect 2020 -4200 2025 -4170
rect 2025 -4200 2055 -4170
rect 2055 -4200 2060 -4170
rect 2020 -4205 2060 -4200
rect 2020 -4240 2060 -4235
rect 2020 -4270 2025 -4240
rect 2025 -4270 2055 -4240
rect 2055 -4270 2060 -4240
rect 2020 -4275 2060 -4270
rect 2020 -4310 2060 -4305
rect 2020 -4340 2025 -4310
rect 2025 -4340 2055 -4310
rect 2055 -4340 2060 -4310
rect 2020 -4345 2060 -4340
rect 2020 -4380 2060 -4375
rect 2020 -4410 2025 -4380
rect 2025 -4410 2055 -4380
rect 2055 -4410 2060 -4380
rect 2020 -4415 2060 -4410
rect 2020 -4445 2060 -4440
rect 2020 -4475 2025 -4445
rect 2025 -4475 2055 -4445
rect 2055 -4475 2060 -4445
rect 2020 -4480 2060 -4475
rect 2370 -1305 2410 -1300
rect 2370 -1335 2375 -1305
rect 2375 -1335 2405 -1305
rect 2405 -1335 2410 -1305
rect 2370 -1340 2410 -1335
rect 2370 -1370 2410 -1365
rect 2370 -1400 2375 -1370
rect 2375 -1400 2405 -1370
rect 2405 -1400 2410 -1370
rect 2370 -1405 2410 -1400
rect 2370 -1440 2410 -1435
rect 2370 -1470 2375 -1440
rect 2375 -1470 2405 -1440
rect 2405 -1470 2410 -1440
rect 2370 -1475 2410 -1470
rect 2370 -1510 2410 -1505
rect 2370 -1540 2375 -1510
rect 2375 -1540 2405 -1510
rect 2405 -1540 2410 -1510
rect 2370 -1545 2410 -1540
rect 2370 -1580 2410 -1575
rect 2370 -1610 2375 -1580
rect 2375 -1610 2405 -1580
rect 2405 -1610 2410 -1580
rect 2370 -1615 2410 -1610
rect 2370 -1645 2410 -1640
rect 2370 -1675 2375 -1645
rect 2375 -1675 2405 -1645
rect 2405 -1675 2410 -1645
rect 2370 -1680 2410 -1675
rect 2370 -1705 2410 -1700
rect 2370 -1735 2375 -1705
rect 2375 -1735 2405 -1705
rect 2405 -1735 2410 -1705
rect 2370 -1740 2410 -1735
rect 2370 -1770 2410 -1765
rect 2370 -1800 2375 -1770
rect 2375 -1800 2405 -1770
rect 2405 -1800 2410 -1770
rect 2370 -1805 2410 -1800
rect 2370 -1840 2410 -1835
rect 2370 -1870 2375 -1840
rect 2375 -1870 2405 -1840
rect 2405 -1870 2410 -1840
rect 2370 -1875 2410 -1870
rect 2370 -1910 2410 -1905
rect 2370 -1940 2375 -1910
rect 2375 -1940 2405 -1910
rect 2405 -1940 2410 -1910
rect 2370 -1945 2410 -1940
rect 2370 -1980 2410 -1975
rect 2370 -2010 2375 -1980
rect 2375 -2010 2405 -1980
rect 2405 -2010 2410 -1980
rect 2370 -2015 2410 -2010
rect 2370 -2045 2410 -2040
rect 2370 -2075 2375 -2045
rect 2375 -2075 2405 -2045
rect 2405 -2075 2410 -2045
rect 2370 -2080 2410 -2075
rect 2370 -2105 2410 -2100
rect 2370 -2135 2375 -2105
rect 2375 -2135 2405 -2105
rect 2405 -2135 2410 -2105
rect 2370 -2140 2410 -2135
rect 2370 -2170 2410 -2165
rect 2370 -2200 2375 -2170
rect 2375 -2200 2405 -2170
rect 2405 -2200 2410 -2170
rect 2370 -2205 2410 -2200
rect 2370 -2240 2410 -2235
rect 2370 -2270 2375 -2240
rect 2375 -2270 2405 -2240
rect 2405 -2270 2410 -2240
rect 2370 -2275 2410 -2270
rect 2370 -2310 2410 -2305
rect 2370 -2340 2375 -2310
rect 2375 -2340 2405 -2310
rect 2405 -2340 2410 -2310
rect 2370 -2345 2410 -2340
rect 2370 -2380 2410 -2375
rect 2370 -2410 2375 -2380
rect 2375 -2410 2405 -2380
rect 2405 -2410 2410 -2380
rect 2370 -2415 2410 -2410
rect 2370 -2445 2410 -2440
rect 2370 -2475 2375 -2445
rect 2375 -2475 2405 -2445
rect 2405 -2475 2410 -2445
rect 2370 -2480 2410 -2475
rect 2370 -2505 2410 -2500
rect 2370 -2535 2375 -2505
rect 2375 -2535 2405 -2505
rect 2405 -2535 2410 -2505
rect 2370 -2540 2410 -2535
rect 2370 -2570 2410 -2565
rect 2370 -2600 2375 -2570
rect 2375 -2600 2405 -2570
rect 2405 -2600 2410 -2570
rect 2370 -2605 2410 -2600
rect 2370 -2640 2410 -2635
rect 2370 -2670 2375 -2640
rect 2375 -2670 2405 -2640
rect 2405 -2670 2410 -2640
rect 2370 -2675 2410 -2670
rect 2370 -2710 2410 -2705
rect 2370 -2740 2375 -2710
rect 2375 -2740 2405 -2710
rect 2405 -2740 2410 -2710
rect 2370 -2745 2410 -2740
rect 2370 -2780 2410 -2775
rect 2370 -2810 2375 -2780
rect 2375 -2810 2405 -2780
rect 2405 -2810 2410 -2780
rect 2370 -2815 2410 -2810
rect 2370 -2845 2410 -2840
rect 2370 -2875 2375 -2845
rect 2375 -2875 2405 -2845
rect 2405 -2875 2410 -2845
rect 2370 -2880 2410 -2875
rect 2370 -2905 2410 -2900
rect 2370 -2935 2375 -2905
rect 2375 -2935 2405 -2905
rect 2405 -2935 2410 -2905
rect 2370 -2940 2410 -2935
rect 2370 -2970 2410 -2965
rect 2370 -3000 2375 -2970
rect 2375 -3000 2405 -2970
rect 2405 -3000 2410 -2970
rect 2370 -3005 2410 -3000
rect 2370 -3040 2410 -3035
rect 2370 -3070 2375 -3040
rect 2375 -3070 2405 -3040
rect 2405 -3070 2410 -3040
rect 2370 -3075 2410 -3070
rect 2370 -3110 2410 -3105
rect 2370 -3140 2375 -3110
rect 2375 -3140 2405 -3110
rect 2405 -3140 2410 -3110
rect 2370 -3145 2410 -3140
rect 2370 -3180 2410 -3175
rect 2370 -3210 2375 -3180
rect 2375 -3210 2405 -3180
rect 2405 -3210 2410 -3180
rect 2370 -3215 2410 -3210
rect 2370 -3245 2410 -3240
rect 2370 -3275 2375 -3245
rect 2375 -3275 2405 -3245
rect 2405 -3275 2410 -3245
rect 2370 -3280 2410 -3275
rect 2370 -3305 2410 -3300
rect 2370 -3335 2375 -3305
rect 2375 -3335 2405 -3305
rect 2405 -3335 2410 -3305
rect 2370 -3340 2410 -3335
rect 2370 -3370 2410 -3365
rect 2370 -3400 2375 -3370
rect 2375 -3400 2405 -3370
rect 2405 -3400 2410 -3370
rect 2370 -3405 2410 -3400
rect 2370 -3440 2410 -3435
rect 2370 -3470 2375 -3440
rect 2375 -3470 2405 -3440
rect 2405 -3470 2410 -3440
rect 2370 -3475 2410 -3470
rect 2370 -3510 2410 -3505
rect 2370 -3540 2375 -3510
rect 2375 -3540 2405 -3510
rect 2405 -3540 2410 -3510
rect 2370 -3545 2410 -3540
rect 2370 -3580 2410 -3575
rect 2370 -3610 2375 -3580
rect 2375 -3610 2405 -3580
rect 2405 -3610 2410 -3580
rect 2370 -3615 2410 -3610
rect 2370 -3645 2410 -3640
rect 2370 -3675 2375 -3645
rect 2375 -3675 2405 -3645
rect 2405 -3675 2410 -3645
rect 2370 -3680 2410 -3675
rect 2370 -3705 2410 -3700
rect 2370 -3735 2375 -3705
rect 2375 -3735 2405 -3705
rect 2405 -3735 2410 -3705
rect 2370 -3740 2410 -3735
rect 2370 -3770 2410 -3765
rect 2370 -3800 2375 -3770
rect 2375 -3800 2405 -3770
rect 2405 -3800 2410 -3770
rect 2370 -3805 2410 -3800
rect 2370 -3840 2410 -3835
rect 2370 -3870 2375 -3840
rect 2375 -3870 2405 -3840
rect 2405 -3870 2410 -3840
rect 2370 -3875 2410 -3870
rect 2370 -3910 2410 -3905
rect 2370 -3940 2375 -3910
rect 2375 -3940 2405 -3910
rect 2405 -3940 2410 -3910
rect 2370 -3945 2410 -3940
rect 2370 -3980 2410 -3975
rect 2370 -4010 2375 -3980
rect 2375 -4010 2405 -3980
rect 2405 -4010 2410 -3980
rect 2370 -4015 2410 -4010
rect 2370 -4045 2410 -4040
rect 2370 -4075 2375 -4045
rect 2375 -4075 2405 -4045
rect 2405 -4075 2410 -4045
rect 2370 -4080 2410 -4075
rect 2370 -4105 2410 -4100
rect 2370 -4135 2375 -4105
rect 2375 -4135 2405 -4105
rect 2405 -4135 2410 -4105
rect 2370 -4140 2410 -4135
rect 2370 -4170 2410 -4165
rect 2370 -4200 2375 -4170
rect 2375 -4200 2405 -4170
rect 2405 -4200 2410 -4170
rect 2370 -4205 2410 -4200
rect 2370 -4240 2410 -4235
rect 2370 -4270 2375 -4240
rect 2375 -4270 2405 -4240
rect 2405 -4270 2410 -4240
rect 2370 -4275 2410 -4270
rect 2370 -4310 2410 -4305
rect 2370 -4340 2375 -4310
rect 2375 -4340 2405 -4310
rect 2405 -4340 2410 -4310
rect 2370 -4345 2410 -4340
rect 2370 -4380 2410 -4375
rect 2370 -4410 2375 -4380
rect 2375 -4410 2405 -4380
rect 2405 -4410 2410 -4380
rect 2370 -4415 2410 -4410
rect 2370 -4445 2410 -4440
rect 2370 -4475 2375 -4445
rect 2375 -4475 2405 -4445
rect 2405 -4475 2410 -4445
rect 2370 -4480 2410 -4475
rect 2720 -1305 2760 -1300
rect 2720 -1335 2725 -1305
rect 2725 -1335 2755 -1305
rect 2755 -1335 2760 -1305
rect 2720 -1340 2760 -1335
rect 2720 -1370 2760 -1365
rect 2720 -1400 2725 -1370
rect 2725 -1400 2755 -1370
rect 2755 -1400 2760 -1370
rect 2720 -1405 2760 -1400
rect 2720 -1440 2760 -1435
rect 2720 -1470 2725 -1440
rect 2725 -1470 2755 -1440
rect 2755 -1470 2760 -1440
rect 2720 -1475 2760 -1470
rect 2720 -1510 2760 -1505
rect 2720 -1540 2725 -1510
rect 2725 -1540 2755 -1510
rect 2755 -1540 2760 -1510
rect 2720 -1545 2760 -1540
rect 2720 -1580 2760 -1575
rect 2720 -1610 2725 -1580
rect 2725 -1610 2755 -1580
rect 2755 -1610 2760 -1580
rect 2720 -1615 2760 -1610
rect 2720 -1645 2760 -1640
rect 2720 -1675 2725 -1645
rect 2725 -1675 2755 -1645
rect 2755 -1675 2760 -1645
rect 2720 -1680 2760 -1675
rect 2720 -1705 2760 -1700
rect 2720 -1735 2725 -1705
rect 2725 -1735 2755 -1705
rect 2755 -1735 2760 -1705
rect 2720 -1740 2760 -1735
rect 2720 -1770 2760 -1765
rect 2720 -1800 2725 -1770
rect 2725 -1800 2755 -1770
rect 2755 -1800 2760 -1770
rect 2720 -1805 2760 -1800
rect 2720 -1840 2760 -1835
rect 2720 -1870 2725 -1840
rect 2725 -1870 2755 -1840
rect 2755 -1870 2760 -1840
rect 2720 -1875 2760 -1870
rect 2720 -1910 2760 -1905
rect 2720 -1940 2725 -1910
rect 2725 -1940 2755 -1910
rect 2755 -1940 2760 -1910
rect 2720 -1945 2760 -1940
rect 2720 -1980 2760 -1975
rect 2720 -2010 2725 -1980
rect 2725 -2010 2755 -1980
rect 2755 -2010 2760 -1980
rect 2720 -2015 2760 -2010
rect 2720 -2045 2760 -2040
rect 2720 -2075 2725 -2045
rect 2725 -2075 2755 -2045
rect 2755 -2075 2760 -2045
rect 2720 -2080 2760 -2075
rect 2720 -2105 2760 -2100
rect 2720 -2135 2725 -2105
rect 2725 -2135 2755 -2105
rect 2755 -2135 2760 -2105
rect 2720 -2140 2760 -2135
rect 2720 -2170 2760 -2165
rect 2720 -2200 2725 -2170
rect 2725 -2200 2755 -2170
rect 2755 -2200 2760 -2170
rect 2720 -2205 2760 -2200
rect 2720 -2240 2760 -2235
rect 2720 -2270 2725 -2240
rect 2725 -2270 2755 -2240
rect 2755 -2270 2760 -2240
rect 2720 -2275 2760 -2270
rect 2720 -2310 2760 -2305
rect 2720 -2340 2725 -2310
rect 2725 -2340 2755 -2310
rect 2755 -2340 2760 -2310
rect 2720 -2345 2760 -2340
rect 2720 -2380 2760 -2375
rect 2720 -2410 2725 -2380
rect 2725 -2410 2755 -2380
rect 2755 -2410 2760 -2380
rect 2720 -2415 2760 -2410
rect 2720 -2445 2760 -2440
rect 2720 -2475 2725 -2445
rect 2725 -2475 2755 -2445
rect 2755 -2475 2760 -2445
rect 2720 -2480 2760 -2475
rect 2720 -2505 2760 -2500
rect 2720 -2535 2725 -2505
rect 2725 -2535 2755 -2505
rect 2755 -2535 2760 -2505
rect 2720 -2540 2760 -2535
rect 2720 -2570 2760 -2565
rect 2720 -2600 2725 -2570
rect 2725 -2600 2755 -2570
rect 2755 -2600 2760 -2570
rect 2720 -2605 2760 -2600
rect 2720 -2640 2760 -2635
rect 2720 -2670 2725 -2640
rect 2725 -2670 2755 -2640
rect 2755 -2670 2760 -2640
rect 2720 -2675 2760 -2670
rect 2720 -2710 2760 -2705
rect 2720 -2740 2725 -2710
rect 2725 -2740 2755 -2710
rect 2755 -2740 2760 -2710
rect 2720 -2745 2760 -2740
rect 2720 -2780 2760 -2775
rect 2720 -2810 2725 -2780
rect 2725 -2810 2755 -2780
rect 2755 -2810 2760 -2780
rect 2720 -2815 2760 -2810
rect 2720 -2845 2760 -2840
rect 2720 -2875 2725 -2845
rect 2725 -2875 2755 -2845
rect 2755 -2875 2760 -2845
rect 2720 -2880 2760 -2875
rect 2720 -2905 2760 -2900
rect 2720 -2935 2725 -2905
rect 2725 -2935 2755 -2905
rect 2755 -2935 2760 -2905
rect 2720 -2940 2760 -2935
rect 2720 -2970 2760 -2965
rect 2720 -3000 2725 -2970
rect 2725 -3000 2755 -2970
rect 2755 -3000 2760 -2970
rect 2720 -3005 2760 -3000
rect 2720 -3040 2760 -3035
rect 2720 -3070 2725 -3040
rect 2725 -3070 2755 -3040
rect 2755 -3070 2760 -3040
rect 2720 -3075 2760 -3070
rect 2720 -3110 2760 -3105
rect 2720 -3140 2725 -3110
rect 2725 -3140 2755 -3110
rect 2755 -3140 2760 -3110
rect 2720 -3145 2760 -3140
rect 2720 -3180 2760 -3175
rect 2720 -3210 2725 -3180
rect 2725 -3210 2755 -3180
rect 2755 -3210 2760 -3180
rect 2720 -3215 2760 -3210
rect 2720 -3245 2760 -3240
rect 2720 -3275 2725 -3245
rect 2725 -3275 2755 -3245
rect 2755 -3275 2760 -3245
rect 2720 -3280 2760 -3275
rect 2720 -3305 2760 -3300
rect 2720 -3335 2725 -3305
rect 2725 -3335 2755 -3305
rect 2755 -3335 2760 -3305
rect 2720 -3340 2760 -3335
rect 2720 -3370 2760 -3365
rect 2720 -3400 2725 -3370
rect 2725 -3400 2755 -3370
rect 2755 -3400 2760 -3370
rect 2720 -3405 2760 -3400
rect 2720 -3440 2760 -3435
rect 2720 -3470 2725 -3440
rect 2725 -3470 2755 -3440
rect 2755 -3470 2760 -3440
rect 2720 -3475 2760 -3470
rect 2720 -3510 2760 -3505
rect 2720 -3540 2725 -3510
rect 2725 -3540 2755 -3510
rect 2755 -3540 2760 -3510
rect 2720 -3545 2760 -3540
rect 2720 -3580 2760 -3575
rect 2720 -3610 2725 -3580
rect 2725 -3610 2755 -3580
rect 2755 -3610 2760 -3580
rect 2720 -3615 2760 -3610
rect 2720 -3645 2760 -3640
rect 2720 -3675 2725 -3645
rect 2725 -3675 2755 -3645
rect 2755 -3675 2760 -3645
rect 2720 -3680 2760 -3675
rect 2720 -3705 2760 -3700
rect 2720 -3735 2725 -3705
rect 2725 -3735 2755 -3705
rect 2755 -3735 2760 -3705
rect 2720 -3740 2760 -3735
rect 2720 -3770 2760 -3765
rect 2720 -3800 2725 -3770
rect 2725 -3800 2755 -3770
rect 2755 -3800 2760 -3770
rect 2720 -3805 2760 -3800
rect 2720 -3840 2760 -3835
rect 2720 -3870 2725 -3840
rect 2725 -3870 2755 -3840
rect 2755 -3870 2760 -3840
rect 2720 -3875 2760 -3870
rect 2720 -3910 2760 -3905
rect 2720 -3940 2725 -3910
rect 2725 -3940 2755 -3910
rect 2755 -3940 2760 -3910
rect 2720 -3945 2760 -3940
rect 2720 -3980 2760 -3975
rect 2720 -4010 2725 -3980
rect 2725 -4010 2755 -3980
rect 2755 -4010 2760 -3980
rect 2720 -4015 2760 -4010
rect 2720 -4045 2760 -4040
rect 2720 -4075 2725 -4045
rect 2725 -4075 2755 -4045
rect 2755 -4075 2760 -4045
rect 2720 -4080 2760 -4075
rect 2720 -4105 2760 -4100
rect 2720 -4135 2725 -4105
rect 2725 -4135 2755 -4105
rect 2755 -4135 2760 -4105
rect 2720 -4140 2760 -4135
rect 2720 -4170 2760 -4165
rect 2720 -4200 2725 -4170
rect 2725 -4200 2755 -4170
rect 2755 -4200 2760 -4170
rect 2720 -4205 2760 -4200
rect 2720 -4240 2760 -4235
rect 2720 -4270 2725 -4240
rect 2725 -4270 2755 -4240
rect 2755 -4270 2760 -4240
rect 2720 -4275 2760 -4270
rect 2720 -4310 2760 -4305
rect 2720 -4340 2725 -4310
rect 2725 -4340 2755 -4310
rect 2755 -4340 2760 -4310
rect 2720 -4345 2760 -4340
rect 2720 -4380 2760 -4375
rect 2720 -4410 2725 -4380
rect 2725 -4410 2755 -4380
rect 2755 -4410 2760 -4380
rect 2720 -4415 2760 -4410
rect 2720 -4445 2760 -4440
rect 2720 -4475 2725 -4445
rect 2725 -4475 2755 -4445
rect 2755 -4475 2760 -4445
rect 2720 -4480 2760 -4475
rect 3070 -1305 3110 -1300
rect 3070 -1335 3075 -1305
rect 3075 -1335 3105 -1305
rect 3105 -1335 3110 -1305
rect 3070 -1340 3110 -1335
rect 3070 -1370 3110 -1365
rect 3070 -1400 3075 -1370
rect 3075 -1400 3105 -1370
rect 3105 -1400 3110 -1370
rect 3070 -1405 3110 -1400
rect 3070 -1440 3110 -1435
rect 3070 -1470 3075 -1440
rect 3075 -1470 3105 -1440
rect 3105 -1470 3110 -1440
rect 3070 -1475 3110 -1470
rect 3070 -1510 3110 -1505
rect 3070 -1540 3075 -1510
rect 3075 -1540 3105 -1510
rect 3105 -1540 3110 -1510
rect 3070 -1545 3110 -1540
rect 3070 -1580 3110 -1575
rect 3070 -1610 3075 -1580
rect 3075 -1610 3105 -1580
rect 3105 -1610 3110 -1580
rect 3070 -1615 3110 -1610
rect 3070 -1645 3110 -1640
rect 3070 -1675 3075 -1645
rect 3075 -1675 3105 -1645
rect 3105 -1675 3110 -1645
rect 3070 -1680 3110 -1675
rect 3070 -1705 3110 -1700
rect 3070 -1735 3075 -1705
rect 3075 -1735 3105 -1705
rect 3105 -1735 3110 -1705
rect 3070 -1740 3110 -1735
rect 3070 -1770 3110 -1765
rect 3070 -1800 3075 -1770
rect 3075 -1800 3105 -1770
rect 3105 -1800 3110 -1770
rect 3070 -1805 3110 -1800
rect 3070 -1840 3110 -1835
rect 3070 -1870 3075 -1840
rect 3075 -1870 3105 -1840
rect 3105 -1870 3110 -1840
rect 3070 -1875 3110 -1870
rect 3070 -1910 3110 -1905
rect 3070 -1940 3075 -1910
rect 3075 -1940 3105 -1910
rect 3105 -1940 3110 -1910
rect 3070 -1945 3110 -1940
rect 3070 -1980 3110 -1975
rect 3070 -2010 3075 -1980
rect 3075 -2010 3105 -1980
rect 3105 -2010 3110 -1980
rect 3070 -2015 3110 -2010
rect 3070 -2045 3110 -2040
rect 3070 -2075 3075 -2045
rect 3075 -2075 3105 -2045
rect 3105 -2075 3110 -2045
rect 3070 -2080 3110 -2075
rect 3070 -2105 3110 -2100
rect 3070 -2135 3075 -2105
rect 3075 -2135 3105 -2105
rect 3105 -2135 3110 -2105
rect 3070 -2140 3110 -2135
rect 3070 -2170 3110 -2165
rect 3070 -2200 3075 -2170
rect 3075 -2200 3105 -2170
rect 3105 -2200 3110 -2170
rect 3070 -2205 3110 -2200
rect 3070 -2240 3110 -2235
rect 3070 -2270 3075 -2240
rect 3075 -2270 3105 -2240
rect 3105 -2270 3110 -2240
rect 3070 -2275 3110 -2270
rect 3070 -2310 3110 -2305
rect 3070 -2340 3075 -2310
rect 3075 -2340 3105 -2310
rect 3105 -2340 3110 -2310
rect 3070 -2345 3110 -2340
rect 3070 -2380 3110 -2375
rect 3070 -2410 3075 -2380
rect 3075 -2410 3105 -2380
rect 3105 -2410 3110 -2380
rect 3070 -2415 3110 -2410
rect 3070 -2445 3110 -2440
rect 3070 -2475 3075 -2445
rect 3075 -2475 3105 -2445
rect 3105 -2475 3110 -2445
rect 3070 -2480 3110 -2475
rect 3070 -2505 3110 -2500
rect 3070 -2535 3075 -2505
rect 3075 -2535 3105 -2505
rect 3105 -2535 3110 -2505
rect 3070 -2540 3110 -2535
rect 3070 -2570 3110 -2565
rect 3070 -2600 3075 -2570
rect 3075 -2600 3105 -2570
rect 3105 -2600 3110 -2570
rect 3070 -2605 3110 -2600
rect 3070 -2640 3110 -2635
rect 3070 -2670 3075 -2640
rect 3075 -2670 3105 -2640
rect 3105 -2670 3110 -2640
rect 3070 -2675 3110 -2670
rect 3070 -2710 3110 -2705
rect 3070 -2740 3075 -2710
rect 3075 -2740 3105 -2710
rect 3105 -2740 3110 -2710
rect 3070 -2745 3110 -2740
rect 3070 -2780 3110 -2775
rect 3070 -2810 3075 -2780
rect 3075 -2810 3105 -2780
rect 3105 -2810 3110 -2780
rect 3070 -2815 3110 -2810
rect 3070 -2845 3110 -2840
rect 3070 -2875 3075 -2845
rect 3075 -2875 3105 -2845
rect 3105 -2875 3110 -2845
rect 3070 -2880 3110 -2875
rect 3070 -2905 3110 -2900
rect 3070 -2935 3075 -2905
rect 3075 -2935 3105 -2905
rect 3105 -2935 3110 -2905
rect 3070 -2940 3110 -2935
rect 3070 -2970 3110 -2965
rect 3070 -3000 3075 -2970
rect 3075 -3000 3105 -2970
rect 3105 -3000 3110 -2970
rect 3070 -3005 3110 -3000
rect 3070 -3040 3110 -3035
rect 3070 -3070 3075 -3040
rect 3075 -3070 3105 -3040
rect 3105 -3070 3110 -3040
rect 3070 -3075 3110 -3070
rect 3070 -3110 3110 -3105
rect 3070 -3140 3075 -3110
rect 3075 -3140 3105 -3110
rect 3105 -3140 3110 -3110
rect 3070 -3145 3110 -3140
rect 3070 -3180 3110 -3175
rect 3070 -3210 3075 -3180
rect 3075 -3210 3105 -3180
rect 3105 -3210 3110 -3180
rect 3070 -3215 3110 -3210
rect 3070 -3245 3110 -3240
rect 3070 -3275 3075 -3245
rect 3075 -3275 3105 -3245
rect 3105 -3275 3110 -3245
rect 3070 -3280 3110 -3275
rect 3070 -3305 3110 -3300
rect 3070 -3335 3075 -3305
rect 3075 -3335 3105 -3305
rect 3105 -3335 3110 -3305
rect 3070 -3340 3110 -3335
rect 3070 -3370 3110 -3365
rect 3070 -3400 3075 -3370
rect 3075 -3400 3105 -3370
rect 3105 -3400 3110 -3370
rect 3070 -3405 3110 -3400
rect 3070 -3440 3110 -3435
rect 3070 -3470 3075 -3440
rect 3075 -3470 3105 -3440
rect 3105 -3470 3110 -3440
rect 3070 -3475 3110 -3470
rect 3070 -3510 3110 -3505
rect 3070 -3540 3075 -3510
rect 3075 -3540 3105 -3510
rect 3105 -3540 3110 -3510
rect 3070 -3545 3110 -3540
rect 3070 -3580 3110 -3575
rect 3070 -3610 3075 -3580
rect 3075 -3610 3105 -3580
rect 3105 -3610 3110 -3580
rect 3070 -3615 3110 -3610
rect 3070 -3645 3110 -3640
rect 3070 -3675 3075 -3645
rect 3075 -3675 3105 -3645
rect 3105 -3675 3110 -3645
rect 3070 -3680 3110 -3675
rect 3070 -3705 3110 -3700
rect 3070 -3735 3075 -3705
rect 3075 -3735 3105 -3705
rect 3105 -3735 3110 -3705
rect 3070 -3740 3110 -3735
rect 3070 -3770 3110 -3765
rect 3070 -3800 3075 -3770
rect 3075 -3800 3105 -3770
rect 3105 -3800 3110 -3770
rect 3070 -3805 3110 -3800
rect 3070 -3840 3110 -3835
rect 3070 -3870 3075 -3840
rect 3075 -3870 3105 -3840
rect 3105 -3870 3110 -3840
rect 3070 -3875 3110 -3870
rect 3070 -3910 3110 -3905
rect 3070 -3940 3075 -3910
rect 3075 -3940 3105 -3910
rect 3105 -3940 3110 -3910
rect 3070 -3945 3110 -3940
rect 3070 -3980 3110 -3975
rect 3070 -4010 3075 -3980
rect 3075 -4010 3105 -3980
rect 3105 -4010 3110 -3980
rect 3070 -4015 3110 -4010
rect 3070 -4045 3110 -4040
rect 3070 -4075 3075 -4045
rect 3075 -4075 3105 -4045
rect 3105 -4075 3110 -4045
rect 3070 -4080 3110 -4075
rect 3070 -4105 3110 -4100
rect 3070 -4135 3075 -4105
rect 3075 -4135 3105 -4105
rect 3105 -4135 3110 -4105
rect 3070 -4140 3110 -4135
rect 3070 -4170 3110 -4165
rect 3070 -4200 3075 -4170
rect 3075 -4200 3105 -4170
rect 3105 -4200 3110 -4170
rect 3070 -4205 3110 -4200
rect 3070 -4240 3110 -4235
rect 3070 -4270 3075 -4240
rect 3075 -4270 3105 -4240
rect 3105 -4270 3110 -4240
rect 3070 -4275 3110 -4270
rect 3070 -4310 3110 -4305
rect 3070 -4340 3075 -4310
rect 3075 -4340 3105 -4310
rect 3105 -4340 3110 -4310
rect 3070 -4345 3110 -4340
rect 3070 -4380 3110 -4375
rect 3070 -4410 3075 -4380
rect 3075 -4410 3105 -4380
rect 3105 -4410 3110 -4380
rect 3070 -4415 3110 -4410
rect 3070 -4445 3110 -4440
rect 3070 -4475 3075 -4445
rect 3075 -4475 3105 -4445
rect 3105 -4475 3110 -4445
rect 3070 -4480 3110 -4475
rect 3420 -1305 3460 -1300
rect 3420 -1335 3425 -1305
rect 3425 -1335 3455 -1305
rect 3455 -1335 3460 -1305
rect 3420 -1340 3460 -1335
rect 3420 -1370 3460 -1365
rect 3420 -1400 3425 -1370
rect 3425 -1400 3455 -1370
rect 3455 -1400 3460 -1370
rect 3420 -1405 3460 -1400
rect 3420 -1440 3460 -1435
rect 3420 -1470 3425 -1440
rect 3425 -1470 3455 -1440
rect 3455 -1470 3460 -1440
rect 3420 -1475 3460 -1470
rect 3420 -1510 3460 -1505
rect 3420 -1540 3425 -1510
rect 3425 -1540 3455 -1510
rect 3455 -1540 3460 -1510
rect 3420 -1545 3460 -1540
rect 3420 -1580 3460 -1575
rect 3420 -1610 3425 -1580
rect 3425 -1610 3455 -1580
rect 3455 -1610 3460 -1580
rect 3420 -1615 3460 -1610
rect 3420 -1645 3460 -1640
rect 3420 -1675 3425 -1645
rect 3425 -1675 3455 -1645
rect 3455 -1675 3460 -1645
rect 3420 -1680 3460 -1675
rect 3420 -1705 3460 -1700
rect 3420 -1735 3425 -1705
rect 3425 -1735 3455 -1705
rect 3455 -1735 3460 -1705
rect 3420 -1740 3460 -1735
rect 3420 -1770 3460 -1765
rect 3420 -1800 3425 -1770
rect 3425 -1800 3455 -1770
rect 3455 -1800 3460 -1770
rect 3420 -1805 3460 -1800
rect 3420 -1840 3460 -1835
rect 3420 -1870 3425 -1840
rect 3425 -1870 3455 -1840
rect 3455 -1870 3460 -1840
rect 3420 -1875 3460 -1870
rect 3420 -1910 3460 -1905
rect 3420 -1940 3425 -1910
rect 3425 -1940 3455 -1910
rect 3455 -1940 3460 -1910
rect 3420 -1945 3460 -1940
rect 3420 -1980 3460 -1975
rect 3420 -2010 3425 -1980
rect 3425 -2010 3455 -1980
rect 3455 -2010 3460 -1980
rect 3420 -2015 3460 -2010
rect 3420 -2045 3460 -2040
rect 3420 -2075 3425 -2045
rect 3425 -2075 3455 -2045
rect 3455 -2075 3460 -2045
rect 3420 -2080 3460 -2075
rect 3420 -2105 3460 -2100
rect 3420 -2135 3425 -2105
rect 3425 -2135 3455 -2105
rect 3455 -2135 3460 -2105
rect 3420 -2140 3460 -2135
rect 3420 -2170 3460 -2165
rect 3420 -2200 3425 -2170
rect 3425 -2200 3455 -2170
rect 3455 -2200 3460 -2170
rect 3420 -2205 3460 -2200
rect 3420 -2240 3460 -2235
rect 3420 -2270 3425 -2240
rect 3425 -2270 3455 -2240
rect 3455 -2270 3460 -2240
rect 3420 -2275 3460 -2270
rect 3420 -2310 3460 -2305
rect 3420 -2340 3425 -2310
rect 3425 -2340 3455 -2310
rect 3455 -2340 3460 -2310
rect 3420 -2345 3460 -2340
rect 3420 -2380 3460 -2375
rect 3420 -2410 3425 -2380
rect 3425 -2410 3455 -2380
rect 3455 -2410 3460 -2380
rect 3420 -2415 3460 -2410
rect 3420 -2445 3460 -2440
rect 3420 -2475 3425 -2445
rect 3425 -2475 3455 -2445
rect 3455 -2475 3460 -2445
rect 3420 -2480 3460 -2475
rect 3420 -2505 3460 -2500
rect 3420 -2535 3425 -2505
rect 3425 -2535 3455 -2505
rect 3455 -2535 3460 -2505
rect 3420 -2540 3460 -2535
rect 3420 -2570 3460 -2565
rect 3420 -2600 3425 -2570
rect 3425 -2600 3455 -2570
rect 3455 -2600 3460 -2570
rect 3420 -2605 3460 -2600
rect 3420 -2640 3460 -2635
rect 3420 -2670 3425 -2640
rect 3425 -2670 3455 -2640
rect 3455 -2670 3460 -2640
rect 3420 -2675 3460 -2670
rect 3420 -2710 3460 -2705
rect 3420 -2740 3425 -2710
rect 3425 -2740 3455 -2710
rect 3455 -2740 3460 -2710
rect 3420 -2745 3460 -2740
rect 3420 -2780 3460 -2775
rect 3420 -2810 3425 -2780
rect 3425 -2810 3455 -2780
rect 3455 -2810 3460 -2780
rect 3420 -2815 3460 -2810
rect 3420 -2845 3460 -2840
rect 3420 -2875 3425 -2845
rect 3425 -2875 3455 -2845
rect 3455 -2875 3460 -2845
rect 3420 -2880 3460 -2875
rect 3420 -2905 3460 -2900
rect 3420 -2935 3425 -2905
rect 3425 -2935 3455 -2905
rect 3455 -2935 3460 -2905
rect 3420 -2940 3460 -2935
rect 3420 -2970 3460 -2965
rect 3420 -3000 3425 -2970
rect 3425 -3000 3455 -2970
rect 3455 -3000 3460 -2970
rect 3420 -3005 3460 -3000
rect 3420 -3040 3460 -3035
rect 3420 -3070 3425 -3040
rect 3425 -3070 3455 -3040
rect 3455 -3070 3460 -3040
rect 3420 -3075 3460 -3070
rect 3420 -3110 3460 -3105
rect 3420 -3140 3425 -3110
rect 3425 -3140 3455 -3110
rect 3455 -3140 3460 -3110
rect 3420 -3145 3460 -3140
rect 3420 -3180 3460 -3175
rect 3420 -3210 3425 -3180
rect 3425 -3210 3455 -3180
rect 3455 -3210 3460 -3180
rect 3420 -3215 3460 -3210
rect 3420 -3245 3460 -3240
rect 3420 -3275 3425 -3245
rect 3425 -3275 3455 -3245
rect 3455 -3275 3460 -3245
rect 3420 -3280 3460 -3275
rect 3420 -3305 3460 -3300
rect 3420 -3335 3425 -3305
rect 3425 -3335 3455 -3305
rect 3455 -3335 3460 -3305
rect 3420 -3340 3460 -3335
rect 3420 -3370 3460 -3365
rect 3420 -3400 3425 -3370
rect 3425 -3400 3455 -3370
rect 3455 -3400 3460 -3370
rect 3420 -3405 3460 -3400
rect 3420 -3440 3460 -3435
rect 3420 -3470 3425 -3440
rect 3425 -3470 3455 -3440
rect 3455 -3470 3460 -3440
rect 3420 -3475 3460 -3470
rect 3420 -3510 3460 -3505
rect 3420 -3540 3425 -3510
rect 3425 -3540 3455 -3510
rect 3455 -3540 3460 -3510
rect 3420 -3545 3460 -3540
rect 3420 -3580 3460 -3575
rect 3420 -3610 3425 -3580
rect 3425 -3610 3455 -3580
rect 3455 -3610 3460 -3580
rect 3420 -3615 3460 -3610
rect 3420 -3645 3460 -3640
rect 3420 -3675 3425 -3645
rect 3425 -3675 3455 -3645
rect 3455 -3675 3460 -3645
rect 3420 -3680 3460 -3675
rect 3420 -3705 3460 -3700
rect 3420 -3735 3425 -3705
rect 3425 -3735 3455 -3705
rect 3455 -3735 3460 -3705
rect 3420 -3740 3460 -3735
rect 3420 -3770 3460 -3765
rect 3420 -3800 3425 -3770
rect 3425 -3800 3455 -3770
rect 3455 -3800 3460 -3770
rect 3420 -3805 3460 -3800
rect 3420 -3840 3460 -3835
rect 3420 -3870 3425 -3840
rect 3425 -3870 3455 -3840
rect 3455 -3870 3460 -3840
rect 3420 -3875 3460 -3870
rect 3420 -3910 3460 -3905
rect 3420 -3940 3425 -3910
rect 3425 -3940 3455 -3910
rect 3455 -3940 3460 -3910
rect 3420 -3945 3460 -3940
rect 3420 -3980 3460 -3975
rect 3420 -4010 3425 -3980
rect 3425 -4010 3455 -3980
rect 3455 -4010 3460 -3980
rect 3420 -4015 3460 -4010
rect 3420 -4045 3460 -4040
rect 3420 -4075 3425 -4045
rect 3425 -4075 3455 -4045
rect 3455 -4075 3460 -4045
rect 3420 -4080 3460 -4075
rect 3420 -4105 3460 -4100
rect 3420 -4135 3425 -4105
rect 3425 -4135 3455 -4105
rect 3455 -4135 3460 -4105
rect 3420 -4140 3460 -4135
rect 3420 -4170 3460 -4165
rect 3420 -4200 3425 -4170
rect 3425 -4200 3455 -4170
rect 3455 -4200 3460 -4170
rect 3420 -4205 3460 -4200
rect 3420 -4240 3460 -4235
rect 3420 -4270 3425 -4240
rect 3425 -4270 3455 -4240
rect 3455 -4270 3460 -4240
rect 3420 -4275 3460 -4270
rect 3420 -4310 3460 -4305
rect 3420 -4340 3425 -4310
rect 3425 -4340 3455 -4310
rect 3455 -4340 3460 -4310
rect 3420 -4345 3460 -4340
rect 3420 -4380 3460 -4375
rect 3420 -4410 3425 -4380
rect 3425 -4410 3455 -4380
rect 3455 -4410 3460 -4380
rect 3420 -4415 3460 -4410
rect 3420 -4445 3460 -4440
rect 3420 -4475 3425 -4445
rect 3425 -4475 3455 -4445
rect 3455 -4475 3460 -4445
rect 3420 -4480 3460 -4475
rect 3770 -1305 3810 -1300
rect 3770 -1335 3775 -1305
rect 3775 -1335 3805 -1305
rect 3805 -1335 3810 -1305
rect 3770 -1340 3810 -1335
rect 3770 -1370 3810 -1365
rect 3770 -1400 3775 -1370
rect 3775 -1400 3805 -1370
rect 3805 -1400 3810 -1370
rect 3770 -1405 3810 -1400
rect 3770 -1440 3810 -1435
rect 3770 -1470 3775 -1440
rect 3775 -1470 3805 -1440
rect 3805 -1470 3810 -1440
rect 3770 -1475 3810 -1470
rect 3770 -1510 3810 -1505
rect 3770 -1540 3775 -1510
rect 3775 -1540 3805 -1510
rect 3805 -1540 3810 -1510
rect 3770 -1545 3810 -1540
rect 3770 -1580 3810 -1575
rect 3770 -1610 3775 -1580
rect 3775 -1610 3805 -1580
rect 3805 -1610 3810 -1580
rect 3770 -1615 3810 -1610
rect 3770 -1645 3810 -1640
rect 3770 -1675 3775 -1645
rect 3775 -1675 3805 -1645
rect 3805 -1675 3810 -1645
rect 3770 -1680 3810 -1675
rect 3770 -1705 3810 -1700
rect 3770 -1735 3775 -1705
rect 3775 -1735 3805 -1705
rect 3805 -1735 3810 -1705
rect 3770 -1740 3810 -1735
rect 3770 -1770 3810 -1765
rect 3770 -1800 3775 -1770
rect 3775 -1800 3805 -1770
rect 3805 -1800 3810 -1770
rect 3770 -1805 3810 -1800
rect 3770 -1840 3810 -1835
rect 3770 -1870 3775 -1840
rect 3775 -1870 3805 -1840
rect 3805 -1870 3810 -1840
rect 3770 -1875 3810 -1870
rect 3770 -1910 3810 -1905
rect 3770 -1940 3775 -1910
rect 3775 -1940 3805 -1910
rect 3805 -1940 3810 -1910
rect 3770 -1945 3810 -1940
rect 3770 -1980 3810 -1975
rect 3770 -2010 3775 -1980
rect 3775 -2010 3805 -1980
rect 3805 -2010 3810 -1980
rect 3770 -2015 3810 -2010
rect 3770 -2045 3810 -2040
rect 3770 -2075 3775 -2045
rect 3775 -2075 3805 -2045
rect 3805 -2075 3810 -2045
rect 3770 -2080 3810 -2075
rect 3770 -2105 3810 -2100
rect 3770 -2135 3775 -2105
rect 3775 -2135 3805 -2105
rect 3805 -2135 3810 -2105
rect 3770 -2140 3810 -2135
rect 3770 -2170 3810 -2165
rect 3770 -2200 3775 -2170
rect 3775 -2200 3805 -2170
rect 3805 -2200 3810 -2170
rect 3770 -2205 3810 -2200
rect 3770 -2240 3810 -2235
rect 3770 -2270 3775 -2240
rect 3775 -2270 3805 -2240
rect 3805 -2270 3810 -2240
rect 3770 -2275 3810 -2270
rect 3770 -2310 3810 -2305
rect 3770 -2340 3775 -2310
rect 3775 -2340 3805 -2310
rect 3805 -2340 3810 -2310
rect 3770 -2345 3810 -2340
rect 3770 -2380 3810 -2375
rect 3770 -2410 3775 -2380
rect 3775 -2410 3805 -2380
rect 3805 -2410 3810 -2380
rect 3770 -2415 3810 -2410
rect 3770 -2445 3810 -2440
rect 3770 -2475 3775 -2445
rect 3775 -2475 3805 -2445
rect 3805 -2475 3810 -2445
rect 3770 -2480 3810 -2475
rect 3770 -2505 3810 -2500
rect 3770 -2535 3775 -2505
rect 3775 -2535 3805 -2505
rect 3805 -2535 3810 -2505
rect 3770 -2540 3810 -2535
rect 3770 -2570 3810 -2565
rect 3770 -2600 3775 -2570
rect 3775 -2600 3805 -2570
rect 3805 -2600 3810 -2570
rect 3770 -2605 3810 -2600
rect 3770 -2640 3810 -2635
rect 3770 -2670 3775 -2640
rect 3775 -2670 3805 -2640
rect 3805 -2670 3810 -2640
rect 3770 -2675 3810 -2670
rect 3770 -2710 3810 -2705
rect 3770 -2740 3775 -2710
rect 3775 -2740 3805 -2710
rect 3805 -2740 3810 -2710
rect 3770 -2745 3810 -2740
rect 3770 -2780 3810 -2775
rect 3770 -2810 3775 -2780
rect 3775 -2810 3805 -2780
rect 3805 -2810 3810 -2780
rect 3770 -2815 3810 -2810
rect 3770 -2845 3810 -2840
rect 3770 -2875 3775 -2845
rect 3775 -2875 3805 -2845
rect 3805 -2875 3810 -2845
rect 3770 -2880 3810 -2875
rect 3770 -2905 3810 -2900
rect 3770 -2935 3775 -2905
rect 3775 -2935 3805 -2905
rect 3805 -2935 3810 -2905
rect 3770 -2940 3810 -2935
rect 3770 -2970 3810 -2965
rect 3770 -3000 3775 -2970
rect 3775 -3000 3805 -2970
rect 3805 -3000 3810 -2970
rect 3770 -3005 3810 -3000
rect 3770 -3040 3810 -3035
rect 3770 -3070 3775 -3040
rect 3775 -3070 3805 -3040
rect 3805 -3070 3810 -3040
rect 3770 -3075 3810 -3070
rect 3770 -3110 3810 -3105
rect 3770 -3140 3775 -3110
rect 3775 -3140 3805 -3110
rect 3805 -3140 3810 -3110
rect 3770 -3145 3810 -3140
rect 3770 -3180 3810 -3175
rect 3770 -3210 3775 -3180
rect 3775 -3210 3805 -3180
rect 3805 -3210 3810 -3180
rect 3770 -3215 3810 -3210
rect 3770 -3245 3810 -3240
rect 3770 -3275 3775 -3245
rect 3775 -3275 3805 -3245
rect 3805 -3275 3810 -3245
rect 3770 -3280 3810 -3275
rect 3770 -3305 3810 -3300
rect 3770 -3335 3775 -3305
rect 3775 -3335 3805 -3305
rect 3805 -3335 3810 -3305
rect 3770 -3340 3810 -3335
rect 3770 -3370 3810 -3365
rect 3770 -3400 3775 -3370
rect 3775 -3400 3805 -3370
rect 3805 -3400 3810 -3370
rect 3770 -3405 3810 -3400
rect 3770 -3440 3810 -3435
rect 3770 -3470 3775 -3440
rect 3775 -3470 3805 -3440
rect 3805 -3470 3810 -3440
rect 3770 -3475 3810 -3470
rect 3770 -3510 3810 -3505
rect 3770 -3540 3775 -3510
rect 3775 -3540 3805 -3510
rect 3805 -3540 3810 -3510
rect 3770 -3545 3810 -3540
rect 3770 -3580 3810 -3575
rect 3770 -3610 3775 -3580
rect 3775 -3610 3805 -3580
rect 3805 -3610 3810 -3580
rect 3770 -3615 3810 -3610
rect 3770 -3645 3810 -3640
rect 3770 -3675 3775 -3645
rect 3775 -3675 3805 -3645
rect 3805 -3675 3810 -3645
rect 3770 -3680 3810 -3675
rect 3770 -3705 3810 -3700
rect 3770 -3735 3775 -3705
rect 3775 -3735 3805 -3705
rect 3805 -3735 3810 -3705
rect 3770 -3740 3810 -3735
rect 3770 -3770 3810 -3765
rect 3770 -3800 3775 -3770
rect 3775 -3800 3805 -3770
rect 3805 -3800 3810 -3770
rect 3770 -3805 3810 -3800
rect 3770 -3840 3810 -3835
rect 3770 -3870 3775 -3840
rect 3775 -3870 3805 -3840
rect 3805 -3870 3810 -3840
rect 3770 -3875 3810 -3870
rect 3770 -3910 3810 -3905
rect 3770 -3940 3775 -3910
rect 3775 -3940 3805 -3910
rect 3805 -3940 3810 -3910
rect 3770 -3945 3810 -3940
rect 3770 -3980 3810 -3975
rect 3770 -4010 3775 -3980
rect 3775 -4010 3805 -3980
rect 3805 -4010 3810 -3980
rect 3770 -4015 3810 -4010
rect 3770 -4045 3810 -4040
rect 3770 -4075 3775 -4045
rect 3775 -4075 3805 -4045
rect 3805 -4075 3810 -4045
rect 3770 -4080 3810 -4075
rect 3770 -4105 3810 -4100
rect 3770 -4135 3775 -4105
rect 3775 -4135 3805 -4105
rect 3805 -4135 3810 -4105
rect 3770 -4140 3810 -4135
rect 3770 -4170 3810 -4165
rect 3770 -4200 3775 -4170
rect 3775 -4200 3805 -4170
rect 3805 -4200 3810 -4170
rect 3770 -4205 3810 -4200
rect 3770 -4240 3810 -4235
rect 3770 -4270 3775 -4240
rect 3775 -4270 3805 -4240
rect 3805 -4270 3810 -4240
rect 3770 -4275 3810 -4270
rect 3770 -4310 3810 -4305
rect 3770 -4340 3775 -4310
rect 3775 -4340 3805 -4310
rect 3805 -4340 3810 -4310
rect 3770 -4345 3810 -4340
rect 3770 -4380 3810 -4375
rect 3770 -4410 3775 -4380
rect 3775 -4410 3805 -4380
rect 3805 -4410 3810 -4380
rect 3770 -4415 3810 -4410
rect 3770 -4445 3810 -4440
rect 3770 -4475 3775 -4445
rect 3775 -4475 3805 -4445
rect 3805 -4475 3810 -4445
rect 3770 -4480 3810 -4475
rect 4120 -1305 4160 -1300
rect 4120 -1335 4125 -1305
rect 4125 -1335 4155 -1305
rect 4155 -1335 4160 -1305
rect 4120 -1340 4160 -1335
rect 4120 -1370 4160 -1365
rect 4120 -1400 4125 -1370
rect 4125 -1400 4155 -1370
rect 4155 -1400 4160 -1370
rect 4120 -1405 4160 -1400
rect 4120 -1440 4160 -1435
rect 4120 -1470 4125 -1440
rect 4125 -1470 4155 -1440
rect 4155 -1470 4160 -1440
rect 4120 -1475 4160 -1470
rect 4120 -1510 4160 -1505
rect 4120 -1540 4125 -1510
rect 4125 -1540 4155 -1510
rect 4155 -1540 4160 -1510
rect 4120 -1545 4160 -1540
rect 4120 -1580 4160 -1575
rect 4120 -1610 4125 -1580
rect 4125 -1610 4155 -1580
rect 4155 -1610 4160 -1580
rect 4120 -1615 4160 -1610
rect 4120 -1645 4160 -1640
rect 4120 -1675 4125 -1645
rect 4125 -1675 4155 -1645
rect 4155 -1675 4160 -1645
rect 4120 -1680 4160 -1675
rect 4120 -1705 4160 -1700
rect 4120 -1735 4125 -1705
rect 4125 -1735 4155 -1705
rect 4155 -1735 4160 -1705
rect 4120 -1740 4160 -1735
rect 4120 -1770 4160 -1765
rect 4120 -1800 4125 -1770
rect 4125 -1800 4155 -1770
rect 4155 -1800 4160 -1770
rect 4120 -1805 4160 -1800
rect 4120 -1840 4160 -1835
rect 4120 -1870 4125 -1840
rect 4125 -1870 4155 -1840
rect 4155 -1870 4160 -1840
rect 4120 -1875 4160 -1870
rect 4120 -1910 4160 -1905
rect 4120 -1940 4125 -1910
rect 4125 -1940 4155 -1910
rect 4155 -1940 4160 -1910
rect 4120 -1945 4160 -1940
rect 4120 -1980 4160 -1975
rect 4120 -2010 4125 -1980
rect 4125 -2010 4155 -1980
rect 4155 -2010 4160 -1980
rect 4120 -2015 4160 -2010
rect 4120 -2045 4160 -2040
rect 4120 -2075 4125 -2045
rect 4125 -2075 4155 -2045
rect 4155 -2075 4160 -2045
rect 4120 -2080 4160 -2075
rect 4120 -2105 4160 -2100
rect 4120 -2135 4125 -2105
rect 4125 -2135 4155 -2105
rect 4155 -2135 4160 -2105
rect 4120 -2140 4160 -2135
rect 4120 -2170 4160 -2165
rect 4120 -2200 4125 -2170
rect 4125 -2200 4155 -2170
rect 4155 -2200 4160 -2170
rect 4120 -2205 4160 -2200
rect 4120 -2240 4160 -2235
rect 4120 -2270 4125 -2240
rect 4125 -2270 4155 -2240
rect 4155 -2270 4160 -2240
rect 4120 -2275 4160 -2270
rect 4120 -2310 4160 -2305
rect 4120 -2340 4125 -2310
rect 4125 -2340 4155 -2310
rect 4155 -2340 4160 -2310
rect 4120 -2345 4160 -2340
rect 4120 -2380 4160 -2375
rect 4120 -2410 4125 -2380
rect 4125 -2410 4155 -2380
rect 4155 -2410 4160 -2380
rect 4120 -2415 4160 -2410
rect 4120 -2445 4160 -2440
rect 4120 -2475 4125 -2445
rect 4125 -2475 4155 -2445
rect 4155 -2475 4160 -2445
rect 4120 -2480 4160 -2475
rect 4120 -2505 4160 -2500
rect 4120 -2535 4125 -2505
rect 4125 -2535 4155 -2505
rect 4155 -2535 4160 -2505
rect 4120 -2540 4160 -2535
rect 4120 -2570 4160 -2565
rect 4120 -2600 4125 -2570
rect 4125 -2600 4155 -2570
rect 4155 -2600 4160 -2570
rect 4120 -2605 4160 -2600
rect 4120 -2640 4160 -2635
rect 4120 -2670 4125 -2640
rect 4125 -2670 4155 -2640
rect 4155 -2670 4160 -2640
rect 4120 -2675 4160 -2670
rect 4120 -2710 4160 -2705
rect 4120 -2740 4125 -2710
rect 4125 -2740 4155 -2710
rect 4155 -2740 4160 -2710
rect 4120 -2745 4160 -2740
rect 4120 -2780 4160 -2775
rect 4120 -2810 4125 -2780
rect 4125 -2810 4155 -2780
rect 4155 -2810 4160 -2780
rect 4120 -2815 4160 -2810
rect 4120 -2845 4160 -2840
rect 4120 -2875 4125 -2845
rect 4125 -2875 4155 -2845
rect 4155 -2875 4160 -2845
rect 4120 -2880 4160 -2875
rect 4120 -2905 4160 -2900
rect 4120 -2935 4125 -2905
rect 4125 -2935 4155 -2905
rect 4155 -2935 4160 -2905
rect 4120 -2940 4160 -2935
rect 4120 -2970 4160 -2965
rect 4120 -3000 4125 -2970
rect 4125 -3000 4155 -2970
rect 4155 -3000 4160 -2970
rect 4120 -3005 4160 -3000
rect 4120 -3040 4160 -3035
rect 4120 -3070 4125 -3040
rect 4125 -3070 4155 -3040
rect 4155 -3070 4160 -3040
rect 4120 -3075 4160 -3070
rect 4120 -3110 4160 -3105
rect 4120 -3140 4125 -3110
rect 4125 -3140 4155 -3110
rect 4155 -3140 4160 -3110
rect 4120 -3145 4160 -3140
rect 4120 -3180 4160 -3175
rect 4120 -3210 4125 -3180
rect 4125 -3210 4155 -3180
rect 4155 -3210 4160 -3180
rect 4120 -3215 4160 -3210
rect 4120 -3245 4160 -3240
rect 4120 -3275 4125 -3245
rect 4125 -3275 4155 -3245
rect 4155 -3275 4160 -3245
rect 4120 -3280 4160 -3275
rect 4120 -3305 4160 -3300
rect 4120 -3335 4125 -3305
rect 4125 -3335 4155 -3305
rect 4155 -3335 4160 -3305
rect 4120 -3340 4160 -3335
rect 4120 -3370 4160 -3365
rect 4120 -3400 4125 -3370
rect 4125 -3400 4155 -3370
rect 4155 -3400 4160 -3370
rect 4120 -3405 4160 -3400
rect 4120 -3440 4160 -3435
rect 4120 -3470 4125 -3440
rect 4125 -3470 4155 -3440
rect 4155 -3470 4160 -3440
rect 4120 -3475 4160 -3470
rect 4120 -3510 4160 -3505
rect 4120 -3540 4125 -3510
rect 4125 -3540 4155 -3510
rect 4155 -3540 4160 -3510
rect 4120 -3545 4160 -3540
rect 4120 -3580 4160 -3575
rect 4120 -3610 4125 -3580
rect 4125 -3610 4155 -3580
rect 4155 -3610 4160 -3580
rect 4120 -3615 4160 -3610
rect 4120 -3645 4160 -3640
rect 4120 -3675 4125 -3645
rect 4125 -3675 4155 -3645
rect 4155 -3675 4160 -3645
rect 4120 -3680 4160 -3675
rect 4120 -3705 4160 -3700
rect 4120 -3735 4125 -3705
rect 4125 -3735 4155 -3705
rect 4155 -3735 4160 -3705
rect 4120 -3740 4160 -3735
rect 4120 -3770 4160 -3765
rect 4120 -3800 4125 -3770
rect 4125 -3800 4155 -3770
rect 4155 -3800 4160 -3770
rect 4120 -3805 4160 -3800
rect 4120 -3840 4160 -3835
rect 4120 -3870 4125 -3840
rect 4125 -3870 4155 -3840
rect 4155 -3870 4160 -3840
rect 4120 -3875 4160 -3870
rect 4120 -3910 4160 -3905
rect 4120 -3940 4125 -3910
rect 4125 -3940 4155 -3910
rect 4155 -3940 4160 -3910
rect 4120 -3945 4160 -3940
rect 4120 -3980 4160 -3975
rect 4120 -4010 4125 -3980
rect 4125 -4010 4155 -3980
rect 4155 -4010 4160 -3980
rect 4120 -4015 4160 -4010
rect 4120 -4045 4160 -4040
rect 4120 -4075 4125 -4045
rect 4125 -4075 4155 -4045
rect 4155 -4075 4160 -4045
rect 4120 -4080 4160 -4075
rect 4120 -4105 4160 -4100
rect 4120 -4135 4125 -4105
rect 4125 -4135 4155 -4105
rect 4155 -4135 4160 -4105
rect 4120 -4140 4160 -4135
rect 4120 -4170 4160 -4165
rect 4120 -4200 4125 -4170
rect 4125 -4200 4155 -4170
rect 4155 -4200 4160 -4170
rect 4120 -4205 4160 -4200
rect 4120 -4240 4160 -4235
rect 4120 -4270 4125 -4240
rect 4125 -4270 4155 -4240
rect 4155 -4270 4160 -4240
rect 4120 -4275 4160 -4270
rect 4120 -4310 4160 -4305
rect 4120 -4340 4125 -4310
rect 4125 -4340 4155 -4310
rect 4155 -4340 4160 -4310
rect 4120 -4345 4160 -4340
rect 4120 -4380 4160 -4375
rect 4120 -4410 4125 -4380
rect 4125 -4410 4155 -4380
rect 4155 -4410 4160 -4380
rect 4120 -4415 4160 -4410
rect 4120 -4445 4160 -4440
rect 4120 -4475 4125 -4445
rect 4125 -4475 4155 -4445
rect 4155 -4475 4160 -4445
rect 4120 -4480 4160 -4475
rect 4470 -1305 4510 -1300
rect 4470 -1335 4475 -1305
rect 4475 -1335 4505 -1305
rect 4505 -1335 4510 -1305
rect 4470 -1340 4510 -1335
rect 4470 -1370 4510 -1365
rect 4470 -1400 4475 -1370
rect 4475 -1400 4505 -1370
rect 4505 -1400 4510 -1370
rect 4470 -1405 4510 -1400
rect 4470 -1440 4510 -1435
rect 4470 -1470 4475 -1440
rect 4475 -1470 4505 -1440
rect 4505 -1470 4510 -1440
rect 4470 -1475 4510 -1470
rect 4470 -1510 4510 -1505
rect 4470 -1540 4475 -1510
rect 4475 -1540 4505 -1510
rect 4505 -1540 4510 -1510
rect 4470 -1545 4510 -1540
rect 4470 -1580 4510 -1575
rect 4470 -1610 4475 -1580
rect 4475 -1610 4505 -1580
rect 4505 -1610 4510 -1580
rect 4470 -1615 4510 -1610
rect 4470 -1645 4510 -1640
rect 4470 -1675 4475 -1645
rect 4475 -1675 4505 -1645
rect 4505 -1675 4510 -1645
rect 4470 -1680 4510 -1675
rect 4470 -1705 4510 -1700
rect 4470 -1735 4475 -1705
rect 4475 -1735 4505 -1705
rect 4505 -1735 4510 -1705
rect 4470 -1740 4510 -1735
rect 4470 -1770 4510 -1765
rect 4470 -1800 4475 -1770
rect 4475 -1800 4505 -1770
rect 4505 -1800 4510 -1770
rect 4470 -1805 4510 -1800
rect 4470 -1840 4510 -1835
rect 4470 -1870 4475 -1840
rect 4475 -1870 4505 -1840
rect 4505 -1870 4510 -1840
rect 4470 -1875 4510 -1870
rect 4470 -1910 4510 -1905
rect 4470 -1940 4475 -1910
rect 4475 -1940 4505 -1910
rect 4505 -1940 4510 -1910
rect 4470 -1945 4510 -1940
rect 4470 -1980 4510 -1975
rect 4470 -2010 4475 -1980
rect 4475 -2010 4505 -1980
rect 4505 -2010 4510 -1980
rect 4470 -2015 4510 -2010
rect 4470 -2045 4510 -2040
rect 4470 -2075 4475 -2045
rect 4475 -2075 4505 -2045
rect 4505 -2075 4510 -2045
rect 4470 -2080 4510 -2075
rect 4470 -2105 4510 -2100
rect 4470 -2135 4475 -2105
rect 4475 -2135 4505 -2105
rect 4505 -2135 4510 -2105
rect 4470 -2140 4510 -2135
rect 4470 -2170 4510 -2165
rect 4470 -2200 4475 -2170
rect 4475 -2200 4505 -2170
rect 4505 -2200 4510 -2170
rect 4470 -2205 4510 -2200
rect 4470 -2240 4510 -2235
rect 4470 -2270 4475 -2240
rect 4475 -2270 4505 -2240
rect 4505 -2270 4510 -2240
rect 4470 -2275 4510 -2270
rect 4470 -2310 4510 -2305
rect 4470 -2340 4475 -2310
rect 4475 -2340 4505 -2310
rect 4505 -2340 4510 -2310
rect 4470 -2345 4510 -2340
rect 4470 -2380 4510 -2375
rect 4470 -2410 4475 -2380
rect 4475 -2410 4505 -2380
rect 4505 -2410 4510 -2380
rect 4470 -2415 4510 -2410
rect 4470 -2445 4510 -2440
rect 4470 -2475 4475 -2445
rect 4475 -2475 4505 -2445
rect 4505 -2475 4510 -2445
rect 4470 -2480 4510 -2475
rect 4470 -2505 4510 -2500
rect 4470 -2535 4475 -2505
rect 4475 -2535 4505 -2505
rect 4505 -2535 4510 -2505
rect 4470 -2540 4510 -2535
rect 4470 -2570 4510 -2565
rect 4470 -2600 4475 -2570
rect 4475 -2600 4505 -2570
rect 4505 -2600 4510 -2570
rect 4470 -2605 4510 -2600
rect 4470 -2640 4510 -2635
rect 4470 -2670 4475 -2640
rect 4475 -2670 4505 -2640
rect 4505 -2670 4510 -2640
rect 4470 -2675 4510 -2670
rect 4470 -2710 4510 -2705
rect 4470 -2740 4475 -2710
rect 4475 -2740 4505 -2710
rect 4505 -2740 4510 -2710
rect 4470 -2745 4510 -2740
rect 4470 -2780 4510 -2775
rect 4470 -2810 4475 -2780
rect 4475 -2810 4505 -2780
rect 4505 -2810 4510 -2780
rect 4470 -2815 4510 -2810
rect 4470 -2845 4510 -2840
rect 4470 -2875 4475 -2845
rect 4475 -2875 4505 -2845
rect 4505 -2875 4510 -2845
rect 4470 -2880 4510 -2875
rect 4470 -2905 4510 -2900
rect 4470 -2935 4475 -2905
rect 4475 -2935 4505 -2905
rect 4505 -2935 4510 -2905
rect 4470 -2940 4510 -2935
rect 4470 -2970 4510 -2965
rect 4470 -3000 4475 -2970
rect 4475 -3000 4505 -2970
rect 4505 -3000 4510 -2970
rect 4470 -3005 4510 -3000
rect 4470 -3040 4510 -3035
rect 4470 -3070 4475 -3040
rect 4475 -3070 4505 -3040
rect 4505 -3070 4510 -3040
rect 4470 -3075 4510 -3070
rect 4470 -3110 4510 -3105
rect 4470 -3140 4475 -3110
rect 4475 -3140 4505 -3110
rect 4505 -3140 4510 -3110
rect 4470 -3145 4510 -3140
rect 4470 -3180 4510 -3175
rect 4470 -3210 4475 -3180
rect 4475 -3210 4505 -3180
rect 4505 -3210 4510 -3180
rect 4470 -3215 4510 -3210
rect 4470 -3245 4510 -3240
rect 4470 -3275 4475 -3245
rect 4475 -3275 4505 -3245
rect 4505 -3275 4510 -3245
rect 4470 -3280 4510 -3275
rect 4470 -3305 4510 -3300
rect 4470 -3335 4475 -3305
rect 4475 -3335 4505 -3305
rect 4505 -3335 4510 -3305
rect 4470 -3340 4510 -3335
rect 4470 -3370 4510 -3365
rect 4470 -3400 4475 -3370
rect 4475 -3400 4505 -3370
rect 4505 -3400 4510 -3370
rect 4470 -3405 4510 -3400
rect 4470 -3440 4510 -3435
rect 4470 -3470 4475 -3440
rect 4475 -3470 4505 -3440
rect 4505 -3470 4510 -3440
rect 4470 -3475 4510 -3470
rect 4470 -3510 4510 -3505
rect 4470 -3540 4475 -3510
rect 4475 -3540 4505 -3510
rect 4505 -3540 4510 -3510
rect 4470 -3545 4510 -3540
rect 4470 -3580 4510 -3575
rect 4470 -3610 4475 -3580
rect 4475 -3610 4505 -3580
rect 4505 -3610 4510 -3580
rect 4470 -3615 4510 -3610
rect 4470 -3645 4510 -3640
rect 4470 -3675 4475 -3645
rect 4475 -3675 4505 -3645
rect 4505 -3675 4510 -3645
rect 4470 -3680 4510 -3675
rect 4470 -3705 4510 -3700
rect 4470 -3735 4475 -3705
rect 4475 -3735 4505 -3705
rect 4505 -3735 4510 -3705
rect 4470 -3740 4510 -3735
rect 4470 -3770 4510 -3765
rect 4470 -3800 4475 -3770
rect 4475 -3800 4505 -3770
rect 4505 -3800 4510 -3770
rect 4470 -3805 4510 -3800
rect 4470 -3840 4510 -3835
rect 4470 -3870 4475 -3840
rect 4475 -3870 4505 -3840
rect 4505 -3870 4510 -3840
rect 4470 -3875 4510 -3870
rect 4470 -3910 4510 -3905
rect 4470 -3940 4475 -3910
rect 4475 -3940 4505 -3910
rect 4505 -3940 4510 -3910
rect 4470 -3945 4510 -3940
rect 4470 -3980 4510 -3975
rect 4470 -4010 4475 -3980
rect 4475 -4010 4505 -3980
rect 4505 -4010 4510 -3980
rect 4470 -4015 4510 -4010
rect 4470 -4045 4510 -4040
rect 4470 -4075 4475 -4045
rect 4475 -4075 4505 -4045
rect 4505 -4075 4510 -4045
rect 4470 -4080 4510 -4075
rect 4470 -4105 4510 -4100
rect 4470 -4135 4475 -4105
rect 4475 -4135 4505 -4105
rect 4505 -4135 4510 -4105
rect 4470 -4140 4510 -4135
rect 4470 -4170 4510 -4165
rect 4470 -4200 4475 -4170
rect 4475 -4200 4505 -4170
rect 4505 -4200 4510 -4170
rect 4470 -4205 4510 -4200
rect 4470 -4240 4510 -4235
rect 4470 -4270 4475 -4240
rect 4475 -4270 4505 -4240
rect 4505 -4270 4510 -4240
rect 4470 -4275 4510 -4270
rect 4470 -4310 4510 -4305
rect 4470 -4340 4475 -4310
rect 4475 -4340 4505 -4310
rect 4505 -4340 4510 -4310
rect 4470 -4345 4510 -4340
rect 4470 -4380 4510 -4375
rect 4470 -4410 4475 -4380
rect 4475 -4410 4505 -4380
rect 4505 -4410 4510 -4380
rect 4470 -4415 4510 -4410
rect 4470 -4445 4510 -4440
rect 4470 -4475 4475 -4445
rect 4475 -4475 4505 -4445
rect 4505 -4475 4510 -4445
rect 4470 -4480 4510 -4475
rect 4820 -1305 4860 -1300
rect 4820 -1335 4825 -1305
rect 4825 -1335 4855 -1305
rect 4855 -1335 4860 -1305
rect 4820 -1340 4860 -1335
rect 4820 -1370 4860 -1365
rect 4820 -1400 4825 -1370
rect 4825 -1400 4855 -1370
rect 4855 -1400 4860 -1370
rect 4820 -1405 4860 -1400
rect 4820 -1440 4860 -1435
rect 4820 -1470 4825 -1440
rect 4825 -1470 4855 -1440
rect 4855 -1470 4860 -1440
rect 4820 -1475 4860 -1470
rect 4820 -1510 4860 -1505
rect 4820 -1540 4825 -1510
rect 4825 -1540 4855 -1510
rect 4855 -1540 4860 -1510
rect 4820 -1545 4860 -1540
rect 4820 -1580 4860 -1575
rect 4820 -1610 4825 -1580
rect 4825 -1610 4855 -1580
rect 4855 -1610 4860 -1580
rect 4820 -1615 4860 -1610
rect 4820 -1645 4860 -1640
rect 4820 -1675 4825 -1645
rect 4825 -1675 4855 -1645
rect 4855 -1675 4860 -1645
rect 4820 -1680 4860 -1675
rect 4820 -1705 4860 -1700
rect 4820 -1735 4825 -1705
rect 4825 -1735 4855 -1705
rect 4855 -1735 4860 -1705
rect 4820 -1740 4860 -1735
rect 4820 -1770 4860 -1765
rect 4820 -1800 4825 -1770
rect 4825 -1800 4855 -1770
rect 4855 -1800 4860 -1770
rect 4820 -1805 4860 -1800
rect 4820 -1840 4860 -1835
rect 4820 -1870 4825 -1840
rect 4825 -1870 4855 -1840
rect 4855 -1870 4860 -1840
rect 4820 -1875 4860 -1870
rect 4820 -1910 4860 -1905
rect 4820 -1940 4825 -1910
rect 4825 -1940 4855 -1910
rect 4855 -1940 4860 -1910
rect 4820 -1945 4860 -1940
rect 4820 -1980 4860 -1975
rect 4820 -2010 4825 -1980
rect 4825 -2010 4855 -1980
rect 4855 -2010 4860 -1980
rect 4820 -2015 4860 -2010
rect 4820 -2045 4860 -2040
rect 4820 -2075 4825 -2045
rect 4825 -2075 4855 -2045
rect 4855 -2075 4860 -2045
rect 4820 -2080 4860 -2075
rect 4820 -2105 4860 -2100
rect 4820 -2135 4825 -2105
rect 4825 -2135 4855 -2105
rect 4855 -2135 4860 -2105
rect 4820 -2140 4860 -2135
rect 4820 -2170 4860 -2165
rect 4820 -2200 4825 -2170
rect 4825 -2200 4855 -2170
rect 4855 -2200 4860 -2170
rect 4820 -2205 4860 -2200
rect 4820 -2240 4860 -2235
rect 4820 -2270 4825 -2240
rect 4825 -2270 4855 -2240
rect 4855 -2270 4860 -2240
rect 4820 -2275 4860 -2270
rect 4820 -2310 4860 -2305
rect 4820 -2340 4825 -2310
rect 4825 -2340 4855 -2310
rect 4855 -2340 4860 -2310
rect 4820 -2345 4860 -2340
rect 4820 -2380 4860 -2375
rect 4820 -2410 4825 -2380
rect 4825 -2410 4855 -2380
rect 4855 -2410 4860 -2380
rect 4820 -2415 4860 -2410
rect 4820 -2445 4860 -2440
rect 4820 -2475 4825 -2445
rect 4825 -2475 4855 -2445
rect 4855 -2475 4860 -2445
rect 4820 -2480 4860 -2475
rect 4820 -2505 4860 -2500
rect 4820 -2535 4825 -2505
rect 4825 -2535 4855 -2505
rect 4855 -2535 4860 -2505
rect 4820 -2540 4860 -2535
rect 4820 -2570 4860 -2565
rect 4820 -2600 4825 -2570
rect 4825 -2600 4855 -2570
rect 4855 -2600 4860 -2570
rect 4820 -2605 4860 -2600
rect 4820 -2640 4860 -2635
rect 4820 -2670 4825 -2640
rect 4825 -2670 4855 -2640
rect 4855 -2670 4860 -2640
rect 4820 -2675 4860 -2670
rect 4820 -2710 4860 -2705
rect 4820 -2740 4825 -2710
rect 4825 -2740 4855 -2710
rect 4855 -2740 4860 -2710
rect 4820 -2745 4860 -2740
rect 4820 -2780 4860 -2775
rect 4820 -2810 4825 -2780
rect 4825 -2810 4855 -2780
rect 4855 -2810 4860 -2780
rect 4820 -2815 4860 -2810
rect 4820 -2845 4860 -2840
rect 4820 -2875 4825 -2845
rect 4825 -2875 4855 -2845
rect 4855 -2875 4860 -2845
rect 4820 -2880 4860 -2875
rect 4820 -2905 4860 -2900
rect 4820 -2935 4825 -2905
rect 4825 -2935 4855 -2905
rect 4855 -2935 4860 -2905
rect 4820 -2940 4860 -2935
rect 4820 -2970 4860 -2965
rect 4820 -3000 4825 -2970
rect 4825 -3000 4855 -2970
rect 4855 -3000 4860 -2970
rect 4820 -3005 4860 -3000
rect 4820 -3040 4860 -3035
rect 4820 -3070 4825 -3040
rect 4825 -3070 4855 -3040
rect 4855 -3070 4860 -3040
rect 4820 -3075 4860 -3070
rect 4820 -3110 4860 -3105
rect 4820 -3140 4825 -3110
rect 4825 -3140 4855 -3110
rect 4855 -3140 4860 -3110
rect 4820 -3145 4860 -3140
rect 4820 -3180 4860 -3175
rect 4820 -3210 4825 -3180
rect 4825 -3210 4855 -3180
rect 4855 -3210 4860 -3180
rect 4820 -3215 4860 -3210
rect 4820 -3245 4860 -3240
rect 4820 -3275 4825 -3245
rect 4825 -3275 4855 -3245
rect 4855 -3275 4860 -3245
rect 4820 -3280 4860 -3275
rect 4820 -3305 4860 -3300
rect 4820 -3335 4825 -3305
rect 4825 -3335 4855 -3305
rect 4855 -3335 4860 -3305
rect 4820 -3340 4860 -3335
rect 4820 -3370 4860 -3365
rect 4820 -3400 4825 -3370
rect 4825 -3400 4855 -3370
rect 4855 -3400 4860 -3370
rect 4820 -3405 4860 -3400
rect 4820 -3440 4860 -3435
rect 4820 -3470 4825 -3440
rect 4825 -3470 4855 -3440
rect 4855 -3470 4860 -3440
rect 4820 -3475 4860 -3470
rect 4820 -3510 4860 -3505
rect 4820 -3540 4825 -3510
rect 4825 -3540 4855 -3510
rect 4855 -3540 4860 -3510
rect 4820 -3545 4860 -3540
rect 4820 -3580 4860 -3575
rect 4820 -3610 4825 -3580
rect 4825 -3610 4855 -3580
rect 4855 -3610 4860 -3580
rect 4820 -3615 4860 -3610
rect 4820 -3645 4860 -3640
rect 4820 -3675 4825 -3645
rect 4825 -3675 4855 -3645
rect 4855 -3675 4860 -3645
rect 4820 -3680 4860 -3675
rect 4820 -3705 4860 -3700
rect 4820 -3735 4825 -3705
rect 4825 -3735 4855 -3705
rect 4855 -3735 4860 -3705
rect 4820 -3740 4860 -3735
rect 4820 -3770 4860 -3765
rect 4820 -3800 4825 -3770
rect 4825 -3800 4855 -3770
rect 4855 -3800 4860 -3770
rect 4820 -3805 4860 -3800
rect 4820 -3840 4860 -3835
rect 4820 -3870 4825 -3840
rect 4825 -3870 4855 -3840
rect 4855 -3870 4860 -3840
rect 4820 -3875 4860 -3870
rect 4820 -3910 4860 -3905
rect 4820 -3940 4825 -3910
rect 4825 -3940 4855 -3910
rect 4855 -3940 4860 -3910
rect 4820 -3945 4860 -3940
rect 4820 -3980 4860 -3975
rect 4820 -4010 4825 -3980
rect 4825 -4010 4855 -3980
rect 4855 -4010 4860 -3980
rect 4820 -4015 4860 -4010
rect 4820 -4045 4860 -4040
rect 4820 -4075 4825 -4045
rect 4825 -4075 4855 -4045
rect 4855 -4075 4860 -4045
rect 4820 -4080 4860 -4075
rect 4820 -4105 4860 -4100
rect 4820 -4135 4825 -4105
rect 4825 -4135 4855 -4105
rect 4855 -4135 4860 -4105
rect 4820 -4140 4860 -4135
rect 4820 -4170 4860 -4165
rect 4820 -4200 4825 -4170
rect 4825 -4200 4855 -4170
rect 4855 -4200 4860 -4170
rect 4820 -4205 4860 -4200
rect 4820 -4240 4860 -4235
rect 4820 -4270 4825 -4240
rect 4825 -4270 4855 -4240
rect 4855 -4270 4860 -4240
rect 4820 -4275 4860 -4270
rect 4820 -4310 4860 -4305
rect 4820 -4340 4825 -4310
rect 4825 -4340 4855 -4310
rect 4855 -4340 4860 -4310
rect 4820 -4345 4860 -4340
rect 4820 -4380 4860 -4375
rect 4820 -4410 4825 -4380
rect 4825 -4410 4855 -4380
rect 4855 -4410 4860 -4380
rect 4820 -4415 4860 -4410
rect 4820 -4445 4860 -4440
rect 4820 -4475 4825 -4445
rect 4825 -4475 4855 -4445
rect 4855 -4475 4860 -4445
rect 4820 -4480 4860 -4475
rect 5170 -1305 5210 -1300
rect 5170 -1335 5175 -1305
rect 5175 -1335 5205 -1305
rect 5205 -1335 5210 -1305
rect 5170 -1340 5210 -1335
rect 5170 -1370 5210 -1365
rect 5170 -1400 5175 -1370
rect 5175 -1400 5205 -1370
rect 5205 -1400 5210 -1370
rect 5170 -1405 5210 -1400
rect 5170 -1440 5210 -1435
rect 5170 -1470 5175 -1440
rect 5175 -1470 5205 -1440
rect 5205 -1470 5210 -1440
rect 5170 -1475 5210 -1470
rect 5170 -1510 5210 -1505
rect 5170 -1540 5175 -1510
rect 5175 -1540 5205 -1510
rect 5205 -1540 5210 -1510
rect 5170 -1545 5210 -1540
rect 5170 -1580 5210 -1575
rect 5170 -1610 5175 -1580
rect 5175 -1610 5205 -1580
rect 5205 -1610 5210 -1580
rect 5170 -1615 5210 -1610
rect 5170 -1645 5210 -1640
rect 5170 -1675 5175 -1645
rect 5175 -1675 5205 -1645
rect 5205 -1675 5210 -1645
rect 5170 -1680 5210 -1675
rect 5170 -1705 5210 -1700
rect 5170 -1735 5175 -1705
rect 5175 -1735 5205 -1705
rect 5205 -1735 5210 -1705
rect 5170 -1740 5210 -1735
rect 5170 -1770 5210 -1765
rect 5170 -1800 5175 -1770
rect 5175 -1800 5205 -1770
rect 5205 -1800 5210 -1770
rect 5170 -1805 5210 -1800
rect 5170 -1840 5210 -1835
rect 5170 -1870 5175 -1840
rect 5175 -1870 5205 -1840
rect 5205 -1870 5210 -1840
rect 5170 -1875 5210 -1870
rect 5170 -1910 5210 -1905
rect 5170 -1940 5175 -1910
rect 5175 -1940 5205 -1910
rect 5205 -1940 5210 -1910
rect 5170 -1945 5210 -1940
rect 5170 -1980 5210 -1975
rect 5170 -2010 5175 -1980
rect 5175 -2010 5205 -1980
rect 5205 -2010 5210 -1980
rect 5170 -2015 5210 -2010
rect 5170 -2045 5210 -2040
rect 5170 -2075 5175 -2045
rect 5175 -2075 5205 -2045
rect 5205 -2075 5210 -2045
rect 5170 -2080 5210 -2075
rect 5170 -2105 5210 -2100
rect 5170 -2135 5175 -2105
rect 5175 -2135 5205 -2105
rect 5205 -2135 5210 -2105
rect 5170 -2140 5210 -2135
rect 5170 -2170 5210 -2165
rect 5170 -2200 5175 -2170
rect 5175 -2200 5205 -2170
rect 5205 -2200 5210 -2170
rect 5170 -2205 5210 -2200
rect 5170 -2240 5210 -2235
rect 5170 -2270 5175 -2240
rect 5175 -2270 5205 -2240
rect 5205 -2270 5210 -2240
rect 5170 -2275 5210 -2270
rect 5170 -2310 5210 -2305
rect 5170 -2340 5175 -2310
rect 5175 -2340 5205 -2310
rect 5205 -2340 5210 -2310
rect 5170 -2345 5210 -2340
rect 5170 -2380 5210 -2375
rect 5170 -2410 5175 -2380
rect 5175 -2410 5205 -2380
rect 5205 -2410 5210 -2380
rect 5170 -2415 5210 -2410
rect 5170 -2445 5210 -2440
rect 5170 -2475 5175 -2445
rect 5175 -2475 5205 -2445
rect 5205 -2475 5210 -2445
rect 5170 -2480 5210 -2475
rect 5170 -2505 5210 -2500
rect 5170 -2535 5175 -2505
rect 5175 -2535 5205 -2505
rect 5205 -2535 5210 -2505
rect 5170 -2540 5210 -2535
rect 5170 -2570 5210 -2565
rect 5170 -2600 5175 -2570
rect 5175 -2600 5205 -2570
rect 5205 -2600 5210 -2570
rect 5170 -2605 5210 -2600
rect 5170 -2640 5210 -2635
rect 5170 -2670 5175 -2640
rect 5175 -2670 5205 -2640
rect 5205 -2670 5210 -2640
rect 5170 -2675 5210 -2670
rect 5170 -2710 5210 -2705
rect 5170 -2740 5175 -2710
rect 5175 -2740 5205 -2710
rect 5205 -2740 5210 -2710
rect 5170 -2745 5210 -2740
rect 5170 -2780 5210 -2775
rect 5170 -2810 5175 -2780
rect 5175 -2810 5205 -2780
rect 5205 -2810 5210 -2780
rect 5170 -2815 5210 -2810
rect 5170 -2845 5210 -2840
rect 5170 -2875 5175 -2845
rect 5175 -2875 5205 -2845
rect 5205 -2875 5210 -2845
rect 5170 -2880 5210 -2875
rect 5170 -2905 5210 -2900
rect 5170 -2935 5175 -2905
rect 5175 -2935 5205 -2905
rect 5205 -2935 5210 -2905
rect 5170 -2940 5210 -2935
rect 5170 -2970 5210 -2965
rect 5170 -3000 5175 -2970
rect 5175 -3000 5205 -2970
rect 5205 -3000 5210 -2970
rect 5170 -3005 5210 -3000
rect 5170 -3040 5210 -3035
rect 5170 -3070 5175 -3040
rect 5175 -3070 5205 -3040
rect 5205 -3070 5210 -3040
rect 5170 -3075 5210 -3070
rect 5170 -3110 5210 -3105
rect 5170 -3140 5175 -3110
rect 5175 -3140 5205 -3110
rect 5205 -3140 5210 -3110
rect 5170 -3145 5210 -3140
rect 5170 -3180 5210 -3175
rect 5170 -3210 5175 -3180
rect 5175 -3210 5205 -3180
rect 5205 -3210 5210 -3180
rect 5170 -3215 5210 -3210
rect 5170 -3245 5210 -3240
rect 5170 -3275 5175 -3245
rect 5175 -3275 5205 -3245
rect 5205 -3275 5210 -3245
rect 5170 -3280 5210 -3275
rect 5170 -3305 5210 -3300
rect 5170 -3335 5175 -3305
rect 5175 -3335 5205 -3305
rect 5205 -3335 5210 -3305
rect 5170 -3340 5210 -3335
rect 5170 -3370 5210 -3365
rect 5170 -3400 5175 -3370
rect 5175 -3400 5205 -3370
rect 5205 -3400 5210 -3370
rect 5170 -3405 5210 -3400
rect 5170 -3440 5210 -3435
rect 5170 -3470 5175 -3440
rect 5175 -3470 5205 -3440
rect 5205 -3470 5210 -3440
rect 5170 -3475 5210 -3470
rect 5170 -3510 5210 -3505
rect 5170 -3540 5175 -3510
rect 5175 -3540 5205 -3510
rect 5205 -3540 5210 -3510
rect 5170 -3545 5210 -3540
rect 5170 -3580 5210 -3575
rect 5170 -3610 5175 -3580
rect 5175 -3610 5205 -3580
rect 5205 -3610 5210 -3580
rect 5170 -3615 5210 -3610
rect 5170 -3645 5210 -3640
rect 5170 -3675 5175 -3645
rect 5175 -3675 5205 -3645
rect 5205 -3675 5210 -3645
rect 5170 -3680 5210 -3675
rect 5170 -3705 5210 -3700
rect 5170 -3735 5175 -3705
rect 5175 -3735 5205 -3705
rect 5205 -3735 5210 -3705
rect 5170 -3740 5210 -3735
rect 5170 -3770 5210 -3765
rect 5170 -3800 5175 -3770
rect 5175 -3800 5205 -3770
rect 5205 -3800 5210 -3770
rect 5170 -3805 5210 -3800
rect 5170 -3840 5210 -3835
rect 5170 -3870 5175 -3840
rect 5175 -3870 5205 -3840
rect 5205 -3870 5210 -3840
rect 5170 -3875 5210 -3870
rect 5170 -3910 5210 -3905
rect 5170 -3940 5175 -3910
rect 5175 -3940 5205 -3910
rect 5205 -3940 5210 -3910
rect 5170 -3945 5210 -3940
rect 5170 -3980 5210 -3975
rect 5170 -4010 5175 -3980
rect 5175 -4010 5205 -3980
rect 5205 -4010 5210 -3980
rect 5170 -4015 5210 -4010
rect 5170 -4045 5210 -4040
rect 5170 -4075 5175 -4045
rect 5175 -4075 5205 -4045
rect 5205 -4075 5210 -4045
rect 5170 -4080 5210 -4075
rect 5170 -4105 5210 -4100
rect 5170 -4135 5175 -4105
rect 5175 -4135 5205 -4105
rect 5205 -4135 5210 -4105
rect 5170 -4140 5210 -4135
rect 5170 -4170 5210 -4165
rect 5170 -4200 5175 -4170
rect 5175 -4200 5205 -4170
rect 5205 -4200 5210 -4170
rect 5170 -4205 5210 -4200
rect 5170 -4240 5210 -4235
rect 5170 -4270 5175 -4240
rect 5175 -4270 5205 -4240
rect 5205 -4270 5210 -4240
rect 5170 -4275 5210 -4270
rect 5170 -4310 5210 -4305
rect 5170 -4340 5175 -4310
rect 5175 -4340 5205 -4310
rect 5205 -4340 5210 -4310
rect 5170 -4345 5210 -4340
rect 5170 -4380 5210 -4375
rect 5170 -4410 5175 -4380
rect 5175 -4410 5205 -4380
rect 5205 -4410 5210 -4380
rect 5170 -4415 5210 -4410
rect 5170 -4445 5210 -4440
rect 5170 -4475 5175 -4445
rect 5175 -4475 5205 -4445
rect 5205 -4475 5210 -4445
rect 5170 -4480 5210 -4475
rect 5520 -1305 5560 -1300
rect 5520 -1335 5525 -1305
rect 5525 -1335 5555 -1305
rect 5555 -1335 5560 -1305
rect 5520 -1340 5560 -1335
rect 5520 -1370 5560 -1365
rect 5520 -1400 5525 -1370
rect 5525 -1400 5555 -1370
rect 5555 -1400 5560 -1370
rect 5520 -1405 5560 -1400
rect 5520 -1440 5560 -1435
rect 5520 -1470 5525 -1440
rect 5525 -1470 5555 -1440
rect 5555 -1470 5560 -1440
rect 5520 -1475 5560 -1470
rect 5520 -1510 5560 -1505
rect 5520 -1540 5525 -1510
rect 5525 -1540 5555 -1510
rect 5555 -1540 5560 -1510
rect 5520 -1545 5560 -1540
rect 5520 -1580 5560 -1575
rect 5520 -1610 5525 -1580
rect 5525 -1610 5555 -1580
rect 5555 -1610 5560 -1580
rect 5520 -1615 5560 -1610
rect 5520 -1645 5560 -1640
rect 5520 -1675 5525 -1645
rect 5525 -1675 5555 -1645
rect 5555 -1675 5560 -1645
rect 5520 -1680 5560 -1675
rect 5520 -1705 5560 -1700
rect 5520 -1735 5525 -1705
rect 5525 -1735 5555 -1705
rect 5555 -1735 5560 -1705
rect 5520 -1740 5560 -1735
rect 5520 -1770 5560 -1765
rect 5520 -1800 5525 -1770
rect 5525 -1800 5555 -1770
rect 5555 -1800 5560 -1770
rect 5520 -1805 5560 -1800
rect 5520 -1840 5560 -1835
rect 5520 -1870 5525 -1840
rect 5525 -1870 5555 -1840
rect 5555 -1870 5560 -1840
rect 5520 -1875 5560 -1870
rect 5520 -1910 5560 -1905
rect 5520 -1940 5525 -1910
rect 5525 -1940 5555 -1910
rect 5555 -1940 5560 -1910
rect 5520 -1945 5560 -1940
rect 5520 -1980 5560 -1975
rect 5520 -2010 5525 -1980
rect 5525 -2010 5555 -1980
rect 5555 -2010 5560 -1980
rect 5520 -2015 5560 -2010
rect 5520 -2045 5560 -2040
rect 5520 -2075 5525 -2045
rect 5525 -2075 5555 -2045
rect 5555 -2075 5560 -2045
rect 5520 -2080 5560 -2075
rect 5520 -2105 5560 -2100
rect 5520 -2135 5525 -2105
rect 5525 -2135 5555 -2105
rect 5555 -2135 5560 -2105
rect 5520 -2140 5560 -2135
rect 5520 -2170 5560 -2165
rect 5520 -2200 5525 -2170
rect 5525 -2200 5555 -2170
rect 5555 -2200 5560 -2170
rect 5520 -2205 5560 -2200
rect 5520 -2240 5560 -2235
rect 5520 -2270 5525 -2240
rect 5525 -2270 5555 -2240
rect 5555 -2270 5560 -2240
rect 5520 -2275 5560 -2270
rect 5520 -2310 5560 -2305
rect 5520 -2340 5525 -2310
rect 5525 -2340 5555 -2310
rect 5555 -2340 5560 -2310
rect 5520 -2345 5560 -2340
rect 5520 -2380 5560 -2375
rect 5520 -2410 5525 -2380
rect 5525 -2410 5555 -2380
rect 5555 -2410 5560 -2380
rect 5520 -2415 5560 -2410
rect 5520 -2445 5560 -2440
rect 5520 -2475 5525 -2445
rect 5525 -2475 5555 -2445
rect 5555 -2475 5560 -2445
rect 5520 -2480 5560 -2475
rect 5520 -2505 5560 -2500
rect 5520 -2535 5525 -2505
rect 5525 -2535 5555 -2505
rect 5555 -2535 5560 -2505
rect 5520 -2540 5560 -2535
rect 5520 -2570 5560 -2565
rect 5520 -2600 5525 -2570
rect 5525 -2600 5555 -2570
rect 5555 -2600 5560 -2570
rect 5520 -2605 5560 -2600
rect 5520 -2640 5560 -2635
rect 5520 -2670 5525 -2640
rect 5525 -2670 5555 -2640
rect 5555 -2670 5560 -2640
rect 5520 -2675 5560 -2670
rect 5520 -2710 5560 -2705
rect 5520 -2740 5525 -2710
rect 5525 -2740 5555 -2710
rect 5555 -2740 5560 -2710
rect 5520 -2745 5560 -2740
rect 5520 -2780 5560 -2775
rect 5520 -2810 5525 -2780
rect 5525 -2810 5555 -2780
rect 5555 -2810 5560 -2780
rect 5520 -2815 5560 -2810
rect 5520 -2845 5560 -2840
rect 5520 -2875 5525 -2845
rect 5525 -2875 5555 -2845
rect 5555 -2875 5560 -2845
rect 5520 -2880 5560 -2875
rect 5520 -2905 5560 -2900
rect 5520 -2935 5525 -2905
rect 5525 -2935 5555 -2905
rect 5555 -2935 5560 -2905
rect 5520 -2940 5560 -2935
rect 5520 -2970 5560 -2965
rect 5520 -3000 5525 -2970
rect 5525 -3000 5555 -2970
rect 5555 -3000 5560 -2970
rect 5520 -3005 5560 -3000
rect 5520 -3040 5560 -3035
rect 5520 -3070 5525 -3040
rect 5525 -3070 5555 -3040
rect 5555 -3070 5560 -3040
rect 5520 -3075 5560 -3070
rect 5520 -3110 5560 -3105
rect 5520 -3140 5525 -3110
rect 5525 -3140 5555 -3110
rect 5555 -3140 5560 -3110
rect 5520 -3145 5560 -3140
rect 5520 -3180 5560 -3175
rect 5520 -3210 5525 -3180
rect 5525 -3210 5555 -3180
rect 5555 -3210 5560 -3180
rect 5520 -3215 5560 -3210
rect 5520 -3245 5560 -3240
rect 5520 -3275 5525 -3245
rect 5525 -3275 5555 -3245
rect 5555 -3275 5560 -3245
rect 5520 -3280 5560 -3275
rect 5520 -3305 5560 -3300
rect 5520 -3335 5525 -3305
rect 5525 -3335 5555 -3305
rect 5555 -3335 5560 -3305
rect 5520 -3340 5560 -3335
rect 5520 -3370 5560 -3365
rect 5520 -3400 5525 -3370
rect 5525 -3400 5555 -3370
rect 5555 -3400 5560 -3370
rect 5520 -3405 5560 -3400
rect 5520 -3440 5560 -3435
rect 5520 -3470 5525 -3440
rect 5525 -3470 5555 -3440
rect 5555 -3470 5560 -3440
rect 5520 -3475 5560 -3470
rect 5520 -3510 5560 -3505
rect 5520 -3540 5525 -3510
rect 5525 -3540 5555 -3510
rect 5555 -3540 5560 -3510
rect 5520 -3545 5560 -3540
rect 5520 -3580 5560 -3575
rect 5520 -3610 5525 -3580
rect 5525 -3610 5555 -3580
rect 5555 -3610 5560 -3580
rect 5520 -3615 5560 -3610
rect 5520 -3645 5560 -3640
rect 5520 -3675 5525 -3645
rect 5525 -3675 5555 -3645
rect 5555 -3675 5560 -3645
rect 5520 -3680 5560 -3675
rect 5520 -3705 5560 -3700
rect 5520 -3735 5525 -3705
rect 5525 -3735 5555 -3705
rect 5555 -3735 5560 -3705
rect 5520 -3740 5560 -3735
rect 5520 -3770 5560 -3765
rect 5520 -3800 5525 -3770
rect 5525 -3800 5555 -3770
rect 5555 -3800 5560 -3770
rect 5520 -3805 5560 -3800
rect 5520 -3840 5560 -3835
rect 5520 -3870 5525 -3840
rect 5525 -3870 5555 -3840
rect 5555 -3870 5560 -3840
rect 5520 -3875 5560 -3870
rect 5520 -3910 5560 -3905
rect 5520 -3940 5525 -3910
rect 5525 -3940 5555 -3910
rect 5555 -3940 5560 -3910
rect 5520 -3945 5560 -3940
rect 5520 -3980 5560 -3975
rect 5520 -4010 5525 -3980
rect 5525 -4010 5555 -3980
rect 5555 -4010 5560 -3980
rect 5520 -4015 5560 -4010
rect 5520 -4045 5560 -4040
rect 5520 -4075 5525 -4045
rect 5525 -4075 5555 -4045
rect 5555 -4075 5560 -4045
rect 5520 -4080 5560 -4075
rect 5520 -4105 5560 -4100
rect 5520 -4135 5525 -4105
rect 5525 -4135 5555 -4105
rect 5555 -4135 5560 -4105
rect 5520 -4140 5560 -4135
rect 5520 -4170 5560 -4165
rect 5520 -4200 5525 -4170
rect 5525 -4200 5555 -4170
rect 5555 -4200 5560 -4170
rect 5520 -4205 5560 -4200
rect 5520 -4240 5560 -4235
rect 5520 -4270 5525 -4240
rect 5525 -4270 5555 -4240
rect 5555 -4270 5560 -4240
rect 5520 -4275 5560 -4270
rect 5520 -4310 5560 -4305
rect 5520 -4340 5525 -4310
rect 5525 -4340 5555 -4310
rect 5555 -4340 5560 -4310
rect 5520 -4345 5560 -4340
rect 5520 -4380 5560 -4375
rect 5520 -4410 5525 -4380
rect 5525 -4410 5555 -4380
rect 5555 -4410 5560 -4380
rect 5520 -4415 5560 -4410
rect 5520 -4445 5560 -4440
rect 5520 -4475 5525 -4445
rect 5525 -4475 5555 -4445
rect 5555 -4475 5560 -4445
rect 5520 -4480 5560 -4475
rect 5870 -1305 5910 -1300
rect 5870 -1335 5875 -1305
rect 5875 -1335 5905 -1305
rect 5905 -1335 5910 -1305
rect 5870 -1340 5910 -1335
rect 5870 -1370 5910 -1365
rect 5870 -1400 5875 -1370
rect 5875 -1400 5905 -1370
rect 5905 -1400 5910 -1370
rect 5870 -1405 5910 -1400
rect 5870 -1440 5910 -1435
rect 5870 -1470 5875 -1440
rect 5875 -1470 5905 -1440
rect 5905 -1470 5910 -1440
rect 5870 -1475 5910 -1470
rect 5870 -1510 5910 -1505
rect 5870 -1540 5875 -1510
rect 5875 -1540 5905 -1510
rect 5905 -1540 5910 -1510
rect 5870 -1545 5910 -1540
rect 5870 -1580 5910 -1575
rect 5870 -1610 5875 -1580
rect 5875 -1610 5905 -1580
rect 5905 -1610 5910 -1580
rect 5870 -1615 5910 -1610
rect 5870 -1645 5910 -1640
rect 5870 -1675 5875 -1645
rect 5875 -1675 5905 -1645
rect 5905 -1675 5910 -1645
rect 5870 -1680 5910 -1675
rect 5870 -1705 5910 -1700
rect 5870 -1735 5875 -1705
rect 5875 -1735 5905 -1705
rect 5905 -1735 5910 -1705
rect 5870 -1740 5910 -1735
rect 5870 -1770 5910 -1765
rect 5870 -1800 5875 -1770
rect 5875 -1800 5905 -1770
rect 5905 -1800 5910 -1770
rect 5870 -1805 5910 -1800
rect 5870 -1840 5910 -1835
rect 5870 -1870 5875 -1840
rect 5875 -1870 5905 -1840
rect 5905 -1870 5910 -1840
rect 5870 -1875 5910 -1870
rect 5870 -1910 5910 -1905
rect 5870 -1940 5875 -1910
rect 5875 -1940 5905 -1910
rect 5905 -1940 5910 -1910
rect 5870 -1945 5910 -1940
rect 5870 -1980 5910 -1975
rect 5870 -2010 5875 -1980
rect 5875 -2010 5905 -1980
rect 5905 -2010 5910 -1980
rect 5870 -2015 5910 -2010
rect 5870 -2045 5910 -2040
rect 5870 -2075 5875 -2045
rect 5875 -2075 5905 -2045
rect 5905 -2075 5910 -2045
rect 5870 -2080 5910 -2075
rect 5870 -2105 5910 -2100
rect 5870 -2135 5875 -2105
rect 5875 -2135 5905 -2105
rect 5905 -2135 5910 -2105
rect 5870 -2140 5910 -2135
rect 5870 -2170 5910 -2165
rect 5870 -2200 5875 -2170
rect 5875 -2200 5905 -2170
rect 5905 -2200 5910 -2170
rect 5870 -2205 5910 -2200
rect 5870 -2240 5910 -2235
rect 5870 -2270 5875 -2240
rect 5875 -2270 5905 -2240
rect 5905 -2270 5910 -2240
rect 5870 -2275 5910 -2270
rect 5870 -2310 5910 -2305
rect 5870 -2340 5875 -2310
rect 5875 -2340 5905 -2310
rect 5905 -2340 5910 -2310
rect 5870 -2345 5910 -2340
rect 5870 -2380 5910 -2375
rect 5870 -2410 5875 -2380
rect 5875 -2410 5905 -2380
rect 5905 -2410 5910 -2380
rect 5870 -2415 5910 -2410
rect 5870 -2445 5910 -2440
rect 5870 -2475 5875 -2445
rect 5875 -2475 5905 -2445
rect 5905 -2475 5910 -2445
rect 5870 -2480 5910 -2475
rect 5870 -2505 5910 -2500
rect 5870 -2535 5875 -2505
rect 5875 -2535 5905 -2505
rect 5905 -2535 5910 -2505
rect 5870 -2540 5910 -2535
rect 5870 -2570 5910 -2565
rect 5870 -2600 5875 -2570
rect 5875 -2600 5905 -2570
rect 5905 -2600 5910 -2570
rect 5870 -2605 5910 -2600
rect 5870 -2640 5910 -2635
rect 5870 -2670 5875 -2640
rect 5875 -2670 5905 -2640
rect 5905 -2670 5910 -2640
rect 5870 -2675 5910 -2670
rect 5870 -2710 5910 -2705
rect 5870 -2740 5875 -2710
rect 5875 -2740 5905 -2710
rect 5905 -2740 5910 -2710
rect 5870 -2745 5910 -2740
rect 5870 -2780 5910 -2775
rect 5870 -2810 5875 -2780
rect 5875 -2810 5905 -2780
rect 5905 -2810 5910 -2780
rect 5870 -2815 5910 -2810
rect 5870 -2845 5910 -2840
rect 5870 -2875 5875 -2845
rect 5875 -2875 5905 -2845
rect 5905 -2875 5910 -2845
rect 5870 -2880 5910 -2875
rect 5870 -2905 5910 -2900
rect 5870 -2935 5875 -2905
rect 5875 -2935 5905 -2905
rect 5905 -2935 5910 -2905
rect 5870 -2940 5910 -2935
rect 5870 -2970 5910 -2965
rect 5870 -3000 5875 -2970
rect 5875 -3000 5905 -2970
rect 5905 -3000 5910 -2970
rect 5870 -3005 5910 -3000
rect 5870 -3040 5910 -3035
rect 5870 -3070 5875 -3040
rect 5875 -3070 5905 -3040
rect 5905 -3070 5910 -3040
rect 5870 -3075 5910 -3070
rect 5870 -3110 5910 -3105
rect 5870 -3140 5875 -3110
rect 5875 -3140 5905 -3110
rect 5905 -3140 5910 -3110
rect 5870 -3145 5910 -3140
rect 5870 -3180 5910 -3175
rect 5870 -3210 5875 -3180
rect 5875 -3210 5905 -3180
rect 5905 -3210 5910 -3180
rect 5870 -3215 5910 -3210
rect 5870 -3245 5910 -3240
rect 5870 -3275 5875 -3245
rect 5875 -3275 5905 -3245
rect 5905 -3275 5910 -3245
rect 5870 -3280 5910 -3275
rect 5870 -3305 5910 -3300
rect 5870 -3335 5875 -3305
rect 5875 -3335 5905 -3305
rect 5905 -3335 5910 -3305
rect 5870 -3340 5910 -3335
rect 5870 -3370 5910 -3365
rect 5870 -3400 5875 -3370
rect 5875 -3400 5905 -3370
rect 5905 -3400 5910 -3370
rect 5870 -3405 5910 -3400
rect 5870 -3440 5910 -3435
rect 5870 -3470 5875 -3440
rect 5875 -3470 5905 -3440
rect 5905 -3470 5910 -3440
rect 5870 -3475 5910 -3470
rect 5870 -3510 5910 -3505
rect 5870 -3540 5875 -3510
rect 5875 -3540 5905 -3510
rect 5905 -3540 5910 -3510
rect 5870 -3545 5910 -3540
rect 5870 -3580 5910 -3575
rect 5870 -3610 5875 -3580
rect 5875 -3610 5905 -3580
rect 5905 -3610 5910 -3580
rect 5870 -3615 5910 -3610
rect 5870 -3645 5910 -3640
rect 5870 -3675 5875 -3645
rect 5875 -3675 5905 -3645
rect 5905 -3675 5910 -3645
rect 5870 -3680 5910 -3675
rect 5870 -3705 5910 -3700
rect 5870 -3735 5875 -3705
rect 5875 -3735 5905 -3705
rect 5905 -3735 5910 -3705
rect 5870 -3740 5910 -3735
rect 5870 -3770 5910 -3765
rect 5870 -3800 5875 -3770
rect 5875 -3800 5905 -3770
rect 5905 -3800 5910 -3770
rect 5870 -3805 5910 -3800
rect 5870 -3840 5910 -3835
rect 5870 -3870 5875 -3840
rect 5875 -3870 5905 -3840
rect 5905 -3870 5910 -3840
rect 5870 -3875 5910 -3870
rect 5870 -3910 5910 -3905
rect 5870 -3940 5875 -3910
rect 5875 -3940 5905 -3910
rect 5905 -3940 5910 -3910
rect 5870 -3945 5910 -3940
rect 5870 -3980 5910 -3975
rect 5870 -4010 5875 -3980
rect 5875 -4010 5905 -3980
rect 5905 -4010 5910 -3980
rect 5870 -4015 5910 -4010
rect 5870 -4045 5910 -4040
rect 5870 -4075 5875 -4045
rect 5875 -4075 5905 -4045
rect 5905 -4075 5910 -4045
rect 5870 -4080 5910 -4075
rect 5870 -4105 5910 -4100
rect 5870 -4135 5875 -4105
rect 5875 -4135 5905 -4105
rect 5905 -4135 5910 -4105
rect 5870 -4140 5910 -4135
rect 5870 -4170 5910 -4165
rect 5870 -4200 5875 -4170
rect 5875 -4200 5905 -4170
rect 5905 -4200 5910 -4170
rect 5870 -4205 5910 -4200
rect 5870 -4240 5910 -4235
rect 5870 -4270 5875 -4240
rect 5875 -4270 5905 -4240
rect 5905 -4270 5910 -4240
rect 5870 -4275 5910 -4270
rect 5870 -4310 5910 -4305
rect 5870 -4340 5875 -4310
rect 5875 -4340 5905 -4310
rect 5905 -4340 5910 -4310
rect 5870 -4345 5910 -4340
rect 5870 -4380 5910 -4375
rect 5870 -4410 5875 -4380
rect 5875 -4410 5905 -4380
rect 5905 -4410 5910 -4380
rect 5870 -4415 5910 -4410
rect 5870 -4445 5910 -4440
rect 5870 -4475 5875 -4445
rect 5875 -4475 5905 -4445
rect 5905 -4475 5910 -4445
rect 5870 -4480 5910 -4475
rect 6220 -1305 6260 -1300
rect 6220 -1335 6225 -1305
rect 6225 -1335 6255 -1305
rect 6255 -1335 6260 -1305
rect 6220 -1340 6260 -1335
rect 6220 -1370 6260 -1365
rect 6220 -1400 6225 -1370
rect 6225 -1400 6255 -1370
rect 6255 -1400 6260 -1370
rect 6220 -1405 6260 -1400
rect 6220 -1440 6260 -1435
rect 6220 -1470 6225 -1440
rect 6225 -1470 6255 -1440
rect 6255 -1470 6260 -1440
rect 6220 -1475 6260 -1470
rect 6220 -1510 6260 -1505
rect 6220 -1540 6225 -1510
rect 6225 -1540 6255 -1510
rect 6255 -1540 6260 -1510
rect 6220 -1545 6260 -1540
rect 6220 -1580 6260 -1575
rect 6220 -1610 6225 -1580
rect 6225 -1610 6255 -1580
rect 6255 -1610 6260 -1580
rect 6220 -1615 6260 -1610
rect 6220 -1645 6260 -1640
rect 6220 -1675 6225 -1645
rect 6225 -1675 6255 -1645
rect 6255 -1675 6260 -1645
rect 6220 -1680 6260 -1675
rect 6220 -1705 6260 -1700
rect 6220 -1735 6225 -1705
rect 6225 -1735 6255 -1705
rect 6255 -1735 6260 -1705
rect 6220 -1740 6260 -1735
rect 6220 -1770 6260 -1765
rect 6220 -1800 6225 -1770
rect 6225 -1800 6255 -1770
rect 6255 -1800 6260 -1770
rect 6220 -1805 6260 -1800
rect 6220 -1840 6260 -1835
rect 6220 -1870 6225 -1840
rect 6225 -1870 6255 -1840
rect 6255 -1870 6260 -1840
rect 6220 -1875 6260 -1870
rect 6220 -1910 6260 -1905
rect 6220 -1940 6225 -1910
rect 6225 -1940 6255 -1910
rect 6255 -1940 6260 -1910
rect 6220 -1945 6260 -1940
rect 6220 -1980 6260 -1975
rect 6220 -2010 6225 -1980
rect 6225 -2010 6255 -1980
rect 6255 -2010 6260 -1980
rect 6220 -2015 6260 -2010
rect 6220 -2045 6260 -2040
rect 6220 -2075 6225 -2045
rect 6225 -2075 6255 -2045
rect 6255 -2075 6260 -2045
rect 6220 -2080 6260 -2075
rect 6220 -2105 6260 -2100
rect 6220 -2135 6225 -2105
rect 6225 -2135 6255 -2105
rect 6255 -2135 6260 -2105
rect 6220 -2140 6260 -2135
rect 6220 -2170 6260 -2165
rect 6220 -2200 6225 -2170
rect 6225 -2200 6255 -2170
rect 6255 -2200 6260 -2170
rect 6220 -2205 6260 -2200
rect 6220 -2240 6260 -2235
rect 6220 -2270 6225 -2240
rect 6225 -2270 6255 -2240
rect 6255 -2270 6260 -2240
rect 6220 -2275 6260 -2270
rect 6220 -2310 6260 -2305
rect 6220 -2340 6225 -2310
rect 6225 -2340 6255 -2310
rect 6255 -2340 6260 -2310
rect 6220 -2345 6260 -2340
rect 6220 -2380 6260 -2375
rect 6220 -2410 6225 -2380
rect 6225 -2410 6255 -2380
rect 6255 -2410 6260 -2380
rect 6220 -2415 6260 -2410
rect 6220 -2445 6260 -2440
rect 6220 -2475 6225 -2445
rect 6225 -2475 6255 -2445
rect 6255 -2475 6260 -2445
rect 6220 -2480 6260 -2475
rect 6220 -2505 6260 -2500
rect 6220 -2535 6225 -2505
rect 6225 -2535 6255 -2505
rect 6255 -2535 6260 -2505
rect 6220 -2540 6260 -2535
rect 6220 -2570 6260 -2565
rect 6220 -2600 6225 -2570
rect 6225 -2600 6255 -2570
rect 6255 -2600 6260 -2570
rect 6220 -2605 6260 -2600
rect 6220 -2640 6260 -2635
rect 6220 -2670 6225 -2640
rect 6225 -2670 6255 -2640
rect 6255 -2670 6260 -2640
rect 6220 -2675 6260 -2670
rect 6220 -2710 6260 -2705
rect 6220 -2740 6225 -2710
rect 6225 -2740 6255 -2710
rect 6255 -2740 6260 -2710
rect 6220 -2745 6260 -2740
rect 6220 -2780 6260 -2775
rect 6220 -2810 6225 -2780
rect 6225 -2810 6255 -2780
rect 6255 -2810 6260 -2780
rect 6220 -2815 6260 -2810
rect 6220 -2845 6260 -2840
rect 6220 -2875 6225 -2845
rect 6225 -2875 6255 -2845
rect 6255 -2875 6260 -2845
rect 6220 -2880 6260 -2875
rect 6220 -2905 6260 -2900
rect 6220 -2935 6225 -2905
rect 6225 -2935 6255 -2905
rect 6255 -2935 6260 -2905
rect 6220 -2940 6260 -2935
rect 6220 -2970 6260 -2965
rect 6220 -3000 6225 -2970
rect 6225 -3000 6255 -2970
rect 6255 -3000 6260 -2970
rect 6220 -3005 6260 -3000
rect 6220 -3040 6260 -3035
rect 6220 -3070 6225 -3040
rect 6225 -3070 6255 -3040
rect 6255 -3070 6260 -3040
rect 6220 -3075 6260 -3070
rect 6220 -3110 6260 -3105
rect 6220 -3140 6225 -3110
rect 6225 -3140 6255 -3110
rect 6255 -3140 6260 -3110
rect 6220 -3145 6260 -3140
rect 6220 -3180 6260 -3175
rect 6220 -3210 6225 -3180
rect 6225 -3210 6255 -3180
rect 6255 -3210 6260 -3180
rect 6220 -3215 6260 -3210
rect 6220 -3245 6260 -3240
rect 6220 -3275 6225 -3245
rect 6225 -3275 6255 -3245
rect 6255 -3275 6260 -3245
rect 6220 -3280 6260 -3275
rect 6220 -3305 6260 -3300
rect 6220 -3335 6225 -3305
rect 6225 -3335 6255 -3305
rect 6255 -3335 6260 -3305
rect 6220 -3340 6260 -3335
rect 6220 -3370 6260 -3365
rect 6220 -3400 6225 -3370
rect 6225 -3400 6255 -3370
rect 6255 -3400 6260 -3370
rect 6220 -3405 6260 -3400
rect 6220 -3440 6260 -3435
rect 6220 -3470 6225 -3440
rect 6225 -3470 6255 -3440
rect 6255 -3470 6260 -3440
rect 6220 -3475 6260 -3470
rect 6220 -3510 6260 -3505
rect 6220 -3540 6225 -3510
rect 6225 -3540 6255 -3510
rect 6255 -3540 6260 -3510
rect 6220 -3545 6260 -3540
rect 6220 -3580 6260 -3575
rect 6220 -3610 6225 -3580
rect 6225 -3610 6255 -3580
rect 6255 -3610 6260 -3580
rect 6220 -3615 6260 -3610
rect 6220 -3645 6260 -3640
rect 6220 -3675 6225 -3645
rect 6225 -3675 6255 -3645
rect 6255 -3675 6260 -3645
rect 6220 -3680 6260 -3675
rect 6220 -3705 6260 -3700
rect 6220 -3735 6225 -3705
rect 6225 -3735 6255 -3705
rect 6255 -3735 6260 -3705
rect 6220 -3740 6260 -3735
rect 6220 -3770 6260 -3765
rect 6220 -3800 6225 -3770
rect 6225 -3800 6255 -3770
rect 6255 -3800 6260 -3770
rect 6220 -3805 6260 -3800
rect 6220 -3840 6260 -3835
rect 6220 -3870 6225 -3840
rect 6225 -3870 6255 -3840
rect 6255 -3870 6260 -3840
rect 6220 -3875 6260 -3870
rect 6220 -3910 6260 -3905
rect 6220 -3940 6225 -3910
rect 6225 -3940 6255 -3910
rect 6255 -3940 6260 -3910
rect 6220 -3945 6260 -3940
rect 6220 -3980 6260 -3975
rect 6220 -4010 6225 -3980
rect 6225 -4010 6255 -3980
rect 6255 -4010 6260 -3980
rect 6220 -4015 6260 -4010
rect 6220 -4045 6260 -4040
rect 6220 -4075 6225 -4045
rect 6225 -4075 6255 -4045
rect 6255 -4075 6260 -4045
rect 6220 -4080 6260 -4075
rect 6220 -4105 6260 -4100
rect 6220 -4135 6225 -4105
rect 6225 -4135 6255 -4105
rect 6255 -4135 6260 -4105
rect 6220 -4140 6260 -4135
rect 6220 -4170 6260 -4165
rect 6220 -4200 6225 -4170
rect 6225 -4200 6255 -4170
rect 6255 -4200 6260 -4170
rect 6220 -4205 6260 -4200
rect 6220 -4240 6260 -4235
rect 6220 -4270 6225 -4240
rect 6225 -4270 6255 -4240
rect 6255 -4270 6260 -4240
rect 6220 -4275 6260 -4270
rect 6220 -4310 6260 -4305
rect 6220 -4340 6225 -4310
rect 6225 -4340 6255 -4310
rect 6255 -4340 6260 -4310
rect 6220 -4345 6260 -4340
rect 6220 -4380 6260 -4375
rect 6220 -4410 6225 -4380
rect 6225 -4410 6255 -4380
rect 6255 -4410 6260 -4380
rect 6220 -4415 6260 -4410
rect 6220 -4445 6260 -4440
rect 6220 -4475 6225 -4445
rect 6225 -4475 6255 -4445
rect 6255 -4475 6260 -4445
rect 6220 -4480 6260 -4475
rect 6570 -1305 6610 -1300
rect 6570 -1335 6575 -1305
rect 6575 -1335 6605 -1305
rect 6605 -1335 6610 -1305
rect 6570 -1340 6610 -1335
rect 6570 -1370 6610 -1365
rect 6570 -1400 6575 -1370
rect 6575 -1400 6605 -1370
rect 6605 -1400 6610 -1370
rect 6570 -1405 6610 -1400
rect 6570 -1440 6610 -1435
rect 6570 -1470 6575 -1440
rect 6575 -1470 6605 -1440
rect 6605 -1470 6610 -1440
rect 6570 -1475 6610 -1470
rect 6570 -1510 6610 -1505
rect 6570 -1540 6575 -1510
rect 6575 -1540 6605 -1510
rect 6605 -1540 6610 -1510
rect 6570 -1545 6610 -1540
rect 6570 -1580 6610 -1575
rect 6570 -1610 6575 -1580
rect 6575 -1610 6605 -1580
rect 6605 -1610 6610 -1580
rect 6570 -1615 6610 -1610
rect 6570 -1645 6610 -1640
rect 6570 -1675 6575 -1645
rect 6575 -1675 6605 -1645
rect 6605 -1675 6610 -1645
rect 6570 -1680 6610 -1675
rect 6570 -1705 6610 -1700
rect 6570 -1735 6575 -1705
rect 6575 -1735 6605 -1705
rect 6605 -1735 6610 -1705
rect 6570 -1740 6610 -1735
rect 6570 -1770 6610 -1765
rect 6570 -1800 6575 -1770
rect 6575 -1800 6605 -1770
rect 6605 -1800 6610 -1770
rect 6570 -1805 6610 -1800
rect 6570 -1840 6610 -1835
rect 6570 -1870 6575 -1840
rect 6575 -1870 6605 -1840
rect 6605 -1870 6610 -1840
rect 6570 -1875 6610 -1870
rect 6570 -1910 6610 -1905
rect 6570 -1940 6575 -1910
rect 6575 -1940 6605 -1910
rect 6605 -1940 6610 -1910
rect 6570 -1945 6610 -1940
rect 6570 -1980 6610 -1975
rect 6570 -2010 6575 -1980
rect 6575 -2010 6605 -1980
rect 6605 -2010 6610 -1980
rect 6570 -2015 6610 -2010
rect 6570 -2045 6610 -2040
rect 6570 -2075 6575 -2045
rect 6575 -2075 6605 -2045
rect 6605 -2075 6610 -2045
rect 6570 -2080 6610 -2075
rect 6570 -2105 6610 -2100
rect 6570 -2135 6575 -2105
rect 6575 -2135 6605 -2105
rect 6605 -2135 6610 -2105
rect 6570 -2140 6610 -2135
rect 6570 -2170 6610 -2165
rect 6570 -2200 6575 -2170
rect 6575 -2200 6605 -2170
rect 6605 -2200 6610 -2170
rect 6570 -2205 6610 -2200
rect 6570 -2240 6610 -2235
rect 6570 -2270 6575 -2240
rect 6575 -2270 6605 -2240
rect 6605 -2270 6610 -2240
rect 6570 -2275 6610 -2270
rect 6570 -2310 6610 -2305
rect 6570 -2340 6575 -2310
rect 6575 -2340 6605 -2310
rect 6605 -2340 6610 -2310
rect 6570 -2345 6610 -2340
rect 6570 -2380 6610 -2375
rect 6570 -2410 6575 -2380
rect 6575 -2410 6605 -2380
rect 6605 -2410 6610 -2380
rect 6570 -2415 6610 -2410
rect 6570 -2445 6610 -2440
rect 6570 -2475 6575 -2445
rect 6575 -2475 6605 -2445
rect 6605 -2475 6610 -2445
rect 6570 -2480 6610 -2475
rect 6570 -2505 6610 -2500
rect 6570 -2535 6575 -2505
rect 6575 -2535 6605 -2505
rect 6605 -2535 6610 -2505
rect 6570 -2540 6610 -2535
rect 6570 -2570 6610 -2565
rect 6570 -2600 6575 -2570
rect 6575 -2600 6605 -2570
rect 6605 -2600 6610 -2570
rect 6570 -2605 6610 -2600
rect 6570 -2640 6610 -2635
rect 6570 -2670 6575 -2640
rect 6575 -2670 6605 -2640
rect 6605 -2670 6610 -2640
rect 6570 -2675 6610 -2670
rect 6570 -2710 6610 -2705
rect 6570 -2740 6575 -2710
rect 6575 -2740 6605 -2710
rect 6605 -2740 6610 -2710
rect 6570 -2745 6610 -2740
rect 6570 -2780 6610 -2775
rect 6570 -2810 6575 -2780
rect 6575 -2810 6605 -2780
rect 6605 -2810 6610 -2780
rect 6570 -2815 6610 -2810
rect 6570 -2845 6610 -2840
rect 6570 -2875 6575 -2845
rect 6575 -2875 6605 -2845
rect 6605 -2875 6610 -2845
rect 6570 -2880 6610 -2875
rect 6570 -2905 6610 -2900
rect 6570 -2935 6575 -2905
rect 6575 -2935 6605 -2905
rect 6605 -2935 6610 -2905
rect 6570 -2940 6610 -2935
rect 6570 -2970 6610 -2965
rect 6570 -3000 6575 -2970
rect 6575 -3000 6605 -2970
rect 6605 -3000 6610 -2970
rect 6570 -3005 6610 -3000
rect 6570 -3040 6610 -3035
rect 6570 -3070 6575 -3040
rect 6575 -3070 6605 -3040
rect 6605 -3070 6610 -3040
rect 6570 -3075 6610 -3070
rect 6570 -3110 6610 -3105
rect 6570 -3140 6575 -3110
rect 6575 -3140 6605 -3110
rect 6605 -3140 6610 -3110
rect 6570 -3145 6610 -3140
rect 6570 -3180 6610 -3175
rect 6570 -3210 6575 -3180
rect 6575 -3210 6605 -3180
rect 6605 -3210 6610 -3180
rect 6570 -3215 6610 -3210
rect 6570 -3245 6610 -3240
rect 6570 -3275 6575 -3245
rect 6575 -3275 6605 -3245
rect 6605 -3275 6610 -3245
rect 6570 -3280 6610 -3275
rect 6570 -3305 6610 -3300
rect 6570 -3335 6575 -3305
rect 6575 -3335 6605 -3305
rect 6605 -3335 6610 -3305
rect 6570 -3340 6610 -3335
rect 6570 -3370 6610 -3365
rect 6570 -3400 6575 -3370
rect 6575 -3400 6605 -3370
rect 6605 -3400 6610 -3370
rect 6570 -3405 6610 -3400
rect 6570 -3440 6610 -3435
rect 6570 -3470 6575 -3440
rect 6575 -3470 6605 -3440
rect 6605 -3470 6610 -3440
rect 6570 -3475 6610 -3470
rect 6570 -3510 6610 -3505
rect 6570 -3540 6575 -3510
rect 6575 -3540 6605 -3510
rect 6605 -3540 6610 -3510
rect 6570 -3545 6610 -3540
rect 6570 -3580 6610 -3575
rect 6570 -3610 6575 -3580
rect 6575 -3610 6605 -3580
rect 6605 -3610 6610 -3580
rect 6570 -3615 6610 -3610
rect 6570 -3645 6610 -3640
rect 6570 -3675 6575 -3645
rect 6575 -3675 6605 -3645
rect 6605 -3675 6610 -3645
rect 6570 -3680 6610 -3675
rect 6570 -3705 6610 -3700
rect 6570 -3735 6575 -3705
rect 6575 -3735 6605 -3705
rect 6605 -3735 6610 -3705
rect 6570 -3740 6610 -3735
rect 6570 -3770 6610 -3765
rect 6570 -3800 6575 -3770
rect 6575 -3800 6605 -3770
rect 6605 -3800 6610 -3770
rect 6570 -3805 6610 -3800
rect 6570 -3840 6610 -3835
rect 6570 -3870 6575 -3840
rect 6575 -3870 6605 -3840
rect 6605 -3870 6610 -3840
rect 6570 -3875 6610 -3870
rect 6570 -3910 6610 -3905
rect 6570 -3940 6575 -3910
rect 6575 -3940 6605 -3910
rect 6605 -3940 6610 -3910
rect 6570 -3945 6610 -3940
rect 6570 -3980 6610 -3975
rect 6570 -4010 6575 -3980
rect 6575 -4010 6605 -3980
rect 6605 -4010 6610 -3980
rect 6570 -4015 6610 -4010
rect 6570 -4045 6610 -4040
rect 6570 -4075 6575 -4045
rect 6575 -4075 6605 -4045
rect 6605 -4075 6610 -4045
rect 6570 -4080 6610 -4075
rect 6570 -4105 6610 -4100
rect 6570 -4135 6575 -4105
rect 6575 -4135 6605 -4105
rect 6605 -4135 6610 -4105
rect 6570 -4140 6610 -4135
rect 6570 -4170 6610 -4165
rect 6570 -4200 6575 -4170
rect 6575 -4200 6605 -4170
rect 6605 -4200 6610 -4170
rect 6570 -4205 6610 -4200
rect 6570 -4240 6610 -4235
rect 6570 -4270 6575 -4240
rect 6575 -4270 6605 -4240
rect 6605 -4270 6610 -4240
rect 6570 -4275 6610 -4270
rect 6570 -4310 6610 -4305
rect 6570 -4340 6575 -4310
rect 6575 -4340 6605 -4310
rect 6605 -4340 6610 -4310
rect 6570 -4345 6610 -4340
rect 6570 -4380 6610 -4375
rect 6570 -4410 6575 -4380
rect 6575 -4410 6605 -4380
rect 6605 -4410 6610 -4380
rect 6570 -4415 6610 -4410
rect 6570 -4445 6610 -4440
rect 6570 -4475 6575 -4445
rect 6575 -4475 6605 -4445
rect 6605 -4475 6610 -4445
rect 6570 -4480 6610 -4475
rect 6920 -1305 6960 -1300
rect 6920 -1335 6925 -1305
rect 6925 -1335 6955 -1305
rect 6955 -1335 6960 -1305
rect 6920 -1340 6960 -1335
rect 6920 -1370 6960 -1365
rect 6920 -1400 6925 -1370
rect 6925 -1400 6955 -1370
rect 6955 -1400 6960 -1370
rect 6920 -1405 6960 -1400
rect 6920 -1440 6960 -1435
rect 6920 -1470 6925 -1440
rect 6925 -1470 6955 -1440
rect 6955 -1470 6960 -1440
rect 6920 -1475 6960 -1470
rect 6920 -1510 6960 -1505
rect 6920 -1540 6925 -1510
rect 6925 -1540 6955 -1510
rect 6955 -1540 6960 -1510
rect 6920 -1545 6960 -1540
rect 6920 -1580 6960 -1575
rect 6920 -1610 6925 -1580
rect 6925 -1610 6955 -1580
rect 6955 -1610 6960 -1580
rect 6920 -1615 6960 -1610
rect 6920 -1645 6960 -1640
rect 6920 -1675 6925 -1645
rect 6925 -1675 6955 -1645
rect 6955 -1675 6960 -1645
rect 6920 -1680 6960 -1675
rect 6920 -1705 6960 -1700
rect 6920 -1735 6925 -1705
rect 6925 -1735 6955 -1705
rect 6955 -1735 6960 -1705
rect 6920 -1740 6960 -1735
rect 6920 -1770 6960 -1765
rect 6920 -1800 6925 -1770
rect 6925 -1800 6955 -1770
rect 6955 -1800 6960 -1770
rect 6920 -1805 6960 -1800
rect 6920 -1840 6960 -1835
rect 6920 -1870 6925 -1840
rect 6925 -1870 6955 -1840
rect 6955 -1870 6960 -1840
rect 6920 -1875 6960 -1870
rect 6920 -1910 6960 -1905
rect 6920 -1940 6925 -1910
rect 6925 -1940 6955 -1910
rect 6955 -1940 6960 -1910
rect 6920 -1945 6960 -1940
rect 6920 -1980 6960 -1975
rect 6920 -2010 6925 -1980
rect 6925 -2010 6955 -1980
rect 6955 -2010 6960 -1980
rect 6920 -2015 6960 -2010
rect 6920 -2045 6960 -2040
rect 6920 -2075 6925 -2045
rect 6925 -2075 6955 -2045
rect 6955 -2075 6960 -2045
rect 6920 -2080 6960 -2075
rect 6920 -2105 6960 -2100
rect 6920 -2135 6925 -2105
rect 6925 -2135 6955 -2105
rect 6955 -2135 6960 -2105
rect 6920 -2140 6960 -2135
rect 6920 -2170 6960 -2165
rect 6920 -2200 6925 -2170
rect 6925 -2200 6955 -2170
rect 6955 -2200 6960 -2170
rect 6920 -2205 6960 -2200
rect 6920 -2240 6960 -2235
rect 6920 -2270 6925 -2240
rect 6925 -2270 6955 -2240
rect 6955 -2270 6960 -2240
rect 6920 -2275 6960 -2270
rect 6920 -2310 6960 -2305
rect 6920 -2340 6925 -2310
rect 6925 -2340 6955 -2310
rect 6955 -2340 6960 -2310
rect 6920 -2345 6960 -2340
rect 6920 -2380 6960 -2375
rect 6920 -2410 6925 -2380
rect 6925 -2410 6955 -2380
rect 6955 -2410 6960 -2380
rect 6920 -2415 6960 -2410
rect 6920 -2445 6960 -2440
rect 6920 -2475 6925 -2445
rect 6925 -2475 6955 -2445
rect 6955 -2475 6960 -2445
rect 6920 -2480 6960 -2475
rect 6920 -2505 6960 -2500
rect 6920 -2535 6925 -2505
rect 6925 -2535 6955 -2505
rect 6955 -2535 6960 -2505
rect 6920 -2540 6960 -2535
rect 6920 -2570 6960 -2565
rect 6920 -2600 6925 -2570
rect 6925 -2600 6955 -2570
rect 6955 -2600 6960 -2570
rect 6920 -2605 6960 -2600
rect 6920 -2640 6960 -2635
rect 6920 -2670 6925 -2640
rect 6925 -2670 6955 -2640
rect 6955 -2670 6960 -2640
rect 6920 -2675 6960 -2670
rect 6920 -2710 6960 -2705
rect 6920 -2740 6925 -2710
rect 6925 -2740 6955 -2710
rect 6955 -2740 6960 -2710
rect 6920 -2745 6960 -2740
rect 6920 -2780 6960 -2775
rect 6920 -2810 6925 -2780
rect 6925 -2810 6955 -2780
rect 6955 -2810 6960 -2780
rect 6920 -2815 6960 -2810
rect 6920 -2845 6960 -2840
rect 6920 -2875 6925 -2845
rect 6925 -2875 6955 -2845
rect 6955 -2875 6960 -2845
rect 6920 -2880 6960 -2875
rect 6920 -2905 6960 -2900
rect 6920 -2935 6925 -2905
rect 6925 -2935 6955 -2905
rect 6955 -2935 6960 -2905
rect 6920 -2940 6960 -2935
rect 6920 -2970 6960 -2965
rect 6920 -3000 6925 -2970
rect 6925 -3000 6955 -2970
rect 6955 -3000 6960 -2970
rect 6920 -3005 6960 -3000
rect 6920 -3040 6960 -3035
rect 6920 -3070 6925 -3040
rect 6925 -3070 6955 -3040
rect 6955 -3070 6960 -3040
rect 6920 -3075 6960 -3070
rect 6920 -3110 6960 -3105
rect 6920 -3140 6925 -3110
rect 6925 -3140 6955 -3110
rect 6955 -3140 6960 -3110
rect 6920 -3145 6960 -3140
rect 6920 -3180 6960 -3175
rect 6920 -3210 6925 -3180
rect 6925 -3210 6955 -3180
rect 6955 -3210 6960 -3180
rect 6920 -3215 6960 -3210
rect 6920 -3245 6960 -3240
rect 6920 -3275 6925 -3245
rect 6925 -3275 6955 -3245
rect 6955 -3275 6960 -3245
rect 6920 -3280 6960 -3275
rect 6920 -3305 6960 -3300
rect 6920 -3335 6925 -3305
rect 6925 -3335 6955 -3305
rect 6955 -3335 6960 -3305
rect 6920 -3340 6960 -3335
rect 6920 -3370 6960 -3365
rect 6920 -3400 6925 -3370
rect 6925 -3400 6955 -3370
rect 6955 -3400 6960 -3370
rect 6920 -3405 6960 -3400
rect 6920 -3440 6960 -3435
rect 6920 -3470 6925 -3440
rect 6925 -3470 6955 -3440
rect 6955 -3470 6960 -3440
rect 6920 -3475 6960 -3470
rect 6920 -3510 6960 -3505
rect 6920 -3540 6925 -3510
rect 6925 -3540 6955 -3510
rect 6955 -3540 6960 -3510
rect 6920 -3545 6960 -3540
rect 6920 -3580 6960 -3575
rect 6920 -3610 6925 -3580
rect 6925 -3610 6955 -3580
rect 6955 -3610 6960 -3580
rect 6920 -3615 6960 -3610
rect 6920 -3645 6960 -3640
rect 6920 -3675 6925 -3645
rect 6925 -3675 6955 -3645
rect 6955 -3675 6960 -3645
rect 6920 -3680 6960 -3675
rect 6920 -3705 6960 -3700
rect 6920 -3735 6925 -3705
rect 6925 -3735 6955 -3705
rect 6955 -3735 6960 -3705
rect 6920 -3740 6960 -3735
rect 6920 -3770 6960 -3765
rect 6920 -3800 6925 -3770
rect 6925 -3800 6955 -3770
rect 6955 -3800 6960 -3770
rect 6920 -3805 6960 -3800
rect 6920 -3840 6960 -3835
rect 6920 -3870 6925 -3840
rect 6925 -3870 6955 -3840
rect 6955 -3870 6960 -3840
rect 6920 -3875 6960 -3870
rect 6920 -3910 6960 -3905
rect 6920 -3940 6925 -3910
rect 6925 -3940 6955 -3910
rect 6955 -3940 6960 -3910
rect 6920 -3945 6960 -3940
rect 6920 -3980 6960 -3975
rect 6920 -4010 6925 -3980
rect 6925 -4010 6955 -3980
rect 6955 -4010 6960 -3980
rect 6920 -4015 6960 -4010
rect 6920 -4045 6960 -4040
rect 6920 -4075 6925 -4045
rect 6925 -4075 6955 -4045
rect 6955 -4075 6960 -4045
rect 6920 -4080 6960 -4075
rect 6920 -4105 6960 -4100
rect 6920 -4135 6925 -4105
rect 6925 -4135 6955 -4105
rect 6955 -4135 6960 -4105
rect 6920 -4140 6960 -4135
rect 6920 -4170 6960 -4165
rect 6920 -4200 6925 -4170
rect 6925 -4200 6955 -4170
rect 6955 -4200 6960 -4170
rect 6920 -4205 6960 -4200
rect 6920 -4240 6960 -4235
rect 6920 -4270 6925 -4240
rect 6925 -4270 6955 -4240
rect 6955 -4270 6960 -4240
rect 6920 -4275 6960 -4270
rect 6920 -4310 6960 -4305
rect 6920 -4340 6925 -4310
rect 6925 -4340 6955 -4310
rect 6955 -4340 6960 -4310
rect 6920 -4345 6960 -4340
rect 6920 -4380 6960 -4375
rect 6920 -4410 6925 -4380
rect 6925 -4410 6955 -4380
rect 6955 -4410 6960 -4380
rect 6920 -4415 6960 -4410
rect 6920 -4445 6960 -4440
rect 6920 -4475 6925 -4445
rect 6925 -4475 6955 -4445
rect 6955 -4475 6960 -4445
rect 6920 -4480 6960 -4475
rect 7270 -1305 7310 -1300
rect 7270 -1335 7275 -1305
rect 7275 -1335 7305 -1305
rect 7305 -1335 7310 -1305
rect 7270 -1340 7310 -1335
rect 7270 -1370 7310 -1365
rect 7270 -1400 7275 -1370
rect 7275 -1400 7305 -1370
rect 7305 -1400 7310 -1370
rect 7270 -1405 7310 -1400
rect 7270 -1440 7310 -1435
rect 7270 -1470 7275 -1440
rect 7275 -1470 7305 -1440
rect 7305 -1470 7310 -1440
rect 7270 -1475 7310 -1470
rect 7270 -1510 7310 -1505
rect 7270 -1540 7275 -1510
rect 7275 -1540 7305 -1510
rect 7305 -1540 7310 -1510
rect 7270 -1545 7310 -1540
rect 7270 -1580 7310 -1575
rect 7270 -1610 7275 -1580
rect 7275 -1610 7305 -1580
rect 7305 -1610 7310 -1580
rect 7270 -1615 7310 -1610
rect 7270 -1645 7310 -1640
rect 7270 -1675 7275 -1645
rect 7275 -1675 7305 -1645
rect 7305 -1675 7310 -1645
rect 7270 -1680 7310 -1675
rect 7270 -1705 7310 -1700
rect 7270 -1735 7275 -1705
rect 7275 -1735 7305 -1705
rect 7305 -1735 7310 -1705
rect 7270 -1740 7310 -1735
rect 7270 -1770 7310 -1765
rect 7270 -1800 7275 -1770
rect 7275 -1800 7305 -1770
rect 7305 -1800 7310 -1770
rect 7270 -1805 7310 -1800
rect 7270 -1840 7310 -1835
rect 7270 -1870 7275 -1840
rect 7275 -1870 7305 -1840
rect 7305 -1870 7310 -1840
rect 7270 -1875 7310 -1870
rect 7270 -1910 7310 -1905
rect 7270 -1940 7275 -1910
rect 7275 -1940 7305 -1910
rect 7305 -1940 7310 -1910
rect 7270 -1945 7310 -1940
rect 7270 -1980 7310 -1975
rect 7270 -2010 7275 -1980
rect 7275 -2010 7305 -1980
rect 7305 -2010 7310 -1980
rect 7270 -2015 7310 -2010
rect 7270 -2045 7310 -2040
rect 7270 -2075 7275 -2045
rect 7275 -2075 7305 -2045
rect 7305 -2075 7310 -2045
rect 7270 -2080 7310 -2075
rect 7270 -2105 7310 -2100
rect 7270 -2135 7275 -2105
rect 7275 -2135 7305 -2105
rect 7305 -2135 7310 -2105
rect 7270 -2140 7310 -2135
rect 7270 -2170 7310 -2165
rect 7270 -2200 7275 -2170
rect 7275 -2200 7305 -2170
rect 7305 -2200 7310 -2170
rect 7270 -2205 7310 -2200
rect 7270 -2240 7310 -2235
rect 7270 -2270 7275 -2240
rect 7275 -2270 7305 -2240
rect 7305 -2270 7310 -2240
rect 7270 -2275 7310 -2270
rect 7270 -2310 7310 -2305
rect 7270 -2340 7275 -2310
rect 7275 -2340 7305 -2310
rect 7305 -2340 7310 -2310
rect 7270 -2345 7310 -2340
rect 7270 -2380 7310 -2375
rect 7270 -2410 7275 -2380
rect 7275 -2410 7305 -2380
rect 7305 -2410 7310 -2380
rect 7270 -2415 7310 -2410
rect 7270 -2445 7310 -2440
rect 7270 -2475 7275 -2445
rect 7275 -2475 7305 -2445
rect 7305 -2475 7310 -2445
rect 7270 -2480 7310 -2475
rect 7270 -2505 7310 -2500
rect 7270 -2535 7275 -2505
rect 7275 -2535 7305 -2505
rect 7305 -2535 7310 -2505
rect 7270 -2540 7310 -2535
rect 7270 -2570 7310 -2565
rect 7270 -2600 7275 -2570
rect 7275 -2600 7305 -2570
rect 7305 -2600 7310 -2570
rect 7270 -2605 7310 -2600
rect 7270 -2640 7310 -2635
rect 7270 -2670 7275 -2640
rect 7275 -2670 7305 -2640
rect 7305 -2670 7310 -2640
rect 7270 -2675 7310 -2670
rect 7270 -2710 7310 -2705
rect 7270 -2740 7275 -2710
rect 7275 -2740 7305 -2710
rect 7305 -2740 7310 -2710
rect 7270 -2745 7310 -2740
rect 7270 -2780 7310 -2775
rect 7270 -2810 7275 -2780
rect 7275 -2810 7305 -2780
rect 7305 -2810 7310 -2780
rect 7270 -2815 7310 -2810
rect 7270 -2845 7310 -2840
rect 7270 -2875 7275 -2845
rect 7275 -2875 7305 -2845
rect 7305 -2875 7310 -2845
rect 7270 -2880 7310 -2875
rect 7270 -2905 7310 -2900
rect 7270 -2935 7275 -2905
rect 7275 -2935 7305 -2905
rect 7305 -2935 7310 -2905
rect 7270 -2940 7310 -2935
rect 7270 -2970 7310 -2965
rect 7270 -3000 7275 -2970
rect 7275 -3000 7305 -2970
rect 7305 -3000 7310 -2970
rect 7270 -3005 7310 -3000
rect 7270 -3040 7310 -3035
rect 7270 -3070 7275 -3040
rect 7275 -3070 7305 -3040
rect 7305 -3070 7310 -3040
rect 7270 -3075 7310 -3070
rect 7270 -3110 7310 -3105
rect 7270 -3140 7275 -3110
rect 7275 -3140 7305 -3110
rect 7305 -3140 7310 -3110
rect 7270 -3145 7310 -3140
rect 7270 -3180 7310 -3175
rect 7270 -3210 7275 -3180
rect 7275 -3210 7305 -3180
rect 7305 -3210 7310 -3180
rect 7270 -3215 7310 -3210
rect 7270 -3245 7310 -3240
rect 7270 -3275 7275 -3245
rect 7275 -3275 7305 -3245
rect 7305 -3275 7310 -3245
rect 7270 -3280 7310 -3275
rect 7270 -3305 7310 -3300
rect 7270 -3335 7275 -3305
rect 7275 -3335 7305 -3305
rect 7305 -3335 7310 -3305
rect 7270 -3340 7310 -3335
rect 7270 -3370 7310 -3365
rect 7270 -3400 7275 -3370
rect 7275 -3400 7305 -3370
rect 7305 -3400 7310 -3370
rect 7270 -3405 7310 -3400
rect 7270 -3440 7310 -3435
rect 7270 -3470 7275 -3440
rect 7275 -3470 7305 -3440
rect 7305 -3470 7310 -3440
rect 7270 -3475 7310 -3470
rect 7270 -3510 7310 -3505
rect 7270 -3540 7275 -3510
rect 7275 -3540 7305 -3510
rect 7305 -3540 7310 -3510
rect 7270 -3545 7310 -3540
rect 7270 -3580 7310 -3575
rect 7270 -3610 7275 -3580
rect 7275 -3610 7305 -3580
rect 7305 -3610 7310 -3580
rect 7270 -3615 7310 -3610
rect 7270 -3645 7310 -3640
rect 7270 -3675 7275 -3645
rect 7275 -3675 7305 -3645
rect 7305 -3675 7310 -3645
rect 7270 -3680 7310 -3675
rect 7270 -3705 7310 -3700
rect 7270 -3735 7275 -3705
rect 7275 -3735 7305 -3705
rect 7305 -3735 7310 -3705
rect 7270 -3740 7310 -3735
rect 7270 -3770 7310 -3765
rect 7270 -3800 7275 -3770
rect 7275 -3800 7305 -3770
rect 7305 -3800 7310 -3770
rect 7270 -3805 7310 -3800
rect 7270 -3840 7310 -3835
rect 7270 -3870 7275 -3840
rect 7275 -3870 7305 -3840
rect 7305 -3870 7310 -3840
rect 7270 -3875 7310 -3870
rect 7270 -3910 7310 -3905
rect 7270 -3940 7275 -3910
rect 7275 -3940 7305 -3910
rect 7305 -3940 7310 -3910
rect 7270 -3945 7310 -3940
rect 7270 -3980 7310 -3975
rect 7270 -4010 7275 -3980
rect 7275 -4010 7305 -3980
rect 7305 -4010 7310 -3980
rect 7270 -4015 7310 -4010
rect 7270 -4045 7310 -4040
rect 7270 -4075 7275 -4045
rect 7275 -4075 7305 -4045
rect 7305 -4075 7310 -4045
rect 7270 -4080 7310 -4075
rect 7270 -4105 7310 -4100
rect 7270 -4135 7275 -4105
rect 7275 -4135 7305 -4105
rect 7305 -4135 7310 -4105
rect 7270 -4140 7310 -4135
rect 7270 -4170 7310 -4165
rect 7270 -4200 7275 -4170
rect 7275 -4200 7305 -4170
rect 7305 -4200 7310 -4170
rect 7270 -4205 7310 -4200
rect 7270 -4240 7310 -4235
rect 7270 -4270 7275 -4240
rect 7275 -4270 7305 -4240
rect 7305 -4270 7310 -4240
rect 7270 -4275 7310 -4270
rect 7270 -4310 7310 -4305
rect 7270 -4340 7275 -4310
rect 7275 -4340 7305 -4310
rect 7305 -4340 7310 -4310
rect 7270 -4345 7310 -4340
rect 7270 -4380 7310 -4375
rect 7270 -4410 7275 -4380
rect 7275 -4410 7305 -4380
rect 7305 -4410 7310 -4380
rect 7270 -4415 7310 -4410
rect 7270 -4445 7310 -4440
rect 7270 -4475 7275 -4445
rect 7275 -4475 7305 -4445
rect 7305 -4475 7310 -4445
rect 7270 -4480 7310 -4475
rect 7620 -1305 7660 -1300
rect 7620 -1335 7625 -1305
rect 7625 -1335 7655 -1305
rect 7655 -1335 7660 -1305
rect 7620 -1340 7660 -1335
rect 7620 -1370 7660 -1365
rect 7620 -1400 7625 -1370
rect 7625 -1400 7655 -1370
rect 7655 -1400 7660 -1370
rect 7620 -1405 7660 -1400
rect 7620 -1440 7660 -1435
rect 7620 -1470 7625 -1440
rect 7625 -1470 7655 -1440
rect 7655 -1470 7660 -1440
rect 7620 -1475 7660 -1470
rect 7620 -1510 7660 -1505
rect 7620 -1540 7625 -1510
rect 7625 -1540 7655 -1510
rect 7655 -1540 7660 -1510
rect 7620 -1545 7660 -1540
rect 7620 -1580 7660 -1575
rect 7620 -1610 7625 -1580
rect 7625 -1610 7655 -1580
rect 7655 -1610 7660 -1580
rect 7620 -1615 7660 -1610
rect 7620 -1645 7660 -1640
rect 7620 -1675 7625 -1645
rect 7625 -1675 7655 -1645
rect 7655 -1675 7660 -1645
rect 7620 -1680 7660 -1675
rect 7620 -1705 7660 -1700
rect 7620 -1735 7625 -1705
rect 7625 -1735 7655 -1705
rect 7655 -1735 7660 -1705
rect 7620 -1740 7660 -1735
rect 7620 -1770 7660 -1765
rect 7620 -1800 7625 -1770
rect 7625 -1800 7655 -1770
rect 7655 -1800 7660 -1770
rect 7620 -1805 7660 -1800
rect 7620 -1840 7660 -1835
rect 7620 -1870 7625 -1840
rect 7625 -1870 7655 -1840
rect 7655 -1870 7660 -1840
rect 7620 -1875 7660 -1870
rect 7620 -1910 7660 -1905
rect 7620 -1940 7625 -1910
rect 7625 -1940 7655 -1910
rect 7655 -1940 7660 -1910
rect 7620 -1945 7660 -1940
rect 7620 -1980 7660 -1975
rect 7620 -2010 7625 -1980
rect 7625 -2010 7655 -1980
rect 7655 -2010 7660 -1980
rect 7620 -2015 7660 -2010
rect 7620 -2045 7660 -2040
rect 7620 -2075 7625 -2045
rect 7625 -2075 7655 -2045
rect 7655 -2075 7660 -2045
rect 7620 -2080 7660 -2075
rect 7620 -2105 7660 -2100
rect 7620 -2135 7625 -2105
rect 7625 -2135 7655 -2105
rect 7655 -2135 7660 -2105
rect 7620 -2140 7660 -2135
rect 7620 -2170 7660 -2165
rect 7620 -2200 7625 -2170
rect 7625 -2200 7655 -2170
rect 7655 -2200 7660 -2170
rect 7620 -2205 7660 -2200
rect 7620 -2240 7660 -2235
rect 7620 -2270 7625 -2240
rect 7625 -2270 7655 -2240
rect 7655 -2270 7660 -2240
rect 7620 -2275 7660 -2270
rect 7620 -2310 7660 -2305
rect 7620 -2340 7625 -2310
rect 7625 -2340 7655 -2310
rect 7655 -2340 7660 -2310
rect 7620 -2345 7660 -2340
rect 7620 -2380 7660 -2375
rect 7620 -2410 7625 -2380
rect 7625 -2410 7655 -2380
rect 7655 -2410 7660 -2380
rect 7620 -2415 7660 -2410
rect 7620 -2445 7660 -2440
rect 7620 -2475 7625 -2445
rect 7625 -2475 7655 -2445
rect 7655 -2475 7660 -2445
rect 7620 -2480 7660 -2475
rect 7620 -2505 7660 -2500
rect 7620 -2535 7625 -2505
rect 7625 -2535 7655 -2505
rect 7655 -2535 7660 -2505
rect 7620 -2540 7660 -2535
rect 7620 -2570 7660 -2565
rect 7620 -2600 7625 -2570
rect 7625 -2600 7655 -2570
rect 7655 -2600 7660 -2570
rect 7620 -2605 7660 -2600
rect 7620 -2640 7660 -2635
rect 7620 -2670 7625 -2640
rect 7625 -2670 7655 -2640
rect 7655 -2670 7660 -2640
rect 7620 -2675 7660 -2670
rect 7620 -2710 7660 -2705
rect 7620 -2740 7625 -2710
rect 7625 -2740 7655 -2710
rect 7655 -2740 7660 -2710
rect 7620 -2745 7660 -2740
rect 7620 -2780 7660 -2775
rect 7620 -2810 7625 -2780
rect 7625 -2810 7655 -2780
rect 7655 -2810 7660 -2780
rect 7620 -2815 7660 -2810
rect 7620 -2845 7660 -2840
rect 7620 -2875 7625 -2845
rect 7625 -2875 7655 -2845
rect 7655 -2875 7660 -2845
rect 7620 -2880 7660 -2875
rect 7620 -2905 7660 -2900
rect 7620 -2935 7625 -2905
rect 7625 -2935 7655 -2905
rect 7655 -2935 7660 -2905
rect 7620 -2940 7660 -2935
rect 7620 -2970 7660 -2965
rect 7620 -3000 7625 -2970
rect 7625 -3000 7655 -2970
rect 7655 -3000 7660 -2970
rect 7620 -3005 7660 -3000
rect 7620 -3040 7660 -3035
rect 7620 -3070 7625 -3040
rect 7625 -3070 7655 -3040
rect 7655 -3070 7660 -3040
rect 7620 -3075 7660 -3070
rect 7620 -3110 7660 -3105
rect 7620 -3140 7625 -3110
rect 7625 -3140 7655 -3110
rect 7655 -3140 7660 -3110
rect 7620 -3145 7660 -3140
rect 7620 -3180 7660 -3175
rect 7620 -3210 7625 -3180
rect 7625 -3210 7655 -3180
rect 7655 -3210 7660 -3180
rect 7620 -3215 7660 -3210
rect 7620 -3245 7660 -3240
rect 7620 -3275 7625 -3245
rect 7625 -3275 7655 -3245
rect 7655 -3275 7660 -3245
rect 7620 -3280 7660 -3275
rect 7620 -3305 7660 -3300
rect 7620 -3335 7625 -3305
rect 7625 -3335 7655 -3305
rect 7655 -3335 7660 -3305
rect 7620 -3340 7660 -3335
rect 7620 -3370 7660 -3365
rect 7620 -3400 7625 -3370
rect 7625 -3400 7655 -3370
rect 7655 -3400 7660 -3370
rect 7620 -3405 7660 -3400
rect 7620 -3440 7660 -3435
rect 7620 -3470 7625 -3440
rect 7625 -3470 7655 -3440
rect 7655 -3470 7660 -3440
rect 7620 -3475 7660 -3470
rect 7620 -3510 7660 -3505
rect 7620 -3540 7625 -3510
rect 7625 -3540 7655 -3510
rect 7655 -3540 7660 -3510
rect 7620 -3545 7660 -3540
rect 7620 -3580 7660 -3575
rect 7620 -3610 7625 -3580
rect 7625 -3610 7655 -3580
rect 7655 -3610 7660 -3580
rect 7620 -3615 7660 -3610
rect 7620 -3645 7660 -3640
rect 7620 -3675 7625 -3645
rect 7625 -3675 7655 -3645
rect 7655 -3675 7660 -3645
rect 7620 -3680 7660 -3675
rect 7620 -3705 7660 -3700
rect 7620 -3735 7625 -3705
rect 7625 -3735 7655 -3705
rect 7655 -3735 7660 -3705
rect 7620 -3740 7660 -3735
rect 7620 -3770 7660 -3765
rect 7620 -3800 7625 -3770
rect 7625 -3800 7655 -3770
rect 7655 -3800 7660 -3770
rect 7620 -3805 7660 -3800
rect 7620 -3840 7660 -3835
rect 7620 -3870 7625 -3840
rect 7625 -3870 7655 -3840
rect 7655 -3870 7660 -3840
rect 7620 -3875 7660 -3870
rect 7620 -3910 7660 -3905
rect 7620 -3940 7625 -3910
rect 7625 -3940 7655 -3910
rect 7655 -3940 7660 -3910
rect 7620 -3945 7660 -3940
rect 7620 -3980 7660 -3975
rect 7620 -4010 7625 -3980
rect 7625 -4010 7655 -3980
rect 7655 -4010 7660 -3980
rect 7620 -4015 7660 -4010
rect 7620 -4045 7660 -4040
rect 7620 -4075 7625 -4045
rect 7625 -4075 7655 -4045
rect 7655 -4075 7660 -4045
rect 7620 -4080 7660 -4075
rect 7620 -4105 7660 -4100
rect 7620 -4135 7625 -4105
rect 7625 -4135 7655 -4105
rect 7655 -4135 7660 -4105
rect 7620 -4140 7660 -4135
rect 7620 -4170 7660 -4165
rect 7620 -4200 7625 -4170
rect 7625 -4200 7655 -4170
rect 7655 -4200 7660 -4170
rect 7620 -4205 7660 -4200
rect 7620 -4240 7660 -4235
rect 7620 -4270 7625 -4240
rect 7625 -4270 7655 -4240
rect 7655 -4270 7660 -4240
rect 7620 -4275 7660 -4270
rect 7620 -4310 7660 -4305
rect 7620 -4340 7625 -4310
rect 7625 -4340 7655 -4310
rect 7655 -4340 7660 -4310
rect 7620 -4345 7660 -4340
rect 7620 -4380 7660 -4375
rect 7620 -4410 7625 -4380
rect 7625 -4410 7655 -4380
rect 7655 -4410 7660 -4380
rect 7620 -4415 7660 -4410
rect 7620 -4445 7660 -4440
rect 7620 -4475 7625 -4445
rect 7625 -4475 7655 -4445
rect 7655 -4475 7660 -4445
rect 7620 -4480 7660 -4475
rect 7970 -1305 8010 -1300
rect 7970 -1335 7975 -1305
rect 7975 -1335 8005 -1305
rect 8005 -1335 8010 -1305
rect 7970 -1340 8010 -1335
rect 7970 -1370 8010 -1365
rect 7970 -1400 7975 -1370
rect 7975 -1400 8005 -1370
rect 8005 -1400 8010 -1370
rect 7970 -1405 8010 -1400
rect 7970 -1440 8010 -1435
rect 7970 -1470 7975 -1440
rect 7975 -1470 8005 -1440
rect 8005 -1470 8010 -1440
rect 7970 -1475 8010 -1470
rect 7970 -1510 8010 -1505
rect 7970 -1540 7975 -1510
rect 7975 -1540 8005 -1510
rect 8005 -1540 8010 -1510
rect 7970 -1545 8010 -1540
rect 7970 -1580 8010 -1575
rect 7970 -1610 7975 -1580
rect 7975 -1610 8005 -1580
rect 8005 -1610 8010 -1580
rect 7970 -1615 8010 -1610
rect 7970 -1645 8010 -1640
rect 7970 -1675 7975 -1645
rect 7975 -1675 8005 -1645
rect 8005 -1675 8010 -1645
rect 7970 -1680 8010 -1675
rect 7970 -1705 8010 -1700
rect 7970 -1735 7975 -1705
rect 7975 -1735 8005 -1705
rect 8005 -1735 8010 -1705
rect 7970 -1740 8010 -1735
rect 7970 -1770 8010 -1765
rect 7970 -1800 7975 -1770
rect 7975 -1800 8005 -1770
rect 8005 -1800 8010 -1770
rect 7970 -1805 8010 -1800
rect 7970 -1840 8010 -1835
rect 7970 -1870 7975 -1840
rect 7975 -1870 8005 -1840
rect 8005 -1870 8010 -1840
rect 7970 -1875 8010 -1870
rect 7970 -1910 8010 -1905
rect 7970 -1940 7975 -1910
rect 7975 -1940 8005 -1910
rect 8005 -1940 8010 -1910
rect 7970 -1945 8010 -1940
rect 7970 -1980 8010 -1975
rect 7970 -2010 7975 -1980
rect 7975 -2010 8005 -1980
rect 8005 -2010 8010 -1980
rect 7970 -2015 8010 -2010
rect 7970 -2045 8010 -2040
rect 7970 -2075 7975 -2045
rect 7975 -2075 8005 -2045
rect 8005 -2075 8010 -2045
rect 7970 -2080 8010 -2075
rect 7970 -2105 8010 -2100
rect 7970 -2135 7975 -2105
rect 7975 -2135 8005 -2105
rect 8005 -2135 8010 -2105
rect 7970 -2140 8010 -2135
rect 7970 -2170 8010 -2165
rect 7970 -2200 7975 -2170
rect 7975 -2200 8005 -2170
rect 8005 -2200 8010 -2170
rect 7970 -2205 8010 -2200
rect 7970 -2240 8010 -2235
rect 7970 -2270 7975 -2240
rect 7975 -2270 8005 -2240
rect 8005 -2270 8010 -2240
rect 7970 -2275 8010 -2270
rect 7970 -2310 8010 -2305
rect 7970 -2340 7975 -2310
rect 7975 -2340 8005 -2310
rect 8005 -2340 8010 -2310
rect 7970 -2345 8010 -2340
rect 7970 -2380 8010 -2375
rect 7970 -2410 7975 -2380
rect 7975 -2410 8005 -2380
rect 8005 -2410 8010 -2380
rect 7970 -2415 8010 -2410
rect 7970 -2445 8010 -2440
rect 7970 -2475 7975 -2445
rect 7975 -2475 8005 -2445
rect 8005 -2475 8010 -2445
rect 7970 -2480 8010 -2475
rect 7970 -2505 8010 -2500
rect 7970 -2535 7975 -2505
rect 7975 -2535 8005 -2505
rect 8005 -2535 8010 -2505
rect 7970 -2540 8010 -2535
rect 7970 -2570 8010 -2565
rect 7970 -2600 7975 -2570
rect 7975 -2600 8005 -2570
rect 8005 -2600 8010 -2570
rect 7970 -2605 8010 -2600
rect 7970 -2640 8010 -2635
rect 7970 -2670 7975 -2640
rect 7975 -2670 8005 -2640
rect 8005 -2670 8010 -2640
rect 7970 -2675 8010 -2670
rect 7970 -2710 8010 -2705
rect 7970 -2740 7975 -2710
rect 7975 -2740 8005 -2710
rect 8005 -2740 8010 -2710
rect 7970 -2745 8010 -2740
rect 7970 -2780 8010 -2775
rect 7970 -2810 7975 -2780
rect 7975 -2810 8005 -2780
rect 8005 -2810 8010 -2780
rect 7970 -2815 8010 -2810
rect 7970 -2845 8010 -2840
rect 7970 -2875 7975 -2845
rect 7975 -2875 8005 -2845
rect 8005 -2875 8010 -2845
rect 7970 -2880 8010 -2875
rect 7970 -2905 8010 -2900
rect 7970 -2935 7975 -2905
rect 7975 -2935 8005 -2905
rect 8005 -2935 8010 -2905
rect 7970 -2940 8010 -2935
rect 7970 -2970 8010 -2965
rect 7970 -3000 7975 -2970
rect 7975 -3000 8005 -2970
rect 8005 -3000 8010 -2970
rect 7970 -3005 8010 -3000
rect 7970 -3040 8010 -3035
rect 7970 -3070 7975 -3040
rect 7975 -3070 8005 -3040
rect 8005 -3070 8010 -3040
rect 7970 -3075 8010 -3070
rect 7970 -3110 8010 -3105
rect 7970 -3140 7975 -3110
rect 7975 -3140 8005 -3110
rect 8005 -3140 8010 -3110
rect 7970 -3145 8010 -3140
rect 7970 -3180 8010 -3175
rect 7970 -3210 7975 -3180
rect 7975 -3210 8005 -3180
rect 8005 -3210 8010 -3180
rect 7970 -3215 8010 -3210
rect 7970 -3245 8010 -3240
rect 7970 -3275 7975 -3245
rect 7975 -3275 8005 -3245
rect 8005 -3275 8010 -3245
rect 7970 -3280 8010 -3275
rect 7970 -3305 8010 -3300
rect 7970 -3335 7975 -3305
rect 7975 -3335 8005 -3305
rect 8005 -3335 8010 -3305
rect 7970 -3340 8010 -3335
rect 7970 -3370 8010 -3365
rect 7970 -3400 7975 -3370
rect 7975 -3400 8005 -3370
rect 8005 -3400 8010 -3370
rect 7970 -3405 8010 -3400
rect 7970 -3440 8010 -3435
rect 7970 -3470 7975 -3440
rect 7975 -3470 8005 -3440
rect 8005 -3470 8010 -3440
rect 7970 -3475 8010 -3470
rect 7970 -3510 8010 -3505
rect 7970 -3540 7975 -3510
rect 7975 -3540 8005 -3510
rect 8005 -3540 8010 -3510
rect 7970 -3545 8010 -3540
rect 7970 -3580 8010 -3575
rect 7970 -3610 7975 -3580
rect 7975 -3610 8005 -3580
rect 8005 -3610 8010 -3580
rect 7970 -3615 8010 -3610
rect 7970 -3645 8010 -3640
rect 7970 -3675 7975 -3645
rect 7975 -3675 8005 -3645
rect 8005 -3675 8010 -3645
rect 7970 -3680 8010 -3675
rect 7970 -3705 8010 -3700
rect 7970 -3735 7975 -3705
rect 7975 -3735 8005 -3705
rect 8005 -3735 8010 -3705
rect 7970 -3740 8010 -3735
rect 7970 -3770 8010 -3765
rect 7970 -3800 7975 -3770
rect 7975 -3800 8005 -3770
rect 8005 -3800 8010 -3770
rect 7970 -3805 8010 -3800
rect 7970 -3840 8010 -3835
rect 7970 -3870 7975 -3840
rect 7975 -3870 8005 -3840
rect 8005 -3870 8010 -3840
rect 7970 -3875 8010 -3870
rect 7970 -3910 8010 -3905
rect 7970 -3940 7975 -3910
rect 7975 -3940 8005 -3910
rect 8005 -3940 8010 -3910
rect 7970 -3945 8010 -3940
rect 7970 -3980 8010 -3975
rect 7970 -4010 7975 -3980
rect 7975 -4010 8005 -3980
rect 8005 -4010 8010 -3980
rect 7970 -4015 8010 -4010
rect 7970 -4045 8010 -4040
rect 7970 -4075 7975 -4045
rect 7975 -4075 8005 -4045
rect 8005 -4075 8010 -4045
rect 7970 -4080 8010 -4075
rect 7970 -4105 8010 -4100
rect 7970 -4135 7975 -4105
rect 7975 -4135 8005 -4105
rect 8005 -4135 8010 -4105
rect 7970 -4140 8010 -4135
rect 7970 -4170 8010 -4165
rect 7970 -4200 7975 -4170
rect 7975 -4200 8005 -4170
rect 8005 -4200 8010 -4170
rect 7970 -4205 8010 -4200
rect 7970 -4240 8010 -4235
rect 7970 -4270 7975 -4240
rect 7975 -4270 8005 -4240
rect 8005 -4270 8010 -4240
rect 7970 -4275 8010 -4270
rect 7970 -4310 8010 -4305
rect 7970 -4340 7975 -4310
rect 7975 -4340 8005 -4310
rect 8005 -4340 8010 -4310
rect 7970 -4345 8010 -4340
rect 7970 -4380 8010 -4375
rect 7970 -4410 7975 -4380
rect 7975 -4410 8005 -4380
rect 8005 -4410 8010 -4380
rect 7970 -4415 8010 -4410
rect 7970 -4445 8010 -4440
rect 7970 -4475 7975 -4445
rect 7975 -4475 8005 -4445
rect 8005 -4475 8010 -4445
rect 7970 -4480 8010 -4475
rect 8320 -1305 8360 -1300
rect 8320 -1335 8325 -1305
rect 8325 -1335 8355 -1305
rect 8355 -1335 8360 -1305
rect 8320 -1340 8360 -1335
rect 8320 -1370 8360 -1365
rect 8320 -1400 8325 -1370
rect 8325 -1400 8355 -1370
rect 8355 -1400 8360 -1370
rect 8320 -1405 8360 -1400
rect 8320 -1440 8360 -1435
rect 8320 -1470 8325 -1440
rect 8325 -1470 8355 -1440
rect 8355 -1470 8360 -1440
rect 8320 -1475 8360 -1470
rect 8320 -1510 8360 -1505
rect 8320 -1540 8325 -1510
rect 8325 -1540 8355 -1510
rect 8355 -1540 8360 -1510
rect 8320 -1545 8360 -1540
rect 8320 -1580 8360 -1575
rect 8320 -1610 8325 -1580
rect 8325 -1610 8355 -1580
rect 8355 -1610 8360 -1580
rect 8320 -1615 8360 -1610
rect 8320 -1645 8360 -1640
rect 8320 -1675 8325 -1645
rect 8325 -1675 8355 -1645
rect 8355 -1675 8360 -1645
rect 8320 -1680 8360 -1675
rect 8320 -1705 8360 -1700
rect 8320 -1735 8325 -1705
rect 8325 -1735 8355 -1705
rect 8355 -1735 8360 -1705
rect 8320 -1740 8360 -1735
rect 8320 -1770 8360 -1765
rect 8320 -1800 8325 -1770
rect 8325 -1800 8355 -1770
rect 8355 -1800 8360 -1770
rect 8320 -1805 8360 -1800
rect 8320 -1840 8360 -1835
rect 8320 -1870 8325 -1840
rect 8325 -1870 8355 -1840
rect 8355 -1870 8360 -1840
rect 8320 -1875 8360 -1870
rect 8320 -1910 8360 -1905
rect 8320 -1940 8325 -1910
rect 8325 -1940 8355 -1910
rect 8355 -1940 8360 -1910
rect 8320 -1945 8360 -1940
rect 8320 -1980 8360 -1975
rect 8320 -2010 8325 -1980
rect 8325 -2010 8355 -1980
rect 8355 -2010 8360 -1980
rect 8320 -2015 8360 -2010
rect 8320 -2045 8360 -2040
rect 8320 -2075 8325 -2045
rect 8325 -2075 8355 -2045
rect 8355 -2075 8360 -2045
rect 8320 -2080 8360 -2075
rect 8320 -2105 8360 -2100
rect 8320 -2135 8325 -2105
rect 8325 -2135 8355 -2105
rect 8355 -2135 8360 -2105
rect 8320 -2140 8360 -2135
rect 8320 -2170 8360 -2165
rect 8320 -2200 8325 -2170
rect 8325 -2200 8355 -2170
rect 8355 -2200 8360 -2170
rect 8320 -2205 8360 -2200
rect 8320 -2240 8360 -2235
rect 8320 -2270 8325 -2240
rect 8325 -2270 8355 -2240
rect 8355 -2270 8360 -2240
rect 8320 -2275 8360 -2270
rect 8320 -2310 8360 -2305
rect 8320 -2340 8325 -2310
rect 8325 -2340 8355 -2310
rect 8355 -2340 8360 -2310
rect 8320 -2345 8360 -2340
rect 8320 -2380 8360 -2375
rect 8320 -2410 8325 -2380
rect 8325 -2410 8355 -2380
rect 8355 -2410 8360 -2380
rect 8320 -2415 8360 -2410
rect 8320 -2445 8360 -2440
rect 8320 -2475 8325 -2445
rect 8325 -2475 8355 -2445
rect 8355 -2475 8360 -2445
rect 8320 -2480 8360 -2475
rect 8320 -2505 8360 -2500
rect 8320 -2535 8325 -2505
rect 8325 -2535 8355 -2505
rect 8355 -2535 8360 -2505
rect 8320 -2540 8360 -2535
rect 8320 -2570 8360 -2565
rect 8320 -2600 8325 -2570
rect 8325 -2600 8355 -2570
rect 8355 -2600 8360 -2570
rect 8320 -2605 8360 -2600
rect 8320 -2640 8360 -2635
rect 8320 -2670 8325 -2640
rect 8325 -2670 8355 -2640
rect 8355 -2670 8360 -2640
rect 8320 -2675 8360 -2670
rect 8320 -2710 8360 -2705
rect 8320 -2740 8325 -2710
rect 8325 -2740 8355 -2710
rect 8355 -2740 8360 -2710
rect 8320 -2745 8360 -2740
rect 8320 -2780 8360 -2775
rect 8320 -2810 8325 -2780
rect 8325 -2810 8355 -2780
rect 8355 -2810 8360 -2780
rect 8320 -2815 8360 -2810
rect 8320 -2845 8360 -2840
rect 8320 -2875 8325 -2845
rect 8325 -2875 8355 -2845
rect 8355 -2875 8360 -2845
rect 8320 -2880 8360 -2875
rect 8320 -2905 8360 -2900
rect 8320 -2935 8325 -2905
rect 8325 -2935 8355 -2905
rect 8355 -2935 8360 -2905
rect 8320 -2940 8360 -2935
rect 8320 -2970 8360 -2965
rect 8320 -3000 8325 -2970
rect 8325 -3000 8355 -2970
rect 8355 -3000 8360 -2970
rect 8320 -3005 8360 -3000
rect 8320 -3040 8360 -3035
rect 8320 -3070 8325 -3040
rect 8325 -3070 8355 -3040
rect 8355 -3070 8360 -3040
rect 8320 -3075 8360 -3070
rect 8320 -3110 8360 -3105
rect 8320 -3140 8325 -3110
rect 8325 -3140 8355 -3110
rect 8355 -3140 8360 -3110
rect 8320 -3145 8360 -3140
rect 8320 -3180 8360 -3175
rect 8320 -3210 8325 -3180
rect 8325 -3210 8355 -3180
rect 8355 -3210 8360 -3180
rect 8320 -3215 8360 -3210
rect 8320 -3245 8360 -3240
rect 8320 -3275 8325 -3245
rect 8325 -3275 8355 -3245
rect 8355 -3275 8360 -3245
rect 8320 -3280 8360 -3275
rect 8320 -3305 8360 -3300
rect 8320 -3335 8325 -3305
rect 8325 -3335 8355 -3305
rect 8355 -3335 8360 -3305
rect 8320 -3340 8360 -3335
rect 8320 -3370 8360 -3365
rect 8320 -3400 8325 -3370
rect 8325 -3400 8355 -3370
rect 8355 -3400 8360 -3370
rect 8320 -3405 8360 -3400
rect 8320 -3440 8360 -3435
rect 8320 -3470 8325 -3440
rect 8325 -3470 8355 -3440
rect 8355 -3470 8360 -3440
rect 8320 -3475 8360 -3470
rect 8320 -3510 8360 -3505
rect 8320 -3540 8325 -3510
rect 8325 -3540 8355 -3510
rect 8355 -3540 8360 -3510
rect 8320 -3545 8360 -3540
rect 8320 -3580 8360 -3575
rect 8320 -3610 8325 -3580
rect 8325 -3610 8355 -3580
rect 8355 -3610 8360 -3580
rect 8320 -3615 8360 -3610
rect 8320 -3645 8360 -3640
rect 8320 -3675 8325 -3645
rect 8325 -3675 8355 -3645
rect 8355 -3675 8360 -3645
rect 8320 -3680 8360 -3675
rect 8320 -3705 8360 -3700
rect 8320 -3735 8325 -3705
rect 8325 -3735 8355 -3705
rect 8355 -3735 8360 -3705
rect 8320 -3740 8360 -3735
rect 8320 -3770 8360 -3765
rect 8320 -3800 8325 -3770
rect 8325 -3800 8355 -3770
rect 8355 -3800 8360 -3770
rect 8320 -3805 8360 -3800
rect 8320 -3840 8360 -3835
rect 8320 -3870 8325 -3840
rect 8325 -3870 8355 -3840
rect 8355 -3870 8360 -3840
rect 8320 -3875 8360 -3870
rect 8320 -3910 8360 -3905
rect 8320 -3940 8325 -3910
rect 8325 -3940 8355 -3910
rect 8355 -3940 8360 -3910
rect 8320 -3945 8360 -3940
rect 8320 -3980 8360 -3975
rect 8320 -4010 8325 -3980
rect 8325 -4010 8355 -3980
rect 8355 -4010 8360 -3980
rect 8320 -4015 8360 -4010
rect 8320 -4045 8360 -4040
rect 8320 -4075 8325 -4045
rect 8325 -4075 8355 -4045
rect 8355 -4075 8360 -4045
rect 8320 -4080 8360 -4075
rect 8320 -4105 8360 -4100
rect 8320 -4135 8325 -4105
rect 8325 -4135 8355 -4105
rect 8355 -4135 8360 -4105
rect 8320 -4140 8360 -4135
rect 8320 -4170 8360 -4165
rect 8320 -4200 8325 -4170
rect 8325 -4200 8355 -4170
rect 8355 -4200 8360 -4170
rect 8320 -4205 8360 -4200
rect 8320 -4240 8360 -4235
rect 8320 -4270 8325 -4240
rect 8325 -4270 8355 -4240
rect 8355 -4270 8360 -4240
rect 8320 -4275 8360 -4270
rect 8320 -4310 8360 -4305
rect 8320 -4340 8325 -4310
rect 8325 -4340 8355 -4310
rect 8355 -4340 8360 -4310
rect 8320 -4345 8360 -4340
rect 8320 -4380 8360 -4375
rect 8320 -4410 8325 -4380
rect 8325 -4410 8355 -4380
rect 8355 -4410 8360 -4380
rect 8320 -4415 8360 -4410
rect 8320 -4445 8360 -4440
rect 8320 -4475 8325 -4445
rect 8325 -4475 8355 -4445
rect 8355 -4475 8360 -4445
rect 8320 -4480 8360 -4475
rect 8670 -1305 8710 -1300
rect 8670 -1335 8675 -1305
rect 8675 -1335 8705 -1305
rect 8705 -1335 8710 -1305
rect 8670 -1340 8710 -1335
rect 8670 -1370 8710 -1365
rect 8670 -1400 8675 -1370
rect 8675 -1400 8705 -1370
rect 8705 -1400 8710 -1370
rect 8670 -1405 8710 -1400
rect 8670 -1440 8710 -1435
rect 8670 -1470 8675 -1440
rect 8675 -1470 8705 -1440
rect 8705 -1470 8710 -1440
rect 8670 -1475 8710 -1470
rect 8670 -1510 8710 -1505
rect 8670 -1540 8675 -1510
rect 8675 -1540 8705 -1510
rect 8705 -1540 8710 -1510
rect 8670 -1545 8710 -1540
rect 8670 -1580 8710 -1575
rect 8670 -1610 8675 -1580
rect 8675 -1610 8705 -1580
rect 8705 -1610 8710 -1580
rect 8670 -1615 8710 -1610
rect 8670 -1645 8710 -1640
rect 8670 -1675 8675 -1645
rect 8675 -1675 8705 -1645
rect 8705 -1675 8710 -1645
rect 8670 -1680 8710 -1675
rect 8670 -1705 8710 -1700
rect 8670 -1735 8675 -1705
rect 8675 -1735 8705 -1705
rect 8705 -1735 8710 -1705
rect 8670 -1740 8710 -1735
rect 8670 -1770 8710 -1765
rect 8670 -1800 8675 -1770
rect 8675 -1800 8705 -1770
rect 8705 -1800 8710 -1770
rect 8670 -1805 8710 -1800
rect 8670 -1840 8710 -1835
rect 8670 -1870 8675 -1840
rect 8675 -1870 8705 -1840
rect 8705 -1870 8710 -1840
rect 8670 -1875 8710 -1870
rect 8670 -1910 8710 -1905
rect 8670 -1940 8675 -1910
rect 8675 -1940 8705 -1910
rect 8705 -1940 8710 -1910
rect 8670 -1945 8710 -1940
rect 8670 -1980 8710 -1975
rect 8670 -2010 8675 -1980
rect 8675 -2010 8705 -1980
rect 8705 -2010 8710 -1980
rect 8670 -2015 8710 -2010
rect 8670 -2045 8710 -2040
rect 8670 -2075 8675 -2045
rect 8675 -2075 8705 -2045
rect 8705 -2075 8710 -2045
rect 8670 -2080 8710 -2075
rect 8670 -2105 8710 -2100
rect 8670 -2135 8675 -2105
rect 8675 -2135 8705 -2105
rect 8705 -2135 8710 -2105
rect 8670 -2140 8710 -2135
rect 8670 -2170 8710 -2165
rect 8670 -2200 8675 -2170
rect 8675 -2200 8705 -2170
rect 8705 -2200 8710 -2170
rect 8670 -2205 8710 -2200
rect 8670 -2240 8710 -2235
rect 8670 -2270 8675 -2240
rect 8675 -2270 8705 -2240
rect 8705 -2270 8710 -2240
rect 8670 -2275 8710 -2270
rect 8670 -2310 8710 -2305
rect 8670 -2340 8675 -2310
rect 8675 -2340 8705 -2310
rect 8705 -2340 8710 -2310
rect 8670 -2345 8710 -2340
rect 8670 -2380 8710 -2375
rect 8670 -2410 8675 -2380
rect 8675 -2410 8705 -2380
rect 8705 -2410 8710 -2380
rect 8670 -2415 8710 -2410
rect 8670 -2445 8710 -2440
rect 8670 -2475 8675 -2445
rect 8675 -2475 8705 -2445
rect 8705 -2475 8710 -2445
rect 8670 -2480 8710 -2475
rect 8670 -2505 8710 -2500
rect 8670 -2535 8675 -2505
rect 8675 -2535 8705 -2505
rect 8705 -2535 8710 -2505
rect 8670 -2540 8710 -2535
rect 8670 -2570 8710 -2565
rect 8670 -2600 8675 -2570
rect 8675 -2600 8705 -2570
rect 8705 -2600 8710 -2570
rect 8670 -2605 8710 -2600
rect 8670 -2640 8710 -2635
rect 8670 -2670 8675 -2640
rect 8675 -2670 8705 -2640
rect 8705 -2670 8710 -2640
rect 8670 -2675 8710 -2670
rect 8670 -2710 8710 -2705
rect 8670 -2740 8675 -2710
rect 8675 -2740 8705 -2710
rect 8705 -2740 8710 -2710
rect 8670 -2745 8710 -2740
rect 8670 -2780 8710 -2775
rect 8670 -2810 8675 -2780
rect 8675 -2810 8705 -2780
rect 8705 -2810 8710 -2780
rect 8670 -2815 8710 -2810
rect 8670 -2845 8710 -2840
rect 8670 -2875 8675 -2845
rect 8675 -2875 8705 -2845
rect 8705 -2875 8710 -2845
rect 8670 -2880 8710 -2875
rect 8670 -2905 8710 -2900
rect 8670 -2935 8675 -2905
rect 8675 -2935 8705 -2905
rect 8705 -2935 8710 -2905
rect 8670 -2940 8710 -2935
rect 8670 -2970 8710 -2965
rect 8670 -3000 8675 -2970
rect 8675 -3000 8705 -2970
rect 8705 -3000 8710 -2970
rect 8670 -3005 8710 -3000
rect 8670 -3040 8710 -3035
rect 8670 -3070 8675 -3040
rect 8675 -3070 8705 -3040
rect 8705 -3070 8710 -3040
rect 8670 -3075 8710 -3070
rect 8670 -3110 8710 -3105
rect 8670 -3140 8675 -3110
rect 8675 -3140 8705 -3110
rect 8705 -3140 8710 -3110
rect 8670 -3145 8710 -3140
rect 8670 -3180 8710 -3175
rect 8670 -3210 8675 -3180
rect 8675 -3210 8705 -3180
rect 8705 -3210 8710 -3180
rect 8670 -3215 8710 -3210
rect 8670 -3245 8710 -3240
rect 8670 -3275 8675 -3245
rect 8675 -3275 8705 -3245
rect 8705 -3275 8710 -3245
rect 8670 -3280 8710 -3275
rect 8670 -3305 8710 -3300
rect 8670 -3335 8675 -3305
rect 8675 -3335 8705 -3305
rect 8705 -3335 8710 -3305
rect 8670 -3340 8710 -3335
rect 8670 -3370 8710 -3365
rect 8670 -3400 8675 -3370
rect 8675 -3400 8705 -3370
rect 8705 -3400 8710 -3370
rect 8670 -3405 8710 -3400
rect 8670 -3440 8710 -3435
rect 8670 -3470 8675 -3440
rect 8675 -3470 8705 -3440
rect 8705 -3470 8710 -3440
rect 8670 -3475 8710 -3470
rect 8670 -3510 8710 -3505
rect 8670 -3540 8675 -3510
rect 8675 -3540 8705 -3510
rect 8705 -3540 8710 -3510
rect 8670 -3545 8710 -3540
rect 8670 -3580 8710 -3575
rect 8670 -3610 8675 -3580
rect 8675 -3610 8705 -3580
rect 8705 -3610 8710 -3580
rect 8670 -3615 8710 -3610
rect 8670 -3645 8710 -3640
rect 8670 -3675 8675 -3645
rect 8675 -3675 8705 -3645
rect 8705 -3675 8710 -3645
rect 8670 -3680 8710 -3675
rect 8670 -3705 8710 -3700
rect 8670 -3735 8675 -3705
rect 8675 -3735 8705 -3705
rect 8705 -3735 8710 -3705
rect 8670 -3740 8710 -3735
rect 8670 -3770 8710 -3765
rect 8670 -3800 8675 -3770
rect 8675 -3800 8705 -3770
rect 8705 -3800 8710 -3770
rect 8670 -3805 8710 -3800
rect 8670 -3840 8710 -3835
rect 8670 -3870 8675 -3840
rect 8675 -3870 8705 -3840
rect 8705 -3870 8710 -3840
rect 8670 -3875 8710 -3870
rect 8670 -3910 8710 -3905
rect 8670 -3940 8675 -3910
rect 8675 -3940 8705 -3910
rect 8705 -3940 8710 -3910
rect 8670 -3945 8710 -3940
rect 8670 -3980 8710 -3975
rect 8670 -4010 8675 -3980
rect 8675 -4010 8705 -3980
rect 8705 -4010 8710 -3980
rect 8670 -4015 8710 -4010
rect 8670 -4045 8710 -4040
rect 8670 -4075 8675 -4045
rect 8675 -4075 8705 -4045
rect 8705 -4075 8710 -4045
rect 8670 -4080 8710 -4075
rect 8670 -4105 8710 -4100
rect 8670 -4135 8675 -4105
rect 8675 -4135 8705 -4105
rect 8705 -4135 8710 -4105
rect 8670 -4140 8710 -4135
rect 8670 -4170 8710 -4165
rect 8670 -4200 8675 -4170
rect 8675 -4200 8705 -4170
rect 8705 -4200 8710 -4170
rect 8670 -4205 8710 -4200
rect 8670 -4240 8710 -4235
rect 8670 -4270 8675 -4240
rect 8675 -4270 8705 -4240
rect 8705 -4270 8710 -4240
rect 8670 -4275 8710 -4270
rect 8670 -4310 8710 -4305
rect 8670 -4340 8675 -4310
rect 8675 -4340 8705 -4310
rect 8705 -4340 8710 -4310
rect 8670 -4345 8710 -4340
rect 8670 -4380 8710 -4375
rect 8670 -4410 8675 -4380
rect 8675 -4410 8705 -4380
rect 8705 -4410 8710 -4380
rect 8670 -4415 8710 -4410
rect 8670 -4445 8710 -4440
rect 8670 -4475 8675 -4445
rect 8675 -4475 8705 -4445
rect 8705 -4475 8710 -4445
rect 8670 -4480 8710 -4475
rect 14825 -1375 14875 -1325
rect 14920 -1375 14970 -1325
rect 15015 -1375 15065 -1325
rect 15115 -1375 15165 -1325
rect 15215 -1375 15265 -1325
rect 15315 -1375 15365 -1325
rect 15410 -1375 15460 -1325
rect 15505 -1375 15555 -1325
rect 15625 -1375 15675 -1325
rect 15720 -1375 15770 -1325
rect 15815 -1375 15865 -1325
rect 15915 -1375 15965 -1325
rect 16015 -1375 16065 -1325
rect 16115 -1375 16165 -1325
rect 16210 -1375 16260 -1325
rect 16305 -1375 16355 -1325
rect 16425 -1375 16475 -1325
rect 16520 -1375 16570 -1325
rect 16615 -1375 16665 -1325
rect 16715 -1375 16765 -1325
rect 16815 -1375 16865 -1325
rect 16915 -1375 16965 -1325
rect 17010 -1375 17060 -1325
rect 17105 -1375 17155 -1325
rect 17225 -1375 17275 -1325
rect 17320 -1375 17370 -1325
rect 17415 -1375 17465 -1325
rect 17515 -1375 17565 -1325
rect 17615 -1375 17665 -1325
rect 17715 -1375 17765 -1325
rect 17810 -1375 17860 -1325
rect 17905 -1375 17955 -1325
rect 14825 -1465 14875 -1415
rect 14920 -1465 14970 -1415
rect 15015 -1465 15065 -1415
rect 15115 -1465 15165 -1415
rect 15215 -1465 15265 -1415
rect 15315 -1465 15365 -1415
rect 15410 -1465 15460 -1415
rect 15505 -1465 15555 -1415
rect 15625 -1465 15675 -1415
rect 15720 -1465 15770 -1415
rect 15815 -1465 15865 -1415
rect 15915 -1465 15965 -1415
rect 16015 -1465 16065 -1415
rect 16115 -1465 16165 -1415
rect 16210 -1465 16260 -1415
rect 16305 -1465 16355 -1415
rect 16425 -1465 16475 -1415
rect 16520 -1465 16570 -1415
rect 16615 -1465 16665 -1415
rect 16715 -1465 16765 -1415
rect 16815 -1465 16865 -1415
rect 16915 -1465 16965 -1415
rect 17010 -1465 17060 -1415
rect 17105 -1465 17155 -1415
rect 17225 -1465 17275 -1415
rect 17320 -1465 17370 -1415
rect 17415 -1465 17465 -1415
rect 17515 -1465 17565 -1415
rect 17615 -1465 17665 -1415
rect 17715 -1465 17765 -1415
rect 17810 -1465 17860 -1415
rect 17905 -1465 17955 -1415
rect 14825 -1565 14875 -1515
rect 14920 -1565 14970 -1515
rect 15015 -1565 15065 -1515
rect 15115 -1565 15165 -1515
rect 15215 -1565 15265 -1515
rect 15315 -1565 15365 -1515
rect 15410 -1565 15460 -1515
rect 15505 -1565 15555 -1515
rect 15625 -1565 15675 -1515
rect 15720 -1565 15770 -1515
rect 15815 -1565 15865 -1515
rect 15915 -1565 15965 -1515
rect 16015 -1565 16065 -1515
rect 16115 -1565 16165 -1515
rect 16210 -1565 16260 -1515
rect 16305 -1565 16355 -1515
rect 16425 -1565 16475 -1515
rect 16520 -1565 16570 -1515
rect 16615 -1565 16665 -1515
rect 16715 -1565 16765 -1515
rect 16815 -1565 16865 -1515
rect 16915 -1565 16965 -1515
rect 17010 -1565 17060 -1515
rect 17105 -1565 17155 -1515
rect 17225 -1565 17275 -1515
rect 17320 -1565 17370 -1515
rect 17415 -1565 17465 -1515
rect 17515 -1565 17565 -1515
rect 17615 -1565 17665 -1515
rect 17715 -1565 17765 -1515
rect 17810 -1565 17860 -1515
rect 17905 -1565 17955 -1515
rect 14825 -1655 14875 -1605
rect 14920 -1655 14970 -1605
rect 15015 -1655 15065 -1605
rect 15115 -1655 15165 -1605
rect 15215 -1655 15265 -1605
rect 15315 -1655 15365 -1605
rect 15410 -1655 15460 -1605
rect 15505 -1655 15555 -1605
rect 15625 -1655 15675 -1605
rect 15720 -1655 15770 -1605
rect 15815 -1655 15865 -1605
rect 15915 -1655 15965 -1605
rect 16015 -1655 16065 -1605
rect 16115 -1655 16165 -1605
rect 16210 -1655 16260 -1605
rect 16305 -1655 16355 -1605
rect 16425 -1655 16475 -1605
rect 16520 -1655 16570 -1605
rect 16615 -1655 16665 -1605
rect 16715 -1655 16765 -1605
rect 16815 -1655 16865 -1605
rect 16915 -1655 16965 -1605
rect 17010 -1655 17060 -1605
rect 17105 -1655 17155 -1605
rect 17225 -1655 17275 -1605
rect 17320 -1655 17370 -1605
rect 17415 -1655 17465 -1605
rect 17515 -1655 17565 -1605
rect 17615 -1655 17665 -1605
rect 17715 -1655 17765 -1605
rect 17810 -1655 17860 -1605
rect 17905 -1655 17955 -1605
rect 14825 -1775 14875 -1725
rect 14920 -1775 14970 -1725
rect 15015 -1775 15065 -1725
rect 15115 -1775 15165 -1725
rect 15215 -1775 15265 -1725
rect 15315 -1775 15365 -1725
rect 15410 -1775 15460 -1725
rect 15505 -1775 15555 -1725
rect 15625 -1775 15675 -1725
rect 15720 -1775 15770 -1725
rect 15815 -1775 15865 -1725
rect 15915 -1775 15965 -1725
rect 16015 -1775 16065 -1725
rect 16115 -1775 16165 -1725
rect 16210 -1775 16260 -1725
rect 16305 -1775 16355 -1725
rect 16425 -1775 16475 -1725
rect 16520 -1775 16570 -1725
rect 16615 -1775 16665 -1725
rect 16715 -1775 16765 -1725
rect 16815 -1775 16865 -1725
rect 16915 -1775 16965 -1725
rect 17010 -1775 17060 -1725
rect 17105 -1775 17155 -1725
rect 17225 -1775 17275 -1725
rect 17320 -1775 17370 -1725
rect 17415 -1775 17465 -1725
rect 17515 -1775 17565 -1725
rect 17615 -1775 17665 -1725
rect 17715 -1775 17765 -1725
rect 17810 -1775 17860 -1725
rect 17905 -1775 17955 -1725
rect 14825 -1865 14875 -1815
rect 14920 -1865 14970 -1815
rect 15015 -1865 15065 -1815
rect 15115 -1865 15165 -1815
rect 15215 -1865 15265 -1815
rect 15315 -1865 15365 -1815
rect 15410 -1865 15460 -1815
rect 15505 -1865 15555 -1815
rect 15625 -1865 15675 -1815
rect 15720 -1865 15770 -1815
rect 15815 -1865 15865 -1815
rect 15915 -1865 15965 -1815
rect 16015 -1865 16065 -1815
rect 16115 -1865 16165 -1815
rect 16210 -1865 16260 -1815
rect 16305 -1865 16355 -1815
rect 16425 -1865 16475 -1815
rect 16520 -1865 16570 -1815
rect 16615 -1865 16665 -1815
rect 16715 -1865 16765 -1815
rect 16815 -1865 16865 -1815
rect 16915 -1865 16965 -1815
rect 17010 -1865 17060 -1815
rect 17105 -1865 17155 -1815
rect 17225 -1865 17275 -1815
rect 17320 -1865 17370 -1815
rect 17415 -1865 17465 -1815
rect 17515 -1865 17565 -1815
rect 17615 -1865 17665 -1815
rect 17715 -1865 17765 -1815
rect 17810 -1865 17860 -1815
rect 17905 -1865 17955 -1815
rect 14825 -1965 14875 -1915
rect 14920 -1965 14970 -1915
rect 15015 -1965 15065 -1915
rect 15115 -1965 15165 -1915
rect 15215 -1965 15265 -1915
rect 15315 -1965 15365 -1915
rect 15410 -1965 15460 -1915
rect 15505 -1965 15555 -1915
rect 15625 -1965 15675 -1915
rect 15720 -1965 15770 -1915
rect 15815 -1965 15865 -1915
rect 15915 -1965 15965 -1915
rect 16015 -1965 16065 -1915
rect 16115 -1965 16165 -1915
rect 16210 -1965 16260 -1915
rect 16305 -1965 16355 -1915
rect 16425 -1965 16475 -1915
rect 16520 -1965 16570 -1915
rect 16615 -1965 16665 -1915
rect 16715 -1965 16765 -1915
rect 16815 -1965 16865 -1915
rect 16915 -1965 16965 -1915
rect 17010 -1965 17060 -1915
rect 17105 -1965 17155 -1915
rect 17225 -1965 17275 -1915
rect 17320 -1965 17370 -1915
rect 17415 -1965 17465 -1915
rect 17515 -1965 17565 -1915
rect 17615 -1965 17665 -1915
rect 17715 -1965 17765 -1915
rect 17810 -1965 17860 -1915
rect 17905 -1965 17955 -1915
rect 14825 -2055 14875 -2005
rect 14920 -2055 14970 -2005
rect 15015 -2055 15065 -2005
rect 15115 -2055 15165 -2005
rect 15215 -2055 15265 -2005
rect 15315 -2055 15365 -2005
rect 15410 -2055 15460 -2005
rect 15505 -2055 15555 -2005
rect 15625 -2055 15675 -2005
rect 15720 -2055 15770 -2005
rect 15815 -2055 15865 -2005
rect 15915 -2055 15965 -2005
rect 16015 -2055 16065 -2005
rect 16115 -2055 16165 -2005
rect 16210 -2055 16260 -2005
rect 16305 -2055 16355 -2005
rect 16425 -2055 16475 -2005
rect 16520 -2055 16570 -2005
rect 16615 -2055 16665 -2005
rect 16715 -2055 16765 -2005
rect 16815 -2055 16865 -2005
rect 16915 -2055 16965 -2005
rect 17010 -2055 17060 -2005
rect 17105 -2055 17155 -2005
rect 17225 -2055 17275 -2005
rect 17320 -2055 17370 -2005
rect 17415 -2055 17465 -2005
rect 17515 -2055 17565 -2005
rect 17615 -2055 17665 -2005
rect 17715 -2055 17765 -2005
rect 17810 -2055 17860 -2005
rect 17905 -2055 17955 -2005
rect 14825 -2175 14875 -2125
rect 14920 -2175 14970 -2125
rect 15015 -2175 15065 -2125
rect 15115 -2175 15165 -2125
rect 15215 -2175 15265 -2125
rect 15315 -2175 15365 -2125
rect 15410 -2175 15460 -2125
rect 15505 -2175 15555 -2125
rect 15625 -2175 15675 -2125
rect 15720 -2175 15770 -2125
rect 15815 -2175 15865 -2125
rect 15915 -2175 15965 -2125
rect 16015 -2175 16065 -2125
rect 16115 -2175 16165 -2125
rect 16210 -2175 16260 -2125
rect 16305 -2175 16355 -2125
rect 16425 -2175 16475 -2125
rect 16520 -2175 16570 -2125
rect 16615 -2175 16665 -2125
rect 16715 -2175 16765 -2125
rect 16815 -2175 16865 -2125
rect 16915 -2175 16965 -2125
rect 17010 -2175 17060 -2125
rect 17105 -2175 17155 -2125
rect 17225 -2175 17275 -2125
rect 17320 -2175 17370 -2125
rect 17415 -2175 17465 -2125
rect 17515 -2175 17565 -2125
rect 17615 -2175 17665 -2125
rect 17715 -2175 17765 -2125
rect 17810 -2175 17860 -2125
rect 17905 -2175 17955 -2125
rect 14825 -2265 14875 -2215
rect 14920 -2265 14970 -2215
rect 15015 -2265 15065 -2215
rect 15115 -2265 15165 -2215
rect 15215 -2265 15265 -2215
rect 15315 -2265 15365 -2215
rect 15410 -2265 15460 -2215
rect 15505 -2265 15555 -2215
rect 15625 -2265 15675 -2215
rect 15720 -2265 15770 -2215
rect 15815 -2265 15865 -2215
rect 15915 -2265 15965 -2215
rect 16015 -2265 16065 -2215
rect 16115 -2265 16165 -2215
rect 16210 -2265 16260 -2215
rect 16305 -2265 16355 -2215
rect 16425 -2265 16475 -2215
rect 16520 -2265 16570 -2215
rect 16615 -2265 16665 -2215
rect 16715 -2265 16765 -2215
rect 16815 -2265 16865 -2215
rect 16915 -2265 16965 -2215
rect 17010 -2265 17060 -2215
rect 17105 -2265 17155 -2215
rect 17225 -2265 17275 -2215
rect 17320 -2265 17370 -2215
rect 17415 -2265 17465 -2215
rect 17515 -2265 17565 -2215
rect 17615 -2265 17665 -2215
rect 17715 -2265 17765 -2215
rect 17810 -2265 17860 -2215
rect 17905 -2265 17955 -2215
rect 14825 -2365 14875 -2315
rect 14920 -2365 14970 -2315
rect 15015 -2365 15065 -2315
rect 15115 -2365 15165 -2315
rect 15215 -2365 15265 -2315
rect 15315 -2365 15365 -2315
rect 15410 -2365 15460 -2315
rect 15505 -2365 15555 -2315
rect 15625 -2365 15675 -2315
rect 15720 -2365 15770 -2315
rect 15815 -2365 15865 -2315
rect 15915 -2365 15965 -2315
rect 16015 -2365 16065 -2315
rect 16115 -2365 16165 -2315
rect 16210 -2365 16260 -2315
rect 16305 -2365 16355 -2315
rect 16425 -2365 16475 -2315
rect 16520 -2365 16570 -2315
rect 16615 -2365 16665 -2315
rect 16715 -2365 16765 -2315
rect 16815 -2365 16865 -2315
rect 16915 -2365 16965 -2315
rect 17010 -2365 17060 -2315
rect 17105 -2365 17155 -2315
rect 17225 -2365 17275 -2315
rect 17320 -2365 17370 -2315
rect 17415 -2365 17465 -2315
rect 17515 -2365 17565 -2315
rect 17615 -2365 17665 -2315
rect 17715 -2365 17765 -2315
rect 17810 -2365 17860 -2315
rect 17905 -2365 17955 -2315
rect 14825 -2455 14875 -2405
rect 14920 -2455 14970 -2405
rect 15015 -2455 15065 -2405
rect 15115 -2455 15165 -2405
rect 15215 -2455 15265 -2405
rect 15315 -2455 15365 -2405
rect 15410 -2455 15460 -2405
rect 15505 -2455 15555 -2405
rect 15625 -2455 15675 -2405
rect 15720 -2455 15770 -2405
rect 15815 -2455 15865 -2405
rect 15915 -2455 15965 -2405
rect 16015 -2455 16065 -2405
rect 16115 -2455 16165 -2405
rect 16210 -2455 16260 -2405
rect 16305 -2455 16355 -2405
rect 16425 -2455 16475 -2405
rect 16520 -2455 16570 -2405
rect 16615 -2455 16665 -2405
rect 16715 -2455 16765 -2405
rect 16815 -2455 16865 -2405
rect 16915 -2455 16965 -2405
rect 17010 -2455 17060 -2405
rect 17105 -2455 17155 -2405
rect 17225 -2455 17275 -2405
rect 17320 -2455 17370 -2405
rect 17415 -2455 17465 -2405
rect 17515 -2455 17565 -2405
rect 17615 -2455 17665 -2405
rect 17715 -2455 17765 -2405
rect 17810 -2455 17860 -2405
rect 17905 -2455 17955 -2405
rect 14825 -2575 14875 -2525
rect 14920 -2575 14970 -2525
rect 15015 -2575 15065 -2525
rect 15115 -2575 15165 -2525
rect 15215 -2575 15265 -2525
rect 15315 -2575 15365 -2525
rect 15410 -2575 15460 -2525
rect 15505 -2575 15555 -2525
rect 15625 -2575 15675 -2525
rect 15720 -2575 15770 -2525
rect 15815 -2575 15865 -2525
rect 15915 -2575 15965 -2525
rect 16015 -2575 16065 -2525
rect 16115 -2575 16165 -2525
rect 16210 -2575 16260 -2525
rect 16305 -2575 16355 -2525
rect 16425 -2575 16475 -2525
rect 16520 -2575 16570 -2525
rect 16615 -2575 16665 -2525
rect 16715 -2575 16765 -2525
rect 16815 -2575 16865 -2525
rect 16915 -2575 16965 -2525
rect 17010 -2575 17060 -2525
rect 17105 -2575 17155 -2525
rect 17225 -2575 17275 -2525
rect 17320 -2575 17370 -2525
rect 17415 -2575 17465 -2525
rect 17515 -2575 17565 -2525
rect 17615 -2575 17665 -2525
rect 17715 -2575 17765 -2525
rect 17810 -2575 17860 -2525
rect 17905 -2575 17955 -2525
rect 14825 -2665 14875 -2615
rect 14920 -2665 14970 -2615
rect 15015 -2665 15065 -2615
rect 15115 -2665 15165 -2615
rect 15215 -2665 15265 -2615
rect 15315 -2665 15365 -2615
rect 15410 -2665 15460 -2615
rect 15505 -2665 15555 -2615
rect 15625 -2665 15675 -2615
rect 15720 -2665 15770 -2615
rect 15815 -2665 15865 -2615
rect 15915 -2665 15965 -2615
rect 16015 -2665 16065 -2615
rect 16115 -2665 16165 -2615
rect 16210 -2665 16260 -2615
rect 16305 -2665 16355 -2615
rect 16425 -2665 16475 -2615
rect 16520 -2665 16570 -2615
rect 16615 -2665 16665 -2615
rect 16715 -2665 16765 -2615
rect 16815 -2665 16865 -2615
rect 16915 -2665 16965 -2615
rect 17010 -2665 17060 -2615
rect 17105 -2665 17155 -2615
rect 17225 -2665 17275 -2615
rect 17320 -2665 17370 -2615
rect 17415 -2665 17465 -2615
rect 17515 -2665 17565 -2615
rect 17615 -2665 17665 -2615
rect 17715 -2665 17765 -2615
rect 17810 -2665 17860 -2615
rect 17905 -2665 17955 -2615
rect 14825 -2765 14875 -2715
rect 14920 -2765 14970 -2715
rect 15015 -2765 15065 -2715
rect 15115 -2765 15165 -2715
rect 15215 -2765 15265 -2715
rect 15315 -2765 15365 -2715
rect 15410 -2765 15460 -2715
rect 15505 -2765 15555 -2715
rect 15625 -2765 15675 -2715
rect 15720 -2765 15770 -2715
rect 15815 -2765 15865 -2715
rect 15915 -2765 15965 -2715
rect 16015 -2765 16065 -2715
rect 16115 -2765 16165 -2715
rect 16210 -2765 16260 -2715
rect 16305 -2765 16355 -2715
rect 16425 -2765 16475 -2715
rect 16520 -2765 16570 -2715
rect 16615 -2765 16665 -2715
rect 16715 -2765 16765 -2715
rect 16815 -2765 16865 -2715
rect 16915 -2765 16965 -2715
rect 17010 -2765 17060 -2715
rect 17105 -2765 17155 -2715
rect 17225 -2765 17275 -2715
rect 17320 -2765 17370 -2715
rect 17415 -2765 17465 -2715
rect 17515 -2765 17565 -2715
rect 17615 -2765 17665 -2715
rect 17715 -2765 17765 -2715
rect 17810 -2765 17860 -2715
rect 17905 -2765 17955 -2715
rect 14825 -2855 14875 -2805
rect 14920 -2855 14970 -2805
rect 15015 -2855 15065 -2805
rect 15115 -2855 15165 -2805
rect 15215 -2855 15265 -2805
rect 15315 -2855 15365 -2805
rect 15410 -2855 15460 -2805
rect 15505 -2855 15555 -2805
rect 15625 -2855 15675 -2805
rect 15720 -2855 15770 -2805
rect 15815 -2855 15865 -2805
rect 15915 -2855 15965 -2805
rect 16015 -2855 16065 -2805
rect 16115 -2855 16165 -2805
rect 16210 -2855 16260 -2805
rect 16305 -2855 16355 -2805
rect 16425 -2855 16475 -2805
rect 16520 -2855 16570 -2805
rect 16615 -2855 16665 -2805
rect 16715 -2855 16765 -2805
rect 16815 -2855 16865 -2805
rect 16915 -2855 16965 -2805
rect 17010 -2855 17060 -2805
rect 17105 -2855 17155 -2805
rect 17225 -2855 17275 -2805
rect 17320 -2855 17370 -2805
rect 17415 -2855 17465 -2805
rect 17515 -2855 17565 -2805
rect 17615 -2855 17665 -2805
rect 17715 -2855 17765 -2805
rect 17810 -2855 17860 -2805
rect 17905 -2855 17955 -2805
rect 14825 -2975 14875 -2925
rect 14920 -2975 14970 -2925
rect 15015 -2975 15065 -2925
rect 15115 -2975 15165 -2925
rect 15215 -2975 15265 -2925
rect 15315 -2975 15365 -2925
rect 15410 -2975 15460 -2925
rect 15505 -2975 15555 -2925
rect 15625 -2975 15675 -2925
rect 15720 -2975 15770 -2925
rect 15815 -2975 15865 -2925
rect 15915 -2975 15965 -2925
rect 16015 -2975 16065 -2925
rect 16115 -2975 16165 -2925
rect 16210 -2975 16260 -2925
rect 16305 -2975 16355 -2925
rect 16425 -2975 16475 -2925
rect 16520 -2975 16570 -2925
rect 16615 -2975 16665 -2925
rect 16715 -2975 16765 -2925
rect 16815 -2975 16865 -2925
rect 16915 -2975 16965 -2925
rect 17010 -2975 17060 -2925
rect 17105 -2975 17155 -2925
rect 17225 -2975 17275 -2925
rect 17320 -2975 17370 -2925
rect 17415 -2975 17465 -2925
rect 17515 -2975 17565 -2925
rect 17615 -2975 17665 -2925
rect 17715 -2975 17765 -2925
rect 17810 -2975 17860 -2925
rect 17905 -2975 17955 -2925
rect 14825 -3065 14875 -3015
rect 14920 -3065 14970 -3015
rect 15015 -3065 15065 -3015
rect 15115 -3065 15165 -3015
rect 15215 -3065 15265 -3015
rect 15315 -3065 15365 -3015
rect 15410 -3065 15460 -3015
rect 15505 -3065 15555 -3015
rect 15625 -3065 15675 -3015
rect 15720 -3065 15770 -3015
rect 15815 -3065 15865 -3015
rect 15915 -3065 15965 -3015
rect 16015 -3065 16065 -3015
rect 16115 -3065 16165 -3015
rect 16210 -3065 16260 -3015
rect 16305 -3065 16355 -3015
rect 16425 -3065 16475 -3015
rect 16520 -3065 16570 -3015
rect 16615 -3065 16665 -3015
rect 16715 -3065 16765 -3015
rect 16815 -3065 16865 -3015
rect 16915 -3065 16965 -3015
rect 17010 -3065 17060 -3015
rect 17105 -3065 17155 -3015
rect 17225 -3065 17275 -3015
rect 17320 -3065 17370 -3015
rect 17415 -3065 17465 -3015
rect 17515 -3065 17565 -3015
rect 17615 -3065 17665 -3015
rect 17715 -3065 17765 -3015
rect 17810 -3065 17860 -3015
rect 17905 -3065 17955 -3015
rect 14825 -3165 14875 -3115
rect 14920 -3165 14970 -3115
rect 15015 -3165 15065 -3115
rect 15115 -3165 15165 -3115
rect 15215 -3165 15265 -3115
rect 15315 -3165 15365 -3115
rect 15410 -3165 15460 -3115
rect 15505 -3165 15555 -3115
rect 15625 -3165 15675 -3115
rect 15720 -3165 15770 -3115
rect 15815 -3165 15865 -3115
rect 15915 -3165 15965 -3115
rect 16015 -3165 16065 -3115
rect 16115 -3165 16165 -3115
rect 16210 -3165 16260 -3115
rect 16305 -3165 16355 -3115
rect 16425 -3165 16475 -3115
rect 16520 -3165 16570 -3115
rect 16615 -3165 16665 -3115
rect 16715 -3165 16765 -3115
rect 16815 -3165 16865 -3115
rect 16915 -3165 16965 -3115
rect 17010 -3165 17060 -3115
rect 17105 -3165 17155 -3115
rect 17225 -3165 17275 -3115
rect 17320 -3165 17370 -3115
rect 17415 -3165 17465 -3115
rect 17515 -3165 17565 -3115
rect 17615 -3165 17665 -3115
rect 17715 -3165 17765 -3115
rect 17810 -3165 17860 -3115
rect 17905 -3165 17955 -3115
rect 14825 -3255 14875 -3205
rect 14920 -3255 14970 -3205
rect 15015 -3255 15065 -3205
rect 15115 -3255 15165 -3205
rect 15215 -3255 15265 -3205
rect 15315 -3255 15365 -3205
rect 15410 -3255 15460 -3205
rect 15505 -3255 15555 -3205
rect 15625 -3255 15675 -3205
rect 15720 -3255 15770 -3205
rect 15815 -3255 15865 -3205
rect 15915 -3255 15965 -3205
rect 16015 -3255 16065 -3205
rect 16115 -3255 16165 -3205
rect 16210 -3255 16260 -3205
rect 16305 -3255 16355 -3205
rect 16425 -3255 16475 -3205
rect 16520 -3255 16570 -3205
rect 16615 -3255 16665 -3205
rect 16715 -3255 16765 -3205
rect 16815 -3255 16865 -3205
rect 16915 -3255 16965 -3205
rect 17010 -3255 17060 -3205
rect 17105 -3255 17155 -3205
rect 17225 -3255 17275 -3205
rect 17320 -3255 17370 -3205
rect 17415 -3255 17465 -3205
rect 17515 -3255 17565 -3205
rect 17615 -3255 17665 -3205
rect 17715 -3255 17765 -3205
rect 17810 -3255 17860 -3205
rect 17905 -3255 17955 -3205
rect 14825 -3375 14875 -3325
rect 14920 -3375 14970 -3325
rect 15015 -3375 15065 -3325
rect 15115 -3375 15165 -3325
rect 15215 -3375 15265 -3325
rect 15315 -3375 15365 -3325
rect 15410 -3375 15460 -3325
rect 15505 -3375 15555 -3325
rect 15625 -3375 15675 -3325
rect 15720 -3375 15770 -3325
rect 15815 -3375 15865 -3325
rect 15915 -3375 15965 -3325
rect 16015 -3375 16065 -3325
rect 16115 -3375 16165 -3325
rect 16210 -3375 16260 -3325
rect 16305 -3375 16355 -3325
rect 16425 -3375 16475 -3325
rect 16520 -3375 16570 -3325
rect 16615 -3375 16665 -3325
rect 16715 -3375 16765 -3325
rect 16815 -3375 16865 -3325
rect 16915 -3375 16965 -3325
rect 17010 -3375 17060 -3325
rect 17105 -3375 17155 -3325
rect 17225 -3375 17275 -3325
rect 17320 -3375 17370 -3325
rect 17415 -3375 17465 -3325
rect 17515 -3375 17565 -3325
rect 17615 -3375 17665 -3325
rect 17715 -3375 17765 -3325
rect 17810 -3375 17860 -3325
rect 17905 -3375 17955 -3325
rect 14825 -3465 14875 -3415
rect 14920 -3465 14970 -3415
rect 15015 -3465 15065 -3415
rect 15115 -3465 15165 -3415
rect 15215 -3465 15265 -3415
rect 15315 -3465 15365 -3415
rect 15410 -3465 15460 -3415
rect 15505 -3465 15555 -3415
rect 15625 -3465 15675 -3415
rect 15720 -3465 15770 -3415
rect 15815 -3465 15865 -3415
rect 15915 -3465 15965 -3415
rect 16015 -3465 16065 -3415
rect 16115 -3465 16165 -3415
rect 16210 -3465 16260 -3415
rect 16305 -3465 16355 -3415
rect 16425 -3465 16475 -3415
rect 16520 -3465 16570 -3415
rect 16615 -3465 16665 -3415
rect 16715 -3465 16765 -3415
rect 16815 -3465 16865 -3415
rect 16915 -3465 16965 -3415
rect 17010 -3465 17060 -3415
rect 17105 -3465 17155 -3415
rect 17225 -3465 17275 -3415
rect 17320 -3465 17370 -3415
rect 17415 -3465 17465 -3415
rect 17515 -3465 17565 -3415
rect 17615 -3465 17665 -3415
rect 17715 -3465 17765 -3415
rect 17810 -3465 17860 -3415
rect 17905 -3465 17955 -3415
rect 14825 -3565 14875 -3515
rect 14920 -3565 14970 -3515
rect 15015 -3565 15065 -3515
rect 15115 -3565 15165 -3515
rect 15215 -3565 15265 -3515
rect 15315 -3565 15365 -3515
rect 15410 -3565 15460 -3515
rect 15505 -3565 15555 -3515
rect 15625 -3565 15675 -3515
rect 15720 -3565 15770 -3515
rect 15815 -3565 15865 -3515
rect 15915 -3565 15965 -3515
rect 16015 -3565 16065 -3515
rect 16115 -3565 16165 -3515
rect 16210 -3565 16260 -3515
rect 16305 -3565 16355 -3515
rect 16425 -3565 16475 -3515
rect 16520 -3565 16570 -3515
rect 16615 -3565 16665 -3515
rect 16715 -3565 16765 -3515
rect 16815 -3565 16865 -3515
rect 16915 -3565 16965 -3515
rect 17010 -3565 17060 -3515
rect 17105 -3565 17155 -3515
rect 17225 -3565 17275 -3515
rect 17320 -3565 17370 -3515
rect 17415 -3565 17465 -3515
rect 17515 -3565 17565 -3515
rect 17615 -3565 17665 -3515
rect 17715 -3565 17765 -3515
rect 17810 -3565 17860 -3515
rect 17905 -3565 17955 -3515
rect 14825 -3655 14875 -3605
rect 14920 -3655 14970 -3605
rect 15015 -3655 15065 -3605
rect 15115 -3655 15165 -3605
rect 15215 -3655 15265 -3605
rect 15315 -3655 15365 -3605
rect 15410 -3655 15460 -3605
rect 15505 -3655 15555 -3605
rect 15625 -3655 15675 -3605
rect 15720 -3655 15770 -3605
rect 15815 -3655 15865 -3605
rect 15915 -3655 15965 -3605
rect 16015 -3655 16065 -3605
rect 16115 -3655 16165 -3605
rect 16210 -3655 16260 -3605
rect 16305 -3655 16355 -3605
rect 16425 -3655 16475 -3605
rect 16520 -3655 16570 -3605
rect 16615 -3655 16665 -3605
rect 16715 -3655 16765 -3605
rect 16815 -3655 16865 -3605
rect 16915 -3655 16965 -3605
rect 17010 -3655 17060 -3605
rect 17105 -3655 17155 -3605
rect 17225 -3655 17275 -3605
rect 17320 -3655 17370 -3605
rect 17415 -3655 17465 -3605
rect 17515 -3655 17565 -3605
rect 17615 -3655 17665 -3605
rect 17715 -3655 17765 -3605
rect 17810 -3655 17860 -3605
rect 17905 -3655 17955 -3605
rect 14825 -3775 14875 -3725
rect 14920 -3775 14970 -3725
rect 15015 -3775 15065 -3725
rect 15115 -3775 15165 -3725
rect 15215 -3775 15265 -3725
rect 15315 -3775 15365 -3725
rect 15410 -3775 15460 -3725
rect 15505 -3775 15555 -3725
rect 15625 -3775 15675 -3725
rect 15720 -3775 15770 -3725
rect 15815 -3775 15865 -3725
rect 15915 -3775 15965 -3725
rect 16015 -3775 16065 -3725
rect 16115 -3775 16165 -3725
rect 16210 -3775 16260 -3725
rect 16305 -3775 16355 -3725
rect 16425 -3775 16475 -3725
rect 16520 -3775 16570 -3725
rect 16615 -3775 16665 -3725
rect 16715 -3775 16765 -3725
rect 16815 -3775 16865 -3725
rect 16915 -3775 16965 -3725
rect 17010 -3775 17060 -3725
rect 17105 -3775 17155 -3725
rect 17225 -3775 17275 -3725
rect 17320 -3775 17370 -3725
rect 17415 -3775 17465 -3725
rect 17515 -3775 17565 -3725
rect 17615 -3775 17665 -3725
rect 17715 -3775 17765 -3725
rect 17810 -3775 17860 -3725
rect 17905 -3775 17955 -3725
rect 14825 -3865 14875 -3815
rect 14920 -3865 14970 -3815
rect 15015 -3865 15065 -3815
rect 15115 -3865 15165 -3815
rect 15215 -3865 15265 -3815
rect 15315 -3865 15365 -3815
rect 15410 -3865 15460 -3815
rect 15505 -3865 15555 -3815
rect 15625 -3865 15675 -3815
rect 15720 -3865 15770 -3815
rect 15815 -3865 15865 -3815
rect 15915 -3865 15965 -3815
rect 16015 -3865 16065 -3815
rect 16115 -3865 16165 -3815
rect 16210 -3865 16260 -3815
rect 16305 -3865 16355 -3815
rect 16425 -3865 16475 -3815
rect 16520 -3865 16570 -3815
rect 16615 -3865 16665 -3815
rect 16715 -3865 16765 -3815
rect 16815 -3865 16865 -3815
rect 16915 -3865 16965 -3815
rect 17010 -3865 17060 -3815
rect 17105 -3865 17155 -3815
rect 17225 -3865 17275 -3815
rect 17320 -3865 17370 -3815
rect 17415 -3865 17465 -3815
rect 17515 -3865 17565 -3815
rect 17615 -3865 17665 -3815
rect 17715 -3865 17765 -3815
rect 17810 -3865 17860 -3815
rect 17905 -3865 17955 -3815
rect 14825 -3965 14875 -3915
rect 14920 -3965 14970 -3915
rect 15015 -3965 15065 -3915
rect 15115 -3965 15165 -3915
rect 15215 -3965 15265 -3915
rect 15315 -3965 15365 -3915
rect 15410 -3965 15460 -3915
rect 15505 -3965 15555 -3915
rect 15625 -3965 15675 -3915
rect 15720 -3965 15770 -3915
rect 15815 -3965 15865 -3915
rect 15915 -3965 15965 -3915
rect 16015 -3965 16065 -3915
rect 16115 -3965 16165 -3915
rect 16210 -3965 16260 -3915
rect 16305 -3965 16355 -3915
rect 16425 -3965 16475 -3915
rect 16520 -3965 16570 -3915
rect 16615 -3965 16665 -3915
rect 16715 -3965 16765 -3915
rect 16815 -3965 16865 -3915
rect 16915 -3965 16965 -3915
rect 17010 -3965 17060 -3915
rect 17105 -3965 17155 -3915
rect 17225 -3965 17275 -3915
rect 17320 -3965 17370 -3915
rect 17415 -3965 17465 -3915
rect 17515 -3965 17565 -3915
rect 17615 -3965 17665 -3915
rect 17715 -3965 17765 -3915
rect 17810 -3965 17860 -3915
rect 17905 -3965 17955 -3915
rect 14825 -4055 14875 -4005
rect 14920 -4055 14970 -4005
rect 15015 -4055 15065 -4005
rect 15115 -4055 15165 -4005
rect 15215 -4055 15265 -4005
rect 15315 -4055 15365 -4005
rect 15410 -4055 15460 -4005
rect 15505 -4055 15555 -4005
rect 15625 -4055 15675 -4005
rect 15720 -4055 15770 -4005
rect 15815 -4055 15865 -4005
rect 15915 -4055 15965 -4005
rect 16015 -4055 16065 -4005
rect 16115 -4055 16165 -4005
rect 16210 -4055 16260 -4005
rect 16305 -4055 16355 -4005
rect 16425 -4055 16475 -4005
rect 16520 -4055 16570 -4005
rect 16615 -4055 16665 -4005
rect 16715 -4055 16765 -4005
rect 16815 -4055 16865 -4005
rect 16915 -4055 16965 -4005
rect 17010 -4055 17060 -4005
rect 17105 -4055 17155 -4005
rect 17225 -4055 17275 -4005
rect 17320 -4055 17370 -4005
rect 17415 -4055 17465 -4005
rect 17515 -4055 17565 -4005
rect 17615 -4055 17665 -4005
rect 17715 -4055 17765 -4005
rect 17810 -4055 17860 -4005
rect 17905 -4055 17955 -4005
rect 14825 -4175 14875 -4125
rect 14920 -4175 14970 -4125
rect 15015 -4175 15065 -4125
rect 15115 -4175 15165 -4125
rect 15215 -4175 15265 -4125
rect 15315 -4175 15365 -4125
rect 15410 -4175 15460 -4125
rect 15505 -4175 15555 -4125
rect 15625 -4175 15675 -4125
rect 15720 -4175 15770 -4125
rect 15815 -4175 15865 -4125
rect 15915 -4175 15965 -4125
rect 16015 -4175 16065 -4125
rect 16115 -4175 16165 -4125
rect 16210 -4175 16260 -4125
rect 16305 -4175 16355 -4125
rect 16425 -4175 16475 -4125
rect 16520 -4175 16570 -4125
rect 16615 -4175 16665 -4125
rect 16715 -4175 16765 -4125
rect 16815 -4175 16865 -4125
rect 16915 -4175 16965 -4125
rect 17010 -4175 17060 -4125
rect 17105 -4175 17155 -4125
rect 17225 -4175 17275 -4125
rect 17320 -4175 17370 -4125
rect 17415 -4175 17465 -4125
rect 17515 -4175 17565 -4125
rect 17615 -4175 17665 -4125
rect 17715 -4175 17765 -4125
rect 17810 -4175 17860 -4125
rect 17905 -4175 17955 -4125
rect 14825 -4265 14875 -4215
rect 14920 -4265 14970 -4215
rect 15015 -4265 15065 -4215
rect 15115 -4265 15165 -4215
rect 15215 -4265 15265 -4215
rect 15315 -4265 15365 -4215
rect 15410 -4265 15460 -4215
rect 15505 -4265 15555 -4215
rect 15625 -4265 15675 -4215
rect 15720 -4265 15770 -4215
rect 15815 -4265 15865 -4215
rect 15915 -4265 15965 -4215
rect 16015 -4265 16065 -4215
rect 16115 -4265 16165 -4215
rect 16210 -4265 16260 -4215
rect 16305 -4265 16355 -4215
rect 16425 -4265 16475 -4215
rect 16520 -4265 16570 -4215
rect 16615 -4265 16665 -4215
rect 16715 -4265 16765 -4215
rect 16815 -4265 16865 -4215
rect 16915 -4265 16965 -4215
rect 17010 -4265 17060 -4215
rect 17105 -4265 17155 -4215
rect 17225 -4265 17275 -4215
rect 17320 -4265 17370 -4215
rect 17415 -4265 17465 -4215
rect 17515 -4265 17565 -4215
rect 17615 -4265 17665 -4215
rect 17715 -4265 17765 -4215
rect 17810 -4265 17860 -4215
rect 17905 -4265 17955 -4215
rect 14825 -4365 14875 -4315
rect 14920 -4365 14970 -4315
rect 15015 -4365 15065 -4315
rect 15115 -4365 15165 -4315
rect 15215 -4365 15265 -4315
rect 15315 -4365 15365 -4315
rect 15410 -4365 15460 -4315
rect 15505 -4365 15555 -4315
rect 15625 -4365 15675 -4315
rect 15720 -4365 15770 -4315
rect 15815 -4365 15865 -4315
rect 15915 -4365 15965 -4315
rect 16015 -4365 16065 -4315
rect 16115 -4365 16165 -4315
rect 16210 -4365 16260 -4315
rect 16305 -4365 16355 -4315
rect 16425 -4365 16475 -4315
rect 16520 -4365 16570 -4315
rect 16615 -4365 16665 -4315
rect 16715 -4365 16765 -4315
rect 16815 -4365 16865 -4315
rect 16915 -4365 16965 -4315
rect 17010 -4365 17060 -4315
rect 17105 -4365 17155 -4315
rect 17225 -4365 17275 -4315
rect 17320 -4365 17370 -4315
rect 17415 -4365 17465 -4315
rect 17515 -4365 17565 -4315
rect 17615 -4365 17665 -4315
rect 17715 -4365 17765 -4315
rect 17810 -4365 17860 -4315
rect 17905 -4365 17955 -4315
rect 14825 -4455 14875 -4405
rect 14920 -4455 14970 -4405
rect 15015 -4455 15065 -4405
rect 15115 -4455 15165 -4405
rect 15215 -4455 15265 -4405
rect 15315 -4455 15365 -4405
rect 15410 -4455 15460 -4405
rect 15505 -4455 15555 -4405
rect 15625 -4455 15675 -4405
rect 15720 -4455 15770 -4405
rect 15815 -4455 15865 -4405
rect 15915 -4455 15965 -4405
rect 16015 -4455 16065 -4405
rect 16115 -4455 16165 -4405
rect 16210 -4455 16260 -4405
rect 16305 -4455 16355 -4405
rect 16425 -4455 16475 -4405
rect 16520 -4455 16570 -4405
rect 16615 -4455 16665 -4405
rect 16715 -4455 16765 -4405
rect 16815 -4455 16865 -4405
rect 16915 -4455 16965 -4405
rect 17010 -4455 17060 -4405
rect 17105 -4455 17155 -4405
rect 17225 -4455 17275 -4405
rect 17320 -4455 17370 -4405
rect 17415 -4455 17465 -4405
rect 17515 -4455 17565 -4405
rect 17615 -4455 17665 -4405
rect 17715 -4455 17765 -4405
rect 17810 -4455 17860 -4405
rect 17905 -4455 17955 -4405
<< mimcap >>
rect -1245 18140 -1045 18215
rect -1245 18100 -1165 18140
rect -1125 18100 -1045 18140
rect -1245 18015 -1045 18100
rect -895 18140 -695 18215
rect -895 18100 -815 18140
rect -775 18100 -695 18140
rect -895 18015 -695 18100
rect -545 18140 -345 18215
rect -545 18100 -465 18140
rect -425 18100 -345 18140
rect -545 18015 -345 18100
rect -195 18140 5 18215
rect -195 18100 -115 18140
rect -75 18100 5 18140
rect -195 18015 5 18100
rect 155 18140 355 18215
rect 155 18100 235 18140
rect 275 18100 355 18140
rect 155 18015 355 18100
rect 505 18140 705 18215
rect 505 18100 585 18140
rect 625 18100 705 18140
rect 505 18015 705 18100
rect 855 18140 1055 18215
rect 855 18100 935 18140
rect 975 18100 1055 18140
rect 855 18015 1055 18100
rect 1205 18140 1405 18215
rect 1205 18100 1285 18140
rect 1325 18100 1405 18140
rect 1205 18015 1405 18100
rect 1555 18140 1755 18215
rect 1555 18100 1635 18140
rect 1675 18100 1755 18140
rect 1555 18015 1755 18100
rect -1245 17790 -1045 17865
rect -1245 17750 -1165 17790
rect -1125 17750 -1045 17790
rect -1245 17665 -1045 17750
rect -895 17790 -695 17865
rect -895 17750 -815 17790
rect -775 17750 -695 17790
rect -895 17665 -695 17750
rect -545 17790 -345 17865
rect -545 17750 -465 17790
rect -425 17750 -345 17790
rect -545 17665 -345 17750
rect -195 17790 5 17865
rect -195 17750 -115 17790
rect -75 17750 5 17790
rect -195 17665 5 17750
rect 155 17790 355 17865
rect 155 17750 235 17790
rect 275 17750 355 17790
rect 155 17665 355 17750
rect 505 17790 705 17865
rect 505 17750 585 17790
rect 625 17750 705 17790
rect 505 17665 705 17750
rect 855 17790 1055 17865
rect 855 17750 935 17790
rect 975 17750 1055 17790
rect 855 17665 1055 17750
rect 1205 17790 1405 17865
rect 1205 17750 1285 17790
rect 1325 17750 1405 17790
rect 1205 17665 1405 17750
rect 1555 17790 1755 17865
rect 1555 17750 1635 17790
rect 1675 17750 1755 17790
rect 1555 17665 1755 17750
rect -1245 17440 -1045 17515
rect -1245 17400 -1165 17440
rect -1125 17400 -1045 17440
rect -1245 17315 -1045 17400
rect -895 17440 -695 17515
rect -895 17400 -815 17440
rect -775 17400 -695 17440
rect -895 17315 -695 17400
rect -545 17440 -345 17515
rect -545 17400 -465 17440
rect -425 17400 -345 17440
rect -545 17315 -345 17400
rect -195 17440 5 17515
rect -195 17400 -115 17440
rect -75 17400 5 17440
rect -195 17315 5 17400
rect 155 17440 355 17515
rect 155 17400 235 17440
rect 275 17400 355 17440
rect 155 17315 355 17400
rect 505 17440 705 17515
rect 505 17400 585 17440
rect 625 17400 705 17440
rect 505 17315 705 17400
rect 855 17440 1055 17515
rect 855 17400 935 17440
rect 975 17400 1055 17440
rect 855 17315 1055 17400
rect 1205 17440 1405 17515
rect 1205 17400 1285 17440
rect 1325 17400 1405 17440
rect 1205 17315 1405 17400
rect 1555 17440 1755 17515
rect 1555 17400 1635 17440
rect 1675 17400 1755 17440
rect 1555 17315 1755 17400
rect 9555 17440 9755 17515
rect 9555 17400 9635 17440
rect 9675 17400 9755 17440
rect 9555 17315 9755 17400
rect 9905 17440 10105 17515
rect 9905 17400 9985 17440
rect 10025 17400 10105 17440
rect 9905 17315 10105 17400
rect 10255 17440 10455 17515
rect 10255 17400 10335 17440
rect 10375 17400 10455 17440
rect 10255 17315 10455 17400
rect 10605 17440 10805 17515
rect 10605 17400 10685 17440
rect 10725 17400 10805 17440
rect 10605 17315 10805 17400
rect 10955 17440 11155 17515
rect 10955 17400 11035 17440
rect 11075 17400 11155 17440
rect 10955 17315 11155 17400
rect 11305 17440 11505 17515
rect 11305 17400 11385 17440
rect 11425 17400 11505 17440
rect 11305 17315 11505 17400
rect 11655 17440 11855 17515
rect 11655 17400 11735 17440
rect 11775 17400 11855 17440
rect 11655 17315 11855 17400
rect 12005 17440 12205 17515
rect 12005 17400 12085 17440
rect 12125 17400 12205 17440
rect 12005 17315 12205 17400
rect 12355 17440 12555 17515
rect 12355 17400 12435 17440
rect 12475 17400 12555 17440
rect 12355 17315 12555 17400
rect 12705 17440 12905 17515
rect 12705 17400 12785 17440
rect 12825 17400 12905 17440
rect 12705 17315 12905 17400
rect 13055 17440 13255 17515
rect 13055 17400 13135 17440
rect 13175 17400 13255 17440
rect 13055 17315 13255 17400
rect 13405 17440 13605 17515
rect 13405 17400 13485 17440
rect 13525 17400 13605 17440
rect 13405 17315 13605 17400
rect 13755 17440 13955 17515
rect 13755 17400 13835 17440
rect 13875 17400 13955 17440
rect 13755 17315 13955 17400
rect 14105 17440 14305 17515
rect 14105 17400 14185 17440
rect 14225 17400 14305 17440
rect 14105 17315 14305 17400
rect 14455 17440 14655 17515
rect 14455 17400 14535 17440
rect 14575 17400 14655 17440
rect 14455 17315 14655 17400
rect -1245 17090 -1045 17165
rect -1245 17050 -1165 17090
rect -1125 17050 -1045 17090
rect -1245 16965 -1045 17050
rect -895 17090 -695 17165
rect -895 17050 -815 17090
rect -775 17050 -695 17090
rect -895 16965 -695 17050
rect -545 17090 -345 17165
rect -545 17050 -465 17090
rect -425 17050 -345 17090
rect -545 16965 -345 17050
rect -195 17090 5 17165
rect -195 17050 -115 17090
rect -75 17050 5 17090
rect -195 16965 5 17050
rect 155 17090 355 17165
rect 155 17050 235 17090
rect 275 17050 355 17090
rect 155 16965 355 17050
rect 505 17090 705 17165
rect 505 17050 585 17090
rect 625 17050 705 17090
rect 505 16965 705 17050
rect 855 17090 1055 17165
rect 855 17050 935 17090
rect 975 17050 1055 17090
rect 855 16965 1055 17050
rect 1205 17090 1405 17165
rect 1205 17050 1285 17090
rect 1325 17050 1405 17090
rect 1205 16965 1405 17050
rect 1555 17090 1755 17165
rect 1555 17050 1635 17090
rect 1675 17050 1755 17090
rect 1555 16965 1755 17050
rect 9555 17090 9755 17165
rect 9555 17050 9635 17090
rect 9675 17050 9755 17090
rect 9555 16965 9755 17050
rect 9905 17090 10105 17165
rect 9905 17050 9985 17090
rect 10025 17050 10105 17090
rect 9905 16965 10105 17050
rect 10255 17090 10455 17165
rect 10255 17050 10335 17090
rect 10375 17050 10455 17090
rect 10255 16965 10455 17050
rect 10605 17090 10805 17165
rect 10605 17050 10685 17090
rect 10725 17050 10805 17090
rect 10605 16965 10805 17050
rect 10955 17090 11155 17165
rect 10955 17050 11035 17090
rect 11075 17050 11155 17090
rect 10955 16965 11155 17050
rect 11305 17090 11505 17165
rect 11305 17050 11385 17090
rect 11425 17050 11505 17090
rect 11305 16965 11505 17050
rect 11655 17090 11855 17165
rect 11655 17050 11735 17090
rect 11775 17050 11855 17090
rect 11655 16965 11855 17050
rect 12005 17090 12205 17165
rect 12005 17050 12085 17090
rect 12125 17050 12205 17090
rect 12005 16965 12205 17050
rect 12355 17090 12555 17165
rect 12355 17050 12435 17090
rect 12475 17050 12555 17090
rect 12355 16965 12555 17050
rect 12705 17090 12905 17165
rect 12705 17050 12785 17090
rect 12825 17050 12905 17090
rect 12705 16965 12905 17050
rect 13055 17090 13255 17165
rect 13055 17050 13135 17090
rect 13175 17050 13255 17090
rect 13055 16965 13255 17050
rect 13405 17090 13605 17165
rect 13405 17050 13485 17090
rect 13525 17050 13605 17090
rect 13405 16965 13605 17050
rect 13755 17090 13955 17165
rect 13755 17050 13835 17090
rect 13875 17050 13955 17090
rect 13755 16965 13955 17050
rect 14105 17090 14305 17165
rect 14105 17050 14185 17090
rect 14225 17050 14305 17090
rect 14105 16965 14305 17050
rect 14455 17090 14655 17165
rect 14455 17050 14535 17090
rect 14575 17050 14655 17090
rect 14455 16965 14655 17050
rect -1245 16740 -1045 16815
rect -1245 16700 -1165 16740
rect -1125 16700 -1045 16740
rect -1245 16615 -1045 16700
rect -895 16740 -695 16815
rect -895 16700 -815 16740
rect -775 16700 -695 16740
rect -895 16615 -695 16700
rect -545 16740 -345 16815
rect -545 16700 -465 16740
rect -425 16700 -345 16740
rect -545 16615 -345 16700
rect -195 16740 5 16815
rect -195 16700 -115 16740
rect -75 16700 5 16740
rect -195 16615 5 16700
rect 155 16740 355 16815
rect 155 16700 235 16740
rect 275 16700 355 16740
rect 155 16615 355 16700
rect 505 16740 705 16815
rect 505 16700 585 16740
rect 625 16700 705 16740
rect 505 16615 705 16700
rect 855 16740 1055 16815
rect 855 16700 935 16740
rect 975 16700 1055 16740
rect 855 16615 1055 16700
rect 1205 16740 1405 16815
rect 1205 16700 1285 16740
rect 1325 16700 1405 16740
rect 1205 16615 1405 16700
rect 1555 16740 1755 16815
rect 1555 16700 1635 16740
rect 1675 16700 1755 16740
rect 1555 16615 1755 16700
rect 9555 16740 9755 16815
rect 9555 16700 9635 16740
rect 9675 16700 9755 16740
rect 9555 16615 9755 16700
rect 9905 16740 10105 16815
rect 9905 16700 9985 16740
rect 10025 16700 10105 16740
rect 9905 16615 10105 16700
rect 10255 16740 10455 16815
rect 10255 16700 10335 16740
rect 10375 16700 10455 16740
rect 10255 16615 10455 16700
rect 10605 16740 10805 16815
rect 10605 16700 10685 16740
rect 10725 16700 10805 16740
rect 10605 16615 10805 16700
rect 10955 16740 11155 16815
rect 10955 16700 11035 16740
rect 11075 16700 11155 16740
rect 10955 16615 11155 16700
rect 11305 16740 11505 16815
rect 11305 16700 11385 16740
rect 11425 16700 11505 16740
rect 11305 16615 11505 16700
rect 11655 16740 11855 16815
rect 11655 16700 11735 16740
rect 11775 16700 11855 16740
rect 11655 16615 11855 16700
rect 12005 16740 12205 16815
rect 12005 16700 12085 16740
rect 12125 16700 12205 16740
rect 12005 16615 12205 16700
rect 12355 16740 12555 16815
rect 12355 16700 12435 16740
rect 12475 16700 12555 16740
rect 12355 16615 12555 16700
rect 12705 16740 12905 16815
rect 12705 16700 12785 16740
rect 12825 16700 12905 16740
rect 12705 16615 12905 16700
rect 13055 16740 13255 16815
rect 13055 16700 13135 16740
rect 13175 16700 13255 16740
rect 13055 16615 13255 16700
rect 13405 16740 13605 16815
rect 13405 16700 13485 16740
rect 13525 16700 13605 16740
rect 13405 16615 13605 16700
rect 13755 16740 13955 16815
rect 13755 16700 13835 16740
rect 13875 16700 13955 16740
rect 13755 16615 13955 16700
rect 14105 16740 14305 16815
rect 14105 16700 14185 16740
rect 14225 16700 14305 16740
rect 14105 16615 14305 16700
rect 14455 16740 14655 16815
rect 14455 16700 14535 16740
rect 14575 16700 14655 16740
rect 14455 16615 14655 16700
rect -1245 16390 -1045 16465
rect -1245 16350 -1165 16390
rect -1125 16350 -1045 16390
rect -1245 16265 -1045 16350
rect -895 16390 -695 16465
rect -895 16350 -815 16390
rect -775 16350 -695 16390
rect -895 16265 -695 16350
rect -545 16390 -345 16465
rect -545 16350 -465 16390
rect -425 16350 -345 16390
rect -545 16265 -345 16350
rect -195 16390 5 16465
rect -195 16350 -115 16390
rect -75 16350 5 16390
rect -195 16265 5 16350
rect 155 16390 355 16465
rect 155 16350 235 16390
rect 275 16350 355 16390
rect 155 16265 355 16350
rect 505 16390 705 16465
rect 505 16350 585 16390
rect 625 16350 705 16390
rect 505 16265 705 16350
rect 855 16390 1055 16465
rect 855 16350 935 16390
rect 975 16350 1055 16390
rect 855 16265 1055 16350
rect 1205 16390 1405 16465
rect 1205 16350 1285 16390
rect 1325 16350 1405 16390
rect 1205 16265 1405 16350
rect 1555 16390 1755 16465
rect 1555 16350 1635 16390
rect 1675 16350 1755 16390
rect 1555 16265 1755 16350
rect 9555 16390 9755 16465
rect 9555 16350 9635 16390
rect 9675 16350 9755 16390
rect 9555 16265 9755 16350
rect 9905 16390 10105 16465
rect 9905 16350 9985 16390
rect 10025 16350 10105 16390
rect 9905 16265 10105 16350
rect 10255 16390 10455 16465
rect 10255 16350 10335 16390
rect 10375 16350 10455 16390
rect 10255 16265 10455 16350
rect 10605 16390 10805 16465
rect 10605 16350 10685 16390
rect 10725 16350 10805 16390
rect 10605 16265 10805 16350
rect 10955 16390 11155 16465
rect 10955 16350 11035 16390
rect 11075 16350 11155 16390
rect 10955 16265 11155 16350
rect 11305 16390 11505 16465
rect 11305 16350 11385 16390
rect 11425 16350 11505 16390
rect 11305 16265 11505 16350
rect 11655 16390 11855 16465
rect 11655 16350 11735 16390
rect 11775 16350 11855 16390
rect 11655 16265 11855 16350
rect 12005 16390 12205 16465
rect 12005 16350 12085 16390
rect 12125 16350 12205 16390
rect 12005 16265 12205 16350
rect 12355 16390 12555 16465
rect 12355 16350 12435 16390
rect 12475 16350 12555 16390
rect 12355 16265 12555 16350
rect 12705 16390 12905 16465
rect 12705 16350 12785 16390
rect 12825 16350 12905 16390
rect 12705 16265 12905 16350
rect 13055 16390 13255 16465
rect 13055 16350 13135 16390
rect 13175 16350 13255 16390
rect 13055 16265 13255 16350
rect 13405 16390 13605 16465
rect 13405 16350 13485 16390
rect 13525 16350 13605 16390
rect 13405 16265 13605 16350
rect 13755 16390 13955 16465
rect 13755 16350 13835 16390
rect 13875 16350 13955 16390
rect 13755 16265 13955 16350
rect 14105 16390 14305 16465
rect 14105 16350 14185 16390
rect 14225 16350 14305 16390
rect 14105 16265 14305 16350
rect 14455 16390 14655 16465
rect 14455 16350 14535 16390
rect 14575 16350 14655 16390
rect 14455 16265 14655 16350
rect -1245 16040 -1045 16115
rect -1245 16000 -1165 16040
rect -1125 16000 -1045 16040
rect -1245 15915 -1045 16000
rect -895 16040 -695 16115
rect -895 16000 -815 16040
rect -775 16000 -695 16040
rect -895 15915 -695 16000
rect -545 16040 -345 16115
rect -545 16000 -465 16040
rect -425 16000 -345 16040
rect -545 15915 -345 16000
rect -195 16040 5 16115
rect -195 16000 -115 16040
rect -75 16000 5 16040
rect -195 15915 5 16000
rect 155 16040 355 16115
rect 155 16000 235 16040
rect 275 16000 355 16040
rect 155 15915 355 16000
rect 505 16040 705 16115
rect 505 16000 585 16040
rect 625 16000 705 16040
rect 505 15915 705 16000
rect 855 16040 1055 16115
rect 855 16000 935 16040
rect 975 16000 1055 16040
rect 855 15915 1055 16000
rect 1205 16040 1405 16115
rect 1205 16000 1285 16040
rect 1325 16000 1405 16040
rect 1205 15915 1405 16000
rect 1555 16040 1755 16115
rect 1555 16000 1635 16040
rect 1675 16000 1755 16040
rect 1555 15915 1755 16000
rect 9555 16040 9755 16115
rect 9555 16000 9635 16040
rect 9675 16000 9755 16040
rect 9555 15915 9755 16000
rect 9905 16040 10105 16115
rect 9905 16000 9985 16040
rect 10025 16000 10105 16040
rect 9905 15915 10105 16000
rect 10255 16040 10455 16115
rect 10255 16000 10335 16040
rect 10375 16000 10455 16040
rect 10255 15915 10455 16000
rect 10605 16040 10805 16115
rect 10605 16000 10685 16040
rect 10725 16000 10805 16040
rect 10605 15915 10805 16000
rect 10955 16040 11155 16115
rect 10955 16000 11035 16040
rect 11075 16000 11155 16040
rect 10955 15915 11155 16000
rect 11305 16040 11505 16115
rect 11305 16000 11385 16040
rect 11425 16000 11505 16040
rect 11305 15915 11505 16000
rect 11655 16040 11855 16115
rect 11655 16000 11735 16040
rect 11775 16000 11855 16040
rect 11655 15915 11855 16000
rect 12005 16040 12205 16115
rect 12005 16000 12085 16040
rect 12125 16000 12205 16040
rect 12005 15915 12205 16000
rect 12355 16040 12555 16115
rect 12355 16000 12435 16040
rect 12475 16000 12555 16040
rect 12355 15915 12555 16000
rect 12705 16040 12905 16115
rect 12705 16000 12785 16040
rect 12825 16000 12905 16040
rect 12705 15915 12905 16000
rect 13055 16040 13255 16115
rect 13055 16000 13135 16040
rect 13175 16000 13255 16040
rect 13055 15915 13255 16000
rect 13405 16040 13605 16115
rect 13405 16000 13485 16040
rect 13525 16000 13605 16040
rect 13405 15915 13605 16000
rect 13755 16040 13955 16115
rect 13755 16000 13835 16040
rect 13875 16000 13955 16040
rect 13755 15915 13955 16000
rect 14105 16040 14305 16115
rect 14105 16000 14185 16040
rect 14225 16000 14305 16040
rect 14105 15915 14305 16000
rect 14455 16040 14655 16115
rect 14455 16000 14535 16040
rect 14575 16000 14655 16040
rect 14455 15915 14655 16000
rect -1245 15690 -1045 15765
rect -1245 15650 -1165 15690
rect -1125 15650 -1045 15690
rect -1245 15565 -1045 15650
rect -895 15690 -695 15765
rect -895 15650 -815 15690
rect -775 15650 -695 15690
rect -895 15565 -695 15650
rect -545 15690 -345 15765
rect -545 15650 -465 15690
rect -425 15650 -345 15690
rect -545 15565 -345 15650
rect -195 15690 5 15765
rect -195 15650 -115 15690
rect -75 15650 5 15690
rect -195 15565 5 15650
rect 155 15690 355 15765
rect 155 15650 235 15690
rect 275 15650 355 15690
rect 155 15565 355 15650
rect 505 15690 705 15765
rect 505 15650 585 15690
rect 625 15650 705 15690
rect 505 15565 705 15650
rect 855 15690 1055 15765
rect 855 15650 935 15690
rect 975 15650 1055 15690
rect 855 15565 1055 15650
rect 1205 15690 1405 15765
rect 1205 15650 1285 15690
rect 1325 15650 1405 15690
rect 1205 15565 1405 15650
rect 1555 15690 1755 15765
rect 1555 15650 1635 15690
rect 1675 15650 1755 15690
rect 1555 15565 1755 15650
rect 9555 15690 9755 15765
rect 9555 15650 9635 15690
rect 9675 15650 9755 15690
rect 9555 15565 9755 15650
rect 9905 15690 10105 15765
rect 9905 15650 9985 15690
rect 10025 15650 10105 15690
rect 9905 15565 10105 15650
rect 10255 15690 10455 15765
rect 10255 15650 10335 15690
rect 10375 15650 10455 15690
rect 10255 15565 10455 15650
rect 10605 15690 10805 15765
rect 10605 15650 10685 15690
rect 10725 15650 10805 15690
rect 10605 15565 10805 15650
rect 10955 15690 11155 15765
rect 10955 15650 11035 15690
rect 11075 15650 11155 15690
rect 10955 15565 11155 15650
rect 11305 15690 11505 15765
rect 11305 15650 11385 15690
rect 11425 15650 11505 15690
rect 11305 15565 11505 15650
rect 11655 15690 11855 15765
rect 11655 15650 11735 15690
rect 11775 15650 11855 15690
rect 11655 15565 11855 15650
rect 12005 15690 12205 15765
rect 12005 15650 12085 15690
rect 12125 15650 12205 15690
rect 12005 15565 12205 15650
rect 12355 15690 12555 15765
rect 12355 15650 12435 15690
rect 12475 15650 12555 15690
rect 12355 15565 12555 15650
rect 12705 15690 12905 15765
rect 12705 15650 12785 15690
rect 12825 15650 12905 15690
rect 12705 15565 12905 15650
rect 13055 15690 13255 15765
rect 13055 15650 13135 15690
rect 13175 15650 13255 15690
rect 13055 15565 13255 15650
rect 13405 15690 13605 15765
rect 13405 15650 13485 15690
rect 13525 15650 13605 15690
rect 13405 15565 13605 15650
rect 13755 15690 13955 15765
rect 13755 15650 13835 15690
rect 13875 15650 13955 15690
rect 13755 15565 13955 15650
rect 14105 15690 14305 15765
rect 14105 15650 14185 15690
rect 14225 15650 14305 15690
rect 14105 15565 14305 15650
rect 14455 15690 14655 15765
rect 14455 15650 14535 15690
rect 14575 15650 14655 15690
rect 14455 15565 14655 15650
rect -1245 15340 -1045 15415
rect -1245 15300 -1165 15340
rect -1125 15300 -1045 15340
rect -1245 15215 -1045 15300
rect -895 15340 -695 15415
rect -895 15300 -815 15340
rect -775 15300 -695 15340
rect -895 15215 -695 15300
rect -545 15340 -345 15415
rect -545 15300 -465 15340
rect -425 15300 -345 15340
rect -545 15215 -345 15300
rect -195 15340 5 15415
rect -195 15300 -115 15340
rect -75 15300 5 15340
rect -195 15215 5 15300
rect 155 15340 355 15415
rect 155 15300 235 15340
rect 275 15300 355 15340
rect 155 15215 355 15300
rect 505 15340 705 15415
rect 505 15300 585 15340
rect 625 15300 705 15340
rect 505 15215 705 15300
rect 855 15340 1055 15415
rect 855 15300 935 15340
rect 975 15300 1055 15340
rect 855 15215 1055 15300
rect 1205 15340 1405 15415
rect 1205 15300 1285 15340
rect 1325 15300 1405 15340
rect 1205 15215 1405 15300
rect 1555 15340 1755 15415
rect 1555 15300 1635 15340
rect 1675 15300 1755 15340
rect 1555 15215 1755 15300
rect 9555 15340 9755 15415
rect 9555 15300 9635 15340
rect 9675 15300 9755 15340
rect 9555 15215 9755 15300
rect 9905 15340 10105 15415
rect 9905 15300 9985 15340
rect 10025 15300 10105 15340
rect 9905 15215 10105 15300
rect 10255 15340 10455 15415
rect 10255 15300 10335 15340
rect 10375 15300 10455 15340
rect 10255 15215 10455 15300
rect 10605 15340 10805 15415
rect 10605 15300 10685 15340
rect 10725 15300 10805 15340
rect 10605 15215 10805 15300
rect 10955 15340 11155 15415
rect 10955 15300 11035 15340
rect 11075 15300 11155 15340
rect 10955 15215 11155 15300
rect 11305 15340 11505 15415
rect 11305 15300 11385 15340
rect 11425 15300 11505 15340
rect 11305 15215 11505 15300
rect 11655 15340 11855 15415
rect 11655 15300 11735 15340
rect 11775 15300 11855 15340
rect 11655 15215 11855 15300
rect 12005 15340 12205 15415
rect 12005 15300 12085 15340
rect 12125 15300 12205 15340
rect 12005 15215 12205 15300
rect 12355 15340 12555 15415
rect 12355 15300 12435 15340
rect 12475 15300 12555 15340
rect 12355 15215 12555 15300
rect 12705 15340 12905 15415
rect 12705 15300 12785 15340
rect 12825 15300 12905 15340
rect 12705 15215 12905 15300
rect 13055 15340 13255 15415
rect 13055 15300 13135 15340
rect 13175 15300 13255 15340
rect 13055 15215 13255 15300
rect 13405 15340 13605 15415
rect 13405 15300 13485 15340
rect 13525 15300 13605 15340
rect 13405 15215 13605 15300
rect 13755 15340 13955 15415
rect 13755 15300 13835 15340
rect 13875 15300 13955 15340
rect 13755 15215 13955 15300
rect 14105 15340 14305 15415
rect 14105 15300 14185 15340
rect 14225 15300 14305 15340
rect 14105 15215 14305 15300
rect 14455 15340 14655 15415
rect 14455 15300 14535 15340
rect 14575 15300 14655 15340
rect 14455 15215 14655 15300
rect -1245 14990 -1045 15065
rect -1245 14950 -1165 14990
rect -1125 14950 -1045 14990
rect -1245 14865 -1045 14950
rect -895 14990 -695 15065
rect -895 14950 -815 14990
rect -775 14950 -695 14990
rect -895 14865 -695 14950
rect -545 14990 -345 15065
rect -545 14950 -465 14990
rect -425 14950 -345 14990
rect -545 14865 -345 14950
rect -195 14990 5 15065
rect -195 14950 -115 14990
rect -75 14950 5 14990
rect -195 14865 5 14950
rect 155 14990 355 15065
rect 155 14950 235 14990
rect 275 14950 355 14990
rect 155 14865 355 14950
rect 505 14990 705 15065
rect 505 14950 585 14990
rect 625 14950 705 14990
rect 505 14865 705 14950
rect 855 14990 1055 15065
rect 855 14950 935 14990
rect 975 14950 1055 14990
rect 855 14865 1055 14950
rect 1205 14990 1405 15065
rect 1205 14950 1285 14990
rect 1325 14950 1405 14990
rect 1205 14865 1405 14950
rect 1555 14990 1755 15065
rect 1555 14950 1635 14990
rect 1675 14950 1755 14990
rect 1555 14865 1755 14950
rect 9555 14990 9755 15065
rect 9555 14950 9635 14990
rect 9675 14950 9755 14990
rect 9555 14865 9755 14950
rect 9905 14990 10105 15065
rect 9905 14950 9985 14990
rect 10025 14950 10105 14990
rect 9905 14865 10105 14950
rect 10255 14990 10455 15065
rect 10255 14950 10335 14990
rect 10375 14950 10455 14990
rect 10255 14865 10455 14950
rect 10605 14990 10805 15065
rect 10605 14950 10685 14990
rect 10725 14950 10805 14990
rect 10605 14865 10805 14950
rect 10955 14990 11155 15065
rect 10955 14950 11035 14990
rect 11075 14950 11155 14990
rect 10955 14865 11155 14950
rect 11305 14990 11505 15065
rect 11305 14950 11385 14990
rect 11425 14950 11505 14990
rect 11305 14865 11505 14950
rect 11655 14990 11855 15065
rect 11655 14950 11735 14990
rect 11775 14950 11855 14990
rect 11655 14865 11855 14950
rect 12005 14990 12205 15065
rect 12005 14950 12085 14990
rect 12125 14950 12205 14990
rect 12005 14865 12205 14950
rect 12355 14990 12555 15065
rect 12355 14950 12435 14990
rect 12475 14950 12555 14990
rect 12355 14865 12555 14950
rect 12705 14990 12905 15065
rect 12705 14950 12785 14990
rect 12825 14950 12905 14990
rect 12705 14865 12905 14950
rect 13055 14990 13255 15065
rect 13055 14950 13135 14990
rect 13175 14950 13255 14990
rect 13055 14865 13255 14950
rect 13405 14990 13605 15065
rect 13405 14950 13485 14990
rect 13525 14950 13605 14990
rect 13405 14865 13605 14950
rect 13755 14990 13955 15065
rect 13755 14950 13835 14990
rect 13875 14950 13955 14990
rect 13755 14865 13955 14950
rect 14105 14990 14305 15065
rect 14105 14950 14185 14990
rect 14225 14950 14305 14990
rect 14105 14865 14305 14950
rect 14455 14990 14655 15065
rect 14455 14950 14535 14990
rect 14575 14950 14655 14990
rect 14455 14865 14655 14950
rect -1245 14640 -1045 14715
rect -1245 14600 -1165 14640
rect -1125 14600 -1045 14640
rect -1245 14515 -1045 14600
rect -895 14640 -695 14715
rect -895 14600 -815 14640
rect -775 14600 -695 14640
rect -895 14515 -695 14600
rect -545 14640 -345 14715
rect -545 14600 -465 14640
rect -425 14600 -345 14640
rect -545 14515 -345 14600
rect -195 14640 5 14715
rect -195 14600 -115 14640
rect -75 14600 5 14640
rect -195 14515 5 14600
rect 155 14640 355 14715
rect 155 14600 235 14640
rect 275 14600 355 14640
rect 155 14515 355 14600
rect 505 14640 705 14715
rect 505 14600 585 14640
rect 625 14600 705 14640
rect 505 14515 705 14600
rect 855 14640 1055 14715
rect 855 14600 935 14640
rect 975 14600 1055 14640
rect 855 14515 1055 14600
rect 1205 14640 1405 14715
rect 1205 14600 1285 14640
rect 1325 14600 1405 14640
rect 1205 14515 1405 14600
rect 1555 14640 1755 14715
rect 1555 14600 1635 14640
rect 1675 14600 1755 14640
rect 1555 14515 1755 14600
rect 9555 14640 9755 14715
rect 9555 14600 9635 14640
rect 9675 14600 9755 14640
rect 9555 14515 9755 14600
rect 9905 14640 10105 14715
rect 9905 14600 9985 14640
rect 10025 14600 10105 14640
rect 9905 14515 10105 14600
rect 10255 14640 10455 14715
rect 10255 14600 10335 14640
rect 10375 14600 10455 14640
rect 10255 14515 10455 14600
rect 10605 14640 10805 14715
rect 10605 14600 10685 14640
rect 10725 14600 10805 14640
rect 10605 14515 10805 14600
rect 10955 14640 11155 14715
rect 10955 14600 11035 14640
rect 11075 14600 11155 14640
rect 10955 14515 11155 14600
rect 11305 14640 11505 14715
rect 11305 14600 11385 14640
rect 11425 14600 11505 14640
rect 11305 14515 11505 14600
rect 11655 14640 11855 14715
rect 11655 14600 11735 14640
rect 11775 14600 11855 14640
rect 11655 14515 11855 14600
rect 12005 14640 12205 14715
rect 12005 14600 12085 14640
rect 12125 14600 12205 14640
rect 12005 14515 12205 14600
rect 12355 14640 12555 14715
rect 12355 14600 12435 14640
rect 12475 14600 12555 14640
rect 12355 14515 12555 14600
rect 12705 14640 12905 14715
rect 12705 14600 12785 14640
rect 12825 14600 12905 14640
rect 12705 14515 12905 14600
rect 13055 14640 13255 14715
rect 13055 14600 13135 14640
rect 13175 14600 13255 14640
rect 13055 14515 13255 14600
rect 13405 14640 13605 14715
rect 13405 14600 13485 14640
rect 13525 14600 13605 14640
rect 13405 14515 13605 14600
rect 13755 14640 13955 14715
rect 13755 14600 13835 14640
rect 13875 14600 13955 14640
rect 13755 14515 13955 14600
rect 14105 14640 14305 14715
rect 14105 14600 14185 14640
rect 14225 14600 14305 14640
rect 14105 14515 14305 14600
rect 14455 14640 14655 14715
rect 14455 14600 14535 14640
rect 14575 14600 14655 14640
rect 14455 14515 14655 14600
rect -1245 14290 -1045 14365
rect -1245 14250 -1165 14290
rect -1125 14250 -1045 14290
rect -1245 14165 -1045 14250
rect -895 14290 -695 14365
rect -895 14250 -815 14290
rect -775 14250 -695 14290
rect -895 14165 -695 14250
rect -545 14290 -345 14365
rect -545 14250 -465 14290
rect -425 14250 -345 14290
rect -545 14165 -345 14250
rect -195 14290 5 14365
rect -195 14250 -115 14290
rect -75 14250 5 14290
rect -195 14165 5 14250
rect 155 14290 355 14365
rect 155 14250 235 14290
rect 275 14250 355 14290
rect 155 14165 355 14250
rect 505 14290 705 14365
rect 505 14250 585 14290
rect 625 14250 705 14290
rect 505 14165 705 14250
rect 855 14290 1055 14365
rect 855 14250 935 14290
rect 975 14250 1055 14290
rect 855 14165 1055 14250
rect 1205 14290 1405 14365
rect 1205 14250 1285 14290
rect 1325 14250 1405 14290
rect 1205 14165 1405 14250
rect 1555 14290 1755 14365
rect 1555 14250 1635 14290
rect 1675 14250 1755 14290
rect 1555 14165 1755 14250
rect 9555 14290 9755 14365
rect 9555 14250 9635 14290
rect 9675 14250 9755 14290
rect 9555 14165 9755 14250
rect 9905 14290 10105 14365
rect 9905 14250 9985 14290
rect 10025 14250 10105 14290
rect 9905 14165 10105 14250
rect 10255 14290 10455 14365
rect 10255 14250 10335 14290
rect 10375 14250 10455 14290
rect 10255 14165 10455 14250
rect 10605 14290 10805 14365
rect 10605 14250 10685 14290
rect 10725 14250 10805 14290
rect 10605 14165 10805 14250
rect 10955 14290 11155 14365
rect 10955 14250 11035 14290
rect 11075 14250 11155 14290
rect 10955 14165 11155 14250
rect 11305 14290 11505 14365
rect 11305 14250 11385 14290
rect 11425 14250 11505 14290
rect 11305 14165 11505 14250
rect 11655 14290 11855 14365
rect 11655 14250 11735 14290
rect 11775 14250 11855 14290
rect 11655 14165 11855 14250
rect 12005 14290 12205 14365
rect 12005 14250 12085 14290
rect 12125 14250 12205 14290
rect 12005 14165 12205 14250
rect 12355 14290 12555 14365
rect 12355 14250 12435 14290
rect 12475 14250 12555 14290
rect 12355 14165 12555 14250
rect 12705 14290 12905 14365
rect 12705 14250 12785 14290
rect 12825 14250 12905 14290
rect 12705 14165 12905 14250
rect 13055 14290 13255 14365
rect 13055 14250 13135 14290
rect 13175 14250 13255 14290
rect 13055 14165 13255 14250
rect 13405 14290 13605 14365
rect 13405 14250 13485 14290
rect 13525 14250 13605 14290
rect 13405 14165 13605 14250
rect 13755 14290 13955 14365
rect 13755 14250 13835 14290
rect 13875 14250 13955 14290
rect 13755 14165 13955 14250
rect 14105 14290 14305 14365
rect 14105 14250 14185 14290
rect 14225 14250 14305 14290
rect 14105 14165 14305 14250
rect 14455 14290 14655 14365
rect 14455 14250 14535 14290
rect 14575 14250 14655 14290
rect 14455 14165 14655 14250
rect -1245 13940 -1045 14015
rect -1245 13900 -1165 13940
rect -1125 13900 -1045 13940
rect -1245 13815 -1045 13900
rect -895 13940 -695 14015
rect -895 13900 -815 13940
rect -775 13900 -695 13940
rect -895 13815 -695 13900
rect -545 13940 -345 14015
rect -545 13900 -465 13940
rect -425 13900 -345 13940
rect -545 13815 -345 13900
rect -195 13940 5 14015
rect -195 13900 -115 13940
rect -75 13900 5 13940
rect -195 13815 5 13900
rect 155 13940 355 14015
rect 155 13900 235 13940
rect 275 13900 355 13940
rect 155 13815 355 13900
rect 505 13940 705 14015
rect 505 13900 585 13940
rect 625 13900 705 13940
rect 505 13815 705 13900
rect 855 13940 1055 14015
rect 855 13900 935 13940
rect 975 13900 1055 13940
rect 855 13815 1055 13900
rect 1205 13940 1405 14015
rect 1205 13900 1285 13940
rect 1325 13900 1405 13940
rect 1205 13815 1405 13900
rect 1555 13940 1755 14015
rect 1555 13900 1635 13940
rect 1675 13900 1755 13940
rect 1555 13815 1755 13900
rect 9555 13940 9755 14015
rect 9555 13900 9635 13940
rect 9675 13900 9755 13940
rect 9555 13815 9755 13900
rect 9905 13940 10105 14015
rect 9905 13900 9985 13940
rect 10025 13900 10105 13940
rect 9905 13815 10105 13900
rect 10255 13940 10455 14015
rect 10255 13900 10335 13940
rect 10375 13900 10455 13940
rect 10255 13815 10455 13900
rect 10605 13940 10805 14015
rect 10605 13900 10685 13940
rect 10725 13900 10805 13940
rect 10605 13815 10805 13900
rect 10955 13940 11155 14015
rect 10955 13900 11035 13940
rect 11075 13900 11155 13940
rect 10955 13815 11155 13900
rect 11305 13940 11505 14015
rect 11305 13900 11385 13940
rect 11425 13900 11505 13940
rect 11305 13815 11505 13900
rect 11655 13940 11855 14015
rect 11655 13900 11735 13940
rect 11775 13900 11855 13940
rect 11655 13815 11855 13900
rect 12005 13940 12205 14015
rect 12005 13900 12085 13940
rect 12125 13900 12205 13940
rect 12005 13815 12205 13900
rect 12355 13940 12555 14015
rect 12355 13900 12435 13940
rect 12475 13900 12555 13940
rect 12355 13815 12555 13900
rect 12705 13940 12905 14015
rect 12705 13900 12785 13940
rect 12825 13900 12905 13940
rect 12705 13815 12905 13900
rect 13055 13940 13255 14015
rect 13055 13900 13135 13940
rect 13175 13900 13255 13940
rect 13055 13815 13255 13900
rect 13405 13940 13605 14015
rect 13405 13900 13485 13940
rect 13525 13900 13605 13940
rect 13405 13815 13605 13900
rect 13755 13940 13955 14015
rect 13755 13900 13835 13940
rect 13875 13900 13955 13940
rect 13755 13815 13955 13900
rect 14105 13940 14305 14015
rect 14105 13900 14185 13940
rect 14225 13900 14305 13940
rect 14105 13815 14305 13900
rect 14455 13940 14655 14015
rect 14455 13900 14535 13940
rect 14575 13900 14655 13940
rect 14455 13815 14655 13900
rect -1245 13590 -1045 13665
rect -1245 13550 -1165 13590
rect -1125 13550 -1045 13590
rect -1245 13465 -1045 13550
rect -895 13590 -695 13665
rect -895 13550 -815 13590
rect -775 13550 -695 13590
rect -895 13465 -695 13550
rect -545 13590 -345 13665
rect -545 13550 -465 13590
rect -425 13550 -345 13590
rect -545 13465 -345 13550
rect -195 13590 5 13665
rect -195 13550 -115 13590
rect -75 13550 5 13590
rect -195 13465 5 13550
rect 155 13590 355 13665
rect 155 13550 235 13590
rect 275 13550 355 13590
rect 155 13465 355 13550
rect 505 13590 705 13665
rect 505 13550 585 13590
rect 625 13550 705 13590
rect 505 13465 705 13550
rect 855 13590 1055 13665
rect 855 13550 935 13590
rect 975 13550 1055 13590
rect 855 13465 1055 13550
rect 1205 13590 1405 13665
rect 1205 13550 1285 13590
rect 1325 13550 1405 13590
rect 1205 13465 1405 13550
rect 1555 13590 1755 13665
rect 1555 13550 1635 13590
rect 1675 13550 1755 13590
rect 1555 13465 1755 13550
rect 9555 13590 9755 13665
rect 9555 13550 9635 13590
rect 9675 13550 9755 13590
rect 9555 13465 9755 13550
rect 9905 13590 10105 13665
rect 9905 13550 9985 13590
rect 10025 13550 10105 13590
rect 9905 13465 10105 13550
rect 10255 13590 10455 13665
rect 10255 13550 10335 13590
rect 10375 13550 10455 13590
rect 10255 13465 10455 13550
rect 10605 13590 10805 13665
rect 10605 13550 10685 13590
rect 10725 13550 10805 13590
rect 10605 13465 10805 13550
rect 10955 13590 11155 13665
rect 10955 13550 11035 13590
rect 11075 13550 11155 13590
rect 10955 13465 11155 13550
rect 11305 13590 11505 13665
rect 11305 13550 11385 13590
rect 11425 13550 11505 13590
rect 11305 13465 11505 13550
rect 11655 13590 11855 13665
rect 11655 13550 11735 13590
rect 11775 13550 11855 13590
rect 11655 13465 11855 13550
rect 12005 13590 12205 13665
rect 12005 13550 12085 13590
rect 12125 13550 12205 13590
rect 12005 13465 12205 13550
rect 12355 13590 12555 13665
rect 12355 13550 12435 13590
rect 12475 13550 12555 13590
rect 12355 13465 12555 13550
rect 12705 13590 12905 13665
rect 12705 13550 12785 13590
rect 12825 13550 12905 13590
rect 12705 13465 12905 13550
rect 13055 13590 13255 13665
rect 13055 13550 13135 13590
rect 13175 13550 13255 13590
rect 13055 13465 13255 13550
rect 13405 13590 13605 13665
rect 13405 13550 13485 13590
rect 13525 13550 13605 13590
rect 13405 13465 13605 13550
rect 13755 13590 13955 13665
rect 13755 13550 13835 13590
rect 13875 13550 13955 13590
rect 13755 13465 13955 13550
rect 14105 13590 14305 13665
rect 14105 13550 14185 13590
rect 14225 13550 14305 13590
rect 14105 13465 14305 13550
rect 14455 13590 14655 13665
rect 14455 13550 14535 13590
rect 14575 13550 14655 13590
rect 14455 13465 14655 13550
rect -1245 13240 -1045 13315
rect -1245 13200 -1165 13240
rect -1125 13200 -1045 13240
rect -1245 13115 -1045 13200
rect -895 13240 -695 13315
rect -895 13200 -815 13240
rect -775 13200 -695 13240
rect -895 13115 -695 13200
rect -545 13240 -345 13315
rect -545 13200 -465 13240
rect -425 13200 -345 13240
rect -545 13115 -345 13200
rect -195 13240 5 13315
rect -195 13200 -115 13240
rect -75 13200 5 13240
rect -195 13115 5 13200
rect 155 13240 355 13315
rect 155 13200 235 13240
rect 275 13200 355 13240
rect 155 13115 355 13200
rect 505 13240 705 13315
rect 505 13200 585 13240
rect 625 13200 705 13240
rect 505 13115 705 13200
rect 855 13240 1055 13315
rect 855 13200 935 13240
rect 975 13200 1055 13240
rect 855 13115 1055 13200
rect 1205 13240 1405 13315
rect 1205 13200 1285 13240
rect 1325 13200 1405 13240
rect 1205 13115 1405 13200
rect 1555 13240 1755 13315
rect 1555 13200 1635 13240
rect 1675 13200 1755 13240
rect 1555 13115 1755 13200
rect 9555 13240 9755 13315
rect 9555 13200 9635 13240
rect 9675 13200 9755 13240
rect 9555 13115 9755 13200
rect 9905 13240 10105 13315
rect 9905 13200 9985 13240
rect 10025 13200 10105 13240
rect 9905 13115 10105 13200
rect 10255 13240 10455 13315
rect 10255 13200 10335 13240
rect 10375 13200 10455 13240
rect 10255 13115 10455 13200
rect 10605 13240 10805 13315
rect 10605 13200 10685 13240
rect 10725 13200 10805 13240
rect 10605 13115 10805 13200
rect 10955 13240 11155 13315
rect 10955 13200 11035 13240
rect 11075 13200 11155 13240
rect 10955 13115 11155 13200
rect 11305 13240 11505 13315
rect 11305 13200 11385 13240
rect 11425 13200 11505 13240
rect 11305 13115 11505 13200
rect 11655 13240 11855 13315
rect 11655 13200 11735 13240
rect 11775 13200 11855 13240
rect 11655 13115 11855 13200
rect 12005 13240 12205 13315
rect 12005 13200 12085 13240
rect 12125 13200 12205 13240
rect 12005 13115 12205 13200
rect 12355 13240 12555 13315
rect 12355 13200 12435 13240
rect 12475 13200 12555 13240
rect 12355 13115 12555 13200
rect 12705 13240 12905 13315
rect 12705 13200 12785 13240
rect 12825 13200 12905 13240
rect 12705 13115 12905 13200
rect 13055 13240 13255 13315
rect 13055 13200 13135 13240
rect 13175 13200 13255 13240
rect 13055 13115 13255 13200
rect 13405 13240 13605 13315
rect 13405 13200 13485 13240
rect 13525 13200 13605 13240
rect 13405 13115 13605 13200
rect 13755 13240 13955 13315
rect 13755 13200 13835 13240
rect 13875 13200 13955 13240
rect 13755 13115 13955 13200
rect 14105 13240 14305 13315
rect 14105 13200 14185 13240
rect 14225 13200 14305 13240
rect 14105 13115 14305 13200
rect 14455 13240 14655 13315
rect 14455 13200 14535 13240
rect 14575 13200 14655 13240
rect 14455 13115 14655 13200
rect -1245 12890 -1045 12965
rect -1245 12850 -1165 12890
rect -1125 12850 -1045 12890
rect -1245 12765 -1045 12850
rect -895 12890 -695 12965
rect -895 12850 -815 12890
rect -775 12850 -695 12890
rect -895 12765 -695 12850
rect -545 12890 -345 12965
rect -545 12850 -465 12890
rect -425 12850 -345 12890
rect -545 12765 -345 12850
rect -195 12890 5 12965
rect -195 12850 -115 12890
rect -75 12850 5 12890
rect -195 12765 5 12850
rect 155 12890 355 12965
rect 155 12850 235 12890
rect 275 12850 355 12890
rect 155 12765 355 12850
rect 505 12890 705 12965
rect 505 12850 585 12890
rect 625 12850 705 12890
rect 505 12765 705 12850
rect 855 12890 1055 12965
rect 855 12850 935 12890
rect 975 12850 1055 12890
rect 855 12765 1055 12850
rect 1205 12890 1405 12965
rect 1205 12850 1285 12890
rect 1325 12850 1405 12890
rect 1205 12765 1405 12850
rect 1555 12890 1755 12965
rect 1555 12850 1635 12890
rect 1675 12850 1755 12890
rect 1555 12765 1755 12850
rect 9555 12890 9755 12965
rect 9555 12850 9635 12890
rect 9675 12850 9755 12890
rect 9555 12765 9755 12850
rect 9905 12890 10105 12965
rect 9905 12850 9985 12890
rect 10025 12850 10105 12890
rect 9905 12765 10105 12850
rect 10255 12890 10455 12965
rect 10255 12850 10335 12890
rect 10375 12850 10455 12890
rect 10255 12765 10455 12850
rect 10605 12890 10805 12965
rect 10605 12850 10685 12890
rect 10725 12850 10805 12890
rect 10605 12765 10805 12850
rect 10955 12890 11155 12965
rect 10955 12850 11035 12890
rect 11075 12850 11155 12890
rect 10955 12765 11155 12850
rect 11305 12890 11505 12965
rect 11305 12850 11385 12890
rect 11425 12850 11505 12890
rect 11305 12765 11505 12850
rect 11655 12890 11855 12965
rect 11655 12850 11735 12890
rect 11775 12850 11855 12890
rect 11655 12765 11855 12850
rect 12005 12890 12205 12965
rect 12005 12850 12085 12890
rect 12125 12850 12205 12890
rect 12005 12765 12205 12850
rect 12355 12890 12555 12965
rect 12355 12850 12435 12890
rect 12475 12850 12555 12890
rect 12355 12765 12555 12850
rect 12705 12890 12905 12965
rect 12705 12850 12785 12890
rect 12825 12850 12905 12890
rect 12705 12765 12905 12850
rect 13055 12890 13255 12965
rect 13055 12850 13135 12890
rect 13175 12850 13255 12890
rect 13055 12765 13255 12850
rect 13405 12890 13605 12965
rect 13405 12850 13485 12890
rect 13525 12850 13605 12890
rect 13405 12765 13605 12850
rect 13755 12890 13955 12965
rect 13755 12850 13835 12890
rect 13875 12850 13955 12890
rect 13755 12765 13955 12850
rect 14105 12890 14305 12965
rect 14105 12850 14185 12890
rect 14225 12850 14305 12890
rect 14105 12765 14305 12850
rect 14455 12890 14655 12965
rect 14455 12850 14535 12890
rect 14575 12850 14655 12890
rect 14455 12765 14655 12850
rect -1245 12540 -1045 12615
rect -1245 12500 -1165 12540
rect -1125 12500 -1045 12540
rect -1245 12415 -1045 12500
rect -895 12540 -695 12615
rect -895 12500 -815 12540
rect -775 12500 -695 12540
rect -895 12415 -695 12500
rect -545 12540 -345 12615
rect -545 12500 -465 12540
rect -425 12500 -345 12540
rect -545 12415 -345 12500
rect -195 12540 5 12615
rect -195 12500 -115 12540
rect -75 12500 5 12540
rect -195 12415 5 12500
rect 155 12540 355 12615
rect 155 12500 235 12540
rect 275 12500 355 12540
rect 155 12415 355 12500
rect 505 12540 705 12615
rect 505 12500 585 12540
rect 625 12500 705 12540
rect 505 12415 705 12500
rect 855 12540 1055 12615
rect 855 12500 935 12540
rect 975 12500 1055 12540
rect 855 12415 1055 12500
rect 1205 12540 1405 12615
rect 1205 12500 1285 12540
rect 1325 12500 1405 12540
rect 1205 12415 1405 12500
rect 1555 12540 1755 12615
rect 1555 12500 1635 12540
rect 1675 12500 1755 12540
rect 1555 12415 1755 12500
rect 9555 12540 9755 12615
rect 9555 12500 9635 12540
rect 9675 12500 9755 12540
rect 9555 12415 9755 12500
rect 9905 12540 10105 12615
rect 9905 12500 9985 12540
rect 10025 12500 10105 12540
rect 9905 12415 10105 12500
rect 10255 12540 10455 12615
rect 10255 12500 10335 12540
rect 10375 12500 10455 12540
rect 10255 12415 10455 12500
rect 10605 12540 10805 12615
rect 10605 12500 10685 12540
rect 10725 12500 10805 12540
rect 10605 12415 10805 12500
rect 10955 12540 11155 12615
rect 10955 12500 11035 12540
rect 11075 12500 11155 12540
rect 10955 12415 11155 12500
rect 11305 12540 11505 12615
rect 11305 12500 11385 12540
rect 11425 12500 11505 12540
rect 11305 12415 11505 12500
rect 11655 12540 11855 12615
rect 11655 12500 11735 12540
rect 11775 12500 11855 12540
rect 11655 12415 11855 12500
rect 12005 12540 12205 12615
rect 12005 12500 12085 12540
rect 12125 12500 12205 12540
rect 12005 12415 12205 12500
rect 12355 12540 12555 12615
rect 12355 12500 12435 12540
rect 12475 12500 12555 12540
rect 12355 12415 12555 12500
rect 12705 12540 12905 12615
rect 12705 12500 12785 12540
rect 12825 12500 12905 12540
rect 12705 12415 12905 12500
rect 13055 12540 13255 12615
rect 13055 12500 13135 12540
rect 13175 12500 13255 12540
rect 13055 12415 13255 12500
rect 13405 12540 13605 12615
rect 13405 12500 13485 12540
rect 13525 12500 13605 12540
rect 13405 12415 13605 12500
rect 13755 12540 13955 12615
rect 13755 12500 13835 12540
rect 13875 12500 13955 12540
rect 13755 12415 13955 12500
rect 14105 12540 14305 12615
rect 14105 12500 14185 12540
rect 14225 12500 14305 12540
rect 14105 12415 14305 12500
rect 14455 12540 14655 12615
rect 14455 12500 14535 12540
rect 14575 12500 14655 12540
rect 14455 12415 14655 12500
rect -1245 12190 -1045 12265
rect -1245 12150 -1165 12190
rect -1125 12150 -1045 12190
rect -1245 12065 -1045 12150
rect -895 12190 -695 12265
rect -895 12150 -815 12190
rect -775 12150 -695 12190
rect -895 12065 -695 12150
rect -545 12190 -345 12265
rect -545 12150 -465 12190
rect -425 12150 -345 12190
rect -545 12065 -345 12150
rect -195 12190 5 12265
rect -195 12150 -115 12190
rect -75 12150 5 12190
rect -195 12065 5 12150
rect 155 12190 355 12265
rect 155 12150 235 12190
rect 275 12150 355 12190
rect 155 12065 355 12150
rect 505 12190 705 12265
rect 505 12150 585 12190
rect 625 12150 705 12190
rect 505 12065 705 12150
rect 855 12190 1055 12265
rect 855 12150 935 12190
rect 975 12150 1055 12190
rect 855 12065 1055 12150
rect 1205 12190 1405 12265
rect 1205 12150 1285 12190
rect 1325 12150 1405 12190
rect 1205 12065 1405 12150
rect 1555 12190 1755 12265
rect 1555 12150 1635 12190
rect 1675 12150 1755 12190
rect 1555 12065 1755 12150
rect 9555 12190 9755 12265
rect 9555 12150 9635 12190
rect 9675 12150 9755 12190
rect 9555 12065 9755 12150
rect 9905 12190 10105 12265
rect 9905 12150 9985 12190
rect 10025 12150 10105 12190
rect 9905 12065 10105 12150
rect 10255 12190 10455 12265
rect 10255 12150 10335 12190
rect 10375 12150 10455 12190
rect 10255 12065 10455 12150
rect 10605 12190 10805 12265
rect 10605 12150 10685 12190
rect 10725 12150 10805 12190
rect 10605 12065 10805 12150
rect 10955 12190 11155 12265
rect 10955 12150 11035 12190
rect 11075 12150 11155 12190
rect 10955 12065 11155 12150
rect 11305 12190 11505 12265
rect 11305 12150 11385 12190
rect 11425 12150 11505 12190
rect 11305 12065 11505 12150
rect 11655 12190 11855 12265
rect 11655 12150 11735 12190
rect 11775 12150 11855 12190
rect 11655 12065 11855 12150
rect 12005 12190 12205 12265
rect 12005 12150 12085 12190
rect 12125 12150 12205 12190
rect 12005 12065 12205 12150
rect 12355 12190 12555 12265
rect 12355 12150 12435 12190
rect 12475 12150 12555 12190
rect 12355 12065 12555 12150
rect 12705 12190 12905 12265
rect 12705 12150 12785 12190
rect 12825 12150 12905 12190
rect 12705 12065 12905 12150
rect 13055 12190 13255 12265
rect 13055 12150 13135 12190
rect 13175 12150 13255 12190
rect 13055 12065 13255 12150
rect 13405 12190 13605 12265
rect 13405 12150 13485 12190
rect 13525 12150 13605 12190
rect 13405 12065 13605 12150
rect 13755 12190 13955 12265
rect 13755 12150 13835 12190
rect 13875 12150 13955 12190
rect 13755 12065 13955 12150
rect 14105 12190 14305 12265
rect 14105 12150 14185 12190
rect 14225 12150 14305 12190
rect 14105 12065 14305 12150
rect 14455 12190 14655 12265
rect 14455 12150 14535 12190
rect 14575 12150 14655 12190
rect 14455 12065 14655 12150
rect -1245 11840 -1045 11915
rect -1245 11800 -1165 11840
rect -1125 11800 -1045 11840
rect -1245 11715 -1045 11800
rect -895 11840 -695 11915
rect -895 11800 -815 11840
rect -775 11800 -695 11840
rect -895 11715 -695 11800
rect -545 11840 -345 11915
rect -545 11800 -465 11840
rect -425 11800 -345 11840
rect -545 11715 -345 11800
rect -195 11840 5 11915
rect -195 11800 -115 11840
rect -75 11800 5 11840
rect -195 11715 5 11800
rect 155 11840 355 11915
rect 155 11800 235 11840
rect 275 11800 355 11840
rect 155 11715 355 11800
rect 505 11840 705 11915
rect 505 11800 585 11840
rect 625 11800 705 11840
rect 505 11715 705 11800
rect 855 11840 1055 11915
rect 855 11800 935 11840
rect 975 11800 1055 11840
rect 855 11715 1055 11800
rect 1205 11840 1405 11915
rect 1205 11800 1285 11840
rect 1325 11800 1405 11840
rect 1205 11715 1405 11800
rect 1555 11840 1755 11915
rect 1555 11800 1635 11840
rect 1675 11800 1755 11840
rect 1555 11715 1755 11800
rect 9555 11840 9755 11915
rect 9555 11800 9635 11840
rect 9675 11800 9755 11840
rect 9555 11715 9755 11800
rect 9905 11840 10105 11915
rect 9905 11800 9985 11840
rect 10025 11800 10105 11840
rect 9905 11715 10105 11800
rect 10255 11840 10455 11915
rect 10255 11800 10335 11840
rect 10375 11800 10455 11840
rect 10255 11715 10455 11800
rect 10605 11840 10805 11915
rect 10605 11800 10685 11840
rect 10725 11800 10805 11840
rect 10605 11715 10805 11800
rect 10955 11840 11155 11915
rect 10955 11800 11035 11840
rect 11075 11800 11155 11840
rect 10955 11715 11155 11800
rect 11305 11840 11505 11915
rect 11305 11800 11385 11840
rect 11425 11800 11505 11840
rect 11305 11715 11505 11800
rect 11655 11840 11855 11915
rect 11655 11800 11735 11840
rect 11775 11800 11855 11840
rect 11655 11715 11855 11800
rect 12005 11840 12205 11915
rect 12005 11800 12085 11840
rect 12125 11800 12205 11840
rect 12005 11715 12205 11800
rect 12355 11840 12555 11915
rect 12355 11800 12435 11840
rect 12475 11800 12555 11840
rect 12355 11715 12555 11800
rect 12705 11840 12905 11915
rect 12705 11800 12785 11840
rect 12825 11800 12905 11840
rect 12705 11715 12905 11800
rect 13055 11840 13255 11915
rect 13055 11800 13135 11840
rect 13175 11800 13255 11840
rect 13055 11715 13255 11800
rect 13405 11840 13605 11915
rect 13405 11800 13485 11840
rect 13525 11800 13605 11840
rect 13405 11715 13605 11800
rect 13755 11840 13955 11915
rect 13755 11800 13835 11840
rect 13875 11800 13955 11840
rect 13755 11715 13955 11800
rect 14105 11840 14305 11915
rect 14105 11800 14185 11840
rect 14225 11800 14305 11840
rect 14105 11715 14305 11800
rect 14455 11840 14655 11915
rect 14455 11800 14535 11840
rect 14575 11800 14655 11840
rect 14455 11715 14655 11800
rect -1245 11490 -1045 11565
rect -1245 11450 -1165 11490
rect -1125 11450 -1045 11490
rect -1245 11365 -1045 11450
rect -895 11490 -695 11565
rect -895 11450 -815 11490
rect -775 11450 -695 11490
rect -895 11365 -695 11450
rect -545 11490 -345 11565
rect -545 11450 -465 11490
rect -425 11450 -345 11490
rect -545 11365 -345 11450
rect -195 11490 5 11565
rect -195 11450 -115 11490
rect -75 11450 5 11490
rect -195 11365 5 11450
rect 155 11490 355 11565
rect 155 11450 235 11490
rect 275 11450 355 11490
rect 155 11365 355 11450
rect 505 11490 705 11565
rect 505 11450 585 11490
rect 625 11450 705 11490
rect 505 11365 705 11450
rect 855 11490 1055 11565
rect 855 11450 935 11490
rect 975 11450 1055 11490
rect 855 11365 1055 11450
rect 1205 11490 1405 11565
rect 1205 11450 1285 11490
rect 1325 11450 1405 11490
rect 1205 11365 1405 11450
rect 1555 11490 1755 11565
rect 1555 11450 1635 11490
rect 1675 11450 1755 11490
rect 1555 11365 1755 11450
rect 9555 11490 9755 11565
rect 9555 11450 9635 11490
rect 9675 11450 9755 11490
rect 9555 11365 9755 11450
rect 9905 11490 10105 11565
rect 9905 11450 9985 11490
rect 10025 11450 10105 11490
rect 9905 11365 10105 11450
rect 10255 11490 10455 11565
rect 10255 11450 10335 11490
rect 10375 11450 10455 11490
rect 10255 11365 10455 11450
rect 10605 11490 10805 11565
rect 10605 11450 10685 11490
rect 10725 11450 10805 11490
rect 10605 11365 10805 11450
rect 10955 11490 11155 11565
rect 10955 11450 11035 11490
rect 11075 11450 11155 11490
rect 10955 11365 11155 11450
rect 11305 11490 11505 11565
rect 11305 11450 11385 11490
rect 11425 11450 11505 11490
rect 11305 11365 11505 11450
rect 11655 11490 11855 11565
rect 11655 11450 11735 11490
rect 11775 11450 11855 11490
rect 11655 11365 11855 11450
rect 12005 11490 12205 11565
rect 12005 11450 12085 11490
rect 12125 11450 12205 11490
rect 12005 11365 12205 11450
rect 12355 11490 12555 11565
rect 12355 11450 12435 11490
rect 12475 11450 12555 11490
rect 12355 11365 12555 11450
rect 12705 11490 12905 11565
rect 12705 11450 12785 11490
rect 12825 11450 12905 11490
rect 12705 11365 12905 11450
rect 13055 11490 13255 11565
rect 13055 11450 13135 11490
rect 13175 11450 13255 11490
rect 13055 11365 13255 11450
rect 13405 11490 13605 11565
rect 13405 11450 13485 11490
rect 13525 11450 13605 11490
rect 13405 11365 13605 11450
rect 13755 11490 13955 11565
rect 13755 11450 13835 11490
rect 13875 11450 13955 11490
rect 13755 11365 13955 11450
rect 14105 11490 14305 11565
rect 14105 11450 14185 11490
rect 14225 11450 14305 11490
rect 14105 11365 14305 11450
rect 14455 11490 14655 11565
rect 14455 11450 14535 11490
rect 14575 11450 14655 11490
rect 14455 11365 14655 11450
rect -1245 11140 -1045 11215
rect -1245 11100 -1165 11140
rect -1125 11100 -1045 11140
rect -1245 11015 -1045 11100
rect -895 11140 -695 11215
rect -895 11100 -815 11140
rect -775 11100 -695 11140
rect -895 11015 -695 11100
rect -545 11140 -345 11215
rect -545 11100 -465 11140
rect -425 11100 -345 11140
rect -545 11015 -345 11100
rect -195 11140 5 11215
rect -195 11100 -115 11140
rect -75 11100 5 11140
rect -195 11015 5 11100
rect 155 11140 355 11215
rect 155 11100 235 11140
rect 275 11100 355 11140
rect 155 11015 355 11100
rect 505 11140 705 11215
rect 505 11100 585 11140
rect 625 11100 705 11140
rect 505 11015 705 11100
rect 855 11140 1055 11215
rect 855 11100 935 11140
rect 975 11100 1055 11140
rect 855 11015 1055 11100
rect 1205 11140 1405 11215
rect 1205 11100 1285 11140
rect 1325 11100 1405 11140
rect 1205 11015 1405 11100
rect 1555 11140 1755 11215
rect 1555 11100 1635 11140
rect 1675 11100 1755 11140
rect 1555 11015 1755 11100
rect 9555 11140 9755 11215
rect 9555 11100 9635 11140
rect 9675 11100 9755 11140
rect 9555 11015 9755 11100
rect 9905 11140 10105 11215
rect 9905 11100 9985 11140
rect 10025 11100 10105 11140
rect 9905 11015 10105 11100
rect 10255 11140 10455 11215
rect 10255 11100 10335 11140
rect 10375 11100 10455 11140
rect 10255 11015 10455 11100
rect 10605 11140 10805 11215
rect 10605 11100 10685 11140
rect 10725 11100 10805 11140
rect 10605 11015 10805 11100
rect 10955 11140 11155 11215
rect 10955 11100 11035 11140
rect 11075 11100 11155 11140
rect 10955 11015 11155 11100
rect 11305 11140 11505 11215
rect 11305 11100 11385 11140
rect 11425 11100 11505 11140
rect 11305 11015 11505 11100
rect 11655 11140 11855 11215
rect 11655 11100 11735 11140
rect 11775 11100 11855 11140
rect 11655 11015 11855 11100
rect 12005 11140 12205 11215
rect 12005 11100 12085 11140
rect 12125 11100 12205 11140
rect 12005 11015 12205 11100
rect 12355 11140 12555 11215
rect 12355 11100 12435 11140
rect 12475 11100 12555 11140
rect 12355 11015 12555 11100
rect 12705 11140 12905 11215
rect 12705 11100 12785 11140
rect 12825 11100 12905 11140
rect 12705 11015 12905 11100
rect 13055 11140 13255 11215
rect 13055 11100 13135 11140
rect 13175 11100 13255 11140
rect 13055 11015 13255 11100
rect 13405 11140 13605 11215
rect 13405 11100 13485 11140
rect 13525 11100 13605 11140
rect 13405 11015 13605 11100
rect 13755 11140 13955 11215
rect 13755 11100 13835 11140
rect 13875 11100 13955 11140
rect 13755 11015 13955 11100
rect 14105 11140 14305 11215
rect 14105 11100 14185 11140
rect 14225 11100 14305 11140
rect 14105 11015 14305 11100
rect 14455 11140 14655 11215
rect 14455 11100 14535 11140
rect 14575 11100 14655 11140
rect 14455 11015 14655 11100
rect -1245 10790 -1045 10865
rect -1245 10750 -1165 10790
rect -1125 10750 -1045 10790
rect -1245 10665 -1045 10750
rect -895 10790 -695 10865
rect -895 10750 -815 10790
rect -775 10750 -695 10790
rect -895 10665 -695 10750
rect -545 10790 -345 10865
rect -545 10750 -465 10790
rect -425 10750 -345 10790
rect -545 10665 -345 10750
rect -195 10790 5 10865
rect -195 10750 -115 10790
rect -75 10750 5 10790
rect -195 10665 5 10750
rect 155 10790 355 10865
rect 155 10750 235 10790
rect 275 10750 355 10790
rect 155 10665 355 10750
rect 505 10790 705 10865
rect 505 10750 585 10790
rect 625 10750 705 10790
rect 505 10665 705 10750
rect 855 10790 1055 10865
rect 855 10750 935 10790
rect 975 10750 1055 10790
rect 855 10665 1055 10750
rect 1205 10790 1405 10865
rect 1205 10750 1285 10790
rect 1325 10750 1405 10790
rect 1205 10665 1405 10750
rect 1555 10790 1755 10865
rect 1555 10750 1635 10790
rect 1675 10750 1755 10790
rect 1555 10665 1755 10750
rect 9555 10790 9755 10865
rect 9555 10750 9635 10790
rect 9675 10750 9755 10790
rect 9555 10665 9755 10750
rect 9905 10790 10105 10865
rect 9905 10750 9985 10790
rect 10025 10750 10105 10790
rect 9905 10665 10105 10750
rect 10255 10790 10455 10865
rect 10255 10750 10335 10790
rect 10375 10750 10455 10790
rect 10255 10665 10455 10750
rect 10605 10790 10805 10865
rect 10605 10750 10685 10790
rect 10725 10750 10805 10790
rect 10605 10665 10805 10750
rect 10955 10790 11155 10865
rect 10955 10750 11035 10790
rect 11075 10750 11155 10790
rect 10955 10665 11155 10750
rect 11305 10790 11505 10865
rect 11305 10750 11385 10790
rect 11425 10750 11505 10790
rect 11305 10665 11505 10750
rect 11655 10790 11855 10865
rect 11655 10750 11735 10790
rect 11775 10750 11855 10790
rect 11655 10665 11855 10750
rect 12005 10790 12205 10865
rect 12005 10750 12085 10790
rect 12125 10750 12205 10790
rect 12005 10665 12205 10750
rect 12355 10790 12555 10865
rect 12355 10750 12435 10790
rect 12475 10750 12555 10790
rect 12355 10665 12555 10750
rect 12705 10790 12905 10865
rect 12705 10750 12785 10790
rect 12825 10750 12905 10790
rect 12705 10665 12905 10750
rect 13055 10790 13255 10865
rect 13055 10750 13135 10790
rect 13175 10750 13255 10790
rect 13055 10665 13255 10750
rect 13405 10790 13605 10865
rect 13405 10750 13485 10790
rect 13525 10750 13605 10790
rect 13405 10665 13605 10750
rect 13755 10790 13955 10865
rect 13755 10750 13835 10790
rect 13875 10750 13955 10790
rect 13755 10665 13955 10750
rect 14105 10790 14305 10865
rect 14105 10750 14185 10790
rect 14225 10750 14305 10790
rect 14105 10665 14305 10750
rect 14455 10790 14655 10865
rect 14455 10750 14535 10790
rect 14575 10750 14655 10790
rect 14455 10665 14655 10750
rect -1245 10440 -1045 10515
rect -1245 10400 -1165 10440
rect -1125 10400 -1045 10440
rect -1245 10315 -1045 10400
rect -895 10440 -695 10515
rect -895 10400 -815 10440
rect -775 10400 -695 10440
rect -895 10315 -695 10400
rect -545 10440 -345 10515
rect -545 10400 -465 10440
rect -425 10400 -345 10440
rect -545 10315 -345 10400
rect -195 10440 5 10515
rect -195 10400 -115 10440
rect -75 10400 5 10440
rect -195 10315 5 10400
rect 155 10440 355 10515
rect 155 10400 235 10440
rect 275 10400 355 10440
rect 155 10315 355 10400
rect 505 10440 705 10515
rect 505 10400 585 10440
rect 625 10400 705 10440
rect 505 10315 705 10400
rect 855 10440 1055 10515
rect 855 10400 935 10440
rect 975 10400 1055 10440
rect 855 10315 1055 10400
rect 1205 10440 1405 10515
rect 1205 10400 1285 10440
rect 1325 10400 1405 10440
rect 1205 10315 1405 10400
rect 1555 10440 1755 10515
rect 1555 10400 1635 10440
rect 1675 10400 1755 10440
rect 1555 10315 1755 10400
rect 9555 10440 9755 10515
rect 9555 10400 9635 10440
rect 9675 10400 9755 10440
rect 9555 10315 9755 10400
rect 9905 10440 10105 10515
rect 9905 10400 9985 10440
rect 10025 10400 10105 10440
rect 9905 10315 10105 10400
rect 10255 10440 10455 10515
rect 10255 10400 10335 10440
rect 10375 10400 10455 10440
rect 10255 10315 10455 10400
rect 10605 10440 10805 10515
rect 10605 10400 10685 10440
rect 10725 10400 10805 10440
rect 10605 10315 10805 10400
rect 10955 10440 11155 10515
rect 10955 10400 11035 10440
rect 11075 10400 11155 10440
rect 10955 10315 11155 10400
rect 11305 10440 11505 10515
rect 11305 10400 11385 10440
rect 11425 10400 11505 10440
rect 11305 10315 11505 10400
rect 11655 10440 11855 10515
rect 11655 10400 11735 10440
rect 11775 10400 11855 10440
rect 11655 10315 11855 10400
rect 12005 10440 12205 10515
rect 12005 10400 12085 10440
rect 12125 10400 12205 10440
rect 12005 10315 12205 10400
rect 12355 10440 12555 10515
rect 12355 10400 12435 10440
rect 12475 10400 12555 10440
rect 12355 10315 12555 10400
rect 12705 10440 12905 10515
rect 12705 10400 12785 10440
rect 12825 10400 12905 10440
rect 12705 10315 12905 10400
rect 13055 10440 13255 10515
rect 13055 10400 13135 10440
rect 13175 10400 13255 10440
rect 13055 10315 13255 10400
rect 13405 10440 13605 10515
rect 13405 10400 13485 10440
rect 13525 10400 13605 10440
rect 13405 10315 13605 10400
rect 13755 10440 13955 10515
rect 13755 10400 13835 10440
rect 13875 10400 13955 10440
rect 13755 10315 13955 10400
rect 14105 10440 14305 10515
rect 14105 10400 14185 10440
rect 14225 10400 14305 10440
rect 14105 10315 14305 10400
rect 14455 10440 14655 10515
rect 14455 10400 14535 10440
rect 14575 10400 14655 10440
rect 14455 10315 14655 10400
rect -1245 10090 -1045 10165
rect -1245 10050 -1165 10090
rect -1125 10050 -1045 10090
rect -1245 9965 -1045 10050
rect -895 10090 -695 10165
rect -895 10050 -815 10090
rect -775 10050 -695 10090
rect -895 9965 -695 10050
rect -545 10090 -345 10165
rect -545 10050 -465 10090
rect -425 10050 -345 10090
rect -545 9965 -345 10050
rect -195 10090 5 10165
rect -195 10050 -115 10090
rect -75 10050 5 10090
rect -195 9965 5 10050
rect 155 10090 355 10165
rect 155 10050 235 10090
rect 275 10050 355 10090
rect 155 9965 355 10050
rect 505 10090 705 10165
rect 505 10050 585 10090
rect 625 10050 705 10090
rect 505 9965 705 10050
rect 855 10090 1055 10165
rect 855 10050 935 10090
rect 975 10050 1055 10090
rect 855 9965 1055 10050
rect 1205 10090 1405 10165
rect 1205 10050 1285 10090
rect 1325 10050 1405 10090
rect 1205 9965 1405 10050
rect 1555 10090 1755 10165
rect 1555 10050 1635 10090
rect 1675 10050 1755 10090
rect 1555 9965 1755 10050
rect 9555 10090 9755 10165
rect 9555 10050 9635 10090
rect 9675 10050 9755 10090
rect 9555 9965 9755 10050
rect 9905 10090 10105 10165
rect 9905 10050 9985 10090
rect 10025 10050 10105 10090
rect 9905 9965 10105 10050
rect 10255 10090 10455 10165
rect 10255 10050 10335 10090
rect 10375 10050 10455 10090
rect 10255 9965 10455 10050
rect 10605 10090 10805 10165
rect 10605 10050 10685 10090
rect 10725 10050 10805 10090
rect 10605 9965 10805 10050
rect 10955 10090 11155 10165
rect 10955 10050 11035 10090
rect 11075 10050 11155 10090
rect 10955 9965 11155 10050
rect 11305 10090 11505 10165
rect 11305 10050 11385 10090
rect 11425 10050 11505 10090
rect 11305 9965 11505 10050
rect 11655 10090 11855 10165
rect 11655 10050 11735 10090
rect 11775 10050 11855 10090
rect 11655 9965 11855 10050
rect 12005 10090 12205 10165
rect 12005 10050 12085 10090
rect 12125 10050 12205 10090
rect 12005 9965 12205 10050
rect 12355 10090 12555 10165
rect 12355 10050 12435 10090
rect 12475 10050 12555 10090
rect 12355 9965 12555 10050
rect 12705 10090 12905 10165
rect 12705 10050 12785 10090
rect 12825 10050 12905 10090
rect 12705 9965 12905 10050
rect 13055 10090 13255 10165
rect 13055 10050 13135 10090
rect 13175 10050 13255 10090
rect 13055 9965 13255 10050
rect 13405 10090 13605 10165
rect 13405 10050 13485 10090
rect 13525 10050 13605 10090
rect 13405 9965 13605 10050
rect 13755 10090 13955 10165
rect 13755 10050 13835 10090
rect 13875 10050 13955 10090
rect 13755 9965 13955 10050
rect 14105 10090 14305 10165
rect 14105 10050 14185 10090
rect 14225 10050 14305 10090
rect 14105 9965 14305 10050
rect 14455 10090 14655 10165
rect 14455 10050 14535 10090
rect 14575 10050 14655 10090
rect 14455 9965 14655 10050
rect 9555 9740 9755 9815
rect 9555 9700 9635 9740
rect 9675 9700 9755 9740
rect 9555 9615 9755 9700
rect 9905 9740 10105 9815
rect 9905 9700 9985 9740
rect 10025 9700 10105 9740
rect 9905 9615 10105 9700
rect 10255 9740 10455 9815
rect 10255 9700 10335 9740
rect 10375 9700 10455 9740
rect 10255 9615 10455 9700
rect 10605 9740 10805 9815
rect 10605 9700 10685 9740
rect 10725 9700 10805 9740
rect 10605 9615 10805 9700
rect 10955 9740 11155 9815
rect 10955 9700 11035 9740
rect 11075 9700 11155 9740
rect 10955 9615 11155 9700
rect 11305 9740 11505 9815
rect 11305 9700 11385 9740
rect 11425 9700 11505 9740
rect 11305 9615 11505 9700
rect 11655 9740 11855 9815
rect 11655 9700 11735 9740
rect 11775 9700 11855 9740
rect 11655 9615 11855 9700
rect 12005 9740 12205 9815
rect 12005 9700 12085 9740
rect 12125 9700 12205 9740
rect 12005 9615 12205 9700
rect 12355 9740 12555 9815
rect 12355 9700 12435 9740
rect 12475 9700 12555 9740
rect 12355 9615 12555 9700
rect 12705 9740 12905 9815
rect 12705 9700 12785 9740
rect 12825 9700 12905 9740
rect 12705 9615 12905 9700
rect 13055 9740 13255 9815
rect 13055 9700 13135 9740
rect 13175 9700 13255 9740
rect 13055 9615 13255 9700
rect 13405 9740 13605 9815
rect 13405 9700 13485 9740
rect 13525 9700 13605 9740
rect 13405 9615 13605 9700
rect 13755 9740 13955 9815
rect 13755 9700 13835 9740
rect 13875 9700 13955 9740
rect 13755 9615 13955 9700
rect 14105 9740 14305 9815
rect 14105 9700 14185 9740
rect 14225 9700 14305 9740
rect 14105 9615 14305 9700
rect 14455 9740 14655 9815
rect 14455 9700 14535 9740
rect 14575 9700 14655 9740
rect 14455 9615 14655 9700
rect 9555 9390 9755 9465
rect 9555 9350 9635 9390
rect 9675 9350 9755 9390
rect 9555 9265 9755 9350
rect 9905 9390 10105 9465
rect 9905 9350 9985 9390
rect 10025 9350 10105 9390
rect 9905 9265 10105 9350
rect 10255 9390 10455 9465
rect 10255 9350 10335 9390
rect 10375 9350 10455 9390
rect 10255 9265 10455 9350
rect 10605 9390 10805 9465
rect 10605 9350 10685 9390
rect 10725 9350 10805 9390
rect 10605 9265 10805 9350
rect 10955 9390 11155 9465
rect 10955 9350 11035 9390
rect 11075 9350 11155 9390
rect 10955 9265 11155 9350
rect 11305 9390 11505 9465
rect 11305 9350 11385 9390
rect 11425 9350 11505 9390
rect 11305 9265 11505 9350
rect 11655 9390 11855 9465
rect 11655 9350 11735 9390
rect 11775 9350 11855 9390
rect 11655 9265 11855 9350
rect 12005 9390 12205 9465
rect 12005 9350 12085 9390
rect 12125 9350 12205 9390
rect 12005 9265 12205 9350
rect 12355 9390 12555 9465
rect 12355 9350 12435 9390
rect 12475 9350 12555 9390
rect 12355 9265 12555 9350
rect 12705 9390 12905 9465
rect 12705 9350 12785 9390
rect 12825 9350 12905 9390
rect 12705 9265 12905 9350
rect 13055 9390 13255 9465
rect 13055 9350 13135 9390
rect 13175 9350 13255 9390
rect 13055 9265 13255 9350
rect 13405 9390 13605 9465
rect 13405 9350 13485 9390
rect 13525 9350 13605 9390
rect 13405 9265 13605 9350
rect 13755 9390 13955 9465
rect 13755 9350 13835 9390
rect 13875 9350 13955 9390
rect 13755 9265 13955 9350
rect 14105 9390 14305 9465
rect 14105 9350 14185 9390
rect 14225 9350 14305 9390
rect 14105 9265 14305 9350
rect 14455 9390 14655 9465
rect 14455 9350 14535 9390
rect 14575 9350 14655 9390
rect 14455 9265 14655 9350
rect 9555 9040 9755 9115
rect 9555 9000 9635 9040
rect 9675 9000 9755 9040
rect 9555 8915 9755 9000
rect 9905 9040 10105 9115
rect 9905 9000 9985 9040
rect 10025 9000 10105 9040
rect 9905 8915 10105 9000
rect 10255 9040 10455 9115
rect 10255 9000 10335 9040
rect 10375 9000 10455 9040
rect 10255 8915 10455 9000
rect 10605 9040 10805 9115
rect 10605 9000 10685 9040
rect 10725 9000 10805 9040
rect 10605 8915 10805 9000
rect 10955 9040 11155 9115
rect 10955 9000 11035 9040
rect 11075 9000 11155 9040
rect 10955 8915 11155 9000
rect 11305 9040 11505 9115
rect 11305 9000 11385 9040
rect 11425 9000 11505 9040
rect 11305 8915 11505 9000
rect 11655 9040 11855 9115
rect 11655 9000 11735 9040
rect 11775 9000 11855 9040
rect 11655 8915 11855 9000
rect 12005 9040 12205 9115
rect 12005 9000 12085 9040
rect 12125 9000 12205 9040
rect 12005 8915 12205 9000
rect 12355 9040 12555 9115
rect 12355 9000 12435 9040
rect 12475 9000 12555 9040
rect 12355 8915 12555 9000
rect 12705 9040 12905 9115
rect 12705 9000 12785 9040
rect 12825 9000 12905 9040
rect 12705 8915 12905 9000
rect 13055 9040 13255 9115
rect 13055 9000 13135 9040
rect 13175 9000 13255 9040
rect 13055 8915 13255 9000
rect 13405 9040 13605 9115
rect 13405 9000 13485 9040
rect 13525 9000 13605 9040
rect 13405 8915 13605 9000
rect 13755 9040 13955 9115
rect 13755 9000 13835 9040
rect 13875 9000 13955 9040
rect 13755 8915 13955 9000
rect 14105 9040 14305 9115
rect 14105 9000 14185 9040
rect 14225 9000 14305 9040
rect 14105 8915 14305 9000
rect 14455 9040 14655 9115
rect 14455 9000 14535 9040
rect 14575 9000 14655 9040
rect 14455 8915 14655 9000
rect 9555 8690 9755 8765
rect 9555 8650 9635 8690
rect 9675 8650 9755 8690
rect 9555 8565 9755 8650
rect 9905 8690 10105 8765
rect 9905 8650 9985 8690
rect 10025 8650 10105 8690
rect 9905 8565 10105 8650
rect 10255 8690 10455 8765
rect 10255 8650 10335 8690
rect 10375 8650 10455 8690
rect 10255 8565 10455 8650
rect 10605 8690 10805 8765
rect 10605 8650 10685 8690
rect 10725 8650 10805 8690
rect 10605 8565 10805 8650
rect 10955 8690 11155 8765
rect 10955 8650 11035 8690
rect 11075 8650 11155 8690
rect 10955 8565 11155 8650
rect 11305 8690 11505 8765
rect 11305 8650 11385 8690
rect 11425 8650 11505 8690
rect 11305 8565 11505 8650
rect 11655 8690 11855 8765
rect 11655 8650 11735 8690
rect 11775 8650 11855 8690
rect 11655 8565 11855 8650
rect 12005 8690 12205 8765
rect 12005 8650 12085 8690
rect 12125 8650 12205 8690
rect 12005 8565 12205 8650
rect 12355 8690 12555 8765
rect 12355 8650 12435 8690
rect 12475 8650 12555 8690
rect 12355 8565 12555 8650
rect 12705 8690 12905 8765
rect 12705 8650 12785 8690
rect 12825 8650 12905 8690
rect 12705 8565 12905 8650
rect 13055 8690 13255 8765
rect 13055 8650 13135 8690
rect 13175 8650 13255 8690
rect 13055 8565 13255 8650
rect 13405 8690 13605 8765
rect 13405 8650 13485 8690
rect 13525 8650 13605 8690
rect 13405 8565 13605 8650
rect 13755 8690 13955 8765
rect 13755 8650 13835 8690
rect 13875 8650 13955 8690
rect 13755 8565 13955 8650
rect 14105 8690 14305 8765
rect 14105 8650 14185 8690
rect 14225 8650 14305 8690
rect 14105 8565 14305 8650
rect 14455 8690 14655 8765
rect 14455 8650 14535 8690
rect 14575 8650 14655 8690
rect 14455 8565 14655 8650
rect 9555 8340 9755 8415
rect 9555 8300 9635 8340
rect 9675 8300 9755 8340
rect 9555 8215 9755 8300
rect 9905 8340 10105 8415
rect 9905 8300 9985 8340
rect 10025 8300 10105 8340
rect 9905 8215 10105 8300
rect 10255 8340 10455 8415
rect 10255 8300 10335 8340
rect 10375 8300 10455 8340
rect 10255 8215 10455 8300
rect 10605 8340 10805 8415
rect 10605 8300 10685 8340
rect 10725 8300 10805 8340
rect 10605 8215 10805 8300
rect 10955 8340 11155 8415
rect 10955 8300 11035 8340
rect 11075 8300 11155 8340
rect 10955 8215 11155 8300
rect 11305 8340 11505 8415
rect 11305 8300 11385 8340
rect 11425 8300 11505 8340
rect 11305 8215 11505 8300
rect 11655 8340 11855 8415
rect 11655 8300 11735 8340
rect 11775 8300 11855 8340
rect 11655 8215 11855 8300
rect 12005 8340 12205 8415
rect 12005 8300 12085 8340
rect 12125 8300 12205 8340
rect 12005 8215 12205 8300
rect 12355 8340 12555 8415
rect 12355 8300 12435 8340
rect 12475 8300 12555 8340
rect 12355 8215 12555 8300
rect 12705 8340 12905 8415
rect 12705 8300 12785 8340
rect 12825 8300 12905 8340
rect 12705 8215 12905 8300
rect 13055 8340 13255 8415
rect 13055 8300 13135 8340
rect 13175 8300 13255 8340
rect 13055 8215 13255 8300
rect 13405 8340 13605 8415
rect 13405 8300 13485 8340
rect 13525 8300 13605 8340
rect 13405 8215 13605 8300
rect 13755 8340 13955 8415
rect 13755 8300 13835 8340
rect 13875 8300 13955 8340
rect 13755 8215 13955 8300
rect 14105 8340 14305 8415
rect 14105 8300 14185 8340
rect 14225 8300 14305 8340
rect 14105 8215 14305 8300
rect 14455 8340 14655 8415
rect 14455 8300 14535 8340
rect 14575 8300 14655 8340
rect 14455 8215 14655 8300
rect 9555 7990 9755 8065
rect 9555 7950 9635 7990
rect 9675 7950 9755 7990
rect 9555 7865 9755 7950
rect 9905 7990 10105 8065
rect 9905 7950 9985 7990
rect 10025 7950 10105 7990
rect 9905 7865 10105 7950
rect 10255 7990 10455 8065
rect 10255 7950 10335 7990
rect 10375 7950 10455 7990
rect 10255 7865 10455 7950
rect 10605 7990 10805 8065
rect 10605 7950 10685 7990
rect 10725 7950 10805 7990
rect 10605 7865 10805 7950
rect 10955 7990 11155 8065
rect 10955 7950 11035 7990
rect 11075 7950 11155 7990
rect 10955 7865 11155 7950
rect 11305 7990 11505 8065
rect 11305 7950 11385 7990
rect 11425 7950 11505 7990
rect 11305 7865 11505 7950
rect 11655 7990 11855 8065
rect 11655 7950 11735 7990
rect 11775 7950 11855 7990
rect 11655 7865 11855 7950
rect 12005 7990 12205 8065
rect 12005 7950 12085 7990
rect 12125 7950 12205 7990
rect 12005 7865 12205 7950
rect 12355 7990 12555 8065
rect 12355 7950 12435 7990
rect 12475 7950 12555 7990
rect 12355 7865 12555 7950
rect 12705 7990 12905 8065
rect 12705 7950 12785 7990
rect 12825 7950 12905 7990
rect 12705 7865 12905 7950
rect 13055 7990 13255 8065
rect 13055 7950 13135 7990
rect 13175 7950 13255 7990
rect 13055 7865 13255 7950
rect 13405 7990 13605 8065
rect 13405 7950 13485 7990
rect 13525 7950 13605 7990
rect 13405 7865 13605 7950
rect 13755 7990 13955 8065
rect 13755 7950 13835 7990
rect 13875 7950 13955 7990
rect 13755 7865 13955 7950
rect 14105 7990 14305 8065
rect 14105 7950 14185 7990
rect 14225 7950 14305 7990
rect 14105 7865 14305 7950
rect 14455 7990 14655 8065
rect 14455 7950 14535 7990
rect 14575 7950 14655 7990
rect 14455 7865 14655 7950
rect 9555 7640 9755 7715
rect 9555 7600 9635 7640
rect 9675 7600 9755 7640
rect 9555 7515 9755 7600
rect 9905 7640 10105 7715
rect 9905 7600 9985 7640
rect 10025 7600 10105 7640
rect 9905 7515 10105 7600
rect 10255 7640 10455 7715
rect 10255 7600 10335 7640
rect 10375 7600 10455 7640
rect 10255 7515 10455 7600
rect 10605 7640 10805 7715
rect 10605 7600 10685 7640
rect 10725 7600 10805 7640
rect 10605 7515 10805 7600
rect 10955 7640 11155 7715
rect 10955 7600 11035 7640
rect 11075 7600 11155 7640
rect 10955 7515 11155 7600
rect 11305 7640 11505 7715
rect 11305 7600 11385 7640
rect 11425 7600 11505 7640
rect 11305 7515 11505 7600
rect 11655 7640 11855 7715
rect 11655 7600 11735 7640
rect 11775 7600 11855 7640
rect 11655 7515 11855 7600
rect 12005 7640 12205 7715
rect 12005 7600 12085 7640
rect 12125 7600 12205 7640
rect 12005 7515 12205 7600
rect 12355 7640 12555 7715
rect 12355 7600 12435 7640
rect 12475 7600 12555 7640
rect 12355 7515 12555 7600
rect 12705 7640 12905 7715
rect 12705 7600 12785 7640
rect 12825 7600 12905 7640
rect 12705 7515 12905 7600
rect 13055 7640 13255 7715
rect 13055 7600 13135 7640
rect 13175 7600 13255 7640
rect 13055 7515 13255 7600
rect 13405 7640 13605 7715
rect 13405 7600 13485 7640
rect 13525 7600 13605 7640
rect 13405 7515 13605 7600
rect 13755 7640 13955 7715
rect 13755 7600 13835 7640
rect 13875 7600 13955 7640
rect 13755 7515 13955 7600
rect 14105 7640 14305 7715
rect 14105 7600 14185 7640
rect 14225 7600 14305 7640
rect 14105 7515 14305 7600
rect 14455 7640 14655 7715
rect 14455 7600 14535 7640
rect 14575 7600 14655 7640
rect 14455 7515 14655 7600
rect 9555 7290 9755 7365
rect 9555 7250 9635 7290
rect 9675 7250 9755 7290
rect 9555 7165 9755 7250
rect 9905 7290 10105 7365
rect 9905 7250 9985 7290
rect 10025 7250 10105 7290
rect 9905 7165 10105 7250
rect 10255 7290 10455 7365
rect 10255 7250 10335 7290
rect 10375 7250 10455 7290
rect 10255 7165 10455 7250
rect 10605 7290 10805 7365
rect 10605 7250 10685 7290
rect 10725 7250 10805 7290
rect 10605 7165 10805 7250
rect 10955 7290 11155 7365
rect 10955 7250 11035 7290
rect 11075 7250 11155 7290
rect 10955 7165 11155 7250
rect 11305 7290 11505 7365
rect 11305 7250 11385 7290
rect 11425 7250 11505 7290
rect 11305 7165 11505 7250
rect 11655 7290 11855 7365
rect 11655 7250 11735 7290
rect 11775 7250 11855 7290
rect 11655 7165 11855 7250
rect 12005 7290 12205 7365
rect 12005 7250 12085 7290
rect 12125 7250 12205 7290
rect 12005 7165 12205 7250
rect 12355 7290 12555 7365
rect 12355 7250 12435 7290
rect 12475 7250 12555 7290
rect 12355 7165 12555 7250
rect 12705 7290 12905 7365
rect 12705 7250 12785 7290
rect 12825 7250 12905 7290
rect 12705 7165 12905 7250
rect 13055 7290 13255 7365
rect 13055 7250 13135 7290
rect 13175 7250 13255 7290
rect 13055 7165 13255 7250
rect 13405 7290 13605 7365
rect 13405 7250 13485 7290
rect 13525 7250 13605 7290
rect 13405 7165 13605 7250
rect 13755 7290 13955 7365
rect 13755 7250 13835 7290
rect 13875 7250 13955 7290
rect 13755 7165 13955 7250
rect 14105 7290 14305 7365
rect 14105 7250 14185 7290
rect 14225 7250 14305 7290
rect 14105 7165 14305 7250
rect 14455 7290 14655 7365
rect 14455 7250 14535 7290
rect 14575 7250 14655 7290
rect 14455 7165 14655 7250
rect 9555 6940 9755 7015
rect 9555 6900 9635 6940
rect 9675 6900 9755 6940
rect 9555 6815 9755 6900
rect 9905 6940 10105 7015
rect 9905 6900 9985 6940
rect 10025 6900 10105 6940
rect 9905 6815 10105 6900
rect 10255 6940 10455 7015
rect 10255 6900 10335 6940
rect 10375 6900 10455 6940
rect 10255 6815 10455 6900
rect 10605 6940 10805 7015
rect 10605 6900 10685 6940
rect 10725 6900 10805 6940
rect 10605 6815 10805 6900
rect 10955 6940 11155 7015
rect 10955 6900 11035 6940
rect 11075 6900 11155 6940
rect 10955 6815 11155 6900
rect 11305 6940 11505 7015
rect 11305 6900 11385 6940
rect 11425 6900 11505 6940
rect 11305 6815 11505 6900
rect 11655 6940 11855 7015
rect 11655 6900 11735 6940
rect 11775 6900 11855 6940
rect 11655 6815 11855 6900
rect 12005 6940 12205 7015
rect 12005 6900 12085 6940
rect 12125 6900 12205 6940
rect 12005 6815 12205 6900
rect 12355 6940 12555 7015
rect 12355 6900 12435 6940
rect 12475 6900 12555 6940
rect 12355 6815 12555 6900
rect 12705 6940 12905 7015
rect 12705 6900 12785 6940
rect 12825 6900 12905 6940
rect 12705 6815 12905 6900
rect 13055 6940 13255 7015
rect 13055 6900 13135 6940
rect 13175 6900 13255 6940
rect 13055 6815 13255 6900
rect 13405 6940 13605 7015
rect 13405 6900 13485 6940
rect 13525 6900 13605 6940
rect 13405 6815 13605 6900
rect 13755 6940 13955 7015
rect 13755 6900 13835 6940
rect 13875 6900 13955 6940
rect 13755 6815 13955 6900
rect 14105 6940 14305 7015
rect 14105 6900 14185 6940
rect 14225 6900 14305 6940
rect 14105 6815 14305 6900
rect 14455 6940 14655 7015
rect 14455 6900 14535 6940
rect 14575 6900 14655 6940
rect 14455 6815 14655 6900
rect 9555 6590 9755 6665
rect 9555 6550 9635 6590
rect 9675 6550 9755 6590
rect 9555 6465 9755 6550
rect 9905 6590 10105 6665
rect 9905 6550 9985 6590
rect 10025 6550 10105 6590
rect 9905 6465 10105 6550
rect 10255 6590 10455 6665
rect 10255 6550 10335 6590
rect 10375 6550 10455 6590
rect 10255 6465 10455 6550
rect 10605 6590 10805 6665
rect 10605 6550 10685 6590
rect 10725 6550 10805 6590
rect 10605 6465 10805 6550
rect 10955 6590 11155 6665
rect 10955 6550 11035 6590
rect 11075 6550 11155 6590
rect 10955 6465 11155 6550
rect 11305 6590 11505 6665
rect 11305 6550 11385 6590
rect 11425 6550 11505 6590
rect 11305 6465 11505 6550
rect 11655 6590 11855 6665
rect 11655 6550 11735 6590
rect 11775 6550 11855 6590
rect 11655 6465 11855 6550
rect 12005 6590 12205 6665
rect 12005 6550 12085 6590
rect 12125 6550 12205 6590
rect 12005 6465 12205 6550
rect 12355 6590 12555 6665
rect 12355 6550 12435 6590
rect 12475 6550 12555 6590
rect 12355 6465 12555 6550
rect 12705 6590 12905 6665
rect 12705 6550 12785 6590
rect 12825 6550 12905 6590
rect 12705 6465 12905 6550
rect 13055 6590 13255 6665
rect 13055 6550 13135 6590
rect 13175 6550 13255 6590
rect 13055 6465 13255 6550
rect 13405 6590 13605 6665
rect 13405 6550 13485 6590
rect 13525 6550 13605 6590
rect 13405 6465 13605 6550
rect 13755 6590 13955 6665
rect 13755 6550 13835 6590
rect 13875 6550 13955 6590
rect 13755 6465 13955 6550
rect 14105 6590 14305 6665
rect 14105 6550 14185 6590
rect 14225 6550 14305 6590
rect 14105 6465 14305 6550
rect 14455 6590 14655 6665
rect 14455 6550 14535 6590
rect 14575 6550 14655 6590
rect 14455 6465 14655 6550
rect 1500 1370 1510 1380
<< mimcapcontact >>
rect -1165 18100 -1125 18140
rect -815 18100 -775 18140
rect -465 18100 -425 18140
rect -115 18100 -75 18140
rect 235 18100 275 18140
rect 585 18100 625 18140
rect 935 18100 975 18140
rect 1285 18100 1325 18140
rect 1635 18100 1675 18140
rect -1165 17750 -1125 17790
rect -815 17750 -775 17790
rect -465 17750 -425 17790
rect -115 17750 -75 17790
rect 235 17750 275 17790
rect 585 17750 625 17790
rect 935 17750 975 17790
rect 1285 17750 1325 17790
rect 1635 17750 1675 17790
rect -1165 17400 -1125 17440
rect -815 17400 -775 17440
rect -465 17400 -425 17440
rect -115 17400 -75 17440
rect 235 17400 275 17440
rect 585 17400 625 17440
rect 935 17400 975 17440
rect 1285 17400 1325 17440
rect 1635 17400 1675 17440
rect 9635 17400 9675 17440
rect 9985 17400 10025 17440
rect 10335 17400 10375 17440
rect 10685 17400 10725 17440
rect 11035 17400 11075 17440
rect 11385 17400 11425 17440
rect 11735 17400 11775 17440
rect 12085 17400 12125 17440
rect 12435 17400 12475 17440
rect 12785 17400 12825 17440
rect 13135 17400 13175 17440
rect 13485 17400 13525 17440
rect 13835 17400 13875 17440
rect 14185 17400 14225 17440
rect 14535 17400 14575 17440
rect -1165 17050 -1125 17090
rect -815 17050 -775 17090
rect -465 17050 -425 17090
rect -115 17050 -75 17090
rect 235 17050 275 17090
rect 585 17050 625 17090
rect 935 17050 975 17090
rect 1285 17050 1325 17090
rect 1635 17050 1675 17090
rect 9635 17050 9675 17090
rect 9985 17050 10025 17090
rect 10335 17050 10375 17090
rect 10685 17050 10725 17090
rect 11035 17050 11075 17090
rect 11385 17050 11425 17090
rect 11735 17050 11775 17090
rect 12085 17050 12125 17090
rect 12435 17050 12475 17090
rect 12785 17050 12825 17090
rect 13135 17050 13175 17090
rect 13485 17050 13525 17090
rect 13835 17050 13875 17090
rect 14185 17050 14225 17090
rect 14535 17050 14575 17090
rect -1165 16700 -1125 16740
rect -815 16700 -775 16740
rect -465 16700 -425 16740
rect -115 16700 -75 16740
rect 235 16700 275 16740
rect 585 16700 625 16740
rect 935 16700 975 16740
rect 1285 16700 1325 16740
rect 1635 16700 1675 16740
rect 9635 16700 9675 16740
rect 9985 16700 10025 16740
rect 10335 16700 10375 16740
rect 10685 16700 10725 16740
rect 11035 16700 11075 16740
rect 11385 16700 11425 16740
rect 11735 16700 11775 16740
rect 12085 16700 12125 16740
rect 12435 16700 12475 16740
rect 12785 16700 12825 16740
rect 13135 16700 13175 16740
rect 13485 16700 13525 16740
rect 13835 16700 13875 16740
rect 14185 16700 14225 16740
rect 14535 16700 14575 16740
rect -1165 16350 -1125 16390
rect -815 16350 -775 16390
rect -465 16350 -425 16390
rect -115 16350 -75 16390
rect 235 16350 275 16390
rect 585 16350 625 16390
rect 935 16350 975 16390
rect 1285 16350 1325 16390
rect 1635 16350 1675 16390
rect 9635 16350 9675 16390
rect 9985 16350 10025 16390
rect 10335 16350 10375 16390
rect 10685 16350 10725 16390
rect 11035 16350 11075 16390
rect 11385 16350 11425 16390
rect 11735 16350 11775 16390
rect 12085 16350 12125 16390
rect 12435 16350 12475 16390
rect 12785 16350 12825 16390
rect 13135 16350 13175 16390
rect 13485 16350 13525 16390
rect 13835 16350 13875 16390
rect 14185 16350 14225 16390
rect 14535 16350 14575 16390
rect -1165 16000 -1125 16040
rect -815 16000 -775 16040
rect -465 16000 -425 16040
rect -115 16000 -75 16040
rect 235 16000 275 16040
rect 585 16000 625 16040
rect 935 16000 975 16040
rect 1285 16000 1325 16040
rect 1635 16000 1675 16040
rect 9635 16000 9675 16040
rect 9985 16000 10025 16040
rect 10335 16000 10375 16040
rect 10685 16000 10725 16040
rect 11035 16000 11075 16040
rect 11385 16000 11425 16040
rect 11735 16000 11775 16040
rect 12085 16000 12125 16040
rect 12435 16000 12475 16040
rect 12785 16000 12825 16040
rect 13135 16000 13175 16040
rect 13485 16000 13525 16040
rect 13835 16000 13875 16040
rect 14185 16000 14225 16040
rect 14535 16000 14575 16040
rect -1165 15650 -1125 15690
rect -815 15650 -775 15690
rect -465 15650 -425 15690
rect -115 15650 -75 15690
rect 235 15650 275 15690
rect 585 15650 625 15690
rect 935 15650 975 15690
rect 1285 15650 1325 15690
rect 1635 15650 1675 15690
rect 9635 15650 9675 15690
rect 9985 15650 10025 15690
rect 10335 15650 10375 15690
rect 10685 15650 10725 15690
rect 11035 15650 11075 15690
rect 11385 15650 11425 15690
rect 11735 15650 11775 15690
rect 12085 15650 12125 15690
rect 12435 15650 12475 15690
rect 12785 15650 12825 15690
rect 13135 15650 13175 15690
rect 13485 15650 13525 15690
rect 13835 15650 13875 15690
rect 14185 15650 14225 15690
rect 14535 15650 14575 15690
rect -1165 15300 -1125 15340
rect -815 15300 -775 15340
rect -465 15300 -425 15340
rect -115 15300 -75 15340
rect 235 15300 275 15340
rect 585 15300 625 15340
rect 935 15300 975 15340
rect 1285 15300 1325 15340
rect 1635 15300 1675 15340
rect 9635 15300 9675 15340
rect 9985 15300 10025 15340
rect 10335 15300 10375 15340
rect 10685 15300 10725 15340
rect 11035 15300 11075 15340
rect 11385 15300 11425 15340
rect 11735 15300 11775 15340
rect 12085 15300 12125 15340
rect 12435 15300 12475 15340
rect 12785 15300 12825 15340
rect 13135 15300 13175 15340
rect 13485 15300 13525 15340
rect 13835 15300 13875 15340
rect 14185 15300 14225 15340
rect 14535 15300 14575 15340
rect -1165 14950 -1125 14990
rect -815 14950 -775 14990
rect -465 14950 -425 14990
rect -115 14950 -75 14990
rect 235 14950 275 14990
rect 585 14950 625 14990
rect 935 14950 975 14990
rect 1285 14950 1325 14990
rect 1635 14950 1675 14990
rect 9635 14950 9675 14990
rect 9985 14950 10025 14990
rect 10335 14950 10375 14990
rect 10685 14950 10725 14990
rect 11035 14950 11075 14990
rect 11385 14950 11425 14990
rect 11735 14950 11775 14990
rect 12085 14950 12125 14990
rect 12435 14950 12475 14990
rect 12785 14950 12825 14990
rect 13135 14950 13175 14990
rect 13485 14950 13525 14990
rect 13835 14950 13875 14990
rect 14185 14950 14225 14990
rect 14535 14950 14575 14990
rect -1165 14600 -1125 14640
rect -815 14600 -775 14640
rect -465 14600 -425 14640
rect -115 14600 -75 14640
rect 235 14600 275 14640
rect 585 14600 625 14640
rect 935 14600 975 14640
rect 1285 14600 1325 14640
rect 1635 14600 1675 14640
rect 9635 14600 9675 14640
rect 9985 14600 10025 14640
rect 10335 14600 10375 14640
rect 10685 14600 10725 14640
rect 11035 14600 11075 14640
rect 11385 14600 11425 14640
rect 11735 14600 11775 14640
rect 12085 14600 12125 14640
rect 12435 14600 12475 14640
rect 12785 14600 12825 14640
rect 13135 14600 13175 14640
rect 13485 14600 13525 14640
rect 13835 14600 13875 14640
rect 14185 14600 14225 14640
rect 14535 14600 14575 14640
rect -1165 14250 -1125 14290
rect -815 14250 -775 14290
rect -465 14250 -425 14290
rect -115 14250 -75 14290
rect 235 14250 275 14290
rect 585 14250 625 14290
rect 935 14250 975 14290
rect 1285 14250 1325 14290
rect 1635 14250 1675 14290
rect 9635 14250 9675 14290
rect 9985 14250 10025 14290
rect 10335 14250 10375 14290
rect 10685 14250 10725 14290
rect 11035 14250 11075 14290
rect 11385 14250 11425 14290
rect 11735 14250 11775 14290
rect 12085 14250 12125 14290
rect 12435 14250 12475 14290
rect 12785 14250 12825 14290
rect 13135 14250 13175 14290
rect 13485 14250 13525 14290
rect 13835 14250 13875 14290
rect 14185 14250 14225 14290
rect 14535 14250 14575 14290
rect -1165 13900 -1125 13940
rect -815 13900 -775 13940
rect -465 13900 -425 13940
rect -115 13900 -75 13940
rect 235 13900 275 13940
rect 585 13900 625 13940
rect 935 13900 975 13940
rect 1285 13900 1325 13940
rect 1635 13900 1675 13940
rect 9635 13900 9675 13940
rect 9985 13900 10025 13940
rect 10335 13900 10375 13940
rect 10685 13900 10725 13940
rect 11035 13900 11075 13940
rect 11385 13900 11425 13940
rect 11735 13900 11775 13940
rect 12085 13900 12125 13940
rect 12435 13900 12475 13940
rect 12785 13900 12825 13940
rect 13135 13900 13175 13940
rect 13485 13900 13525 13940
rect 13835 13900 13875 13940
rect 14185 13900 14225 13940
rect 14535 13900 14575 13940
rect -1165 13550 -1125 13590
rect -815 13550 -775 13590
rect -465 13550 -425 13590
rect -115 13550 -75 13590
rect 235 13550 275 13590
rect 585 13550 625 13590
rect 935 13550 975 13590
rect 1285 13550 1325 13590
rect 1635 13550 1675 13590
rect 9635 13550 9675 13590
rect 9985 13550 10025 13590
rect 10335 13550 10375 13590
rect 10685 13550 10725 13590
rect 11035 13550 11075 13590
rect 11385 13550 11425 13590
rect 11735 13550 11775 13590
rect 12085 13550 12125 13590
rect 12435 13550 12475 13590
rect 12785 13550 12825 13590
rect 13135 13550 13175 13590
rect 13485 13550 13525 13590
rect 13835 13550 13875 13590
rect 14185 13550 14225 13590
rect 14535 13550 14575 13590
rect -1165 13200 -1125 13240
rect -815 13200 -775 13240
rect -465 13200 -425 13240
rect -115 13200 -75 13240
rect 235 13200 275 13240
rect 585 13200 625 13240
rect 935 13200 975 13240
rect 1285 13200 1325 13240
rect 1635 13200 1675 13240
rect 9635 13200 9675 13240
rect 9985 13200 10025 13240
rect 10335 13200 10375 13240
rect 10685 13200 10725 13240
rect 11035 13200 11075 13240
rect 11385 13200 11425 13240
rect 11735 13200 11775 13240
rect 12085 13200 12125 13240
rect 12435 13200 12475 13240
rect 12785 13200 12825 13240
rect 13135 13200 13175 13240
rect 13485 13200 13525 13240
rect 13835 13200 13875 13240
rect 14185 13200 14225 13240
rect 14535 13200 14575 13240
rect -1165 12850 -1125 12890
rect -815 12850 -775 12890
rect -465 12850 -425 12890
rect -115 12850 -75 12890
rect 235 12850 275 12890
rect 585 12850 625 12890
rect 935 12850 975 12890
rect 1285 12850 1325 12890
rect 1635 12850 1675 12890
rect 9635 12850 9675 12890
rect 9985 12850 10025 12890
rect 10335 12850 10375 12890
rect 10685 12850 10725 12890
rect 11035 12850 11075 12890
rect 11385 12850 11425 12890
rect 11735 12850 11775 12890
rect 12085 12850 12125 12890
rect 12435 12850 12475 12890
rect 12785 12850 12825 12890
rect 13135 12850 13175 12890
rect 13485 12850 13525 12890
rect 13835 12850 13875 12890
rect 14185 12850 14225 12890
rect 14535 12850 14575 12890
rect -1165 12500 -1125 12540
rect -815 12500 -775 12540
rect -465 12500 -425 12540
rect -115 12500 -75 12540
rect 235 12500 275 12540
rect 585 12500 625 12540
rect 935 12500 975 12540
rect 1285 12500 1325 12540
rect 1635 12500 1675 12540
rect 9635 12500 9675 12540
rect 9985 12500 10025 12540
rect 10335 12500 10375 12540
rect 10685 12500 10725 12540
rect 11035 12500 11075 12540
rect 11385 12500 11425 12540
rect 11735 12500 11775 12540
rect 12085 12500 12125 12540
rect 12435 12500 12475 12540
rect 12785 12500 12825 12540
rect 13135 12500 13175 12540
rect 13485 12500 13525 12540
rect 13835 12500 13875 12540
rect 14185 12500 14225 12540
rect 14535 12500 14575 12540
rect -1165 12150 -1125 12190
rect -815 12150 -775 12190
rect -465 12150 -425 12190
rect -115 12150 -75 12190
rect 235 12150 275 12190
rect 585 12150 625 12190
rect 935 12150 975 12190
rect 1285 12150 1325 12190
rect 1635 12150 1675 12190
rect 9635 12150 9675 12190
rect 9985 12150 10025 12190
rect 10335 12150 10375 12190
rect 10685 12150 10725 12190
rect 11035 12150 11075 12190
rect 11385 12150 11425 12190
rect 11735 12150 11775 12190
rect 12085 12150 12125 12190
rect 12435 12150 12475 12190
rect 12785 12150 12825 12190
rect 13135 12150 13175 12190
rect 13485 12150 13525 12190
rect 13835 12150 13875 12190
rect 14185 12150 14225 12190
rect 14535 12150 14575 12190
rect -1165 11800 -1125 11840
rect -815 11800 -775 11840
rect -465 11800 -425 11840
rect -115 11800 -75 11840
rect 235 11800 275 11840
rect 585 11800 625 11840
rect 935 11800 975 11840
rect 1285 11800 1325 11840
rect 1635 11800 1675 11840
rect 9635 11800 9675 11840
rect 9985 11800 10025 11840
rect 10335 11800 10375 11840
rect 10685 11800 10725 11840
rect 11035 11800 11075 11840
rect 11385 11800 11425 11840
rect 11735 11800 11775 11840
rect 12085 11800 12125 11840
rect 12435 11800 12475 11840
rect 12785 11800 12825 11840
rect 13135 11800 13175 11840
rect 13485 11800 13525 11840
rect 13835 11800 13875 11840
rect 14185 11800 14225 11840
rect 14535 11800 14575 11840
rect -1165 11450 -1125 11490
rect -815 11450 -775 11490
rect -465 11450 -425 11490
rect -115 11450 -75 11490
rect 235 11450 275 11490
rect 585 11450 625 11490
rect 935 11450 975 11490
rect 1285 11450 1325 11490
rect 1635 11450 1675 11490
rect 9635 11450 9675 11490
rect 9985 11450 10025 11490
rect 10335 11450 10375 11490
rect 10685 11450 10725 11490
rect 11035 11450 11075 11490
rect 11385 11450 11425 11490
rect 11735 11450 11775 11490
rect 12085 11450 12125 11490
rect 12435 11450 12475 11490
rect 12785 11450 12825 11490
rect 13135 11450 13175 11490
rect 13485 11450 13525 11490
rect 13835 11450 13875 11490
rect 14185 11450 14225 11490
rect 14535 11450 14575 11490
rect -1165 11100 -1125 11140
rect -815 11100 -775 11140
rect -465 11100 -425 11140
rect -115 11100 -75 11140
rect 235 11100 275 11140
rect 585 11100 625 11140
rect 935 11100 975 11140
rect 1285 11100 1325 11140
rect 1635 11100 1675 11140
rect 9635 11100 9675 11140
rect 9985 11100 10025 11140
rect 10335 11100 10375 11140
rect 10685 11100 10725 11140
rect 11035 11100 11075 11140
rect 11385 11100 11425 11140
rect 11735 11100 11775 11140
rect 12085 11100 12125 11140
rect 12435 11100 12475 11140
rect 12785 11100 12825 11140
rect 13135 11100 13175 11140
rect 13485 11100 13525 11140
rect 13835 11100 13875 11140
rect 14185 11100 14225 11140
rect 14535 11100 14575 11140
rect -1165 10750 -1125 10790
rect -815 10750 -775 10790
rect -465 10750 -425 10790
rect -115 10750 -75 10790
rect 235 10750 275 10790
rect 585 10750 625 10790
rect 935 10750 975 10790
rect 1285 10750 1325 10790
rect 1635 10750 1675 10790
rect 9635 10750 9675 10790
rect 9985 10750 10025 10790
rect 10335 10750 10375 10790
rect 10685 10750 10725 10790
rect 11035 10750 11075 10790
rect 11385 10750 11425 10790
rect 11735 10750 11775 10790
rect 12085 10750 12125 10790
rect 12435 10750 12475 10790
rect 12785 10750 12825 10790
rect 13135 10750 13175 10790
rect 13485 10750 13525 10790
rect 13835 10750 13875 10790
rect 14185 10750 14225 10790
rect 14535 10750 14575 10790
rect -1165 10400 -1125 10440
rect -815 10400 -775 10440
rect -465 10400 -425 10440
rect -115 10400 -75 10440
rect 235 10400 275 10440
rect 585 10400 625 10440
rect 935 10400 975 10440
rect 1285 10400 1325 10440
rect 1635 10400 1675 10440
rect 9635 10400 9675 10440
rect 9985 10400 10025 10440
rect 10335 10400 10375 10440
rect 10685 10400 10725 10440
rect 11035 10400 11075 10440
rect 11385 10400 11425 10440
rect 11735 10400 11775 10440
rect 12085 10400 12125 10440
rect 12435 10400 12475 10440
rect 12785 10400 12825 10440
rect 13135 10400 13175 10440
rect 13485 10400 13525 10440
rect 13835 10400 13875 10440
rect 14185 10400 14225 10440
rect 14535 10400 14575 10440
rect -1165 10050 -1125 10090
rect -815 10050 -775 10090
rect -465 10050 -425 10090
rect -115 10050 -75 10090
rect 235 10050 275 10090
rect 585 10050 625 10090
rect 935 10050 975 10090
rect 1285 10050 1325 10090
rect 1635 10050 1675 10090
rect 9635 10050 9675 10090
rect 9985 10050 10025 10090
rect 10335 10050 10375 10090
rect 10685 10050 10725 10090
rect 11035 10050 11075 10090
rect 11385 10050 11425 10090
rect 11735 10050 11775 10090
rect 12085 10050 12125 10090
rect 12435 10050 12475 10090
rect 12785 10050 12825 10090
rect 13135 10050 13175 10090
rect 13485 10050 13525 10090
rect 13835 10050 13875 10090
rect 14185 10050 14225 10090
rect 14535 10050 14575 10090
rect 9635 9700 9675 9740
rect 9985 9700 10025 9740
rect 10335 9700 10375 9740
rect 10685 9700 10725 9740
rect 11035 9700 11075 9740
rect 11385 9700 11425 9740
rect 11735 9700 11775 9740
rect 12085 9700 12125 9740
rect 12435 9700 12475 9740
rect 12785 9700 12825 9740
rect 13135 9700 13175 9740
rect 13485 9700 13525 9740
rect 13835 9700 13875 9740
rect 14185 9700 14225 9740
rect 14535 9700 14575 9740
rect 9635 9350 9675 9390
rect 9985 9350 10025 9390
rect 10335 9350 10375 9390
rect 10685 9350 10725 9390
rect 11035 9350 11075 9390
rect 11385 9350 11425 9390
rect 11735 9350 11775 9390
rect 12085 9350 12125 9390
rect 12435 9350 12475 9390
rect 12785 9350 12825 9390
rect 13135 9350 13175 9390
rect 13485 9350 13525 9390
rect 13835 9350 13875 9390
rect 14185 9350 14225 9390
rect 14535 9350 14575 9390
rect 9635 9000 9675 9040
rect 9985 9000 10025 9040
rect 10335 9000 10375 9040
rect 10685 9000 10725 9040
rect 11035 9000 11075 9040
rect 11385 9000 11425 9040
rect 11735 9000 11775 9040
rect 12085 9000 12125 9040
rect 12435 9000 12475 9040
rect 12785 9000 12825 9040
rect 13135 9000 13175 9040
rect 13485 9000 13525 9040
rect 13835 9000 13875 9040
rect 14185 9000 14225 9040
rect 14535 9000 14575 9040
rect 9635 8650 9675 8690
rect 9985 8650 10025 8690
rect 10335 8650 10375 8690
rect 10685 8650 10725 8690
rect 11035 8650 11075 8690
rect 11385 8650 11425 8690
rect 11735 8650 11775 8690
rect 12085 8650 12125 8690
rect 12435 8650 12475 8690
rect 12785 8650 12825 8690
rect 13135 8650 13175 8690
rect 13485 8650 13525 8690
rect 13835 8650 13875 8690
rect 14185 8650 14225 8690
rect 14535 8650 14575 8690
rect 9635 8300 9675 8340
rect 9985 8300 10025 8340
rect 10335 8300 10375 8340
rect 10685 8300 10725 8340
rect 11035 8300 11075 8340
rect 11385 8300 11425 8340
rect 11735 8300 11775 8340
rect 12085 8300 12125 8340
rect 12435 8300 12475 8340
rect 12785 8300 12825 8340
rect 13135 8300 13175 8340
rect 13485 8300 13525 8340
rect 13835 8300 13875 8340
rect 14185 8300 14225 8340
rect 14535 8300 14575 8340
rect 9635 7950 9675 7990
rect 9985 7950 10025 7990
rect 10335 7950 10375 7990
rect 10685 7950 10725 7990
rect 11035 7950 11075 7990
rect 11385 7950 11425 7990
rect 11735 7950 11775 7990
rect 12085 7950 12125 7990
rect 12435 7950 12475 7990
rect 12785 7950 12825 7990
rect 13135 7950 13175 7990
rect 13485 7950 13525 7990
rect 13835 7950 13875 7990
rect 14185 7950 14225 7990
rect 14535 7950 14575 7990
rect 9635 7600 9675 7640
rect 9985 7600 10025 7640
rect 10335 7600 10375 7640
rect 10685 7600 10725 7640
rect 11035 7600 11075 7640
rect 11385 7600 11425 7640
rect 11735 7600 11775 7640
rect 12085 7600 12125 7640
rect 12435 7600 12475 7640
rect 12785 7600 12825 7640
rect 13135 7600 13175 7640
rect 13485 7600 13525 7640
rect 13835 7600 13875 7640
rect 14185 7600 14225 7640
rect 14535 7600 14575 7640
rect 9635 7250 9675 7290
rect 9985 7250 10025 7290
rect 10335 7250 10375 7290
rect 10685 7250 10725 7290
rect 11035 7250 11075 7290
rect 11385 7250 11425 7290
rect 11735 7250 11775 7290
rect 12085 7250 12125 7290
rect 12435 7250 12475 7290
rect 12785 7250 12825 7290
rect 13135 7250 13175 7290
rect 13485 7250 13525 7290
rect 13835 7250 13875 7290
rect 14185 7250 14225 7290
rect 14535 7250 14575 7290
rect 9635 6900 9675 6940
rect 9985 6900 10025 6940
rect 10335 6900 10375 6940
rect 10685 6900 10725 6940
rect 11035 6900 11075 6940
rect 11385 6900 11425 6940
rect 11735 6900 11775 6940
rect 12085 6900 12125 6940
rect 12435 6900 12475 6940
rect 12785 6900 12825 6940
rect 13135 6900 13175 6940
rect 13485 6900 13525 6940
rect 13835 6900 13875 6940
rect 14185 6900 14225 6940
rect 14535 6900 14575 6940
rect 9635 6550 9675 6590
rect 9985 6550 10025 6590
rect 10335 6550 10375 6590
rect 10685 6550 10725 6590
rect 11035 6550 11075 6590
rect 11385 6550 11425 6590
rect 11735 6550 11775 6590
rect 12085 6550 12125 6590
rect 12435 6550 12475 6590
rect 12785 6550 12825 6590
rect 13135 6550 13175 6590
rect 13485 6550 13525 6590
rect 13835 6550 13875 6590
rect 14185 6550 14225 6590
rect 14535 6550 14575 6590
<< metal4 >>
rect 2320 20915 17990 20925
rect 2320 20875 2330 20915
rect 2370 20875 6700 20915
rect 6740 20890 17990 20915
rect 6740 20875 14825 20890
rect 2320 20850 14825 20875
rect 2320 20810 2330 20850
rect 2370 20810 6700 20850
rect 6740 20840 14825 20850
rect 14875 20840 14920 20890
rect 14970 20840 15015 20890
rect 15065 20840 15115 20890
rect 15165 20840 15215 20890
rect 15265 20840 15315 20890
rect 15365 20840 15410 20890
rect 15460 20840 15505 20890
rect 15555 20840 15625 20890
rect 15675 20840 15720 20890
rect 15770 20840 15815 20890
rect 15865 20840 15915 20890
rect 15965 20840 16015 20890
rect 16065 20840 16115 20890
rect 16165 20840 16210 20890
rect 16260 20840 16305 20890
rect 16355 20840 16425 20890
rect 16475 20840 16520 20890
rect 16570 20840 16615 20890
rect 16665 20840 16715 20890
rect 16765 20840 16815 20890
rect 16865 20840 16915 20890
rect 16965 20840 17010 20890
rect 17060 20840 17105 20890
rect 17155 20840 17225 20890
rect 17275 20840 17320 20890
rect 17370 20840 17415 20890
rect 17465 20840 17515 20890
rect 17565 20840 17615 20890
rect 17665 20840 17715 20890
rect 17765 20840 17810 20890
rect 17860 20840 17905 20890
rect 17955 20840 17990 20890
rect 6740 20810 17990 20840
rect 2320 20800 17990 20810
rect 2320 20780 14825 20800
rect 2320 20740 2330 20780
rect 2370 20740 6700 20780
rect 6740 20750 14825 20780
rect 14875 20750 14920 20800
rect 14970 20750 15015 20800
rect 15065 20750 15115 20800
rect 15165 20750 15215 20800
rect 15265 20750 15315 20800
rect 15365 20750 15410 20800
rect 15460 20750 15505 20800
rect 15555 20750 15625 20800
rect 15675 20750 15720 20800
rect 15770 20750 15815 20800
rect 15865 20750 15915 20800
rect 15965 20750 16015 20800
rect 16065 20750 16115 20800
rect 16165 20750 16210 20800
rect 16260 20750 16305 20800
rect 16355 20750 16425 20800
rect 16475 20750 16520 20800
rect 16570 20750 16615 20800
rect 16665 20750 16715 20800
rect 16765 20750 16815 20800
rect 16865 20750 16915 20800
rect 16965 20750 17010 20800
rect 17060 20750 17105 20800
rect 17155 20750 17225 20800
rect 17275 20750 17320 20800
rect 17370 20750 17415 20800
rect 17465 20750 17515 20800
rect 17565 20750 17615 20800
rect 17665 20750 17715 20800
rect 17765 20750 17810 20800
rect 17860 20750 17905 20800
rect 17955 20750 17990 20800
rect 6740 20740 17990 20750
rect 2320 20710 17990 20740
rect 2320 20670 2330 20710
rect 2370 20670 6700 20710
rect 6740 20700 17990 20710
rect 6740 20670 14825 20700
rect 2320 20650 14825 20670
rect 14875 20650 14920 20700
rect 14970 20650 15015 20700
rect 15065 20650 15115 20700
rect 15165 20650 15215 20700
rect 15265 20650 15315 20700
rect 15365 20650 15410 20700
rect 15460 20650 15505 20700
rect 15555 20650 15625 20700
rect 15675 20650 15720 20700
rect 15770 20650 15815 20700
rect 15865 20650 15915 20700
rect 15965 20650 16015 20700
rect 16065 20650 16115 20700
rect 16165 20650 16210 20700
rect 16260 20650 16305 20700
rect 16355 20650 16425 20700
rect 16475 20650 16520 20700
rect 16570 20650 16615 20700
rect 16665 20650 16715 20700
rect 16765 20650 16815 20700
rect 16865 20650 16915 20700
rect 16965 20650 17010 20700
rect 17060 20650 17105 20700
rect 17155 20650 17225 20700
rect 17275 20650 17320 20700
rect 17370 20650 17415 20700
rect 17465 20650 17515 20700
rect 17565 20650 17615 20700
rect 17665 20650 17715 20700
rect 17765 20650 17810 20700
rect 17860 20650 17905 20700
rect 17955 20650 17990 20700
rect 2320 20640 17990 20650
rect 2320 20600 2330 20640
rect 2370 20600 6700 20640
rect 6740 20610 17990 20640
rect 6740 20600 14825 20610
rect 2320 20575 14825 20600
rect 2320 20535 2330 20575
rect 2370 20535 6700 20575
rect 6740 20560 14825 20575
rect 14875 20560 14920 20610
rect 14970 20560 15015 20610
rect 15065 20560 15115 20610
rect 15165 20560 15215 20610
rect 15265 20560 15315 20610
rect 15365 20560 15410 20610
rect 15460 20560 15505 20610
rect 15555 20560 15625 20610
rect 15675 20560 15720 20610
rect 15770 20560 15815 20610
rect 15865 20560 15915 20610
rect 15965 20560 16015 20610
rect 16065 20560 16115 20610
rect 16165 20560 16210 20610
rect 16260 20560 16305 20610
rect 16355 20560 16425 20610
rect 16475 20560 16520 20610
rect 16570 20560 16615 20610
rect 16665 20560 16715 20610
rect 16765 20560 16815 20610
rect 16865 20560 16915 20610
rect 16965 20560 17010 20610
rect 17060 20560 17105 20610
rect 17155 20560 17225 20610
rect 17275 20560 17320 20610
rect 17370 20560 17415 20610
rect 17465 20560 17515 20610
rect 17565 20560 17615 20610
rect 17665 20560 17715 20610
rect 17765 20560 17810 20610
rect 17860 20560 17905 20610
rect 17955 20560 17990 20610
rect 6740 20535 17990 20560
rect 2320 20515 17990 20535
rect 2320 20475 2330 20515
rect 2370 20475 6700 20515
rect 6740 20490 17990 20515
rect 6740 20475 14825 20490
rect 2320 20450 14825 20475
rect 2320 20410 2330 20450
rect 2370 20410 6700 20450
rect 6740 20440 14825 20450
rect 14875 20440 14920 20490
rect 14970 20440 15015 20490
rect 15065 20440 15115 20490
rect 15165 20440 15215 20490
rect 15265 20440 15315 20490
rect 15365 20440 15410 20490
rect 15460 20440 15505 20490
rect 15555 20440 15625 20490
rect 15675 20440 15720 20490
rect 15770 20440 15815 20490
rect 15865 20440 15915 20490
rect 15965 20440 16015 20490
rect 16065 20440 16115 20490
rect 16165 20440 16210 20490
rect 16260 20440 16305 20490
rect 16355 20440 16425 20490
rect 16475 20440 16520 20490
rect 16570 20440 16615 20490
rect 16665 20440 16715 20490
rect 16765 20440 16815 20490
rect 16865 20440 16915 20490
rect 16965 20440 17010 20490
rect 17060 20440 17105 20490
rect 17155 20440 17225 20490
rect 17275 20440 17320 20490
rect 17370 20440 17415 20490
rect 17465 20440 17515 20490
rect 17565 20440 17615 20490
rect 17665 20440 17715 20490
rect 17765 20440 17810 20490
rect 17860 20440 17905 20490
rect 17955 20440 17990 20490
rect 6740 20410 17990 20440
rect 2320 20400 17990 20410
rect 2320 20380 14825 20400
rect 2320 20340 2330 20380
rect 2370 20340 6700 20380
rect 6740 20350 14825 20380
rect 14875 20350 14920 20400
rect 14970 20350 15015 20400
rect 15065 20350 15115 20400
rect 15165 20350 15215 20400
rect 15265 20350 15315 20400
rect 15365 20350 15410 20400
rect 15460 20350 15505 20400
rect 15555 20350 15625 20400
rect 15675 20350 15720 20400
rect 15770 20350 15815 20400
rect 15865 20350 15915 20400
rect 15965 20350 16015 20400
rect 16065 20350 16115 20400
rect 16165 20350 16210 20400
rect 16260 20350 16305 20400
rect 16355 20350 16425 20400
rect 16475 20350 16520 20400
rect 16570 20350 16615 20400
rect 16665 20350 16715 20400
rect 16765 20350 16815 20400
rect 16865 20350 16915 20400
rect 16965 20350 17010 20400
rect 17060 20350 17105 20400
rect 17155 20350 17225 20400
rect 17275 20350 17320 20400
rect 17370 20350 17415 20400
rect 17465 20350 17515 20400
rect 17565 20350 17615 20400
rect 17665 20350 17715 20400
rect 17765 20350 17810 20400
rect 17860 20350 17905 20400
rect 17955 20350 17990 20400
rect 6740 20340 17990 20350
rect 2320 20310 17990 20340
rect 2320 20270 2330 20310
rect 2370 20270 6700 20310
rect 6740 20300 17990 20310
rect 6740 20270 14825 20300
rect 2320 20250 14825 20270
rect 14875 20250 14920 20300
rect 14970 20250 15015 20300
rect 15065 20250 15115 20300
rect 15165 20250 15215 20300
rect 15265 20250 15315 20300
rect 15365 20250 15410 20300
rect 15460 20250 15505 20300
rect 15555 20250 15625 20300
rect 15675 20250 15720 20300
rect 15770 20250 15815 20300
rect 15865 20250 15915 20300
rect 15965 20250 16015 20300
rect 16065 20250 16115 20300
rect 16165 20250 16210 20300
rect 16260 20250 16305 20300
rect 16355 20250 16425 20300
rect 16475 20250 16520 20300
rect 16570 20250 16615 20300
rect 16665 20250 16715 20300
rect 16765 20250 16815 20300
rect 16865 20250 16915 20300
rect 16965 20250 17010 20300
rect 17060 20250 17105 20300
rect 17155 20250 17225 20300
rect 17275 20250 17320 20300
rect 17370 20250 17415 20300
rect 17465 20250 17515 20300
rect 17565 20250 17615 20300
rect 17665 20250 17715 20300
rect 17765 20250 17810 20300
rect 17860 20250 17905 20300
rect 17955 20250 17990 20300
rect 2320 20240 17990 20250
rect 2320 20200 2330 20240
rect 2370 20200 6700 20240
rect 6740 20210 17990 20240
rect 6740 20200 14825 20210
rect 2320 20175 14825 20200
rect 2320 20135 2330 20175
rect 2370 20135 6700 20175
rect 6740 20160 14825 20175
rect 14875 20160 14920 20210
rect 14970 20160 15015 20210
rect 15065 20160 15115 20210
rect 15165 20160 15215 20210
rect 15265 20160 15315 20210
rect 15365 20160 15410 20210
rect 15460 20160 15505 20210
rect 15555 20160 15625 20210
rect 15675 20160 15720 20210
rect 15770 20160 15815 20210
rect 15865 20160 15915 20210
rect 15965 20160 16015 20210
rect 16065 20160 16115 20210
rect 16165 20160 16210 20210
rect 16260 20160 16305 20210
rect 16355 20160 16425 20210
rect 16475 20160 16520 20210
rect 16570 20160 16615 20210
rect 16665 20160 16715 20210
rect 16765 20160 16815 20210
rect 16865 20160 16915 20210
rect 16965 20160 17010 20210
rect 17060 20160 17105 20210
rect 17155 20160 17225 20210
rect 17275 20160 17320 20210
rect 17370 20160 17415 20210
rect 17465 20160 17515 20210
rect 17565 20160 17615 20210
rect 17665 20160 17715 20210
rect 17765 20160 17810 20210
rect 17860 20160 17905 20210
rect 17955 20160 17990 20210
rect 6740 20135 17990 20160
rect 2320 20115 17990 20135
rect 2320 20075 2330 20115
rect 2370 20075 6700 20115
rect 6740 20090 17990 20115
rect 6740 20075 14825 20090
rect 2320 20050 14825 20075
rect 2320 20010 2330 20050
rect 2370 20010 6700 20050
rect 6740 20040 14825 20050
rect 14875 20040 14920 20090
rect 14970 20040 15015 20090
rect 15065 20040 15115 20090
rect 15165 20040 15215 20090
rect 15265 20040 15315 20090
rect 15365 20040 15410 20090
rect 15460 20040 15505 20090
rect 15555 20040 15625 20090
rect 15675 20040 15720 20090
rect 15770 20040 15815 20090
rect 15865 20040 15915 20090
rect 15965 20040 16015 20090
rect 16065 20040 16115 20090
rect 16165 20040 16210 20090
rect 16260 20040 16305 20090
rect 16355 20040 16425 20090
rect 16475 20040 16520 20090
rect 16570 20040 16615 20090
rect 16665 20040 16715 20090
rect 16765 20040 16815 20090
rect 16865 20040 16915 20090
rect 16965 20040 17010 20090
rect 17060 20040 17105 20090
rect 17155 20040 17225 20090
rect 17275 20040 17320 20090
rect 17370 20040 17415 20090
rect 17465 20040 17515 20090
rect 17565 20040 17615 20090
rect 17665 20040 17715 20090
rect 17765 20040 17810 20090
rect 17860 20040 17905 20090
rect 17955 20040 17990 20090
rect 6740 20010 17990 20040
rect 2320 20000 17990 20010
rect 2320 19980 14825 20000
rect 2320 19940 2330 19980
rect 2370 19940 6700 19980
rect 6740 19950 14825 19980
rect 14875 19950 14920 20000
rect 14970 19950 15015 20000
rect 15065 19950 15115 20000
rect 15165 19950 15215 20000
rect 15265 19950 15315 20000
rect 15365 19950 15410 20000
rect 15460 19950 15505 20000
rect 15555 19950 15625 20000
rect 15675 19950 15720 20000
rect 15770 19950 15815 20000
rect 15865 19950 15915 20000
rect 15965 19950 16015 20000
rect 16065 19950 16115 20000
rect 16165 19950 16210 20000
rect 16260 19950 16305 20000
rect 16355 19950 16425 20000
rect 16475 19950 16520 20000
rect 16570 19950 16615 20000
rect 16665 19950 16715 20000
rect 16765 19950 16815 20000
rect 16865 19950 16915 20000
rect 16965 19950 17010 20000
rect 17060 19950 17105 20000
rect 17155 19950 17225 20000
rect 17275 19950 17320 20000
rect 17370 19950 17415 20000
rect 17465 19950 17515 20000
rect 17565 19950 17615 20000
rect 17665 19950 17715 20000
rect 17765 19950 17810 20000
rect 17860 19950 17905 20000
rect 17955 19950 17990 20000
rect 6740 19940 17990 19950
rect 2320 19910 17990 19940
rect 2320 19870 2330 19910
rect 2370 19870 6700 19910
rect 6740 19900 17990 19910
rect 6740 19870 14825 19900
rect 2320 19850 14825 19870
rect 14875 19850 14920 19900
rect 14970 19850 15015 19900
rect 15065 19850 15115 19900
rect 15165 19850 15215 19900
rect 15265 19850 15315 19900
rect 15365 19850 15410 19900
rect 15460 19850 15505 19900
rect 15555 19850 15625 19900
rect 15675 19850 15720 19900
rect 15770 19850 15815 19900
rect 15865 19850 15915 19900
rect 15965 19850 16015 19900
rect 16065 19850 16115 19900
rect 16165 19850 16210 19900
rect 16260 19850 16305 19900
rect 16355 19850 16425 19900
rect 16475 19850 16520 19900
rect 16570 19850 16615 19900
rect 16665 19850 16715 19900
rect 16765 19850 16815 19900
rect 16865 19850 16915 19900
rect 16965 19850 17010 19900
rect 17060 19850 17105 19900
rect 17155 19850 17225 19900
rect 17275 19850 17320 19900
rect 17370 19850 17415 19900
rect 17465 19850 17515 19900
rect 17565 19850 17615 19900
rect 17665 19850 17715 19900
rect 17765 19850 17810 19900
rect 17860 19850 17905 19900
rect 17955 19850 17990 19900
rect 2320 19840 17990 19850
rect 2320 19800 2330 19840
rect 2370 19800 6700 19840
rect 6740 19810 17990 19840
rect 6740 19800 14825 19810
rect 2320 19775 14825 19800
rect 2320 19735 2330 19775
rect 2370 19735 6700 19775
rect 6740 19760 14825 19775
rect 14875 19760 14920 19810
rect 14970 19760 15015 19810
rect 15065 19760 15115 19810
rect 15165 19760 15215 19810
rect 15265 19760 15315 19810
rect 15365 19760 15410 19810
rect 15460 19760 15505 19810
rect 15555 19760 15625 19810
rect 15675 19760 15720 19810
rect 15770 19760 15815 19810
rect 15865 19760 15915 19810
rect 15965 19760 16015 19810
rect 16065 19760 16115 19810
rect 16165 19760 16210 19810
rect 16260 19760 16305 19810
rect 16355 19760 16425 19810
rect 16475 19760 16520 19810
rect 16570 19760 16615 19810
rect 16665 19760 16715 19810
rect 16765 19760 16815 19810
rect 16865 19760 16915 19810
rect 16965 19760 17010 19810
rect 17060 19760 17105 19810
rect 17155 19760 17225 19810
rect 17275 19760 17320 19810
rect 17370 19760 17415 19810
rect 17465 19760 17515 19810
rect 17565 19760 17615 19810
rect 17665 19760 17715 19810
rect 17765 19760 17810 19810
rect 17860 19760 17905 19810
rect 17955 19760 17990 19810
rect 6740 19735 17990 19760
rect 2320 19715 17990 19735
rect 2320 19675 2330 19715
rect 2370 19675 6700 19715
rect 6740 19690 17990 19715
rect 6740 19675 14825 19690
rect 2320 19650 14825 19675
rect 2320 19610 2330 19650
rect 2370 19610 6700 19650
rect 6740 19640 14825 19650
rect 14875 19640 14920 19690
rect 14970 19640 15015 19690
rect 15065 19640 15115 19690
rect 15165 19640 15215 19690
rect 15265 19640 15315 19690
rect 15365 19640 15410 19690
rect 15460 19640 15505 19690
rect 15555 19640 15625 19690
rect 15675 19640 15720 19690
rect 15770 19640 15815 19690
rect 15865 19640 15915 19690
rect 15965 19640 16015 19690
rect 16065 19640 16115 19690
rect 16165 19640 16210 19690
rect 16260 19640 16305 19690
rect 16355 19640 16425 19690
rect 16475 19640 16520 19690
rect 16570 19640 16615 19690
rect 16665 19640 16715 19690
rect 16765 19640 16815 19690
rect 16865 19640 16915 19690
rect 16965 19640 17010 19690
rect 17060 19640 17105 19690
rect 17155 19640 17225 19690
rect 17275 19640 17320 19690
rect 17370 19640 17415 19690
rect 17465 19640 17515 19690
rect 17565 19640 17615 19690
rect 17665 19640 17715 19690
rect 17765 19640 17810 19690
rect 17860 19640 17905 19690
rect 17955 19640 17990 19690
rect 6740 19610 17990 19640
rect 2320 19600 17990 19610
rect 2320 19580 14825 19600
rect 2320 19540 2330 19580
rect 2370 19540 6700 19580
rect 6740 19550 14825 19580
rect 14875 19550 14920 19600
rect 14970 19550 15015 19600
rect 15065 19550 15115 19600
rect 15165 19550 15215 19600
rect 15265 19550 15315 19600
rect 15365 19550 15410 19600
rect 15460 19550 15505 19600
rect 15555 19550 15625 19600
rect 15675 19550 15720 19600
rect 15770 19550 15815 19600
rect 15865 19550 15915 19600
rect 15965 19550 16015 19600
rect 16065 19550 16115 19600
rect 16165 19550 16210 19600
rect 16260 19550 16305 19600
rect 16355 19550 16425 19600
rect 16475 19550 16520 19600
rect 16570 19550 16615 19600
rect 16665 19550 16715 19600
rect 16765 19550 16815 19600
rect 16865 19550 16915 19600
rect 16965 19550 17010 19600
rect 17060 19550 17105 19600
rect 17155 19550 17225 19600
rect 17275 19550 17320 19600
rect 17370 19550 17415 19600
rect 17465 19550 17515 19600
rect 17565 19550 17615 19600
rect 17665 19550 17715 19600
rect 17765 19550 17810 19600
rect 17860 19550 17905 19600
rect 17955 19550 17990 19600
rect 6740 19540 17990 19550
rect 2320 19510 17990 19540
rect 2320 19470 2330 19510
rect 2370 19470 6700 19510
rect 6740 19500 17990 19510
rect 6740 19470 14825 19500
rect 2320 19450 14825 19470
rect 14875 19450 14920 19500
rect 14970 19450 15015 19500
rect 15065 19450 15115 19500
rect 15165 19450 15215 19500
rect 15265 19450 15315 19500
rect 15365 19450 15410 19500
rect 15460 19450 15505 19500
rect 15555 19450 15625 19500
rect 15675 19450 15720 19500
rect 15770 19450 15815 19500
rect 15865 19450 15915 19500
rect 15965 19450 16015 19500
rect 16065 19450 16115 19500
rect 16165 19450 16210 19500
rect 16260 19450 16305 19500
rect 16355 19450 16425 19500
rect 16475 19450 16520 19500
rect 16570 19450 16615 19500
rect 16665 19450 16715 19500
rect 16765 19450 16815 19500
rect 16865 19450 16915 19500
rect 16965 19450 17010 19500
rect 17060 19450 17105 19500
rect 17155 19450 17225 19500
rect 17275 19450 17320 19500
rect 17370 19450 17415 19500
rect 17465 19450 17515 19500
rect 17565 19450 17615 19500
rect 17665 19450 17715 19500
rect 17765 19450 17810 19500
rect 17860 19450 17905 19500
rect 17955 19450 17990 19500
rect 2320 19440 17990 19450
rect 2320 19400 2330 19440
rect 2370 19400 6700 19440
rect 6740 19410 17990 19440
rect 6740 19400 14825 19410
rect 2320 19375 14825 19400
rect 2320 19335 2330 19375
rect 2370 19335 6700 19375
rect 6740 19360 14825 19375
rect 14875 19360 14920 19410
rect 14970 19360 15015 19410
rect 15065 19360 15115 19410
rect 15165 19360 15215 19410
rect 15265 19360 15315 19410
rect 15365 19360 15410 19410
rect 15460 19360 15505 19410
rect 15555 19360 15625 19410
rect 15675 19360 15720 19410
rect 15770 19360 15815 19410
rect 15865 19360 15915 19410
rect 15965 19360 16015 19410
rect 16065 19360 16115 19410
rect 16165 19360 16210 19410
rect 16260 19360 16305 19410
rect 16355 19360 16425 19410
rect 16475 19360 16520 19410
rect 16570 19360 16615 19410
rect 16665 19360 16715 19410
rect 16765 19360 16815 19410
rect 16865 19360 16915 19410
rect 16965 19360 17010 19410
rect 17060 19360 17105 19410
rect 17155 19360 17225 19410
rect 17275 19360 17320 19410
rect 17370 19360 17415 19410
rect 17465 19360 17515 19410
rect 17565 19360 17615 19410
rect 17665 19360 17715 19410
rect 17765 19360 17810 19410
rect 17860 19360 17905 19410
rect 17955 19360 17990 19410
rect 6740 19335 17990 19360
rect 2320 19315 17990 19335
rect 2320 19275 2330 19315
rect 2370 19275 6700 19315
rect 6740 19290 17990 19315
rect 6740 19275 14825 19290
rect 2320 19250 14825 19275
rect 2320 19210 2330 19250
rect 2370 19210 6700 19250
rect 6740 19240 14825 19250
rect 14875 19240 14920 19290
rect 14970 19240 15015 19290
rect 15065 19240 15115 19290
rect 15165 19240 15215 19290
rect 15265 19240 15315 19290
rect 15365 19240 15410 19290
rect 15460 19240 15505 19290
rect 15555 19240 15625 19290
rect 15675 19240 15720 19290
rect 15770 19240 15815 19290
rect 15865 19240 15915 19290
rect 15965 19240 16015 19290
rect 16065 19240 16115 19290
rect 16165 19240 16210 19290
rect 16260 19240 16305 19290
rect 16355 19240 16425 19290
rect 16475 19240 16520 19290
rect 16570 19240 16615 19290
rect 16665 19240 16715 19290
rect 16765 19240 16815 19290
rect 16865 19240 16915 19290
rect 16965 19240 17010 19290
rect 17060 19240 17105 19290
rect 17155 19240 17225 19290
rect 17275 19240 17320 19290
rect 17370 19240 17415 19290
rect 17465 19240 17515 19290
rect 17565 19240 17615 19290
rect 17665 19240 17715 19290
rect 17765 19240 17810 19290
rect 17860 19240 17905 19290
rect 17955 19240 17990 19290
rect 6740 19210 17990 19240
rect 2320 19200 17990 19210
rect 2320 19180 14825 19200
rect 2320 19140 2330 19180
rect 2370 19140 6700 19180
rect 6740 19150 14825 19180
rect 14875 19150 14920 19200
rect 14970 19150 15015 19200
rect 15065 19150 15115 19200
rect 15165 19150 15215 19200
rect 15265 19150 15315 19200
rect 15365 19150 15410 19200
rect 15460 19150 15505 19200
rect 15555 19150 15625 19200
rect 15675 19150 15720 19200
rect 15770 19150 15815 19200
rect 15865 19150 15915 19200
rect 15965 19150 16015 19200
rect 16065 19150 16115 19200
rect 16165 19150 16210 19200
rect 16260 19150 16305 19200
rect 16355 19150 16425 19200
rect 16475 19150 16520 19200
rect 16570 19150 16615 19200
rect 16665 19150 16715 19200
rect 16765 19150 16815 19200
rect 16865 19150 16915 19200
rect 16965 19150 17010 19200
rect 17060 19150 17105 19200
rect 17155 19150 17225 19200
rect 17275 19150 17320 19200
rect 17370 19150 17415 19200
rect 17465 19150 17515 19200
rect 17565 19150 17615 19200
rect 17665 19150 17715 19200
rect 17765 19150 17810 19200
rect 17860 19150 17905 19200
rect 17955 19150 17990 19200
rect 6740 19140 17990 19150
rect 2320 19110 17990 19140
rect 2320 19070 2330 19110
rect 2370 19070 6700 19110
rect 6740 19100 17990 19110
rect 6740 19070 14825 19100
rect 2320 19050 14825 19070
rect 14875 19050 14920 19100
rect 14970 19050 15015 19100
rect 15065 19050 15115 19100
rect 15165 19050 15215 19100
rect 15265 19050 15315 19100
rect 15365 19050 15410 19100
rect 15460 19050 15505 19100
rect 15555 19050 15625 19100
rect 15675 19050 15720 19100
rect 15770 19050 15815 19100
rect 15865 19050 15915 19100
rect 15965 19050 16015 19100
rect 16065 19050 16115 19100
rect 16165 19050 16210 19100
rect 16260 19050 16305 19100
rect 16355 19050 16425 19100
rect 16475 19050 16520 19100
rect 16570 19050 16615 19100
rect 16665 19050 16715 19100
rect 16765 19050 16815 19100
rect 16865 19050 16915 19100
rect 16965 19050 17010 19100
rect 17060 19050 17105 19100
rect 17155 19050 17225 19100
rect 17275 19050 17320 19100
rect 17370 19050 17415 19100
rect 17465 19050 17515 19100
rect 17565 19050 17615 19100
rect 17665 19050 17715 19100
rect 17765 19050 17810 19100
rect 17860 19050 17905 19100
rect 17955 19050 17990 19100
rect 2320 19040 17990 19050
rect 2320 19000 2330 19040
rect 2370 19000 6700 19040
rect 6740 19010 17990 19040
rect 6740 19000 14825 19010
rect 2320 18975 14825 19000
rect 2320 18935 2330 18975
rect 2370 18935 6700 18975
rect 6740 18960 14825 18975
rect 14875 18960 14920 19010
rect 14970 18960 15015 19010
rect 15065 18960 15115 19010
rect 15165 18960 15215 19010
rect 15265 18960 15315 19010
rect 15365 18960 15410 19010
rect 15460 18960 15505 19010
rect 15555 18960 15625 19010
rect 15675 18960 15720 19010
rect 15770 18960 15815 19010
rect 15865 18960 15915 19010
rect 15965 18960 16015 19010
rect 16065 18960 16115 19010
rect 16165 18960 16210 19010
rect 16260 18960 16305 19010
rect 16355 18960 16425 19010
rect 16475 18960 16520 19010
rect 16570 18960 16615 19010
rect 16665 18960 16715 19010
rect 16765 18960 16815 19010
rect 16865 18960 16915 19010
rect 16965 18960 17010 19010
rect 17060 18960 17105 19010
rect 17155 18960 17225 19010
rect 17275 18960 17320 19010
rect 17370 18960 17415 19010
rect 17465 18960 17515 19010
rect 17565 18960 17615 19010
rect 17665 18960 17715 19010
rect 17765 18960 17810 19010
rect 17860 18960 17905 19010
rect 17955 18960 17990 19010
rect 6740 18935 17990 18960
rect 2320 18915 17990 18935
rect 2320 18875 2330 18915
rect 2370 18875 6700 18915
rect 6740 18890 17990 18915
rect 6740 18875 14825 18890
rect 2320 18850 14825 18875
rect 2320 18810 2330 18850
rect 2370 18810 6700 18850
rect 6740 18840 14825 18850
rect 14875 18840 14920 18890
rect 14970 18840 15015 18890
rect 15065 18840 15115 18890
rect 15165 18840 15215 18890
rect 15265 18840 15315 18890
rect 15365 18840 15410 18890
rect 15460 18840 15505 18890
rect 15555 18840 15625 18890
rect 15675 18840 15720 18890
rect 15770 18840 15815 18890
rect 15865 18840 15915 18890
rect 15965 18840 16015 18890
rect 16065 18840 16115 18890
rect 16165 18840 16210 18890
rect 16260 18840 16305 18890
rect 16355 18840 16425 18890
rect 16475 18840 16520 18890
rect 16570 18840 16615 18890
rect 16665 18840 16715 18890
rect 16765 18840 16815 18890
rect 16865 18840 16915 18890
rect 16965 18840 17010 18890
rect 17060 18840 17105 18890
rect 17155 18840 17225 18890
rect 17275 18840 17320 18890
rect 17370 18840 17415 18890
rect 17465 18840 17515 18890
rect 17565 18840 17615 18890
rect 17665 18840 17715 18890
rect 17765 18840 17810 18890
rect 17860 18840 17905 18890
rect 17955 18840 17990 18890
rect 6740 18810 17990 18840
rect 2320 18800 17990 18810
rect 2320 18780 14825 18800
rect 2320 18740 2330 18780
rect 2370 18740 6700 18780
rect 6740 18750 14825 18780
rect 14875 18750 14920 18800
rect 14970 18750 15015 18800
rect 15065 18750 15115 18800
rect 15165 18750 15215 18800
rect 15265 18750 15315 18800
rect 15365 18750 15410 18800
rect 15460 18750 15505 18800
rect 15555 18750 15625 18800
rect 15675 18750 15720 18800
rect 15770 18750 15815 18800
rect 15865 18750 15915 18800
rect 15965 18750 16015 18800
rect 16065 18750 16115 18800
rect 16165 18750 16210 18800
rect 16260 18750 16305 18800
rect 16355 18750 16425 18800
rect 16475 18750 16520 18800
rect 16570 18750 16615 18800
rect 16665 18750 16715 18800
rect 16765 18750 16815 18800
rect 16865 18750 16915 18800
rect 16965 18750 17010 18800
rect 17060 18750 17105 18800
rect 17155 18750 17225 18800
rect 17275 18750 17320 18800
rect 17370 18750 17415 18800
rect 17465 18750 17515 18800
rect 17565 18750 17615 18800
rect 17665 18750 17715 18800
rect 17765 18750 17810 18800
rect 17860 18750 17905 18800
rect 17955 18750 17990 18800
rect 6740 18740 17990 18750
rect 2320 18710 17990 18740
rect 2320 18670 2330 18710
rect 2370 18670 6700 18710
rect 6740 18700 17990 18710
rect 6740 18670 14825 18700
rect 2320 18650 14825 18670
rect 14875 18650 14920 18700
rect 14970 18650 15015 18700
rect 15065 18650 15115 18700
rect 15165 18650 15215 18700
rect 15265 18650 15315 18700
rect 15365 18650 15410 18700
rect 15460 18650 15505 18700
rect 15555 18650 15625 18700
rect 15675 18650 15720 18700
rect 15770 18650 15815 18700
rect 15865 18650 15915 18700
rect 15965 18650 16015 18700
rect 16065 18650 16115 18700
rect 16165 18650 16210 18700
rect 16260 18650 16305 18700
rect 16355 18650 16425 18700
rect 16475 18650 16520 18700
rect 16570 18650 16615 18700
rect 16665 18650 16715 18700
rect 16765 18650 16815 18700
rect 16865 18650 16915 18700
rect 16965 18650 17010 18700
rect 17060 18650 17105 18700
rect 17155 18650 17225 18700
rect 17275 18650 17320 18700
rect 17370 18650 17415 18700
rect 17465 18650 17515 18700
rect 17565 18650 17615 18700
rect 17665 18650 17715 18700
rect 17765 18650 17810 18700
rect 17860 18650 17905 18700
rect 17955 18650 17990 18700
rect 2320 18640 17990 18650
rect 2320 18600 2330 18640
rect 2370 18600 6700 18640
rect 6740 18610 17990 18640
rect 6740 18600 14825 18610
rect 2320 18575 14825 18600
rect 2320 18535 2330 18575
rect 2370 18535 6700 18575
rect 6740 18560 14825 18575
rect 14875 18560 14920 18610
rect 14970 18560 15015 18610
rect 15065 18560 15115 18610
rect 15165 18560 15215 18610
rect 15265 18560 15315 18610
rect 15365 18560 15410 18610
rect 15460 18560 15505 18610
rect 15555 18560 15625 18610
rect 15675 18560 15720 18610
rect 15770 18560 15815 18610
rect 15865 18560 15915 18610
rect 15965 18560 16015 18610
rect 16065 18560 16115 18610
rect 16165 18560 16210 18610
rect 16260 18560 16305 18610
rect 16355 18560 16425 18610
rect 16475 18560 16520 18610
rect 16570 18560 16615 18610
rect 16665 18560 16715 18610
rect 16765 18560 16815 18610
rect 16865 18560 16915 18610
rect 16965 18560 17010 18610
rect 17060 18560 17105 18610
rect 17155 18560 17225 18610
rect 17275 18560 17320 18610
rect 17370 18560 17415 18610
rect 17465 18560 17515 18610
rect 17565 18560 17615 18610
rect 17665 18560 17715 18610
rect 17765 18560 17810 18610
rect 17860 18560 17905 18610
rect 17955 18560 17990 18610
rect 6740 18535 17990 18560
rect 2320 18515 17990 18535
rect 2320 18475 2330 18515
rect 2370 18475 6700 18515
rect 6740 18490 17990 18515
rect 6740 18475 14825 18490
rect 2320 18450 14825 18475
rect 2320 18410 2330 18450
rect 2370 18410 6700 18450
rect 6740 18440 14825 18450
rect 14875 18440 14920 18490
rect 14970 18440 15015 18490
rect 15065 18440 15115 18490
rect 15165 18440 15215 18490
rect 15265 18440 15315 18490
rect 15365 18440 15410 18490
rect 15460 18440 15505 18490
rect 15555 18440 15625 18490
rect 15675 18440 15720 18490
rect 15770 18440 15815 18490
rect 15865 18440 15915 18490
rect 15965 18440 16015 18490
rect 16065 18440 16115 18490
rect 16165 18440 16210 18490
rect 16260 18440 16305 18490
rect 16355 18440 16425 18490
rect 16475 18440 16520 18490
rect 16570 18440 16615 18490
rect 16665 18440 16715 18490
rect 16765 18440 16815 18490
rect 16865 18440 16915 18490
rect 16965 18440 17010 18490
rect 17060 18440 17105 18490
rect 17155 18440 17225 18490
rect 17275 18440 17320 18490
rect 17370 18440 17415 18490
rect 17465 18440 17515 18490
rect 17565 18440 17615 18490
rect 17665 18440 17715 18490
rect 17765 18440 17810 18490
rect 17860 18440 17905 18490
rect 17955 18440 17990 18490
rect 6740 18410 17990 18440
rect 2320 18400 17990 18410
rect 2320 18380 14825 18400
rect 2320 18340 2330 18380
rect 2370 18340 6700 18380
rect 6740 18350 14825 18380
rect 14875 18350 14920 18400
rect 14970 18350 15015 18400
rect 15065 18350 15115 18400
rect 15165 18350 15215 18400
rect 15265 18350 15315 18400
rect 15365 18350 15410 18400
rect 15460 18350 15505 18400
rect 15555 18350 15625 18400
rect 15675 18350 15720 18400
rect 15770 18350 15815 18400
rect 15865 18350 15915 18400
rect 15965 18350 16015 18400
rect 16065 18350 16115 18400
rect 16165 18350 16210 18400
rect 16260 18350 16305 18400
rect 16355 18350 16425 18400
rect 16475 18350 16520 18400
rect 16570 18350 16615 18400
rect 16665 18350 16715 18400
rect 16765 18350 16815 18400
rect 16865 18350 16915 18400
rect 16965 18350 17010 18400
rect 17060 18350 17105 18400
rect 17155 18350 17225 18400
rect 17275 18350 17320 18400
rect 17370 18350 17415 18400
rect 17465 18350 17515 18400
rect 17565 18350 17615 18400
rect 17665 18350 17715 18400
rect 17765 18350 17810 18400
rect 17860 18350 17905 18400
rect 17955 18350 17990 18400
rect 6740 18340 17990 18350
rect 2320 18310 17990 18340
rect 2320 18270 2330 18310
rect 2370 18270 6700 18310
rect 6740 18300 17990 18310
rect 6740 18270 14825 18300
rect 2320 18250 14825 18270
rect 14875 18250 14920 18300
rect 14970 18250 15015 18300
rect 15065 18250 15115 18300
rect 15165 18250 15215 18300
rect 15265 18250 15315 18300
rect 15365 18250 15410 18300
rect 15460 18250 15505 18300
rect 15555 18250 15625 18300
rect 15675 18250 15720 18300
rect 15770 18250 15815 18300
rect 15865 18250 15915 18300
rect 15965 18250 16015 18300
rect 16065 18250 16115 18300
rect 16165 18250 16210 18300
rect 16260 18250 16305 18300
rect 16355 18250 16425 18300
rect 16475 18250 16520 18300
rect 16570 18250 16615 18300
rect 16665 18250 16715 18300
rect 16765 18250 16815 18300
rect 16865 18250 16915 18300
rect 16965 18250 17010 18300
rect 17060 18250 17105 18300
rect 17155 18250 17225 18300
rect 17275 18250 17320 18300
rect 17370 18250 17415 18300
rect 17465 18250 17515 18300
rect 17565 18250 17615 18300
rect 17665 18250 17715 18300
rect 17765 18250 17810 18300
rect 17860 18250 17905 18300
rect 17955 18250 17990 18300
rect 2320 18240 17990 18250
rect 2320 18200 2330 18240
rect 2370 18200 6700 18240
rect 6740 18210 17990 18240
rect 6740 18200 14825 18210
rect 2320 18175 14825 18200
rect 2320 18145 2330 18175
rect -1170 18140 2330 18145
rect -1170 18100 -1165 18140
rect -1125 18100 -815 18140
rect -775 18100 -465 18140
rect -425 18100 -115 18140
rect -75 18100 235 18140
rect 275 18100 585 18140
rect 625 18100 935 18140
rect 975 18100 1285 18140
rect 1325 18100 1635 18140
rect 1675 18135 2330 18140
rect 2370 18135 6700 18175
rect 6740 18160 14825 18175
rect 14875 18160 14920 18210
rect 14970 18160 15015 18210
rect 15065 18160 15115 18210
rect 15165 18160 15215 18210
rect 15265 18160 15315 18210
rect 15365 18160 15410 18210
rect 15460 18160 15505 18210
rect 15555 18160 15625 18210
rect 15675 18160 15720 18210
rect 15770 18160 15815 18210
rect 15865 18160 15915 18210
rect 15965 18160 16015 18210
rect 16065 18160 16115 18210
rect 16165 18160 16210 18210
rect 16260 18160 16305 18210
rect 16355 18160 16425 18210
rect 16475 18160 16520 18210
rect 16570 18160 16615 18210
rect 16665 18160 16715 18210
rect 16765 18160 16815 18210
rect 16865 18160 16915 18210
rect 16965 18160 17010 18210
rect 17060 18160 17105 18210
rect 17155 18160 17225 18210
rect 17275 18160 17320 18210
rect 17370 18160 17415 18210
rect 17465 18160 17515 18210
rect 17565 18160 17615 18210
rect 17665 18160 17715 18210
rect 17765 18160 17810 18210
rect 17860 18160 17905 18210
rect 17955 18160 17990 18210
rect 6740 18135 17990 18160
rect 1675 18115 17990 18135
rect 1675 18100 2330 18115
rect -1170 18095 2330 18100
rect 230 17795 280 18095
rect 2320 18075 2330 18095
rect 2370 18075 6700 18115
rect 6740 18090 17990 18115
rect 6740 18075 14825 18090
rect 2320 18050 14825 18075
rect 2320 18010 2330 18050
rect 2370 18010 6700 18050
rect 6740 18040 14825 18050
rect 14875 18040 14920 18090
rect 14970 18040 15015 18090
rect 15065 18040 15115 18090
rect 15165 18040 15215 18090
rect 15265 18040 15315 18090
rect 15365 18040 15410 18090
rect 15460 18040 15505 18090
rect 15555 18040 15625 18090
rect 15675 18040 15720 18090
rect 15770 18040 15815 18090
rect 15865 18040 15915 18090
rect 15965 18040 16015 18090
rect 16065 18040 16115 18090
rect 16165 18040 16210 18090
rect 16260 18040 16305 18090
rect 16355 18040 16425 18090
rect 16475 18040 16520 18090
rect 16570 18040 16615 18090
rect 16665 18040 16715 18090
rect 16765 18040 16815 18090
rect 16865 18040 16915 18090
rect 16965 18040 17010 18090
rect 17060 18040 17105 18090
rect 17155 18040 17225 18090
rect 17275 18040 17320 18090
rect 17370 18040 17415 18090
rect 17465 18040 17515 18090
rect 17565 18040 17615 18090
rect 17665 18040 17715 18090
rect 17765 18040 17810 18090
rect 17860 18040 17905 18090
rect 17955 18040 17990 18090
rect 6740 18010 17990 18040
rect 2320 18000 17990 18010
rect 2320 17980 14825 18000
rect 2320 17940 2330 17980
rect 2370 17940 6700 17980
rect 6740 17950 14825 17980
rect 14875 17950 14920 18000
rect 14970 17950 15015 18000
rect 15065 17950 15115 18000
rect 15165 17950 15215 18000
rect 15265 17950 15315 18000
rect 15365 17950 15410 18000
rect 15460 17950 15505 18000
rect 15555 17950 15625 18000
rect 15675 17950 15720 18000
rect 15770 17950 15815 18000
rect 15865 17950 15915 18000
rect 15965 17950 16015 18000
rect 16065 17950 16115 18000
rect 16165 17950 16210 18000
rect 16260 17950 16305 18000
rect 16355 17950 16425 18000
rect 16475 17950 16520 18000
rect 16570 17950 16615 18000
rect 16665 17950 16715 18000
rect 16765 17950 16815 18000
rect 16865 17950 16915 18000
rect 16965 17950 17010 18000
rect 17060 17950 17105 18000
rect 17155 17950 17225 18000
rect 17275 17950 17320 18000
rect 17370 17950 17415 18000
rect 17465 17950 17515 18000
rect 17565 17950 17615 18000
rect 17665 17950 17715 18000
rect 17765 17950 17810 18000
rect 17860 17950 17905 18000
rect 17955 17950 17990 18000
rect 6740 17940 17990 17950
rect 2320 17910 17990 17940
rect 2320 17870 2330 17910
rect 2370 17870 6700 17910
rect 6740 17900 17990 17910
rect 6740 17870 14825 17900
rect 2320 17850 14825 17870
rect 14875 17850 14920 17900
rect 14970 17850 15015 17900
rect 15065 17850 15115 17900
rect 15165 17850 15215 17900
rect 15265 17850 15315 17900
rect 15365 17850 15410 17900
rect 15460 17850 15505 17900
rect 15555 17850 15625 17900
rect 15675 17850 15720 17900
rect 15770 17850 15815 17900
rect 15865 17850 15915 17900
rect 15965 17850 16015 17900
rect 16065 17850 16115 17900
rect 16165 17850 16210 17900
rect 16260 17850 16305 17900
rect 16355 17850 16425 17900
rect 16475 17850 16520 17900
rect 16570 17850 16615 17900
rect 16665 17850 16715 17900
rect 16765 17850 16815 17900
rect 16865 17850 16915 17900
rect 16965 17850 17010 17900
rect 17060 17850 17105 17900
rect 17155 17850 17225 17900
rect 17275 17850 17320 17900
rect 17370 17850 17415 17900
rect 17465 17850 17515 17900
rect 17565 17850 17615 17900
rect 17665 17850 17715 17900
rect 17765 17850 17810 17900
rect 17860 17850 17905 17900
rect 17955 17850 17990 17900
rect 2320 17840 17990 17850
rect 2320 17800 2330 17840
rect 2370 17800 6700 17840
rect 6740 17810 17990 17840
rect 6740 17800 14825 17810
rect -1170 17790 1680 17795
rect -1170 17750 -1165 17790
rect -1125 17750 -815 17790
rect -775 17750 -465 17790
rect -425 17750 -115 17790
rect -75 17750 235 17790
rect 275 17750 585 17790
rect 625 17750 935 17790
rect 975 17750 1285 17790
rect 1325 17750 1635 17790
rect 1675 17750 1680 17790
rect -1170 17745 1680 17750
rect 2320 17775 14825 17800
rect 230 17445 280 17745
rect 2320 17735 2330 17775
rect 2370 17735 6700 17775
rect 6740 17760 14825 17775
rect 14875 17760 14920 17810
rect 14970 17760 15015 17810
rect 15065 17760 15115 17810
rect 15165 17760 15215 17810
rect 15265 17760 15315 17810
rect 15365 17760 15410 17810
rect 15460 17760 15505 17810
rect 15555 17760 15625 17810
rect 15675 17760 15720 17810
rect 15770 17760 15815 17810
rect 15865 17760 15915 17810
rect 15965 17760 16015 17810
rect 16065 17760 16115 17810
rect 16165 17760 16210 17810
rect 16260 17760 16305 17810
rect 16355 17760 16425 17810
rect 16475 17760 16520 17810
rect 16570 17760 16615 17810
rect 16665 17760 16715 17810
rect 16765 17760 16815 17810
rect 16865 17760 16915 17810
rect 16965 17760 17010 17810
rect 17060 17760 17105 17810
rect 17155 17760 17225 17810
rect 17275 17760 17320 17810
rect 17370 17760 17415 17810
rect 17465 17760 17515 17810
rect 17565 17760 17615 17810
rect 17665 17760 17715 17810
rect 17765 17760 17810 17810
rect 17860 17760 17905 17810
rect 17955 17760 17990 17810
rect 6740 17735 17990 17760
rect 2320 17725 17990 17735
rect -1170 17440 1680 17445
rect -1170 17400 -1165 17440
rect -1125 17400 -815 17440
rect -775 17400 -465 17440
rect -425 17400 -115 17440
rect -75 17400 235 17440
rect 275 17400 585 17440
rect 625 17400 935 17440
rect 975 17400 1285 17440
rect 1325 17400 1635 17440
rect 1675 17400 1680 17440
rect -1170 17395 1680 17400
rect 9630 17440 14580 17445
rect 9630 17400 9635 17440
rect 9675 17400 9985 17440
rect 10025 17400 10335 17440
rect 10375 17400 10685 17440
rect 10725 17400 11035 17440
rect 11075 17400 11385 17440
rect 11425 17400 11735 17440
rect 11775 17400 12085 17440
rect 12125 17400 12435 17440
rect 12475 17400 12785 17440
rect 12825 17400 13135 17440
rect 13175 17400 13485 17440
rect 13525 17400 13835 17440
rect 13875 17400 14185 17440
rect 14225 17400 14535 17440
rect 14575 17400 14580 17440
rect 9630 17395 14580 17400
rect 230 17095 280 17395
rect 12080 17095 12130 17395
rect -1170 17090 1680 17095
rect -1170 17050 -1165 17090
rect -1125 17050 -815 17090
rect -775 17050 -465 17090
rect -425 17050 -115 17090
rect -75 17050 235 17090
rect 275 17050 585 17090
rect 625 17050 935 17090
rect 975 17050 1285 17090
rect 1325 17050 1635 17090
rect 1675 17050 1680 17090
rect -1170 17045 1680 17050
rect 9630 17090 14580 17095
rect 9630 17050 9635 17090
rect 9675 17050 9985 17090
rect 10025 17050 10335 17090
rect 10375 17050 10685 17090
rect 10725 17050 11035 17090
rect 11075 17050 11385 17090
rect 11425 17050 11735 17090
rect 11775 17050 12085 17090
rect 12125 17050 12435 17090
rect 12475 17050 12785 17090
rect 12825 17050 13135 17090
rect 13175 17050 13485 17090
rect 13525 17050 13835 17090
rect 13875 17050 14185 17090
rect 14225 17050 14535 17090
rect 14575 17050 14580 17090
rect 9630 17045 14580 17050
rect 230 16745 280 17045
rect 12080 16745 12130 17045
rect -1170 16740 1680 16745
rect -1170 16700 -1165 16740
rect -1125 16700 -815 16740
rect -775 16700 -465 16740
rect -425 16700 -115 16740
rect -75 16700 235 16740
rect 275 16700 585 16740
rect 625 16700 935 16740
rect 975 16700 1285 16740
rect 1325 16700 1635 16740
rect 1675 16700 1680 16740
rect -1170 16695 1680 16700
rect 9630 16740 14580 16745
rect 9630 16700 9635 16740
rect 9675 16700 9985 16740
rect 10025 16700 10335 16740
rect 10375 16700 10685 16740
rect 10725 16700 11035 16740
rect 11075 16700 11385 16740
rect 11425 16700 11735 16740
rect 11775 16700 12085 16740
rect 12125 16700 12435 16740
rect 12475 16700 12785 16740
rect 12825 16700 13135 16740
rect 13175 16700 13485 16740
rect 13525 16700 13835 16740
rect 13875 16700 14185 16740
rect 14225 16700 14535 16740
rect 14575 16700 14580 16740
rect 9630 16695 14580 16700
rect 230 16395 280 16695
rect 12080 16395 12130 16695
rect -1170 16390 1680 16395
rect -1170 16350 -1165 16390
rect -1125 16350 -815 16390
rect -775 16350 -465 16390
rect -425 16350 -115 16390
rect -75 16350 235 16390
rect 275 16350 585 16390
rect 625 16350 935 16390
rect 975 16350 1285 16390
rect 1325 16350 1635 16390
rect 1675 16350 1680 16390
rect -1170 16345 1680 16350
rect 9630 16390 14580 16395
rect 9630 16350 9635 16390
rect 9675 16350 9985 16390
rect 10025 16350 10335 16390
rect 10375 16350 10685 16390
rect 10725 16350 11035 16390
rect 11075 16350 11385 16390
rect 11425 16350 11735 16390
rect 11775 16350 12085 16390
rect 12125 16350 12435 16390
rect 12475 16350 12785 16390
rect 12825 16350 13135 16390
rect 13175 16350 13485 16390
rect 13525 16350 13835 16390
rect 13875 16350 14185 16390
rect 14225 16350 14535 16390
rect 14575 16350 14580 16390
rect 9630 16345 14580 16350
rect 230 16045 280 16345
rect 12080 16045 12130 16345
rect -1170 16040 1680 16045
rect -1170 16000 -1165 16040
rect -1125 16000 -815 16040
rect -775 16000 -465 16040
rect -425 16000 -115 16040
rect -75 16000 235 16040
rect 275 16000 585 16040
rect 625 16000 935 16040
rect 975 16000 1285 16040
rect 1325 16000 1635 16040
rect 1675 16000 1680 16040
rect -1170 15995 1680 16000
rect 9630 16040 14580 16045
rect 9630 16000 9635 16040
rect 9675 16000 9985 16040
rect 10025 16000 10335 16040
rect 10375 16000 10685 16040
rect 10725 16000 11035 16040
rect 11075 16000 11385 16040
rect 11425 16000 11735 16040
rect 11775 16000 12085 16040
rect 12125 16000 12435 16040
rect 12475 16000 12785 16040
rect 12825 16000 13135 16040
rect 13175 16000 13485 16040
rect 13525 16000 13835 16040
rect 13875 16000 14185 16040
rect 14225 16000 14535 16040
rect 14575 16000 14580 16040
rect 9630 15995 14580 16000
rect 230 15695 280 15995
rect 12080 15695 12130 15995
rect -1170 15690 1680 15695
rect -1170 15650 -1165 15690
rect -1125 15650 -815 15690
rect -775 15650 -465 15690
rect -425 15650 -115 15690
rect -75 15650 235 15690
rect 275 15650 585 15690
rect 625 15650 935 15690
rect 975 15650 1285 15690
rect 1325 15650 1635 15690
rect 1675 15650 1680 15690
rect -1170 15645 1680 15650
rect 9630 15690 14580 15695
rect 9630 15650 9635 15690
rect 9675 15650 9985 15690
rect 10025 15650 10335 15690
rect 10375 15650 10685 15690
rect 10725 15650 11035 15690
rect 11075 15650 11385 15690
rect 11425 15650 11735 15690
rect 11775 15650 12085 15690
rect 12125 15650 12435 15690
rect 12475 15650 12785 15690
rect 12825 15650 13135 15690
rect 13175 15650 13485 15690
rect 13525 15650 13835 15690
rect 13875 15650 14185 15690
rect 14225 15650 14535 15690
rect 14575 15650 14580 15690
rect 9630 15645 14580 15650
rect 230 15345 280 15645
rect 12080 15345 12130 15645
rect -1170 15340 1680 15345
rect -1170 15300 -1165 15340
rect -1125 15300 -815 15340
rect -775 15300 -465 15340
rect -425 15300 -115 15340
rect -75 15300 235 15340
rect 275 15300 585 15340
rect 625 15300 935 15340
rect 975 15300 1285 15340
rect 1325 15300 1635 15340
rect 1675 15300 1680 15340
rect -1170 15295 1680 15300
rect 9630 15340 14580 15345
rect 9630 15300 9635 15340
rect 9675 15300 9985 15340
rect 10025 15300 10335 15340
rect 10375 15300 10685 15340
rect 10725 15300 11035 15340
rect 11075 15300 11385 15340
rect 11425 15300 11735 15340
rect 11775 15300 12085 15340
rect 12125 15300 12435 15340
rect 12475 15300 12785 15340
rect 12825 15300 13135 15340
rect 13175 15300 13485 15340
rect 13525 15300 13835 15340
rect 13875 15300 14185 15340
rect 14225 15300 14535 15340
rect 14575 15300 14580 15340
rect 9630 15295 14580 15300
rect 230 14995 280 15295
rect 12080 14995 12130 15295
rect -1170 14990 1680 14995
rect -1170 14950 -1165 14990
rect -1125 14950 -815 14990
rect -775 14950 -465 14990
rect -425 14950 -115 14990
rect -75 14950 235 14990
rect 275 14950 585 14990
rect 625 14950 935 14990
rect 975 14950 1285 14990
rect 1325 14950 1635 14990
rect 1675 14950 1680 14990
rect -1170 14945 1680 14950
rect 9630 14990 14580 14995
rect 9630 14950 9635 14990
rect 9675 14950 9985 14990
rect 10025 14950 10335 14990
rect 10375 14950 10685 14990
rect 10725 14950 11035 14990
rect 11075 14950 11385 14990
rect 11425 14950 11735 14990
rect 11775 14950 12085 14990
rect 12125 14950 12435 14990
rect 12475 14950 12785 14990
rect 12825 14950 13135 14990
rect 13175 14950 13485 14990
rect 13525 14950 13835 14990
rect 13875 14950 14185 14990
rect 14225 14950 14535 14990
rect 14575 14950 14580 14990
rect 9630 14945 14580 14950
rect 230 14645 280 14945
rect 12080 14645 12130 14945
rect -1170 14640 1680 14645
rect -1170 14600 -1165 14640
rect -1125 14600 -815 14640
rect -775 14600 -465 14640
rect -425 14600 -115 14640
rect -75 14600 235 14640
rect 275 14600 585 14640
rect 625 14600 935 14640
rect 975 14600 1285 14640
rect 1325 14600 1635 14640
rect 1675 14600 1680 14640
rect -1170 14595 1680 14600
rect 9630 14640 14580 14645
rect 9630 14600 9635 14640
rect 9675 14600 9985 14640
rect 10025 14600 10335 14640
rect 10375 14600 10685 14640
rect 10725 14600 11035 14640
rect 11075 14600 11385 14640
rect 11425 14600 11735 14640
rect 11775 14600 12085 14640
rect 12125 14600 12435 14640
rect 12475 14600 12785 14640
rect 12825 14600 13135 14640
rect 13175 14600 13485 14640
rect 13525 14600 13835 14640
rect 13875 14600 14185 14640
rect 14225 14600 14535 14640
rect 14575 14600 14580 14640
rect 9630 14595 14580 14600
rect 230 14295 280 14595
rect 12080 14295 12130 14595
rect -1170 14290 1680 14295
rect -1170 14250 -1165 14290
rect -1125 14250 -815 14290
rect -775 14250 -465 14290
rect -425 14250 -115 14290
rect -75 14250 235 14290
rect 275 14250 585 14290
rect 625 14250 935 14290
rect 975 14250 1285 14290
rect 1325 14250 1635 14290
rect 1675 14250 1680 14290
rect -1170 14245 1680 14250
rect 9630 14290 14580 14295
rect 9630 14250 9635 14290
rect 9675 14250 9985 14290
rect 10025 14250 10335 14290
rect 10375 14250 10685 14290
rect 10725 14250 11035 14290
rect 11075 14250 11385 14290
rect 11425 14250 11735 14290
rect 11775 14250 12085 14290
rect 12125 14250 12435 14290
rect 12475 14250 12785 14290
rect 12825 14250 13135 14290
rect 13175 14250 13485 14290
rect 13525 14250 13835 14290
rect 13875 14250 14185 14290
rect 14225 14250 14535 14290
rect 14575 14250 14580 14290
rect 9630 14245 14580 14250
rect 230 13945 280 14245
rect 12080 13945 12130 14245
rect -1170 13940 1680 13945
rect -1170 13900 -1165 13940
rect -1125 13900 -815 13940
rect -775 13900 -465 13940
rect -425 13900 -115 13940
rect -75 13900 235 13940
rect 275 13900 585 13940
rect 625 13900 935 13940
rect 975 13900 1285 13940
rect 1325 13900 1635 13940
rect 1675 13900 1680 13940
rect -1170 13895 1680 13900
rect 9630 13940 14580 13945
rect 9630 13900 9635 13940
rect 9675 13900 9985 13940
rect 10025 13900 10335 13940
rect 10375 13900 10685 13940
rect 10725 13900 11035 13940
rect 11075 13900 11385 13940
rect 11425 13900 11735 13940
rect 11775 13900 12085 13940
rect 12125 13900 12435 13940
rect 12475 13900 12785 13940
rect 12825 13900 13135 13940
rect 13175 13900 13485 13940
rect 13525 13900 13835 13940
rect 13875 13900 14185 13940
rect 14225 13900 14535 13940
rect 14575 13900 14580 13940
rect 9630 13895 14580 13900
rect 230 13595 280 13895
rect 12080 13595 12130 13895
rect -1170 13590 1680 13595
rect -1170 13550 -1165 13590
rect -1125 13550 -815 13590
rect -775 13550 -465 13590
rect -425 13550 -115 13590
rect -75 13550 235 13590
rect 275 13550 585 13590
rect 625 13550 935 13590
rect 975 13550 1285 13590
rect 1325 13550 1635 13590
rect 1675 13550 1680 13590
rect -1170 13545 1680 13550
rect 9630 13590 14580 13595
rect 9630 13550 9635 13590
rect 9675 13550 9985 13590
rect 10025 13550 10335 13590
rect 10375 13550 10685 13590
rect 10725 13550 11035 13590
rect 11075 13550 11385 13590
rect 11425 13550 11735 13590
rect 11775 13550 12085 13590
rect 12125 13550 12435 13590
rect 12475 13550 12785 13590
rect 12825 13550 13135 13590
rect 13175 13550 13485 13590
rect 13525 13550 13835 13590
rect 13875 13550 14185 13590
rect 14225 13550 14535 13590
rect 14575 13550 14580 13590
rect 9630 13545 14580 13550
rect 230 13245 280 13545
rect 12080 13245 12130 13545
rect -1170 13240 1680 13245
rect -1170 13200 -1165 13240
rect -1125 13200 -815 13240
rect -775 13200 -465 13240
rect -425 13200 -115 13240
rect -75 13200 235 13240
rect 275 13200 585 13240
rect 625 13200 935 13240
rect 975 13200 1285 13240
rect 1325 13200 1635 13240
rect 1675 13200 1680 13240
rect -1170 13195 1680 13200
rect 9630 13240 14580 13245
rect 9630 13200 9635 13240
rect 9675 13200 9985 13240
rect 10025 13200 10335 13240
rect 10375 13200 10685 13240
rect 10725 13200 11035 13240
rect 11075 13200 11385 13240
rect 11425 13200 11735 13240
rect 11775 13200 12085 13240
rect 12125 13200 12435 13240
rect 12475 13200 12785 13240
rect 12825 13200 13135 13240
rect 13175 13200 13485 13240
rect 13525 13200 13835 13240
rect 13875 13200 14185 13240
rect 14225 13200 14535 13240
rect 14575 13200 14580 13240
rect 9630 13195 14580 13200
rect 230 12895 280 13195
rect 12080 12895 12130 13195
rect -1170 12890 1680 12895
rect -1170 12850 -1165 12890
rect -1125 12850 -815 12890
rect -775 12850 -465 12890
rect -425 12850 -115 12890
rect -75 12850 235 12890
rect 275 12850 585 12890
rect 625 12850 935 12890
rect 975 12850 1285 12890
rect 1325 12850 1635 12890
rect 1675 12850 1680 12890
rect -1170 12845 1680 12850
rect 9630 12890 14580 12895
rect 9630 12850 9635 12890
rect 9675 12850 9985 12890
rect 10025 12850 10335 12890
rect 10375 12850 10685 12890
rect 10725 12850 11035 12890
rect 11075 12850 11385 12890
rect 11425 12850 11735 12890
rect 11775 12850 12085 12890
rect 12125 12850 12435 12890
rect 12475 12850 12785 12890
rect 12825 12850 13135 12890
rect 13175 12850 13485 12890
rect 13525 12850 13835 12890
rect 13875 12850 14185 12890
rect 14225 12850 14535 12890
rect 14575 12850 14580 12890
rect 9630 12845 14580 12850
rect 230 12545 280 12845
rect 12080 12545 12130 12845
rect -1170 12540 1680 12545
rect -1170 12500 -1165 12540
rect -1125 12500 -815 12540
rect -775 12500 -465 12540
rect -425 12500 -115 12540
rect -75 12500 235 12540
rect 275 12500 585 12540
rect 625 12500 935 12540
rect 975 12500 1285 12540
rect 1325 12500 1635 12540
rect 1675 12500 1680 12540
rect -1170 12495 1680 12500
rect 9630 12540 14580 12545
rect 9630 12500 9635 12540
rect 9675 12500 9985 12540
rect 10025 12500 10335 12540
rect 10375 12500 10685 12540
rect 10725 12500 11035 12540
rect 11075 12500 11385 12540
rect 11425 12500 11735 12540
rect 11775 12500 12085 12540
rect 12125 12500 12435 12540
rect 12475 12500 12785 12540
rect 12825 12500 13135 12540
rect 13175 12500 13485 12540
rect 13525 12500 13835 12540
rect 13875 12500 14185 12540
rect 14225 12500 14535 12540
rect 14575 12500 14580 12540
rect 9630 12495 14580 12500
rect 230 12195 280 12495
rect 12080 12195 12130 12495
rect -1170 12190 1680 12195
rect -1170 12150 -1165 12190
rect -1125 12150 -815 12190
rect -775 12150 -465 12190
rect -425 12150 -115 12190
rect -75 12150 235 12190
rect 275 12150 585 12190
rect 625 12150 935 12190
rect 975 12150 1285 12190
rect 1325 12150 1635 12190
rect 1675 12150 1680 12190
rect -1170 12145 1680 12150
rect 9630 12190 14580 12195
rect 9630 12150 9635 12190
rect 9675 12150 9985 12190
rect 10025 12150 10335 12190
rect 10375 12150 10685 12190
rect 10725 12150 11035 12190
rect 11075 12150 11385 12190
rect 11425 12150 11735 12190
rect 11775 12150 12085 12190
rect 12125 12150 12435 12190
rect 12475 12150 12785 12190
rect 12825 12150 13135 12190
rect 13175 12150 13485 12190
rect 13525 12150 13835 12190
rect 13875 12150 14185 12190
rect 14225 12150 14535 12190
rect 14575 12150 14580 12190
rect 9630 12145 14580 12150
rect 230 11845 280 12145
rect 12080 11845 12130 12145
rect -1170 11840 1680 11845
rect -1170 11800 -1165 11840
rect -1125 11800 -815 11840
rect -775 11800 -465 11840
rect -425 11800 -115 11840
rect -75 11800 235 11840
rect 275 11800 585 11840
rect 625 11800 935 11840
rect 975 11800 1285 11840
rect 1325 11800 1635 11840
rect 1675 11800 1680 11840
rect -1170 11795 1680 11800
rect 9630 11840 14580 11845
rect 9630 11800 9635 11840
rect 9675 11800 9985 11840
rect 10025 11800 10335 11840
rect 10375 11800 10685 11840
rect 10725 11800 11035 11840
rect 11075 11800 11385 11840
rect 11425 11800 11735 11840
rect 11775 11800 12085 11840
rect 12125 11800 12435 11840
rect 12475 11800 12785 11840
rect 12825 11800 13135 11840
rect 13175 11800 13485 11840
rect 13525 11800 13835 11840
rect 13875 11800 14185 11840
rect 14225 11800 14535 11840
rect 14575 11800 14580 11840
rect 9630 11795 14580 11800
rect 230 11495 280 11795
rect 12080 11495 12130 11795
rect -1170 11490 1680 11495
rect -1170 11450 -1165 11490
rect -1125 11450 -815 11490
rect -775 11450 -465 11490
rect -425 11450 -115 11490
rect -75 11450 235 11490
rect 275 11450 585 11490
rect 625 11450 935 11490
rect 975 11450 1285 11490
rect 1325 11450 1635 11490
rect 1675 11450 1680 11490
rect -1170 11445 1680 11450
rect 9630 11490 14580 11495
rect 9630 11450 9635 11490
rect 9675 11450 9985 11490
rect 10025 11450 10335 11490
rect 10375 11450 10685 11490
rect 10725 11450 11035 11490
rect 11075 11450 11385 11490
rect 11425 11450 11735 11490
rect 11775 11450 12085 11490
rect 12125 11450 12435 11490
rect 12475 11450 12785 11490
rect 12825 11450 13135 11490
rect 13175 11450 13485 11490
rect 13525 11450 13835 11490
rect 13875 11450 14185 11490
rect 14225 11450 14535 11490
rect 14575 11450 14580 11490
rect 9630 11445 14580 11450
rect 230 11145 280 11445
rect 12080 11145 12130 11445
rect -1170 11140 1680 11145
rect -1170 11100 -1165 11140
rect -1125 11100 -815 11140
rect -775 11100 -465 11140
rect -425 11100 -115 11140
rect -75 11100 235 11140
rect 275 11100 585 11140
rect 625 11100 935 11140
rect 975 11100 1285 11140
rect 1325 11100 1635 11140
rect 1675 11100 1680 11140
rect -1170 11095 1680 11100
rect 9630 11140 14580 11145
rect 9630 11100 9635 11140
rect 9675 11100 9985 11140
rect 10025 11100 10335 11140
rect 10375 11100 10685 11140
rect 10725 11100 11035 11140
rect 11075 11100 11385 11140
rect 11425 11100 11735 11140
rect 11775 11100 12085 11140
rect 12125 11100 12435 11140
rect 12475 11100 12785 11140
rect 12825 11100 13135 11140
rect 13175 11100 13485 11140
rect 13525 11100 13835 11140
rect 13875 11100 14185 11140
rect 14225 11100 14535 11140
rect 14575 11100 14580 11140
rect 9630 11095 14580 11100
rect 230 10795 280 11095
rect 12080 10795 12130 11095
rect -1170 10790 1680 10795
rect -1170 10750 -1165 10790
rect -1125 10750 -815 10790
rect -775 10750 -465 10790
rect -425 10750 -115 10790
rect -75 10750 235 10790
rect 275 10750 585 10790
rect 625 10750 935 10790
rect 975 10750 1285 10790
rect 1325 10750 1635 10790
rect 1675 10750 1680 10790
rect -1170 10745 1680 10750
rect 9630 10790 14580 10795
rect 9630 10750 9635 10790
rect 9675 10750 9985 10790
rect 10025 10750 10335 10790
rect 10375 10750 10685 10790
rect 10725 10750 11035 10790
rect 11075 10750 11385 10790
rect 11425 10750 11735 10790
rect 11775 10750 12085 10790
rect 12125 10750 12435 10790
rect 12475 10750 12785 10790
rect 12825 10750 13135 10790
rect 13175 10750 13485 10790
rect 13525 10750 13835 10790
rect 13875 10750 14185 10790
rect 14225 10750 14535 10790
rect 14575 10750 14580 10790
rect 9630 10745 14580 10750
rect 230 10445 280 10745
rect 12080 10445 12130 10745
rect -1170 10440 1680 10445
rect -1170 10400 -1165 10440
rect -1125 10400 -815 10440
rect -775 10400 -465 10440
rect -425 10400 -115 10440
rect -75 10400 235 10440
rect 275 10400 585 10440
rect 625 10400 935 10440
rect 975 10400 1285 10440
rect 1325 10400 1635 10440
rect 1675 10400 1680 10440
rect -1170 10395 1680 10400
rect 9630 10440 14580 10445
rect 9630 10400 9635 10440
rect 9675 10400 9985 10440
rect 10025 10400 10335 10440
rect 10375 10400 10685 10440
rect 10725 10400 11035 10440
rect 11075 10400 11385 10440
rect 11425 10400 11735 10440
rect 11775 10400 12085 10440
rect 12125 10400 12435 10440
rect 12475 10400 12785 10440
rect 12825 10400 13135 10440
rect 13175 10400 13485 10440
rect 13525 10400 13835 10440
rect 13875 10400 14185 10440
rect 14225 10400 14535 10440
rect 14575 10400 14580 10440
rect 9630 10395 14580 10400
rect 230 10095 280 10395
rect 12080 10095 12130 10395
rect -1170 10090 1680 10095
rect -1170 10050 -1165 10090
rect -1125 10050 -815 10090
rect -775 10050 -465 10090
rect -425 10050 -115 10090
rect -75 10050 235 10090
rect 275 10050 585 10090
rect 625 10050 935 10090
rect 975 10050 1285 10090
rect 1325 10050 1635 10090
rect 1675 10050 1680 10090
rect -1170 10045 1680 10050
rect 9630 10090 14580 10095
rect 9630 10050 9635 10090
rect 9675 10050 9985 10090
rect 10025 10050 10335 10090
rect 10375 10050 10685 10090
rect 10725 10050 11035 10090
rect 11075 10050 11385 10090
rect 11425 10050 11735 10090
rect 11775 10050 12085 10090
rect 12125 10050 12435 10090
rect 12475 10050 12785 10090
rect 12825 10050 13135 10090
rect 13175 10050 13485 10090
rect 13525 10050 13835 10090
rect 13875 10050 14185 10090
rect 14225 10050 14535 10090
rect 14575 10050 14580 10090
rect 9630 10045 14580 10050
rect 12080 9745 12130 10045
rect 9630 9740 14580 9745
rect 9630 9700 9635 9740
rect 9675 9700 9985 9740
rect 10025 9700 10335 9740
rect 10375 9700 10685 9740
rect 10725 9700 11035 9740
rect 11075 9700 11385 9740
rect 11425 9700 11735 9740
rect 11775 9700 12085 9740
rect 12125 9700 12435 9740
rect 12475 9700 12785 9740
rect 12825 9700 13135 9740
rect 13175 9700 13485 9740
rect 13525 9700 13835 9740
rect 13875 9700 14185 9740
rect 14225 9700 14535 9740
rect 14575 9700 14580 9740
rect 9630 9695 14580 9700
rect -4840 9640 9100 9650
rect -4840 9615 -80 9640
rect -4840 9565 -4805 9615
rect -4755 9565 -4710 9615
rect -4660 9565 -4615 9615
rect -4565 9565 -4515 9615
rect -4465 9565 -4415 9615
rect -4365 9565 -4315 9615
rect -4265 9565 -4220 9615
rect -4170 9565 -4125 9615
rect -4075 9565 -4005 9615
rect -3955 9565 -3910 9615
rect -3860 9565 -3815 9615
rect -3765 9565 -3715 9615
rect -3665 9565 -3615 9615
rect -3565 9565 -3515 9615
rect -3465 9565 -3420 9615
rect -3370 9565 -3325 9615
rect -3275 9565 -3205 9615
rect -3155 9565 -3110 9615
rect -3060 9565 -3015 9615
rect -2965 9565 -2915 9615
rect -2865 9565 -2815 9615
rect -2765 9565 -2715 9615
rect -2665 9565 -2620 9615
rect -2570 9565 -2525 9615
rect -2475 9565 -2405 9615
rect -2355 9565 -2310 9615
rect -2260 9565 -2215 9615
rect -2165 9565 -2115 9615
rect -2065 9565 -2015 9615
rect -1965 9565 -1915 9615
rect -1865 9565 -1820 9615
rect -1770 9565 -1725 9615
rect -1675 9600 -80 9615
rect -40 9600 270 9640
rect 310 9600 620 9640
rect 660 9600 1320 9640
rect 1360 9600 1670 9640
rect 1710 9600 2385 9640
rect 2425 9600 3235 9640
rect 3275 9600 5645 9640
rect 5685 9600 6300 9640
rect 6340 9600 6590 9640
rect 6630 9600 7270 9640
rect 7310 9600 7620 9640
rect 7660 9600 8320 9640
rect 8360 9600 8670 9640
rect 8710 9600 9020 9640
rect 9060 9600 9100 9640
rect -1675 9575 9100 9600
rect -1675 9565 -80 9575
rect -4840 9535 -80 9565
rect -40 9535 270 9575
rect 310 9535 620 9575
rect 660 9535 1320 9575
rect 1360 9535 1670 9575
rect 1710 9535 2385 9575
rect 2425 9535 3235 9575
rect 3275 9535 5645 9575
rect 5685 9535 6300 9575
rect 6340 9535 6590 9575
rect 6630 9535 7270 9575
rect 7310 9535 7620 9575
rect 7660 9535 8320 9575
rect 8360 9535 8670 9575
rect 8710 9535 9020 9575
rect 9060 9535 9100 9575
rect -4840 9525 9100 9535
rect -4840 9475 -4805 9525
rect -4755 9475 -4710 9525
rect -4660 9475 -4615 9525
rect -4565 9475 -4515 9525
rect -4465 9475 -4415 9525
rect -4365 9475 -4315 9525
rect -4265 9475 -4220 9525
rect -4170 9475 -4125 9525
rect -4075 9475 -4005 9525
rect -3955 9475 -3910 9525
rect -3860 9475 -3815 9525
rect -3765 9475 -3715 9525
rect -3665 9475 -3615 9525
rect -3565 9475 -3515 9525
rect -3465 9475 -3420 9525
rect -3370 9475 -3325 9525
rect -3275 9475 -3205 9525
rect -3155 9475 -3110 9525
rect -3060 9475 -3015 9525
rect -2965 9475 -2915 9525
rect -2865 9475 -2815 9525
rect -2765 9475 -2715 9525
rect -2665 9475 -2620 9525
rect -2570 9475 -2525 9525
rect -2475 9475 -2405 9525
rect -2355 9475 -2310 9525
rect -2260 9475 -2215 9525
rect -2165 9475 -2115 9525
rect -2065 9475 -2015 9525
rect -1965 9475 -1915 9525
rect -1865 9475 -1820 9525
rect -1770 9475 -1725 9525
rect -1675 9505 9100 9525
rect -1675 9475 -80 9505
rect -4840 9465 -80 9475
rect -40 9465 270 9505
rect 310 9465 620 9505
rect 660 9465 1320 9505
rect 1360 9465 1670 9505
rect 1710 9465 2385 9505
rect 2425 9465 3235 9505
rect 3275 9465 5645 9505
rect 5685 9465 6300 9505
rect 6340 9465 6590 9505
rect 6630 9465 7270 9505
rect 7310 9465 7620 9505
rect 7660 9465 8320 9505
rect 8360 9465 8670 9505
rect 8710 9465 9020 9505
rect 9060 9465 9100 9505
rect -4840 9435 9100 9465
rect -4840 9425 -80 9435
rect -4840 9375 -4805 9425
rect -4755 9375 -4710 9425
rect -4660 9375 -4615 9425
rect -4565 9375 -4515 9425
rect -4465 9375 -4415 9425
rect -4365 9375 -4315 9425
rect -4265 9375 -4220 9425
rect -4170 9375 -4125 9425
rect -4075 9375 -4005 9425
rect -3955 9375 -3910 9425
rect -3860 9375 -3815 9425
rect -3765 9375 -3715 9425
rect -3665 9375 -3615 9425
rect -3565 9375 -3515 9425
rect -3465 9375 -3420 9425
rect -3370 9375 -3325 9425
rect -3275 9375 -3205 9425
rect -3155 9375 -3110 9425
rect -3060 9375 -3015 9425
rect -2965 9375 -2915 9425
rect -2865 9375 -2815 9425
rect -2765 9375 -2715 9425
rect -2665 9375 -2620 9425
rect -2570 9375 -2525 9425
rect -2475 9375 -2405 9425
rect -2355 9375 -2310 9425
rect -2260 9375 -2215 9425
rect -2165 9375 -2115 9425
rect -2065 9375 -2015 9425
rect -1965 9375 -1915 9425
rect -1865 9375 -1820 9425
rect -1770 9375 -1725 9425
rect -1675 9395 -80 9425
rect -40 9395 270 9435
rect 310 9395 620 9435
rect 660 9395 1320 9435
rect 1360 9395 1670 9435
rect 1710 9395 2385 9435
rect 2425 9395 3235 9435
rect 3275 9395 5645 9435
rect 5685 9395 6300 9435
rect 6340 9395 6590 9435
rect 6630 9395 7270 9435
rect 7310 9395 7620 9435
rect 7660 9395 8320 9435
rect 8360 9395 8670 9435
rect 8710 9395 9020 9435
rect 9060 9395 9100 9435
rect 12080 9395 12130 9695
rect 14790 9615 20720 9650
rect 14790 9565 14825 9615
rect 14875 9565 14920 9615
rect 14970 9565 15015 9615
rect 15065 9565 15115 9615
rect 15165 9565 15215 9615
rect 15265 9565 15315 9615
rect 15365 9565 15410 9615
rect 15460 9565 15505 9615
rect 15555 9565 15625 9615
rect 15675 9565 15720 9615
rect 15770 9565 15815 9615
rect 15865 9565 15915 9615
rect 15965 9565 16015 9615
rect 16065 9565 16115 9615
rect 16165 9565 16210 9615
rect 16260 9565 16305 9615
rect 16355 9565 16425 9615
rect 16475 9565 16520 9615
rect 16570 9565 16615 9615
rect 16665 9565 16715 9615
rect 16765 9565 16815 9615
rect 16865 9565 16915 9615
rect 16965 9565 17010 9615
rect 17060 9565 17105 9615
rect 17155 9565 17225 9615
rect 17275 9565 17320 9615
rect 17370 9565 17415 9615
rect 17465 9565 17515 9615
rect 17565 9565 17615 9615
rect 17665 9565 17715 9615
rect 17765 9565 17810 9615
rect 17860 9565 17905 9615
rect 17955 9565 20720 9615
rect 14790 9525 20720 9565
rect 14790 9475 14825 9525
rect 14875 9475 14920 9525
rect 14970 9475 15015 9525
rect 15065 9475 15115 9525
rect 15165 9475 15215 9525
rect 15265 9475 15315 9525
rect 15365 9475 15410 9525
rect 15460 9475 15505 9525
rect 15555 9475 15625 9525
rect 15675 9475 15720 9525
rect 15770 9475 15815 9525
rect 15865 9475 15915 9525
rect 15965 9475 16015 9525
rect 16065 9475 16115 9525
rect 16165 9475 16210 9525
rect 16260 9475 16305 9525
rect 16355 9475 16425 9525
rect 16475 9475 16520 9525
rect 16570 9475 16615 9525
rect 16665 9475 16715 9525
rect 16765 9475 16815 9525
rect 16865 9475 16915 9525
rect 16965 9475 17010 9525
rect 17060 9475 17105 9525
rect 17155 9475 17225 9525
rect 17275 9475 17320 9525
rect 17370 9475 17415 9525
rect 17465 9475 17515 9525
rect 17565 9475 17615 9525
rect 17665 9475 17715 9525
rect 17765 9475 17810 9525
rect 17860 9475 17905 9525
rect 17955 9475 20720 9525
rect 14790 9425 20720 9475
rect -1675 9375 9100 9395
rect -4840 9365 9100 9375
rect -4840 9335 -80 9365
rect -4840 9285 -4805 9335
rect -4755 9285 -4710 9335
rect -4660 9285 -4615 9335
rect -4565 9285 -4515 9335
rect -4465 9285 -4415 9335
rect -4365 9285 -4315 9335
rect -4265 9285 -4220 9335
rect -4170 9285 -4125 9335
rect -4075 9285 -4005 9335
rect -3955 9285 -3910 9335
rect -3860 9285 -3815 9335
rect -3765 9285 -3715 9335
rect -3665 9285 -3615 9335
rect -3565 9285 -3515 9335
rect -3465 9285 -3420 9335
rect -3370 9285 -3325 9335
rect -3275 9285 -3205 9335
rect -3155 9285 -3110 9335
rect -3060 9285 -3015 9335
rect -2965 9285 -2915 9335
rect -2865 9285 -2815 9335
rect -2765 9285 -2715 9335
rect -2665 9285 -2620 9335
rect -2570 9285 -2525 9335
rect -2475 9285 -2405 9335
rect -2355 9285 -2310 9335
rect -2260 9285 -2215 9335
rect -2165 9285 -2115 9335
rect -2065 9285 -2015 9335
rect -1965 9285 -1915 9335
rect -1865 9285 -1820 9335
rect -1770 9285 -1725 9335
rect -1675 9325 -80 9335
rect -40 9325 270 9365
rect 310 9325 620 9365
rect 660 9325 1320 9365
rect 1360 9325 1670 9365
rect 1710 9325 2385 9365
rect 2425 9325 3235 9365
rect 3275 9325 5645 9365
rect 5685 9325 6300 9365
rect 6340 9325 6590 9365
rect 6630 9325 7270 9365
rect 7310 9325 7620 9365
rect 7660 9325 8320 9365
rect 8360 9325 8670 9365
rect 8710 9325 9020 9365
rect 9060 9325 9100 9365
rect 9630 9390 14580 9395
rect 9630 9350 9635 9390
rect 9675 9350 9985 9390
rect 10025 9350 10335 9390
rect 10375 9350 10685 9390
rect 10725 9350 11035 9390
rect 11075 9350 11385 9390
rect 11425 9350 11735 9390
rect 11775 9350 12085 9390
rect 12125 9350 12435 9390
rect 12475 9350 12785 9390
rect 12825 9350 13135 9390
rect 13175 9350 13485 9390
rect 13525 9350 13835 9390
rect 13875 9350 14185 9390
rect 14225 9350 14535 9390
rect 14575 9350 14580 9390
rect 9630 9345 14580 9350
rect 14790 9375 14825 9425
rect 14875 9375 14920 9425
rect 14970 9375 15015 9425
rect 15065 9375 15115 9425
rect 15165 9375 15215 9425
rect 15265 9375 15315 9425
rect 15365 9375 15410 9425
rect 15460 9375 15505 9425
rect 15555 9375 15625 9425
rect 15675 9375 15720 9425
rect 15770 9375 15815 9425
rect 15865 9375 15915 9425
rect 15965 9375 16015 9425
rect 16065 9375 16115 9425
rect 16165 9375 16210 9425
rect 16260 9375 16305 9425
rect 16355 9375 16425 9425
rect 16475 9375 16520 9425
rect 16570 9375 16615 9425
rect 16665 9375 16715 9425
rect 16765 9375 16815 9425
rect 16865 9375 16915 9425
rect 16965 9375 17010 9425
rect 17060 9375 17105 9425
rect 17155 9375 17225 9425
rect 17275 9375 17320 9425
rect 17370 9375 17415 9425
rect 17465 9375 17515 9425
rect 17565 9375 17615 9425
rect 17665 9375 17715 9425
rect 17765 9375 17810 9425
rect 17860 9375 17905 9425
rect 17955 9375 20720 9425
rect -1675 9300 9100 9325
rect -1675 9285 -80 9300
rect -4840 9260 -80 9285
rect -40 9260 270 9300
rect 310 9260 620 9300
rect 660 9260 1320 9300
rect 1360 9260 1670 9300
rect 1710 9260 2385 9300
rect 2425 9260 3235 9300
rect 3275 9260 5645 9300
rect 5685 9260 6300 9300
rect 6340 9260 6590 9300
rect 6630 9260 7270 9300
rect 7310 9260 7620 9300
rect 7660 9260 8320 9300
rect 8360 9260 8670 9300
rect 8710 9260 9020 9300
rect 9060 9260 9100 9300
rect -4840 9240 9100 9260
rect -4840 9215 -80 9240
rect -4840 9165 -4805 9215
rect -4755 9165 -4710 9215
rect -4660 9165 -4615 9215
rect -4565 9165 -4515 9215
rect -4465 9165 -4415 9215
rect -4365 9165 -4315 9215
rect -4265 9165 -4220 9215
rect -4170 9165 -4125 9215
rect -4075 9165 -4005 9215
rect -3955 9165 -3910 9215
rect -3860 9165 -3815 9215
rect -3765 9165 -3715 9215
rect -3665 9165 -3615 9215
rect -3565 9165 -3515 9215
rect -3465 9165 -3420 9215
rect -3370 9165 -3325 9215
rect -3275 9165 -3205 9215
rect -3155 9165 -3110 9215
rect -3060 9165 -3015 9215
rect -2965 9165 -2915 9215
rect -2865 9165 -2815 9215
rect -2765 9165 -2715 9215
rect -2665 9165 -2620 9215
rect -2570 9165 -2525 9215
rect -2475 9165 -2405 9215
rect -2355 9165 -2310 9215
rect -2260 9165 -2215 9215
rect -2165 9165 -2115 9215
rect -2065 9165 -2015 9215
rect -1965 9165 -1915 9215
rect -1865 9165 -1820 9215
rect -1770 9165 -1725 9215
rect -1675 9200 -80 9215
rect -40 9200 270 9240
rect 310 9200 620 9240
rect 660 9200 1320 9240
rect 1360 9200 1670 9240
rect 1710 9200 2385 9240
rect 2425 9200 3235 9240
rect 3275 9200 5645 9240
rect 5685 9200 6300 9240
rect 6340 9200 6590 9240
rect 6630 9200 7270 9240
rect 7310 9200 7620 9240
rect 7660 9200 8320 9240
rect 8360 9200 8670 9240
rect 8710 9200 9020 9240
rect 9060 9200 9100 9240
rect -1675 9175 9100 9200
rect -1675 9165 -80 9175
rect -4840 9135 -80 9165
rect -40 9135 270 9175
rect 310 9135 620 9175
rect 660 9135 1320 9175
rect 1360 9135 1670 9175
rect 1710 9135 2385 9175
rect 2425 9135 3235 9175
rect 3275 9135 5645 9175
rect 5685 9135 6300 9175
rect 6340 9135 6590 9175
rect 6630 9135 7270 9175
rect 7310 9135 7620 9175
rect 7660 9135 8320 9175
rect 8360 9135 8670 9175
rect 8710 9135 9020 9175
rect 9060 9135 9100 9175
rect -4840 9125 9100 9135
rect -4840 9075 -4805 9125
rect -4755 9075 -4710 9125
rect -4660 9075 -4615 9125
rect -4565 9075 -4515 9125
rect -4465 9075 -4415 9125
rect -4365 9075 -4315 9125
rect -4265 9075 -4220 9125
rect -4170 9075 -4125 9125
rect -4075 9075 -4005 9125
rect -3955 9075 -3910 9125
rect -3860 9075 -3815 9125
rect -3765 9075 -3715 9125
rect -3665 9075 -3615 9125
rect -3565 9075 -3515 9125
rect -3465 9075 -3420 9125
rect -3370 9075 -3325 9125
rect -3275 9075 -3205 9125
rect -3155 9075 -3110 9125
rect -3060 9075 -3015 9125
rect -2965 9075 -2915 9125
rect -2865 9075 -2815 9125
rect -2765 9075 -2715 9125
rect -2665 9075 -2620 9125
rect -2570 9075 -2525 9125
rect -2475 9075 -2405 9125
rect -2355 9075 -2310 9125
rect -2260 9075 -2215 9125
rect -2165 9075 -2115 9125
rect -2065 9075 -2015 9125
rect -1965 9075 -1915 9125
rect -1865 9075 -1820 9125
rect -1770 9075 -1725 9125
rect -1675 9105 9100 9125
rect -1675 9075 -80 9105
rect -4840 9065 -80 9075
rect -40 9065 270 9105
rect 310 9065 620 9105
rect 660 9065 1320 9105
rect 1360 9065 1670 9105
rect 1710 9065 2385 9105
rect 2425 9065 3235 9105
rect 3275 9065 5645 9105
rect 5685 9065 6300 9105
rect 6340 9065 6590 9105
rect 6630 9065 7270 9105
rect 7310 9065 7620 9105
rect 7660 9065 8320 9105
rect 8360 9065 8670 9105
rect 8710 9065 9020 9105
rect 9060 9065 9100 9105
rect -4840 9035 9100 9065
rect 12080 9045 12130 9345
rect 14790 9335 20720 9375
rect 14790 9285 14825 9335
rect 14875 9285 14920 9335
rect 14970 9285 15015 9335
rect 15065 9285 15115 9335
rect 15165 9285 15215 9335
rect 15265 9285 15315 9335
rect 15365 9285 15410 9335
rect 15460 9285 15505 9335
rect 15555 9285 15625 9335
rect 15675 9285 15720 9335
rect 15770 9285 15815 9335
rect 15865 9285 15915 9335
rect 15965 9285 16015 9335
rect 16065 9285 16115 9335
rect 16165 9285 16210 9335
rect 16260 9285 16305 9335
rect 16355 9285 16425 9335
rect 16475 9285 16520 9335
rect 16570 9285 16615 9335
rect 16665 9285 16715 9335
rect 16765 9285 16815 9335
rect 16865 9285 16915 9335
rect 16965 9285 17010 9335
rect 17060 9285 17105 9335
rect 17155 9285 17225 9335
rect 17275 9285 17320 9335
rect 17370 9285 17415 9335
rect 17465 9285 17515 9335
rect 17565 9285 17615 9335
rect 17665 9285 17715 9335
rect 17765 9285 17810 9335
rect 17860 9285 17905 9335
rect 17955 9285 20720 9335
rect 14790 9215 20720 9285
rect 14790 9165 14825 9215
rect 14875 9165 14920 9215
rect 14970 9165 15015 9215
rect 15065 9165 15115 9215
rect 15165 9165 15215 9215
rect 15265 9165 15315 9215
rect 15365 9165 15410 9215
rect 15460 9165 15505 9215
rect 15555 9165 15625 9215
rect 15675 9165 15720 9215
rect 15770 9165 15815 9215
rect 15865 9165 15915 9215
rect 15965 9165 16015 9215
rect 16065 9165 16115 9215
rect 16165 9165 16210 9215
rect 16260 9165 16305 9215
rect 16355 9165 16425 9215
rect 16475 9165 16520 9215
rect 16570 9165 16615 9215
rect 16665 9165 16715 9215
rect 16765 9165 16815 9215
rect 16865 9165 16915 9215
rect 16965 9165 17010 9215
rect 17060 9165 17105 9215
rect 17155 9165 17225 9215
rect 17275 9165 17320 9215
rect 17370 9165 17415 9215
rect 17465 9165 17515 9215
rect 17565 9165 17615 9215
rect 17665 9165 17715 9215
rect 17765 9165 17810 9215
rect 17860 9165 17905 9215
rect 17955 9165 20720 9215
rect 14790 9125 20720 9165
rect 14790 9075 14825 9125
rect 14875 9075 14920 9125
rect 14970 9075 15015 9125
rect 15065 9075 15115 9125
rect 15165 9075 15215 9125
rect 15265 9075 15315 9125
rect 15365 9075 15410 9125
rect 15460 9075 15505 9125
rect 15555 9075 15625 9125
rect 15675 9075 15720 9125
rect 15770 9075 15815 9125
rect 15865 9075 15915 9125
rect 15965 9075 16015 9125
rect 16065 9075 16115 9125
rect 16165 9075 16210 9125
rect 16260 9075 16305 9125
rect 16355 9075 16425 9125
rect 16475 9075 16520 9125
rect 16570 9075 16615 9125
rect 16665 9075 16715 9125
rect 16765 9075 16815 9125
rect 16865 9075 16915 9125
rect 16965 9075 17010 9125
rect 17060 9075 17105 9125
rect 17155 9075 17225 9125
rect 17275 9075 17320 9125
rect 17370 9075 17415 9125
rect 17465 9075 17515 9125
rect 17565 9075 17615 9125
rect 17665 9075 17715 9125
rect 17765 9075 17810 9125
rect 17860 9075 17905 9125
rect 17955 9075 20720 9125
rect -4840 9025 -80 9035
rect -4840 8975 -4805 9025
rect -4755 8975 -4710 9025
rect -4660 8975 -4615 9025
rect -4565 8975 -4515 9025
rect -4465 8975 -4415 9025
rect -4365 8975 -4315 9025
rect -4265 8975 -4220 9025
rect -4170 8975 -4125 9025
rect -4075 8975 -4005 9025
rect -3955 8975 -3910 9025
rect -3860 8975 -3815 9025
rect -3765 8975 -3715 9025
rect -3665 8975 -3615 9025
rect -3565 8975 -3515 9025
rect -3465 8975 -3420 9025
rect -3370 8975 -3325 9025
rect -3275 8975 -3205 9025
rect -3155 8975 -3110 9025
rect -3060 8975 -3015 9025
rect -2965 8975 -2915 9025
rect -2865 8975 -2815 9025
rect -2765 8975 -2715 9025
rect -2665 8975 -2620 9025
rect -2570 8975 -2525 9025
rect -2475 8975 -2405 9025
rect -2355 8975 -2310 9025
rect -2260 8975 -2215 9025
rect -2165 8975 -2115 9025
rect -2065 8975 -2015 9025
rect -1965 8975 -1915 9025
rect -1865 8975 -1820 9025
rect -1770 8975 -1725 9025
rect -1675 8995 -80 9025
rect -40 8995 270 9035
rect 310 8995 620 9035
rect 660 8995 1320 9035
rect 1360 8995 1670 9035
rect 1710 8995 2385 9035
rect 2425 8995 3235 9035
rect 3275 8995 5645 9035
rect 5685 8995 6300 9035
rect 6340 8995 6590 9035
rect 6630 8995 7270 9035
rect 7310 8995 7620 9035
rect 7660 8995 8320 9035
rect 8360 8995 8670 9035
rect 8710 8995 9020 9035
rect 9060 8995 9100 9035
rect 9630 9040 14580 9045
rect 9630 9000 9635 9040
rect 9675 9000 9985 9040
rect 10025 9000 10335 9040
rect 10375 9000 10685 9040
rect 10725 9000 11035 9040
rect 11075 9000 11385 9040
rect 11425 9000 11735 9040
rect 11775 9000 12085 9040
rect 12125 9000 12435 9040
rect 12475 9000 12785 9040
rect 12825 9000 13135 9040
rect 13175 9000 13485 9040
rect 13525 9000 13835 9040
rect 13875 9000 14185 9040
rect 14225 9000 14535 9040
rect 14575 9000 14580 9040
rect 9630 8995 14580 9000
rect 14790 9025 20720 9075
rect -1675 8975 9100 8995
rect -4840 8965 9100 8975
rect -4840 8935 -80 8965
rect -4840 8885 -4805 8935
rect -4755 8885 -4710 8935
rect -4660 8885 -4615 8935
rect -4565 8885 -4515 8935
rect -4465 8885 -4415 8935
rect -4365 8885 -4315 8935
rect -4265 8885 -4220 8935
rect -4170 8885 -4125 8935
rect -4075 8885 -4005 8935
rect -3955 8885 -3910 8935
rect -3860 8885 -3815 8935
rect -3765 8885 -3715 8935
rect -3665 8885 -3615 8935
rect -3565 8885 -3515 8935
rect -3465 8885 -3420 8935
rect -3370 8885 -3325 8935
rect -3275 8885 -3205 8935
rect -3155 8885 -3110 8935
rect -3060 8885 -3015 8935
rect -2965 8885 -2915 8935
rect -2865 8885 -2815 8935
rect -2765 8885 -2715 8935
rect -2665 8885 -2620 8935
rect -2570 8885 -2525 8935
rect -2475 8885 -2405 8935
rect -2355 8885 -2310 8935
rect -2260 8885 -2215 8935
rect -2165 8885 -2115 8935
rect -2065 8885 -2015 8935
rect -1965 8885 -1915 8935
rect -1865 8885 -1820 8935
rect -1770 8885 -1725 8935
rect -1675 8925 -80 8935
rect -40 8925 270 8965
rect 310 8925 620 8965
rect 660 8925 1320 8965
rect 1360 8925 1670 8965
rect 1710 8925 2385 8965
rect 2425 8925 3235 8965
rect 3275 8925 5645 8965
rect 5685 8925 6300 8965
rect 6340 8925 6590 8965
rect 6630 8925 7270 8965
rect 7310 8925 7620 8965
rect 7660 8925 8320 8965
rect 8360 8925 8670 8965
rect 8710 8925 9020 8965
rect 9060 8925 9100 8965
rect -1675 8900 9100 8925
rect -1675 8885 -80 8900
rect -4840 8860 -80 8885
rect -40 8860 270 8900
rect 310 8860 620 8900
rect 660 8860 1320 8900
rect 1360 8860 1670 8900
rect 1710 8860 2385 8900
rect 2425 8860 3235 8900
rect 3275 8860 5645 8900
rect 5685 8860 6300 8900
rect 6340 8860 6590 8900
rect 6630 8860 7270 8900
rect 7310 8860 7620 8900
rect 7660 8860 8320 8900
rect 8360 8860 8670 8900
rect 8710 8860 9020 8900
rect 9060 8860 9100 8900
rect -4840 8840 9100 8860
rect -4840 8815 -80 8840
rect -4840 8765 -4805 8815
rect -4755 8765 -4710 8815
rect -4660 8765 -4615 8815
rect -4565 8765 -4515 8815
rect -4465 8765 -4415 8815
rect -4365 8765 -4315 8815
rect -4265 8765 -4220 8815
rect -4170 8765 -4125 8815
rect -4075 8765 -4005 8815
rect -3955 8765 -3910 8815
rect -3860 8765 -3815 8815
rect -3765 8765 -3715 8815
rect -3665 8765 -3615 8815
rect -3565 8765 -3515 8815
rect -3465 8765 -3420 8815
rect -3370 8765 -3325 8815
rect -3275 8765 -3205 8815
rect -3155 8765 -3110 8815
rect -3060 8765 -3015 8815
rect -2965 8765 -2915 8815
rect -2865 8765 -2815 8815
rect -2765 8765 -2715 8815
rect -2665 8765 -2620 8815
rect -2570 8765 -2525 8815
rect -2475 8765 -2405 8815
rect -2355 8765 -2310 8815
rect -2260 8765 -2215 8815
rect -2165 8765 -2115 8815
rect -2065 8765 -2015 8815
rect -1965 8765 -1915 8815
rect -1865 8765 -1820 8815
rect -1770 8765 -1725 8815
rect -1675 8800 -80 8815
rect -40 8800 270 8840
rect 310 8800 620 8840
rect 660 8800 1320 8840
rect 1360 8800 1670 8840
rect 1710 8800 2385 8840
rect 2425 8800 3235 8840
rect 3275 8800 5645 8840
rect 5685 8800 6300 8840
rect 6340 8800 6590 8840
rect 6630 8800 7270 8840
rect 7310 8800 7620 8840
rect 7660 8800 8320 8840
rect 8360 8800 8670 8840
rect 8710 8800 9020 8840
rect 9060 8800 9100 8840
rect -1675 8775 9100 8800
rect -1675 8765 -80 8775
rect -4840 8735 -80 8765
rect -40 8735 270 8775
rect 310 8735 620 8775
rect 660 8735 1320 8775
rect 1360 8735 1670 8775
rect 1710 8735 2385 8775
rect 2425 8735 3235 8775
rect 3275 8735 5645 8775
rect 5685 8735 6300 8775
rect 6340 8735 6590 8775
rect 6630 8735 7270 8775
rect 7310 8735 7620 8775
rect 7660 8735 8320 8775
rect 8360 8735 8670 8775
rect 8710 8735 9020 8775
rect 9060 8735 9100 8775
rect -4840 8725 9100 8735
rect -4840 8675 -4805 8725
rect -4755 8675 -4710 8725
rect -4660 8675 -4615 8725
rect -4565 8675 -4515 8725
rect -4465 8675 -4415 8725
rect -4365 8675 -4315 8725
rect -4265 8675 -4220 8725
rect -4170 8675 -4125 8725
rect -4075 8675 -4005 8725
rect -3955 8675 -3910 8725
rect -3860 8675 -3815 8725
rect -3765 8675 -3715 8725
rect -3665 8675 -3615 8725
rect -3565 8675 -3515 8725
rect -3465 8675 -3420 8725
rect -3370 8675 -3325 8725
rect -3275 8675 -3205 8725
rect -3155 8675 -3110 8725
rect -3060 8675 -3015 8725
rect -2965 8675 -2915 8725
rect -2865 8675 -2815 8725
rect -2765 8675 -2715 8725
rect -2665 8675 -2620 8725
rect -2570 8675 -2525 8725
rect -2475 8675 -2405 8725
rect -2355 8675 -2310 8725
rect -2260 8675 -2215 8725
rect -2165 8675 -2115 8725
rect -2065 8675 -2015 8725
rect -1965 8675 -1915 8725
rect -1865 8675 -1820 8725
rect -1770 8675 -1725 8725
rect -1675 8705 9100 8725
rect -1675 8675 -80 8705
rect -4840 8665 -80 8675
rect -40 8665 270 8705
rect 310 8665 620 8705
rect 660 8665 1320 8705
rect 1360 8665 1670 8705
rect 1710 8665 2385 8705
rect 2425 8665 3235 8705
rect 3275 8665 5645 8705
rect 5685 8665 6300 8705
rect 6340 8665 6590 8705
rect 6630 8665 7270 8705
rect 7310 8665 7620 8705
rect 7660 8665 8320 8705
rect 8360 8665 8670 8705
rect 8710 8665 9020 8705
rect 9060 8665 9100 8705
rect 12080 8695 12130 8995
rect 14790 8975 14825 9025
rect 14875 8975 14920 9025
rect 14970 8975 15015 9025
rect 15065 8975 15115 9025
rect 15165 8975 15215 9025
rect 15265 8975 15315 9025
rect 15365 8975 15410 9025
rect 15460 8975 15505 9025
rect 15555 8975 15625 9025
rect 15675 8975 15720 9025
rect 15770 8975 15815 9025
rect 15865 8975 15915 9025
rect 15965 8975 16015 9025
rect 16065 8975 16115 9025
rect 16165 8975 16210 9025
rect 16260 8975 16305 9025
rect 16355 8975 16425 9025
rect 16475 8975 16520 9025
rect 16570 8975 16615 9025
rect 16665 8975 16715 9025
rect 16765 8975 16815 9025
rect 16865 8975 16915 9025
rect 16965 8975 17010 9025
rect 17060 8975 17105 9025
rect 17155 8975 17225 9025
rect 17275 8975 17320 9025
rect 17370 8975 17415 9025
rect 17465 8975 17515 9025
rect 17565 8975 17615 9025
rect 17665 8975 17715 9025
rect 17765 8975 17810 9025
rect 17860 8975 17905 9025
rect 17955 8975 20720 9025
rect 14790 8935 20720 8975
rect 14790 8885 14825 8935
rect 14875 8885 14920 8935
rect 14970 8885 15015 8935
rect 15065 8885 15115 8935
rect 15165 8885 15215 8935
rect 15265 8885 15315 8935
rect 15365 8885 15410 8935
rect 15460 8885 15505 8935
rect 15555 8885 15625 8935
rect 15675 8885 15720 8935
rect 15770 8885 15815 8935
rect 15865 8885 15915 8935
rect 15965 8885 16015 8935
rect 16065 8885 16115 8935
rect 16165 8885 16210 8935
rect 16260 8885 16305 8935
rect 16355 8885 16425 8935
rect 16475 8885 16520 8935
rect 16570 8885 16615 8935
rect 16665 8885 16715 8935
rect 16765 8885 16815 8935
rect 16865 8885 16915 8935
rect 16965 8885 17010 8935
rect 17060 8885 17105 8935
rect 17155 8885 17225 8935
rect 17275 8885 17320 8935
rect 17370 8885 17415 8935
rect 17465 8885 17515 8935
rect 17565 8885 17615 8935
rect 17665 8885 17715 8935
rect 17765 8885 17810 8935
rect 17860 8885 17905 8935
rect 17955 8885 20720 8935
rect 14790 8815 20720 8885
rect 14790 8765 14825 8815
rect 14875 8765 14920 8815
rect 14970 8765 15015 8815
rect 15065 8765 15115 8815
rect 15165 8765 15215 8815
rect 15265 8765 15315 8815
rect 15365 8765 15410 8815
rect 15460 8765 15505 8815
rect 15555 8765 15625 8815
rect 15675 8765 15720 8815
rect 15770 8765 15815 8815
rect 15865 8765 15915 8815
rect 15965 8765 16015 8815
rect 16065 8765 16115 8815
rect 16165 8765 16210 8815
rect 16260 8765 16305 8815
rect 16355 8765 16425 8815
rect 16475 8765 16520 8815
rect 16570 8765 16615 8815
rect 16665 8765 16715 8815
rect 16765 8765 16815 8815
rect 16865 8765 16915 8815
rect 16965 8765 17010 8815
rect 17060 8765 17105 8815
rect 17155 8765 17225 8815
rect 17275 8765 17320 8815
rect 17370 8765 17415 8815
rect 17465 8765 17515 8815
rect 17565 8765 17615 8815
rect 17665 8765 17715 8815
rect 17765 8765 17810 8815
rect 17860 8765 17905 8815
rect 17955 8765 20720 8815
rect 14790 8725 20720 8765
rect -4840 8635 9100 8665
rect 9630 8690 14580 8695
rect 9630 8650 9635 8690
rect 9675 8650 9985 8690
rect 10025 8650 10335 8690
rect 10375 8650 10685 8690
rect 10725 8650 11035 8690
rect 11075 8650 11385 8690
rect 11425 8650 11735 8690
rect 11775 8650 12085 8690
rect 12125 8650 12435 8690
rect 12475 8650 12785 8690
rect 12825 8650 13135 8690
rect 13175 8650 13485 8690
rect 13525 8650 13835 8690
rect 13875 8650 14185 8690
rect 14225 8650 14535 8690
rect 14575 8650 14580 8690
rect 9630 8645 14580 8650
rect 14790 8675 14825 8725
rect 14875 8675 14920 8725
rect 14970 8675 15015 8725
rect 15065 8675 15115 8725
rect 15165 8675 15215 8725
rect 15265 8675 15315 8725
rect 15365 8675 15410 8725
rect 15460 8675 15505 8725
rect 15555 8675 15625 8725
rect 15675 8675 15720 8725
rect 15770 8675 15815 8725
rect 15865 8675 15915 8725
rect 15965 8675 16015 8725
rect 16065 8675 16115 8725
rect 16165 8675 16210 8725
rect 16260 8675 16305 8725
rect 16355 8675 16425 8725
rect 16475 8675 16520 8725
rect 16570 8675 16615 8725
rect 16665 8675 16715 8725
rect 16765 8675 16815 8725
rect 16865 8675 16915 8725
rect 16965 8675 17010 8725
rect 17060 8675 17105 8725
rect 17155 8675 17225 8725
rect 17275 8675 17320 8725
rect 17370 8675 17415 8725
rect 17465 8675 17515 8725
rect 17565 8675 17615 8725
rect 17665 8675 17715 8725
rect 17765 8675 17810 8725
rect 17860 8675 17905 8725
rect 17955 8675 20720 8725
rect -4840 8625 -80 8635
rect -4840 8575 -4805 8625
rect -4755 8575 -4710 8625
rect -4660 8575 -4615 8625
rect -4565 8575 -4515 8625
rect -4465 8575 -4415 8625
rect -4365 8575 -4315 8625
rect -4265 8575 -4220 8625
rect -4170 8575 -4125 8625
rect -4075 8575 -4005 8625
rect -3955 8575 -3910 8625
rect -3860 8575 -3815 8625
rect -3765 8575 -3715 8625
rect -3665 8575 -3615 8625
rect -3565 8575 -3515 8625
rect -3465 8575 -3420 8625
rect -3370 8575 -3325 8625
rect -3275 8575 -3205 8625
rect -3155 8575 -3110 8625
rect -3060 8575 -3015 8625
rect -2965 8575 -2915 8625
rect -2865 8575 -2815 8625
rect -2765 8575 -2715 8625
rect -2665 8575 -2620 8625
rect -2570 8575 -2525 8625
rect -2475 8575 -2405 8625
rect -2355 8575 -2310 8625
rect -2260 8575 -2215 8625
rect -2165 8575 -2115 8625
rect -2065 8575 -2015 8625
rect -1965 8575 -1915 8625
rect -1865 8575 -1820 8625
rect -1770 8575 -1725 8625
rect -1675 8595 -80 8625
rect -40 8595 270 8635
rect 310 8595 620 8635
rect 660 8595 1320 8635
rect 1360 8595 1670 8635
rect 1710 8595 2385 8635
rect 2425 8595 3235 8635
rect 3275 8595 5645 8635
rect 5685 8595 6300 8635
rect 6340 8595 6590 8635
rect 6630 8595 7270 8635
rect 7310 8595 7620 8635
rect 7660 8595 8320 8635
rect 8360 8595 8670 8635
rect 8710 8595 9020 8635
rect 9060 8595 9100 8635
rect -1675 8575 9100 8595
rect -4840 8565 9100 8575
rect -4840 8535 -80 8565
rect -4840 8485 -4805 8535
rect -4755 8485 -4710 8535
rect -4660 8485 -4615 8535
rect -4565 8485 -4515 8535
rect -4465 8485 -4415 8535
rect -4365 8485 -4315 8535
rect -4265 8485 -4220 8535
rect -4170 8485 -4125 8535
rect -4075 8485 -4005 8535
rect -3955 8485 -3910 8535
rect -3860 8485 -3815 8535
rect -3765 8485 -3715 8535
rect -3665 8485 -3615 8535
rect -3565 8485 -3515 8535
rect -3465 8485 -3420 8535
rect -3370 8485 -3325 8535
rect -3275 8485 -3205 8535
rect -3155 8485 -3110 8535
rect -3060 8485 -3015 8535
rect -2965 8485 -2915 8535
rect -2865 8485 -2815 8535
rect -2765 8485 -2715 8535
rect -2665 8485 -2620 8535
rect -2570 8485 -2525 8535
rect -2475 8485 -2405 8535
rect -2355 8485 -2310 8535
rect -2260 8485 -2215 8535
rect -2165 8485 -2115 8535
rect -2065 8485 -2015 8535
rect -1965 8485 -1915 8535
rect -1865 8485 -1820 8535
rect -1770 8485 -1725 8535
rect -1675 8525 -80 8535
rect -40 8525 270 8565
rect 310 8525 620 8565
rect 660 8525 1320 8565
rect 1360 8525 1670 8565
rect 1710 8525 2385 8565
rect 2425 8525 3235 8565
rect 3275 8525 5645 8565
rect 5685 8525 6300 8565
rect 6340 8525 6590 8565
rect 6630 8525 7270 8565
rect 7310 8525 7620 8565
rect 7660 8525 8320 8565
rect 8360 8525 8670 8565
rect 8710 8525 9020 8565
rect 9060 8525 9100 8565
rect -1675 8500 9100 8525
rect -1675 8485 -80 8500
rect -4840 8460 -80 8485
rect -40 8460 270 8500
rect 310 8460 620 8500
rect 660 8460 1320 8500
rect 1360 8460 1670 8500
rect 1710 8460 2385 8500
rect 2425 8460 3235 8500
rect 3275 8460 5645 8500
rect 5685 8460 6300 8500
rect 6340 8460 6590 8500
rect 6630 8460 7270 8500
rect 7310 8460 7620 8500
rect 7660 8460 8320 8500
rect 8360 8460 8670 8500
rect 8710 8460 9020 8500
rect 9060 8460 9100 8500
rect -4840 8440 9100 8460
rect -4840 8415 -80 8440
rect -4840 8365 -4805 8415
rect -4755 8365 -4710 8415
rect -4660 8365 -4615 8415
rect -4565 8365 -4515 8415
rect -4465 8365 -4415 8415
rect -4365 8365 -4315 8415
rect -4265 8365 -4220 8415
rect -4170 8365 -4125 8415
rect -4075 8365 -4005 8415
rect -3955 8365 -3910 8415
rect -3860 8365 -3815 8415
rect -3765 8365 -3715 8415
rect -3665 8365 -3615 8415
rect -3565 8365 -3515 8415
rect -3465 8365 -3420 8415
rect -3370 8365 -3325 8415
rect -3275 8365 -3205 8415
rect -3155 8365 -3110 8415
rect -3060 8365 -3015 8415
rect -2965 8365 -2915 8415
rect -2865 8365 -2815 8415
rect -2765 8365 -2715 8415
rect -2665 8365 -2620 8415
rect -2570 8365 -2525 8415
rect -2475 8365 -2405 8415
rect -2355 8365 -2310 8415
rect -2260 8365 -2215 8415
rect -2165 8365 -2115 8415
rect -2065 8365 -2015 8415
rect -1965 8365 -1915 8415
rect -1865 8365 -1820 8415
rect -1770 8365 -1725 8415
rect -1675 8400 -80 8415
rect -40 8400 270 8440
rect 310 8400 620 8440
rect 660 8400 1320 8440
rect 1360 8400 1670 8440
rect 1710 8400 2385 8440
rect 2425 8400 3235 8440
rect 3275 8400 5645 8440
rect 5685 8400 6300 8440
rect 6340 8400 6590 8440
rect 6630 8400 7270 8440
rect 7310 8400 7620 8440
rect 7660 8400 8320 8440
rect 8360 8400 8670 8440
rect 8710 8400 9020 8440
rect 9060 8400 9100 8440
rect -1675 8375 9100 8400
rect -1675 8365 -80 8375
rect -4840 8335 -80 8365
rect -40 8335 270 8375
rect 310 8335 620 8375
rect 660 8335 1320 8375
rect 1360 8335 1670 8375
rect 1710 8335 2385 8375
rect 2425 8335 3235 8375
rect 3275 8335 5645 8375
rect 5685 8335 6300 8375
rect 6340 8335 6590 8375
rect 6630 8335 7270 8375
rect 7310 8335 7620 8375
rect 7660 8335 8320 8375
rect 8360 8335 8670 8375
rect 8710 8335 9020 8375
rect 9060 8335 9100 8375
rect 12080 8345 12130 8645
rect 14790 8625 20720 8675
rect 14790 8575 14825 8625
rect 14875 8575 14920 8625
rect 14970 8575 15015 8625
rect 15065 8575 15115 8625
rect 15165 8575 15215 8625
rect 15265 8575 15315 8625
rect 15365 8575 15410 8625
rect 15460 8575 15505 8625
rect 15555 8575 15625 8625
rect 15675 8575 15720 8625
rect 15770 8575 15815 8625
rect 15865 8575 15915 8625
rect 15965 8575 16015 8625
rect 16065 8575 16115 8625
rect 16165 8575 16210 8625
rect 16260 8575 16305 8625
rect 16355 8575 16425 8625
rect 16475 8575 16520 8625
rect 16570 8575 16615 8625
rect 16665 8575 16715 8625
rect 16765 8575 16815 8625
rect 16865 8575 16915 8625
rect 16965 8575 17010 8625
rect 17060 8575 17105 8625
rect 17155 8575 17225 8625
rect 17275 8575 17320 8625
rect 17370 8575 17415 8625
rect 17465 8575 17515 8625
rect 17565 8575 17615 8625
rect 17665 8575 17715 8625
rect 17765 8575 17810 8625
rect 17860 8575 17905 8625
rect 17955 8575 20720 8625
rect 14790 8535 20720 8575
rect 14790 8485 14825 8535
rect 14875 8485 14920 8535
rect 14970 8485 15015 8535
rect 15065 8485 15115 8535
rect 15165 8485 15215 8535
rect 15265 8485 15315 8535
rect 15365 8485 15410 8535
rect 15460 8485 15505 8535
rect 15555 8485 15625 8535
rect 15675 8485 15720 8535
rect 15770 8485 15815 8535
rect 15865 8485 15915 8535
rect 15965 8485 16015 8535
rect 16065 8485 16115 8535
rect 16165 8485 16210 8535
rect 16260 8485 16305 8535
rect 16355 8485 16425 8535
rect 16475 8485 16520 8535
rect 16570 8485 16615 8535
rect 16665 8485 16715 8535
rect 16765 8485 16815 8535
rect 16865 8485 16915 8535
rect 16965 8485 17010 8535
rect 17060 8485 17105 8535
rect 17155 8485 17225 8535
rect 17275 8485 17320 8535
rect 17370 8485 17415 8535
rect 17465 8485 17515 8535
rect 17565 8485 17615 8535
rect 17665 8485 17715 8535
rect 17765 8485 17810 8535
rect 17860 8485 17905 8535
rect 17955 8485 20720 8535
rect 14790 8415 20720 8485
rect 14790 8365 14825 8415
rect 14875 8365 14920 8415
rect 14970 8365 15015 8415
rect 15065 8365 15115 8415
rect 15165 8365 15215 8415
rect 15265 8365 15315 8415
rect 15365 8365 15410 8415
rect 15460 8365 15505 8415
rect 15555 8365 15625 8415
rect 15675 8365 15720 8415
rect 15770 8365 15815 8415
rect 15865 8365 15915 8415
rect 15965 8365 16015 8415
rect 16065 8365 16115 8415
rect 16165 8365 16210 8415
rect 16260 8365 16305 8415
rect 16355 8365 16425 8415
rect 16475 8365 16520 8415
rect 16570 8365 16615 8415
rect 16665 8365 16715 8415
rect 16765 8365 16815 8415
rect 16865 8365 16915 8415
rect 16965 8365 17010 8415
rect 17060 8365 17105 8415
rect 17155 8365 17225 8415
rect 17275 8365 17320 8415
rect 17370 8365 17415 8415
rect 17465 8365 17515 8415
rect 17565 8365 17615 8415
rect 17665 8365 17715 8415
rect 17765 8365 17810 8415
rect 17860 8365 17905 8415
rect 17955 8365 20720 8415
rect -4840 8325 9100 8335
rect -4840 8275 -4805 8325
rect -4755 8275 -4710 8325
rect -4660 8275 -4615 8325
rect -4565 8275 -4515 8325
rect -4465 8275 -4415 8325
rect -4365 8275 -4315 8325
rect -4265 8275 -4220 8325
rect -4170 8275 -4125 8325
rect -4075 8275 -4005 8325
rect -3955 8275 -3910 8325
rect -3860 8275 -3815 8325
rect -3765 8275 -3715 8325
rect -3665 8275 -3615 8325
rect -3565 8275 -3515 8325
rect -3465 8275 -3420 8325
rect -3370 8275 -3325 8325
rect -3275 8275 -3205 8325
rect -3155 8275 -3110 8325
rect -3060 8275 -3015 8325
rect -2965 8275 -2915 8325
rect -2865 8275 -2815 8325
rect -2765 8275 -2715 8325
rect -2665 8275 -2620 8325
rect -2570 8275 -2525 8325
rect -2475 8275 -2405 8325
rect -2355 8275 -2310 8325
rect -2260 8275 -2215 8325
rect -2165 8275 -2115 8325
rect -2065 8275 -2015 8325
rect -1965 8275 -1915 8325
rect -1865 8275 -1820 8325
rect -1770 8275 -1725 8325
rect -1675 8305 9100 8325
rect -1675 8275 -80 8305
rect -4840 8265 -80 8275
rect -40 8265 270 8305
rect 310 8265 620 8305
rect 660 8265 1320 8305
rect 1360 8265 1670 8305
rect 1710 8265 2385 8305
rect 2425 8265 3235 8305
rect 3275 8265 5645 8305
rect 5685 8265 6300 8305
rect 6340 8265 6590 8305
rect 6630 8265 7270 8305
rect 7310 8265 7620 8305
rect 7660 8265 8320 8305
rect 8360 8265 8670 8305
rect 8710 8265 9020 8305
rect 9060 8265 9100 8305
rect 9630 8340 14580 8345
rect 9630 8300 9635 8340
rect 9675 8300 9985 8340
rect 10025 8300 10335 8340
rect 10375 8300 10685 8340
rect 10725 8300 11035 8340
rect 11075 8300 11385 8340
rect 11425 8300 11735 8340
rect 11775 8300 12085 8340
rect 12125 8300 12435 8340
rect 12475 8300 12785 8340
rect 12825 8300 13135 8340
rect 13175 8300 13485 8340
rect 13525 8300 13835 8340
rect 13875 8300 14185 8340
rect 14225 8300 14535 8340
rect 14575 8300 14580 8340
rect 9630 8295 14580 8300
rect 14790 8325 20720 8365
rect -4840 8235 9100 8265
rect -4840 8225 -80 8235
rect -4840 8175 -4805 8225
rect -4755 8175 -4710 8225
rect -4660 8175 -4615 8225
rect -4565 8175 -4515 8225
rect -4465 8175 -4415 8225
rect -4365 8175 -4315 8225
rect -4265 8175 -4220 8225
rect -4170 8175 -4125 8225
rect -4075 8175 -4005 8225
rect -3955 8175 -3910 8225
rect -3860 8175 -3815 8225
rect -3765 8175 -3715 8225
rect -3665 8175 -3615 8225
rect -3565 8175 -3515 8225
rect -3465 8175 -3420 8225
rect -3370 8175 -3325 8225
rect -3275 8175 -3205 8225
rect -3155 8175 -3110 8225
rect -3060 8175 -3015 8225
rect -2965 8175 -2915 8225
rect -2865 8175 -2815 8225
rect -2765 8175 -2715 8225
rect -2665 8175 -2620 8225
rect -2570 8175 -2525 8225
rect -2475 8175 -2405 8225
rect -2355 8175 -2310 8225
rect -2260 8175 -2215 8225
rect -2165 8175 -2115 8225
rect -2065 8175 -2015 8225
rect -1965 8175 -1915 8225
rect -1865 8175 -1820 8225
rect -1770 8175 -1725 8225
rect -1675 8195 -80 8225
rect -40 8195 270 8235
rect 310 8195 620 8235
rect 660 8195 1320 8235
rect 1360 8195 1670 8235
rect 1710 8195 2385 8235
rect 2425 8195 3235 8235
rect 3275 8195 5645 8235
rect 5685 8195 6300 8235
rect 6340 8195 6590 8235
rect 6630 8195 7270 8235
rect 7310 8195 7620 8235
rect 7660 8195 8320 8235
rect 8360 8195 8670 8235
rect 8710 8195 9020 8235
rect 9060 8195 9100 8235
rect -1675 8175 9100 8195
rect -4840 8165 9100 8175
rect -4840 8135 -80 8165
rect -4840 8085 -4805 8135
rect -4755 8085 -4710 8135
rect -4660 8085 -4615 8135
rect -4565 8085 -4515 8135
rect -4465 8085 -4415 8135
rect -4365 8085 -4315 8135
rect -4265 8085 -4220 8135
rect -4170 8085 -4125 8135
rect -4075 8085 -4005 8135
rect -3955 8085 -3910 8135
rect -3860 8085 -3815 8135
rect -3765 8085 -3715 8135
rect -3665 8085 -3615 8135
rect -3565 8085 -3515 8135
rect -3465 8085 -3420 8135
rect -3370 8085 -3325 8135
rect -3275 8085 -3205 8135
rect -3155 8085 -3110 8135
rect -3060 8085 -3015 8135
rect -2965 8085 -2915 8135
rect -2865 8085 -2815 8135
rect -2765 8085 -2715 8135
rect -2665 8085 -2620 8135
rect -2570 8085 -2525 8135
rect -2475 8085 -2405 8135
rect -2355 8085 -2310 8135
rect -2260 8085 -2215 8135
rect -2165 8085 -2115 8135
rect -2065 8085 -2015 8135
rect -1965 8085 -1915 8135
rect -1865 8085 -1820 8135
rect -1770 8085 -1725 8135
rect -1675 8125 -80 8135
rect -40 8125 270 8165
rect 310 8125 620 8165
rect 660 8125 1320 8165
rect 1360 8125 1670 8165
rect 1710 8125 2385 8165
rect 2425 8125 3235 8165
rect 3275 8125 5645 8165
rect 5685 8125 6300 8165
rect 6340 8125 6590 8165
rect 6630 8125 7270 8165
rect 7310 8125 7620 8165
rect 7660 8125 8320 8165
rect 8360 8125 8670 8165
rect 8710 8125 9020 8165
rect 9060 8125 9100 8165
rect -1675 8100 9100 8125
rect -1675 8085 -80 8100
rect -4840 8060 -80 8085
rect -40 8060 270 8100
rect 310 8060 620 8100
rect 660 8060 1320 8100
rect 1360 8060 1670 8100
rect 1710 8060 2385 8100
rect 2425 8060 3235 8100
rect 3275 8060 5645 8100
rect 5685 8060 6300 8100
rect 6340 8060 6590 8100
rect 6630 8060 7270 8100
rect 7310 8060 7620 8100
rect 7660 8060 8320 8100
rect 8360 8060 8670 8100
rect 8710 8060 9020 8100
rect 9060 8060 9100 8100
rect -4840 8040 9100 8060
rect -4840 8015 -80 8040
rect -4840 7965 -4805 8015
rect -4755 7965 -4710 8015
rect -4660 7965 -4615 8015
rect -4565 7965 -4515 8015
rect -4465 7965 -4415 8015
rect -4365 7965 -4315 8015
rect -4265 7965 -4220 8015
rect -4170 7965 -4125 8015
rect -4075 7965 -4005 8015
rect -3955 7965 -3910 8015
rect -3860 7965 -3815 8015
rect -3765 7965 -3715 8015
rect -3665 7965 -3615 8015
rect -3565 7965 -3515 8015
rect -3465 7965 -3420 8015
rect -3370 7965 -3325 8015
rect -3275 7965 -3205 8015
rect -3155 7965 -3110 8015
rect -3060 7965 -3015 8015
rect -2965 7965 -2915 8015
rect -2865 7965 -2815 8015
rect -2765 7965 -2715 8015
rect -2665 7965 -2620 8015
rect -2570 7965 -2525 8015
rect -2475 7965 -2405 8015
rect -2355 7965 -2310 8015
rect -2260 7965 -2215 8015
rect -2165 7965 -2115 8015
rect -2065 7965 -2015 8015
rect -1965 7965 -1915 8015
rect -1865 7965 -1820 8015
rect -1770 7965 -1725 8015
rect -1675 8000 -80 8015
rect -40 8000 270 8040
rect 310 8000 620 8040
rect 660 8000 1320 8040
rect 1360 8000 1670 8040
rect 1710 8000 2385 8040
rect 2425 8000 3235 8040
rect 3275 8000 5645 8040
rect 5685 8000 6300 8040
rect 6340 8000 6590 8040
rect 6630 8000 7270 8040
rect 7310 8000 7620 8040
rect 7660 8000 8320 8040
rect 8360 8000 8670 8040
rect 8710 8000 9020 8040
rect 9060 8000 9100 8040
rect -1675 7975 9100 8000
rect 12080 7995 12130 8295
rect 14790 8275 14825 8325
rect 14875 8275 14920 8325
rect 14970 8275 15015 8325
rect 15065 8275 15115 8325
rect 15165 8275 15215 8325
rect 15265 8275 15315 8325
rect 15365 8275 15410 8325
rect 15460 8275 15505 8325
rect 15555 8275 15625 8325
rect 15675 8275 15720 8325
rect 15770 8275 15815 8325
rect 15865 8275 15915 8325
rect 15965 8275 16015 8325
rect 16065 8275 16115 8325
rect 16165 8275 16210 8325
rect 16260 8275 16305 8325
rect 16355 8275 16425 8325
rect 16475 8275 16520 8325
rect 16570 8275 16615 8325
rect 16665 8275 16715 8325
rect 16765 8275 16815 8325
rect 16865 8275 16915 8325
rect 16965 8275 17010 8325
rect 17060 8275 17105 8325
rect 17155 8275 17225 8325
rect 17275 8275 17320 8325
rect 17370 8275 17415 8325
rect 17465 8275 17515 8325
rect 17565 8275 17615 8325
rect 17665 8275 17715 8325
rect 17765 8275 17810 8325
rect 17860 8275 17905 8325
rect 17955 8275 20720 8325
rect 14790 8225 20720 8275
rect 14790 8175 14825 8225
rect 14875 8175 14920 8225
rect 14970 8175 15015 8225
rect 15065 8175 15115 8225
rect 15165 8175 15215 8225
rect 15265 8175 15315 8225
rect 15365 8175 15410 8225
rect 15460 8175 15505 8225
rect 15555 8175 15625 8225
rect 15675 8175 15720 8225
rect 15770 8175 15815 8225
rect 15865 8175 15915 8225
rect 15965 8175 16015 8225
rect 16065 8175 16115 8225
rect 16165 8175 16210 8225
rect 16260 8175 16305 8225
rect 16355 8175 16425 8225
rect 16475 8175 16520 8225
rect 16570 8175 16615 8225
rect 16665 8175 16715 8225
rect 16765 8175 16815 8225
rect 16865 8175 16915 8225
rect 16965 8175 17010 8225
rect 17060 8175 17105 8225
rect 17155 8175 17225 8225
rect 17275 8175 17320 8225
rect 17370 8175 17415 8225
rect 17465 8175 17515 8225
rect 17565 8175 17615 8225
rect 17665 8175 17715 8225
rect 17765 8175 17810 8225
rect 17860 8175 17905 8225
rect 17955 8175 20720 8225
rect 14790 8135 20720 8175
rect 14790 8085 14825 8135
rect 14875 8085 14920 8135
rect 14970 8085 15015 8135
rect 15065 8085 15115 8135
rect 15165 8085 15215 8135
rect 15265 8085 15315 8135
rect 15365 8085 15410 8135
rect 15460 8085 15505 8135
rect 15555 8085 15625 8135
rect 15675 8085 15720 8135
rect 15770 8085 15815 8135
rect 15865 8085 15915 8135
rect 15965 8085 16015 8135
rect 16065 8085 16115 8135
rect 16165 8085 16210 8135
rect 16260 8085 16305 8135
rect 16355 8085 16425 8135
rect 16475 8085 16520 8135
rect 16570 8085 16615 8135
rect 16665 8085 16715 8135
rect 16765 8085 16815 8135
rect 16865 8085 16915 8135
rect 16965 8085 17010 8135
rect 17060 8085 17105 8135
rect 17155 8085 17225 8135
rect 17275 8085 17320 8135
rect 17370 8085 17415 8135
rect 17465 8085 17515 8135
rect 17565 8085 17615 8135
rect 17665 8085 17715 8135
rect 17765 8085 17810 8135
rect 17860 8085 17905 8135
rect 17955 8085 20720 8135
rect 14790 8015 20720 8085
rect -1675 7965 -80 7975
rect -4840 7935 -80 7965
rect -40 7935 270 7975
rect 310 7935 620 7975
rect 660 7935 1320 7975
rect 1360 7935 1670 7975
rect 1710 7935 2385 7975
rect 2425 7935 3235 7975
rect 3275 7935 5645 7975
rect 5685 7935 6300 7975
rect 6340 7935 6590 7975
rect 6630 7935 7270 7975
rect 7310 7935 7620 7975
rect 7660 7935 8320 7975
rect 8360 7935 8670 7975
rect 8710 7935 9020 7975
rect 9060 7935 9100 7975
rect 9630 7990 14580 7995
rect 9630 7950 9635 7990
rect 9675 7950 9985 7990
rect 10025 7950 10335 7990
rect 10375 7950 10685 7990
rect 10725 7950 11035 7990
rect 11075 7950 11385 7990
rect 11425 7950 11735 7990
rect 11775 7950 12085 7990
rect 12125 7950 12435 7990
rect 12475 7950 12785 7990
rect 12825 7950 13135 7990
rect 13175 7950 13485 7990
rect 13525 7950 13835 7990
rect 13875 7950 14185 7990
rect 14225 7950 14535 7990
rect 14575 7950 14580 7990
rect 9630 7945 14580 7950
rect 14790 7965 14825 8015
rect 14875 7965 14920 8015
rect 14970 7965 15015 8015
rect 15065 7965 15115 8015
rect 15165 7965 15215 8015
rect 15265 7965 15315 8015
rect 15365 7965 15410 8015
rect 15460 7965 15505 8015
rect 15555 7965 15625 8015
rect 15675 7965 15720 8015
rect 15770 7965 15815 8015
rect 15865 7965 15915 8015
rect 15965 7965 16015 8015
rect 16065 7965 16115 8015
rect 16165 7965 16210 8015
rect 16260 7965 16305 8015
rect 16355 7965 16425 8015
rect 16475 7965 16520 8015
rect 16570 7965 16615 8015
rect 16665 7965 16715 8015
rect 16765 7965 16815 8015
rect 16865 7965 16915 8015
rect 16965 7965 17010 8015
rect 17060 7965 17105 8015
rect 17155 7965 17225 8015
rect 17275 7965 17320 8015
rect 17370 7965 17415 8015
rect 17465 7965 17515 8015
rect 17565 7965 17615 8015
rect 17665 7965 17715 8015
rect 17765 7965 17810 8015
rect 17860 7965 17905 8015
rect 17955 7965 20720 8015
rect -4840 7925 9100 7935
rect -4840 7875 -4805 7925
rect -4755 7875 -4710 7925
rect -4660 7875 -4615 7925
rect -4565 7875 -4515 7925
rect -4465 7875 -4415 7925
rect -4365 7875 -4315 7925
rect -4265 7875 -4220 7925
rect -4170 7875 -4125 7925
rect -4075 7875 -4005 7925
rect -3955 7875 -3910 7925
rect -3860 7875 -3815 7925
rect -3765 7875 -3715 7925
rect -3665 7875 -3615 7925
rect -3565 7875 -3515 7925
rect -3465 7875 -3420 7925
rect -3370 7875 -3325 7925
rect -3275 7875 -3205 7925
rect -3155 7875 -3110 7925
rect -3060 7875 -3015 7925
rect -2965 7875 -2915 7925
rect -2865 7875 -2815 7925
rect -2765 7875 -2715 7925
rect -2665 7875 -2620 7925
rect -2570 7875 -2525 7925
rect -2475 7875 -2405 7925
rect -2355 7875 -2310 7925
rect -2260 7875 -2215 7925
rect -2165 7875 -2115 7925
rect -2065 7875 -2015 7925
rect -1965 7875 -1915 7925
rect -1865 7875 -1820 7925
rect -1770 7875 -1725 7925
rect -1675 7905 9100 7925
rect -1675 7875 -80 7905
rect -4840 7865 -80 7875
rect -40 7865 270 7905
rect 310 7865 620 7905
rect 660 7865 1320 7905
rect 1360 7865 1670 7905
rect 1710 7865 2385 7905
rect 2425 7865 3235 7905
rect 3275 7865 5645 7905
rect 5685 7865 6300 7905
rect 6340 7865 6590 7905
rect 6630 7865 7270 7905
rect 7310 7865 7620 7905
rect 7660 7865 8320 7905
rect 8360 7865 8670 7905
rect 8710 7865 9020 7905
rect 9060 7865 9100 7905
rect -4840 7835 9100 7865
rect -4840 7825 -80 7835
rect -4840 7775 -4805 7825
rect -4755 7775 -4710 7825
rect -4660 7775 -4615 7825
rect -4565 7775 -4515 7825
rect -4465 7775 -4415 7825
rect -4365 7775 -4315 7825
rect -4265 7775 -4220 7825
rect -4170 7775 -4125 7825
rect -4075 7775 -4005 7825
rect -3955 7775 -3910 7825
rect -3860 7775 -3815 7825
rect -3765 7775 -3715 7825
rect -3665 7775 -3615 7825
rect -3565 7775 -3515 7825
rect -3465 7775 -3420 7825
rect -3370 7775 -3325 7825
rect -3275 7775 -3205 7825
rect -3155 7775 -3110 7825
rect -3060 7775 -3015 7825
rect -2965 7775 -2915 7825
rect -2865 7775 -2815 7825
rect -2765 7775 -2715 7825
rect -2665 7775 -2620 7825
rect -2570 7775 -2525 7825
rect -2475 7775 -2405 7825
rect -2355 7775 -2310 7825
rect -2260 7775 -2215 7825
rect -2165 7775 -2115 7825
rect -2065 7775 -2015 7825
rect -1965 7775 -1915 7825
rect -1865 7775 -1820 7825
rect -1770 7775 -1725 7825
rect -1675 7795 -80 7825
rect -40 7795 270 7835
rect 310 7795 620 7835
rect 660 7795 1320 7835
rect 1360 7795 1670 7835
rect 1710 7795 2385 7835
rect 2425 7795 3235 7835
rect 3275 7795 5645 7835
rect 5685 7795 6300 7835
rect 6340 7795 6590 7835
rect 6630 7795 7270 7835
rect 7310 7795 7620 7835
rect 7660 7795 8320 7835
rect 8360 7795 8670 7835
rect 8710 7795 9020 7835
rect 9060 7795 9100 7835
rect -1675 7775 9100 7795
rect -4840 7765 9100 7775
rect -4840 7735 -80 7765
rect -4840 7685 -4805 7735
rect -4755 7685 -4710 7735
rect -4660 7685 -4615 7735
rect -4565 7685 -4515 7735
rect -4465 7685 -4415 7735
rect -4365 7685 -4315 7735
rect -4265 7685 -4220 7735
rect -4170 7685 -4125 7735
rect -4075 7685 -4005 7735
rect -3955 7685 -3910 7735
rect -3860 7685 -3815 7735
rect -3765 7685 -3715 7735
rect -3665 7685 -3615 7735
rect -3565 7685 -3515 7735
rect -3465 7685 -3420 7735
rect -3370 7685 -3325 7735
rect -3275 7685 -3205 7735
rect -3155 7685 -3110 7735
rect -3060 7685 -3015 7735
rect -2965 7685 -2915 7735
rect -2865 7685 -2815 7735
rect -2765 7685 -2715 7735
rect -2665 7685 -2620 7735
rect -2570 7685 -2525 7735
rect -2475 7685 -2405 7735
rect -2355 7685 -2310 7735
rect -2260 7685 -2215 7735
rect -2165 7685 -2115 7735
rect -2065 7685 -2015 7735
rect -1965 7685 -1915 7735
rect -1865 7685 -1820 7735
rect -1770 7685 -1725 7735
rect -1675 7725 -80 7735
rect -40 7725 270 7765
rect 310 7725 620 7765
rect 660 7725 1320 7765
rect 1360 7725 1670 7765
rect 1710 7725 2385 7765
rect 2425 7725 3235 7765
rect 3275 7725 5645 7765
rect 5685 7725 6300 7765
rect 6340 7725 6590 7765
rect 6630 7725 7270 7765
rect 7310 7725 7620 7765
rect 7660 7725 8320 7765
rect 8360 7725 8670 7765
rect 8710 7725 9020 7765
rect 9060 7725 9100 7765
rect -1675 7700 9100 7725
rect -1675 7685 -80 7700
rect -4840 7660 -80 7685
rect -40 7660 270 7700
rect 310 7660 620 7700
rect 660 7660 1320 7700
rect 1360 7660 1670 7700
rect 1710 7660 2385 7700
rect 2425 7660 3235 7700
rect 3275 7660 5645 7700
rect 5685 7660 6300 7700
rect 6340 7660 6590 7700
rect 6630 7660 7270 7700
rect 7310 7660 7620 7700
rect 7660 7660 8320 7700
rect 8360 7660 8670 7700
rect 8710 7660 9020 7700
rect 9060 7660 9100 7700
rect -4840 7640 9100 7660
rect 12080 7645 12130 7945
rect 14790 7925 20720 7965
rect 14790 7875 14825 7925
rect 14875 7875 14920 7925
rect 14970 7875 15015 7925
rect 15065 7875 15115 7925
rect 15165 7875 15215 7925
rect 15265 7875 15315 7925
rect 15365 7875 15410 7925
rect 15460 7875 15505 7925
rect 15555 7875 15625 7925
rect 15675 7875 15720 7925
rect 15770 7875 15815 7925
rect 15865 7875 15915 7925
rect 15965 7875 16015 7925
rect 16065 7875 16115 7925
rect 16165 7875 16210 7925
rect 16260 7875 16305 7925
rect 16355 7875 16425 7925
rect 16475 7875 16520 7925
rect 16570 7875 16615 7925
rect 16665 7875 16715 7925
rect 16765 7875 16815 7925
rect 16865 7875 16915 7925
rect 16965 7875 17010 7925
rect 17060 7875 17105 7925
rect 17155 7875 17225 7925
rect 17275 7875 17320 7925
rect 17370 7875 17415 7925
rect 17465 7875 17515 7925
rect 17565 7875 17615 7925
rect 17665 7875 17715 7925
rect 17765 7875 17810 7925
rect 17860 7875 17905 7925
rect 17955 7875 20720 7925
rect 14790 7825 20720 7875
rect 14790 7775 14825 7825
rect 14875 7775 14920 7825
rect 14970 7775 15015 7825
rect 15065 7775 15115 7825
rect 15165 7775 15215 7825
rect 15265 7775 15315 7825
rect 15365 7775 15410 7825
rect 15460 7775 15505 7825
rect 15555 7775 15625 7825
rect 15675 7775 15720 7825
rect 15770 7775 15815 7825
rect 15865 7775 15915 7825
rect 15965 7775 16015 7825
rect 16065 7775 16115 7825
rect 16165 7775 16210 7825
rect 16260 7775 16305 7825
rect 16355 7775 16425 7825
rect 16475 7775 16520 7825
rect 16570 7775 16615 7825
rect 16665 7775 16715 7825
rect 16765 7775 16815 7825
rect 16865 7775 16915 7825
rect 16965 7775 17010 7825
rect 17060 7775 17105 7825
rect 17155 7775 17225 7825
rect 17275 7775 17320 7825
rect 17370 7775 17415 7825
rect 17465 7775 17515 7825
rect 17565 7775 17615 7825
rect 17665 7775 17715 7825
rect 17765 7775 17810 7825
rect 17860 7775 17905 7825
rect 17955 7775 20720 7825
rect 14790 7735 20720 7775
rect 14790 7685 14825 7735
rect 14875 7685 14920 7735
rect 14970 7685 15015 7735
rect 15065 7685 15115 7735
rect 15165 7685 15215 7735
rect 15265 7685 15315 7735
rect 15365 7685 15410 7735
rect 15460 7685 15505 7735
rect 15555 7685 15625 7735
rect 15675 7685 15720 7735
rect 15770 7685 15815 7735
rect 15865 7685 15915 7735
rect 15965 7685 16015 7735
rect 16065 7685 16115 7735
rect 16165 7685 16210 7735
rect 16260 7685 16305 7735
rect 16355 7685 16425 7735
rect 16475 7685 16520 7735
rect 16570 7685 16615 7735
rect 16665 7685 16715 7735
rect 16765 7685 16815 7735
rect 16865 7685 16915 7735
rect 16965 7685 17010 7735
rect 17060 7685 17105 7735
rect 17155 7685 17225 7735
rect 17275 7685 17320 7735
rect 17370 7685 17415 7735
rect 17465 7685 17515 7735
rect 17565 7685 17615 7735
rect 17665 7685 17715 7735
rect 17765 7685 17810 7735
rect 17860 7685 17905 7735
rect 17955 7685 20720 7735
rect -4840 7615 -80 7640
rect -4840 7565 -4805 7615
rect -4755 7565 -4710 7615
rect -4660 7565 -4615 7615
rect -4565 7565 -4515 7615
rect -4465 7565 -4415 7615
rect -4365 7565 -4315 7615
rect -4265 7565 -4220 7615
rect -4170 7565 -4125 7615
rect -4075 7565 -4005 7615
rect -3955 7565 -3910 7615
rect -3860 7565 -3815 7615
rect -3765 7565 -3715 7615
rect -3665 7565 -3615 7615
rect -3565 7565 -3515 7615
rect -3465 7565 -3420 7615
rect -3370 7565 -3325 7615
rect -3275 7565 -3205 7615
rect -3155 7565 -3110 7615
rect -3060 7565 -3015 7615
rect -2965 7565 -2915 7615
rect -2865 7565 -2815 7615
rect -2765 7565 -2715 7615
rect -2665 7565 -2620 7615
rect -2570 7565 -2525 7615
rect -2475 7565 -2405 7615
rect -2355 7565 -2310 7615
rect -2260 7565 -2215 7615
rect -2165 7565 -2115 7615
rect -2065 7565 -2015 7615
rect -1965 7565 -1915 7615
rect -1865 7565 -1820 7615
rect -1770 7565 -1725 7615
rect -1675 7600 -80 7615
rect -40 7600 270 7640
rect 310 7600 620 7640
rect 660 7600 1320 7640
rect 1360 7600 1670 7640
rect 1710 7600 2385 7640
rect 2425 7600 3235 7640
rect 3275 7600 5645 7640
rect 5685 7600 6300 7640
rect 6340 7600 6590 7640
rect 6630 7600 7270 7640
rect 7310 7600 7620 7640
rect 7660 7600 8320 7640
rect 8360 7600 8670 7640
rect 8710 7600 9020 7640
rect 9060 7600 9100 7640
rect -1675 7575 9100 7600
rect 9630 7640 14580 7645
rect 9630 7600 9635 7640
rect 9675 7600 9985 7640
rect 10025 7600 10335 7640
rect 10375 7600 10685 7640
rect 10725 7600 11035 7640
rect 11075 7600 11385 7640
rect 11425 7600 11735 7640
rect 11775 7600 12085 7640
rect 12125 7600 12435 7640
rect 12475 7600 12785 7640
rect 12825 7600 13135 7640
rect 13175 7600 13485 7640
rect 13525 7600 13835 7640
rect 13875 7600 14185 7640
rect 14225 7600 14535 7640
rect 14575 7600 14580 7640
rect 9630 7595 14580 7600
rect 14790 7615 20720 7685
rect -1675 7565 -80 7575
rect -4840 7535 -80 7565
rect -40 7535 270 7575
rect 310 7535 620 7575
rect 660 7535 1320 7575
rect 1360 7535 1670 7575
rect 1710 7535 2385 7575
rect 2425 7535 3235 7575
rect 3275 7535 5645 7575
rect 5685 7535 6300 7575
rect 6340 7535 6590 7575
rect 6630 7535 7270 7575
rect 7310 7535 7620 7575
rect 7660 7535 8320 7575
rect 8360 7535 8670 7575
rect 8710 7535 9020 7575
rect 9060 7535 9100 7575
rect -4840 7525 9100 7535
rect -4840 7475 -4805 7525
rect -4755 7475 -4710 7525
rect -4660 7475 -4615 7525
rect -4565 7475 -4515 7525
rect -4465 7475 -4415 7525
rect -4365 7475 -4315 7525
rect -4265 7475 -4220 7525
rect -4170 7475 -4125 7525
rect -4075 7475 -4005 7525
rect -3955 7475 -3910 7525
rect -3860 7475 -3815 7525
rect -3765 7475 -3715 7525
rect -3665 7475 -3615 7525
rect -3565 7475 -3515 7525
rect -3465 7475 -3420 7525
rect -3370 7475 -3325 7525
rect -3275 7475 -3205 7525
rect -3155 7475 -3110 7525
rect -3060 7475 -3015 7525
rect -2965 7475 -2915 7525
rect -2865 7475 -2815 7525
rect -2765 7475 -2715 7525
rect -2665 7475 -2620 7525
rect -2570 7475 -2525 7525
rect -2475 7475 -2405 7525
rect -2355 7475 -2310 7525
rect -2260 7475 -2215 7525
rect -2165 7475 -2115 7525
rect -2065 7475 -2015 7525
rect -1965 7475 -1915 7525
rect -1865 7475 -1820 7525
rect -1770 7475 -1725 7525
rect -1675 7505 9100 7525
rect -1675 7475 -80 7505
rect -4840 7465 -80 7475
rect -40 7465 270 7505
rect 310 7465 620 7505
rect 660 7465 1320 7505
rect 1360 7465 1670 7505
rect 1710 7465 2385 7505
rect 2425 7465 3235 7505
rect 3275 7465 5645 7505
rect 5685 7465 6300 7505
rect 6340 7465 6590 7505
rect 6630 7465 7270 7505
rect 7310 7465 7620 7505
rect 7660 7465 8320 7505
rect 8360 7465 8670 7505
rect 8710 7465 9020 7505
rect 9060 7465 9100 7505
rect -4840 7435 9100 7465
rect -4840 7425 -80 7435
rect -4840 7375 -4805 7425
rect -4755 7375 -4710 7425
rect -4660 7375 -4615 7425
rect -4565 7375 -4515 7425
rect -4465 7375 -4415 7425
rect -4365 7375 -4315 7425
rect -4265 7375 -4220 7425
rect -4170 7375 -4125 7425
rect -4075 7375 -4005 7425
rect -3955 7375 -3910 7425
rect -3860 7375 -3815 7425
rect -3765 7375 -3715 7425
rect -3665 7375 -3615 7425
rect -3565 7375 -3515 7425
rect -3465 7375 -3420 7425
rect -3370 7375 -3325 7425
rect -3275 7375 -3205 7425
rect -3155 7375 -3110 7425
rect -3060 7375 -3015 7425
rect -2965 7375 -2915 7425
rect -2865 7375 -2815 7425
rect -2765 7375 -2715 7425
rect -2665 7375 -2620 7425
rect -2570 7375 -2525 7425
rect -2475 7375 -2405 7425
rect -2355 7375 -2310 7425
rect -2260 7375 -2215 7425
rect -2165 7375 -2115 7425
rect -2065 7375 -2015 7425
rect -1965 7375 -1915 7425
rect -1865 7375 -1820 7425
rect -1770 7375 -1725 7425
rect -1675 7395 -80 7425
rect -40 7395 270 7435
rect 310 7395 620 7435
rect 660 7395 1320 7435
rect 1360 7395 1670 7435
rect 1710 7395 2385 7435
rect 2425 7395 3235 7435
rect 3275 7395 5645 7435
rect 5685 7395 6300 7435
rect 6340 7395 6590 7435
rect 6630 7395 7270 7435
rect 7310 7395 7620 7435
rect 7660 7395 8320 7435
rect 8360 7395 8670 7435
rect 8710 7395 9020 7435
rect 9060 7395 9100 7435
rect -1675 7375 9100 7395
rect -4840 7365 9100 7375
rect -4840 7335 -80 7365
rect -4840 7285 -4805 7335
rect -4755 7285 -4710 7335
rect -4660 7285 -4615 7335
rect -4565 7285 -4515 7335
rect -4465 7285 -4415 7335
rect -4365 7285 -4315 7335
rect -4265 7285 -4220 7335
rect -4170 7285 -4125 7335
rect -4075 7285 -4005 7335
rect -3955 7285 -3910 7335
rect -3860 7285 -3815 7335
rect -3765 7285 -3715 7335
rect -3665 7285 -3615 7335
rect -3565 7285 -3515 7335
rect -3465 7285 -3420 7335
rect -3370 7285 -3325 7335
rect -3275 7285 -3205 7335
rect -3155 7285 -3110 7335
rect -3060 7285 -3015 7335
rect -2965 7285 -2915 7335
rect -2865 7285 -2815 7335
rect -2765 7285 -2715 7335
rect -2665 7285 -2620 7335
rect -2570 7285 -2525 7335
rect -2475 7285 -2405 7335
rect -2355 7285 -2310 7335
rect -2260 7285 -2215 7335
rect -2165 7285 -2115 7335
rect -2065 7285 -2015 7335
rect -1965 7285 -1915 7335
rect -1865 7285 -1820 7335
rect -1770 7285 -1725 7335
rect -1675 7325 -80 7335
rect -40 7325 270 7365
rect 310 7325 620 7365
rect 660 7325 1320 7365
rect 1360 7325 1670 7365
rect 1710 7325 2385 7365
rect 2425 7325 3235 7365
rect 3275 7325 5645 7365
rect 5685 7325 6300 7365
rect 6340 7325 6590 7365
rect 6630 7325 7270 7365
rect 7310 7325 7620 7365
rect 7660 7325 8320 7365
rect 8360 7325 8670 7365
rect 8710 7325 9020 7365
rect 9060 7325 9100 7365
rect -1675 7300 9100 7325
rect -1675 7285 -80 7300
rect -4840 7260 -80 7285
rect -40 7260 270 7300
rect 310 7260 620 7300
rect 660 7260 1320 7300
rect 1360 7260 1670 7300
rect 1710 7260 2385 7300
rect 2425 7260 3235 7300
rect 3275 7260 5645 7300
rect 5685 7260 6300 7300
rect 6340 7260 6590 7300
rect 6630 7260 7270 7300
rect 7310 7260 7620 7300
rect 7660 7260 8320 7300
rect 8360 7260 8670 7300
rect 8710 7260 9020 7300
rect 9060 7260 9100 7300
rect 12080 7295 12130 7595
rect 14790 7565 14825 7615
rect 14875 7565 14920 7615
rect 14970 7565 15015 7615
rect 15065 7565 15115 7615
rect 15165 7565 15215 7615
rect 15265 7565 15315 7615
rect 15365 7565 15410 7615
rect 15460 7565 15505 7615
rect 15555 7565 15625 7615
rect 15675 7565 15720 7615
rect 15770 7565 15815 7615
rect 15865 7565 15915 7615
rect 15965 7565 16015 7615
rect 16065 7565 16115 7615
rect 16165 7565 16210 7615
rect 16260 7565 16305 7615
rect 16355 7565 16425 7615
rect 16475 7565 16520 7615
rect 16570 7565 16615 7615
rect 16665 7565 16715 7615
rect 16765 7565 16815 7615
rect 16865 7565 16915 7615
rect 16965 7565 17010 7615
rect 17060 7565 17105 7615
rect 17155 7565 17225 7615
rect 17275 7565 17320 7615
rect 17370 7565 17415 7615
rect 17465 7565 17515 7615
rect 17565 7565 17615 7615
rect 17665 7565 17715 7615
rect 17765 7565 17810 7615
rect 17860 7565 17905 7615
rect 17955 7565 20720 7615
rect 14790 7525 20720 7565
rect 14790 7475 14825 7525
rect 14875 7475 14920 7525
rect 14970 7475 15015 7525
rect 15065 7475 15115 7525
rect 15165 7475 15215 7525
rect 15265 7475 15315 7525
rect 15365 7475 15410 7525
rect 15460 7475 15505 7525
rect 15555 7475 15625 7525
rect 15675 7475 15720 7525
rect 15770 7475 15815 7525
rect 15865 7475 15915 7525
rect 15965 7475 16015 7525
rect 16065 7475 16115 7525
rect 16165 7475 16210 7525
rect 16260 7475 16305 7525
rect 16355 7475 16425 7525
rect 16475 7475 16520 7525
rect 16570 7475 16615 7525
rect 16665 7475 16715 7525
rect 16765 7475 16815 7525
rect 16865 7475 16915 7525
rect 16965 7475 17010 7525
rect 17060 7475 17105 7525
rect 17155 7475 17225 7525
rect 17275 7475 17320 7525
rect 17370 7475 17415 7525
rect 17465 7475 17515 7525
rect 17565 7475 17615 7525
rect 17665 7475 17715 7525
rect 17765 7475 17810 7525
rect 17860 7475 17905 7525
rect 17955 7475 20720 7525
rect 14790 7425 20720 7475
rect 14790 7375 14825 7425
rect 14875 7375 14920 7425
rect 14970 7375 15015 7425
rect 15065 7375 15115 7425
rect 15165 7375 15215 7425
rect 15265 7375 15315 7425
rect 15365 7375 15410 7425
rect 15460 7375 15505 7425
rect 15555 7375 15625 7425
rect 15675 7375 15720 7425
rect 15770 7375 15815 7425
rect 15865 7375 15915 7425
rect 15965 7375 16015 7425
rect 16065 7375 16115 7425
rect 16165 7375 16210 7425
rect 16260 7375 16305 7425
rect 16355 7375 16425 7425
rect 16475 7375 16520 7425
rect 16570 7375 16615 7425
rect 16665 7375 16715 7425
rect 16765 7375 16815 7425
rect 16865 7375 16915 7425
rect 16965 7375 17010 7425
rect 17060 7375 17105 7425
rect 17155 7375 17225 7425
rect 17275 7375 17320 7425
rect 17370 7375 17415 7425
rect 17465 7375 17515 7425
rect 17565 7375 17615 7425
rect 17665 7375 17715 7425
rect 17765 7375 17810 7425
rect 17860 7375 17905 7425
rect 17955 7375 20720 7425
rect 14790 7335 20720 7375
rect -4840 7240 9100 7260
rect 9630 7290 14580 7295
rect 9630 7250 9635 7290
rect 9675 7250 9985 7290
rect 10025 7250 10335 7290
rect 10375 7250 10685 7290
rect 10725 7250 11035 7290
rect 11075 7250 11385 7290
rect 11425 7250 11735 7290
rect 11775 7250 12085 7290
rect 12125 7250 12435 7290
rect 12475 7250 12785 7290
rect 12825 7250 13135 7290
rect 13175 7250 13485 7290
rect 13525 7250 13835 7290
rect 13875 7250 14185 7290
rect 14225 7250 14535 7290
rect 14575 7250 14580 7290
rect 9630 7245 14580 7250
rect 14790 7285 14825 7335
rect 14875 7285 14920 7335
rect 14970 7285 15015 7335
rect 15065 7285 15115 7335
rect 15165 7285 15215 7335
rect 15265 7285 15315 7335
rect 15365 7285 15410 7335
rect 15460 7285 15505 7335
rect 15555 7285 15625 7335
rect 15675 7285 15720 7335
rect 15770 7285 15815 7335
rect 15865 7285 15915 7335
rect 15965 7285 16015 7335
rect 16065 7285 16115 7335
rect 16165 7285 16210 7335
rect 16260 7285 16305 7335
rect 16355 7285 16425 7335
rect 16475 7285 16520 7335
rect 16570 7285 16615 7335
rect 16665 7285 16715 7335
rect 16765 7285 16815 7335
rect 16865 7285 16915 7335
rect 16965 7285 17010 7335
rect 17060 7285 17105 7335
rect 17155 7285 17225 7335
rect 17275 7285 17320 7335
rect 17370 7285 17415 7335
rect 17465 7285 17515 7335
rect 17565 7285 17615 7335
rect 17665 7285 17715 7335
rect 17765 7285 17810 7335
rect 17860 7285 17905 7335
rect 17955 7285 20720 7335
rect -4840 7215 -80 7240
rect -4840 7165 -4805 7215
rect -4755 7165 -4710 7215
rect -4660 7165 -4615 7215
rect -4565 7165 -4515 7215
rect -4465 7165 -4415 7215
rect -4365 7165 -4315 7215
rect -4265 7165 -4220 7215
rect -4170 7165 -4125 7215
rect -4075 7165 -4005 7215
rect -3955 7165 -3910 7215
rect -3860 7165 -3815 7215
rect -3765 7165 -3715 7215
rect -3665 7165 -3615 7215
rect -3565 7165 -3515 7215
rect -3465 7165 -3420 7215
rect -3370 7165 -3325 7215
rect -3275 7165 -3205 7215
rect -3155 7165 -3110 7215
rect -3060 7165 -3015 7215
rect -2965 7165 -2915 7215
rect -2865 7165 -2815 7215
rect -2765 7165 -2715 7215
rect -2665 7165 -2620 7215
rect -2570 7165 -2525 7215
rect -2475 7165 -2405 7215
rect -2355 7165 -2310 7215
rect -2260 7165 -2215 7215
rect -2165 7165 -2115 7215
rect -2065 7165 -2015 7215
rect -1965 7165 -1915 7215
rect -1865 7165 -1820 7215
rect -1770 7165 -1725 7215
rect -1675 7200 -80 7215
rect -40 7200 270 7240
rect 310 7200 620 7240
rect 660 7200 1320 7240
rect 1360 7200 1670 7240
rect 1710 7200 2385 7240
rect 2425 7200 3235 7240
rect 3275 7200 5645 7240
rect 5685 7200 6300 7240
rect 6340 7200 6590 7240
rect 6630 7200 7270 7240
rect 7310 7200 7620 7240
rect 7660 7200 8320 7240
rect 8360 7200 8670 7240
rect 8710 7200 9020 7240
rect 9060 7200 9100 7240
rect -1675 7175 9100 7200
rect -1675 7165 -80 7175
rect -4840 7135 -80 7165
rect -40 7135 270 7175
rect 310 7135 620 7175
rect 660 7135 1320 7175
rect 1360 7135 1670 7175
rect 1710 7135 2385 7175
rect 2425 7135 3235 7175
rect 3275 7135 5645 7175
rect 5685 7135 6300 7175
rect 6340 7135 6590 7175
rect 6630 7135 7270 7175
rect 7310 7135 7620 7175
rect 7660 7135 8320 7175
rect 8360 7135 8670 7175
rect 8710 7135 9020 7175
rect 9060 7135 9100 7175
rect -4840 7125 9100 7135
rect -4840 7075 -4805 7125
rect -4755 7075 -4710 7125
rect -4660 7075 -4615 7125
rect -4565 7075 -4515 7125
rect -4465 7075 -4415 7125
rect -4365 7075 -4315 7125
rect -4265 7075 -4220 7125
rect -4170 7075 -4125 7125
rect -4075 7075 -4005 7125
rect -3955 7075 -3910 7125
rect -3860 7075 -3815 7125
rect -3765 7075 -3715 7125
rect -3665 7075 -3615 7125
rect -3565 7075 -3515 7125
rect -3465 7075 -3420 7125
rect -3370 7075 -3325 7125
rect -3275 7075 -3205 7125
rect -3155 7075 -3110 7125
rect -3060 7075 -3015 7125
rect -2965 7075 -2915 7125
rect -2865 7075 -2815 7125
rect -2765 7075 -2715 7125
rect -2665 7075 -2620 7125
rect -2570 7075 -2525 7125
rect -2475 7075 -2405 7125
rect -2355 7075 -2310 7125
rect -2260 7075 -2215 7125
rect -2165 7075 -2115 7125
rect -2065 7075 -2015 7125
rect -1965 7075 -1915 7125
rect -1865 7075 -1820 7125
rect -1770 7075 -1725 7125
rect -1675 7105 9100 7125
rect -1675 7075 -80 7105
rect -4840 7065 -80 7075
rect -40 7065 270 7105
rect 310 7065 620 7105
rect 660 7065 1320 7105
rect 1360 7065 1670 7105
rect 1710 7065 2385 7105
rect 2425 7065 3235 7105
rect 3275 7065 5645 7105
rect 5685 7065 6300 7105
rect 6340 7065 6590 7105
rect 6630 7065 7270 7105
rect 7310 7065 7620 7105
rect 7660 7065 8320 7105
rect 8360 7065 8670 7105
rect 8710 7065 9020 7105
rect 9060 7065 9100 7105
rect -4840 7035 9100 7065
rect -4840 7025 -80 7035
rect -4840 6975 -4805 7025
rect -4755 6975 -4710 7025
rect -4660 6975 -4615 7025
rect -4565 6975 -4515 7025
rect -4465 6975 -4415 7025
rect -4365 6975 -4315 7025
rect -4265 6975 -4220 7025
rect -4170 6975 -4125 7025
rect -4075 6975 -4005 7025
rect -3955 6975 -3910 7025
rect -3860 6975 -3815 7025
rect -3765 6975 -3715 7025
rect -3665 6975 -3615 7025
rect -3565 6975 -3515 7025
rect -3465 6975 -3420 7025
rect -3370 6975 -3325 7025
rect -3275 6975 -3205 7025
rect -3155 6975 -3110 7025
rect -3060 6975 -3015 7025
rect -2965 6975 -2915 7025
rect -2865 6975 -2815 7025
rect -2765 6975 -2715 7025
rect -2665 6975 -2620 7025
rect -2570 6975 -2525 7025
rect -2475 6975 -2405 7025
rect -2355 6975 -2310 7025
rect -2260 6975 -2215 7025
rect -2165 6975 -2115 7025
rect -2065 6975 -2015 7025
rect -1965 6975 -1915 7025
rect -1865 6975 -1820 7025
rect -1770 6975 -1725 7025
rect -1675 6995 -80 7025
rect -40 6995 270 7035
rect 310 6995 620 7035
rect 660 6995 1320 7035
rect 1360 6995 1670 7035
rect 1710 6995 2385 7035
rect 2425 6995 3235 7035
rect 3275 6995 5645 7035
rect 5685 6995 6300 7035
rect 6340 6995 6590 7035
rect 6630 6995 7270 7035
rect 7310 6995 7620 7035
rect 7660 6995 8320 7035
rect 8360 6995 8670 7035
rect 8710 6995 9020 7035
rect 9060 6995 9100 7035
rect -1675 6975 9100 6995
rect -4840 6965 9100 6975
rect -4840 6935 -80 6965
rect -4840 6885 -4805 6935
rect -4755 6885 -4710 6935
rect -4660 6885 -4615 6935
rect -4565 6885 -4515 6935
rect -4465 6885 -4415 6935
rect -4365 6885 -4315 6935
rect -4265 6885 -4220 6935
rect -4170 6885 -4125 6935
rect -4075 6885 -4005 6935
rect -3955 6885 -3910 6935
rect -3860 6885 -3815 6935
rect -3765 6885 -3715 6935
rect -3665 6885 -3615 6935
rect -3565 6885 -3515 6935
rect -3465 6885 -3420 6935
rect -3370 6885 -3325 6935
rect -3275 6885 -3205 6935
rect -3155 6885 -3110 6935
rect -3060 6885 -3015 6935
rect -2965 6885 -2915 6935
rect -2865 6885 -2815 6935
rect -2765 6885 -2715 6935
rect -2665 6885 -2620 6935
rect -2570 6885 -2525 6935
rect -2475 6885 -2405 6935
rect -2355 6885 -2310 6935
rect -2260 6885 -2215 6935
rect -2165 6885 -2115 6935
rect -2065 6885 -2015 6935
rect -1965 6885 -1915 6935
rect -1865 6885 -1820 6935
rect -1770 6885 -1725 6935
rect -1675 6925 -80 6935
rect -40 6925 270 6965
rect 310 6925 620 6965
rect 660 6925 1320 6965
rect 1360 6925 1670 6965
rect 1710 6925 2385 6965
rect 2425 6925 3235 6965
rect 3275 6925 5645 6965
rect 5685 6925 6300 6965
rect 6340 6925 6590 6965
rect 6630 6925 7270 6965
rect 7310 6925 7620 6965
rect 7660 6925 8320 6965
rect 8360 6925 8670 6965
rect 8710 6925 9020 6965
rect 9060 6925 9100 6965
rect 12080 6945 12130 7245
rect 14790 7215 20720 7285
rect 14790 7165 14825 7215
rect 14875 7165 14920 7215
rect 14970 7165 15015 7215
rect 15065 7165 15115 7215
rect 15165 7165 15215 7215
rect 15265 7165 15315 7215
rect 15365 7165 15410 7215
rect 15460 7165 15505 7215
rect 15555 7165 15625 7215
rect 15675 7165 15720 7215
rect 15770 7165 15815 7215
rect 15865 7165 15915 7215
rect 15965 7165 16015 7215
rect 16065 7165 16115 7215
rect 16165 7165 16210 7215
rect 16260 7165 16305 7215
rect 16355 7165 16425 7215
rect 16475 7165 16520 7215
rect 16570 7165 16615 7215
rect 16665 7165 16715 7215
rect 16765 7165 16815 7215
rect 16865 7165 16915 7215
rect 16965 7165 17010 7215
rect 17060 7165 17105 7215
rect 17155 7165 17225 7215
rect 17275 7165 17320 7215
rect 17370 7165 17415 7215
rect 17465 7165 17515 7215
rect 17565 7165 17615 7215
rect 17665 7165 17715 7215
rect 17765 7165 17810 7215
rect 17860 7165 17905 7215
rect 17955 7165 20720 7215
rect 14790 7125 20720 7165
rect 14790 7075 14825 7125
rect 14875 7075 14920 7125
rect 14970 7075 15015 7125
rect 15065 7075 15115 7125
rect 15165 7075 15215 7125
rect 15265 7075 15315 7125
rect 15365 7075 15410 7125
rect 15460 7075 15505 7125
rect 15555 7075 15625 7125
rect 15675 7075 15720 7125
rect 15770 7075 15815 7125
rect 15865 7075 15915 7125
rect 15965 7075 16015 7125
rect 16065 7075 16115 7125
rect 16165 7075 16210 7125
rect 16260 7075 16305 7125
rect 16355 7075 16425 7125
rect 16475 7075 16520 7125
rect 16570 7075 16615 7125
rect 16665 7075 16715 7125
rect 16765 7075 16815 7125
rect 16865 7075 16915 7125
rect 16965 7075 17010 7125
rect 17060 7075 17105 7125
rect 17155 7075 17225 7125
rect 17275 7075 17320 7125
rect 17370 7075 17415 7125
rect 17465 7075 17515 7125
rect 17565 7075 17615 7125
rect 17665 7075 17715 7125
rect 17765 7075 17810 7125
rect 17860 7075 17905 7125
rect 17955 7075 20720 7125
rect 14790 7025 20720 7075
rect 14790 6975 14825 7025
rect 14875 6975 14920 7025
rect 14970 6975 15015 7025
rect 15065 6975 15115 7025
rect 15165 6975 15215 7025
rect 15265 6975 15315 7025
rect 15365 6975 15410 7025
rect 15460 6975 15505 7025
rect 15555 6975 15625 7025
rect 15675 6975 15720 7025
rect 15770 6975 15815 7025
rect 15865 6975 15915 7025
rect 15965 6975 16015 7025
rect 16065 6975 16115 7025
rect 16165 6975 16210 7025
rect 16260 6975 16305 7025
rect 16355 6975 16425 7025
rect 16475 6975 16520 7025
rect 16570 6975 16615 7025
rect 16665 6975 16715 7025
rect 16765 6975 16815 7025
rect 16865 6975 16915 7025
rect 16965 6975 17010 7025
rect 17060 6975 17105 7025
rect 17155 6975 17225 7025
rect 17275 6975 17320 7025
rect 17370 6975 17415 7025
rect 17465 6975 17515 7025
rect 17565 6975 17615 7025
rect 17665 6975 17715 7025
rect 17765 6975 17810 7025
rect 17860 6975 17905 7025
rect 17955 6975 20720 7025
rect -1675 6900 9100 6925
rect -1675 6885 -80 6900
rect -4840 6860 -80 6885
rect -40 6860 270 6900
rect 310 6860 620 6900
rect 660 6860 1320 6900
rect 1360 6860 1670 6900
rect 1710 6860 2385 6900
rect 2425 6860 3235 6900
rect 3275 6860 5645 6900
rect 5685 6860 6300 6900
rect 6340 6860 6590 6900
rect 6630 6860 7270 6900
rect 7310 6860 7620 6900
rect 7660 6860 8320 6900
rect 8360 6860 8670 6900
rect 8710 6860 9020 6900
rect 9060 6860 9100 6900
rect 9630 6940 14580 6945
rect 9630 6900 9635 6940
rect 9675 6900 9985 6940
rect 10025 6900 10335 6940
rect 10375 6900 10685 6940
rect 10725 6900 11035 6940
rect 11075 6900 11385 6940
rect 11425 6900 11735 6940
rect 11775 6900 12085 6940
rect 12125 6900 12435 6940
rect 12475 6900 12785 6940
rect 12825 6900 13135 6940
rect 13175 6900 13485 6940
rect 13525 6900 13835 6940
rect 13875 6900 14185 6940
rect 14225 6900 14535 6940
rect 14575 6900 14580 6940
rect 9630 6895 14580 6900
rect 14790 6935 20720 6975
rect -4840 6840 9100 6860
rect -4840 6815 -80 6840
rect -4840 6765 -4805 6815
rect -4755 6765 -4710 6815
rect -4660 6765 -4615 6815
rect -4565 6765 -4515 6815
rect -4465 6765 -4415 6815
rect -4365 6765 -4315 6815
rect -4265 6765 -4220 6815
rect -4170 6765 -4125 6815
rect -4075 6765 -4005 6815
rect -3955 6765 -3910 6815
rect -3860 6765 -3815 6815
rect -3765 6765 -3715 6815
rect -3665 6765 -3615 6815
rect -3565 6765 -3515 6815
rect -3465 6765 -3420 6815
rect -3370 6765 -3325 6815
rect -3275 6765 -3205 6815
rect -3155 6765 -3110 6815
rect -3060 6765 -3015 6815
rect -2965 6765 -2915 6815
rect -2865 6765 -2815 6815
rect -2765 6765 -2715 6815
rect -2665 6765 -2620 6815
rect -2570 6765 -2525 6815
rect -2475 6765 -2405 6815
rect -2355 6765 -2310 6815
rect -2260 6765 -2215 6815
rect -2165 6765 -2115 6815
rect -2065 6765 -2015 6815
rect -1965 6765 -1915 6815
rect -1865 6765 -1820 6815
rect -1770 6765 -1725 6815
rect -1675 6800 -80 6815
rect -40 6800 270 6840
rect 310 6800 620 6840
rect 660 6800 1320 6840
rect 1360 6800 1670 6840
rect 1710 6800 2385 6840
rect 2425 6800 3235 6840
rect 3275 6800 5645 6840
rect 5685 6800 6300 6840
rect 6340 6800 6590 6840
rect 6630 6800 7270 6840
rect 7310 6800 7620 6840
rect 7660 6800 8320 6840
rect 8360 6800 8670 6840
rect 8710 6800 9020 6840
rect 9060 6800 9100 6840
rect -1675 6775 9100 6800
rect -1675 6765 -80 6775
rect -4840 6735 -80 6765
rect -40 6735 270 6775
rect 310 6735 620 6775
rect 660 6735 1320 6775
rect 1360 6735 1670 6775
rect 1710 6735 2385 6775
rect 2425 6735 3235 6775
rect 3275 6735 5645 6775
rect 5685 6735 6300 6775
rect 6340 6735 6590 6775
rect 6630 6735 7270 6775
rect 7310 6735 7620 6775
rect 7660 6735 8320 6775
rect 8360 6735 8670 6775
rect 8710 6735 9020 6775
rect 9060 6735 9100 6775
rect -4840 6725 9100 6735
rect -4840 6675 -4805 6725
rect -4755 6675 -4710 6725
rect -4660 6675 -4615 6725
rect -4565 6675 -4515 6725
rect -4465 6675 -4415 6725
rect -4365 6675 -4315 6725
rect -4265 6675 -4220 6725
rect -4170 6675 -4125 6725
rect -4075 6675 -4005 6725
rect -3955 6675 -3910 6725
rect -3860 6675 -3815 6725
rect -3765 6675 -3715 6725
rect -3665 6675 -3615 6725
rect -3565 6675 -3515 6725
rect -3465 6675 -3420 6725
rect -3370 6675 -3325 6725
rect -3275 6675 -3205 6725
rect -3155 6675 -3110 6725
rect -3060 6675 -3015 6725
rect -2965 6675 -2915 6725
rect -2865 6675 -2815 6725
rect -2765 6675 -2715 6725
rect -2665 6675 -2620 6725
rect -2570 6675 -2525 6725
rect -2475 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6705 9100 6725
rect -1675 6675 -80 6705
rect -4840 6665 -80 6675
rect -40 6665 270 6705
rect 310 6665 620 6705
rect 660 6665 1320 6705
rect 1360 6665 1670 6705
rect 1710 6665 2385 6705
rect 2425 6665 3235 6705
rect 3275 6665 5645 6705
rect 5685 6665 6300 6705
rect 6340 6665 6590 6705
rect 6630 6665 7270 6705
rect 7310 6665 7620 6705
rect 7660 6665 8320 6705
rect 8360 6665 8670 6705
rect 8710 6665 9020 6705
rect 9060 6665 9100 6705
rect -4840 6635 9100 6665
rect -4840 6625 -80 6635
rect -4840 6575 -4805 6625
rect -4755 6575 -4710 6625
rect -4660 6575 -4615 6625
rect -4565 6575 -4515 6625
rect -4465 6575 -4415 6625
rect -4365 6575 -4315 6625
rect -4265 6575 -4220 6625
rect -4170 6575 -4125 6625
rect -4075 6575 -4005 6625
rect -3955 6575 -3910 6625
rect -3860 6575 -3815 6625
rect -3765 6575 -3715 6625
rect -3665 6575 -3615 6625
rect -3565 6575 -3515 6625
rect -3465 6575 -3420 6625
rect -3370 6575 -3325 6625
rect -3275 6575 -3205 6625
rect -3155 6575 -3110 6625
rect -3060 6575 -3015 6625
rect -2965 6575 -2915 6625
rect -2865 6575 -2815 6625
rect -2765 6575 -2715 6625
rect -2665 6575 -2620 6625
rect -2570 6575 -2525 6625
rect -2475 6575 -2405 6625
rect -2355 6575 -2310 6625
rect -2260 6575 -2215 6625
rect -2165 6575 -2115 6625
rect -2065 6575 -2015 6625
rect -1965 6575 -1915 6625
rect -1865 6575 -1820 6625
rect -1770 6575 -1725 6625
rect -1675 6595 -80 6625
rect -40 6595 270 6635
rect 310 6595 620 6635
rect 660 6595 1320 6635
rect 1360 6595 1670 6635
rect 1710 6595 2385 6635
rect 2425 6595 3235 6635
rect 3275 6595 5645 6635
rect 5685 6595 6300 6635
rect 6340 6595 6590 6635
rect 6630 6595 7270 6635
rect 7310 6595 7620 6635
rect 7660 6595 8320 6635
rect 8360 6595 8670 6635
rect 8710 6595 9020 6635
rect 9060 6595 9100 6635
rect 12080 6595 12130 6895
rect 14790 6885 14825 6935
rect 14875 6885 14920 6935
rect 14970 6885 15015 6935
rect 15065 6885 15115 6935
rect 15165 6885 15215 6935
rect 15265 6885 15315 6935
rect 15365 6885 15410 6935
rect 15460 6885 15505 6935
rect 15555 6885 15625 6935
rect 15675 6885 15720 6935
rect 15770 6885 15815 6935
rect 15865 6885 15915 6935
rect 15965 6885 16015 6935
rect 16065 6885 16115 6935
rect 16165 6885 16210 6935
rect 16260 6885 16305 6935
rect 16355 6885 16425 6935
rect 16475 6885 16520 6935
rect 16570 6885 16615 6935
rect 16665 6885 16715 6935
rect 16765 6885 16815 6935
rect 16865 6885 16915 6935
rect 16965 6885 17010 6935
rect 17060 6885 17105 6935
rect 17155 6885 17225 6935
rect 17275 6885 17320 6935
rect 17370 6885 17415 6935
rect 17465 6885 17515 6935
rect 17565 6885 17615 6935
rect 17665 6885 17715 6935
rect 17765 6885 17810 6935
rect 17860 6885 17905 6935
rect 17955 6885 20720 6935
rect 14790 6815 20720 6885
rect 14790 6765 14825 6815
rect 14875 6765 14920 6815
rect 14970 6765 15015 6815
rect 15065 6765 15115 6815
rect 15165 6765 15215 6815
rect 15265 6765 15315 6815
rect 15365 6765 15410 6815
rect 15460 6765 15505 6815
rect 15555 6765 15625 6815
rect 15675 6765 15720 6815
rect 15770 6765 15815 6815
rect 15865 6765 15915 6815
rect 15965 6765 16015 6815
rect 16065 6765 16115 6815
rect 16165 6765 16210 6815
rect 16260 6765 16305 6815
rect 16355 6765 16425 6815
rect 16475 6765 16520 6815
rect 16570 6765 16615 6815
rect 16665 6765 16715 6815
rect 16765 6765 16815 6815
rect 16865 6765 16915 6815
rect 16965 6765 17010 6815
rect 17060 6765 17105 6815
rect 17155 6765 17225 6815
rect 17275 6765 17320 6815
rect 17370 6765 17415 6815
rect 17465 6765 17515 6815
rect 17565 6765 17615 6815
rect 17665 6765 17715 6815
rect 17765 6765 17810 6815
rect 17860 6765 17905 6815
rect 17955 6765 20720 6815
rect 14790 6725 20720 6765
rect 14790 6675 14825 6725
rect 14875 6675 14920 6725
rect 14970 6675 15015 6725
rect 15065 6675 15115 6725
rect 15165 6675 15215 6725
rect 15265 6675 15315 6725
rect 15365 6675 15410 6725
rect 15460 6675 15505 6725
rect 15555 6675 15625 6725
rect 15675 6675 15720 6725
rect 15770 6675 15815 6725
rect 15865 6675 15915 6725
rect 15965 6675 16015 6725
rect 16065 6675 16115 6725
rect 16165 6675 16210 6725
rect 16260 6675 16305 6725
rect 16355 6675 16425 6725
rect 16475 6675 16520 6725
rect 16570 6675 16615 6725
rect 16665 6675 16715 6725
rect 16765 6675 16815 6725
rect 16865 6675 16915 6725
rect 16965 6675 17010 6725
rect 17060 6675 17105 6725
rect 17155 6675 17225 6725
rect 17275 6675 17320 6725
rect 17370 6675 17415 6725
rect 17465 6675 17515 6725
rect 17565 6675 17615 6725
rect 17665 6675 17715 6725
rect 17765 6675 17810 6725
rect 17860 6675 17905 6725
rect 17955 6675 20720 6725
rect 14790 6625 20720 6675
rect -1675 6590 14580 6595
rect -1675 6575 9635 6590
rect -4840 6565 9635 6575
rect -4840 6535 -80 6565
rect -4840 6485 -4805 6535
rect -4755 6485 -4710 6535
rect -4660 6485 -4615 6535
rect -4565 6485 -4515 6535
rect -4465 6485 -4415 6535
rect -4365 6485 -4315 6535
rect -4265 6485 -4220 6535
rect -4170 6485 -4125 6535
rect -4075 6485 -4005 6535
rect -3955 6485 -3910 6535
rect -3860 6485 -3815 6535
rect -3765 6485 -3715 6535
rect -3665 6485 -3615 6535
rect -3565 6485 -3515 6535
rect -3465 6485 -3420 6535
rect -3370 6485 -3325 6535
rect -3275 6485 -3205 6535
rect -3155 6485 -3110 6535
rect -3060 6485 -3015 6535
rect -2965 6485 -2915 6535
rect -2865 6485 -2815 6535
rect -2765 6485 -2715 6535
rect -2665 6485 -2620 6535
rect -2570 6485 -2525 6535
rect -2475 6485 -2405 6535
rect -2355 6485 -2310 6535
rect -2260 6485 -2215 6535
rect -2165 6485 -2115 6535
rect -2065 6485 -2015 6535
rect -1965 6485 -1915 6535
rect -1865 6485 -1820 6535
rect -1770 6485 -1725 6535
rect -1675 6525 -80 6535
rect -40 6525 270 6565
rect 310 6525 620 6565
rect 660 6525 1320 6565
rect 1360 6525 1670 6565
rect 1710 6525 2385 6565
rect 2425 6525 3235 6565
rect 3275 6525 5645 6565
rect 5685 6525 6300 6565
rect 6340 6525 6590 6565
rect 6630 6525 7270 6565
rect 7310 6525 7620 6565
rect 7660 6525 8320 6565
rect 8360 6525 8670 6565
rect 8710 6525 9020 6565
rect 9060 6550 9635 6565
rect 9675 6550 9985 6590
rect 10025 6550 10335 6590
rect 10375 6550 10685 6590
rect 10725 6550 11035 6590
rect 11075 6550 11385 6590
rect 11425 6550 11735 6590
rect 11775 6550 12085 6590
rect 12125 6550 12435 6590
rect 12475 6550 12785 6590
rect 12825 6550 13135 6590
rect 13175 6550 13485 6590
rect 13525 6550 13835 6590
rect 13875 6550 14185 6590
rect 14225 6550 14535 6590
rect 14575 6550 14580 6590
rect 9060 6545 14580 6550
rect 14790 6575 14825 6625
rect 14875 6575 14920 6625
rect 14970 6575 15015 6625
rect 15065 6575 15115 6625
rect 15165 6575 15215 6625
rect 15265 6575 15315 6625
rect 15365 6575 15410 6625
rect 15460 6575 15505 6625
rect 15555 6575 15625 6625
rect 15675 6575 15720 6625
rect 15770 6575 15815 6625
rect 15865 6575 15915 6625
rect 15965 6575 16015 6625
rect 16065 6575 16115 6625
rect 16165 6575 16210 6625
rect 16260 6575 16305 6625
rect 16355 6575 16425 6625
rect 16475 6575 16520 6625
rect 16570 6575 16615 6625
rect 16665 6575 16715 6625
rect 16765 6575 16815 6625
rect 16865 6575 16915 6625
rect 16965 6575 17010 6625
rect 17060 6575 17105 6625
rect 17155 6575 17225 6625
rect 17275 6575 17320 6625
rect 17370 6575 17415 6625
rect 17465 6575 17515 6625
rect 17565 6575 17615 6625
rect 17665 6575 17715 6625
rect 17765 6575 17810 6625
rect 17860 6575 17905 6625
rect 17955 6575 20720 6625
rect 9060 6525 9100 6545
rect -1675 6500 9100 6525
rect -1675 6485 -80 6500
rect -4840 6460 -80 6485
rect -40 6460 270 6500
rect 310 6460 620 6500
rect 660 6460 1320 6500
rect 1360 6460 1670 6500
rect 1710 6460 2385 6500
rect 2425 6460 3235 6500
rect 3275 6460 5645 6500
rect 5685 6460 6300 6500
rect 6340 6460 6590 6500
rect 6630 6460 7270 6500
rect 7310 6460 7620 6500
rect 7660 6460 8320 6500
rect 8360 6460 8670 6500
rect 8710 6460 9020 6500
rect 9060 6460 9100 6500
rect -4840 6450 9100 6460
rect 14790 6535 20720 6575
rect 14790 6485 14825 6535
rect 14875 6485 14920 6535
rect 14970 6485 15015 6535
rect 15065 6485 15115 6535
rect 15165 6485 15215 6535
rect 15265 6485 15315 6535
rect 15365 6485 15410 6535
rect 15460 6485 15505 6535
rect 15555 6485 15625 6535
rect 15675 6485 15720 6535
rect 15770 6485 15815 6535
rect 15865 6485 15915 6535
rect 15965 6485 16015 6535
rect 16065 6485 16115 6535
rect 16165 6485 16210 6535
rect 16260 6485 16305 6535
rect 16355 6485 16425 6535
rect 16475 6485 16520 6535
rect 16570 6485 16615 6535
rect 16665 6485 16715 6535
rect 16765 6485 16815 6535
rect 16865 6485 16915 6535
rect 16965 6485 17010 6535
rect 17060 6485 17105 6535
rect 17155 6485 17225 6535
rect 17275 6485 17320 6535
rect 17370 6485 17415 6535
rect 17465 6485 17515 6535
rect 17565 6485 17615 6535
rect 17665 6485 17715 6535
rect 17765 6485 17810 6535
rect 17860 6485 17905 6535
rect 17955 6485 20720 6535
rect 14790 6450 20720 6485
rect 1500 1370 1510 1380
rect -120 -1300 17990 -1290
rect -120 -1340 -80 -1300
rect -40 -1340 270 -1300
rect 310 -1340 620 -1300
rect 660 -1340 970 -1300
rect 1010 -1340 1320 -1300
rect 1360 -1340 1670 -1300
rect 1710 -1340 2020 -1300
rect 2060 -1340 2370 -1300
rect 2410 -1340 2720 -1300
rect 2760 -1340 3070 -1300
rect 3110 -1340 3420 -1300
rect 3460 -1340 3770 -1300
rect 3810 -1340 4120 -1300
rect 4160 -1340 4470 -1300
rect 4510 -1340 4820 -1300
rect 4860 -1340 5170 -1300
rect 5210 -1340 5520 -1300
rect 5560 -1340 5870 -1300
rect 5910 -1340 6220 -1300
rect 6260 -1340 6570 -1300
rect 6610 -1340 6920 -1300
rect 6960 -1340 7270 -1300
rect 7310 -1340 7620 -1300
rect 7660 -1340 7970 -1300
rect 8010 -1340 8320 -1300
rect 8360 -1340 8670 -1300
rect 8710 -1325 17990 -1300
rect 8710 -1340 14825 -1325
rect -120 -1365 14825 -1340
rect -120 -1405 -80 -1365
rect -40 -1405 270 -1365
rect 310 -1405 620 -1365
rect 660 -1405 970 -1365
rect 1010 -1405 1320 -1365
rect 1360 -1405 1670 -1365
rect 1710 -1405 2020 -1365
rect 2060 -1405 2370 -1365
rect 2410 -1405 2720 -1365
rect 2760 -1405 3070 -1365
rect 3110 -1405 3420 -1365
rect 3460 -1405 3770 -1365
rect 3810 -1405 4120 -1365
rect 4160 -1405 4470 -1365
rect 4510 -1405 4820 -1365
rect 4860 -1405 5170 -1365
rect 5210 -1405 5520 -1365
rect 5560 -1405 5870 -1365
rect 5910 -1405 6220 -1365
rect 6260 -1405 6570 -1365
rect 6610 -1405 6920 -1365
rect 6960 -1405 7270 -1365
rect 7310 -1405 7620 -1365
rect 7660 -1405 7970 -1365
rect 8010 -1405 8320 -1365
rect 8360 -1405 8670 -1365
rect 8710 -1375 14825 -1365
rect 14875 -1375 14920 -1325
rect 14970 -1375 15015 -1325
rect 15065 -1375 15115 -1325
rect 15165 -1375 15215 -1325
rect 15265 -1375 15315 -1325
rect 15365 -1375 15410 -1325
rect 15460 -1375 15505 -1325
rect 15555 -1375 15625 -1325
rect 15675 -1375 15720 -1325
rect 15770 -1375 15815 -1325
rect 15865 -1375 15915 -1325
rect 15965 -1375 16015 -1325
rect 16065 -1375 16115 -1325
rect 16165 -1375 16210 -1325
rect 16260 -1375 16305 -1325
rect 16355 -1375 16425 -1325
rect 16475 -1375 16520 -1325
rect 16570 -1375 16615 -1325
rect 16665 -1375 16715 -1325
rect 16765 -1375 16815 -1325
rect 16865 -1375 16915 -1325
rect 16965 -1375 17010 -1325
rect 17060 -1375 17105 -1325
rect 17155 -1375 17225 -1325
rect 17275 -1375 17320 -1325
rect 17370 -1375 17415 -1325
rect 17465 -1375 17515 -1325
rect 17565 -1375 17615 -1325
rect 17665 -1375 17715 -1325
rect 17765 -1375 17810 -1325
rect 17860 -1375 17905 -1325
rect 17955 -1375 17990 -1325
rect 8710 -1405 17990 -1375
rect -120 -1415 17990 -1405
rect -120 -1435 14825 -1415
rect -120 -1475 -80 -1435
rect -40 -1475 270 -1435
rect 310 -1475 620 -1435
rect 660 -1475 970 -1435
rect 1010 -1475 1320 -1435
rect 1360 -1475 1670 -1435
rect 1710 -1475 2020 -1435
rect 2060 -1475 2370 -1435
rect 2410 -1475 2720 -1435
rect 2760 -1475 3070 -1435
rect 3110 -1475 3420 -1435
rect 3460 -1475 3770 -1435
rect 3810 -1475 4120 -1435
rect 4160 -1475 4470 -1435
rect 4510 -1475 4820 -1435
rect 4860 -1475 5170 -1435
rect 5210 -1475 5520 -1435
rect 5560 -1475 5870 -1435
rect 5910 -1475 6220 -1435
rect 6260 -1475 6570 -1435
rect 6610 -1475 6920 -1435
rect 6960 -1475 7270 -1435
rect 7310 -1475 7620 -1435
rect 7660 -1475 7970 -1435
rect 8010 -1475 8320 -1435
rect 8360 -1475 8670 -1435
rect 8710 -1465 14825 -1435
rect 14875 -1465 14920 -1415
rect 14970 -1465 15015 -1415
rect 15065 -1465 15115 -1415
rect 15165 -1465 15215 -1415
rect 15265 -1465 15315 -1415
rect 15365 -1465 15410 -1415
rect 15460 -1465 15505 -1415
rect 15555 -1465 15625 -1415
rect 15675 -1465 15720 -1415
rect 15770 -1465 15815 -1415
rect 15865 -1465 15915 -1415
rect 15965 -1465 16015 -1415
rect 16065 -1465 16115 -1415
rect 16165 -1465 16210 -1415
rect 16260 -1465 16305 -1415
rect 16355 -1465 16425 -1415
rect 16475 -1465 16520 -1415
rect 16570 -1465 16615 -1415
rect 16665 -1465 16715 -1415
rect 16765 -1465 16815 -1415
rect 16865 -1465 16915 -1415
rect 16965 -1465 17010 -1415
rect 17060 -1465 17105 -1415
rect 17155 -1465 17225 -1415
rect 17275 -1465 17320 -1415
rect 17370 -1465 17415 -1415
rect 17465 -1465 17515 -1415
rect 17565 -1465 17615 -1415
rect 17665 -1465 17715 -1415
rect 17765 -1465 17810 -1415
rect 17860 -1465 17905 -1415
rect 17955 -1465 17990 -1415
rect 8710 -1475 17990 -1465
rect -120 -1505 17990 -1475
rect -120 -1545 -80 -1505
rect -40 -1545 270 -1505
rect 310 -1545 620 -1505
rect 660 -1545 970 -1505
rect 1010 -1545 1320 -1505
rect 1360 -1545 1670 -1505
rect 1710 -1545 2020 -1505
rect 2060 -1545 2370 -1505
rect 2410 -1545 2720 -1505
rect 2760 -1545 3070 -1505
rect 3110 -1545 3420 -1505
rect 3460 -1545 3770 -1505
rect 3810 -1545 4120 -1505
rect 4160 -1545 4470 -1505
rect 4510 -1545 4820 -1505
rect 4860 -1545 5170 -1505
rect 5210 -1545 5520 -1505
rect 5560 -1545 5870 -1505
rect 5910 -1545 6220 -1505
rect 6260 -1545 6570 -1505
rect 6610 -1545 6920 -1505
rect 6960 -1545 7270 -1505
rect 7310 -1545 7620 -1505
rect 7660 -1545 7970 -1505
rect 8010 -1545 8320 -1505
rect 8360 -1545 8670 -1505
rect 8710 -1515 17990 -1505
rect 8710 -1545 14825 -1515
rect -120 -1565 14825 -1545
rect 14875 -1565 14920 -1515
rect 14970 -1565 15015 -1515
rect 15065 -1565 15115 -1515
rect 15165 -1565 15215 -1515
rect 15265 -1565 15315 -1515
rect 15365 -1565 15410 -1515
rect 15460 -1565 15505 -1515
rect 15555 -1565 15625 -1515
rect 15675 -1565 15720 -1515
rect 15770 -1565 15815 -1515
rect 15865 -1565 15915 -1515
rect 15965 -1565 16015 -1515
rect 16065 -1565 16115 -1515
rect 16165 -1565 16210 -1515
rect 16260 -1565 16305 -1515
rect 16355 -1565 16425 -1515
rect 16475 -1565 16520 -1515
rect 16570 -1565 16615 -1515
rect 16665 -1565 16715 -1515
rect 16765 -1565 16815 -1515
rect 16865 -1565 16915 -1515
rect 16965 -1565 17010 -1515
rect 17060 -1565 17105 -1515
rect 17155 -1565 17225 -1515
rect 17275 -1565 17320 -1515
rect 17370 -1565 17415 -1515
rect 17465 -1565 17515 -1515
rect 17565 -1565 17615 -1515
rect 17665 -1565 17715 -1515
rect 17765 -1565 17810 -1515
rect 17860 -1565 17905 -1515
rect 17955 -1565 17990 -1515
rect -120 -1575 17990 -1565
rect -120 -1615 -80 -1575
rect -40 -1615 270 -1575
rect 310 -1615 620 -1575
rect 660 -1615 970 -1575
rect 1010 -1615 1320 -1575
rect 1360 -1615 1670 -1575
rect 1710 -1615 2020 -1575
rect 2060 -1615 2370 -1575
rect 2410 -1615 2720 -1575
rect 2760 -1615 3070 -1575
rect 3110 -1615 3420 -1575
rect 3460 -1615 3770 -1575
rect 3810 -1615 4120 -1575
rect 4160 -1615 4470 -1575
rect 4510 -1615 4820 -1575
rect 4860 -1615 5170 -1575
rect 5210 -1615 5520 -1575
rect 5560 -1615 5870 -1575
rect 5910 -1615 6220 -1575
rect 6260 -1615 6570 -1575
rect 6610 -1615 6920 -1575
rect 6960 -1615 7270 -1575
rect 7310 -1615 7620 -1575
rect 7660 -1615 7970 -1575
rect 8010 -1615 8320 -1575
rect 8360 -1615 8670 -1575
rect 8710 -1605 17990 -1575
rect 8710 -1615 14825 -1605
rect -120 -1640 14825 -1615
rect -120 -1680 -80 -1640
rect -40 -1680 270 -1640
rect 310 -1680 620 -1640
rect 660 -1680 970 -1640
rect 1010 -1680 1320 -1640
rect 1360 -1680 1670 -1640
rect 1710 -1680 2020 -1640
rect 2060 -1680 2370 -1640
rect 2410 -1680 2720 -1640
rect 2760 -1680 3070 -1640
rect 3110 -1680 3420 -1640
rect 3460 -1680 3770 -1640
rect 3810 -1680 4120 -1640
rect 4160 -1680 4470 -1640
rect 4510 -1680 4820 -1640
rect 4860 -1680 5170 -1640
rect 5210 -1680 5520 -1640
rect 5560 -1680 5870 -1640
rect 5910 -1680 6220 -1640
rect 6260 -1680 6570 -1640
rect 6610 -1680 6920 -1640
rect 6960 -1680 7270 -1640
rect 7310 -1680 7620 -1640
rect 7660 -1680 7970 -1640
rect 8010 -1680 8320 -1640
rect 8360 -1680 8670 -1640
rect 8710 -1655 14825 -1640
rect 14875 -1655 14920 -1605
rect 14970 -1655 15015 -1605
rect 15065 -1655 15115 -1605
rect 15165 -1655 15215 -1605
rect 15265 -1655 15315 -1605
rect 15365 -1655 15410 -1605
rect 15460 -1655 15505 -1605
rect 15555 -1655 15625 -1605
rect 15675 -1655 15720 -1605
rect 15770 -1655 15815 -1605
rect 15865 -1655 15915 -1605
rect 15965 -1655 16015 -1605
rect 16065 -1655 16115 -1605
rect 16165 -1655 16210 -1605
rect 16260 -1655 16305 -1605
rect 16355 -1655 16425 -1605
rect 16475 -1655 16520 -1605
rect 16570 -1655 16615 -1605
rect 16665 -1655 16715 -1605
rect 16765 -1655 16815 -1605
rect 16865 -1655 16915 -1605
rect 16965 -1655 17010 -1605
rect 17060 -1655 17105 -1605
rect 17155 -1655 17225 -1605
rect 17275 -1655 17320 -1605
rect 17370 -1655 17415 -1605
rect 17465 -1655 17515 -1605
rect 17565 -1655 17615 -1605
rect 17665 -1655 17715 -1605
rect 17765 -1655 17810 -1605
rect 17860 -1655 17905 -1605
rect 17955 -1655 17990 -1605
rect 8710 -1680 17990 -1655
rect -120 -1700 17990 -1680
rect -120 -1740 -80 -1700
rect -40 -1740 270 -1700
rect 310 -1740 620 -1700
rect 660 -1740 970 -1700
rect 1010 -1740 1320 -1700
rect 1360 -1740 1670 -1700
rect 1710 -1740 2020 -1700
rect 2060 -1740 2370 -1700
rect 2410 -1740 2720 -1700
rect 2760 -1740 3070 -1700
rect 3110 -1740 3420 -1700
rect 3460 -1740 3770 -1700
rect 3810 -1740 4120 -1700
rect 4160 -1740 4470 -1700
rect 4510 -1740 4820 -1700
rect 4860 -1740 5170 -1700
rect 5210 -1740 5520 -1700
rect 5560 -1740 5870 -1700
rect 5910 -1740 6220 -1700
rect 6260 -1740 6570 -1700
rect 6610 -1740 6920 -1700
rect 6960 -1740 7270 -1700
rect 7310 -1740 7620 -1700
rect 7660 -1740 7970 -1700
rect 8010 -1740 8320 -1700
rect 8360 -1740 8670 -1700
rect 8710 -1725 17990 -1700
rect 8710 -1740 14825 -1725
rect -120 -1765 14825 -1740
rect -120 -1805 -80 -1765
rect -40 -1805 270 -1765
rect 310 -1805 620 -1765
rect 660 -1805 970 -1765
rect 1010 -1805 1320 -1765
rect 1360 -1805 1670 -1765
rect 1710 -1805 2020 -1765
rect 2060 -1805 2370 -1765
rect 2410 -1805 2720 -1765
rect 2760 -1805 3070 -1765
rect 3110 -1805 3420 -1765
rect 3460 -1805 3770 -1765
rect 3810 -1805 4120 -1765
rect 4160 -1805 4470 -1765
rect 4510 -1805 4820 -1765
rect 4860 -1805 5170 -1765
rect 5210 -1805 5520 -1765
rect 5560 -1805 5870 -1765
rect 5910 -1805 6220 -1765
rect 6260 -1805 6570 -1765
rect 6610 -1805 6920 -1765
rect 6960 -1805 7270 -1765
rect 7310 -1805 7620 -1765
rect 7660 -1805 7970 -1765
rect 8010 -1805 8320 -1765
rect 8360 -1805 8670 -1765
rect 8710 -1775 14825 -1765
rect 14875 -1775 14920 -1725
rect 14970 -1775 15015 -1725
rect 15065 -1775 15115 -1725
rect 15165 -1775 15215 -1725
rect 15265 -1775 15315 -1725
rect 15365 -1775 15410 -1725
rect 15460 -1775 15505 -1725
rect 15555 -1775 15625 -1725
rect 15675 -1775 15720 -1725
rect 15770 -1775 15815 -1725
rect 15865 -1775 15915 -1725
rect 15965 -1775 16015 -1725
rect 16065 -1775 16115 -1725
rect 16165 -1775 16210 -1725
rect 16260 -1775 16305 -1725
rect 16355 -1775 16425 -1725
rect 16475 -1775 16520 -1725
rect 16570 -1775 16615 -1725
rect 16665 -1775 16715 -1725
rect 16765 -1775 16815 -1725
rect 16865 -1775 16915 -1725
rect 16965 -1775 17010 -1725
rect 17060 -1775 17105 -1725
rect 17155 -1775 17225 -1725
rect 17275 -1775 17320 -1725
rect 17370 -1775 17415 -1725
rect 17465 -1775 17515 -1725
rect 17565 -1775 17615 -1725
rect 17665 -1775 17715 -1725
rect 17765 -1775 17810 -1725
rect 17860 -1775 17905 -1725
rect 17955 -1775 17990 -1725
rect 8710 -1805 17990 -1775
rect -120 -1815 17990 -1805
rect -120 -1835 14825 -1815
rect -120 -1875 -80 -1835
rect -40 -1875 270 -1835
rect 310 -1875 620 -1835
rect 660 -1875 970 -1835
rect 1010 -1875 1320 -1835
rect 1360 -1875 1670 -1835
rect 1710 -1875 2020 -1835
rect 2060 -1875 2370 -1835
rect 2410 -1875 2720 -1835
rect 2760 -1875 3070 -1835
rect 3110 -1875 3420 -1835
rect 3460 -1875 3770 -1835
rect 3810 -1875 4120 -1835
rect 4160 -1875 4470 -1835
rect 4510 -1875 4820 -1835
rect 4860 -1875 5170 -1835
rect 5210 -1875 5520 -1835
rect 5560 -1875 5870 -1835
rect 5910 -1875 6220 -1835
rect 6260 -1875 6570 -1835
rect 6610 -1875 6920 -1835
rect 6960 -1875 7270 -1835
rect 7310 -1875 7620 -1835
rect 7660 -1875 7970 -1835
rect 8010 -1875 8320 -1835
rect 8360 -1875 8670 -1835
rect 8710 -1865 14825 -1835
rect 14875 -1865 14920 -1815
rect 14970 -1865 15015 -1815
rect 15065 -1865 15115 -1815
rect 15165 -1865 15215 -1815
rect 15265 -1865 15315 -1815
rect 15365 -1865 15410 -1815
rect 15460 -1865 15505 -1815
rect 15555 -1865 15625 -1815
rect 15675 -1865 15720 -1815
rect 15770 -1865 15815 -1815
rect 15865 -1865 15915 -1815
rect 15965 -1865 16015 -1815
rect 16065 -1865 16115 -1815
rect 16165 -1865 16210 -1815
rect 16260 -1865 16305 -1815
rect 16355 -1865 16425 -1815
rect 16475 -1865 16520 -1815
rect 16570 -1865 16615 -1815
rect 16665 -1865 16715 -1815
rect 16765 -1865 16815 -1815
rect 16865 -1865 16915 -1815
rect 16965 -1865 17010 -1815
rect 17060 -1865 17105 -1815
rect 17155 -1865 17225 -1815
rect 17275 -1865 17320 -1815
rect 17370 -1865 17415 -1815
rect 17465 -1865 17515 -1815
rect 17565 -1865 17615 -1815
rect 17665 -1865 17715 -1815
rect 17765 -1865 17810 -1815
rect 17860 -1865 17905 -1815
rect 17955 -1865 17990 -1815
rect 8710 -1875 17990 -1865
rect -120 -1905 17990 -1875
rect -120 -1945 -80 -1905
rect -40 -1945 270 -1905
rect 310 -1945 620 -1905
rect 660 -1945 970 -1905
rect 1010 -1945 1320 -1905
rect 1360 -1945 1670 -1905
rect 1710 -1945 2020 -1905
rect 2060 -1945 2370 -1905
rect 2410 -1945 2720 -1905
rect 2760 -1945 3070 -1905
rect 3110 -1945 3420 -1905
rect 3460 -1945 3770 -1905
rect 3810 -1945 4120 -1905
rect 4160 -1945 4470 -1905
rect 4510 -1945 4820 -1905
rect 4860 -1945 5170 -1905
rect 5210 -1945 5520 -1905
rect 5560 -1945 5870 -1905
rect 5910 -1945 6220 -1905
rect 6260 -1945 6570 -1905
rect 6610 -1945 6920 -1905
rect 6960 -1945 7270 -1905
rect 7310 -1945 7620 -1905
rect 7660 -1945 7970 -1905
rect 8010 -1945 8320 -1905
rect 8360 -1945 8670 -1905
rect 8710 -1915 17990 -1905
rect 8710 -1945 14825 -1915
rect -120 -1965 14825 -1945
rect 14875 -1965 14920 -1915
rect 14970 -1965 15015 -1915
rect 15065 -1965 15115 -1915
rect 15165 -1965 15215 -1915
rect 15265 -1965 15315 -1915
rect 15365 -1965 15410 -1915
rect 15460 -1965 15505 -1915
rect 15555 -1965 15625 -1915
rect 15675 -1965 15720 -1915
rect 15770 -1965 15815 -1915
rect 15865 -1965 15915 -1915
rect 15965 -1965 16015 -1915
rect 16065 -1965 16115 -1915
rect 16165 -1965 16210 -1915
rect 16260 -1965 16305 -1915
rect 16355 -1965 16425 -1915
rect 16475 -1965 16520 -1915
rect 16570 -1965 16615 -1915
rect 16665 -1965 16715 -1915
rect 16765 -1965 16815 -1915
rect 16865 -1965 16915 -1915
rect 16965 -1965 17010 -1915
rect 17060 -1965 17105 -1915
rect 17155 -1965 17225 -1915
rect 17275 -1965 17320 -1915
rect 17370 -1965 17415 -1915
rect 17465 -1965 17515 -1915
rect 17565 -1965 17615 -1915
rect 17665 -1965 17715 -1915
rect 17765 -1965 17810 -1915
rect 17860 -1965 17905 -1915
rect 17955 -1965 17990 -1915
rect -120 -1975 17990 -1965
rect -120 -2015 -80 -1975
rect -40 -2015 270 -1975
rect 310 -2015 620 -1975
rect 660 -2015 970 -1975
rect 1010 -2015 1320 -1975
rect 1360 -2015 1670 -1975
rect 1710 -2015 2020 -1975
rect 2060 -2015 2370 -1975
rect 2410 -2015 2720 -1975
rect 2760 -2015 3070 -1975
rect 3110 -2015 3420 -1975
rect 3460 -2015 3770 -1975
rect 3810 -2015 4120 -1975
rect 4160 -2015 4470 -1975
rect 4510 -2015 4820 -1975
rect 4860 -2015 5170 -1975
rect 5210 -2015 5520 -1975
rect 5560 -2015 5870 -1975
rect 5910 -2015 6220 -1975
rect 6260 -2015 6570 -1975
rect 6610 -2015 6920 -1975
rect 6960 -2015 7270 -1975
rect 7310 -2015 7620 -1975
rect 7660 -2015 7970 -1975
rect 8010 -2015 8320 -1975
rect 8360 -2015 8670 -1975
rect 8710 -2005 17990 -1975
rect 8710 -2015 14825 -2005
rect -120 -2040 14825 -2015
rect -120 -2080 -80 -2040
rect -40 -2080 270 -2040
rect 310 -2080 620 -2040
rect 660 -2080 970 -2040
rect 1010 -2080 1320 -2040
rect 1360 -2080 1670 -2040
rect 1710 -2080 2020 -2040
rect 2060 -2080 2370 -2040
rect 2410 -2080 2720 -2040
rect 2760 -2080 3070 -2040
rect 3110 -2080 3420 -2040
rect 3460 -2080 3770 -2040
rect 3810 -2080 4120 -2040
rect 4160 -2080 4470 -2040
rect 4510 -2080 4820 -2040
rect 4860 -2080 5170 -2040
rect 5210 -2080 5520 -2040
rect 5560 -2080 5870 -2040
rect 5910 -2080 6220 -2040
rect 6260 -2080 6570 -2040
rect 6610 -2080 6920 -2040
rect 6960 -2080 7270 -2040
rect 7310 -2080 7620 -2040
rect 7660 -2080 7970 -2040
rect 8010 -2080 8320 -2040
rect 8360 -2080 8670 -2040
rect 8710 -2055 14825 -2040
rect 14875 -2055 14920 -2005
rect 14970 -2055 15015 -2005
rect 15065 -2055 15115 -2005
rect 15165 -2055 15215 -2005
rect 15265 -2055 15315 -2005
rect 15365 -2055 15410 -2005
rect 15460 -2055 15505 -2005
rect 15555 -2055 15625 -2005
rect 15675 -2055 15720 -2005
rect 15770 -2055 15815 -2005
rect 15865 -2055 15915 -2005
rect 15965 -2055 16015 -2005
rect 16065 -2055 16115 -2005
rect 16165 -2055 16210 -2005
rect 16260 -2055 16305 -2005
rect 16355 -2055 16425 -2005
rect 16475 -2055 16520 -2005
rect 16570 -2055 16615 -2005
rect 16665 -2055 16715 -2005
rect 16765 -2055 16815 -2005
rect 16865 -2055 16915 -2005
rect 16965 -2055 17010 -2005
rect 17060 -2055 17105 -2005
rect 17155 -2055 17225 -2005
rect 17275 -2055 17320 -2005
rect 17370 -2055 17415 -2005
rect 17465 -2055 17515 -2005
rect 17565 -2055 17615 -2005
rect 17665 -2055 17715 -2005
rect 17765 -2055 17810 -2005
rect 17860 -2055 17905 -2005
rect 17955 -2055 17990 -2005
rect 8710 -2080 17990 -2055
rect -120 -2100 17990 -2080
rect -120 -2140 -80 -2100
rect -40 -2140 270 -2100
rect 310 -2140 620 -2100
rect 660 -2140 970 -2100
rect 1010 -2140 1320 -2100
rect 1360 -2140 1670 -2100
rect 1710 -2140 2020 -2100
rect 2060 -2140 2370 -2100
rect 2410 -2140 2720 -2100
rect 2760 -2140 3070 -2100
rect 3110 -2140 3420 -2100
rect 3460 -2140 3770 -2100
rect 3810 -2140 4120 -2100
rect 4160 -2140 4470 -2100
rect 4510 -2140 4820 -2100
rect 4860 -2140 5170 -2100
rect 5210 -2140 5520 -2100
rect 5560 -2140 5870 -2100
rect 5910 -2140 6220 -2100
rect 6260 -2140 6570 -2100
rect 6610 -2140 6920 -2100
rect 6960 -2140 7270 -2100
rect 7310 -2140 7620 -2100
rect 7660 -2140 7970 -2100
rect 8010 -2140 8320 -2100
rect 8360 -2140 8670 -2100
rect 8710 -2125 17990 -2100
rect 8710 -2140 14825 -2125
rect -120 -2165 14825 -2140
rect -120 -2205 -80 -2165
rect -40 -2205 270 -2165
rect 310 -2205 620 -2165
rect 660 -2205 970 -2165
rect 1010 -2205 1320 -2165
rect 1360 -2205 1670 -2165
rect 1710 -2205 2020 -2165
rect 2060 -2205 2370 -2165
rect 2410 -2205 2720 -2165
rect 2760 -2205 3070 -2165
rect 3110 -2205 3420 -2165
rect 3460 -2205 3770 -2165
rect 3810 -2205 4120 -2165
rect 4160 -2205 4470 -2165
rect 4510 -2205 4820 -2165
rect 4860 -2205 5170 -2165
rect 5210 -2205 5520 -2165
rect 5560 -2205 5870 -2165
rect 5910 -2205 6220 -2165
rect 6260 -2205 6570 -2165
rect 6610 -2205 6920 -2165
rect 6960 -2205 7270 -2165
rect 7310 -2205 7620 -2165
rect 7660 -2205 7970 -2165
rect 8010 -2205 8320 -2165
rect 8360 -2205 8670 -2165
rect 8710 -2175 14825 -2165
rect 14875 -2175 14920 -2125
rect 14970 -2175 15015 -2125
rect 15065 -2175 15115 -2125
rect 15165 -2175 15215 -2125
rect 15265 -2175 15315 -2125
rect 15365 -2175 15410 -2125
rect 15460 -2175 15505 -2125
rect 15555 -2175 15625 -2125
rect 15675 -2175 15720 -2125
rect 15770 -2175 15815 -2125
rect 15865 -2175 15915 -2125
rect 15965 -2175 16015 -2125
rect 16065 -2175 16115 -2125
rect 16165 -2175 16210 -2125
rect 16260 -2175 16305 -2125
rect 16355 -2175 16425 -2125
rect 16475 -2175 16520 -2125
rect 16570 -2175 16615 -2125
rect 16665 -2175 16715 -2125
rect 16765 -2175 16815 -2125
rect 16865 -2175 16915 -2125
rect 16965 -2175 17010 -2125
rect 17060 -2175 17105 -2125
rect 17155 -2175 17225 -2125
rect 17275 -2175 17320 -2125
rect 17370 -2175 17415 -2125
rect 17465 -2175 17515 -2125
rect 17565 -2175 17615 -2125
rect 17665 -2175 17715 -2125
rect 17765 -2175 17810 -2125
rect 17860 -2175 17905 -2125
rect 17955 -2175 17990 -2125
rect 8710 -2205 17990 -2175
rect -120 -2215 17990 -2205
rect -120 -2235 14825 -2215
rect -120 -2275 -80 -2235
rect -40 -2275 270 -2235
rect 310 -2275 620 -2235
rect 660 -2275 970 -2235
rect 1010 -2275 1320 -2235
rect 1360 -2275 1670 -2235
rect 1710 -2275 2020 -2235
rect 2060 -2275 2370 -2235
rect 2410 -2275 2720 -2235
rect 2760 -2275 3070 -2235
rect 3110 -2275 3420 -2235
rect 3460 -2275 3770 -2235
rect 3810 -2275 4120 -2235
rect 4160 -2275 4470 -2235
rect 4510 -2275 4820 -2235
rect 4860 -2275 5170 -2235
rect 5210 -2275 5520 -2235
rect 5560 -2275 5870 -2235
rect 5910 -2275 6220 -2235
rect 6260 -2275 6570 -2235
rect 6610 -2275 6920 -2235
rect 6960 -2275 7270 -2235
rect 7310 -2275 7620 -2235
rect 7660 -2275 7970 -2235
rect 8010 -2275 8320 -2235
rect 8360 -2275 8670 -2235
rect 8710 -2265 14825 -2235
rect 14875 -2265 14920 -2215
rect 14970 -2265 15015 -2215
rect 15065 -2265 15115 -2215
rect 15165 -2265 15215 -2215
rect 15265 -2265 15315 -2215
rect 15365 -2265 15410 -2215
rect 15460 -2265 15505 -2215
rect 15555 -2265 15625 -2215
rect 15675 -2265 15720 -2215
rect 15770 -2265 15815 -2215
rect 15865 -2265 15915 -2215
rect 15965 -2265 16015 -2215
rect 16065 -2265 16115 -2215
rect 16165 -2265 16210 -2215
rect 16260 -2265 16305 -2215
rect 16355 -2265 16425 -2215
rect 16475 -2265 16520 -2215
rect 16570 -2265 16615 -2215
rect 16665 -2265 16715 -2215
rect 16765 -2265 16815 -2215
rect 16865 -2265 16915 -2215
rect 16965 -2265 17010 -2215
rect 17060 -2265 17105 -2215
rect 17155 -2265 17225 -2215
rect 17275 -2265 17320 -2215
rect 17370 -2265 17415 -2215
rect 17465 -2265 17515 -2215
rect 17565 -2265 17615 -2215
rect 17665 -2265 17715 -2215
rect 17765 -2265 17810 -2215
rect 17860 -2265 17905 -2215
rect 17955 -2265 17990 -2215
rect 8710 -2275 17990 -2265
rect -120 -2305 17990 -2275
rect -120 -2345 -80 -2305
rect -40 -2345 270 -2305
rect 310 -2345 620 -2305
rect 660 -2345 970 -2305
rect 1010 -2345 1320 -2305
rect 1360 -2345 1670 -2305
rect 1710 -2345 2020 -2305
rect 2060 -2345 2370 -2305
rect 2410 -2345 2720 -2305
rect 2760 -2345 3070 -2305
rect 3110 -2345 3420 -2305
rect 3460 -2345 3770 -2305
rect 3810 -2345 4120 -2305
rect 4160 -2345 4470 -2305
rect 4510 -2345 4820 -2305
rect 4860 -2345 5170 -2305
rect 5210 -2345 5520 -2305
rect 5560 -2345 5870 -2305
rect 5910 -2345 6220 -2305
rect 6260 -2345 6570 -2305
rect 6610 -2345 6920 -2305
rect 6960 -2345 7270 -2305
rect 7310 -2345 7620 -2305
rect 7660 -2345 7970 -2305
rect 8010 -2345 8320 -2305
rect 8360 -2345 8670 -2305
rect 8710 -2315 17990 -2305
rect 8710 -2345 14825 -2315
rect -120 -2365 14825 -2345
rect 14875 -2365 14920 -2315
rect 14970 -2365 15015 -2315
rect 15065 -2365 15115 -2315
rect 15165 -2365 15215 -2315
rect 15265 -2365 15315 -2315
rect 15365 -2365 15410 -2315
rect 15460 -2365 15505 -2315
rect 15555 -2365 15625 -2315
rect 15675 -2365 15720 -2315
rect 15770 -2365 15815 -2315
rect 15865 -2365 15915 -2315
rect 15965 -2365 16015 -2315
rect 16065 -2365 16115 -2315
rect 16165 -2365 16210 -2315
rect 16260 -2365 16305 -2315
rect 16355 -2365 16425 -2315
rect 16475 -2365 16520 -2315
rect 16570 -2365 16615 -2315
rect 16665 -2365 16715 -2315
rect 16765 -2365 16815 -2315
rect 16865 -2365 16915 -2315
rect 16965 -2365 17010 -2315
rect 17060 -2365 17105 -2315
rect 17155 -2365 17225 -2315
rect 17275 -2365 17320 -2315
rect 17370 -2365 17415 -2315
rect 17465 -2365 17515 -2315
rect 17565 -2365 17615 -2315
rect 17665 -2365 17715 -2315
rect 17765 -2365 17810 -2315
rect 17860 -2365 17905 -2315
rect 17955 -2365 17990 -2315
rect -120 -2375 17990 -2365
rect -120 -2415 -80 -2375
rect -40 -2415 270 -2375
rect 310 -2415 620 -2375
rect 660 -2415 970 -2375
rect 1010 -2415 1320 -2375
rect 1360 -2415 1670 -2375
rect 1710 -2415 2020 -2375
rect 2060 -2415 2370 -2375
rect 2410 -2415 2720 -2375
rect 2760 -2415 3070 -2375
rect 3110 -2415 3420 -2375
rect 3460 -2415 3770 -2375
rect 3810 -2415 4120 -2375
rect 4160 -2415 4470 -2375
rect 4510 -2415 4820 -2375
rect 4860 -2415 5170 -2375
rect 5210 -2415 5520 -2375
rect 5560 -2415 5870 -2375
rect 5910 -2415 6220 -2375
rect 6260 -2415 6570 -2375
rect 6610 -2415 6920 -2375
rect 6960 -2415 7270 -2375
rect 7310 -2415 7620 -2375
rect 7660 -2415 7970 -2375
rect 8010 -2415 8320 -2375
rect 8360 -2415 8670 -2375
rect 8710 -2405 17990 -2375
rect 8710 -2415 14825 -2405
rect -120 -2440 14825 -2415
rect -120 -2480 -80 -2440
rect -40 -2480 270 -2440
rect 310 -2480 620 -2440
rect 660 -2480 970 -2440
rect 1010 -2480 1320 -2440
rect 1360 -2480 1670 -2440
rect 1710 -2480 2020 -2440
rect 2060 -2480 2370 -2440
rect 2410 -2480 2720 -2440
rect 2760 -2480 3070 -2440
rect 3110 -2480 3420 -2440
rect 3460 -2480 3770 -2440
rect 3810 -2480 4120 -2440
rect 4160 -2480 4470 -2440
rect 4510 -2480 4820 -2440
rect 4860 -2480 5170 -2440
rect 5210 -2480 5520 -2440
rect 5560 -2480 5870 -2440
rect 5910 -2480 6220 -2440
rect 6260 -2480 6570 -2440
rect 6610 -2480 6920 -2440
rect 6960 -2480 7270 -2440
rect 7310 -2480 7620 -2440
rect 7660 -2480 7970 -2440
rect 8010 -2480 8320 -2440
rect 8360 -2480 8670 -2440
rect 8710 -2455 14825 -2440
rect 14875 -2455 14920 -2405
rect 14970 -2455 15015 -2405
rect 15065 -2455 15115 -2405
rect 15165 -2455 15215 -2405
rect 15265 -2455 15315 -2405
rect 15365 -2455 15410 -2405
rect 15460 -2455 15505 -2405
rect 15555 -2455 15625 -2405
rect 15675 -2455 15720 -2405
rect 15770 -2455 15815 -2405
rect 15865 -2455 15915 -2405
rect 15965 -2455 16015 -2405
rect 16065 -2455 16115 -2405
rect 16165 -2455 16210 -2405
rect 16260 -2455 16305 -2405
rect 16355 -2455 16425 -2405
rect 16475 -2455 16520 -2405
rect 16570 -2455 16615 -2405
rect 16665 -2455 16715 -2405
rect 16765 -2455 16815 -2405
rect 16865 -2455 16915 -2405
rect 16965 -2455 17010 -2405
rect 17060 -2455 17105 -2405
rect 17155 -2455 17225 -2405
rect 17275 -2455 17320 -2405
rect 17370 -2455 17415 -2405
rect 17465 -2455 17515 -2405
rect 17565 -2455 17615 -2405
rect 17665 -2455 17715 -2405
rect 17765 -2455 17810 -2405
rect 17860 -2455 17905 -2405
rect 17955 -2455 17990 -2405
rect 8710 -2480 17990 -2455
rect -120 -2500 17990 -2480
rect -120 -2540 -80 -2500
rect -40 -2540 270 -2500
rect 310 -2540 620 -2500
rect 660 -2540 970 -2500
rect 1010 -2540 1320 -2500
rect 1360 -2540 1670 -2500
rect 1710 -2540 2020 -2500
rect 2060 -2540 2370 -2500
rect 2410 -2540 2720 -2500
rect 2760 -2540 3070 -2500
rect 3110 -2540 3420 -2500
rect 3460 -2540 3770 -2500
rect 3810 -2540 4120 -2500
rect 4160 -2540 4470 -2500
rect 4510 -2540 4820 -2500
rect 4860 -2540 5170 -2500
rect 5210 -2540 5520 -2500
rect 5560 -2540 5870 -2500
rect 5910 -2540 6220 -2500
rect 6260 -2540 6570 -2500
rect 6610 -2540 6920 -2500
rect 6960 -2540 7270 -2500
rect 7310 -2540 7620 -2500
rect 7660 -2540 7970 -2500
rect 8010 -2540 8320 -2500
rect 8360 -2540 8670 -2500
rect 8710 -2525 17990 -2500
rect 8710 -2540 14825 -2525
rect -120 -2565 14825 -2540
rect -120 -2605 -80 -2565
rect -40 -2605 270 -2565
rect 310 -2605 620 -2565
rect 660 -2605 970 -2565
rect 1010 -2605 1320 -2565
rect 1360 -2605 1670 -2565
rect 1710 -2605 2020 -2565
rect 2060 -2605 2370 -2565
rect 2410 -2605 2720 -2565
rect 2760 -2605 3070 -2565
rect 3110 -2605 3420 -2565
rect 3460 -2605 3770 -2565
rect 3810 -2605 4120 -2565
rect 4160 -2605 4470 -2565
rect 4510 -2605 4820 -2565
rect 4860 -2605 5170 -2565
rect 5210 -2605 5520 -2565
rect 5560 -2605 5870 -2565
rect 5910 -2605 6220 -2565
rect 6260 -2605 6570 -2565
rect 6610 -2605 6920 -2565
rect 6960 -2605 7270 -2565
rect 7310 -2605 7620 -2565
rect 7660 -2605 7970 -2565
rect 8010 -2605 8320 -2565
rect 8360 -2605 8670 -2565
rect 8710 -2575 14825 -2565
rect 14875 -2575 14920 -2525
rect 14970 -2575 15015 -2525
rect 15065 -2575 15115 -2525
rect 15165 -2575 15215 -2525
rect 15265 -2575 15315 -2525
rect 15365 -2575 15410 -2525
rect 15460 -2575 15505 -2525
rect 15555 -2575 15625 -2525
rect 15675 -2575 15720 -2525
rect 15770 -2575 15815 -2525
rect 15865 -2575 15915 -2525
rect 15965 -2575 16015 -2525
rect 16065 -2575 16115 -2525
rect 16165 -2575 16210 -2525
rect 16260 -2575 16305 -2525
rect 16355 -2575 16425 -2525
rect 16475 -2575 16520 -2525
rect 16570 -2575 16615 -2525
rect 16665 -2575 16715 -2525
rect 16765 -2575 16815 -2525
rect 16865 -2575 16915 -2525
rect 16965 -2575 17010 -2525
rect 17060 -2575 17105 -2525
rect 17155 -2575 17225 -2525
rect 17275 -2575 17320 -2525
rect 17370 -2575 17415 -2525
rect 17465 -2575 17515 -2525
rect 17565 -2575 17615 -2525
rect 17665 -2575 17715 -2525
rect 17765 -2575 17810 -2525
rect 17860 -2575 17905 -2525
rect 17955 -2575 17990 -2525
rect 8710 -2605 17990 -2575
rect -120 -2615 17990 -2605
rect -120 -2635 14825 -2615
rect -120 -2675 -80 -2635
rect -40 -2675 270 -2635
rect 310 -2675 620 -2635
rect 660 -2675 970 -2635
rect 1010 -2675 1320 -2635
rect 1360 -2675 1670 -2635
rect 1710 -2675 2020 -2635
rect 2060 -2675 2370 -2635
rect 2410 -2675 2720 -2635
rect 2760 -2675 3070 -2635
rect 3110 -2675 3420 -2635
rect 3460 -2675 3770 -2635
rect 3810 -2675 4120 -2635
rect 4160 -2675 4470 -2635
rect 4510 -2675 4820 -2635
rect 4860 -2675 5170 -2635
rect 5210 -2675 5520 -2635
rect 5560 -2675 5870 -2635
rect 5910 -2675 6220 -2635
rect 6260 -2675 6570 -2635
rect 6610 -2675 6920 -2635
rect 6960 -2675 7270 -2635
rect 7310 -2675 7620 -2635
rect 7660 -2675 7970 -2635
rect 8010 -2675 8320 -2635
rect 8360 -2675 8670 -2635
rect 8710 -2665 14825 -2635
rect 14875 -2665 14920 -2615
rect 14970 -2665 15015 -2615
rect 15065 -2665 15115 -2615
rect 15165 -2665 15215 -2615
rect 15265 -2665 15315 -2615
rect 15365 -2665 15410 -2615
rect 15460 -2665 15505 -2615
rect 15555 -2665 15625 -2615
rect 15675 -2665 15720 -2615
rect 15770 -2665 15815 -2615
rect 15865 -2665 15915 -2615
rect 15965 -2665 16015 -2615
rect 16065 -2665 16115 -2615
rect 16165 -2665 16210 -2615
rect 16260 -2665 16305 -2615
rect 16355 -2665 16425 -2615
rect 16475 -2665 16520 -2615
rect 16570 -2665 16615 -2615
rect 16665 -2665 16715 -2615
rect 16765 -2665 16815 -2615
rect 16865 -2665 16915 -2615
rect 16965 -2665 17010 -2615
rect 17060 -2665 17105 -2615
rect 17155 -2665 17225 -2615
rect 17275 -2665 17320 -2615
rect 17370 -2665 17415 -2615
rect 17465 -2665 17515 -2615
rect 17565 -2665 17615 -2615
rect 17665 -2665 17715 -2615
rect 17765 -2665 17810 -2615
rect 17860 -2665 17905 -2615
rect 17955 -2665 17990 -2615
rect 8710 -2675 17990 -2665
rect -120 -2705 17990 -2675
rect -120 -2745 -80 -2705
rect -40 -2745 270 -2705
rect 310 -2745 620 -2705
rect 660 -2745 970 -2705
rect 1010 -2745 1320 -2705
rect 1360 -2745 1670 -2705
rect 1710 -2745 2020 -2705
rect 2060 -2745 2370 -2705
rect 2410 -2745 2720 -2705
rect 2760 -2745 3070 -2705
rect 3110 -2745 3420 -2705
rect 3460 -2745 3770 -2705
rect 3810 -2745 4120 -2705
rect 4160 -2745 4470 -2705
rect 4510 -2745 4820 -2705
rect 4860 -2745 5170 -2705
rect 5210 -2745 5520 -2705
rect 5560 -2745 5870 -2705
rect 5910 -2745 6220 -2705
rect 6260 -2745 6570 -2705
rect 6610 -2745 6920 -2705
rect 6960 -2745 7270 -2705
rect 7310 -2745 7620 -2705
rect 7660 -2745 7970 -2705
rect 8010 -2745 8320 -2705
rect 8360 -2745 8670 -2705
rect 8710 -2715 17990 -2705
rect 8710 -2745 14825 -2715
rect -120 -2765 14825 -2745
rect 14875 -2765 14920 -2715
rect 14970 -2765 15015 -2715
rect 15065 -2765 15115 -2715
rect 15165 -2765 15215 -2715
rect 15265 -2765 15315 -2715
rect 15365 -2765 15410 -2715
rect 15460 -2765 15505 -2715
rect 15555 -2765 15625 -2715
rect 15675 -2765 15720 -2715
rect 15770 -2765 15815 -2715
rect 15865 -2765 15915 -2715
rect 15965 -2765 16015 -2715
rect 16065 -2765 16115 -2715
rect 16165 -2765 16210 -2715
rect 16260 -2765 16305 -2715
rect 16355 -2765 16425 -2715
rect 16475 -2765 16520 -2715
rect 16570 -2765 16615 -2715
rect 16665 -2765 16715 -2715
rect 16765 -2765 16815 -2715
rect 16865 -2765 16915 -2715
rect 16965 -2765 17010 -2715
rect 17060 -2765 17105 -2715
rect 17155 -2765 17225 -2715
rect 17275 -2765 17320 -2715
rect 17370 -2765 17415 -2715
rect 17465 -2765 17515 -2715
rect 17565 -2765 17615 -2715
rect 17665 -2765 17715 -2715
rect 17765 -2765 17810 -2715
rect 17860 -2765 17905 -2715
rect 17955 -2765 17990 -2715
rect -120 -2775 17990 -2765
rect -120 -2815 -80 -2775
rect -40 -2815 270 -2775
rect 310 -2815 620 -2775
rect 660 -2815 970 -2775
rect 1010 -2815 1320 -2775
rect 1360 -2815 1670 -2775
rect 1710 -2815 2020 -2775
rect 2060 -2815 2370 -2775
rect 2410 -2815 2720 -2775
rect 2760 -2815 3070 -2775
rect 3110 -2815 3420 -2775
rect 3460 -2815 3770 -2775
rect 3810 -2815 4120 -2775
rect 4160 -2815 4470 -2775
rect 4510 -2815 4820 -2775
rect 4860 -2815 5170 -2775
rect 5210 -2815 5520 -2775
rect 5560 -2815 5870 -2775
rect 5910 -2815 6220 -2775
rect 6260 -2815 6570 -2775
rect 6610 -2815 6920 -2775
rect 6960 -2815 7270 -2775
rect 7310 -2815 7620 -2775
rect 7660 -2815 7970 -2775
rect 8010 -2815 8320 -2775
rect 8360 -2815 8670 -2775
rect 8710 -2805 17990 -2775
rect 8710 -2815 14825 -2805
rect -120 -2840 14825 -2815
rect -120 -2880 -80 -2840
rect -40 -2880 270 -2840
rect 310 -2880 620 -2840
rect 660 -2880 970 -2840
rect 1010 -2880 1320 -2840
rect 1360 -2880 1670 -2840
rect 1710 -2880 2020 -2840
rect 2060 -2880 2370 -2840
rect 2410 -2880 2720 -2840
rect 2760 -2880 3070 -2840
rect 3110 -2880 3420 -2840
rect 3460 -2880 3770 -2840
rect 3810 -2880 4120 -2840
rect 4160 -2880 4470 -2840
rect 4510 -2880 4820 -2840
rect 4860 -2880 5170 -2840
rect 5210 -2880 5520 -2840
rect 5560 -2880 5870 -2840
rect 5910 -2880 6220 -2840
rect 6260 -2880 6570 -2840
rect 6610 -2880 6920 -2840
rect 6960 -2880 7270 -2840
rect 7310 -2880 7620 -2840
rect 7660 -2880 7970 -2840
rect 8010 -2880 8320 -2840
rect 8360 -2880 8670 -2840
rect 8710 -2855 14825 -2840
rect 14875 -2855 14920 -2805
rect 14970 -2855 15015 -2805
rect 15065 -2855 15115 -2805
rect 15165 -2855 15215 -2805
rect 15265 -2855 15315 -2805
rect 15365 -2855 15410 -2805
rect 15460 -2855 15505 -2805
rect 15555 -2855 15625 -2805
rect 15675 -2855 15720 -2805
rect 15770 -2855 15815 -2805
rect 15865 -2855 15915 -2805
rect 15965 -2855 16015 -2805
rect 16065 -2855 16115 -2805
rect 16165 -2855 16210 -2805
rect 16260 -2855 16305 -2805
rect 16355 -2855 16425 -2805
rect 16475 -2855 16520 -2805
rect 16570 -2855 16615 -2805
rect 16665 -2855 16715 -2805
rect 16765 -2855 16815 -2805
rect 16865 -2855 16915 -2805
rect 16965 -2855 17010 -2805
rect 17060 -2855 17105 -2805
rect 17155 -2855 17225 -2805
rect 17275 -2855 17320 -2805
rect 17370 -2855 17415 -2805
rect 17465 -2855 17515 -2805
rect 17565 -2855 17615 -2805
rect 17665 -2855 17715 -2805
rect 17765 -2855 17810 -2805
rect 17860 -2855 17905 -2805
rect 17955 -2855 17990 -2805
rect 8710 -2880 17990 -2855
rect -120 -2900 17990 -2880
rect -120 -2940 -80 -2900
rect -40 -2940 270 -2900
rect 310 -2940 620 -2900
rect 660 -2940 970 -2900
rect 1010 -2940 1320 -2900
rect 1360 -2940 1670 -2900
rect 1710 -2940 2020 -2900
rect 2060 -2940 2370 -2900
rect 2410 -2940 2720 -2900
rect 2760 -2940 3070 -2900
rect 3110 -2940 3420 -2900
rect 3460 -2940 3770 -2900
rect 3810 -2940 4120 -2900
rect 4160 -2940 4470 -2900
rect 4510 -2940 4820 -2900
rect 4860 -2940 5170 -2900
rect 5210 -2940 5520 -2900
rect 5560 -2940 5870 -2900
rect 5910 -2940 6220 -2900
rect 6260 -2940 6570 -2900
rect 6610 -2940 6920 -2900
rect 6960 -2940 7270 -2900
rect 7310 -2940 7620 -2900
rect 7660 -2940 7970 -2900
rect 8010 -2940 8320 -2900
rect 8360 -2940 8670 -2900
rect 8710 -2925 17990 -2900
rect 8710 -2940 14825 -2925
rect -120 -2965 14825 -2940
rect -120 -3005 -80 -2965
rect -40 -3005 270 -2965
rect 310 -3005 620 -2965
rect 660 -3005 970 -2965
rect 1010 -3005 1320 -2965
rect 1360 -3005 1670 -2965
rect 1710 -3005 2020 -2965
rect 2060 -3005 2370 -2965
rect 2410 -3005 2720 -2965
rect 2760 -3005 3070 -2965
rect 3110 -3005 3420 -2965
rect 3460 -3005 3770 -2965
rect 3810 -3005 4120 -2965
rect 4160 -3005 4470 -2965
rect 4510 -3005 4820 -2965
rect 4860 -3005 5170 -2965
rect 5210 -3005 5520 -2965
rect 5560 -3005 5870 -2965
rect 5910 -3005 6220 -2965
rect 6260 -3005 6570 -2965
rect 6610 -3005 6920 -2965
rect 6960 -3005 7270 -2965
rect 7310 -3005 7620 -2965
rect 7660 -3005 7970 -2965
rect 8010 -3005 8320 -2965
rect 8360 -3005 8670 -2965
rect 8710 -2975 14825 -2965
rect 14875 -2975 14920 -2925
rect 14970 -2975 15015 -2925
rect 15065 -2975 15115 -2925
rect 15165 -2975 15215 -2925
rect 15265 -2975 15315 -2925
rect 15365 -2975 15410 -2925
rect 15460 -2975 15505 -2925
rect 15555 -2975 15625 -2925
rect 15675 -2975 15720 -2925
rect 15770 -2975 15815 -2925
rect 15865 -2975 15915 -2925
rect 15965 -2975 16015 -2925
rect 16065 -2975 16115 -2925
rect 16165 -2975 16210 -2925
rect 16260 -2975 16305 -2925
rect 16355 -2975 16425 -2925
rect 16475 -2975 16520 -2925
rect 16570 -2975 16615 -2925
rect 16665 -2975 16715 -2925
rect 16765 -2975 16815 -2925
rect 16865 -2975 16915 -2925
rect 16965 -2975 17010 -2925
rect 17060 -2975 17105 -2925
rect 17155 -2975 17225 -2925
rect 17275 -2975 17320 -2925
rect 17370 -2975 17415 -2925
rect 17465 -2975 17515 -2925
rect 17565 -2975 17615 -2925
rect 17665 -2975 17715 -2925
rect 17765 -2975 17810 -2925
rect 17860 -2975 17905 -2925
rect 17955 -2975 17990 -2925
rect 8710 -3005 17990 -2975
rect -120 -3015 17990 -3005
rect -120 -3035 14825 -3015
rect -120 -3075 -80 -3035
rect -40 -3075 270 -3035
rect 310 -3075 620 -3035
rect 660 -3075 970 -3035
rect 1010 -3075 1320 -3035
rect 1360 -3075 1670 -3035
rect 1710 -3075 2020 -3035
rect 2060 -3075 2370 -3035
rect 2410 -3075 2720 -3035
rect 2760 -3075 3070 -3035
rect 3110 -3075 3420 -3035
rect 3460 -3075 3770 -3035
rect 3810 -3075 4120 -3035
rect 4160 -3075 4470 -3035
rect 4510 -3075 4820 -3035
rect 4860 -3075 5170 -3035
rect 5210 -3075 5520 -3035
rect 5560 -3075 5870 -3035
rect 5910 -3075 6220 -3035
rect 6260 -3075 6570 -3035
rect 6610 -3075 6920 -3035
rect 6960 -3075 7270 -3035
rect 7310 -3075 7620 -3035
rect 7660 -3075 7970 -3035
rect 8010 -3075 8320 -3035
rect 8360 -3075 8670 -3035
rect 8710 -3065 14825 -3035
rect 14875 -3065 14920 -3015
rect 14970 -3065 15015 -3015
rect 15065 -3065 15115 -3015
rect 15165 -3065 15215 -3015
rect 15265 -3065 15315 -3015
rect 15365 -3065 15410 -3015
rect 15460 -3065 15505 -3015
rect 15555 -3065 15625 -3015
rect 15675 -3065 15720 -3015
rect 15770 -3065 15815 -3015
rect 15865 -3065 15915 -3015
rect 15965 -3065 16015 -3015
rect 16065 -3065 16115 -3015
rect 16165 -3065 16210 -3015
rect 16260 -3065 16305 -3015
rect 16355 -3065 16425 -3015
rect 16475 -3065 16520 -3015
rect 16570 -3065 16615 -3015
rect 16665 -3065 16715 -3015
rect 16765 -3065 16815 -3015
rect 16865 -3065 16915 -3015
rect 16965 -3065 17010 -3015
rect 17060 -3065 17105 -3015
rect 17155 -3065 17225 -3015
rect 17275 -3065 17320 -3015
rect 17370 -3065 17415 -3015
rect 17465 -3065 17515 -3015
rect 17565 -3065 17615 -3015
rect 17665 -3065 17715 -3015
rect 17765 -3065 17810 -3015
rect 17860 -3065 17905 -3015
rect 17955 -3065 17990 -3015
rect 8710 -3075 17990 -3065
rect -120 -3105 17990 -3075
rect -120 -3145 -80 -3105
rect -40 -3145 270 -3105
rect 310 -3145 620 -3105
rect 660 -3145 970 -3105
rect 1010 -3145 1320 -3105
rect 1360 -3145 1670 -3105
rect 1710 -3145 2020 -3105
rect 2060 -3145 2370 -3105
rect 2410 -3145 2720 -3105
rect 2760 -3145 3070 -3105
rect 3110 -3145 3420 -3105
rect 3460 -3145 3770 -3105
rect 3810 -3145 4120 -3105
rect 4160 -3145 4470 -3105
rect 4510 -3145 4820 -3105
rect 4860 -3145 5170 -3105
rect 5210 -3145 5520 -3105
rect 5560 -3145 5870 -3105
rect 5910 -3145 6220 -3105
rect 6260 -3145 6570 -3105
rect 6610 -3145 6920 -3105
rect 6960 -3145 7270 -3105
rect 7310 -3145 7620 -3105
rect 7660 -3145 7970 -3105
rect 8010 -3145 8320 -3105
rect 8360 -3145 8670 -3105
rect 8710 -3115 17990 -3105
rect 8710 -3145 14825 -3115
rect -120 -3165 14825 -3145
rect 14875 -3165 14920 -3115
rect 14970 -3165 15015 -3115
rect 15065 -3165 15115 -3115
rect 15165 -3165 15215 -3115
rect 15265 -3165 15315 -3115
rect 15365 -3165 15410 -3115
rect 15460 -3165 15505 -3115
rect 15555 -3165 15625 -3115
rect 15675 -3165 15720 -3115
rect 15770 -3165 15815 -3115
rect 15865 -3165 15915 -3115
rect 15965 -3165 16015 -3115
rect 16065 -3165 16115 -3115
rect 16165 -3165 16210 -3115
rect 16260 -3165 16305 -3115
rect 16355 -3165 16425 -3115
rect 16475 -3165 16520 -3115
rect 16570 -3165 16615 -3115
rect 16665 -3165 16715 -3115
rect 16765 -3165 16815 -3115
rect 16865 -3165 16915 -3115
rect 16965 -3165 17010 -3115
rect 17060 -3165 17105 -3115
rect 17155 -3165 17225 -3115
rect 17275 -3165 17320 -3115
rect 17370 -3165 17415 -3115
rect 17465 -3165 17515 -3115
rect 17565 -3165 17615 -3115
rect 17665 -3165 17715 -3115
rect 17765 -3165 17810 -3115
rect 17860 -3165 17905 -3115
rect 17955 -3165 17990 -3115
rect -120 -3175 17990 -3165
rect -120 -3215 -80 -3175
rect -40 -3215 270 -3175
rect 310 -3215 620 -3175
rect 660 -3215 970 -3175
rect 1010 -3215 1320 -3175
rect 1360 -3215 1670 -3175
rect 1710 -3215 2020 -3175
rect 2060 -3215 2370 -3175
rect 2410 -3215 2720 -3175
rect 2760 -3215 3070 -3175
rect 3110 -3215 3420 -3175
rect 3460 -3215 3770 -3175
rect 3810 -3215 4120 -3175
rect 4160 -3215 4470 -3175
rect 4510 -3215 4820 -3175
rect 4860 -3215 5170 -3175
rect 5210 -3215 5520 -3175
rect 5560 -3215 5870 -3175
rect 5910 -3215 6220 -3175
rect 6260 -3215 6570 -3175
rect 6610 -3215 6920 -3175
rect 6960 -3215 7270 -3175
rect 7310 -3215 7620 -3175
rect 7660 -3215 7970 -3175
rect 8010 -3215 8320 -3175
rect 8360 -3215 8670 -3175
rect 8710 -3205 17990 -3175
rect 8710 -3215 14825 -3205
rect -120 -3240 14825 -3215
rect -120 -3280 -80 -3240
rect -40 -3280 270 -3240
rect 310 -3280 620 -3240
rect 660 -3280 970 -3240
rect 1010 -3280 1320 -3240
rect 1360 -3280 1670 -3240
rect 1710 -3280 2020 -3240
rect 2060 -3280 2370 -3240
rect 2410 -3280 2720 -3240
rect 2760 -3280 3070 -3240
rect 3110 -3280 3420 -3240
rect 3460 -3280 3770 -3240
rect 3810 -3280 4120 -3240
rect 4160 -3280 4470 -3240
rect 4510 -3280 4820 -3240
rect 4860 -3280 5170 -3240
rect 5210 -3280 5520 -3240
rect 5560 -3280 5870 -3240
rect 5910 -3280 6220 -3240
rect 6260 -3280 6570 -3240
rect 6610 -3280 6920 -3240
rect 6960 -3280 7270 -3240
rect 7310 -3280 7620 -3240
rect 7660 -3280 7970 -3240
rect 8010 -3280 8320 -3240
rect 8360 -3280 8670 -3240
rect 8710 -3255 14825 -3240
rect 14875 -3255 14920 -3205
rect 14970 -3255 15015 -3205
rect 15065 -3255 15115 -3205
rect 15165 -3255 15215 -3205
rect 15265 -3255 15315 -3205
rect 15365 -3255 15410 -3205
rect 15460 -3255 15505 -3205
rect 15555 -3255 15625 -3205
rect 15675 -3255 15720 -3205
rect 15770 -3255 15815 -3205
rect 15865 -3255 15915 -3205
rect 15965 -3255 16015 -3205
rect 16065 -3255 16115 -3205
rect 16165 -3255 16210 -3205
rect 16260 -3255 16305 -3205
rect 16355 -3255 16425 -3205
rect 16475 -3255 16520 -3205
rect 16570 -3255 16615 -3205
rect 16665 -3255 16715 -3205
rect 16765 -3255 16815 -3205
rect 16865 -3255 16915 -3205
rect 16965 -3255 17010 -3205
rect 17060 -3255 17105 -3205
rect 17155 -3255 17225 -3205
rect 17275 -3255 17320 -3205
rect 17370 -3255 17415 -3205
rect 17465 -3255 17515 -3205
rect 17565 -3255 17615 -3205
rect 17665 -3255 17715 -3205
rect 17765 -3255 17810 -3205
rect 17860 -3255 17905 -3205
rect 17955 -3255 17990 -3205
rect 8710 -3280 17990 -3255
rect -120 -3300 17990 -3280
rect -120 -3340 -80 -3300
rect -40 -3340 270 -3300
rect 310 -3340 620 -3300
rect 660 -3340 970 -3300
rect 1010 -3340 1320 -3300
rect 1360 -3340 1670 -3300
rect 1710 -3340 2020 -3300
rect 2060 -3340 2370 -3300
rect 2410 -3340 2720 -3300
rect 2760 -3340 3070 -3300
rect 3110 -3340 3420 -3300
rect 3460 -3340 3770 -3300
rect 3810 -3340 4120 -3300
rect 4160 -3340 4470 -3300
rect 4510 -3340 4820 -3300
rect 4860 -3340 5170 -3300
rect 5210 -3340 5520 -3300
rect 5560 -3340 5870 -3300
rect 5910 -3340 6220 -3300
rect 6260 -3340 6570 -3300
rect 6610 -3340 6920 -3300
rect 6960 -3340 7270 -3300
rect 7310 -3340 7620 -3300
rect 7660 -3340 7970 -3300
rect 8010 -3340 8320 -3300
rect 8360 -3340 8670 -3300
rect 8710 -3325 17990 -3300
rect 8710 -3340 14825 -3325
rect -120 -3365 14825 -3340
rect -120 -3405 -80 -3365
rect -40 -3405 270 -3365
rect 310 -3405 620 -3365
rect 660 -3405 970 -3365
rect 1010 -3405 1320 -3365
rect 1360 -3405 1670 -3365
rect 1710 -3405 2020 -3365
rect 2060 -3405 2370 -3365
rect 2410 -3405 2720 -3365
rect 2760 -3405 3070 -3365
rect 3110 -3405 3420 -3365
rect 3460 -3405 3770 -3365
rect 3810 -3405 4120 -3365
rect 4160 -3405 4470 -3365
rect 4510 -3405 4820 -3365
rect 4860 -3405 5170 -3365
rect 5210 -3405 5520 -3365
rect 5560 -3405 5870 -3365
rect 5910 -3405 6220 -3365
rect 6260 -3405 6570 -3365
rect 6610 -3405 6920 -3365
rect 6960 -3405 7270 -3365
rect 7310 -3405 7620 -3365
rect 7660 -3405 7970 -3365
rect 8010 -3405 8320 -3365
rect 8360 -3405 8670 -3365
rect 8710 -3375 14825 -3365
rect 14875 -3375 14920 -3325
rect 14970 -3375 15015 -3325
rect 15065 -3375 15115 -3325
rect 15165 -3375 15215 -3325
rect 15265 -3375 15315 -3325
rect 15365 -3375 15410 -3325
rect 15460 -3375 15505 -3325
rect 15555 -3375 15625 -3325
rect 15675 -3375 15720 -3325
rect 15770 -3375 15815 -3325
rect 15865 -3375 15915 -3325
rect 15965 -3375 16015 -3325
rect 16065 -3375 16115 -3325
rect 16165 -3375 16210 -3325
rect 16260 -3375 16305 -3325
rect 16355 -3375 16425 -3325
rect 16475 -3375 16520 -3325
rect 16570 -3375 16615 -3325
rect 16665 -3375 16715 -3325
rect 16765 -3375 16815 -3325
rect 16865 -3375 16915 -3325
rect 16965 -3375 17010 -3325
rect 17060 -3375 17105 -3325
rect 17155 -3375 17225 -3325
rect 17275 -3375 17320 -3325
rect 17370 -3375 17415 -3325
rect 17465 -3375 17515 -3325
rect 17565 -3375 17615 -3325
rect 17665 -3375 17715 -3325
rect 17765 -3375 17810 -3325
rect 17860 -3375 17905 -3325
rect 17955 -3375 17990 -3325
rect 8710 -3405 17990 -3375
rect -120 -3415 17990 -3405
rect -120 -3435 14825 -3415
rect -120 -3475 -80 -3435
rect -40 -3475 270 -3435
rect 310 -3475 620 -3435
rect 660 -3475 970 -3435
rect 1010 -3475 1320 -3435
rect 1360 -3475 1670 -3435
rect 1710 -3475 2020 -3435
rect 2060 -3475 2370 -3435
rect 2410 -3475 2720 -3435
rect 2760 -3475 3070 -3435
rect 3110 -3475 3420 -3435
rect 3460 -3475 3770 -3435
rect 3810 -3475 4120 -3435
rect 4160 -3475 4470 -3435
rect 4510 -3475 4820 -3435
rect 4860 -3475 5170 -3435
rect 5210 -3475 5520 -3435
rect 5560 -3475 5870 -3435
rect 5910 -3475 6220 -3435
rect 6260 -3475 6570 -3435
rect 6610 -3475 6920 -3435
rect 6960 -3475 7270 -3435
rect 7310 -3475 7620 -3435
rect 7660 -3475 7970 -3435
rect 8010 -3475 8320 -3435
rect 8360 -3475 8670 -3435
rect 8710 -3465 14825 -3435
rect 14875 -3465 14920 -3415
rect 14970 -3465 15015 -3415
rect 15065 -3465 15115 -3415
rect 15165 -3465 15215 -3415
rect 15265 -3465 15315 -3415
rect 15365 -3465 15410 -3415
rect 15460 -3465 15505 -3415
rect 15555 -3465 15625 -3415
rect 15675 -3465 15720 -3415
rect 15770 -3465 15815 -3415
rect 15865 -3465 15915 -3415
rect 15965 -3465 16015 -3415
rect 16065 -3465 16115 -3415
rect 16165 -3465 16210 -3415
rect 16260 -3465 16305 -3415
rect 16355 -3465 16425 -3415
rect 16475 -3465 16520 -3415
rect 16570 -3465 16615 -3415
rect 16665 -3465 16715 -3415
rect 16765 -3465 16815 -3415
rect 16865 -3465 16915 -3415
rect 16965 -3465 17010 -3415
rect 17060 -3465 17105 -3415
rect 17155 -3465 17225 -3415
rect 17275 -3465 17320 -3415
rect 17370 -3465 17415 -3415
rect 17465 -3465 17515 -3415
rect 17565 -3465 17615 -3415
rect 17665 -3465 17715 -3415
rect 17765 -3465 17810 -3415
rect 17860 -3465 17905 -3415
rect 17955 -3465 17990 -3415
rect 8710 -3475 17990 -3465
rect -120 -3505 17990 -3475
rect -120 -3545 -80 -3505
rect -40 -3545 270 -3505
rect 310 -3545 620 -3505
rect 660 -3545 970 -3505
rect 1010 -3545 1320 -3505
rect 1360 -3545 1670 -3505
rect 1710 -3545 2020 -3505
rect 2060 -3545 2370 -3505
rect 2410 -3545 2720 -3505
rect 2760 -3545 3070 -3505
rect 3110 -3545 3420 -3505
rect 3460 -3545 3770 -3505
rect 3810 -3545 4120 -3505
rect 4160 -3545 4470 -3505
rect 4510 -3545 4820 -3505
rect 4860 -3545 5170 -3505
rect 5210 -3545 5520 -3505
rect 5560 -3545 5870 -3505
rect 5910 -3545 6220 -3505
rect 6260 -3545 6570 -3505
rect 6610 -3545 6920 -3505
rect 6960 -3545 7270 -3505
rect 7310 -3545 7620 -3505
rect 7660 -3545 7970 -3505
rect 8010 -3545 8320 -3505
rect 8360 -3545 8670 -3505
rect 8710 -3515 17990 -3505
rect 8710 -3545 14825 -3515
rect -120 -3565 14825 -3545
rect 14875 -3565 14920 -3515
rect 14970 -3565 15015 -3515
rect 15065 -3565 15115 -3515
rect 15165 -3565 15215 -3515
rect 15265 -3565 15315 -3515
rect 15365 -3565 15410 -3515
rect 15460 -3565 15505 -3515
rect 15555 -3565 15625 -3515
rect 15675 -3565 15720 -3515
rect 15770 -3565 15815 -3515
rect 15865 -3565 15915 -3515
rect 15965 -3565 16015 -3515
rect 16065 -3565 16115 -3515
rect 16165 -3565 16210 -3515
rect 16260 -3565 16305 -3515
rect 16355 -3565 16425 -3515
rect 16475 -3565 16520 -3515
rect 16570 -3565 16615 -3515
rect 16665 -3565 16715 -3515
rect 16765 -3565 16815 -3515
rect 16865 -3565 16915 -3515
rect 16965 -3565 17010 -3515
rect 17060 -3565 17105 -3515
rect 17155 -3565 17225 -3515
rect 17275 -3565 17320 -3515
rect 17370 -3565 17415 -3515
rect 17465 -3565 17515 -3515
rect 17565 -3565 17615 -3515
rect 17665 -3565 17715 -3515
rect 17765 -3565 17810 -3515
rect 17860 -3565 17905 -3515
rect 17955 -3565 17990 -3515
rect -120 -3575 17990 -3565
rect -120 -3615 -80 -3575
rect -40 -3615 270 -3575
rect 310 -3615 620 -3575
rect 660 -3615 970 -3575
rect 1010 -3615 1320 -3575
rect 1360 -3615 1670 -3575
rect 1710 -3615 2020 -3575
rect 2060 -3615 2370 -3575
rect 2410 -3615 2720 -3575
rect 2760 -3615 3070 -3575
rect 3110 -3615 3420 -3575
rect 3460 -3615 3770 -3575
rect 3810 -3615 4120 -3575
rect 4160 -3615 4470 -3575
rect 4510 -3615 4820 -3575
rect 4860 -3615 5170 -3575
rect 5210 -3615 5520 -3575
rect 5560 -3615 5870 -3575
rect 5910 -3615 6220 -3575
rect 6260 -3615 6570 -3575
rect 6610 -3615 6920 -3575
rect 6960 -3615 7270 -3575
rect 7310 -3615 7620 -3575
rect 7660 -3615 7970 -3575
rect 8010 -3615 8320 -3575
rect 8360 -3615 8670 -3575
rect 8710 -3605 17990 -3575
rect 8710 -3615 14825 -3605
rect -120 -3640 14825 -3615
rect -120 -3680 -80 -3640
rect -40 -3680 270 -3640
rect 310 -3680 620 -3640
rect 660 -3680 970 -3640
rect 1010 -3680 1320 -3640
rect 1360 -3680 1670 -3640
rect 1710 -3680 2020 -3640
rect 2060 -3680 2370 -3640
rect 2410 -3680 2720 -3640
rect 2760 -3680 3070 -3640
rect 3110 -3680 3420 -3640
rect 3460 -3680 3770 -3640
rect 3810 -3680 4120 -3640
rect 4160 -3680 4470 -3640
rect 4510 -3680 4820 -3640
rect 4860 -3680 5170 -3640
rect 5210 -3680 5520 -3640
rect 5560 -3680 5870 -3640
rect 5910 -3680 6220 -3640
rect 6260 -3680 6570 -3640
rect 6610 -3680 6920 -3640
rect 6960 -3680 7270 -3640
rect 7310 -3680 7620 -3640
rect 7660 -3680 7970 -3640
rect 8010 -3680 8320 -3640
rect 8360 -3680 8670 -3640
rect 8710 -3655 14825 -3640
rect 14875 -3655 14920 -3605
rect 14970 -3655 15015 -3605
rect 15065 -3655 15115 -3605
rect 15165 -3655 15215 -3605
rect 15265 -3655 15315 -3605
rect 15365 -3655 15410 -3605
rect 15460 -3655 15505 -3605
rect 15555 -3655 15625 -3605
rect 15675 -3655 15720 -3605
rect 15770 -3655 15815 -3605
rect 15865 -3655 15915 -3605
rect 15965 -3655 16015 -3605
rect 16065 -3655 16115 -3605
rect 16165 -3655 16210 -3605
rect 16260 -3655 16305 -3605
rect 16355 -3655 16425 -3605
rect 16475 -3655 16520 -3605
rect 16570 -3655 16615 -3605
rect 16665 -3655 16715 -3605
rect 16765 -3655 16815 -3605
rect 16865 -3655 16915 -3605
rect 16965 -3655 17010 -3605
rect 17060 -3655 17105 -3605
rect 17155 -3655 17225 -3605
rect 17275 -3655 17320 -3605
rect 17370 -3655 17415 -3605
rect 17465 -3655 17515 -3605
rect 17565 -3655 17615 -3605
rect 17665 -3655 17715 -3605
rect 17765 -3655 17810 -3605
rect 17860 -3655 17905 -3605
rect 17955 -3655 17990 -3605
rect 8710 -3680 17990 -3655
rect -120 -3700 17990 -3680
rect -120 -3740 -80 -3700
rect -40 -3740 270 -3700
rect 310 -3740 620 -3700
rect 660 -3740 970 -3700
rect 1010 -3740 1320 -3700
rect 1360 -3740 1670 -3700
rect 1710 -3740 2020 -3700
rect 2060 -3740 2370 -3700
rect 2410 -3740 2720 -3700
rect 2760 -3740 3070 -3700
rect 3110 -3740 3420 -3700
rect 3460 -3740 3770 -3700
rect 3810 -3740 4120 -3700
rect 4160 -3740 4470 -3700
rect 4510 -3740 4820 -3700
rect 4860 -3740 5170 -3700
rect 5210 -3740 5520 -3700
rect 5560 -3740 5870 -3700
rect 5910 -3740 6220 -3700
rect 6260 -3740 6570 -3700
rect 6610 -3740 6920 -3700
rect 6960 -3740 7270 -3700
rect 7310 -3740 7620 -3700
rect 7660 -3740 7970 -3700
rect 8010 -3740 8320 -3700
rect 8360 -3740 8670 -3700
rect 8710 -3725 17990 -3700
rect 8710 -3740 14825 -3725
rect -120 -3765 14825 -3740
rect -120 -3805 -80 -3765
rect -40 -3805 270 -3765
rect 310 -3805 620 -3765
rect 660 -3805 970 -3765
rect 1010 -3805 1320 -3765
rect 1360 -3805 1670 -3765
rect 1710 -3805 2020 -3765
rect 2060 -3805 2370 -3765
rect 2410 -3805 2720 -3765
rect 2760 -3805 3070 -3765
rect 3110 -3805 3420 -3765
rect 3460 -3805 3770 -3765
rect 3810 -3805 4120 -3765
rect 4160 -3805 4470 -3765
rect 4510 -3805 4820 -3765
rect 4860 -3805 5170 -3765
rect 5210 -3805 5520 -3765
rect 5560 -3805 5870 -3765
rect 5910 -3805 6220 -3765
rect 6260 -3805 6570 -3765
rect 6610 -3805 6920 -3765
rect 6960 -3805 7270 -3765
rect 7310 -3805 7620 -3765
rect 7660 -3805 7970 -3765
rect 8010 -3805 8320 -3765
rect 8360 -3805 8670 -3765
rect 8710 -3775 14825 -3765
rect 14875 -3775 14920 -3725
rect 14970 -3775 15015 -3725
rect 15065 -3775 15115 -3725
rect 15165 -3775 15215 -3725
rect 15265 -3775 15315 -3725
rect 15365 -3775 15410 -3725
rect 15460 -3775 15505 -3725
rect 15555 -3775 15625 -3725
rect 15675 -3775 15720 -3725
rect 15770 -3775 15815 -3725
rect 15865 -3775 15915 -3725
rect 15965 -3775 16015 -3725
rect 16065 -3775 16115 -3725
rect 16165 -3775 16210 -3725
rect 16260 -3775 16305 -3725
rect 16355 -3775 16425 -3725
rect 16475 -3775 16520 -3725
rect 16570 -3775 16615 -3725
rect 16665 -3775 16715 -3725
rect 16765 -3775 16815 -3725
rect 16865 -3775 16915 -3725
rect 16965 -3775 17010 -3725
rect 17060 -3775 17105 -3725
rect 17155 -3775 17225 -3725
rect 17275 -3775 17320 -3725
rect 17370 -3775 17415 -3725
rect 17465 -3775 17515 -3725
rect 17565 -3775 17615 -3725
rect 17665 -3775 17715 -3725
rect 17765 -3775 17810 -3725
rect 17860 -3775 17905 -3725
rect 17955 -3775 17990 -3725
rect 8710 -3805 17990 -3775
rect -120 -3815 17990 -3805
rect -120 -3835 14825 -3815
rect -120 -3875 -80 -3835
rect -40 -3875 270 -3835
rect 310 -3875 620 -3835
rect 660 -3875 970 -3835
rect 1010 -3875 1320 -3835
rect 1360 -3875 1670 -3835
rect 1710 -3875 2020 -3835
rect 2060 -3875 2370 -3835
rect 2410 -3875 2720 -3835
rect 2760 -3875 3070 -3835
rect 3110 -3875 3420 -3835
rect 3460 -3875 3770 -3835
rect 3810 -3875 4120 -3835
rect 4160 -3875 4470 -3835
rect 4510 -3875 4820 -3835
rect 4860 -3875 5170 -3835
rect 5210 -3875 5520 -3835
rect 5560 -3875 5870 -3835
rect 5910 -3875 6220 -3835
rect 6260 -3875 6570 -3835
rect 6610 -3875 6920 -3835
rect 6960 -3875 7270 -3835
rect 7310 -3875 7620 -3835
rect 7660 -3875 7970 -3835
rect 8010 -3875 8320 -3835
rect 8360 -3875 8670 -3835
rect 8710 -3865 14825 -3835
rect 14875 -3865 14920 -3815
rect 14970 -3865 15015 -3815
rect 15065 -3865 15115 -3815
rect 15165 -3865 15215 -3815
rect 15265 -3865 15315 -3815
rect 15365 -3865 15410 -3815
rect 15460 -3865 15505 -3815
rect 15555 -3865 15625 -3815
rect 15675 -3865 15720 -3815
rect 15770 -3865 15815 -3815
rect 15865 -3865 15915 -3815
rect 15965 -3865 16015 -3815
rect 16065 -3865 16115 -3815
rect 16165 -3865 16210 -3815
rect 16260 -3865 16305 -3815
rect 16355 -3865 16425 -3815
rect 16475 -3865 16520 -3815
rect 16570 -3865 16615 -3815
rect 16665 -3865 16715 -3815
rect 16765 -3865 16815 -3815
rect 16865 -3865 16915 -3815
rect 16965 -3865 17010 -3815
rect 17060 -3865 17105 -3815
rect 17155 -3865 17225 -3815
rect 17275 -3865 17320 -3815
rect 17370 -3865 17415 -3815
rect 17465 -3865 17515 -3815
rect 17565 -3865 17615 -3815
rect 17665 -3865 17715 -3815
rect 17765 -3865 17810 -3815
rect 17860 -3865 17905 -3815
rect 17955 -3865 17990 -3815
rect 8710 -3875 17990 -3865
rect -120 -3905 17990 -3875
rect -120 -3945 -80 -3905
rect -40 -3945 270 -3905
rect 310 -3945 620 -3905
rect 660 -3945 970 -3905
rect 1010 -3945 1320 -3905
rect 1360 -3945 1670 -3905
rect 1710 -3945 2020 -3905
rect 2060 -3945 2370 -3905
rect 2410 -3945 2720 -3905
rect 2760 -3945 3070 -3905
rect 3110 -3945 3420 -3905
rect 3460 -3945 3770 -3905
rect 3810 -3945 4120 -3905
rect 4160 -3945 4470 -3905
rect 4510 -3945 4820 -3905
rect 4860 -3945 5170 -3905
rect 5210 -3945 5520 -3905
rect 5560 -3945 5870 -3905
rect 5910 -3945 6220 -3905
rect 6260 -3945 6570 -3905
rect 6610 -3945 6920 -3905
rect 6960 -3945 7270 -3905
rect 7310 -3945 7620 -3905
rect 7660 -3945 7970 -3905
rect 8010 -3945 8320 -3905
rect 8360 -3945 8670 -3905
rect 8710 -3915 17990 -3905
rect 8710 -3945 14825 -3915
rect -120 -3965 14825 -3945
rect 14875 -3965 14920 -3915
rect 14970 -3965 15015 -3915
rect 15065 -3965 15115 -3915
rect 15165 -3965 15215 -3915
rect 15265 -3965 15315 -3915
rect 15365 -3965 15410 -3915
rect 15460 -3965 15505 -3915
rect 15555 -3965 15625 -3915
rect 15675 -3965 15720 -3915
rect 15770 -3965 15815 -3915
rect 15865 -3965 15915 -3915
rect 15965 -3965 16015 -3915
rect 16065 -3965 16115 -3915
rect 16165 -3965 16210 -3915
rect 16260 -3965 16305 -3915
rect 16355 -3965 16425 -3915
rect 16475 -3965 16520 -3915
rect 16570 -3965 16615 -3915
rect 16665 -3965 16715 -3915
rect 16765 -3965 16815 -3915
rect 16865 -3965 16915 -3915
rect 16965 -3965 17010 -3915
rect 17060 -3965 17105 -3915
rect 17155 -3965 17225 -3915
rect 17275 -3965 17320 -3915
rect 17370 -3965 17415 -3915
rect 17465 -3965 17515 -3915
rect 17565 -3965 17615 -3915
rect 17665 -3965 17715 -3915
rect 17765 -3965 17810 -3915
rect 17860 -3965 17905 -3915
rect 17955 -3965 17990 -3915
rect -120 -3975 17990 -3965
rect -120 -4015 -80 -3975
rect -40 -4015 270 -3975
rect 310 -4015 620 -3975
rect 660 -4015 970 -3975
rect 1010 -4015 1320 -3975
rect 1360 -4015 1670 -3975
rect 1710 -4015 2020 -3975
rect 2060 -4015 2370 -3975
rect 2410 -4015 2720 -3975
rect 2760 -4015 3070 -3975
rect 3110 -4015 3420 -3975
rect 3460 -4015 3770 -3975
rect 3810 -4015 4120 -3975
rect 4160 -4015 4470 -3975
rect 4510 -4015 4820 -3975
rect 4860 -4015 5170 -3975
rect 5210 -4015 5520 -3975
rect 5560 -4015 5870 -3975
rect 5910 -4015 6220 -3975
rect 6260 -4015 6570 -3975
rect 6610 -4015 6920 -3975
rect 6960 -4015 7270 -3975
rect 7310 -4015 7620 -3975
rect 7660 -4015 7970 -3975
rect 8010 -4015 8320 -3975
rect 8360 -4015 8670 -3975
rect 8710 -4005 17990 -3975
rect 8710 -4015 14825 -4005
rect -120 -4040 14825 -4015
rect -120 -4080 -80 -4040
rect -40 -4080 270 -4040
rect 310 -4080 620 -4040
rect 660 -4080 970 -4040
rect 1010 -4080 1320 -4040
rect 1360 -4080 1670 -4040
rect 1710 -4080 2020 -4040
rect 2060 -4080 2370 -4040
rect 2410 -4080 2720 -4040
rect 2760 -4080 3070 -4040
rect 3110 -4080 3420 -4040
rect 3460 -4080 3770 -4040
rect 3810 -4080 4120 -4040
rect 4160 -4080 4470 -4040
rect 4510 -4080 4820 -4040
rect 4860 -4080 5170 -4040
rect 5210 -4080 5520 -4040
rect 5560 -4080 5870 -4040
rect 5910 -4080 6220 -4040
rect 6260 -4080 6570 -4040
rect 6610 -4080 6920 -4040
rect 6960 -4080 7270 -4040
rect 7310 -4080 7620 -4040
rect 7660 -4080 7970 -4040
rect 8010 -4080 8320 -4040
rect 8360 -4080 8670 -4040
rect 8710 -4055 14825 -4040
rect 14875 -4055 14920 -4005
rect 14970 -4055 15015 -4005
rect 15065 -4055 15115 -4005
rect 15165 -4055 15215 -4005
rect 15265 -4055 15315 -4005
rect 15365 -4055 15410 -4005
rect 15460 -4055 15505 -4005
rect 15555 -4055 15625 -4005
rect 15675 -4055 15720 -4005
rect 15770 -4055 15815 -4005
rect 15865 -4055 15915 -4005
rect 15965 -4055 16015 -4005
rect 16065 -4055 16115 -4005
rect 16165 -4055 16210 -4005
rect 16260 -4055 16305 -4005
rect 16355 -4055 16425 -4005
rect 16475 -4055 16520 -4005
rect 16570 -4055 16615 -4005
rect 16665 -4055 16715 -4005
rect 16765 -4055 16815 -4005
rect 16865 -4055 16915 -4005
rect 16965 -4055 17010 -4005
rect 17060 -4055 17105 -4005
rect 17155 -4055 17225 -4005
rect 17275 -4055 17320 -4005
rect 17370 -4055 17415 -4005
rect 17465 -4055 17515 -4005
rect 17565 -4055 17615 -4005
rect 17665 -4055 17715 -4005
rect 17765 -4055 17810 -4005
rect 17860 -4055 17905 -4005
rect 17955 -4055 17990 -4005
rect 8710 -4080 17990 -4055
rect -120 -4100 17990 -4080
rect -120 -4140 -80 -4100
rect -40 -4140 270 -4100
rect 310 -4140 620 -4100
rect 660 -4140 970 -4100
rect 1010 -4140 1320 -4100
rect 1360 -4140 1670 -4100
rect 1710 -4140 2020 -4100
rect 2060 -4140 2370 -4100
rect 2410 -4140 2720 -4100
rect 2760 -4140 3070 -4100
rect 3110 -4140 3420 -4100
rect 3460 -4140 3770 -4100
rect 3810 -4140 4120 -4100
rect 4160 -4140 4470 -4100
rect 4510 -4140 4820 -4100
rect 4860 -4140 5170 -4100
rect 5210 -4140 5520 -4100
rect 5560 -4140 5870 -4100
rect 5910 -4140 6220 -4100
rect 6260 -4140 6570 -4100
rect 6610 -4140 6920 -4100
rect 6960 -4140 7270 -4100
rect 7310 -4140 7620 -4100
rect 7660 -4140 7970 -4100
rect 8010 -4140 8320 -4100
rect 8360 -4140 8670 -4100
rect 8710 -4125 17990 -4100
rect 8710 -4140 14825 -4125
rect -120 -4165 14825 -4140
rect -120 -4205 -80 -4165
rect -40 -4205 270 -4165
rect 310 -4205 620 -4165
rect 660 -4205 970 -4165
rect 1010 -4205 1320 -4165
rect 1360 -4205 1670 -4165
rect 1710 -4205 2020 -4165
rect 2060 -4205 2370 -4165
rect 2410 -4205 2720 -4165
rect 2760 -4205 3070 -4165
rect 3110 -4205 3420 -4165
rect 3460 -4205 3770 -4165
rect 3810 -4205 4120 -4165
rect 4160 -4205 4470 -4165
rect 4510 -4205 4820 -4165
rect 4860 -4205 5170 -4165
rect 5210 -4205 5520 -4165
rect 5560 -4205 5870 -4165
rect 5910 -4205 6220 -4165
rect 6260 -4205 6570 -4165
rect 6610 -4205 6920 -4165
rect 6960 -4205 7270 -4165
rect 7310 -4205 7620 -4165
rect 7660 -4205 7970 -4165
rect 8010 -4205 8320 -4165
rect 8360 -4205 8670 -4165
rect 8710 -4175 14825 -4165
rect 14875 -4175 14920 -4125
rect 14970 -4175 15015 -4125
rect 15065 -4175 15115 -4125
rect 15165 -4175 15215 -4125
rect 15265 -4175 15315 -4125
rect 15365 -4175 15410 -4125
rect 15460 -4175 15505 -4125
rect 15555 -4175 15625 -4125
rect 15675 -4175 15720 -4125
rect 15770 -4175 15815 -4125
rect 15865 -4175 15915 -4125
rect 15965 -4175 16015 -4125
rect 16065 -4175 16115 -4125
rect 16165 -4175 16210 -4125
rect 16260 -4175 16305 -4125
rect 16355 -4175 16425 -4125
rect 16475 -4175 16520 -4125
rect 16570 -4175 16615 -4125
rect 16665 -4175 16715 -4125
rect 16765 -4175 16815 -4125
rect 16865 -4175 16915 -4125
rect 16965 -4175 17010 -4125
rect 17060 -4175 17105 -4125
rect 17155 -4175 17225 -4125
rect 17275 -4175 17320 -4125
rect 17370 -4175 17415 -4125
rect 17465 -4175 17515 -4125
rect 17565 -4175 17615 -4125
rect 17665 -4175 17715 -4125
rect 17765 -4175 17810 -4125
rect 17860 -4175 17905 -4125
rect 17955 -4175 17990 -4125
rect 8710 -4205 17990 -4175
rect -120 -4215 17990 -4205
rect -120 -4235 14825 -4215
rect -120 -4275 -80 -4235
rect -40 -4275 270 -4235
rect 310 -4275 620 -4235
rect 660 -4275 970 -4235
rect 1010 -4275 1320 -4235
rect 1360 -4275 1670 -4235
rect 1710 -4275 2020 -4235
rect 2060 -4275 2370 -4235
rect 2410 -4275 2720 -4235
rect 2760 -4275 3070 -4235
rect 3110 -4275 3420 -4235
rect 3460 -4275 3770 -4235
rect 3810 -4275 4120 -4235
rect 4160 -4275 4470 -4235
rect 4510 -4275 4820 -4235
rect 4860 -4275 5170 -4235
rect 5210 -4275 5520 -4235
rect 5560 -4275 5870 -4235
rect 5910 -4275 6220 -4235
rect 6260 -4275 6570 -4235
rect 6610 -4275 6920 -4235
rect 6960 -4275 7270 -4235
rect 7310 -4275 7620 -4235
rect 7660 -4275 7970 -4235
rect 8010 -4275 8320 -4235
rect 8360 -4275 8670 -4235
rect 8710 -4265 14825 -4235
rect 14875 -4265 14920 -4215
rect 14970 -4265 15015 -4215
rect 15065 -4265 15115 -4215
rect 15165 -4265 15215 -4215
rect 15265 -4265 15315 -4215
rect 15365 -4265 15410 -4215
rect 15460 -4265 15505 -4215
rect 15555 -4265 15625 -4215
rect 15675 -4265 15720 -4215
rect 15770 -4265 15815 -4215
rect 15865 -4265 15915 -4215
rect 15965 -4265 16015 -4215
rect 16065 -4265 16115 -4215
rect 16165 -4265 16210 -4215
rect 16260 -4265 16305 -4215
rect 16355 -4265 16425 -4215
rect 16475 -4265 16520 -4215
rect 16570 -4265 16615 -4215
rect 16665 -4265 16715 -4215
rect 16765 -4265 16815 -4215
rect 16865 -4265 16915 -4215
rect 16965 -4265 17010 -4215
rect 17060 -4265 17105 -4215
rect 17155 -4265 17225 -4215
rect 17275 -4265 17320 -4215
rect 17370 -4265 17415 -4215
rect 17465 -4265 17515 -4215
rect 17565 -4265 17615 -4215
rect 17665 -4265 17715 -4215
rect 17765 -4265 17810 -4215
rect 17860 -4265 17905 -4215
rect 17955 -4265 17990 -4215
rect 8710 -4275 17990 -4265
rect -120 -4305 17990 -4275
rect -120 -4345 -80 -4305
rect -40 -4345 270 -4305
rect 310 -4345 620 -4305
rect 660 -4345 970 -4305
rect 1010 -4345 1320 -4305
rect 1360 -4345 1670 -4305
rect 1710 -4345 2020 -4305
rect 2060 -4345 2370 -4305
rect 2410 -4345 2720 -4305
rect 2760 -4345 3070 -4305
rect 3110 -4345 3420 -4305
rect 3460 -4345 3770 -4305
rect 3810 -4345 4120 -4305
rect 4160 -4345 4470 -4305
rect 4510 -4345 4820 -4305
rect 4860 -4345 5170 -4305
rect 5210 -4345 5520 -4305
rect 5560 -4345 5870 -4305
rect 5910 -4345 6220 -4305
rect 6260 -4345 6570 -4305
rect 6610 -4345 6920 -4305
rect 6960 -4345 7270 -4305
rect 7310 -4345 7620 -4305
rect 7660 -4345 7970 -4305
rect 8010 -4345 8320 -4305
rect 8360 -4345 8670 -4305
rect 8710 -4315 17990 -4305
rect 8710 -4345 14825 -4315
rect -120 -4365 14825 -4345
rect 14875 -4365 14920 -4315
rect 14970 -4365 15015 -4315
rect 15065 -4365 15115 -4315
rect 15165 -4365 15215 -4315
rect 15265 -4365 15315 -4315
rect 15365 -4365 15410 -4315
rect 15460 -4365 15505 -4315
rect 15555 -4365 15625 -4315
rect 15675 -4365 15720 -4315
rect 15770 -4365 15815 -4315
rect 15865 -4365 15915 -4315
rect 15965 -4365 16015 -4315
rect 16065 -4365 16115 -4315
rect 16165 -4365 16210 -4315
rect 16260 -4365 16305 -4315
rect 16355 -4365 16425 -4315
rect 16475 -4365 16520 -4315
rect 16570 -4365 16615 -4315
rect 16665 -4365 16715 -4315
rect 16765 -4365 16815 -4315
rect 16865 -4365 16915 -4315
rect 16965 -4365 17010 -4315
rect 17060 -4365 17105 -4315
rect 17155 -4365 17225 -4315
rect 17275 -4365 17320 -4315
rect 17370 -4365 17415 -4315
rect 17465 -4365 17515 -4315
rect 17565 -4365 17615 -4315
rect 17665 -4365 17715 -4315
rect 17765 -4365 17810 -4315
rect 17860 -4365 17905 -4315
rect 17955 -4365 17990 -4315
rect -120 -4375 17990 -4365
rect -120 -4415 -80 -4375
rect -40 -4415 270 -4375
rect 310 -4415 620 -4375
rect 660 -4415 970 -4375
rect 1010 -4415 1320 -4375
rect 1360 -4415 1670 -4375
rect 1710 -4415 2020 -4375
rect 2060 -4415 2370 -4375
rect 2410 -4415 2720 -4375
rect 2760 -4415 3070 -4375
rect 3110 -4415 3420 -4375
rect 3460 -4415 3770 -4375
rect 3810 -4415 4120 -4375
rect 4160 -4415 4470 -4375
rect 4510 -4415 4820 -4375
rect 4860 -4415 5170 -4375
rect 5210 -4415 5520 -4375
rect 5560 -4415 5870 -4375
rect 5910 -4415 6220 -4375
rect 6260 -4415 6570 -4375
rect 6610 -4415 6920 -4375
rect 6960 -4415 7270 -4375
rect 7310 -4415 7620 -4375
rect 7660 -4415 7970 -4375
rect 8010 -4415 8320 -4375
rect 8360 -4415 8670 -4375
rect 8710 -4405 17990 -4375
rect 8710 -4415 14825 -4405
rect -120 -4440 14825 -4415
rect -120 -4480 -80 -4440
rect -40 -4480 270 -4440
rect 310 -4480 620 -4440
rect 660 -4480 970 -4440
rect 1010 -4480 1320 -4440
rect 1360 -4480 1670 -4440
rect 1710 -4480 2020 -4440
rect 2060 -4480 2370 -4440
rect 2410 -4480 2720 -4440
rect 2760 -4480 3070 -4440
rect 3110 -4480 3420 -4440
rect 3460 -4480 3770 -4440
rect 3810 -4480 4120 -4440
rect 4160 -4480 4470 -4440
rect 4510 -4480 4820 -4440
rect 4860 -4480 5170 -4440
rect 5210 -4480 5520 -4440
rect 5560 -4480 5870 -4440
rect 5910 -4480 6220 -4440
rect 6260 -4480 6570 -4440
rect 6610 -4480 6920 -4440
rect 6960 -4480 7270 -4440
rect 7310 -4480 7620 -4440
rect 7660 -4480 7970 -4440
rect 8010 -4480 8320 -4440
rect 8360 -4480 8670 -4440
rect 8710 -4455 14825 -4440
rect 14875 -4455 14920 -4405
rect 14970 -4455 15015 -4405
rect 15065 -4455 15115 -4405
rect 15165 -4455 15215 -4405
rect 15265 -4455 15315 -4405
rect 15365 -4455 15410 -4405
rect 15460 -4455 15505 -4405
rect 15555 -4455 15625 -4405
rect 15675 -4455 15720 -4405
rect 15770 -4455 15815 -4405
rect 15865 -4455 15915 -4405
rect 15965 -4455 16015 -4405
rect 16065 -4455 16115 -4405
rect 16165 -4455 16210 -4405
rect 16260 -4455 16305 -4405
rect 16355 -4455 16425 -4405
rect 16475 -4455 16520 -4405
rect 16570 -4455 16615 -4405
rect 16665 -4455 16715 -4405
rect 16765 -4455 16815 -4405
rect 16865 -4455 16915 -4405
rect 16965 -4455 17010 -4405
rect 17060 -4455 17105 -4405
rect 17155 -4455 17225 -4405
rect 17275 -4455 17320 -4405
rect 17370 -4455 17415 -4405
rect 17465 -4455 17515 -4405
rect 17565 -4455 17615 -4405
rect 17665 -4455 17715 -4405
rect 17765 -4455 17810 -4405
rect 17860 -4455 17905 -4405
rect 17955 -4455 17990 -4405
rect 8710 -4480 17990 -4455
rect -120 -4490 17990 -4480
use bgr_11  bgr_11_0
timestamp 1754058664
transform -1 0 22290 0 -1 11485
box 15665 -6150 19905 1755
use two_stage_opamp_dummy_magic_24  two_stage_opamp_dummy_magic_24_0
timestamp 1754061271
transform 1 0 -52410 0 1 100
box 52060 -1500 61740 6110
<< labels >>
flabel metal3 -2040 10155 -2040 10155 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 5375 1755 5375 1755 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 3605 1755 3605 1755 7 FreeSans 400 0 -160 0 VIN+
port 5 w
flabel metal2 6875 920 6875 920 5 FreeSans 400 0 0 -160 VOUT-
port 4 s
flabel metal2 2060 920 2060 920 5 FreeSans 400 0 0 -160 VOUT+
port 3 s
flabel metal4 20720 6650 20720 6650 3 FreeSans 800 0 320 0 GNDA
port 2 e
<< end >>
