magic
tech sky130A
timestamp 1738239539
<< nwell >>
rect 2765 -4430 3815 -3910
<< nmos >>
rect 2835 -4735 2850 -4685
rect 2900 -4735 2915 -4685
rect 2965 -4735 2980 -4685
rect 3030 -4735 3045 -4685
rect 3195 -4735 3210 -4685
rect 3260 -4735 3275 -4685
rect 3325 -4735 3340 -4685
rect 3390 -4735 3405 -4685
rect 3535 -4735 3550 -4685
rect 3600 -4735 3615 -4685
rect 3665 -4735 3680 -4685
rect 3730 -4735 3745 -4685
rect 3345 -5115 3395 -4865
rect 3445 -5115 3495 -4865
rect 3545 -5115 3595 -4865
rect 3645 -5115 3695 -4865
<< pmos >>
rect 2850 -4215 2900 -3965
rect 2950 -4215 3000 -3965
rect 3050 -4215 3100 -3965
rect 3150 -4215 3200 -3965
rect 3250 -4215 3300 -3965
rect 3350 -4215 3400 -3965
rect 3450 -4215 3500 -3965
rect 3550 -4215 3600 -3965
rect 2835 -4405 2850 -4305
rect 2900 -4405 2915 -4305
rect 2965 -4405 2980 -4305
rect 3030 -4405 3045 -4305
rect 3195 -4405 3210 -4305
rect 3260 -4405 3275 -4305
rect 3325 -4405 3340 -4305
rect 3390 -4405 3405 -4305
rect 3535 -4405 3550 -4305
rect 3600 -4405 3615 -4305
rect 3665 -4405 3680 -4305
rect 3730 -4405 3745 -4305
<< ndiff >>
rect 2785 -4700 2835 -4685
rect 2785 -4720 2800 -4700
rect 2820 -4720 2835 -4700
rect 2785 -4735 2835 -4720
rect 2850 -4700 2900 -4685
rect 2850 -4720 2865 -4700
rect 2885 -4720 2900 -4700
rect 2850 -4735 2900 -4720
rect 2915 -4700 2965 -4685
rect 2915 -4720 2930 -4700
rect 2950 -4720 2965 -4700
rect 2915 -4735 2965 -4720
rect 2980 -4700 3030 -4685
rect 2980 -4720 2995 -4700
rect 3015 -4720 3030 -4700
rect 2980 -4735 3030 -4720
rect 3045 -4700 3095 -4685
rect 3045 -4720 3060 -4700
rect 3080 -4720 3095 -4700
rect 3045 -4735 3095 -4720
rect 3145 -4700 3195 -4685
rect 3145 -4720 3160 -4700
rect 3180 -4720 3195 -4700
rect 3145 -4735 3195 -4720
rect 3210 -4700 3260 -4685
rect 3210 -4720 3225 -4700
rect 3245 -4720 3260 -4700
rect 3210 -4735 3260 -4720
rect 3275 -4700 3325 -4685
rect 3275 -4720 3290 -4700
rect 3310 -4720 3325 -4700
rect 3275 -4735 3325 -4720
rect 3340 -4700 3390 -4685
rect 3340 -4720 3355 -4700
rect 3375 -4720 3390 -4700
rect 3340 -4735 3390 -4720
rect 3405 -4700 3455 -4685
rect 3405 -4720 3420 -4700
rect 3440 -4720 3455 -4700
rect 3405 -4735 3455 -4720
rect 3485 -4700 3535 -4685
rect 3485 -4720 3500 -4700
rect 3520 -4720 3535 -4700
rect 3485 -4735 3535 -4720
rect 3550 -4700 3600 -4685
rect 3550 -4720 3565 -4700
rect 3585 -4720 3600 -4700
rect 3550 -4735 3600 -4720
rect 3615 -4700 3665 -4685
rect 3615 -4720 3630 -4700
rect 3650 -4720 3665 -4700
rect 3615 -4735 3665 -4720
rect 3680 -4700 3730 -4685
rect 3680 -4720 3695 -4700
rect 3715 -4720 3730 -4700
rect 3680 -4735 3730 -4720
rect 3745 -4700 3795 -4685
rect 3745 -4720 3760 -4700
rect 3780 -4720 3795 -4700
rect 3745 -4735 3795 -4720
rect 3295 -4880 3345 -4865
rect 3295 -5100 3310 -4880
rect 3330 -5100 3345 -4880
rect 3295 -5115 3345 -5100
rect 3395 -4880 3445 -4865
rect 3395 -5100 3410 -4880
rect 3430 -5100 3445 -4880
rect 3395 -5115 3445 -5100
rect 3495 -4880 3545 -4865
rect 3495 -5100 3510 -4880
rect 3530 -5100 3545 -4880
rect 3495 -5115 3545 -5100
rect 3595 -4880 3645 -4865
rect 3595 -5100 3610 -4880
rect 3630 -5100 3645 -4880
rect 3595 -5115 3645 -5100
rect 3695 -4880 3745 -4865
rect 3695 -5100 3710 -4880
rect 3730 -5100 3745 -4880
rect 3695 -5115 3745 -5100
<< pdiff >>
rect 2800 -3980 2850 -3965
rect 2800 -4200 2815 -3980
rect 2835 -4200 2850 -3980
rect 2800 -4215 2850 -4200
rect 2900 -3980 2950 -3965
rect 2900 -4200 2915 -3980
rect 2935 -4200 2950 -3980
rect 2900 -4215 2950 -4200
rect 3000 -3980 3050 -3965
rect 3000 -4200 3015 -3980
rect 3035 -4200 3050 -3980
rect 3000 -4215 3050 -4200
rect 3100 -3980 3150 -3965
rect 3100 -4200 3115 -3980
rect 3135 -4200 3150 -3980
rect 3100 -4215 3150 -4200
rect 3200 -3980 3250 -3965
rect 3200 -4200 3215 -3980
rect 3235 -4200 3250 -3980
rect 3200 -4215 3250 -4200
rect 3300 -3980 3350 -3965
rect 3300 -4200 3315 -3980
rect 3335 -4200 3350 -3980
rect 3300 -4215 3350 -4200
rect 3400 -3980 3450 -3965
rect 3400 -4200 3415 -3980
rect 3435 -4200 3450 -3980
rect 3400 -4215 3450 -4200
rect 3500 -3980 3550 -3965
rect 3500 -4200 3515 -3980
rect 3535 -4200 3550 -3980
rect 3500 -4215 3550 -4200
rect 3600 -3980 3650 -3965
rect 3600 -4200 3615 -3980
rect 3635 -4200 3650 -3980
rect 3600 -4215 3650 -4200
rect 2785 -4320 2835 -4305
rect 2785 -4390 2800 -4320
rect 2820 -4390 2835 -4320
rect 2785 -4405 2835 -4390
rect 2850 -4320 2900 -4305
rect 2850 -4390 2865 -4320
rect 2885 -4390 2900 -4320
rect 2850 -4405 2900 -4390
rect 2915 -4320 2965 -4305
rect 2915 -4390 2930 -4320
rect 2950 -4390 2965 -4320
rect 2915 -4405 2965 -4390
rect 2980 -4320 3030 -4305
rect 2980 -4390 2995 -4320
rect 3015 -4390 3030 -4320
rect 2980 -4405 3030 -4390
rect 3045 -4320 3095 -4305
rect 3045 -4390 3060 -4320
rect 3080 -4390 3095 -4320
rect 3045 -4405 3095 -4390
rect 3145 -4320 3195 -4305
rect 3145 -4390 3160 -4320
rect 3180 -4390 3195 -4320
rect 3145 -4405 3195 -4390
rect 3210 -4320 3260 -4305
rect 3210 -4390 3225 -4320
rect 3245 -4390 3260 -4320
rect 3210 -4405 3260 -4390
rect 3275 -4320 3325 -4305
rect 3275 -4390 3290 -4320
rect 3310 -4390 3325 -4320
rect 3275 -4405 3325 -4390
rect 3340 -4320 3390 -4305
rect 3340 -4390 3355 -4320
rect 3375 -4390 3390 -4320
rect 3340 -4405 3390 -4390
rect 3405 -4320 3455 -4305
rect 3405 -4390 3420 -4320
rect 3440 -4390 3455 -4320
rect 3405 -4405 3455 -4390
rect 3485 -4320 3535 -4305
rect 3485 -4390 3500 -4320
rect 3520 -4390 3535 -4320
rect 3485 -4405 3535 -4390
rect 3550 -4320 3600 -4305
rect 3550 -4390 3565 -4320
rect 3585 -4390 3600 -4320
rect 3550 -4405 3600 -4390
rect 3615 -4320 3665 -4305
rect 3615 -4390 3630 -4320
rect 3650 -4390 3665 -4320
rect 3615 -4405 3665 -4390
rect 3680 -4320 3730 -4305
rect 3680 -4390 3695 -4320
rect 3715 -4390 3730 -4320
rect 3680 -4405 3730 -4390
rect 3745 -4320 3795 -4305
rect 3745 -4390 3760 -4320
rect 3780 -4390 3795 -4320
rect 3745 -4405 3795 -4390
<< ndiffc >>
rect 2800 -4720 2820 -4700
rect 2865 -4720 2885 -4700
rect 2930 -4720 2950 -4700
rect 2995 -4720 3015 -4700
rect 3060 -4720 3080 -4700
rect 3160 -4720 3180 -4700
rect 3225 -4720 3245 -4700
rect 3290 -4720 3310 -4700
rect 3355 -4720 3375 -4700
rect 3420 -4720 3440 -4700
rect 3500 -4720 3520 -4700
rect 3565 -4720 3585 -4700
rect 3630 -4720 3650 -4700
rect 3695 -4720 3715 -4700
rect 3760 -4720 3780 -4700
rect 3310 -5100 3330 -4880
rect 3410 -5100 3430 -4880
rect 3510 -5100 3530 -4880
rect 3610 -5100 3630 -4880
rect 3710 -5100 3730 -4880
<< pdiffc >>
rect 2815 -4200 2835 -3980
rect 2915 -4200 2935 -3980
rect 3015 -4200 3035 -3980
rect 3115 -4200 3135 -3980
rect 3215 -4200 3235 -3980
rect 3315 -4200 3335 -3980
rect 3415 -4200 3435 -3980
rect 3515 -4200 3535 -3980
rect 3615 -4200 3635 -3980
rect 2800 -4390 2820 -4320
rect 2865 -4390 2885 -4320
rect 2930 -4390 2950 -4320
rect 2995 -4390 3015 -4320
rect 3060 -4390 3080 -4320
rect 3160 -4390 3180 -4320
rect 3225 -4390 3245 -4320
rect 3290 -4390 3310 -4320
rect 3355 -4390 3375 -4320
rect 3420 -4390 3440 -4320
rect 3500 -4390 3520 -4320
rect 3565 -4390 3585 -4320
rect 3630 -4390 3650 -4320
rect 3695 -4390 3715 -4320
rect 3760 -4390 3780 -4320
<< psubdiff >>
rect 2915 -4780 2965 -4765
rect 2915 -4800 2930 -4780
rect 2950 -4800 2965 -4780
rect 2915 -4815 2965 -4800
rect 2975 -5250 3025 -5200
<< nsubdiff >>
rect 3695 -3980 3745 -3965
rect 3695 -4200 3710 -3980
rect 3730 -4200 3745 -3980
rect 3695 -4215 3745 -4200
<< psubdiffcont >>
rect 2930 -4800 2950 -4780
<< nsubdiffcont >>
rect 3710 -4200 3730 -3980
<< poly >>
rect 2255 -3690 2415 -3675
rect 2255 -4170 2310 -4160
rect 2255 -4175 2280 -4170
rect 2270 -4190 2280 -4175
rect 2300 -4190 2310 -4170
rect 2270 -4200 2310 -4190
rect 2400 -4280 2415 -3690
rect 2830 -3920 2870 -3910
rect 2830 -3940 2840 -3920
rect 2860 -3940 2870 -3920
rect 3205 -3920 3245 -3910
rect 3205 -3940 3215 -3920
rect 3235 -3940 3245 -3920
rect 3585 -3920 3625 -3910
rect 3585 -3940 3595 -3920
rect 3615 -3940 3625 -3920
rect 2830 -3950 3625 -3940
rect 2850 -3955 3600 -3950
rect 2850 -3965 2900 -3955
rect 2950 -3965 3000 -3955
rect 3050 -3965 3100 -3955
rect 3150 -3965 3200 -3955
rect 3250 -3965 3300 -3955
rect 3350 -3965 3400 -3955
rect 3450 -3965 3500 -3955
rect 3550 -3965 3600 -3955
rect 2850 -4230 2900 -4215
rect 2950 -4230 3000 -4215
rect 3050 -4230 3100 -4215
rect 3150 -4230 3200 -4215
rect 3250 -4230 3300 -4215
rect 3350 -4230 3400 -4215
rect 3450 -4230 3500 -4215
rect 3550 -4230 3600 -4215
rect 2400 -4295 2915 -4280
rect 2430 -4440 2470 -4430
rect 2430 -4455 2440 -4440
rect 2255 -4460 2440 -4455
rect 2460 -4460 2470 -4440
rect 2255 -4470 2470 -4460
rect 2525 -4590 2540 -4295
rect 2835 -4305 2850 -4295
rect 2900 -4305 2915 -4295
rect 2965 -4305 2980 -4290
rect 3030 -4305 3045 -4290
rect 3195 -4305 3210 -4290
rect 3260 -4305 3275 -4290
rect 3325 -4305 3340 -4290
rect 3390 -4305 3405 -4290
rect 3535 -4305 3550 -4290
rect 3600 -4305 3615 -4290
rect 3665 -4305 3680 -4290
rect 3730 -4305 3745 -4290
rect 2835 -4420 2850 -4405
rect 2900 -4420 2915 -4405
rect 2590 -4440 2630 -4430
rect 2590 -4460 2600 -4440
rect 2620 -4445 2630 -4440
rect 2965 -4445 2980 -4405
rect 3030 -4445 3045 -4405
rect 3195 -4415 3210 -4405
rect 3260 -4415 3275 -4405
rect 3325 -4415 3340 -4405
rect 3390 -4415 3405 -4405
rect 3195 -4420 3405 -4415
rect 3535 -4415 3550 -4405
rect 3600 -4415 3615 -4405
rect 3665 -4415 3680 -4405
rect 3730 -4415 3745 -4405
rect 3165 -4430 3440 -4420
rect 2620 -4455 3140 -4445
rect 2620 -4460 3110 -4455
rect 2590 -4470 2630 -4460
rect 3100 -4475 3110 -4460
rect 3130 -4475 3140 -4455
rect 3165 -4450 3175 -4430
rect 3195 -4435 3410 -4430
rect 3195 -4450 3205 -4435
rect 3165 -4460 3205 -4450
rect 3400 -4450 3410 -4435
rect 3430 -4450 3440 -4430
rect 3400 -4460 3440 -4450
rect 3535 -4430 3885 -4415
rect 3535 -4450 3545 -4430
rect 3565 -4450 3575 -4430
rect 3535 -4460 3575 -4450
rect 3100 -4485 3140 -4475
rect 2930 -4535 2970 -4525
rect 2930 -4555 2940 -4535
rect 2960 -4550 2970 -4535
rect 2960 -4555 3550 -4550
rect 2930 -4565 3550 -4555
rect 2525 -4605 3275 -4590
rect 2800 -4640 2840 -4630
rect 2800 -4660 2810 -4640
rect 2830 -4655 2840 -4640
rect 3040 -4640 3080 -4630
rect 3040 -4655 3050 -4640
rect 2830 -4660 3050 -4655
rect 3070 -4660 3080 -4640
rect 2800 -4670 3080 -4660
rect 2835 -4675 3045 -4670
rect 2835 -4685 2850 -4675
rect 2900 -4685 2915 -4675
rect 2965 -4685 2980 -4675
rect 3030 -4685 3045 -4675
rect 3195 -4685 3210 -4605
rect 3260 -4685 3275 -4605
rect 3535 -4660 3550 -4565
rect 3325 -4685 3340 -4670
rect 3390 -4685 3405 -4670
rect 3535 -4675 3845 -4660
rect 3535 -4685 3550 -4675
rect 3600 -4685 3615 -4675
rect 3665 -4685 3680 -4675
rect 3730 -4685 3745 -4675
rect 2835 -4750 2850 -4735
rect 2900 -4750 2915 -4735
rect 2965 -4750 2980 -4735
rect 3030 -4750 3045 -4735
rect 3195 -4750 3210 -4735
rect 3260 -4750 3275 -4735
rect 3090 -4770 3130 -4760
rect 3090 -4790 3100 -4770
rect 3120 -4775 3130 -4770
rect 3325 -4775 3340 -4735
rect 3390 -4775 3405 -4735
rect 3535 -4750 3550 -4735
rect 3600 -4750 3615 -4735
rect 3665 -4750 3680 -4735
rect 3730 -4750 3745 -4735
rect 3120 -4790 3405 -4775
rect 3090 -4800 3130 -4790
rect 3345 -4865 3395 -4850
rect 3445 -4865 3495 -4850
rect 3545 -4865 3595 -4850
rect 3645 -4865 3695 -4850
rect 3345 -5125 3395 -5115
rect 3445 -5125 3495 -5115
rect 3545 -5125 3595 -5115
rect 3645 -5125 3695 -5115
rect 3345 -5135 3695 -5125
rect 3345 -5140 3360 -5135
rect 3350 -5155 3360 -5140
rect 3380 -5140 3660 -5135
rect 3380 -5155 3390 -5140
rect 3350 -5165 3390 -5155
rect 3650 -5155 3660 -5140
rect 3680 -5140 3695 -5135
rect 3680 -5155 3690 -5140
rect 3650 -5165 3690 -5155
rect 3830 -5295 3845 -4675
rect 3450 -5310 3845 -5295
rect 3260 -5406 3300 -5396
rect 3260 -5426 3270 -5406
rect 3290 -5421 3300 -5406
rect 3450 -5421 3465 -5310
rect 3870 -5335 3885 -4430
rect 3695 -5350 3885 -5335
rect 3695 -5396 3710 -5350
rect 3290 -5426 3465 -5421
rect 3260 -5436 3465 -5426
rect 3690 -5406 3730 -5396
rect 3690 -5426 3700 -5406
rect 3720 -5426 3730 -5406
rect 3690 -5436 3730 -5426
<< polycont >>
rect 2280 -4190 2300 -4170
rect 2840 -3940 2860 -3920
rect 3215 -3940 3235 -3920
rect 3595 -3940 3615 -3920
rect 2440 -4460 2460 -4440
rect 2600 -4460 2620 -4440
rect 3110 -4475 3130 -4455
rect 3175 -4450 3195 -4430
rect 3410 -4450 3430 -4430
rect 3545 -4450 3565 -4430
rect 2940 -4555 2960 -4535
rect 2810 -4660 2830 -4640
rect 3050 -4660 3070 -4640
rect 3100 -4790 3120 -4770
rect 3360 -5155 3380 -5135
rect 3660 -5155 3680 -5135
rect 3270 -5426 3290 -5406
rect 3700 -5426 3720 -5406
<< xpolycontact >>
rect 2765 -5150 2985 -4865
rect 3020 -5150 3240 -4865
rect 2635 -5436 2855 -5401
rect 2925 -5436 3145 -5401
rect 3780 -5436 4000 -5401
rect 4098 -5436 4318 -5401
<< xpolyres >>
rect 2985 -5150 3020 -4865
rect 2855 -5436 2925 -5401
rect 4000 -5436 4098 -5401
<< locali >>
rect 2495 -3640 3245 -3620
rect 2270 -4170 2310 -4160
rect 2270 -4190 2280 -4170
rect 2300 -4190 2310 -4170
rect 2270 -4200 2310 -4190
rect 2290 -5540 2310 -4200
rect 2430 -4440 2470 -4430
rect 2430 -4460 2440 -4440
rect 2460 -4450 2470 -4440
rect 2495 -4450 2515 -3640
rect 2830 -3920 2870 -3910
rect 2830 -3925 2840 -3920
rect 2695 -3940 2840 -3925
rect 2860 -3925 2870 -3920
rect 3205 -3920 3245 -3910
rect 3205 -3925 3215 -3920
rect 2860 -3940 3215 -3925
rect 3235 -3925 3245 -3920
rect 3585 -3920 3625 -3910
rect 3585 -3925 3595 -3920
rect 3235 -3940 3595 -3925
rect 3615 -3925 3625 -3920
rect 3615 -3940 3635 -3925
rect 2695 -3945 3635 -3940
rect 2590 -4440 2630 -4430
rect 2590 -4450 2600 -4440
rect 2460 -4460 2600 -4450
rect 2620 -4460 2630 -4440
rect 2430 -4470 2630 -4460
rect 2695 -4865 2715 -3945
rect 2815 -3950 2870 -3945
rect 3205 -3950 3245 -3945
rect 3585 -3950 3635 -3945
rect 2815 -3970 2835 -3950
rect 3215 -3970 3235 -3950
rect 3615 -3970 3635 -3950
rect 2800 -3980 2845 -3970
rect 2800 -4200 2815 -3980
rect 2835 -4200 2845 -3980
rect 2800 -4210 2845 -4200
rect 2905 -3980 2945 -3970
rect 2905 -4200 2915 -3980
rect 2935 -4200 2945 -3980
rect 2905 -4210 2945 -4200
rect 3005 -3980 3045 -3970
rect 3005 -4200 3015 -3980
rect 3035 -4200 3045 -3980
rect 3005 -4210 3045 -4200
rect 3105 -3980 3145 -3970
rect 3105 -4200 3115 -3980
rect 3135 -4200 3145 -3980
rect 3105 -4210 3145 -4200
rect 3205 -3980 3245 -3970
rect 3205 -4200 3215 -3980
rect 3235 -4200 3245 -3980
rect 3205 -4210 3245 -4200
rect 3305 -3980 3345 -3970
rect 3305 -4200 3315 -3980
rect 3335 -4200 3345 -3980
rect 3305 -4210 3345 -4200
rect 3405 -3980 3445 -3970
rect 3405 -4200 3415 -3980
rect 3435 -4200 3445 -3980
rect 3405 -4210 3445 -4200
rect 3505 -3980 3545 -3970
rect 3505 -4200 3515 -3980
rect 3535 -4200 3545 -3980
rect 3505 -4210 3545 -4200
rect 3605 -3980 3645 -3970
rect 3605 -4200 3615 -3980
rect 3635 -4200 3645 -3980
rect 3605 -4210 3645 -4200
rect 3700 -3980 3740 -3970
rect 3700 -4200 3710 -3980
rect 3730 -4200 3740 -3980
rect 3700 -4210 3740 -4200
rect 3015 -4230 3035 -4210
rect 3415 -4230 3435 -4210
rect 2880 -4250 3435 -4230
rect 2880 -4270 2900 -4250
rect 2800 -4290 3080 -4270
rect 2800 -4310 2820 -4290
rect 2930 -4310 2950 -4290
rect 3060 -4310 3080 -4290
rect 3500 -4290 3780 -4270
rect 3500 -4310 3520 -4290
rect 3630 -4310 3650 -4290
rect 3760 -4310 3780 -4290
rect 2790 -4320 2830 -4310
rect 2790 -4390 2800 -4320
rect 2820 -4390 2830 -4320
rect 2790 -4400 2830 -4390
rect 2855 -4320 2895 -4310
rect 2855 -4390 2865 -4320
rect 2885 -4390 2895 -4320
rect 2855 -4400 2895 -4390
rect 2920 -4320 2960 -4310
rect 2920 -4390 2930 -4320
rect 2950 -4390 2960 -4320
rect 2920 -4400 2960 -4390
rect 2985 -4320 3025 -4310
rect 2985 -4390 2995 -4320
rect 3015 -4390 3025 -4320
rect 2985 -4400 3025 -4390
rect 3050 -4320 3095 -4310
rect 3050 -4390 3060 -4320
rect 3080 -4390 3095 -4320
rect 3050 -4400 3095 -4390
rect 3150 -4320 3190 -4310
rect 3150 -4390 3160 -4320
rect 3180 -4390 3190 -4320
rect 3150 -4400 3190 -4390
rect 3215 -4320 3255 -4310
rect 3215 -4390 3225 -4320
rect 3245 -4390 3255 -4320
rect 3215 -4400 3255 -4390
rect 3280 -4320 3320 -4310
rect 3280 -4390 3290 -4320
rect 3310 -4390 3320 -4320
rect 3280 -4400 3320 -4390
rect 3345 -4320 3390 -4310
rect 3345 -4390 3355 -4320
rect 3375 -4390 3390 -4320
rect 3345 -4400 3390 -4390
rect 3410 -4320 3450 -4310
rect 3410 -4390 3420 -4320
rect 3440 -4390 3450 -4320
rect 3410 -4400 3450 -4390
rect 3490 -4320 3530 -4310
rect 3490 -4390 3500 -4320
rect 3520 -4390 3530 -4320
rect 3490 -4400 3530 -4390
rect 3555 -4320 3595 -4310
rect 3555 -4390 3565 -4320
rect 3585 -4390 3595 -4320
rect 3555 -4400 3595 -4390
rect 3620 -4320 3660 -4310
rect 3620 -4390 3630 -4320
rect 3650 -4390 3660 -4320
rect 3620 -4400 3660 -4390
rect 3685 -4320 3725 -4310
rect 3685 -4390 3695 -4320
rect 3715 -4390 3725 -4320
rect 3685 -4400 3725 -4390
rect 3750 -4320 3790 -4310
rect 3750 -4390 3760 -4320
rect 3780 -4390 3790 -4320
rect 3750 -4400 3790 -4390
rect 2865 -4485 2885 -4400
rect 2995 -4485 3015 -4400
rect 3160 -4420 3185 -4400
rect 3165 -4430 3205 -4420
rect 3100 -4455 3140 -4445
rect 3100 -4475 3110 -4455
rect 3130 -4475 3140 -4455
rect 3165 -4450 3175 -4430
rect 3195 -4450 3205 -4430
rect 3165 -4460 3205 -4450
rect 3100 -4485 3140 -4475
rect 3170 -4485 3190 -4460
rect 2810 -4510 2885 -4485
rect 2940 -4505 3015 -4485
rect 2810 -4630 2830 -4510
rect 2940 -4525 2960 -4505
rect 2930 -4535 2970 -4525
rect 2930 -4555 2940 -4535
rect 2960 -4555 2970 -4535
rect 2930 -4565 2970 -4555
rect 2800 -4640 2840 -4630
rect 2800 -4660 2810 -4640
rect 2830 -4660 2840 -4640
rect 2800 -4670 2840 -4660
rect 2800 -4690 2820 -4670
rect 2930 -4690 2950 -4565
rect 3040 -4640 3080 -4630
rect 3040 -4660 3050 -4640
rect 3070 -4660 3080 -4640
rect 3040 -4670 3080 -4660
rect 3060 -4690 3080 -4670
rect 2790 -4700 2830 -4690
rect 2790 -4720 2800 -4700
rect 2820 -4720 2830 -4700
rect 2790 -4730 2830 -4720
rect 2855 -4700 2895 -4690
rect 2855 -4720 2865 -4700
rect 2885 -4720 2895 -4700
rect 2855 -4730 2895 -4720
rect 2920 -4700 2960 -4690
rect 2920 -4720 2930 -4700
rect 2950 -4720 2960 -4700
rect 2920 -4730 2960 -4720
rect 2985 -4700 3025 -4690
rect 2985 -4720 2995 -4700
rect 3015 -4720 3025 -4700
rect 2985 -4730 3025 -4720
rect 3050 -4700 3090 -4690
rect 3050 -4720 3060 -4700
rect 3080 -4720 3090 -4700
rect 3050 -4730 3090 -4720
rect 2865 -4780 2885 -4730
rect 2920 -4780 2960 -4770
rect 2995 -4780 3015 -4730
rect 3110 -4760 3130 -4485
rect 3170 -4505 3245 -4485
rect 3225 -4690 3245 -4505
rect 3290 -4495 3310 -4400
rect 3420 -4420 3440 -4400
rect 3760 -4420 3780 -4400
rect 3400 -4430 3440 -4420
rect 3400 -4450 3410 -4430
rect 3430 -4450 3440 -4430
rect 3400 -4460 3440 -4450
rect 3535 -4430 3575 -4420
rect 3535 -4450 3545 -4430
rect 3565 -4450 3575 -4430
rect 3760 -4440 3895 -4420
rect 3535 -4460 3575 -4450
rect 3535 -4495 3555 -4460
rect 3290 -4515 3555 -4495
rect 3355 -4690 3375 -4515
rect 3150 -4700 3190 -4690
rect 3150 -4720 3160 -4700
rect 3180 -4720 3190 -4700
rect 3150 -4730 3190 -4720
rect 3215 -4700 3255 -4690
rect 3215 -4720 3225 -4700
rect 3245 -4720 3255 -4700
rect 3215 -4730 3255 -4720
rect 3280 -4700 3320 -4690
rect 3280 -4720 3290 -4700
rect 3310 -4720 3320 -4700
rect 3280 -4730 3320 -4720
rect 3345 -4700 3385 -4690
rect 3345 -4720 3355 -4700
rect 3375 -4720 3385 -4700
rect 3345 -4730 3385 -4720
rect 3410 -4700 3450 -4690
rect 3410 -4720 3420 -4700
rect 3440 -4720 3450 -4700
rect 3410 -4730 3450 -4720
rect 3490 -4700 3530 -4690
rect 3490 -4720 3500 -4700
rect 3520 -4720 3530 -4700
rect 3490 -4730 3530 -4720
rect 3555 -4700 3595 -4690
rect 3555 -4720 3565 -4700
rect 3585 -4720 3595 -4700
rect 3555 -4730 3595 -4720
rect 3620 -4700 3660 -4690
rect 3620 -4720 3630 -4700
rect 3650 -4720 3660 -4700
rect 3620 -4730 3660 -4720
rect 3685 -4700 3725 -4690
rect 3685 -4720 3695 -4700
rect 3715 -4720 3725 -4700
rect 3685 -4730 3725 -4720
rect 3750 -4700 3790 -4690
rect 3750 -4720 3760 -4700
rect 3780 -4720 3790 -4700
rect 3750 -4730 3790 -4720
rect 2865 -4800 2930 -4780
rect 2950 -4800 3015 -4780
rect 3090 -4770 3130 -4760
rect 3160 -4750 3180 -4730
rect 3290 -4750 3310 -4730
rect 3420 -4750 3440 -4730
rect 3160 -4770 3440 -4750
rect 3500 -4750 3520 -4730
rect 3630 -4750 3650 -4730
rect 3760 -4750 3780 -4730
rect 3500 -4755 3780 -4750
rect 3090 -4790 3100 -4770
rect 3120 -4790 3130 -4770
rect 3090 -4800 3130 -4790
rect 2920 -4810 2960 -4800
rect 3290 -4830 3310 -4770
rect 3500 -4775 3855 -4755
rect 3290 -4850 3530 -4830
rect 2695 -4885 2765 -4865
rect 3510 -4870 3530 -4850
rect 3300 -4880 3340 -4870
rect 3300 -5100 3310 -4880
rect 3330 -5100 3340 -4880
rect 3300 -5110 3340 -5100
rect 3400 -4880 3440 -4870
rect 3400 -5100 3410 -4880
rect 3430 -5100 3440 -4880
rect 3400 -5110 3440 -5100
rect 3500 -4880 3540 -4870
rect 3500 -5100 3510 -4880
rect 3530 -5100 3540 -4880
rect 3500 -5110 3540 -5100
rect 3600 -4880 3640 -4870
rect 3600 -5100 3610 -4880
rect 3630 -5100 3640 -4880
rect 3600 -5110 3640 -5100
rect 3700 -4880 3740 -4870
rect 3700 -5100 3710 -4880
rect 3730 -5100 3740 -4880
rect 3700 -5110 3740 -5100
rect 3310 -5130 3330 -5110
rect 3350 -5130 3390 -5125
rect 3650 -5130 3690 -5125
rect 3710 -5130 3730 -5110
rect 3240 -5135 3730 -5130
rect 3240 -5150 3360 -5135
rect 3350 -5155 3360 -5150
rect 3380 -5150 3660 -5135
rect 3380 -5155 3390 -5150
rect 3350 -5165 3390 -5155
rect 3650 -5155 3660 -5150
rect 3680 -5150 3730 -5135
rect 3680 -5155 3690 -5150
rect 3650 -5165 3690 -5155
rect 2980 -5215 3020 -5205
rect 2980 -5235 2990 -5215
rect 3010 -5235 3020 -5215
rect 2980 -5245 3020 -5235
rect 3835 -5315 3855 -4775
rect 3495 -5335 3855 -5315
rect 2440 -5436 2635 -5416
rect 3260 -5406 3300 -5396
rect 3260 -5416 3270 -5406
rect 3145 -5426 3270 -5416
rect 3290 -5426 3300 -5406
rect 3145 -5436 3300 -5426
rect 2440 -5456 2460 -5436
rect 3495 -5456 3515 -5335
rect 3875 -5355 3895 -4440
rect 2420 -5466 2470 -5456
rect 2420 -5496 2430 -5466
rect 2460 -5496 2470 -5466
rect 2420 -5506 2470 -5496
rect 3385 -5466 3515 -5456
rect 3385 -5501 3395 -5466
rect 3430 -5476 3515 -5466
rect 3430 -5501 3440 -5476
rect 3385 -5511 3440 -5501
rect 3495 -5540 3515 -5476
rect 3575 -5375 3895 -5355
rect 3575 -5456 3595 -5375
rect 3690 -5401 3730 -5396
rect 3690 -5406 3780 -5401
rect 3690 -5426 3700 -5406
rect 3720 -5421 3780 -5406
rect 3720 -5426 3730 -5421
rect 3690 -5436 3730 -5426
rect 4318 -5436 4635 -5416
rect 4615 -5456 4635 -5436
rect 3575 -5466 3690 -5456
rect 3575 -5476 3645 -5466
rect 3575 -5540 3595 -5476
rect 3635 -5501 3645 -5476
rect 3680 -5501 3690 -5466
rect 3635 -5511 3690 -5501
rect 4605 -5466 4655 -5456
rect 4605 -5496 4615 -5466
rect 4645 -5496 4655 -5466
rect 4605 -5506 4655 -5496
rect 2290 -5560 3595 -5540
<< viali >>
rect 2915 -4200 2935 -3980
rect 3115 -4200 3135 -3980
rect 3315 -4200 3335 -3980
rect 3515 -4200 3535 -3980
rect 3710 -4200 3730 -3980
rect 3225 -4390 3245 -4320
rect 3355 -4390 3375 -4320
rect 3565 -4390 3585 -4320
rect 3695 -4390 3715 -4320
rect 2865 -4720 2885 -4700
rect 2995 -4720 3015 -4700
rect 3565 -4720 3585 -4700
rect 3695 -4720 3715 -4700
rect 2930 -4800 2950 -4780
rect 3410 -5100 3430 -4880
rect 3610 -5100 3630 -4880
rect 2990 -5235 3010 -5215
rect 2430 -5496 2460 -5466
rect 3395 -5501 3430 -5466
rect 3645 -5501 3680 -5466
rect 4615 -5496 4645 -5466
<< metal1 >>
rect 2255 -3910 2915 -3845
rect 2255 -3980 3815 -3910
rect 2255 -4200 2915 -3980
rect 2935 -4200 3115 -3980
rect 3135 -4200 3315 -3980
rect 3335 -4200 3515 -3980
rect 3535 -4200 3710 -3980
rect 3730 -4200 3815 -3980
rect 2255 -4320 3815 -4200
rect 2255 -4390 3225 -4320
rect 3245 -4390 3355 -4320
rect 3375 -4390 3565 -4320
rect 3585 -4390 3695 -4320
rect 3715 -4390 3815 -4320
rect 2255 -4430 3815 -4390
rect 2255 -4480 2915 -4430
rect 2255 -4645 2915 -4610
rect 2255 -4700 3815 -4645
rect 2255 -4720 2865 -4700
rect 2885 -4720 2995 -4700
rect 3015 -4720 3565 -4700
rect 3585 -4720 3695 -4700
rect 3715 -4720 3815 -4700
rect 2255 -4780 3815 -4720
rect 2255 -4800 2930 -4780
rect 2950 -4800 3815 -4780
rect 2255 -4880 3815 -4800
rect 2255 -4965 3410 -4880
rect 2745 -5100 3410 -4965
rect 3430 -5100 3610 -4880
rect 3630 -5100 3815 -4880
rect 2745 -5215 3815 -5100
rect 2745 -5235 2990 -5215
rect 3010 -5235 3815 -5215
rect 2745 -5275 3815 -5235
rect 2420 -5466 2470 -5456
rect 2420 -5496 2430 -5466
rect 2460 -5496 2470 -5466
rect 2420 -5506 2470 -5496
rect 3385 -5466 3440 -5456
rect 3385 -5501 3395 -5466
rect 3430 -5501 3440 -5466
rect 3385 -5511 3440 -5501
rect 3635 -5466 3690 -5456
rect 3635 -5501 3645 -5466
rect 3680 -5501 3690 -5466
rect 3635 -5511 3690 -5501
rect 4605 -5466 4655 -5456
rect 4605 -5496 4615 -5466
rect 4645 -5496 4655 -5466
rect 4605 -5506 4655 -5496
<< via1 >>
rect 2430 -5496 2460 -5466
rect 3395 -5501 3430 -5466
rect 3645 -5501 3680 -5466
rect 4615 -5496 4645 -5466
<< metal2 >>
rect 2420 -5466 2470 -5456
rect 2420 -5496 2430 -5466
rect 2460 -5496 2470 -5466
rect 2420 -5506 2470 -5496
rect 3385 -5466 3440 -5456
rect 3385 -5501 3395 -5466
rect 3430 -5501 3440 -5466
rect 3385 -5511 3440 -5501
rect 3635 -5466 3690 -5456
rect 3635 -5501 3645 -5466
rect 3680 -5501 3690 -5466
rect 3635 -5511 3690 -5501
rect 4605 -5466 4655 -5456
rect 4605 -5496 4615 -5466
rect 4645 -5496 4655 -5466
rect 4605 -5506 4655 -5496
<< via2 >>
rect 2430 -5496 2460 -5466
rect 3395 -5501 3430 -5466
rect 3645 -5501 3680 -5466
rect 4615 -5496 4645 -5466
<< metal3 >>
rect 2420 -5466 2470 -5456
rect 2420 -5496 2430 -5466
rect 2460 -5496 2470 -5466
rect 2420 -5506 2470 -5496
rect 2425 -5631 2470 -5506
rect 3385 -5466 3440 -5456
rect 3385 -5501 3395 -5466
rect 3430 -5501 3440 -5466
rect 3385 -5511 3440 -5501
rect 3635 -5466 3690 -5456
rect 3635 -5501 3645 -5466
rect 3680 -5501 3690 -5466
rect 3635 -5511 3690 -5501
rect 4605 -5466 4655 -5456
rect 4605 -5496 4615 -5466
rect 4645 -5496 4655 -5466
rect 4605 -5506 4655 -5496
rect 4605 -5631 4650 -5506
rect 2425 -6661 3455 -5631
rect 3620 -6661 4650 -5631
<< via3 >>
rect 3395 -5501 3430 -5466
rect 3645 -5501 3680 -5466
<< mimcap >>
rect 2440 -5656 3440 -5646
rect 2440 -5691 3395 -5656
rect 3430 -5691 3440 -5656
rect 2440 -6646 3440 -5691
rect 3635 -5656 4635 -5646
rect 3635 -5691 3645 -5656
rect 3680 -5691 4635 -5656
rect 3635 -6646 4635 -5691
<< mimcapcontact >>
rect 3395 -5691 3430 -5656
rect 3645 -5691 3680 -5656
<< metal4 >>
rect 3385 -5466 3440 -5456
rect 3385 -5501 3395 -5466
rect 3430 -5501 3440 -5466
rect 3385 -5656 3440 -5501
rect 3385 -5691 3395 -5656
rect 3430 -5691 3440 -5656
rect 3385 -5696 3440 -5691
rect 3635 -5466 3690 -5456
rect 3635 -5501 3645 -5466
rect 3680 -5501 3690 -5466
rect 3635 -5656 3690 -5501
rect 3635 -5691 3645 -5656
rect 3680 -5691 3690 -5656
rect 3635 -5696 3690 -5691
<< labels >>
flabel locali 3530 -4830 3530 -4830 2 FreeSans 400 0 0 0 v_common_n
flabel locali 3435 -4250 3435 -4250 4 FreeSans 400 0 0 0 v_common_p
flabel locali 3245 -4530 3245 -4530 3 FreeSans 160 0 80 0 n_left
flabel locali 3375 -4530 3375 -4530 3 FreeSans 160 0 80 0 n_right
flabel locali 3015 -4505 3015 -4505 3 FreeSans 160 0 80 0 p_right
flabel locali 2810 -4510 2810 -4510 7 FreeSans 160 0 -80 0 p_left
flabel locali 3290 -5150 3290 -5150 5 FreeSans 160 0 0 -80 n_bias
flabel locali 2695 -4050 2695 -4050 7 FreeSans 160 0 -80 0 p_bias
<< end >>
