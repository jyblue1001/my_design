magic
tech sky130A
timestamp 1739021450
<< nwell >>
rect 8350 2165 10840 2355
<< nmos >>
rect 8530 1905 8590 2005
rect 8640 1905 8700 2005
rect 8750 1905 8810 2005
rect 8860 1905 8920 2005
rect 8970 1905 9030 2005
rect 9080 1905 9140 2005
rect 9290 1905 9350 2005
rect 9400 1905 9460 2005
rect 9510 1905 9570 2005
rect 9620 1905 9680 2005
rect 9730 1905 9790 2005
rect 9840 1905 9900 2005
rect 10050 1905 10110 2005
rect 10160 1905 10220 2005
rect 10270 1905 10330 2005
rect 10380 1905 10440 2005
rect 10490 1905 10550 2005
rect 10600 1905 10660 2005
<< pmos >>
rect 8470 2235 8530 2335
rect 8580 2235 8640 2335
rect 8690 2235 8750 2335
rect 8800 2235 8860 2335
rect 8910 2235 8970 2335
rect 9020 2235 9080 2335
rect 9130 2235 9190 2335
rect 9240 2235 9300 2335
rect 9350 2235 9410 2335
rect 9460 2235 9520 2335
rect 9670 2235 9730 2335
rect 9780 2235 9840 2335
rect 9890 2235 9950 2335
rect 10000 2235 10060 2335
rect 10110 2235 10170 2335
rect 10220 2235 10280 2335
rect 10330 2235 10390 2335
rect 10440 2235 10500 2335
rect 10550 2235 10610 2335
rect 10660 2235 10720 2335
<< ndiff >>
rect 8480 1990 8530 2005
rect 8480 1920 8495 1990
rect 8515 1920 8530 1990
rect 8480 1905 8530 1920
rect 8590 1990 8640 2005
rect 8590 1920 8605 1990
rect 8625 1920 8640 1990
rect 8590 1905 8640 1920
rect 8700 1990 8750 2005
rect 8700 1920 8715 1990
rect 8735 1920 8750 1990
rect 8700 1905 8750 1920
rect 8810 1990 8860 2005
rect 8810 1920 8825 1990
rect 8845 1920 8860 1990
rect 8810 1905 8860 1920
rect 8920 1990 8970 2005
rect 8920 1920 8935 1990
rect 8955 1920 8970 1990
rect 8920 1905 8970 1920
rect 9030 1990 9080 2005
rect 9030 1920 9045 1990
rect 9065 1920 9080 1990
rect 9030 1905 9080 1920
rect 9140 1990 9190 2005
rect 9240 1990 9290 2005
rect 9140 1920 9155 1990
rect 9175 1920 9190 1990
rect 9240 1920 9255 1990
rect 9275 1920 9290 1990
rect 9140 1905 9190 1920
rect 9240 1905 9290 1920
rect 9350 1990 9400 2005
rect 9350 1920 9365 1990
rect 9385 1920 9400 1990
rect 9350 1905 9400 1920
rect 9460 1990 9510 2005
rect 9460 1920 9475 1990
rect 9495 1920 9510 1990
rect 9460 1905 9510 1920
rect 9570 1990 9620 2005
rect 9570 1920 9585 1990
rect 9605 1920 9620 1990
rect 9570 1905 9620 1920
rect 9680 1990 9730 2005
rect 9680 1920 9695 1990
rect 9715 1920 9730 1990
rect 9680 1905 9730 1920
rect 9790 1990 9840 2005
rect 9790 1920 9805 1990
rect 9825 1920 9840 1990
rect 9790 1905 9840 1920
rect 9900 1990 9950 2005
rect 10000 1990 10050 2005
rect 9900 1920 9915 1990
rect 9935 1920 9950 1990
rect 10000 1920 10015 1990
rect 10035 1920 10050 1990
rect 9900 1905 9950 1920
rect 10000 1905 10050 1920
rect 10110 1990 10160 2005
rect 10110 1920 10125 1990
rect 10145 1920 10160 1990
rect 10110 1905 10160 1920
rect 10220 1990 10270 2005
rect 10220 1920 10235 1990
rect 10255 1920 10270 1990
rect 10220 1905 10270 1920
rect 10330 1990 10380 2005
rect 10330 1920 10345 1990
rect 10365 1920 10380 1990
rect 10330 1905 10380 1920
rect 10440 1990 10490 2005
rect 10440 1920 10455 1990
rect 10475 1920 10490 1990
rect 10440 1905 10490 1920
rect 10550 1990 10600 2005
rect 10550 1920 10565 1990
rect 10585 1920 10600 1990
rect 10550 1905 10600 1920
rect 10660 1990 10710 2005
rect 10660 1920 10675 1990
rect 10695 1920 10710 1990
rect 10660 1905 10710 1920
<< pdiff >>
rect 8420 2320 8470 2335
rect 8420 2250 8435 2320
rect 8455 2250 8470 2320
rect 8420 2235 8470 2250
rect 8530 2320 8580 2335
rect 8530 2250 8545 2320
rect 8565 2250 8580 2320
rect 8530 2235 8580 2250
rect 8640 2320 8690 2335
rect 8640 2250 8655 2320
rect 8675 2250 8690 2320
rect 8640 2235 8690 2250
rect 8750 2320 8800 2335
rect 8750 2250 8765 2320
rect 8785 2250 8800 2320
rect 8750 2235 8800 2250
rect 8860 2320 8910 2335
rect 8860 2250 8875 2320
rect 8895 2250 8910 2320
rect 8860 2235 8910 2250
rect 8970 2320 9020 2335
rect 8970 2250 8985 2320
rect 9005 2250 9020 2320
rect 8970 2235 9020 2250
rect 9080 2320 9130 2335
rect 9080 2250 9095 2320
rect 9115 2250 9130 2320
rect 9080 2235 9130 2250
rect 9190 2320 9240 2335
rect 9190 2250 9205 2320
rect 9225 2250 9240 2320
rect 9190 2235 9240 2250
rect 9300 2320 9350 2335
rect 9300 2250 9315 2320
rect 9335 2250 9350 2320
rect 9300 2235 9350 2250
rect 9410 2320 9460 2335
rect 9410 2250 9425 2320
rect 9445 2250 9460 2320
rect 9410 2235 9460 2250
rect 9520 2320 9570 2335
rect 9620 2320 9670 2335
rect 9520 2250 9535 2320
rect 9555 2250 9570 2320
rect 9620 2250 9635 2320
rect 9655 2250 9670 2320
rect 9520 2235 9570 2250
rect 9620 2235 9670 2250
rect 9730 2320 9780 2335
rect 9730 2250 9745 2320
rect 9765 2250 9780 2320
rect 9730 2235 9780 2250
rect 9840 2320 9890 2335
rect 9840 2250 9855 2320
rect 9875 2250 9890 2320
rect 9840 2235 9890 2250
rect 9950 2320 10000 2335
rect 9950 2250 9965 2320
rect 9985 2250 10000 2320
rect 9950 2235 10000 2250
rect 10060 2320 10110 2335
rect 10060 2250 10075 2320
rect 10095 2250 10110 2320
rect 10060 2235 10110 2250
rect 10170 2320 10220 2335
rect 10170 2250 10185 2320
rect 10205 2250 10220 2320
rect 10170 2235 10220 2250
rect 10280 2320 10330 2335
rect 10280 2250 10295 2320
rect 10315 2250 10330 2320
rect 10280 2235 10330 2250
rect 10390 2320 10440 2335
rect 10390 2250 10405 2320
rect 10425 2250 10440 2320
rect 10390 2235 10440 2250
rect 10500 2320 10550 2335
rect 10500 2250 10515 2320
rect 10535 2250 10550 2320
rect 10500 2235 10550 2250
rect 10610 2320 10660 2335
rect 10610 2250 10625 2320
rect 10645 2250 10660 2320
rect 10610 2235 10660 2250
rect 10720 2320 10770 2335
rect 10720 2250 10735 2320
rect 10755 2250 10770 2320
rect 10720 2235 10770 2250
<< ndiffc >>
rect 8495 1920 8515 1990
rect 8605 1920 8625 1990
rect 8715 1920 8735 1990
rect 8825 1920 8845 1990
rect 8935 1920 8955 1990
rect 9045 1920 9065 1990
rect 9155 1920 9175 1990
rect 9255 1920 9275 1990
rect 9365 1920 9385 1990
rect 9475 1920 9495 1990
rect 9585 1920 9605 1990
rect 9695 1920 9715 1990
rect 9805 1920 9825 1990
rect 9915 1920 9935 1990
rect 10015 1920 10035 1990
rect 10125 1920 10145 1990
rect 10235 1920 10255 1990
rect 10345 1920 10365 1990
rect 10455 1920 10475 1990
rect 10565 1920 10585 1990
rect 10675 1920 10695 1990
<< pdiffc >>
rect 8435 2250 8455 2320
rect 8545 2250 8565 2320
rect 8655 2250 8675 2320
rect 8765 2250 8785 2320
rect 8875 2250 8895 2320
rect 8985 2250 9005 2320
rect 9095 2250 9115 2320
rect 9205 2250 9225 2320
rect 9315 2250 9335 2320
rect 9425 2250 9445 2320
rect 9535 2250 9555 2320
rect 9635 2250 9655 2320
rect 9745 2250 9765 2320
rect 9855 2250 9875 2320
rect 9965 2250 9985 2320
rect 10075 2250 10095 2320
rect 10185 2250 10205 2320
rect 10295 2250 10315 2320
rect 10405 2250 10425 2320
rect 10515 2250 10535 2320
rect 10625 2250 10645 2320
rect 10735 2250 10755 2320
<< psubdiff >>
rect 8430 1990 8480 2005
rect 8430 1920 8445 1990
rect 8465 1920 8480 1990
rect 8430 1905 8480 1920
rect 9190 1990 9240 2005
rect 9190 1920 9205 1990
rect 9225 1920 9240 1990
rect 9190 1905 9240 1920
rect 9950 1990 10000 2005
rect 9950 1920 9965 1990
rect 9985 1920 10000 1990
rect 9950 1905 10000 1920
rect 10710 1990 10760 2005
rect 10710 1920 10725 1990
rect 10745 1920 10760 1990
rect 10710 1905 10760 1920
<< nsubdiff >>
rect 8370 2320 8420 2335
rect 8370 2250 8385 2320
rect 8405 2250 8420 2320
rect 8370 2235 8420 2250
rect 9570 2320 9620 2335
rect 9570 2250 9585 2320
rect 9605 2250 9620 2320
rect 9570 2235 9620 2250
rect 10770 2320 10820 2335
rect 10770 2250 10785 2320
rect 10805 2250 10820 2320
rect 10770 2235 10820 2250
<< psubdiffcont >>
rect 8445 1920 8465 1990
rect 9205 1920 9225 1990
rect 9965 1920 9985 1990
rect 10725 1920 10745 1990
<< nsubdiffcont >>
rect 8385 2250 8405 2320
rect 9585 2250 9605 2320
rect 10785 2250 10805 2320
<< poly >>
rect 10555 2405 10610 2415
rect 10555 2370 10565 2405
rect 10600 2370 10610 2405
rect 10555 2360 10610 2370
rect 8470 2335 8530 2350
rect 8580 2335 8640 2350
rect 8690 2335 8750 2350
rect 8800 2335 8860 2350
rect 8910 2335 8970 2350
rect 9020 2335 9080 2350
rect 9130 2335 9190 2350
rect 9240 2335 9300 2350
rect 9350 2335 9410 2350
rect 9460 2335 9520 2350
rect 9670 2335 9730 2350
rect 9780 2345 10610 2360
rect 9780 2335 9840 2345
rect 9890 2335 9950 2345
rect 10000 2335 10060 2345
rect 10110 2335 10170 2345
rect 10220 2335 10280 2345
rect 10330 2335 10390 2345
rect 10440 2335 10500 2345
rect 10550 2335 10610 2345
rect 10660 2335 10720 2350
rect 8470 2225 8530 2235
rect 8425 2210 8530 2225
rect 8425 2190 8435 2210
rect 8455 2205 8530 2210
rect 8580 2225 8640 2235
rect 8690 2225 8750 2235
rect 8800 2225 8860 2235
rect 8910 2225 8970 2235
rect 9020 2225 9080 2235
rect 9130 2225 9190 2235
rect 9240 2225 9300 2235
rect 9350 2225 9410 2235
rect 8580 2205 9410 2225
rect 9460 2225 9520 2235
rect 9670 2225 9730 2235
rect 9460 2210 9730 2225
rect 9780 2220 9840 2235
rect 9890 2220 9950 2235
rect 10000 2220 10060 2235
rect 10110 2220 10170 2235
rect 10220 2220 10280 2235
rect 10330 2220 10390 2235
rect 10440 2220 10500 2235
rect 10550 2220 10610 2235
rect 10660 2225 10720 2235
rect 10660 2210 10765 2225
rect 8455 2190 8465 2205
rect 8425 2180 8465 2190
rect 9575 2190 9585 2210
rect 9605 2190 9615 2210
rect 9575 2180 9615 2190
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 8485 2050 8525 2060
rect 8485 2030 8495 2050
rect 8515 2030 8525 2050
rect 8650 2050 8690 2060
rect 8650 2030 8660 2050
rect 8680 2030 8690 2050
rect 8760 2050 8800 2060
rect 8760 2030 8770 2050
rect 8790 2030 8800 2050
rect 8870 2050 8910 2060
rect 8870 2030 8880 2050
rect 8900 2030 8910 2050
rect 8980 2050 9020 2060
rect 8980 2030 8990 2050
rect 9010 2030 9020 2050
rect 9195 2050 9235 2060
rect 9195 2030 9205 2050
rect 9225 2030 9235 2050
rect 9955 2050 9995 2060
rect 9955 2030 9965 2050
rect 9985 2030 9995 2050
rect 10665 2050 10705 2060
rect 10665 2030 10675 2050
rect 10695 2030 10705 2050
rect 8485 2015 8590 2030
rect 8530 2005 8590 2015
rect 8640 2015 9030 2030
rect 8640 2005 8700 2015
rect 8750 2005 8810 2015
rect 8860 2005 8920 2015
rect 8970 2005 9030 2015
rect 9080 2015 9350 2030
rect 9080 2005 9140 2015
rect 9290 2005 9350 2015
rect 9400 2015 9790 2030
rect 9400 2005 9460 2015
rect 9510 2005 9570 2015
rect 9620 2005 9680 2015
rect 9730 2005 9790 2015
rect 9840 2015 10110 2030
rect 9840 2005 9900 2015
rect 10050 2005 10110 2015
rect 10160 2005 10220 2020
rect 10270 2005 10330 2020
rect 10380 2005 10440 2020
rect 10490 2005 10550 2020
rect 10600 2015 10705 2030
rect 10600 2005 10660 2015
rect 8530 1890 8590 1905
rect 8640 1890 8700 1905
rect 8750 1890 8810 1905
rect 8860 1890 8920 1905
rect 8970 1865 9030 1905
rect 9080 1890 9140 1905
rect 9290 1890 9350 1905
rect 9400 1865 9460 1905
rect 9510 1890 9570 1905
rect 9620 1890 9680 1905
rect 9730 1890 9790 1905
rect 9840 1890 9900 1905
rect 10050 1890 10110 1905
rect 10160 1895 10220 1905
rect 10270 1895 10330 1905
rect 10380 1895 10440 1905
rect 10490 1895 10550 1905
rect 10160 1880 10550 1895
rect 10600 1890 10660 1905
rect 8970 1850 9460 1865
rect 10495 1870 10550 1880
rect 10495 1835 10505 1870
rect 10540 1835 10550 1870
rect 10495 1825 10550 1835
<< polycont >>
rect 10565 2370 10600 2405
rect 8435 2190 8455 2210
rect 9585 2190 9605 2210
rect 10735 2190 10755 2210
rect 8495 2030 8515 2050
rect 8660 2030 8680 2050
rect 8770 2030 8790 2050
rect 8880 2030 8900 2050
rect 8990 2030 9010 2050
rect 9205 2030 9225 2050
rect 9965 2030 9985 2050
rect 10675 2030 10695 2050
rect 10505 1835 10540 1870
<< locali >>
rect 8205 2785 10905 2795
rect 8205 2750 10860 2785
rect 10895 2750 10905 2785
rect 8205 2740 10905 2750
rect 10555 2405 10905 2415
rect 10555 2370 10565 2405
rect 10600 2370 10860 2405
rect 10895 2370 10905 2405
rect 10555 2360 10905 2370
rect 8375 2320 8465 2330
rect 8375 2250 8385 2320
rect 8405 2250 8435 2320
rect 8455 2250 8465 2320
rect 8375 2240 8465 2250
rect 8425 2210 8465 2240
rect 8425 2190 8435 2210
rect 8455 2190 8465 2210
rect 8425 2180 8465 2190
rect 8535 2320 8575 2330
rect 8535 2250 8545 2320
rect 8565 2250 8575 2320
rect 8535 2210 8575 2250
rect 8645 2320 8685 2330
rect 8645 2250 8655 2320
rect 8675 2250 8685 2320
rect 8645 2240 8685 2250
rect 8755 2320 8795 2330
rect 8755 2250 8765 2320
rect 8785 2250 8795 2320
rect 8755 2210 8795 2250
rect 8865 2320 8905 2330
rect 8865 2250 8875 2320
rect 8895 2250 8905 2320
rect 8865 2240 8905 2250
rect 8975 2320 9015 2330
rect 8975 2250 8985 2320
rect 9005 2250 9015 2320
rect 8975 2210 9015 2250
rect 9085 2320 9125 2330
rect 9085 2250 9095 2320
rect 9115 2250 9125 2320
rect 9085 2240 9125 2250
rect 9195 2320 9235 2330
rect 9195 2250 9205 2320
rect 9225 2250 9235 2320
rect 9195 2210 9235 2250
rect 9305 2320 9345 2330
rect 9305 2250 9315 2320
rect 9335 2250 9345 2320
rect 9305 2240 9345 2250
rect 9415 2320 9455 2330
rect 9415 2250 9425 2320
rect 9445 2250 9455 2320
rect 9415 2210 9455 2250
rect 9525 2320 9665 2330
rect 9525 2250 9535 2320
rect 9555 2250 9585 2320
rect 9605 2250 9635 2320
rect 9655 2250 9665 2320
rect 9525 2240 9665 2250
rect 9735 2320 9775 2330
rect 9735 2250 9745 2320
rect 9765 2250 9775 2320
rect 8535 2170 9455 2210
rect 9575 2210 9615 2240
rect 9575 2190 9585 2210
rect 9605 2190 9615 2210
rect 9575 2180 9615 2190
rect 9735 2215 9775 2250
rect 9845 2320 9885 2330
rect 9845 2250 9855 2320
rect 9875 2250 9885 2320
rect 9845 2240 9885 2250
rect 9955 2320 9995 2330
rect 9955 2250 9965 2320
rect 9985 2250 9995 2320
rect 9955 2215 9995 2250
rect 10065 2320 10105 2330
rect 10065 2250 10075 2320
rect 10095 2250 10105 2320
rect 10065 2240 10105 2250
rect 10175 2320 10215 2330
rect 10175 2250 10185 2320
rect 10205 2250 10215 2320
rect 10175 2215 10215 2250
rect 10285 2320 10325 2330
rect 10285 2250 10295 2320
rect 10315 2250 10325 2320
rect 10285 2240 10325 2250
rect 10395 2320 10435 2330
rect 10395 2250 10405 2320
rect 10425 2250 10435 2320
rect 10395 2215 10435 2250
rect 10505 2320 10545 2330
rect 10505 2250 10515 2320
rect 10535 2250 10545 2320
rect 10505 2240 10545 2250
rect 10615 2320 10655 2330
rect 10615 2250 10625 2320
rect 10645 2250 10655 2320
rect 10615 2215 10655 2250
rect 9735 2175 10655 2215
rect 10725 2320 10815 2330
rect 10725 2250 10735 2320
rect 10755 2250 10785 2320
rect 10805 2250 10815 2320
rect 10725 2240 10815 2250
rect 10725 2210 10765 2240
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 8155 2080 8635 2100
rect 8595 2060 8635 2080
rect 9355 2060 9395 2170
rect 10555 2060 10595 2175
rect 8485 2050 8525 2060
rect 8485 2030 8495 2050
rect 8515 2030 8525 2050
rect 8485 2000 8525 2030
rect 8435 1990 8525 2000
rect 8435 1920 8445 1990
rect 8465 1920 8495 1990
rect 8515 1920 8525 1990
rect 8435 1910 8525 1920
rect 8595 2050 9075 2060
rect 8595 2030 8660 2050
rect 8680 2030 8770 2050
rect 8790 2030 8880 2050
rect 8900 2030 8990 2050
rect 9010 2030 9075 2050
rect 8595 2020 9075 2030
rect 8595 1990 8635 2020
rect 8595 1920 8605 1990
rect 8625 1920 8635 1990
rect 8595 1910 8635 1920
rect 8705 1990 8745 2000
rect 8705 1920 8715 1990
rect 8735 1920 8745 1990
rect 8705 1910 8745 1920
rect 8815 1990 8855 2020
rect 8815 1920 8825 1990
rect 8845 1920 8855 1990
rect 8815 1910 8855 1920
rect 8925 1990 8965 2000
rect 8925 1920 8935 1990
rect 8955 1920 8965 1990
rect 8925 1910 8965 1920
rect 9035 1990 9075 2020
rect 9195 2050 9235 2060
rect 9195 2030 9205 2050
rect 9225 2030 9235 2050
rect 9195 2000 9235 2030
rect 9355 2020 9835 2060
rect 9035 1920 9045 1990
rect 9065 1920 9075 1990
rect 9035 1910 9075 1920
rect 9145 1990 9285 2000
rect 9145 1920 9155 1990
rect 9175 1920 9205 1990
rect 9225 1920 9255 1990
rect 9275 1920 9285 1990
rect 9145 1910 9285 1920
rect 9355 1990 9395 2020
rect 9355 1920 9365 1990
rect 9385 1920 9395 1990
rect 9355 1910 9395 1920
rect 9465 1990 9505 2000
rect 9465 1920 9475 1990
rect 9495 1920 9505 1990
rect 9465 1910 9505 1920
rect 9575 1990 9615 2020
rect 9575 1920 9585 1990
rect 9605 1920 9615 1990
rect 9575 1910 9615 1920
rect 9685 1990 9725 2000
rect 9685 1920 9695 1990
rect 9715 1920 9725 1990
rect 9685 1910 9725 1920
rect 9795 1990 9835 2020
rect 9955 2050 9995 2060
rect 9955 2030 9965 2050
rect 9985 2030 9995 2050
rect 9955 2000 9995 2030
rect 10115 2020 10595 2060
rect 9795 1920 9805 1990
rect 9825 1920 9835 1990
rect 9795 1910 9835 1920
rect 9905 1990 10045 2000
rect 9905 1920 9915 1990
rect 9935 1920 9965 1990
rect 9985 1920 10015 1990
rect 10035 1920 10045 1990
rect 9905 1910 10045 1920
rect 10115 1990 10155 2020
rect 10115 1920 10125 1990
rect 10145 1920 10155 1990
rect 10115 1910 10155 1920
rect 10225 1990 10265 2000
rect 10225 1920 10235 1990
rect 10255 1920 10265 1990
rect 10225 1910 10265 1920
rect 10335 1990 10375 2020
rect 10335 1920 10345 1990
rect 10365 1920 10375 1990
rect 10335 1910 10375 1920
rect 10445 1990 10485 2000
rect 10445 1920 10455 1990
rect 10475 1920 10485 1990
rect 10445 1910 10485 1920
rect 10555 1990 10595 2020
rect 10555 1920 10565 1990
rect 10585 1920 10595 1990
rect 10555 1910 10595 1920
rect 10665 2050 10705 2060
rect 10665 2030 10675 2050
rect 10695 2030 10705 2050
rect 10665 2000 10705 2030
rect 10665 1990 10755 2000
rect 10665 1920 10675 1990
rect 10695 1920 10725 1990
rect 10745 1920 10755 1990
rect 10665 1910 10755 1920
rect 10495 1870 10885 1880
rect 10495 1835 10505 1870
rect 10540 1835 10840 1870
rect 10875 1835 10885 1870
rect 10495 1825 10885 1835
rect 8190 1650 10885 1660
rect 8190 1615 10840 1650
rect 10875 1615 10885 1650
rect 8190 1605 10885 1615
<< viali >>
rect 10860 2750 10895 2785
rect 10860 2370 10895 2405
rect 8385 2250 8405 2320
rect 8435 2250 8455 2320
rect 8655 2250 8675 2320
rect 8875 2250 8895 2320
rect 9095 2250 9115 2320
rect 9315 2250 9335 2320
rect 9535 2250 9555 2320
rect 9585 2250 9605 2320
rect 9635 2250 9655 2320
rect 9855 2250 9875 2320
rect 10075 2250 10095 2320
rect 10295 2250 10315 2320
rect 10515 2250 10535 2320
rect 10735 2250 10755 2320
rect 10785 2250 10805 2320
rect 8445 1920 8465 1990
rect 8495 1920 8515 1990
rect 8715 1920 8735 1990
rect 8935 1920 8955 1990
rect 9155 1920 9175 1990
rect 9205 1920 9225 1990
rect 9255 1920 9275 1990
rect 9475 1920 9495 1990
rect 9695 1920 9715 1990
rect 9915 1920 9935 1990
rect 9965 1920 9985 1990
rect 10015 1920 10035 1990
rect 10235 1920 10255 1990
rect 10455 1920 10475 1990
rect 10675 1920 10695 1990
rect 10725 1920 10745 1990
rect 10840 1835 10875 1870
rect 10840 1615 10875 1650
<< metal1 >>
rect 10850 2785 10905 2795
rect 10850 2750 10860 2785
rect 10895 2750 10905 2785
rect 10850 2740 10905 2750
rect 10850 2405 10905 2415
rect 10850 2370 10860 2405
rect 10895 2370 10905 2405
rect 10850 2360 10905 2370
rect 8370 2330 10820 2335
rect 8340 2320 10820 2330
rect 8340 2250 8385 2320
rect 8405 2250 8435 2320
rect 8455 2250 8655 2320
rect 8675 2250 8875 2320
rect 8895 2250 9095 2320
rect 9115 2250 9315 2320
rect 9335 2250 9535 2320
rect 9555 2250 9585 2320
rect 9605 2250 9635 2320
rect 9655 2250 9855 2320
rect 9875 2250 10075 2320
rect 10095 2250 10295 2320
rect 10315 2250 10515 2320
rect 10535 2250 10735 2320
rect 10755 2250 10785 2320
rect 10805 2250 10820 2320
rect 8340 2240 10820 2250
rect 8370 2235 10820 2240
rect 8340 1990 10760 2005
rect 8340 1920 8445 1990
rect 8465 1920 8495 1990
rect 8515 1920 8715 1990
rect 8735 1920 8935 1990
rect 8955 1920 9155 1990
rect 9175 1920 9205 1990
rect 9225 1920 9255 1990
rect 9275 1920 9475 1990
rect 9495 1920 9695 1990
rect 9715 1920 9915 1990
rect 9935 1920 9965 1990
rect 9985 1920 10015 1990
rect 10035 1920 10235 1990
rect 10255 1920 10455 1990
rect 10475 1920 10675 1990
rect 10695 1920 10725 1990
rect 10745 1920 10760 1990
rect 8340 1905 10760 1920
rect 10830 1870 10885 1880
rect 10830 1835 10840 1870
rect 10875 1835 10885 1870
rect 10830 1825 10885 1835
rect 10830 1650 10885 1660
rect 10830 1615 10840 1650
rect 10875 1615 10885 1650
rect 10830 1605 10885 1615
<< via1 >>
rect 10860 2750 10895 2785
rect 10860 2370 10895 2405
rect 10840 1835 10875 1870
rect 10840 1615 10875 1650
<< metal2 >>
rect 10850 2785 10905 2795
rect 10850 2750 10860 2785
rect 10895 2750 10905 2785
rect 10850 2740 10905 2750
rect 10850 2405 10905 2415
rect 10850 2370 10860 2405
rect 10895 2370 10905 2405
rect 10850 2360 10905 2370
rect 10830 1870 10885 1880
rect 10830 1835 10840 1870
rect 10875 1835 10885 1870
rect 10830 1825 10885 1835
rect 10830 1650 10885 1660
rect 10830 1615 10840 1650
rect 10875 1615 10885 1650
rect 10830 1605 10885 1615
<< via2 >>
rect 10860 2750 10895 2785
rect 10860 2370 10895 2405
rect 10840 1835 10875 1870
rect 10840 1615 10875 1650
<< metal3 >>
rect 10850 2785 11655 2795
rect 10850 2750 10860 2785
rect 10895 2750 11655 2785
rect 10850 2740 11655 2750
rect 10850 2405 10905 2415
rect 10850 2370 10860 2405
rect 10895 2370 10905 2405
rect 10850 2360 10905 2370
rect 11025 2345 11655 2740
rect 10830 1870 10885 1880
rect 10830 1835 10840 1870
rect 10875 1835 10885 1870
rect 10830 1825 10885 1835
rect 11005 1660 11295 1895
rect 10830 1650 11295 1660
rect 10830 1615 10840 1650
rect 10875 1615 11295 1650
rect 10830 1605 11295 1615
<< via3 >>
rect 10860 2370 10895 2405
rect 10840 1835 10875 1870
<< mimcap >>
rect 11040 2405 11640 2780
rect 11040 2370 11050 2405
rect 11085 2370 11640 2405
rect 11040 2360 11640 2370
rect 11020 1870 11280 1880
rect 11020 1835 11030 1870
rect 11065 1835 11280 1870
rect 11020 1620 11280 1835
<< mimcapcontact >>
rect 11050 2370 11085 2405
rect 11030 1835 11065 1870
<< metal4 >>
rect 10850 2405 11095 2415
rect 10850 2370 10860 2405
rect 10895 2370 11050 2405
rect 11085 2370 11095 2405
rect 10850 2360 11095 2370
rect 10830 1870 11075 1880
rect 10830 1835 10840 1870
rect 10875 1835 11030 1870
rect 11065 1835 11075 1870
rect 10830 1825 11075 1835
<< labels >>
flabel locali 8155 2090 8155 2090 7 FreeSans 400 0 -200 0 I_IN
flabel metal1 8340 1950 8340 1950 7 FreeSans 400 0 -200 0 GNDA
flabel metal1 8340 2285 8340 2285 7 FreeSans 400 0 -200 0 VDDA
flabel locali 9355 2110 9355 2110 7 FreeSans 400 0 -200 0 x
flabel poly 8915 2205 8915 2205 5 FreeSans 400 0 0 -200 opamp_out
flabel poly 10200 2360 10200 2360 1 FreeSans 400 0 0 200 UP_input
flabel poly 10355 1880 10355 1880 5 FreeSans 400 0 0 -200 DOWN_input
flabel locali 8190 1630 8190 1630 7 FreeSans 400 0 -200 0 DOWN
flabel locali 8205 2770 8205 2770 7 FreeSans 400 0 -200 0 UP_b
<< end >>
