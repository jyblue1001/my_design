* NGSPICE file created from charge_pump_cell.ext - technology: sky130A

**.subckt charge_pump_cell
X0 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X1 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X2 a_17540_4470# I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X3 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X4 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X5 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X6 a_18600_3120# a_18310_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 a_20050_3120# a_19470_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X8 I_IN I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X9 a_17800_2610# I_IN a_17540_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X10 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X11 a_19470_3120# w_17500_3540# a_19050_3120# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X12 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X13 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X14 a_18310_3120# a_18020_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X15 a_20050_3120# a_19470_3120# I_IN w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 I_IN I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X17 a_18890_3120# a_18600_3120# sky130_fd_pr__cap_mim_m3_1 l=6 w=4.2
X18 w_17500_3540# DOWN_PFD a_19050_3120# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X19 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X20 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X21 a_18020_3120# UP_PFD w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X22 a_17800_2610# I_IN I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X23 a_18890_3120# a_18600_3120# OPAMP_out w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X24 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X25 a_17800_2610# I_IN I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X26 a_19760_3120# a_19470_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X28 a_18310_3120# a_18020_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X29 a_20050_3120# a_19760_3120# I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X30 a_17800_2610# DOWN_PFD a_19050_3120# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X31 a_17800_2610# a_20050_3120# a_19460_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X32 a_19460_4470# a_20050_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X33 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X34 a_18020_3120# UP_PFD a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X35 a_20050_3120# a_19760_3120# sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
X36 a_19460_4470# a_20050_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X37 a_18890_3120# a_18310_3120# OPAMP_out a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 a_19760_3120# a_19470_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X40 a_17800_2610# a_20050_3120# a_19460_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X41 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X42 a_18890_3120# a_18310_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X43 a_18600_3120# a_18310_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X44 a_19470_3120# a_17800_2610# a_19050_3120# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X45 a_17540_4470# I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X46 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X47 a_17800_2610# I_IN a_17540_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
**.ends

