* PEX produced on Tue Jul 15 03:05:21 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_12.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_12 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t189 bgr_7_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_14_0.Vb3.t1 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_7_0.V_TOP.t9 VDDA.t289 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t2 GNDA.t284 GNDA.t285 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X4 GNDA.t6 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 two_stage_opamp_dummy_magic_14_0.V_source.t29 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 VOUT+.t19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VDDA.t78 two_stage_opamp_dummy_magic_14_0.X.t25 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X7 VOUT+.t20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 GNDA.t95 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 VOUT-.t3 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X9 VDDA.t83 bgr_7_0.V_TOP.t14 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X10 VDDA.t288 VDDA.t286 two_stage_opamp_dummy_magic_14_0.err_amp_out.t0 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X11 VOUT+.t21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GNDA.t283 GNDA.t281 VDDA.t361 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X13 bgr_7_0.Vin+.t5 bgr_7_0.V_TOP.t15 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 two_stage_opamp_dummy_magic_14_0.X.t26 GNDA.t305 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X15 VDDA.t135 bgr_7_0.V_mir1.t17 bgr_7_0.1st_Vout_1.t5 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X16 VOUT+.t22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 bgr_7_0.1st_Vout_2.t11 bgr_7_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 two_stage_opamp_dummy_magic_14_0.X.t22 two_stage_opamp_dummy_magic_14_0.Vb2.t11 two_stage_opamp_dummy_magic_14_0.VD3.t19 two_stage_opamp_dummy_magic_14_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X19 GNDA.t42 two_stage_opamp_dummy_magic_14_0.Y.t25 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X20 VOUT+.t23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 bgr_7_0.1st_Vout_2.t2 bgr_7_0.V_CUR_REF_REG.t3 bgr_7_0.V_p_2.t4 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X22 VOUT+.t24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 VOUT+.t25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 a_7460_23988.t0 bgr_7_0.Vin+.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=6
X25 two_stage_opamp_dummy_magic_14_0.VD2.t16 GNDA.t279 GNDA.t280 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X26 VDDA.t309 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t2 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X27 two_stage_opamp_dummy_magic_14_0.VD1.t13 two_stage_opamp_dummy_magic_14_0.Vb1.t12 two_stage_opamp_dummy_magic_14_0.X.t1 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X28 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t5 GNDA.t277 GNDA.t278 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X29 VOUT+.t26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 two_stage_opamp_dummy_magic_14_0.VD1.t12 two_stage_opamp_dummy_magic_14_0.Vb1.t13 two_stage_opamp_dummy_magic_14_0.X.t18 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X31 bgr_7_0.1st_Vout_2.t12 bgr_7_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 two_stage_opamp_dummy_magic_14_0.VD2.t5 two_stage_opamp_dummy_magic_14_0.Vb1.t14 two_stage_opamp_dummy_magic_14_0.Y.t13 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X33 GNDA.t308 a_6930_22564.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X34 VDDA.t285 VDDA.t283 VDDA.t285 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0 ps=0 w=2 l=0.15
X35 GNDA.t276 GNDA.t275 two_stage_opamp_dummy_magic_14_0.Y.t23 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X36 VDDA.t303 bgr_7_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X37 VOUT-.t20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT-.t21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT-.t22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT+.t27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 bgr_7_0.1st_Vout_1.t11 bgr_7_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 bgr_7_0.1st_Vout_2.t4 bgr_7_0.V_mir2.t17 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X43 VDDA.t76 bgr_7_0.V_TOP.t16 bgr_7_0.Vin-.t6 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X44 bgr_7_0.1st_Vout_1.t8 bgr_7_0.Vin+.t6 bgr_7_0.V_p_1.t10 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X45 GNDA.t148 VDDA.t412 bgr_7_0.V_p_2.t5 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X46 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_14_0.X.t27 VDDA.t32 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X47 VOUT+.t28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 bgr_7_0.cap_res2.t20 bgr_7_0.PFET_GATE_10uA.t6 GNDA.t124 sky130_fd_pr__res_high_po_0p35 l=2.05
X49 bgr_7_0.1st_Vout_1.t12 bgr_7_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VOUT-.t0 two_stage_opamp_dummy_magic_14_0.X.t28 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X51 two_stage_opamp_dummy_magic_14_0.V_source.t2 VIN-.t0 two_stage_opamp_dummy_magic_14_0.VD1.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X52 VOUT+.t29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VOUT-.t23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 two_stage_opamp_dummy_magic_14_0.V_source.t34 two_stage_opamp_dummy_magic_14_0.Vb1.t15 two_stage_opamp_dummy_magic_14_0.Vb1_2.t4 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X55 two_stage_opamp_dummy_magic_14_0.VD4.t37 two_stage_opamp_dummy_magic_14_0.Vb3.t8 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X56 two_stage_opamp_dummy_magic_14_0.V_source.t38 VIN+.t0 two_stage_opamp_dummy_magic_14_0.VD2.t20 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X57 VOUT-.t24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VOUT-.t25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VDDA.t36 two_stage_opamp_dummy_magic_14_0.Y.t26 VOUT+.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X60 two_stage_opamp_dummy_magic_14_0.err_amp_out.t2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t5 GNDA.t30 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X61 two_stage_opamp_dummy_magic_14_0.V_source.t28 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X62 VDDA.t394 bgr_7_0.1st_Vout_1.t13 bgr_7_0.V_TOP.t13 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X63 bgr_7_0.V_TOP.t17 VDDA.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 VOUT-.t26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 GNDA.t274 GNDA.t272 bgr_7_0.NFET_GATE_10uA.t0 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X66 bgr_7_0.START_UP.t5 bgr_7_0.V_TOP.t18 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X67 VOUT-.t27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 bgr_7_0.NFET_GATE_10uA.t6 GNDA.t187 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X69 VDDA.t355 two_stage_opamp_dummy_magic_14_0.Vb3.t9 two_stage_opamp_dummy_magic_14_0.VD3.t37 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X70 bgr_7_0.1st_Vout_1.t10 bgr_7_0.Vin+.t7 bgr_7_0.V_p_1.t9 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X71 VOUT-.t28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 GNDA.t132 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 two_stage_opamp_dummy_magic_14_0.V_source.t27 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X73 VOUT+.t30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 VDDA.t389 two_stage_opamp_dummy_magic_14_0.X.t29 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X75 bgr_7_0.1st_Vout_1.t14 bgr_7_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_14_0.Y.t27 VDDA.t94 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X77 two_stage_opamp_dummy_magic_14_0.V_err_p.t2 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X78 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t3 VIN-.t1 two_stage_opamp_dummy_magic_14_0.V_p_mir.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X79 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_14_0.Y.t28 VDDA.t84 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X80 bgr_7_0.V_TOP.t19 VDDA.t155 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 bgr_7_0.V_mir2.t11 bgr_7_0.V_mir2.t10 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 VDDA.t271 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X83 VOUT-.t29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT+.t10 a_5980_2720.t1 GNDA.t123 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X85 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 bgr_7_0.PFET_GATE_10uA.t11 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X86 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t9 VDDA.t280 VDDA.t282 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X87 VDDA.t365 bgr_7_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 VDDA.t364 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X88 GNDA.t62 two_stage_opamp_dummy_magic_14_0.Y.t29 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X89 VOUT+.t31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 bgr_7_0.V_TOP.t20 VDDA.t156 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 GNDA.t134 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 two_stage_opamp_dummy_magic_14_0.V_source.t26 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X92 bgr_7_0.1st_Vout_2.t1 bgr_7_0.V_CUR_REF_REG.t4 bgr_7_0.V_p_2.t3 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X93 two_stage_opamp_dummy_magic_14_0.VD4.t19 two_stage_opamp_dummy_magic_14_0.Vb2.t12 two_stage_opamp_dummy_magic_14_0.Y.t2 two_stage_opamp_dummy_magic_14_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X94 VOUT+.t2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X95 VOUT-.t30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT-.t31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT-.t32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 two_stage_opamp_dummy_magic_14_0.VD2.t8 two_stage_opamp_dummy_magic_14_0.Vb1.t16 two_stage_opamp_dummy_magic_14_0.Y.t14 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X99 two_stage_opamp_dummy_magic_14_0.V_source.t25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X100 VOUT-.t18 a_14010_2720.t1 GNDA.t307 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X101 bgr_7_0.PFET_GATE_10uA.t5 bgr_7_0.1st_Vout_2.t13 VDDA.t293 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X102 VOUT-.t33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 bgr_7_0.V_TOP.t21 VDDA.t150 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 bgr_7_0.START_UP_NFET1.t0 bgr_7_0.START_UP_NFET1 GNDA.t295 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X105 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_14_0.Vb3.t6 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X106 two_stage_opamp_dummy_magic_14_0.VD3.t17 two_stage_opamp_dummy_magic_14_0.Vb2.t13 two_stage_opamp_dummy_magic_14_0.X.t5 two_stage_opamp_dummy_magic_14_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X107 VOUT+.t32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 two_stage_opamp_dummy_magic_14_0.V_source.t6 VIN-.t2 two_stage_opamp_dummy_magic_14_0.VD1.t3 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X109 bgr_7_0.V_CUR_REF_REG.t1 VDDA.t277 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X110 VOUT-.t9 VDDA.t274 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X111 two_stage_opamp_dummy_magic_14_0.V_source.t8 VIN-.t3 two_stage_opamp_dummy_magic_14_0.VD1.t14 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X112 VOUT+.t33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 bgr_7_0.V_TOP.t22 VDDA.t151 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 GNDA.t185 bgr_7_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X115 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 bgr_7_0.NFET_GATE_10uA.t8 GNDA.t183 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_14_0.VD4.t17 two_stage_opamp_dummy_magic_14_0.Vb2.t14 two_stage_opamp_dummy_magic_14_0.Y.t1 two_stage_opamp_dummy_magic_14_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 two_stage_opamp_dummy_magic_14_0.V_source.t3 VIN+.t1 two_stage_opamp_dummy_magic_14_0.VD2.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X118 VDDA.t123 two_stage_opamp_dummy_magic_14_0.Y.t30 VOUT+.t6 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X119 GNDA.t271 GNDA.t269 two_stage_opamp_dummy_magic_14_0.VD2.t15 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X120 VOUT-.t34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 two_stage_opamp_dummy_magic_14_0.V_source.t24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X122 VOUT-.t35 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT-.t36 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT-.t37 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 bgr_7_0.1st_Vout_2.t14 bgr_7_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT+.t34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT+.t35 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 two_stage_opamp_dummy_magic_14_0.Vb1.t4 two_stage_opamp_dummy_magic_14_0.Vb1.t3 two_stage_opamp_dummy_magic_14_0.Vb1_2.t3 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X129 VOUT+.t36 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT+.t37 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VOUT+.t38 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 GNDA.t129 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_14_0.V_source.t23 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X133 a_12530_23988.t1 bgr_7_0.Vin-.t7 GNDA.t312 sky130_fd_pr__res_xhigh_po_0p35 l=6
X134 two_stage_opamp_dummy_magic_14_0.VD3.t15 two_stage_opamp_dummy_magic_14_0.Vb2.t15 two_stage_opamp_dummy_magic_14_0.X.t0 two_stage_opamp_dummy_magic_14_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X135 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_14_0.Y.t31 VDDA.t106 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X136 VOUT-.t38 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT-.t39 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 bgr_7_0.1st_Vout_2.t0 bgr_7_0.V_mir2.t18 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X139 two_stage_opamp_dummy_magic_14_0.V_err_p.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t4 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X140 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 two_stage_opamp_dummy_magic_14_0.X.t30 GNDA.t141 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X141 VOUT-.t40 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 GNDA.t303 two_stage_opamp_dummy_magic_14_0.Y.t32 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X143 VOUT-.t41 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 bgr_7_0.1st_Vout_2.t15 bgr_7_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t270 VDDA.t268 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0 ps=0 w=2 l=0.15
X146 VOUT-.t42 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT+.t39 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT-.t43 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t40 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VOUT+.t41 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 bgr_7_0.1st_Vout_1.t15 bgr_7_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VOUT+.t42 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 bgr_7_0.V_mir1.t3 bgr_7_0.Vin-.t8 bgr_7_0.V_p_1.t4 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X154 bgr_7_0.V_mir1.t16 bgr_7_0.V_mir1.t15 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X155 two_stage_opamp_dummy_magic_14_0.VD2.t4 two_stage_opamp_dummy_magic_14_0.Vb1.t17 two_stage_opamp_dummy_magic_14_0.Y.t12 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X156 GNDA.t1 a_7580_22380.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=6
X157 VOUT-.t44 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT-.t45 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VOUT+.t43 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VOUT-.t46 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT-.t47 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT-.t48 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VDDA.t353 two_stage_opamp_dummy_magic_14_0.Vb3.t10 two_stage_opamp_dummy_magic_14_0.VD4.t36 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X164 bgr_7_0.V_TOP.t23 VDDA.t152 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VDDA.t267 VDDA.t265 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X166 VOUT-.t49 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT-.t50 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 GNDA.t103 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 VOUT+.t8 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X169 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 bgr_7_0.PFET_GATE_10uA.t13 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X170 VOUT-.t5 two_stage_opamp_dummy_magic_14_0.X.t31 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X171 VOUT+.t44 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VOUT+.t45 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 two_stage_opamp_dummy_magic_14_0.V_source.t40 VIN+.t2 two_stage_opamp_dummy_magic_14_0.VD2.t21 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X174 bgr_7_0.V_mir1.t1 bgr_7_0.Vin-.t9 bgr_7_0.V_p_1.t3 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X175 two_stage_opamp_dummy_magic_14_0.X.t24 two_stage_opamp_dummy_magic_14_0.Vb1.t18 two_stage_opamp_dummy_magic_14_0.VD1.t11 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X176 VOUT+.t46 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 two_stage_opamp_dummy_magic_14_0.VD3.t36 two_stage_opamp_dummy_magic_14_0.Vb3.t11 VDDA.t351 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X178 VOUT+.t47 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 two_stage_opamp_dummy_magic_14_0.VD3.t13 two_stage_opamp_dummy_magic_14_0.Vb2.t16 two_stage_opamp_dummy_magic_14_0.X.t21 two_stage_opamp_dummy_magic_14_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X180 two_stage_opamp_dummy_magic_14_0.Vb1.t11 GNDA.t267 GNDA.t268 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X181 bgr_7_0.START_UP.t4 bgr_7_0.V_TOP.t24 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X182 VOUT-.t51 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 bgr_7_0.PFET_GATE_10uA.t4 bgr_7_0.1st_Vout_2.t16 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X184 VDDA.t38 bgr_7_0.V_mir1.t18 bgr_7_0.1st_Vout_1.t4 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X185 VOUT+.t48 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VOUT+.t49 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VOUT-.t52 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VDDA.t63 two_stage_opamp_dummy_magic_14_0.X.t32 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X189 VOUT-.t53 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 two_stage_opamp_dummy_magic_14_0.Vb2.t7 bgr_7_0.NFET_GATE_10uA.t9 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X191 VDDA.t349 two_stage_opamp_dummy_magic_14_0.Vb3.t12 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t10 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X192 GNDA.t179 bgr_7_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_14_0.Vb2.t6 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_14_0.Y.t33 VDDA.t401 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X194 VOUT+.t50 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 bgr_7_0.V_TOP.t25 VDDA.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 GNDA.t177 bgr_7_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_14_0.Vb2.t5 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X197 two_stage_opamp_dummy_magic_14_0.Y.t5 two_stage_opamp_dummy_magic_14_0.Vb2.t17 two_stage_opamp_dummy_magic_14_0.VD4.t15 two_stage_opamp_dummy_magic_14_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X198 VDDA.t264 VDDA.t262 VOUT-.t8 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X199 VOUT+.t51 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 VOUT-.t54 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 GNDA.t137 VDDA.t259 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X202 GNDA.t86 two_stage_opamp_dummy_magic_14_0.Y.t34 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X203 VOUT+.t52 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT+.t53 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VOUT+.t54 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT+.t55 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VDDA.t72 bgr_7_0.V_TOP.t26 bgr_7_0.Vin+.t4 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X208 bgr_7_0.1st_Vout_2.t5 bgr_7_0.V_mir2.t19 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X209 VOUT-.t55 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 a_14010_2720.t0 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X211 bgr_7_0.V_TOP.t12 bgr_7_0.1st_Vout_1.t16 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X212 VOUT-.t56 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT-.t57 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT-.t58 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VOUT+.t56 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 bgr_7_0.PFET_GATE_10uA.t14 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X217 VOUT-.t59 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 two_stage_opamp_dummy_magic_14_0.X.t7 two_stage_opamp_dummy_magic_14_0.Vb2.t18 two_stage_opamp_dummy_magic_14_0.VD3.t11 two_stage_opamp_dummy_magic_14_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X219 a_14330_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 GNDA.t300 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X220 VOUT+.t57 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VOUT+.t58 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 bgr_7_0.1st_Vout_2.t17 bgr_7_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 a_6810_23838.t0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X224 two_stage_opamp_dummy_magic_14_0.Y.t6 two_stage_opamp_dummy_magic_14_0.Vb2.t19 two_stage_opamp_dummy_magic_14_0.VD4.t13 two_stage_opamp_dummy_magic_14_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X225 bgr_7_0.Vin+.t1 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t100 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X226 VOUT+.t59 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t60 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT-.t60 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT-.t61 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_7_0.1st_Vout_2.t18 bgr_7_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 bgr_7_0.Vin+.t3 bgr_7_0.V_TOP.t27 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X232 VOUT-.t13 two_stage_opamp_dummy_magic_14_0.X.t33 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X233 VOUT-.t62 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VDDA.t258 VDDA.t256 bgr_7_0.PFET_GATE_10uA.t8 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X235 VOUT+.t61 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VDDA.t51 bgr_7_0.V_TOP.t28 bgr_7_0.Vin+.t2 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X237 two_stage_opamp_dummy_magic_14_0.V_source.t35 VIN+.t3 two_stage_opamp_dummy_magic_14_0.VD2.t18 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X238 VOUT+.t62 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 two_stage_opamp_dummy_magic_14_0.X.t19 two_stage_opamp_dummy_magic_14_0.Vb1.t19 two_stage_opamp_dummy_magic_14_0.VD1.t10 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X240 bgr_7_0.1st_Vout_1.t17 bgr_7_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 GNDA.t291 a_12410_22380.t1 GNDA.t290 sky130_fd_pr__res_xhigh_po_0p35 l=6
X242 GNDA.t175 bgr_7_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_14_0.Vb3.t5 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X243 VOUT-.t63 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT-.t64 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_14_0.Y.t16 GNDA.t99 sky130_fd_pr__res_high_po_1p41 l=1.41
X246 VOUT+.t63 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 bgr_7_0.cap_res1.t0 bgr_7_0.V_TOP.t0 GNDA.t50 sky130_fd_pr__res_high_po_0p35 l=2.05
X248 two_stage_opamp_dummy_magic_14_0.Vb3.t3 bgr_7_0.NFET_GATE_10uA.t13 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X249 bgr_7_0.V_mir2.t9 bgr_7_0.V_mir2.t8 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X250 VDDA.t255 VDDA.t253 bgr_7_0.V_TOP.t8 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X251 two_stage_opamp_dummy_magic_14_0.X.t6 two_stage_opamp_dummy_magic_14_0.Vb2.t20 two_stage_opamp_dummy_magic_14_0.VD3.t9 two_stage_opamp_dummy_magic_14_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 VOUT+.t64 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VOUT+.t65 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VDDA.t360 GNDA.t264 GNDA.t266 GNDA.t265 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X255 bgr_7_0.1st_Vout_1.t18 bgr_7_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VOUT-.t65 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_14_0.Y.t35 VDDA.t377 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X258 VOUT+.t66 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 bgr_7_0.V_TOP.t29 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X260 bgr_7_0.1st_Vout_2.t19 bgr_7_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_14_0.VD1.t20 VIN-.t4 two_stage_opamp_dummy_magic_14_0.V_source.t37 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X262 VOUT-.t66 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 GNDA.t299 a_13060_22630.t1 GNDA.t298 sky130_fd_pr__res_xhigh_po_0p35 l=4
X264 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 two_stage_opamp_dummy_magic_14_0.X.t34 GNDA.t310 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X265 VDDA.t397 two_stage_opamp_dummy_magic_14_0.X.t35 VOUT-.t17 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X266 VOUT+.t67 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 bgr_7_0.1st_Vout_1.t3 bgr_7_0.V_mir1.t19 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 VOUT+.t0 two_stage_opamp_dummy_magic_14_0.Y.t36 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X269 a_5420_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t0 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X270 bgr_7_0.1st_Vout_1.t19 bgr_7_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 two_stage_opamp_dummy_magic_14_0.X.t4 two_stage_opamp_dummy_magic_14_0.Vb2.t21 two_stage_opamp_dummy_magic_14_0.VD3.t7 two_stage_opamp_dummy_magic_14_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X272 VOUT-.t67 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 two_stage_opamp_dummy_magic_14_0.VD4.t27 VDDA.t235 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X274 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 VDDA.t241 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X275 VDDA.t246 VDDA.t244 bgr_7_0.NFET_GATE_10uA.t1 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X276 two_stage_opamp_dummy_magic_14_0.Vb1_2.t2 two_stage_opamp_dummy_magic_14_0.Vb1.t1 two_stage_opamp_dummy_magic_14_0.Vb1.t2 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X277 VDDA.t379 bgr_7_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X278 two_stage_opamp_dummy_magic_14_0.Y.t7 two_stage_opamp_dummy_magic_14_0.Vb2.t22 two_stage_opamp_dummy_magic_14_0.VD4.t11 two_stage_opamp_dummy_magic_14_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X279 two_stage_opamp_dummy_magic_14_0.VD2.t10 two_stage_opamp_dummy_magic_14_0.Vb1.t20 two_stage_opamp_dummy_magic_14_0.Y.t17 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X280 VOUT+.t68 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 two_stage_opamp_dummy_magic_14_0.V_p_mir.t5 GNDA.t262 GNDA.t263 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X282 VOUT+.t69 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 bgr_7_0.1st_Vout_1.t20 bgr_7_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 GNDA.t26 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 VOUT-.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X285 bgr_7_0.V_p_2.t7 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 bgr_7_0.V_mir2.t16 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X286 two_stage_opamp_dummy_magic_14_0.V_source.t11 two_stage_opamp_dummy_magic_14_0.err_amp_out.t4 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X287 VDDA.t347 two_stage_opamp_dummy_magic_14_0.Vb3.t13 two_stage_opamp_dummy_magic_14_0.VD3.t35 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X288 VDDA.t305 bgr_7_0.V_TOP.t30 bgr_7_0.START_UP.t3 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X289 VOUT+.t70 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 VOUT-.t68 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT-.t69 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VOUT+.t71 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 VOUT+.t72 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 bgr_7_0.V_TOP.t31 VDDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 bgr_7_0.V_TOP.t3 bgr_7_0.1st_Vout_1.t21 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X296 GNDA.t296 two_stage_opamp_dummy_magic_14_0.X.t36 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X297 VOUT+.t73 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VDDA.t249 VDDA.t247 GNDA.t11 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X299 VDDA.t252 VDDA.t250 two_stage_opamp_dummy_magic_14_0.VD3.t21 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X300 two_stage_opamp_dummy_magic_14_0.X.t14 two_stage_opamp_dummy_magic_14_0.Vb2.t23 two_stage_opamp_dummy_magic_14_0.VD3.t5 two_stage_opamp_dummy_magic_14_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X301 VDDA.t240 VDDA.t238 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X302 GNDA.t261 GNDA.t259 VOUT-.t11 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X303 VOUT-.t70 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 two_stage_opamp_dummy_magic_14_0.X.t9 two_stage_opamp_dummy_magic_14_0.Vb1.t21 two_stage_opamp_dummy_magic_14_0.VD1.t9 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X305 VOUT-.t71 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 bgr_7_0.V_TOP.t5 bgr_7_0.1st_Vout_1.t22 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 two_stage_opamp_dummy_magic_14_0.Y.t19 two_stage_opamp_dummy_magic_14_0.Vb1.t22 two_stage_opamp_dummy_magic_14_0.VD2.t13 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X308 VOUT+.t74 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT+.t75 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VOUT+.t76 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 bgr_7_0.NFET_GATE_10uA.t4 bgr_7_0.NFET_GATE_10uA.t3 GNDA.t171 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X312 GNDA.t169 bgr_7_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_14_0.Vb3.t2 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X313 VOUT+.t77 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 bgr_7_0.V_TOP.t32 VDDA.t307 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VDDA.t234 VDDA.t232 VDDA.t234 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X316 two_stage_opamp_dummy_magic_14_0.VD4.t9 two_stage_opamp_dummy_magic_14_0.Vb2.t24 two_stage_opamp_dummy_magic_14_0.Y.t0 two_stage_opamp_dummy_magic_14_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X317 VDDA.t126 two_stage_opamp_dummy_magic_14_0.X.t37 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X318 bgr_7_0.1st_Vout_2.t20 bgr_7_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT-.t72 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT-.t73 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT-.t74 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT+.t78 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 two_stage_opamp_dummy_magic_14_0.VD1.t15 VIN-.t5 two_stage_opamp_dummy_magic_14_0.V_source.t9 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X324 GNDA.t258 GNDA.t257 two_stage_opamp_dummy_magic_14_0.Vb1.t10 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X325 VDDA.t2 bgr_7_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 two_stage_opamp_dummy_magic_14_0.X.t38 GNDA.t309 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X327 VOUT-.t75 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VDDA.t388 two_stage_opamp_dummy_magic_14_0.X.t39 VOUT-.t16 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X329 bgr_7_0.1st_Vout_1.t23 bgr_7_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 bgr_7_0.V_mir1.t14 bgr_7_0.V_mir1.t13 VDDA.t363 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X331 VOUT+.t3 two_stage_opamp_dummy_magic_14_0.Y.t37 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X332 GNDA.t130 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_14_0.V_source.t22 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X333 VDDA.t11 bgr_7_0.V_TOP.t33 bgr_7_0.START_UP.t2 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X334 two_stage_opamp_dummy_magic_14_0.V_p_mir.t3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X335 VOUT-.t76 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 bgr_7_0.1st_Vout_2.t21 bgr_7_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 VOUT+.t79 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VOUT+.t80 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 a_7460_23988.t1 a_7580_22380.t1 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=6
X340 bgr_7_0.V_p_2.t2 bgr_7_0.V_CUR_REF_REG.t5 bgr_7_0.1st_Vout_2.t6 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X341 VOUT-.t77 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT+.t81 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 two_stage_opamp_dummy_magic_14_0.VD3.t3 two_stage_opamp_dummy_magic_14_0.Vb2.t25 two_stage_opamp_dummy_magic_14_0.X.t23 two_stage_opamp_dummy_magic_14_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X344 a_14450_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 GNDA.t122 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X345 two_stage_opamp_dummy_magic_14_0.V_source.t21 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X346 GNDA.t256 GNDA.t254 VDDA.t359 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X347 bgr_7_0.1st_Vout_2.t22 bgr_7_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 two_stage_opamp_dummy_magic_14_0.VD4.t7 two_stage_opamp_dummy_magic_14_0.Vb2.t26 two_stage_opamp_dummy_magic_14_0.Y.t8 two_stage_opamp_dummy_magic_14_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X349 bgr_7_0.1st_Vout_1.t9 bgr_7_0.Vin+.t8 bgr_7_0.V_p_1.t8 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X350 VDDA.t163 bgr_7_0.V_mir2.t20 bgr_7_0.1st_Vout_2.t7 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X351 two_stage_opamp_dummy_magic_14_0.VD4.t35 two_stage_opamp_dummy_magic_14_0.Vb3.t14 VDDA.t345 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X352 VOUT-.t78 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 VOUT-.t79 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 GNDA.t118 two_stage_opamp_dummy_magic_14_0.X.t40 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X355 bgr_7_0.1st_Vout_1.t24 bgr_7_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 GNDA.t191 GNDA.t253 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X357 bgr_7_0.NFET_GATE_10uA.t2 bgr_7_0.PFET_GATE_10uA.t17 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X358 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_14_0.Y.t38 GNDA.t101 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X359 VOUT-.t80 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 bgr_7_0.1st_Vout_2.t23 bgr_7_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 GNDA.t167 bgr_7_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_14_0.Vb2.t4 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X362 two_stage_opamp_dummy_magic_14_0.Vb2.t3 bgr_7_0.NFET_GATE_10uA.t16 GNDA.t165 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X363 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_14_0.Y.t39 GNDA.t128 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X364 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 GNDA.t250 GNDA.t252 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X365 VOUT+.t82 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 GNDA.t191 GNDA.t190 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X367 GNDA.t249 GNDA.t247 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X368 GNDA.t246 GNDA.t244 two_stage_opamp_dummy_magic_14_0.Vb2.t9 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X369 two_stage_opamp_dummy_magic_14_0.V_source.t10 VIN+.t4 two_stage_opamp_dummy_magic_14_0.VD2.t7 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X370 VOUT-.t81 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X372 VOUT+.t83 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 bgr_7_0.PFET_GATE_10uA.t7 VDDA.t229 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X374 two_stage_opamp_dummy_magic_14_0.X.t10 two_stage_opamp_dummy_magic_14_0.Vb1.t23 two_stage_opamp_dummy_magic_14_0.VD1.t8 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X375 VOUT+.t84 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 bgr_7_0.1st_Vout_1.t2 bgr_7_0.V_mir1.t20 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X377 two_stage_opamp_dummy_magic_14_0.X.t13 two_stage_opamp_dummy_magic_14_0.Vb1.t24 two_stage_opamp_dummy_magic_14_0.VD1.t7 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X378 two_stage_opamp_dummy_magic_14_0.Vb2_2.t2 two_stage_opamp_dummy_magic_14_0.Vb2.t27 VDDA.t146 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X379 VOUT-.t82 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VOUT-.t10 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X381 two_stage_opamp_dummy_magic_14_0.Y.t18 two_stage_opamp_dummy_magic_14_0.Vb1.t25 two_stage_opamp_dummy_magic_14_0.VD2.t11 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X382 bgr_7_0.V_p_2.t1 bgr_7_0.V_CUR_REF_REG.t6 bgr_7_0.1st_Vout_2.t10 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X383 VOUT-.t83 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VOUT+.t85 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 GNDA.t191 GNDA.t240 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X386 VOUT-.t84 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t127 two_stage_opamp_dummy_magic_14_0.X.t41 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X388 VOUT+.t86 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 GNDA.t191 GNDA.t239 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X390 VOUT-.t85 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 two_stage_opamp_dummy_magic_14_0.VD1.t21 VIN-.t6 two_stage_opamp_dummy_magic_14_0.V_source.t39 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X392 a_5540_5524.t1 two_stage_opamp_dummy_magic_14_0.V_tot.t3 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X393 VDDA.t44 bgr_7_0.V_mir2.t6 bgr_7_0.V_mir2.t7 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X394 two_stage_opamp_dummy_magic_14_0.VD2.t2 VIN+.t5 two_stage_opamp_dummy_magic_14_0.V_source.t4 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X395 VDDA.t343 two_stage_opamp_dummy_magic_14_0.Vb3.t15 two_stage_opamp_dummy_magic_14_0.VD4.t34 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X396 VOUT+.t9 two_stage_opamp_dummy_magic_14_0.Y.t40 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X397 VOUT+.t87 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 VOUT+.t88 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VOUT+.t89 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 GNDA.t53 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_14_0.V_source.t20 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X401 GNDA.t238 GNDA.t237 two_stage_opamp_dummy_magic_14_0.err_amp_out.t1 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X402 VOUT+.t90 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 VDDA.t42 bgr_7_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_14_0.Vb1.t0 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X404 bgr_7_0.V_p_2.t0 bgr_7_0.V_CUR_REF_REG.t7 bgr_7_0.1st_Vout_2.t9 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X405 two_stage_opamp_dummy_magic_14_0.VD4.t25 two_stage_opamp_dummy_magic_14_0.VD4.t23 two_stage_opamp_dummy_magic_14_0.Y.t10 two_stage_opamp_dummy_magic_14_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X406 VOUT+.t91 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 a_13180_23838.t0 bgr_7_0.V_CUR_REF_REG.t0 GNDA.t89 sky130_fd_pr__res_xhigh_po_0p35 l=4
X408 two_stage_opamp_dummy_magic_14_0.VD3.t34 two_stage_opamp_dummy_magic_14_0.Vb3.t16 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X409 VOUT-.t86 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 bgr_7_0.V_TOP.t34 VDDA.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VOUT-.t87 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 VOUT-.t88 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT-.t89 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT-.t90 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 two_stage_opamp_dummy_magic_14_0.V_source.t19 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X416 VOUT-.t91 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT+.t92 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 bgr_7_0.V_TOP.t35 VDDA.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_14_0.X.t42 VDDA.t112 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X420 VDDA.t34 bgr_7_0.1st_Vout_2.t24 bgr_7_0.PFET_GATE_10uA.t3 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X421 two_stage_opamp_dummy_magic_14_0.err_amp_out.t3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_14_0.V_err_p.t3 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X422 GNDA.t236 GNDA.t235 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t4 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X423 VOUT+.t93 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VDDA.t170 two_stage_opamp_dummy_magic_14_0.Y.t41 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X425 VOUT-.t92 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT+.t94 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_14_0.Y.t42 GNDA.t120 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X428 VOUT+.t95 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VOUT+.t96 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 bgr_7_0.PFET_GATE_10uA.t19 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X431 two_stage_opamp_dummy_magic_14_0.VD3.t27 two_stage_opamp_dummy_magic_14_0.VD3.t25 two_stage_opamp_dummy_magic_14_0.X.t11 two_stage_opamp_dummy_magic_14_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X432 VOUT-.t93 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VOUT-.t94 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t27 bgr_7_0.PFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X435 VOUT-.t95 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VOUT-.t96 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X438 two_stage_opamp_dummy_magic_14_0.X.t17 GNDA.t233 GNDA.t234 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X439 two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 two_stage_opamp_dummy_magic_14_0.X.t15 GNDA.t146 sky130_fd_pr__res_high_po_1p41 l=1.41
X440 VOUT-.t97 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 bgr_7_0.V_TOP.t36 VDDA.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VOUT-.t98 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 two_stage_opamp_dummy_magic_14_0.Y.t24 two_stage_opamp_dummy_magic_14_0.Vb1.t26 two_stage_opamp_dummy_magic_14_0.VD2.t17 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X444 bgr_7_0.Vin-.t5 bgr_7_0.V_TOP.t37 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X445 two_stage_opamp_dummy_magic_14_0.Y.t3 two_stage_opamp_dummy_magic_14_0.Vb2.t28 two_stage_opamp_dummy_magic_14_0.VD4.t5 two_stage_opamp_dummy_magic_14_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X446 VOUT-.t99 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 VDDA.t228 VDDA.t225 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X448 VOUT+.t97 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VOUT+.t98 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 VDDA.t339 two_stage_opamp_dummy_magic_14_0.Vb3.t17 two_stage_opamp_dummy_magic_14_0.VD4.t33 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X451 VOUT+.t99 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 GNDA.t163 bgr_7_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X453 bgr_7_0.1st_Vout_1.t1 bgr_7_0.V_mir1.t21 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X454 two_stage_opamp_dummy_magic_14_0.Vb2.t8 GNDA.t230 GNDA.t232 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X455 VOUT+.t100 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 VOUT+.t101 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 VOUT+.t102 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 bgr_7_0.1st_Vout_1.t25 bgr_7_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 GNDA.t143 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 VOUT+.t14 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X460 VOUT-.t100 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 bgr_7_0.1st_Vout_2.t25 bgr_7_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_14_0.VD1.t1 VIN-.t7 two_stage_opamp_dummy_magic_14_0.V_source.t1 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X463 VDDA.t367 two_stage_opamp_dummy_magic_14_0.X.t43 VOUT-.t12 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X464 VOUT+.t103 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 two_stage_opamp_dummy_magic_14_0.VD1.t16 VIN-.t8 two_stage_opamp_dummy_magic_14_0.V_source.t30 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X466 two_stage_opamp_dummy_magic_14_0.VD2.t3 VIN+.t6 two_stage_opamp_dummy_magic_14_0.V_source.t5 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X467 VOUT-.t101 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VOUT+.t18 two_stage_opamp_dummy_magic_14_0.Y.t43 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X469 GNDA.t117 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t4 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X470 bgr_7_0.1st_Vout_1.t26 bgr_7_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 GNDA.t114 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_14_0.V_source.t18 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X472 VOUT-.t102 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT-.t103 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT-.t104 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 a_14450_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t2 GNDA.t75 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X476 VOUT-.t105 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 bgr_7_0.V_TOP.t38 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X478 VOUT+.t104 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 GNDA.t229 GNDA.t227 VOUT+.t16 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X480 VDDA.t5 bgr_7_0.V_mir2.t4 bgr_7_0.V_mir2.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X481 VOUT+.t105 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VDDA.t125 bgr_7_0.V_mir1.t11 bgr_7_0.V_mir1.t12 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X483 VDDA.t209 VDDA.t206 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X484 two_stage_opamp_dummy_magic_14_0.V_source.t17 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X485 bgr_7_0.V_p_1.t2 bgr_7_0.Vin-.t10 bgr_7_0.V_mir1.t4 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X486 VDDA.t337 two_stage_opamp_dummy_magic_14_0.Vb3.t18 two_stage_opamp_dummy_magic_14_0.VD4.t32 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X487 two_stage_opamp_dummy_magic_14_0.Vb2.t10 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.t8 two_stage_opamp_dummy_magic_14_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X488 VOUT+.t106 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 bgr_7_0.1st_Vout_1.t27 bgr_7_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_14_0.X.t44 VDDA.t117 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X491 bgr_7_0.1st_Vout_2.t26 bgr_7_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VDDA.t391 two_stage_opamp_dummy_magic_14_0.Y.t44 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X493 VDDA.t158 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 two_stage_opamp_dummy_magic_14_0.V_err_p.t1 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X494 two_stage_opamp_dummy_magic_14_0.V_p_mir.t1 VIN+.t7 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t7 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X495 GNDA.t107 two_stage_opamp_dummy_magic_14_0.X.t45 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X496 VOUT+.t107 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VOUT+.t108 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 bgr_7_0.V_TOP.t7 VDDA.t222 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X499 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 two_stage_opamp_dummy_magic_14_0.Y.t45 GNDA.t311 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X500 VOUT+.t109 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 bgr_7_0.1st_Vout_1.t28 bgr_7_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 two_stage_opamp_dummy_magic_14_0.V_source.t16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X503 VOUT-.t106 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VDDA.t221 VDDA.t219 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X505 VDDA.t218 VDDA.t216 two_stage_opamp_dummy_magic_14_0.Vb2_2.t9 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X506 bgr_7_0.V_p_1.t1 bgr_7_0.Vin-.t11 bgr_7_0.V_mir1.t2 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X507 VOUT+.t110 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT-.t107 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT+.t111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT+.t112 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT+.t113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 bgr_7_0.1st_Vout_1.t29 bgr_7_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 two_stage_opamp_dummy_magic_14_0.Vb3.t0 GNDA.t224 GNDA.t226 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X514 VOUT+.t114 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 bgr_7_0.Vin-.t1 bgr_7_0.START_UP.t6 bgr_7_0.V_TOP.t4 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X516 two_stage_opamp_dummy_magic_14_0.Y.t11 two_stage_opamp_dummy_magic_14_0.Vb1.t27 two_stage_opamp_dummy_magic_14_0.VD2.t1 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X517 bgr_7_0.V_TOP.t2 bgr_7_0.START_UP.t7 bgr_7_0.Vin-.t0 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X518 VOUT-.t108 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT+.t115 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT+.t116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VDDA.t81 bgr_7_0.1st_Vout_2.t27 bgr_7_0.PFET_GATE_10uA.t2 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X522 bgr_7_0.V_mir1.t10 bgr_7_0.V_mir1.t9 VDDA.t297 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X523 VOUT-.t109 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 a_5540_5524.t0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X525 VOUT-.t110 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 VOUT-.t111 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 GNDA.t191 GNDA.t216 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X528 bgr_7_0.START_UP.t1 bgr_7_0.START_UP.t0 bgr_7_0.START_UP_NFET1.t0 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X529 two_stage_opamp_dummy_magic_14_0.VD4.t31 two_stage_opamp_dummy_magic_14_0.Vb3.t19 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X530 bgr_7_0.V_p_2.t10 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 bgr_7_0.V_mir2.t15 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X531 two_stage_opamp_dummy_magic_14_0.VD1.t19 GNDA.t217 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X532 VOUT+.t13 VDDA.t213 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X533 VOUT+.t7 two_stage_opamp_dummy_magic_14_0.Y.t46 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X534 two_stage_opamp_dummy_magic_14_0.VD2.t6 VIN+.t8 two_stage_opamp_dummy_magic_14_0.V_source.t7 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X535 GNDA.t223 GNDA.t220 GNDA.t222 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X536 GNDA.t215 GNDA.t214 two_stage_opamp_dummy_magic_14_0.X.t16 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X537 VOUT+.t117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VOUT+.t118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VDDA.t333 two_stage_opamp_dummy_magic_14_0.Vb3.t20 two_stage_opamp_dummy_magic_14_0.VD3.t33 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X540 VOUT-.t112 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 bgr_7_0.1st_Vout_2.t28 bgr_7_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT-.t113 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VOUT+.t119 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 two_stage_opamp_dummy_magic_14_0.Vb1_2.t1 two_stage_opamp_dummy_magic_14_0.Vb1.t7 two_stage_opamp_dummy_magic_14_0.Vb1.t8 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X545 VDDA.t93 bgr_7_0.V_mir2.t21 bgr_7_0.1st_Vout_2.t3 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X546 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 bgr_7_0.PFET_GATE_10uA.t21 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X547 VOUT-.t114 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 bgr_7_0.V_p_1.t0 bgr_7_0.Vin-.t12 bgr_7_0.V_mir1.t0 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X549 GNDA.t191 GNDA.t207 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X550 bgr_7_0.1st_Vout_2.t29 bgr_7_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VOUT-.t115 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 VOUT-.t116 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_14_0.V_source.t15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X554 VOUT+.t120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT+.t15 GNDA.t204 GNDA.t206 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X556 VDDA.t139 two_stage_opamp_dummy_magic_14_0.Y.t47 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X557 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t1 VDDA.t210 VDDA.t212 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X558 VOUT-.t117 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VOUT+.t121 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 bgr_7_0.1st_Vout_1.t30 bgr_7_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 GNDA.t213 GNDA.t212 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X562 GNDA.t60 VDDA.t203 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X563 a_6810_23838.t1 a_6930_22564.t1 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X564 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 two_stage_opamp_dummy_magic_14_0.Y.t48 GNDA.t51 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X565 VOUT+.t122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 GNDA.t191 GNDA.t208 bgr_7_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X567 VOUT+.t123 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 bgr_7_0.1st_Vout_2.t30 bgr_7_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT+.t11 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 GNDA.t136 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X570 VOUT+.t124 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 GNDA.t161 bgr_7_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 bgr_7_0.Vin-.t4 bgr_7_0.V_TOP.t39 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X573 a_12530_23988.t0 a_12410_22380.t0 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=6
X574 two_stage_opamp_dummy_magic_14_0.Vb3.t4 bgr_7_0.NFET_GATE_10uA.t19 GNDA.t159 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X575 two_stage_opamp_dummy_magic_14_0.VD4.t30 two_stage_opamp_dummy_magic_14_0.Vb3.t21 VDDA.t331 VDDA.t330 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X576 bgr_7_0.1st_Vout_2.t31 bgr_7_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VOUT-.t118 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t313 bgr_7_0.V_mir2.t2 bgr_7_0.V_mir2.t3 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X579 VOUT+.t125 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 bgr_7_0.1st_Vout_1.t31 bgr_7_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_7_0.1st_Vout_2.t32 bgr_7_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 bgr_7_0.V_p_1.t5 VDDA.t413 GNDA.t77 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X583 VDDA.t329 two_stage_opamp_dummy_magic_14_0.Vb3.t22 two_stage_opamp_dummy_magic_14_0.VD3.t32 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X584 VDDA.t202 VDDA.t200 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X585 VOUT+.t126 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 bgr_7_0.PFET_GATE_10uA.t22 VDDA.t315 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X587 VOUT-.t119 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 VOUT-.t120 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 a_13180_23838.t1 a_13060_22630.t0 GNDA.t144 sky130_fd_pr__res_xhigh_po_0p35 l=4
X590 VDDA.t383 two_stage_opamp_dummy_magic_14_0.X.t46 VOUT-.t14 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X591 VOUT+.t127 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 a_14330_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t1 GNDA.t41 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X593 VOUT+.t128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VOUT+.t129 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 two_stage_opamp_dummy_magic_14_0.VD2.t19 VIN+.t9 two_stage_opamp_dummy_magic_14_0.V_source.t36 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X596 two_stage_opamp_dummy_magic_14_0.VD1.t6 two_stage_opamp_dummy_magic_14_0.Vb1.t28 two_stage_opamp_dummy_magic_14_0.X.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X597 bgr_7_0.V_p_1.t7 bgr_7_0.Vin+.t9 bgr_7_0.1st_Vout_1.t7 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X598 VDDA.t108 bgr_7_0.V_mir1.t22 bgr_7_0.1st_Vout_1.t0 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X599 bgr_7_0.V_TOP.t40 VDDA.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 two_stage_opamp_dummy_magic_14_0.VD4.t29 two_stage_opamp_dummy_magic_14_0.Vb3.t23 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X601 two_stage_opamp_dummy_magic_14_0.Vb2_2.t1 two_stage_opamp_dummy_magic_14_0.Vb2.t0 two_stage_opamp_dummy_magic_14_0.Vb2.t1 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X602 VOUT-.t121 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VOUT-.t122 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT-.t123 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_14_0.X.t47 VDDA.t147 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X606 VOUT-.t124 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VDDA.t121 two_stage_opamp_dummy_magic_14_0.Y.t49 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X608 GNDA.t211 GNDA.t209 two_stage_opamp_dummy_magic_14_0.VD1.t18 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X609 VOUT+.t130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VOUT+.t131 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 VDDA.t410 bgr_7_0.PFET_GATE_10uA.t23 bgr_7_0.V_CUR_REF_REG.t2 VDDA.t409 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X612 VOUT-.t2 two_stage_opamp_dummy_magic_14_0.X.t48 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X613 GNDA.t140 two_stage_opamp_dummy_magic_14_0.X.t49 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X614 bgr_7_0.V_TOP.t41 VDDA.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 bgr_7_0.V_p_1.t6 bgr_7_0.Vin+.t10 bgr_7_0.1st_Vout_1.t6 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X616 VDDA.t199 VDDA.t197 bgr_7_0.V_TOP.t6 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X617 VOUT-.t125 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_14_0.Vb2.t2 bgr_7_0.NFET_GATE_10uA.t20 GNDA.t157 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X619 GNDA.t155 bgr_7_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X620 VOUT-.t126 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 VOUT-.t127 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 two_stage_opamp_dummy_magic_14_0.VD3.t20 VDDA.t194 VDDA.t196 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X623 VDDA.t193 VDDA.t191 VOUT+.t12 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X624 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 bgr_7_0.NFET_GATE_10uA.t22 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X625 bgr_7_0.V_TOP.t42 VDDA.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X627 bgr_7_0.V_TOP.t43 VDDA.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 VOUT-.t128 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_14_0.Vb1.t6 two_stage_opamp_dummy_magic_14_0.Vb1.t5 two_stage_opamp_dummy_magic_14_0.Vb1_2.t0 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X630 VOUT-.t129 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VDDA.t299 bgr_7_0.V_mir2.t22 bgr_7_0.1st_Vout_2.t8 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X632 two_stage_opamp_dummy_magic_14_0.VD4.t3 two_stage_opamp_dummy_magic_14_0.Vb2.t29 two_stage_opamp_dummy_magic_14_0.Y.t9 two_stage_opamp_dummy_magic_14_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X633 two_stage_opamp_dummy_magic_14_0.Y.t21 two_stage_opamp_dummy_magic_14_0.Vb1.t29 two_stage_opamp_dummy_magic_14_0.VD2.t14 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X634 VOUT-.t130 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VDDA.t98 bgr_7_0.1st_Vout_1.t32 bgr_7_0.V_TOP.t1 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X636 VOUT+.t132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 VOUT-.t131 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VOUT-.t132 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 GNDA.t203 GNDA.t201 two_stage_opamp_dummy_magic_14_0.V_source.t33 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X640 a_5420_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X641 VOUT+.t133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VOUT+.t134 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 VDDA.t190 VDDA.t188 GNDA.t9 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X644 bgr_7_0.V_TOP.t44 VDDA.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 a_5980_2720.t0 GNDA.t81 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X646 two_stage_opamp_dummy_magic_14_0.VD3.t31 two_stage_opamp_dummy_magic_14_0.Vb3.t24 VDDA.t325 VDDA.t324 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X647 VOUT-.t133 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 VDDA.t149 two_stage_opamp_dummy_magic_14_0.X.t50 VOUT-.t6 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X649 VOUT-.t4 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 GNDA.t106 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X650 two_stage_opamp_dummy_magic_14_0.VD3.t1 two_stage_opamp_dummy_magic_14_0.Vb2.t30 two_stage_opamp_dummy_magic_14_0.X.t20 two_stage_opamp_dummy_magic_14_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X651 bgr_7_0.V_TOP.t45 VDDA.t166 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 bgr_7_0.V_mir2.t1 bgr_7_0.V_mir2.t0 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X653 VDDA.t137 bgr_7_0.V_mir1.t7 bgr_7_0.V_mir1.t8 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X654 two_stage_opamp_dummy_magic_14_0.Vb1.t9 VDDA.t185 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X655 VOUT-.t134 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 two_stage_opamp_dummy_magic_14_0.VD1.t5 two_stage_opamp_dummy_magic_14_0.Vb1.t30 two_stage_opamp_dummy_magic_14_0.X.t3 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X657 VOUT-.t135 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 VOUT-.t136 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 bgr_7_0.V_mir2.t14 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 bgr_7_0.V_p_2.t9 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X660 VOUT+.t135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VOUT+.t136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_7_0.PFET_GATE_10uA.t9 VDDA.t414 GNDA.t78 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X663 VOUT+.t137 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 bgr_7_0.1st_Vout_1.t33 bgr_7_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 two_stage_opamp_dummy_magic_14_0.VD3.t30 two_stage_opamp_dummy_magic_14_0.Vb3.t25 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X666 VOUT-.t137 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 VDDA.t168 bgr_7_0.V_TOP.t46 bgr_7_0.Vin-.t3 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X668 VDDA.t358 GNDA.t198 GNDA.t200 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X669 VDDA.t390 two_stage_opamp_dummy_magic_14_0.Y.t50 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X670 VOUT+.t138 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VOUT-.t7 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X672 two_stage_opamp_dummy_magic_14_0.V_source.t0 VIN-.t9 two_stage_opamp_dummy_magic_14_0.VD1.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X673 VOUT-.t138 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 bgr_7_0.PFET_GATE_10uA.t1 bgr_7_0.1st_Vout_2.t33 VDDA.t376 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X675 VOUT-.t15 two_stage_opamp_dummy_magic_14_0.X.t51 VDDA.t385 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X676 GNDA.t84 two_stage_opamp_dummy_magic_14_0.X.t52 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X677 VOUT+.t139 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 VDDA.t21 bgr_7_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X679 VDDA.t400 two_stage_opamp_dummy_magic_14_0.Y.t51 VOUT+.t17 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X680 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 VDDA.t182 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X681 GNDA.t197 GNDA.t196 two_stage_opamp_dummy_magic_14_0.V_p_mir.t4 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X682 VOUT-.t139 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VDDA.t114 two_stage_opamp_dummy_magic_14_0.Y.t52 VOUT+.t4 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X684 VDDA.t321 two_stage_opamp_dummy_magic_14_0.Vb3.t26 two_stage_opamp_dummy_magic_14_0.VD4.t28 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X685 VOUT-.t140 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 VOUT+.t140 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 VDDA.t7 bgr_7_0.1st_Vout_2.t34 bgr_7_0.PFET_GATE_10uA.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X688 VOUT+.t141 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT+.t142 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 two_stage_opamp_dummy_magic_14_0.Y.t22 GNDA.t193 GNDA.t195 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X691 VOUT+.t143 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VOUT+.t144 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_7_0.1st_Vout_1.t34 bgr_7_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 GNDA.t44 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_14_0.V_source.t14 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X695 bgr_7_0.1st_Vout_2.t35 bgr_7_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 VOUT-.t141 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 GNDA.t46 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_14_0.V_source.t13 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X698 bgr_7_0.V_mir2.t13 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 bgr_7_0.V_p_2.t6 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X699 two_stage_opamp_dummy_magic_14_0.VD3.t29 two_stage_opamp_dummy_magic_14_0.Vb3.t27 VDDA.t319 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X700 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 bgr_7_0.NFET_GATE_10uA.t23 GNDA.t151 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X701 VOUT-.t142 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 VOUT-.t143 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 GNDA.t191 GNDA.t192 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X704 VOUT-.t144 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_14_0.X.t53 GNDA.t304 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X706 VOUT+.t145 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 bgr_7_0.1st_Vout_1.t35 bgr_7_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT-.t145 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VDDA.t371 bgr_7_0.1st_Vout_1.t36 bgr_7_0.V_TOP.t11 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X710 GNDA.t82 two_stage_opamp_dummy_magic_14_0.Y.t53 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X711 GNDA.t79 VDDA.t415 bgr_7_0.V_TOP.t10 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X712 bgr_7_0.V_TOP.t47 VDDA.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 two_stage_opamp_dummy_magic_14_0.VD2.t12 VIN+.t10 two_stage_opamp_dummy_magic_14_0.V_source.t32 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X714 VOUT-.t146 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VDDA.t100 bgr_7_0.V_TOP.t48 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X716 VDDA.t181 VDDA.t179 two_stage_opamp_dummy_magic_14_0.VD4.t26 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X717 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t5 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X718 VOUT+.t146 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VOUT+.t147 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT+.t148 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VOUT-.t147 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.t3 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X723 two_stage_opamp_dummy_magic_14_0.Y.t20 two_stage_opamp_dummy_magic_14_0.VD4.t20 two_stage_opamp_dummy_magic_14_0.VD4.t22 two_stage_opamp_dummy_magic_14_0.VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X724 two_stage_opamp_dummy_magic_14_0.VD1.t4 two_stage_opamp_dummy_magic_14_0.Vb1.t31 two_stage_opamp_dummy_magic_14_0.X.t8 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X725 VOUT-.t148 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 bgr_7_0.V_mir2.t12 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 bgr_7_0.V_p_2.t8 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X727 two_stage_opamp_dummy_magic_14_0.VD2.t9 two_stage_opamp_dummy_magic_14_0.Vb1.t32 two_stage_opamp_dummy_magic_14_0.Y.t15 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X728 VOUT+.t149 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VOUT+.t150 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 VOUT-.t149 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT+.t151 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 VOUT-.t150 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 VOUT-.t151 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_14_0.X.t54 VDDA.t374 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X735 VOUT+.t152 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VOUT-.t152 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VOUT-.t153 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 VDDA.t317 two_stage_opamp_dummy_magic_14_0.Vb3.t28 two_stage_opamp_dummy_magic_14_0.VD3.t28 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X739 two_stage_opamp_dummy_magic_14_0.V_source.t31 VIN-.t10 two_stage_opamp_dummy_magic_14_0.VD1.t17 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X740 bgr_7_0.V_TOP.t49 VDDA.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 VDDA.t176 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X742 two_stage_opamp_dummy_magic_14_0.Vb3.t7 two_stage_opamp_dummy_magic_14_0.Vb2.t31 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X743 two_stage_opamp_dummy_magic_14_0.X.t12 two_stage_opamp_dummy_magic_14_0.VD3.t22 two_stage_opamp_dummy_magic_14_0.VD3.t24 two_stage_opamp_dummy_magic_14_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X744 VOUT+.t153 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VDDA.t119 two_stage_opamp_dummy_magic_14_0.Y.t54 VOUT+.t5 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X746 VOUT-.t154 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT+.t154 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 VOUT-.t155 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 bgr_7_0.1st_Vout_2.t36 bgr_7_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_14_0.V_source.t12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 GNDA.t111 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X751 GNDA.t112 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_14_0.V_p_mir.t2 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X752 VDDA.t9 bgr_7_0.V_mir1.t5 bgr_7_0.V_mir1.t6 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X753 VOUT+.t155 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_14_0.Y.t4 two_stage_opamp_dummy_magic_14_0.Vb2.t32 two_stage_opamp_dummy_magic_14_0.VD4.t1 two_stage_opamp_dummy_magic_14_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X755 VOUT+.t156 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VOUT-.t156 two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_7_0.NFET_GATE_10uA.n19 bgr_7_0.NFET_GATE_10uA.t3 384.967
R1 bgr_7_0.NFET_GATE_10uA.n10 bgr_7_0.NFET_GATE_10uA.t10 369.534
R2 bgr_7_0.NFET_GATE_10uA.n9 bgr_7_0.NFET_GATE_10uA.t22 369.534
R3 bgr_7_0.NFET_GATE_10uA.n7 bgr_7_0.NFET_GATE_10uA.t7 369.534
R4 bgr_7_0.NFET_GATE_10uA.n4 bgr_7_0.NFET_GATE_10uA.t16 369.534
R5 bgr_7_0.NFET_GATE_10uA.n1 bgr_7_0.NFET_GATE_10uA.t12 369.534
R6 bgr_7_0.NFET_GATE_10uA.t3 bgr_7_0.NFET_GATE_10uA.n18 369.534
R7 bgr_7_0.NFET_GATE_10uA bgr_7_0.NFET_GATE_10uA.n20 366.147
R8 bgr_7_0.NFET_GATE_10uA.n12 bgr_7_0.NFET_GATE_10uA.t9 192.8
R9 bgr_7_0.NFET_GATE_10uA.n11 bgr_7_0.NFET_GATE_10uA.t17 192.8
R10 bgr_7_0.NFET_GATE_10uA.n10 bgr_7_0.NFET_GATE_10uA.t23 192.8
R11 bgr_7_0.NFET_GATE_10uA.n9 bgr_7_0.NFET_GATE_10uA.t11 192.8
R12 bgr_7_0.NFET_GATE_10uA.n7 bgr_7_0.NFET_GATE_10uA.t20 192.8
R13 bgr_7_0.NFET_GATE_10uA.n4 bgr_7_0.NFET_GATE_10uA.t21 192.8
R14 bgr_7_0.NFET_GATE_10uA.n5 bgr_7_0.NFET_GATE_10uA.t8 192.8
R15 bgr_7_0.NFET_GATE_10uA.n6 bgr_7_0.NFET_GATE_10uA.t15 192.8
R16 bgr_7_0.NFET_GATE_10uA.n3 bgr_7_0.NFET_GATE_10uA.t19 192.8
R17 bgr_7_0.NFET_GATE_10uA.n2 bgr_7_0.NFET_GATE_10uA.t5 192.8
R18 bgr_7_0.NFET_GATE_10uA.n1 bgr_7_0.NFET_GATE_10uA.t13 192.8
R19 bgr_7_0.NFET_GATE_10uA.n18 bgr_7_0.NFET_GATE_10uA.t18 192.8
R20 bgr_7_0.NFET_GATE_10uA.n17 bgr_7_0.NFET_GATE_10uA.t6 192.8
R21 bgr_7_0.NFET_GATE_10uA.n16 bgr_7_0.NFET_GATE_10uA.t14 192.8
R22 bgr_7_0.NFET_GATE_10uA.n12 bgr_7_0.NFET_GATE_10uA.n11 176.733
R23 bgr_7_0.NFET_GATE_10uA.n11 bgr_7_0.NFET_GATE_10uA.n10 176.733
R24 bgr_7_0.NFET_GATE_10uA.n5 bgr_7_0.NFET_GATE_10uA.n4 176.733
R25 bgr_7_0.NFET_GATE_10uA.n6 bgr_7_0.NFET_GATE_10uA.n5 176.733
R26 bgr_7_0.NFET_GATE_10uA.n3 bgr_7_0.NFET_GATE_10uA.n2 176.733
R27 bgr_7_0.NFET_GATE_10uA.n2 bgr_7_0.NFET_GATE_10uA.n1 176.733
R28 bgr_7_0.NFET_GATE_10uA.n18 bgr_7_0.NFET_GATE_10uA.n17 176.733
R29 bgr_7_0.NFET_GATE_10uA.n17 bgr_7_0.NFET_GATE_10uA.n16 176.733
R30 bgr_7_0.NFET_GATE_10uA.n14 bgr_7_0.NFET_GATE_10uA.n13 169.852
R31 bgr_7_0.NFET_GATE_10uA.n14 bgr_7_0.NFET_GATE_10uA.n8 169.852
R32 bgr_7_0.NFET_GATE_10uA.n15 bgr_7_0.NFET_GATE_10uA.n14 166.133
R33 bgr_7_0.NFET_GATE_10uA.n19 bgr_7_0.NFET_GATE_10uA.n0 126.877
R34 bgr_7_0.NFET_GATE_10uA.n13 bgr_7_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_7_0.NFET_GATE_10uA.n13 bgr_7_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_7_0.NFET_GATE_10uA.n8 bgr_7_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_7_0.NFET_GATE_10uA.n8 bgr_7_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_7_0.NFET_GATE_10uA.n15 bgr_7_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_7_0.NFET_GATE_10uA.n16 bgr_7_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_7_0.NFET_GATE_10uA.n20 bgr_7_0.NFET_GATE_10uA.t1 39.4005
R41 bgr_7_0.NFET_GATE_10uA.n20 bgr_7_0.NFET_GATE_10uA.t2 39.4005
R42 bgr_7_0.NFET_GATE_10uA bgr_7_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_7_0.NFET_GATE_10uA.n0 bgr_7_0.NFET_GATE_10uA.t0 24.0005
R44 bgr_7_0.NFET_GATE_10uA.n0 bgr_7_0.NFET_GATE_10uA.t4 24.0005
R45 two_stage_opamp_dummy_magic_14_0.Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb3.t12 650.511
R46 two_stage_opamp_dummy_magic_14_0.Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb3.t15 611.739
R47 two_stage_opamp_dummy_magic_14_0.Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb3.t23 611.739
R48 two_stage_opamp_dummy_magic_14_0.Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb3.t28 611.739
R49 two_stage_opamp_dummy_magic_14_0.Vb3.n6 two_stage_opamp_dummy_magic_14_0.Vb3.t11 611.739
R50 two_stage_opamp_dummy_magic_14_0.Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb3.t19 421.75
R51 two_stage_opamp_dummy_magic_14_0.Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb3.t17 421.75
R52 two_stage_opamp_dummy_magic_14_0.Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb3.t21 421.75
R53 two_stage_opamp_dummy_magic_14_0.Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb3.t26 421.75
R54 two_stage_opamp_dummy_magic_14_0.Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb3.t18 421.75
R55 two_stage_opamp_dummy_magic_14_0.Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb3.t14 421.75
R56 two_stage_opamp_dummy_magic_14_0.Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb3.t10 421.75
R57 two_stage_opamp_dummy_magic_14_0.Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb3.t8 421.75
R58 two_stage_opamp_dummy_magic_14_0.Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb3.t25 421.75
R59 two_stage_opamp_dummy_magic_14_0.Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb3.t13 421.75
R60 two_stage_opamp_dummy_magic_14_0.Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb3.t16 421.75
R61 two_stage_opamp_dummy_magic_14_0.Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb3.t20 421.75
R62 two_stage_opamp_dummy_magic_14_0.Vb3.n6 two_stage_opamp_dummy_magic_14_0.Vb3.t9 421.75
R63 two_stage_opamp_dummy_magic_14_0.Vb3.n7 two_stage_opamp_dummy_magic_14_0.Vb3.t27 421.75
R64 two_stage_opamp_dummy_magic_14_0.Vb3.n8 two_stage_opamp_dummy_magic_14_0.Vb3.t22 421.75
R65 two_stage_opamp_dummy_magic_14_0.Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb3.t24 421.75
R66 two_stage_opamp_dummy_magic_14_0.Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb3.n23 176.685
R67 two_stage_opamp_dummy_magic_14_0.Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb3.n14 176.124
R68 two_stage_opamp_dummy_magic_14_0.Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_14_0.Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb3.n20 167.094
R70 two_stage_opamp_dummy_magic_14_0.Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb3.n21 167.094
R71 two_stage_opamp_dummy_magic_14_0.Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb3.n15 167.094
R72 two_stage_opamp_dummy_magic_14_0.Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb3.n16 167.094
R73 two_stage_opamp_dummy_magic_14_0.Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb3.n17 167.094
R74 two_stage_opamp_dummy_magic_14_0.Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb3.n10 167.094
R75 two_stage_opamp_dummy_magic_14_0.Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb3.n11 167.094
R76 two_stage_opamp_dummy_magic_14_0.Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb3.n12 167.094
R77 two_stage_opamp_dummy_magic_14_0.Vb3.n7 two_stage_opamp_dummy_magic_14_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_14_0.Vb3.n8 two_stage_opamp_dummy_magic_14_0.Vb3.n7 167.094
R79 two_stage_opamp_dummy_magic_14_0.Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb3.n8 167.094
R80 two_stage_opamp_dummy_magic_14_0.Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb3.n5 161.631
R81 two_stage_opamp_dummy_magic_14_0.Vb3.n2 two_stage_opamp_dummy_magic_14_0.Vb3.n0 139.639
R82 two_stage_opamp_dummy_magic_14_0.Vb3.n2 two_stage_opamp_dummy_magic_14_0.Vb3.n1 139.638
R83 two_stage_opamp_dummy_magic_14_0.Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb3.n3 134.577
R84 two_stage_opamp_dummy_magic_14_0.Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb3.n22 49.8072
R85 two_stage_opamp_dummy_magic_14_0.Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb3.n18 49.8072
R86 two_stage_opamp_dummy_magic_14_0.Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb3.n13 49.8072
R87 two_stage_opamp_dummy_magic_14_0.Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb3.n9 49.8072
R88 bgr_7_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb3.n26 48.0943
R89 bgr_7_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb3.n4 41.063
R90 two_stage_opamp_dummy_magic_14_0.Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb3.t1 24.0005
R91 two_stage_opamp_dummy_magic_14_0.Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb3.t3 24.0005
R92 two_stage_opamp_dummy_magic_14_0.Vb3.n1 two_stage_opamp_dummy_magic_14_0.Vb3.t5 24.0005
R93 two_stage_opamp_dummy_magic_14_0.Vb3.n1 two_stage_opamp_dummy_magic_14_0.Vb3.t0 24.0005
R94 two_stage_opamp_dummy_magic_14_0.Vb3.n0 two_stage_opamp_dummy_magic_14_0.Vb3.t2 24.0005
R95 two_stage_opamp_dummy_magic_14_0.Vb3.n0 two_stage_opamp_dummy_magic_14_0.Vb3.t4 24.0005
R96 two_stage_opamp_dummy_magic_14_0.Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb3.n24 13.7349
R97 two_stage_opamp_dummy_magic_14_0.Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb3.t6 11.2576
R98 two_stage_opamp_dummy_magic_14_0.Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb3.t7 11.2576
R99 two_stage_opamp_dummy_magic_14_0.Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb3.n2 4.5005
R100 two_stage_opamp_dummy_magic_14_0.Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb3.n25 1.438
R101 GNDA.n2166 GNDA.n99 89432.2
R102 GNDA.n2164 GNDA.n99 87364.4
R103 GNDA.n2415 GNDA.n88 21966.8
R104 GNDA.n2629 GNDA.n10 21966.8
R105 GNDA.n2170 GNDA.n91 14422.9
R106 GNDA.n2631 GNDA.n2630 14422.9
R107 GNDA.n2169 GNDA.n92 13534.7
R108 GNDA.n98 GNDA.n97 13528.5
R109 GNDA.n96 GNDA.n7 13200
R110 GNDA.n2171 GNDA.n7 12089.3
R111 GNDA.n2632 GNDA.n7 12089.3
R112 GNDA.n2164 GNDA.n2163 11953.3
R113 GNDA.n2163 GNDA.n100 11949.5
R114 GNDA.n97 GNDA.n96 11178.4
R115 GNDA.n168 GNDA.n100 10235.4
R116 GNDA.n97 GNDA.n8 9632.43
R117 GNDA.n9 GNDA.n8 9001.83
R118 GNDA.n2165 GNDA.n94 8901.32
R119 GNDA.n168 GNDA.n94 8812.35
R120 GNDA.n2167 GNDA.n2166 8661.12
R121 GNDA.n2631 GNDA.n8 7750.87
R122 GNDA.n2170 GNDA.n2169 7548.93
R123 GNDA.n2169 GNDA.n2168 6567.6
R124 GNDA.n99 GNDA.n93 5523.81
R125 GNDA.n98 GNDA.n92 4761.61
R126 GNDA.n2165 GNDA.n2164 4106.67
R127 GNDA.n2163 GNDA.n2162 3974.19
R128 GNDA.n170 GNDA.n100 3962.24
R129 GNDA.n96 GNDA.n92 3961.87
R130 GNDA.n2168 GNDA.n91 2972.3
R131 GNDA.n2167 GNDA.n94 2531.14
R132 GNDA.n2168 GNDA.n93 2522.64
R133 GNDA.n2630 GNDA.n9 2503.88
R134 GNDA.n2167 GNDA.n98 2315.79
R135 GNDA.n2632 GNDA.n2631 1986.41
R136 GNDA.n2171 GNDA.n2170 1986.41
R137 GNDA.t41 GNDA.n88 1966.49
R138 GNDA.n2166 GNDA.n2165 1863.53
R139 GNDA.n2168 GNDA.n2167 1693.44
R140 GNDA.n2167 GNDA.n95 1647.44
R141 GNDA.t15 GNDA.t81 1622.45
R142 GNDA.n169 GNDA.n95 1397
R143 GNDA.n1262 GNDA.n1067 1336.64
R144 GNDA.t147 GNDA.n170 1225.15
R145 GNDA.n1237 GNDA.n1236 1214.72
R146 GNDA.n1236 GNDA.n1235 1214.72
R147 GNDA.n1235 GNDA.n1206 1214.72
R148 GNDA.n1229 GNDA.n1206 1214.72
R149 GNDA.n1229 GNDA.n238 1214.72
R150 GNDA.n1218 GNDA.n237 1214.72
R151 GNDA.n1222 GNDA.n1218 1214.72
R152 GNDA.n1222 GNDA.n1221 1214.72
R153 GNDA.n1221 GNDA.n1220 1214.72
R154 GNDA.n1220 GNDA.n236 1214.72
R155 GNDA.n1139 GNDA.n1104 1214.72
R156 GNDA.n1139 GNDA.n1138 1214.72
R157 GNDA.n1138 GNDA.n1137 1214.72
R158 GNDA.n1137 GNDA.n1112 1214.72
R159 GNDA.n1112 GNDA.n230 1214.72
R160 GNDA.n1129 GNDA.n229 1214.72
R161 GNDA.n1129 GNDA.n1128 1214.72
R162 GNDA.n1128 GNDA.n1127 1214.72
R163 GNDA.n1127 GNDA.n1123 1214.72
R164 GNDA.n1123 GNDA.n228 1214.72
R165 GNDA.n2023 GNDA.n2022 1212.88
R166 GNDA.n2136 GNDA.n2135 1185.07
R167 GNDA.n2135 GNDA.n128 1185.07
R168 GNDA.n170 GNDA.n169 937.1
R169 GNDA.n91 GNDA.t146 927.827
R170 GNDA.n2629 GNDA.t15 845.198
R171 GNDA.n169 GNDA.n168 832.433
R172 GNDA.t191 GNDA.n238 823.313
R173 GNDA.t191 GNDA.n230 823.313
R174 GNDA.n2630 GNDA.t99 803.766
R175 GNDA.n2305 GNDA.t264 762.534
R176 GNDA.n2173 GNDA.t254 762.534
R177 GNDA.n2615 GNDA.t281 762.534
R178 GNDA.n2617 GNDA.t198 762.534
R179 GNDA.t50 GNDA.n93 744.481
R180 GNDA.t146 GNDA.n88 726.957
R181 GNDA.n2627 GNDA.n2626 692.506
R182 GNDA.n2611 GNDA.n2610 692.506
R183 GNDA.n2301 GNDA.n2300 692.506
R184 GNDA.n2212 GNDA.n2211 692.506
R185 GNDA.n2599 GNDA.n2598 692.506
R186 GNDA.n2538 GNDA.n2535 692.506
R187 GNDA.n2289 GNDA.n2288 692.506
R188 GNDA.n2253 GNDA.n2252 692.506
R189 GNDA.n2387 GNDA.n2382 691.179
R190 GNDA.n2460 GNDA.n57 691.179
R191 GNDA.n2132 GNDA.n2131 686.717
R192 GNDA.n46 GNDA.n45 686.717
R193 GNDA.n2471 GNDA.n2470 686.717
R194 GNDA.n2482 GNDA.n2481 686.717
R195 GNDA.n2441 GNDA.n2440 686.717
R196 GNDA.n2424 GNDA.n2423 686.717
R197 GNDA.n2414 GNDA.n2413 686.717
R198 GNDA.n2458 GNDA.n2457 686.717
R199 GNDA.n2381 GNDA.n2380 686.717
R200 GNDA.n2313 GNDA.n2312 686.717
R201 GNDA.n2347 GNDA.n2346 686.717
R202 GNDA.n2641 GNDA.n2640 686.717
R203 GNDA.n65 GNDA.n64 686.717
R204 GNDA.n2024 GNDA.n2023 686.717
R205 GNDA.n2024 GNDA.n171 686.717
R206 GNDA.n2354 GNDA.n2353 686.717
R207 GNDA.n2320 GNDA.n2319 686.717
R208 GNDA.n2365 GNDA.n2364 686.717
R209 GNDA.n2402 GNDA.n2395 686.717
R210 GNDA.n2490 GNDA.n2489 686.717
R211 GNDA.n2501 GNDA.n2494 686.717
R212 GNDA.n2433 GNDA.n68 686.717
R213 GNDA.n53 GNDA.n52 686.717
R214 GNDA.n2123 GNDA.n136 686.717
R215 GNDA.n216 GNDA.n209 686.717
R216 GNDA.n2321 GNDA.t220 682.201
R217 GNDA.n1094 GNDA.n1093 669.307
R218 GNDA.n2355 GNDA.t201 650.067
R219 GNDA.n2391 GNDA.t196 650.067
R220 GNDA.n2448 GNDA.t262 650.067
R221 GNDA.n2432 GNDA.t237 650.067
R222 GNDA.n54 GNDA.t284 650.067
R223 GNDA.t99 GNDA.n2629 629.755
R224 GNDA.n2394 GNDA.t217 627.976
R225 GNDA.n2491 GNDA.t269 627.976
R226 GNDA.n309 GNDA.n206 585.001
R227 GNDA.n1931 GNDA.n1930 585.001
R228 GNDA.n1957 GNDA.n1956 585.001
R229 GNDA.n1943 GNDA.n306 585.001
R230 GNDA.n1940 GNDA.n1939 585.001
R231 GNDA.n2031 GNDA.n2030 585.001
R232 GNDA.n2019 GNDA.n189 585
R233 GNDA.n2018 GNDA.n193 585
R234 GNDA.n2018 GNDA.n2017 585
R235 GNDA.n2012 GNDA.n192 585
R236 GNDA.n2016 GNDA.n192 585
R237 GNDA.n2014 GNDA.n2013 585
R238 GNDA.n2015 GNDA.n2014 585
R239 GNDA.n2011 GNDA.n195 585
R240 GNDA.n195 GNDA.n194 585
R241 GNDA.n2010 GNDA.n2009 585
R242 GNDA.n2009 GNDA.n139 585
R243 GNDA.n2008 GNDA.n196 585
R244 GNDA.n2008 GNDA.n138 585
R245 GNDA.n2007 GNDA.n198 585
R246 GNDA.n2007 GNDA.n2006 585
R247 GNDA.n2001 GNDA.n197 585
R248 GNDA.n2005 GNDA.n197 585
R249 GNDA.n2003 GNDA.n2002 585
R250 GNDA.n2004 GNDA.n2003 585
R251 GNDA.n2000 GNDA.n200 585
R252 GNDA.n200 GNDA.n199 585
R253 GNDA.n1999 GNDA.n1998 585
R254 GNDA.n1998 GNDA.n1997 585
R255 GNDA.n2022 GNDA.n2021 585
R256 GNDA.n626 GNDA.n625 585
R257 GNDA.n1038 GNDA.n622 585
R258 GNDA.n622 GNDA.n621 585
R259 GNDA.n1040 GNDA.n1039 585
R260 GNDA.n1041 GNDA.n1040 585
R261 GNDA.n623 GNDA.n620 585
R262 GNDA.n1042 GNDA.n620 585
R263 GNDA.n1044 GNDA.n619 585
R264 GNDA.n1044 GNDA.n1043 585
R265 GNDA.n1046 GNDA.n1045 585
R266 GNDA.n1045 GNDA.n232 585
R267 GNDA.n1047 GNDA.n618 585
R268 GNDA.n618 GNDA.n233 585
R269 GNDA.n1049 GNDA.n1048 585
R270 GNDA.n1050 GNDA.n1049 585
R271 GNDA.n617 GNDA.n616 585
R272 GNDA.n1051 GNDA.n617 585
R273 GNDA.n1054 GNDA.n1053 585
R274 GNDA.n1053 GNDA.n1052 585
R275 GNDA.n1055 GNDA.n523 585
R276 GNDA.n523 GNDA.n521 585
R277 GNDA.n1057 GNDA.n1056 585
R278 GNDA.n1058 GNDA.n1057 585
R279 GNDA.n1035 GNDA.n231 585
R280 GNDA.n1288 GNDA.n1287 585
R281 GNDA.n1290 GNDA.n1059 585
R282 GNDA.n1282 GNDA.n1060 585
R283 GNDA.n1286 GNDA.n1060 585
R284 GNDA.n1284 GNDA.n1283 585
R285 GNDA.n1285 GNDA.n1284 585
R286 GNDA.n1281 GNDA.n1062 585
R287 GNDA.n1062 GNDA.n1061 585
R288 GNDA.n1280 GNDA.n1279 585
R289 GNDA.n1279 GNDA.n1278 585
R290 GNDA.n1277 GNDA.n1063 585
R291 GNDA.n1277 GNDA.n234 585
R292 GNDA.n1276 GNDA.n1275 585
R293 GNDA.n1276 GNDA.n235 585
R294 GNDA.n1274 GNDA.n1064 585
R295 GNDA.n1270 GNDA.n1064 585
R296 GNDA.n1273 GNDA.n1272 585
R297 GNDA.n1272 GNDA.n1271 585
R298 GNDA.n1066 GNDA.n1065 585
R299 GNDA.n1269 GNDA.n1066 585
R300 GNDA.n1267 GNDA.n1266 585
R301 GNDA.n1268 GNDA.n1267 585
R302 GNDA.n1265 GNDA.n1068 585
R303 GNDA.n1068 GNDA.n1067 585
R304 GNDA.n1389 GNDA.n1388 585
R305 GNDA.n1389 GNDA.n236 585
R306 GNDA.n497 GNDA.n496 585
R307 GNDA.n1220 GNDA.n496 585
R308 GNDA.n1219 GNDA.n1216 585
R309 GNDA.n1221 GNDA.n1219 585
R310 GNDA.n1224 GNDA.n1215 585
R311 GNDA.n1222 GNDA.n1215 585
R312 GNDA.n1225 GNDA.n1214 585
R313 GNDA.n1218 GNDA.n1214 585
R314 GNDA.n1226 GNDA.n1213 585
R315 GNDA.n1213 GNDA.n237 585
R316 GNDA.n1212 GNDA.n1210 585
R317 GNDA.n1212 GNDA.n238 585
R318 GNDA.n1231 GNDA.n1209 585
R319 GNDA.n1229 GNDA.n1209 585
R320 GNDA.n1232 GNDA.n1208 585
R321 GNDA.n1208 GNDA.n1206 585
R322 GNDA.n1233 GNDA.n1205 585
R323 GNDA.n1235 GNDA.n1205 585
R324 GNDA.n1204 GNDA.n1083 585
R325 GNDA.n1236 GNDA.n1204 585
R326 GNDA.n1239 GNDA.n1082 585
R327 GNDA.n1237 GNDA.n1082 585
R328 GNDA.n1239 GNDA.n1238 585
R329 GNDA.n1238 GNDA.n1237 585
R330 GNDA.n1084 GNDA.n1083 585
R331 GNDA.n1236 GNDA.n1084 585
R332 GNDA.n1234 GNDA.n1233 585
R333 GNDA.n1235 GNDA.n1234 585
R334 GNDA.n1232 GNDA.n1207 585
R335 GNDA.n1207 GNDA.n1206 585
R336 GNDA.n1231 GNDA.n1230 585
R337 GNDA.n1230 GNDA.n1229 585
R338 GNDA.n1228 GNDA.n1210 585
R339 GNDA.n1228 GNDA.n238 585
R340 GNDA.n1227 GNDA.n1226 585
R341 GNDA.n1227 GNDA.n237 585
R342 GNDA.n1225 GNDA.n1211 585
R343 GNDA.n1218 GNDA.n1211 585
R344 GNDA.n1224 GNDA.n1223 585
R345 GNDA.n1223 GNDA.n1222 585
R346 GNDA.n1217 GNDA.n1216 585
R347 GNDA.n1221 GNDA.n1217 585
R348 GNDA.n498 GNDA.n497 585
R349 GNDA.n1220 GNDA.n498 585
R350 GNDA.n1388 GNDA.n1387 585
R351 GNDA.n1387 GNDA.n236 585
R352 GNDA.n571 GNDA.n570 585
R353 GNDA.n572 GNDA.n568 585
R354 GNDA.n567 GNDA.n565 585
R355 GNDA.n578 GNDA.n564 585
R356 GNDA.n579 GNDA.n563 585
R357 GNDA.n580 GNDA.n561 585
R358 GNDA.n560 GNDA.n557 585
R359 GNDA.n585 GNDA.n556 585
R360 GNDA.n586 GNDA.n555 585
R361 GNDA.n553 GNDA.n551 585
R362 GNDA.n590 GNDA.n550 585
R363 GNDA.n591 GNDA.n548 585
R364 GNDA.n592 GNDA.n591 585
R365 GNDA.n590 GNDA.n589 585
R366 GNDA.n588 GNDA.n551 585
R367 GNDA.n588 GNDA.n239 585
R368 GNDA.n587 GNDA.n586 585
R369 GNDA.n585 GNDA.n584 585
R370 GNDA.n583 GNDA.n557 585
R371 GNDA.n581 GNDA.n580 585
R372 GNDA.n579 GNDA.n558 585
R373 GNDA.n578 GNDA.n577 585
R374 GNDA.n575 GNDA.n565 585
R375 GNDA.n573 GNDA.n572 585
R376 GNDA.n571 GNDA.n293 585
R377 GNDA.n293 GNDA.n239 585
R378 GNDA.n1844 GNDA.n1843 585
R379 GNDA.n1780 GNDA.n1779 585
R380 GNDA.n1782 GNDA.n1781 585
R381 GNDA.n1836 GNDA.n1835 585
R382 GNDA.n1834 GNDA.n1833 585
R383 GNDA.n1832 GNDA.n1786 585
R384 GNDA.n1785 GNDA.n1784 585
R385 GNDA.n1826 GNDA.n1825 585
R386 GNDA.n1824 GNDA.n1823 585
R387 GNDA.n1822 GNDA.n1789 585
R388 GNDA.n1788 GNDA.n300 585
R389 GNDA.n1960 GNDA.n297 585
R390 GNDA.n1817 GNDA.n297 585
R391 GNDA.n1819 GNDA.n1788 585
R392 GNDA.n1822 GNDA.n1821 585
R393 GNDA.n1823 GNDA.n1787 585
R394 GNDA.n1827 GNDA.n1826 585
R395 GNDA.n1829 GNDA.n1784 585
R396 GNDA.n1832 GNDA.n1831 585
R397 GNDA.n1833 GNDA.n1783 585
R398 GNDA.n1837 GNDA.n1836 585
R399 GNDA.n1839 GNDA.n1782 585
R400 GNDA.n1840 GNDA.n1779 585
R401 GNDA.n1843 GNDA.n1842 585
R402 GNDA.n1927 GNDA.n319 585
R403 GNDA.n1925 GNDA.n1924 585
R404 GNDA.n321 GNDA.n320 585
R405 GNDA.n1669 GNDA.n1668 585
R406 GNDA.n1674 GNDA.n1666 585
R407 GNDA.n1675 GNDA.n1664 585
R408 GNDA.n1676 GNDA.n1663 585
R409 GNDA.n1661 GNDA.n1659 585
R410 GNDA.n1681 GNDA.n1658 585
R411 GNDA.n1682 GNDA.n1656 585
R412 GNDA.n1655 GNDA.n1627 585
R413 GNDA.n1687 GNDA.n1625 585
R414 GNDA.n1687 GNDA.n1686 585
R415 GNDA.n1684 GNDA.n1627 585
R416 GNDA.n1683 GNDA.n1682 585
R417 GNDA.n1681 GNDA.n1680 585
R418 GNDA.n1679 GNDA.n1659 585
R419 GNDA.n1677 GNDA.n1676 585
R420 GNDA.n1675 GNDA.n1660 585
R421 GNDA.n1674 GNDA.n1673 585
R422 GNDA.n1671 GNDA.n1669 585
R423 GNDA.n322 GNDA.n321 585
R424 GNDA.n1924 GNDA.n1923 585
R425 GNDA.n1921 GNDA.n319 585
R426 GNDA.n1969 GNDA.n287 585
R427 GNDA.n1970 GNDA.n278 585
R428 GNDA.n1973 GNDA.n277 585
R429 GNDA.n1974 GNDA.n276 585
R430 GNDA.n1977 GNDA.n275 585
R431 GNDA.n1978 GNDA.n274 585
R432 GNDA.n1981 GNDA.n273 585
R433 GNDA.n1983 GNDA.n272 585
R434 GNDA.n1984 GNDA.n271 585
R435 GNDA.n1985 GNDA.n270 585
R436 GNDA.n279 GNDA.n262 585
R437 GNDA.n1991 GNDA.n258 585
R438 GNDA.n1991 GNDA.n1990 585
R439 GNDA.n264 GNDA.n262 585
R440 GNDA.n1986 GNDA.n1985 585
R441 GNDA.n1984 GNDA.n269 585
R442 GNDA.n1983 GNDA.n1982 585
R443 GNDA.n1981 GNDA.n1980 585
R444 GNDA.n1979 GNDA.n1978 585
R445 GNDA.n1977 GNDA.n1976 585
R446 GNDA.n1975 GNDA.n1974 585
R447 GNDA.n1973 GNDA.n1972 585
R448 GNDA.n1971 GNDA.n1970 585
R449 GNDA.n1969 GNDA.n1968 585
R450 GNDA.n1489 GNDA.n1488 585
R451 GNDA.n1489 GNDA.n228 585
R452 GNDA.n471 GNDA.n470 585
R453 GNDA.n1123 GNDA.n470 585
R454 GNDA.n1125 GNDA.n1122 585
R455 GNDA.n1127 GNDA.n1122 585
R456 GNDA.n1124 GNDA.n1121 585
R457 GNDA.n1128 GNDA.n1121 585
R458 GNDA.n1120 GNDA.n1118 585
R459 GNDA.n1129 GNDA.n1120 585
R460 GNDA.n1119 GNDA.n1116 585
R461 GNDA.n1119 GNDA.n229 585
R462 GNDA.n1133 GNDA.n1115 585
R463 GNDA.n1115 GNDA.n230 585
R464 GNDA.n1134 GNDA.n1114 585
R465 GNDA.n1114 GNDA.n1112 585
R466 GNDA.n1135 GNDA.n1111 585
R467 GNDA.n1137 GNDA.n1111 585
R468 GNDA.n1110 GNDA.n1108 585
R469 GNDA.n1138 GNDA.n1110 585
R470 GNDA.n1141 GNDA.n1107 585
R471 GNDA.n1139 GNDA.n1107 585
R472 GNDA.n1143 GNDA.n1142 585
R473 GNDA.n1143 GNDA.n1104 585
R474 GNDA.n1142 GNDA.n1103 585
R475 GNDA.n1104 GNDA.n1103 585
R476 GNDA.n1141 GNDA.n1140 585
R477 GNDA.n1140 GNDA.n1139 585
R478 GNDA.n1109 GNDA.n1108 585
R479 GNDA.n1138 GNDA.n1109 585
R480 GNDA.n1136 GNDA.n1135 585
R481 GNDA.n1137 GNDA.n1136 585
R482 GNDA.n1134 GNDA.n1113 585
R483 GNDA.n1113 GNDA.n1112 585
R484 GNDA.n1133 GNDA.n1132 585
R485 GNDA.n1132 GNDA.n230 585
R486 GNDA.n1131 GNDA.n1116 585
R487 GNDA.n1131 GNDA.n229 585
R488 GNDA.n1130 GNDA.n1118 585
R489 GNDA.n1130 GNDA.n1129 585
R490 GNDA.n1124 GNDA.n1117 585
R491 GNDA.n1128 GNDA.n1117 585
R492 GNDA.n1126 GNDA.n1125 585
R493 GNDA.n1127 GNDA.n1126 585
R494 GNDA.n472 GNDA.n471 585
R495 GNDA.n1123 GNDA.n472 585
R496 GNDA.n1488 GNDA.n1487 585
R497 GNDA.n1487 GNDA.n228 585
R498 GNDA.n1173 GNDA.n1172 585
R499 GNDA.n1174 GNDA.n1173 585
R500 GNDA.n1171 GNDA.n1106 585
R501 GNDA.n1106 GNDA.n1105 585
R502 GNDA.n1170 GNDA.n1169 585
R503 GNDA.n1169 GNDA.n1168 585
R504 GNDA.n1145 GNDA.n1144 585
R505 GNDA.n1167 GNDA.n1145 585
R506 GNDA.n1165 GNDA.n1164 585
R507 GNDA.n1166 GNDA.n1165 585
R508 GNDA.n1163 GNDA.n1147 585
R509 GNDA.n1147 GNDA.n1146 585
R510 GNDA.n1162 GNDA.n1161 585
R511 GNDA.n1161 GNDA.n1160 585
R512 GNDA.n1149 GNDA.n1148 585
R513 GNDA.n1159 GNDA.n1149 585
R514 GNDA.n1157 GNDA.n1156 585
R515 GNDA.n1158 GNDA.n1157 585
R516 GNDA.n1155 GNDA.n1151 585
R517 GNDA.n1151 GNDA.n1150 585
R518 GNDA.n1154 GNDA.n1153 585
R519 GNDA.n1153 GNDA.n1152 585
R520 GNDA.n427 GNDA.n426 585
R521 GNDA.n426 GNDA.n227 585
R522 GNDA.n1201 GNDA.n1081 585
R523 GNDA.n1202 GNDA.n1201 585
R524 GNDA.n1200 GNDA.n1199 585
R525 GNDA.n1200 GNDA.n1085 585
R526 GNDA.n1198 GNDA.n1086 585
R527 GNDA.n1194 GNDA.n1086 585
R528 GNDA.n1197 GNDA.n1196 585
R529 GNDA.n1196 GNDA.n1195 585
R530 GNDA.n1088 GNDA.n1087 585
R531 GNDA.n1193 GNDA.n1088 585
R532 GNDA.n1191 GNDA.n1190 585
R533 GNDA.n1192 GNDA.n1191 585
R534 GNDA.n1188 GNDA.n1089 585
R535 GNDA.n1184 GNDA.n1089 585
R536 GNDA.n1187 GNDA.n1186 585
R537 GNDA.n1186 GNDA.n1185 585
R538 GNDA.n1099 GNDA.n1098 585
R539 GNDA.n1183 GNDA.n1099 585
R540 GNDA.n1181 GNDA.n1180 585
R541 GNDA.n1182 GNDA.n1181 585
R542 GNDA.n1179 GNDA.n1101 585
R543 GNDA.n1101 GNDA.n1100 585
R544 GNDA.n1178 GNDA.n1177 585
R545 GNDA.n1177 GNDA.n1176 585
R546 GNDA.n1264 GNDA.n1263 585
R547 GNDA.n1263 GNDA.n1262 585
R548 GNDA.n1070 GNDA.n1069 585
R549 GNDA.n1261 GNDA.n1070 585
R550 GNDA.n1259 GNDA.n1258 585
R551 GNDA.n1260 GNDA.n1259 585
R552 GNDA.n1257 GNDA.n1072 585
R553 GNDA.n1072 GNDA.n1071 585
R554 GNDA.n1256 GNDA.n1255 585
R555 GNDA.n1255 GNDA.n1254 585
R556 GNDA.n1074 GNDA.n1073 585
R557 GNDA.n1253 GNDA.n1074 585
R558 GNDA.n1251 GNDA.n1250 585
R559 GNDA.n1252 GNDA.n1251 585
R560 GNDA.n1249 GNDA.n1076 585
R561 GNDA.n1076 GNDA.n1075 585
R562 GNDA.n1248 GNDA.n1247 585
R563 GNDA.n1247 GNDA.n1246 585
R564 GNDA.n1078 GNDA.n1077 585
R565 GNDA.n1245 GNDA.n1078 585
R566 GNDA.n1243 GNDA.n1242 585
R567 GNDA.n1244 GNDA.n1243 585
R568 GNDA.n1241 GNDA.n1080 585
R569 GNDA.n1080 GNDA.n1079 585
R570 GNDA.n1095 GNDA.n1090 585
R571 GNDA.n1097 GNDA.n1096 585
R572 GNDA.n1096 GNDA.t191 585
R573 GNDA.n1994 GNDA.n1993 585
R574 GNDA.n259 GNDA.n257 585
R575 GNDA.n755 GNDA.n754 585
R576 GNDA.n757 GNDA.n756 585
R577 GNDA.n759 GNDA.n758 585
R578 GNDA.n761 GNDA.n760 585
R579 GNDA.n763 GNDA.n762 585
R580 GNDA.n765 GNDA.n764 585
R581 GNDA.n767 GNDA.n766 585
R582 GNDA.n769 GNDA.n768 585
R583 GNDA.n771 GNDA.n770 585
R584 GNDA.n773 GNDA.n772 585
R585 GNDA.n547 GNDA.n546 585
R586 GNDA.n545 GNDA.n544 585
R587 GNDA.n543 GNDA.n542 585
R588 GNDA.n541 GNDA.n540 585
R589 GNDA.n539 GNDA.n538 585
R590 GNDA.n537 GNDA.n536 585
R591 GNDA.n535 GNDA.n534 585
R592 GNDA.n533 GNDA.n532 585
R593 GNDA.n531 GNDA.n530 585
R594 GNDA.n529 GNDA.n528 585
R595 GNDA.n527 GNDA.n526 585
R596 GNDA.n263 GNDA.n260 585
R597 GNDA.n615 GNDA.n522 585
R598 GNDA.n614 GNDA.n613 585
R599 GNDA.n612 GNDA.n611 585
R600 GNDA.n610 GNDA.n609 585
R601 GNDA.n608 GNDA.n607 585
R602 GNDA.n606 GNDA.n605 585
R603 GNDA.n604 GNDA.n603 585
R604 GNDA.n602 GNDA.n601 585
R605 GNDA.n600 GNDA.n599 585
R606 GNDA.n598 GNDA.n597 585
R607 GNDA.n596 GNDA.n595 585
R608 GNDA.n594 GNDA.n593 585
R609 GNDA.n1490 GNDA.n261 585
R610 GNDA.n1490 GNDA.n469 585
R611 GNDA.n1585 GNDA.n428 585
R612 GNDA.n1572 GNDA.n429 585
R613 GNDA.n1581 GNDA.n1580 585
R614 GNDA.n448 GNDA.n446 585
R615 GNDA.n1497 GNDA.n1496 585
R616 GNDA.n1501 GNDA.n1500 585
R617 GNDA.n1503 GNDA.n1502 585
R618 GNDA.n1510 GNDA.n1509 585
R619 GNDA.n1508 GNDA.n1494 585
R620 GNDA.n1516 GNDA.n1515 585
R621 GNDA.n1518 GNDA.n1517 585
R622 GNDA.n1492 GNDA.n1491 585
R623 GNDA.n1390 GNDA.n495 585
R624 GNDA.n1390 GNDA.n469 585
R625 GNDA.n1486 GNDA.n261 585
R626 GNDA.n1486 GNDA.n469 585
R627 GNDA.n1485 GNDA.n1484 585
R628 GNDA.n1482 GNDA.n1481 585
R629 GNDA.n1480 GNDA.n1479 585
R630 GNDA.n1396 GNDA.n475 585
R631 GNDA.n1398 GNDA.n1397 585
R632 GNDA.n1402 GNDA.n1401 585
R633 GNDA.n1404 GNDA.n1403 585
R634 GNDA.n1411 GNDA.n1410 585
R635 GNDA.n1409 GNDA.n1394 585
R636 GNDA.n1417 GNDA.n1416 585
R637 GNDA.n1419 GNDA.n1418 585
R638 GNDA.n1392 GNDA.n1391 585
R639 GNDA.n1386 GNDA.n495 585
R640 GNDA.n1386 GNDA.n469 585
R641 GNDA.n1385 GNDA.n1384 585
R642 GNDA.n1382 GNDA.n1381 585
R643 GNDA.n1380 GNDA.n1379 585
R644 GNDA.n1296 GNDA.n501 585
R645 GNDA.n1298 GNDA.n1297 585
R646 GNDA.n1302 GNDA.n1301 585
R647 GNDA.n1304 GNDA.n1303 585
R648 GNDA.n1311 GNDA.n1310 585
R649 GNDA.n1309 GNDA.n1294 585
R650 GNDA.n1317 GNDA.n1316 585
R651 GNDA.n1319 GNDA.n1318 585
R652 GNDA.n1292 GNDA.n1291 585
R653 GNDA.n1690 GNDA.n1689 585
R654 GNDA.n1692 GNDA.n1623 585
R655 GNDA.n1694 GNDA.n1693 585
R656 GNDA.n1695 GNDA.n1622 585
R657 GNDA.n1697 GNDA.n1696 585
R658 GNDA.n1699 GNDA.n1620 585
R659 GNDA.n1701 GNDA.n1700 585
R660 GNDA.n1702 GNDA.n1619 585
R661 GNDA.n1704 GNDA.n1703 585
R662 GNDA.n1706 GNDA.n1617 585
R663 GNDA.n1708 GNDA.n1707 585
R664 GNDA.n1709 GNDA.n1616 585
R665 GNDA.n1962 GNDA.n1961 585
R666 GNDA.n1634 GNDA.n298 585
R667 GNDA.n1636 GNDA.n1635 585
R668 GNDA.n1638 GNDA.n1632 585
R669 GNDA.n1640 GNDA.n1639 585
R670 GNDA.n1641 GNDA.n1631 585
R671 GNDA.n1643 GNDA.n1642 585
R672 GNDA.n1645 GNDA.n1629 585
R673 GNDA.n1647 GNDA.n1646 585
R674 GNDA.n1648 GNDA.n1628 585
R675 GNDA.n1650 GNDA.n1649 585
R676 GNDA.n1652 GNDA.n1626 585
R677 GNDA.n202 GNDA.n201 585
R678 GNDA.n1798 GNDA.n1797 585
R679 GNDA.n1800 GNDA.n1799 585
R680 GNDA.n1802 GNDA.n1794 585
R681 GNDA.n1804 GNDA.n1803 585
R682 GNDA.n1805 GNDA.n1793 585
R683 GNDA.n1807 GNDA.n1806 585
R684 GNDA.n1809 GNDA.n1791 585
R685 GNDA.n1811 GNDA.n1810 585
R686 GNDA.n1812 GNDA.n1790 585
R687 GNDA.n1814 GNDA.n1813 585
R688 GNDA.n1816 GNDA.n296 585
R689 GNDA.n291 GNDA.n290 585
R690 GNDA.n1966 GNDA.n291 585
R691 GNDA.n912 GNDA.n911 585
R692 GNDA.n909 GNDA.n753 585
R693 GNDA.n800 GNDA.n799 585
R694 GNDA.n904 GNDA.n903 585
R695 GNDA.n902 GNDA.n901 585
R696 GNDA.n828 GNDA.n804 585
R697 GNDA.n830 GNDA.n829 585
R698 GNDA.n835 GNDA.n834 585
R699 GNDA.n833 GNDA.n826 585
R700 GNDA.n841 GNDA.n840 585
R701 GNDA.n843 GNDA.n842 585
R702 GNDA.n824 GNDA.n823 585
R703 GNDA.n1964 GNDA.n292 585
R704 GNDA.n1966 GNDA.n292 585
R705 GNDA.n1967 GNDA.n290 585
R706 GNDA.n1967 GNDA.n1966 585
R707 GNDA.n633 GNDA.n289 585
R708 GNDA.n746 GNDA.n745 585
R709 GNDA.n635 GNDA.n632 585
R710 GNDA.n740 GNDA.n739 585
R711 GNDA.n738 GNDA.n737 585
R712 GNDA.n663 GNDA.n639 585
R713 GNDA.n665 GNDA.n664 585
R714 GNDA.n670 GNDA.n669 585
R715 GNDA.n668 GNDA.n661 585
R716 GNDA.n676 GNDA.n675 585
R717 GNDA.n678 GNDA.n677 585
R718 GNDA.n659 GNDA.n658 585
R719 GNDA.n1965 GNDA.n1964 585
R720 GNDA.n1966 GNDA.n1965 585
R721 GNDA.n991 GNDA.n294 585
R722 GNDA.n992 GNDA.n928 585
R723 GNDA.n1002 GNDA.n1001 585
R724 GNDA.n1004 GNDA.n926 585
R725 GNDA.n1007 GNDA.n1006 585
R726 GNDA.n1008 GNDA.n922 585
R727 GNDA.n1017 GNDA.n1016 585
R728 GNDA.n1019 GNDA.n921 585
R729 GNDA.n1022 GNDA.n1021 585
R730 GNDA.n1023 GNDA.n915 585
R731 GNDA.n1032 GNDA.n1031 585
R732 GNDA.n1034 GNDA.n624 585
R733 GNDA.n1711 GNDA.n1710 585
R734 GNDA.n1713 GNDA.n1615 585
R735 GNDA.n1716 GNDA.n1715 585
R736 GNDA.n1717 GNDA.n1614 585
R737 GNDA.n1719 GNDA.n1718 585
R738 GNDA.n1721 GNDA.n1613 585
R739 GNDA.n1724 GNDA.n1723 585
R740 GNDA.n1725 GNDA.n1612 585
R741 GNDA.n1727 GNDA.n1726 585
R742 GNDA.n1729 GNDA.n1611 585
R743 GNDA.n1730 GNDA.n411 585
R744 GNDA.n1610 GNDA.n410 585
R745 GNDA.n775 GNDA.n774 585
R746 GNDA.n777 GNDA.n776 585
R747 GNDA.n779 GNDA.n778 585
R748 GNDA.n781 GNDA.n780 585
R749 GNDA.n783 GNDA.n782 585
R750 GNDA.n785 GNDA.n784 585
R751 GNDA.n787 GNDA.n786 585
R752 GNDA.n789 GNDA.n788 585
R753 GNDA.n791 GNDA.n790 585
R754 GNDA.n793 GNDA.n792 585
R755 GNDA.n795 GNDA.n794 585
R756 GNDA.n1610 GNDA.n423 585
R757 GNDA.n1608 GNDA.n1607 585
R758 GNDA.n1606 GNDA.n425 585
R759 GNDA.n1605 GNDA.n424 585
R760 GNDA.n1610 GNDA.n424 585
R761 GNDA.n1604 GNDA.n1603 585
R762 GNDA.n1602 GNDA.n1601 585
R763 GNDA.n1600 GNDA.n1599 585
R764 GNDA.n1598 GNDA.n1597 585
R765 GNDA.n1596 GNDA.n1595 585
R766 GNDA.n1594 GNDA.n1593 585
R767 GNDA.n1592 GNDA.n1591 585
R768 GNDA.n1590 GNDA.n1589 585
R769 GNDA.n1588 GNDA.n1587 585
R770 GNDA.n1587 GNDA.n1586 585
R771 GNDA.n2221 GNDA.n2220 585
R772 GNDA.n2250 GNDA.n2219 585
R773 GNDA.n2254 GNDA.n2219 585
R774 GNDA.n2249 GNDA.n2248 585
R775 GNDA.n2247 GNDA.n2246 585
R776 GNDA.n2245 GNDA.n2244 585
R777 GNDA.n2243 GNDA.n2242 585
R778 GNDA.n2241 GNDA.n2240 585
R779 GNDA.n2239 GNDA.n2238 585
R780 GNDA.n2237 GNDA.n2236 585
R781 GNDA.n2235 GNDA.n2234 585
R782 GNDA.n2233 GNDA.n2232 585
R783 GNDA.n2231 GNDA.n2196 585
R784 GNDA.n2256 GNDA.n2255 585
R785 GNDA.n2255 GNDA.n2254 585
R786 GNDA.n63 GNDA.n59 585
R787 GNDA.n61 GNDA.n58 585
R788 GNDA.n66 GNDA.n58 585
R789 GNDA.n2639 GNDA.n5 585
R790 GNDA.n2644 GNDA.n2643 585
R791 GNDA.n2643 GNDA.n2642 585
R792 GNDA.n2345 GNDA.n2344 585
R793 GNDA.n2350 GNDA.n2343 585
R794 GNDA.n2343 GNDA.n2172 585
R795 GNDA.n2352 GNDA.n2351 585
R796 GNDA.n2311 GNDA.n2310 585
R797 GNDA.n2316 GNDA.n2309 585
R798 GNDA.n2309 GNDA.n6 585
R799 GNDA.n2318 GNDA.n2317 585
R800 GNDA.n2185 GNDA.n2184 585
R801 GNDA.n2286 GNDA.n2183 585
R802 GNDA.n2290 GNDA.n2183 585
R803 GNDA.n2285 GNDA.n2284 585
R804 GNDA.n2283 GNDA.n2282 585
R805 GNDA.n2281 GNDA.n2280 585
R806 GNDA.n2279 GNDA.n2278 585
R807 GNDA.n2277 GNDA.n2276 585
R808 GNDA.n2275 GNDA.n2274 585
R809 GNDA.n2273 GNDA.n2272 585
R810 GNDA.n2271 GNDA.n2270 585
R811 GNDA.n2269 GNDA.n2268 585
R812 GNDA.n2267 GNDA.n2266 585
R813 GNDA.n2264 GNDA.n2182 585
R814 GNDA.n2290 GNDA.n2182 585
R815 GNDA.n2537 GNDA.n2536 585
R816 GNDA.n2534 GNDA.n2533 585
R817 GNDA.n2533 GNDA.n2503 585
R818 GNDA.n2542 GNDA.n2541 585
R819 GNDA.n2544 GNDA.n2532 585
R820 GNDA.n2547 GNDA.n2546 585
R821 GNDA.n2530 GNDA.n2529 585
R822 GNDA.n2552 GNDA.n2551 585
R823 GNDA.n2554 GNDA.n2528 585
R824 GNDA.n2557 GNDA.n2556 585
R825 GNDA.n2526 GNDA.n2525 585
R826 GNDA.n2562 GNDA.n2561 585
R827 GNDA.n2564 GNDA.n2524 585
R828 GNDA.n2566 GNDA.n2565 585
R829 GNDA.n2565 GNDA.n2503 585
R830 GNDA.n2513 GNDA.n2512 585
R831 GNDA.n2596 GNDA.n2511 585
R832 GNDA.n2600 GNDA.n2511 585
R833 GNDA.n2595 GNDA.n2594 585
R834 GNDA.n2593 GNDA.n2592 585
R835 GNDA.n2591 GNDA.n2590 585
R836 GNDA.n2589 GNDA.n2588 585
R837 GNDA.n2587 GNDA.n2586 585
R838 GNDA.n2585 GNDA.n2584 585
R839 GNDA.n2583 GNDA.n2582 585
R840 GNDA.n2581 GNDA.n2580 585
R841 GNDA.n2579 GNDA.n2578 585
R842 GNDA.n2577 GNDA.n2576 585
R843 GNDA.n2574 GNDA.n2510 585
R844 GNDA.n2600 GNDA.n2510 585
R845 GNDA.n2201 GNDA.n2200 585
R846 GNDA.n2209 GNDA.n2199 585
R847 GNDA.n2213 GNDA.n2199 585
R848 GNDA.n2208 GNDA.n2207 585
R849 GNDA.n2206 GNDA.n2205 585
R850 GNDA.n2203 GNDA.n2198 585
R851 GNDA.n2213 GNDA.n2198 585
R852 GNDA.n2379 GNDA.n2373 585
R853 GNDA.n2377 GNDA.n2376 585
R854 GNDA.n2375 GNDA.n2371 585
R855 GNDA.n2390 GNDA.n2389 585
R856 GNDA.n2389 GNDA.n2388 585
R857 GNDA.n2456 GNDA.n2446 585
R858 GNDA.n2454 GNDA.n2453 585
R859 GNDA.n2452 GNDA.n2451 585
R860 GNDA.n2449 GNDA.n2444 585
R861 GNDA.n2459 GNDA.n2444 585
R862 GNDA.n2293 GNDA.n2292 585
R863 GNDA.n2298 GNDA.n2291 585
R864 GNDA.n2302 GNDA.n2291 585
R865 GNDA.n2297 GNDA.n2296 585
R866 GNDA.n2295 GNDA.n2175 585
R867 GNDA.n2304 GNDA.n2303 585
R868 GNDA.n2303 GNDA.n2302 585
R869 GNDA.n2603 GNDA.n2602 585
R870 GNDA.n2608 GNDA.n2601 585
R871 GNDA.n2612 GNDA.n2601 585
R872 GNDA.n2607 GNDA.n2606 585
R873 GNDA.n2605 GNDA.n30 585
R874 GNDA.n2614 GNDA.n2613 585
R875 GNDA.n2613 GNDA.n2612 585
R876 GNDA.n15 GNDA.n14 585
R877 GNDA.n2624 GNDA.n13 585
R878 GNDA.n2628 GNDA.n13 585
R879 GNDA.n2623 GNDA.n2622 585
R880 GNDA.n2621 GNDA.n2620 585
R881 GNDA.n2618 GNDA.n12 585
R882 GNDA.n2628 GNDA.n12 585
R883 GNDA.n2363 GNDA.n2362 585
R884 GNDA.n2401 GNDA.n2400 585
R885 GNDA.n2386 GNDA.n2385 585
R886 GNDA.n2461 GNDA.n56 585
R887 GNDA.n2488 GNDA.n2487 585
R888 GNDA.n2500 GNDA.n2499 585
R889 GNDA.n2361 GNDA.n89 585
R890 GNDA.n2415 GNDA.n89 585
R891 GNDA.n2397 GNDA.n2396 585
R892 GNDA.n2396 GNDA.n67 585
R893 GNDA.n2384 GNDA.n69 585
R894 GNDA.n2442 GNDA.n69 585
R895 GNDA.n2463 GNDA.n2462 585
R896 GNDA.n2462 GNDA.n34 585
R897 GNDA.n2486 GNDA.n2484 585
R898 GNDA.n2484 GNDA.n2483 585
R899 GNDA.n2496 GNDA.n2495 585
R900 GNDA.n2495 GNDA.n10 585
R901 GNDA.n2412 GNDA.n87 585
R902 GNDA.n2417 GNDA.n2416 585
R903 GNDA.n2416 GNDA.n2415 585
R904 GNDA.n2425 GNDA.n2421 585
R905 GNDA.n2427 GNDA.n2426 585
R906 GNDA.n2426 GNDA.n67 585
R907 GNDA.n2439 GNDA.n71 585
R908 GNDA.n2437 GNDA.n70 585
R909 GNDA.n2442 GNDA.n70 585
R910 GNDA.n2436 GNDA.n2435 585
R911 GNDA.n2480 GNDA.n37 585
R912 GNDA.n2478 GNDA.n36 585
R913 GNDA.n2483 GNDA.n36 585
R914 GNDA.n2472 GNDA.n2468 585
R915 GNDA.n2474 GNDA.n2473 585
R916 GNDA.n2473 GNDA.n10 585
R917 GNDA.n44 GNDA.n43 585
R918 GNDA.n49 GNDA.n42 585
R919 GNDA.n42 GNDA.n34 585
R920 GNDA.n51 GNDA.n50 585
R921 GNDA.n2126 GNDA.n135 585
R922 GNDA.n2129 GNDA.n2128 585
R923 GNDA.n2130 GNDA.n2129 585
R924 GNDA.n2121 GNDA.n2120 585
R925 GNDA.n1928 GNDA.n318 585
R926 GNDA.n1929 GNDA.n1928 585
R927 GNDA.n1735 GNDA.n1734 585
R928 GNDA.n1736 GNDA.n1735 585
R929 GNDA.n1740 GNDA.n1739 585
R930 GNDA.n1739 GNDA.n1738 585
R931 GNDA.n339 GNDA.n338 585
R932 GNDA.n1737 GNDA.n338 585
R933 GNDA.n1748 GNDA.n1747 585
R934 GNDA.n1749 GNDA.n1748 585
R935 GNDA.n337 GNDA.n336 585
R936 GNDA.n1750 GNDA.n337 585
R937 GNDA.n1753 GNDA.n1752 585
R938 GNDA.n1752 GNDA.n1751 585
R939 GNDA.n333 GNDA.n328 585
R940 GNDA.n328 GNDA.n327 585
R941 GNDA.n1763 GNDA.n1762 585
R942 GNDA.n1764 GNDA.n1763 585
R943 GNDA.n330 GNDA.n325 585
R944 GNDA.n1765 GNDA.n325 585
R945 GNDA.n1767 GNDA.n326 585
R946 GNDA.n1767 GNDA.n1766 585
R947 GNDA.n1771 GNDA.n1770 585
R948 GNDA.n1770 GNDA.n1769 585
R949 GNDA.n1773 GNDA.n317 585
R950 GNDA.n1768 GNDA.n317 585
R951 GNDA.n1845 GNDA.n1778 585
R952 GNDA.n1847 GNDA.n1845 585
R953 GNDA.n1920 GNDA.n318 585
R954 GNDA.n1920 GNDA.n308 585
R955 GNDA.n1919 GNDA.n1917 585
R956 GNDA.n1919 GNDA.n1918 585
R957 GNDA.n126 GNDA.n124 585
R958 GNDA.n2137 GNDA.n126 585
R959 GNDA.n2152 GNDA.n2151 585
R960 GNDA.n2151 GNDA.n2150 585
R961 GNDA.n2139 GNDA.n127 585
R962 GNDA.n2149 GNDA.n127 585
R963 GNDA.n2147 GNDA.n2146 585
R964 GNDA.n2148 GNDA.n2147 585
R965 GNDA.n2142 GNDA.n101 585
R966 GNDA.n2138 GNDA.n101 585
R967 GNDA.n2160 GNDA.n2159 585
R968 GNDA.n2161 GNDA.n2160 585
R969 GNDA.n103 GNDA.n102 585
R970 GNDA.n1850 GNDA.n102 585
R971 GNDA.n1855 GNDA.n1854 585
R972 GNDA.n1856 GNDA.n1855 585
R973 GNDA.n1777 GNDA.n1776 585
R974 GNDA.n1857 GNDA.n1777 585
R975 GNDA.n1860 GNDA.n1859 585
R976 GNDA.n1859 GNDA.n1858 585
R977 GNDA.n1849 GNDA.n1846 585
R978 GNDA.n1849 GNDA.n1848 585
R979 GNDA.n1778 GNDA.n172 585
R980 GNDA.n1938 GNDA.n172 585
R981 GNDA.n2093 GNDA.n2092 585
R982 GNDA.n2094 GNDA.n2093 585
R983 GNDA.n165 GNDA.n163 585
R984 GNDA.n2095 GNDA.n165 585
R985 GNDA.n2110 GNDA.n2109 585
R986 GNDA.n2109 GNDA.n2108 585
R987 GNDA.n2097 GNDA.n166 585
R988 GNDA.n2107 GNDA.n166 585
R989 GNDA.n2105 GNDA.n2104 585
R990 GNDA.n2106 GNDA.n2105 585
R991 GNDA.n2100 GNDA.n140 585
R992 GNDA.n2096 GNDA.n140 585
R993 GNDA.n2118 GNDA.n2117 585
R994 GNDA.n2119 GNDA.n2118 585
R995 GNDA.n142 GNDA.n141 585
R996 GNDA.n178 GNDA.n141 585
R997 GNDA.n183 GNDA.n182 585
R998 GNDA.n184 GNDA.n183 585
R999 GNDA.n176 GNDA.n175 585
R1000 GNDA.n185 GNDA.n176 585
R1001 GNDA.n2035 GNDA.n2034 585
R1002 GNDA.n2034 GNDA.n2033 585
R1003 GNDA.n190 GNDA.n177 585
R1004 GNDA.n2032 GNDA.n177 585
R1005 GNDA.n222 GNDA.n129 585
R1006 GNDA.n223 GNDA.n222 585
R1007 GNDA.n221 GNDA.n220 585
R1008 GNDA.n219 GNDA.n212 585
R1009 GNDA.n214 GNDA.n213 585
R1010 GNDA.t191 GNDA.n236 512.884
R1011 GNDA.t191 GNDA.n228 512.884
R1012 GNDA.n2257 GNDA.t259 505.467
R1013 GNDA.n2573 GNDA.t204 505.467
R1014 GNDA.n2567 GNDA.t227 505.467
R1015 GNDA.n2263 GNDA.t241 505.467
R1016 GNDA.n2366 GNDA.t209 499.442
R1017 GNDA.n2493 GNDA.t279 499.442
R1018 GNDA.n2418 GNDA.t214 499.442
R1019 GNDA.n2428 GNDA.t233 499.442
R1020 GNDA.n2477 GNDA.t275 499.442
R1021 GNDA.n2475 GNDA.t193 499.442
R1022 GNDA.n1 GNDA.t257 499.442
R1023 GNDA.n2645 GNDA.t267 499.442
R1024 GNDA.n73 GNDA.t235 489.401
R1025 GNDA.n2464 GNDA.t277 489.401
R1026 GNDA.n171 GNDA.t147 433.382
R1027 GNDA.n2442 GNDA.n67 431.902
R1028 GNDA.n2483 GNDA.n34 431.902
R1029 GNDA.n310 GNDA.t244 409.067
R1030 GNDA.n1932 GNDA.t250 409.067
R1031 GNDA.n1955 GNDA.t272 409.067
R1032 GNDA.n1944 GNDA.t224 409.067
R1033 GNDA.n1941 GNDA.t247 409.067
R1034 GNDA.n2029 GNDA.t230 409.067
R1035 GNDA.t191 GNDA.n237 391.411
R1036 GNDA.t191 GNDA.n229 391.411
R1037 GNDA.n2290 GNDA.n90 368.587
R1038 GNDA.n2503 GNDA.n2502 368.587
R1039 GNDA.n2415 GNDA.t210 364.418
R1040 GNDA.t218 GNDA.n67 364.418
R1041 GNDA.t115 GNDA.n2442 364.418
R1042 GNDA.t133 GNDA.n34 364.418
R1043 GNDA.n2483 GNDA.t270 364.418
R1044 GNDA.t194 GNDA.n10 364.418
R1045 GNDA.t191 GNDA.n204 172.876
R1046 GNDA.n1958 GNDA.t191 172.876
R1047 GNDA.n307 GNDA.t191 172.615
R1048 GNDA.t191 GNDA.n137 172.615
R1049 GNDA.n95 GNDA.n9 309.122
R1050 GNDA.t10 GNDA.t218 296.933
R1051 GNDA.t93 GNDA.t64 296.933
R1052 GNDA.t191 GNDA.t92 294.625
R1053 GNDA.n2252 GNDA.n2251 267.125
R1054 GNDA.n2230 GNDA.n2195 267.125
R1055 GNDA.n2300 GNDA.n2299 267.125
R1056 GNDA.n2294 GNDA.n2174 267.125
R1057 GNDA.n2211 GNDA.n2210 267.125
R1058 GNDA.n2204 GNDA.n2202 267.125
R1059 GNDA.n2610 GNDA.n2609 267.125
R1060 GNDA.n2604 GNDA.n29 267.125
R1061 GNDA.n2626 GNDA.n2625 267.125
R1062 GNDA.n2619 GNDA.n16 267.125
R1063 GNDA.n2598 GNDA.n2597 267.125
R1064 GNDA.n2575 GNDA.n2522 267.125
R1065 GNDA.n2539 GNDA.n2538 267.125
R1066 GNDA.n2560 GNDA.n2523 267.125
R1067 GNDA.n2288 GNDA.n2287 267.125
R1068 GNDA.n2265 GNDA.n2194 267.125
R1069 GNDA.n1610 GNDA.n416 264.301
R1070 GNDA.n2020 GNDA.n191 264.301
R1071 GNDA.n1037 GNDA.n1036 264.301
R1072 GNDA.n1289 GNDA.n520 264.301
R1073 GNDA.n1733 GNDA.n1732 264.301
R1074 GNDA.n797 GNDA.n796 264.301
R1075 GNDA.n1173 GNDA.n1143 259.416
R1076 GNDA.n1994 GNDA.n258 259.416
R1077 GNDA.n1690 GNDA.n1625 259.416
R1078 GNDA.n1961 GNDA.n1960 259.416
R1079 GNDA.n548 GNDA.n547 259.416
R1080 GNDA.n1201 GNDA.n1082 259.416
R1081 GNDA.n1057 GNDA.n522 259.416
R1082 GNDA.n1998 GNDA.n202 259.416
R1083 GNDA.n1263 GNDA.n1068 259.416
R1084 GNDA.n1557 GNDA.n1556 258.334
R1085 GNDA.n880 GNDA.n821 258.334
R1086 GNDA.n392 GNDA.n390 258.334
R1087 GNDA.n1899 GNDA.n1898 258.334
R1088 GNDA.n715 GNDA.n656 258.334
R1089 GNDA.n1458 GNDA.n1457 258.334
R1090 GNDA.n976 GNDA.n934 258.334
R1091 GNDA.n2074 GNDA.n2073 258.334
R1092 GNDA.n1358 GNDA.n1357 258.334
R1093 GNDA.n569 GNDA.n205 254.34
R1094 GNDA.n566 GNDA.n205 254.34
R1095 GNDA.n562 GNDA.n205 254.34
R1096 GNDA.n559 GNDA.n205 254.34
R1097 GNDA.n554 GNDA.n205 254.34
R1098 GNDA.n549 GNDA.n205 254.34
R1099 GNDA.n525 GNDA.n239 254.34
R1100 GNDA.n552 GNDA.n239 254.34
R1101 GNDA.n582 GNDA.n239 254.34
R1102 GNDA.n576 GNDA.n239 254.34
R1103 GNDA.n574 GNDA.n239 254.34
R1104 GNDA.n1958 GNDA.n305 254.34
R1105 GNDA.n1958 GNDA.n304 254.34
R1106 GNDA.n1958 GNDA.n303 254.34
R1107 GNDA.n1958 GNDA.n302 254.34
R1108 GNDA.n1958 GNDA.n301 254.34
R1109 GNDA.n1959 GNDA.n1958 254.34
R1110 GNDA.n1818 GNDA.n137 254.34
R1111 GNDA.n1820 GNDA.n137 254.34
R1112 GNDA.n1828 GNDA.n137 254.34
R1113 GNDA.n1830 GNDA.n137 254.34
R1114 GNDA.n1838 GNDA.n137 254.34
R1115 GNDA.n1841 GNDA.n137 254.34
R1116 GNDA.n1926 GNDA.n204 254.34
R1117 GNDA.n1667 GNDA.n204 254.34
R1118 GNDA.n1665 GNDA.n204 254.34
R1119 GNDA.n1662 GNDA.n204 254.34
R1120 GNDA.n1657 GNDA.n204 254.34
R1121 GNDA.n1654 GNDA.n204 254.34
R1122 GNDA.n1685 GNDA.n307 254.34
R1123 GNDA.n1653 GNDA.n307 254.34
R1124 GNDA.n1678 GNDA.n307 254.34
R1125 GNDA.n1672 GNDA.n307 254.34
R1126 GNDA.n1670 GNDA.n307 254.34
R1127 GNDA.n1922 GNDA.n307 254.34
R1128 GNDA.n286 GNDA.n285 254.34
R1129 GNDA.n285 GNDA.n284 254.34
R1130 GNDA.n285 GNDA.n283 254.34
R1131 GNDA.n285 GNDA.n282 254.34
R1132 GNDA.n285 GNDA.n281 254.34
R1133 GNDA.n285 GNDA.n280 254.34
R1134 GNDA.n1989 GNDA.n1988 254.34
R1135 GNDA.n1988 GNDA.n1987 254.34
R1136 GNDA.n1988 GNDA.n268 254.34
R1137 GNDA.n1988 GNDA.n267 254.34
R1138 GNDA.n1988 GNDA.n266 254.34
R1139 GNDA.n1988 GNDA.n265 254.34
R1140 GNDA.n1996 GNDA.n1995 254.34
R1141 GNDA.n1996 GNDA.n256 254.34
R1142 GNDA.n1996 GNDA.n255 254.34
R1143 GNDA.n1996 GNDA.n254 254.34
R1144 GNDA.n1996 GNDA.n253 254.34
R1145 GNDA.n1996 GNDA.n252 254.34
R1146 GNDA.n1996 GNDA.n251 254.34
R1147 GNDA.n1996 GNDA.n250 254.34
R1148 GNDA.n1996 GNDA.n249 254.34
R1149 GNDA.n1996 GNDA.n248 254.34
R1150 GNDA.n1996 GNDA.n247 254.34
R1151 GNDA.n1996 GNDA.n246 254.34
R1152 GNDA.n1996 GNDA.n245 254.34
R1153 GNDA.n1996 GNDA.n244 254.34
R1154 GNDA.n1996 GNDA.n243 254.34
R1155 GNDA.n1996 GNDA.n242 254.34
R1156 GNDA.n1996 GNDA.n241 254.34
R1157 GNDA.n1996 GNDA.n240 254.34
R1158 GNDA.n1584 GNDA.n1583 254.34
R1159 GNDA.n1583 GNDA.n1582 254.34
R1160 GNDA.n1583 GNDA.n445 254.34
R1161 GNDA.n1583 GNDA.n444 254.34
R1162 GNDA.n1583 GNDA.n443 254.34
R1163 GNDA.n1583 GNDA.n442 254.34
R1164 GNDA.n1583 GNDA.n441 254.34
R1165 GNDA.n1583 GNDA.n440 254.34
R1166 GNDA.n1583 GNDA.n439 254.34
R1167 GNDA.n1583 GNDA.n438 254.34
R1168 GNDA.n1583 GNDA.n437 254.34
R1169 GNDA.n1583 GNDA.n436 254.34
R1170 GNDA.n1583 GNDA.n435 254.34
R1171 GNDA.n1583 GNDA.n434 254.34
R1172 GNDA.n1583 GNDA.n433 254.34
R1173 GNDA.n1583 GNDA.n432 254.34
R1174 GNDA.n1583 GNDA.n431 254.34
R1175 GNDA.n1583 GNDA.n430 254.34
R1176 GNDA.n1691 GNDA.n224 254.34
R1177 GNDA.n1624 GNDA.n224 254.34
R1178 GNDA.n1698 GNDA.n224 254.34
R1179 GNDA.n1621 GNDA.n224 254.34
R1180 GNDA.n1705 GNDA.n224 254.34
R1181 GNDA.n1618 GNDA.n224 254.34
R1182 GNDA.n299 GNDA.n224 254.34
R1183 GNDA.n1637 GNDA.n224 254.34
R1184 GNDA.n1633 GNDA.n224 254.34
R1185 GNDA.n1644 GNDA.n224 254.34
R1186 GNDA.n1630 GNDA.n224 254.34
R1187 GNDA.n1651 GNDA.n224 254.34
R1188 GNDA.n1796 GNDA.n224 254.34
R1189 GNDA.n1801 GNDA.n224 254.34
R1190 GNDA.n1795 GNDA.n224 254.34
R1191 GNDA.n1808 GNDA.n224 254.34
R1192 GNDA.n1792 GNDA.n224 254.34
R1193 GNDA.n1815 GNDA.n224 254.34
R1194 GNDA.n914 GNDA.n913 254.34
R1195 GNDA.n914 GNDA.n752 254.34
R1196 GNDA.n914 GNDA.n751 254.34
R1197 GNDA.n914 GNDA.n750 254.34
R1198 GNDA.n914 GNDA.n749 254.34
R1199 GNDA.n914 GNDA.n748 254.34
R1200 GNDA.n914 GNDA.n747 254.34
R1201 GNDA.n914 GNDA.n631 254.34
R1202 GNDA.n914 GNDA.n630 254.34
R1203 GNDA.n914 GNDA.n629 254.34
R1204 GNDA.n914 GNDA.n628 254.34
R1205 GNDA.n914 GNDA.n627 254.34
R1206 GNDA.n927 GNDA.n914 254.34
R1207 GNDA.n1003 GNDA.n914 254.34
R1208 GNDA.n1005 GNDA.n914 254.34
R1209 GNDA.n1018 GNDA.n914 254.34
R1210 GNDA.n1020 GNDA.n914 254.34
R1211 GNDA.n1033 GNDA.n914 254.34
R1212 GNDA.n1712 GNDA.n1610 254.34
R1213 GNDA.n1714 GNDA.n1610 254.34
R1214 GNDA.n1720 GNDA.n1610 254.34
R1215 GNDA.n1722 GNDA.n1610 254.34
R1216 GNDA.n1728 GNDA.n1610 254.34
R1217 GNDA.n1731 GNDA.n1610 254.34
R1218 GNDA.n1610 GNDA.n417 254.34
R1219 GNDA.n1610 GNDA.n418 254.34
R1220 GNDA.n1610 GNDA.n419 254.34
R1221 GNDA.n1610 GNDA.n420 254.34
R1222 GNDA.n1610 GNDA.n421 254.34
R1223 GNDA.n1610 GNDA.n422 254.34
R1224 GNDA.n1610 GNDA.n1609 254.34
R1225 GNDA.n1610 GNDA.n412 254.34
R1226 GNDA.n1610 GNDA.n413 254.34
R1227 GNDA.n1610 GNDA.n414 254.34
R1228 GNDA.n1610 GNDA.n415 254.34
R1229 GNDA.n1094 GNDA.t191 250.349
R1230 GNDA.n1608 GNDA.n426 249.663
R1231 GNDA.n774 GNDA.n773 249.663
R1232 GNDA.n1711 GNDA.n1616 249.663
R1233 GNDA.n1686 GNDA.n1652 249.663
R1234 GNDA.n1990 GNDA.n263 249.663
R1235 GNDA.n1177 GNDA.n1103 249.663
R1236 GNDA.n593 GNDA.n592 249.663
R1237 GNDA.n1817 GNDA.n1816 249.663
R1238 GNDA.n1238 GNDA.n1080 249.663
R1239 GNDA.n2129 GNDA.n135 246.25
R1240 GNDA.n2129 GNDA.n2120 246.25
R1241 GNDA.n44 GNDA.n42 246.25
R1242 GNDA.n51 GNDA.n42 246.25
R1243 GNDA.n2473 GNDA.n2472 246.25
R1244 GNDA.n37 GNDA.n36 246.25
R1245 GNDA.n71 GNDA.n70 246.25
R1246 GNDA.n2435 GNDA.n70 246.25
R1247 GNDA.n2426 GNDA.n2425 246.25
R1248 GNDA.n2416 GNDA.n87 246.25
R1249 GNDA.n2500 GNDA.n2495 246.25
R1250 GNDA.n2488 GNDA.n2484 246.25
R1251 GNDA.n2462 GNDA.n2461 246.25
R1252 GNDA.n2386 GNDA.n69 246.25
R1253 GNDA.n2401 GNDA.n2396 246.25
R1254 GNDA.n2363 GNDA.n89 246.25
R1255 GNDA.n14 GNDA.n13 246.25
R1256 GNDA.n2622 GNDA.n13 246.25
R1257 GNDA.n2620 GNDA.n12 246.25
R1258 GNDA.n2602 GNDA.n2601 246.25
R1259 GNDA.n2606 GNDA.n2601 246.25
R1260 GNDA.n2613 GNDA.n30 246.25
R1261 GNDA.n2292 GNDA.n2291 246.25
R1262 GNDA.n2296 GNDA.n2291 246.25
R1263 GNDA.n2303 GNDA.n2175 246.25
R1264 GNDA.n2453 GNDA.n2446 246.25
R1265 GNDA.n2451 GNDA.n2444 246.25
R1266 GNDA.n2376 GNDA.n2373 246.25
R1267 GNDA.n2389 GNDA.n2371 246.25
R1268 GNDA.n2200 GNDA.n2199 246.25
R1269 GNDA.n2207 GNDA.n2199 246.25
R1270 GNDA.n2205 GNDA.n2198 246.25
R1271 GNDA.n2512 GNDA.n2511 246.25
R1272 GNDA.n2594 GNDA.n2511 246.25
R1273 GNDA.n2592 GNDA.n2591 246.25
R1274 GNDA.n2588 GNDA.n2587 246.25
R1275 GNDA.n2584 GNDA.n2583 246.25
R1276 GNDA.n2580 GNDA.n2579 246.25
R1277 GNDA.n2576 GNDA.n2510 246.25
R1278 GNDA.n2536 GNDA.n2533 246.25
R1279 GNDA.n2542 GNDA.n2533 246.25
R1280 GNDA.n2546 GNDA.n2544 246.25
R1281 GNDA.n2552 GNDA.n2529 246.25
R1282 GNDA.n2556 GNDA.n2554 246.25
R1283 GNDA.n2562 GNDA.n2525 246.25
R1284 GNDA.n2565 GNDA.n2564 246.25
R1285 GNDA.n2184 GNDA.n2183 246.25
R1286 GNDA.n2284 GNDA.n2183 246.25
R1287 GNDA.n2282 GNDA.n2281 246.25
R1288 GNDA.n2278 GNDA.n2277 246.25
R1289 GNDA.n2274 GNDA.n2273 246.25
R1290 GNDA.n2270 GNDA.n2269 246.25
R1291 GNDA.n2266 GNDA.n2182 246.25
R1292 GNDA.n2311 GNDA.n2309 246.25
R1293 GNDA.n2318 GNDA.n2309 246.25
R1294 GNDA.n2345 GNDA.n2343 246.25
R1295 GNDA.n2352 GNDA.n2343 246.25
R1296 GNDA.n2643 GNDA.n5 246.25
R1297 GNDA.n59 GNDA.n58 246.25
R1298 GNDA.n2220 GNDA.n2219 246.25
R1299 GNDA.n2248 GNDA.n2219 246.25
R1300 GNDA.n2246 GNDA.n2245 246.25
R1301 GNDA.n2242 GNDA.n2241 246.25
R1302 GNDA.n2238 GNDA.n2237 246.25
R1303 GNDA.n2234 GNDA.n2233 246.25
R1304 GNDA.n2255 GNDA.n2196 246.25
R1305 GNDA.n222 GNDA.n221 246.25
R1306 GNDA.n213 GNDA.n212 246.25
R1307 GNDA.n2025 GNDA.n2024 241.643
R1308 GNDA.n2254 GNDA.n2253 241.643
R1309 GNDA.n2254 GNDA.n2214 241.643
R1310 GNDA.n2254 GNDA.n2215 241.643
R1311 GNDA.n2254 GNDA.n2216 241.643
R1312 GNDA.n2254 GNDA.n2217 241.643
R1313 GNDA.n2254 GNDA.n2218 241.643
R1314 GNDA.n66 GNDA.n65 241.643
R1315 GNDA.n2642 GNDA.n2641 241.643
R1316 GNDA.n2346 GNDA.n2172 241.643
R1317 GNDA.n2353 GNDA.n2172 241.643
R1318 GNDA.n2312 GNDA.n6 241.643
R1319 GNDA.n2319 GNDA.n6 241.643
R1320 GNDA.n2290 GNDA.n2289 241.643
R1321 GNDA.n2290 GNDA.n2177 241.643
R1322 GNDA.n2290 GNDA.n2178 241.643
R1323 GNDA.n2290 GNDA.n2179 241.643
R1324 GNDA.n2290 GNDA.n2180 241.643
R1325 GNDA.n2290 GNDA.n2181 241.643
R1326 GNDA.n2535 GNDA.n2503 241.643
R1327 GNDA.n2543 GNDA.n2503 241.643
R1328 GNDA.n2545 GNDA.n2503 241.643
R1329 GNDA.n2553 GNDA.n2503 241.643
R1330 GNDA.n2555 GNDA.n2503 241.643
R1331 GNDA.n2563 GNDA.n2503 241.643
R1332 GNDA.n2600 GNDA.n2599 241.643
R1333 GNDA.n2600 GNDA.n2505 241.643
R1334 GNDA.n2600 GNDA.n2506 241.643
R1335 GNDA.n2600 GNDA.n2507 241.643
R1336 GNDA.n2600 GNDA.n2508 241.643
R1337 GNDA.n2600 GNDA.n2509 241.643
R1338 GNDA.n2213 GNDA.n2212 241.643
R1339 GNDA.n2213 GNDA.n2197 241.643
R1340 GNDA.n2388 GNDA.n2381 241.643
R1341 GNDA.n2388 GNDA.n2372 241.643
R1342 GNDA.n2459 GNDA.n2458 241.643
R1343 GNDA.n2459 GNDA.n2445 241.643
R1344 GNDA.n2302 GNDA.n2301 241.643
R1345 GNDA.n2302 GNDA.n2176 241.643
R1346 GNDA.n2612 GNDA.n2611 241.643
R1347 GNDA.n2612 GNDA.n2504 241.643
R1348 GNDA.n2628 GNDA.n2627 241.643
R1349 GNDA.n2628 GNDA.n11 241.643
R1350 GNDA.n2364 GNDA.n90 241.643
R1351 GNDA.n2403 GNDA.n2402 241.643
R1352 GNDA.n2388 GNDA.n2387 241.643
R1353 GNDA.n2460 GNDA.n2459 241.643
R1354 GNDA.n2489 GNDA.n33 241.643
R1355 GNDA.n2502 GNDA.n2501 241.643
R1356 GNDA.n2415 GNDA.n2414 241.643
R1357 GNDA.n2424 GNDA.n67 241.643
R1358 GNDA.n2442 GNDA.n2441 241.643
R1359 GNDA.n2442 GNDA.n68 241.643
R1360 GNDA.n2483 GNDA.n2482 241.643
R1361 GNDA.n2471 GNDA.n10 241.643
R1362 GNDA.n45 GNDA.n34 241.643
R1363 GNDA.n52 GNDA.n34 241.643
R1364 GNDA.n2131 GNDA.n2130 241.643
R1365 GNDA.n2130 GNDA.n136 241.643
R1366 GNDA.n223 GNDA.n208 241.643
R1367 GNDA.n223 GNDA.n209 241.643
R1368 GNDA.n76 GNDA.n74 206.052
R1369 GNDA.n19 GNDA.n17 206.052
R1370 GNDA.n82 GNDA.n81 205.488
R1371 GNDA.n80 GNDA.n79 205.488
R1372 GNDA.n78 GNDA.n77 205.488
R1373 GNDA.n76 GNDA.n75 205.488
R1374 GNDA.n25 GNDA.n24 205.488
R1375 GNDA.n23 GNDA.n22 205.488
R1376 GNDA.n21 GNDA.n20 205.488
R1377 GNDA.n19 GNDA.n18 205.488
R1378 GNDA.n84 GNDA.n83 200.988
R1379 GNDA.n27 GNDA.n26 200.988
R1380 GNDA.n1096 GNDA.n1095 197
R1381 GNDA.n1491 GNDA.n1490 197
R1382 GNDA.n823 GNDA.n291 197
R1383 GNDA.n1928 GNDA.n317 197
R1384 GNDA.n1849 GNDA.n1845 197
R1385 GNDA.n658 GNDA.n292 197
R1386 GNDA.n1391 GNDA.n1390 197
R1387 GNDA.n1035 GNDA.n1034 197
R1388 GNDA.n2021 GNDA.n177 197
R1389 GNDA.n1291 GNDA.n1290 197
R1390 GNDA.n1586 GNDA.n1585 187.249
R1391 GNDA.n912 GNDA.n423 187.249
R1392 GNDA.n1735 GNDA.n410 187.249
R1393 GNDA.n1920 GNDA.n1919 187.249
R1394 GNDA.n1967 GNDA.n289 187.249
R1395 GNDA.n1486 GNDA.n1485 187.249
R1396 GNDA.n1965 GNDA.n294 187.249
R1397 GNDA.n2093 GNDA.n172 187.249
R1398 GNDA.n1386 GNDA.n1385 187.249
R1399 GNDA.n2132 GNDA.n134 185
R1400 GNDA.n2124 GNDA.n2123 185
R1401 GNDA.n2348 GNDA.n2347 185
R1402 GNDA.n2314 GNDA.n2313 185
R1403 GNDA.n2361 GNDA.n2360 185
R1404 GNDA.n2398 GNDA.n2397 185
R1405 GNDA.n2380 GNDA.n2374 185
R1406 GNDA.n2457 GNDA.n2447 185
R1407 GNDA.n2486 GNDA.n2485 185
R1408 GNDA.n2497 GNDA.n2496 185
R1409 GNDA.n2299 GNDA.n2298 185
R1410 GNDA.n2297 GNDA.n2294 185
R1411 GNDA.n2210 GNDA.n2209 185
R1412 GNDA.n2208 GNDA.n2202 185
R1413 GNDA.n2413 GNDA.n2411 185
R1414 GNDA.n2423 GNDA.n2422 185
R1415 GNDA.n2440 GNDA.n72 185
R1416 GNDA.n2384 GNDA.n2383 185
R1417 GNDA.n47 GNDA.n46 185
R1418 GNDA.n2463 GNDA.n55 185
R1419 GNDA.n2481 GNDA.n38 185
R1420 GNDA.n2470 GNDA.n2469 185
R1421 GNDA.n64 GNDA.n60 185
R1422 GNDA.n2640 GNDA.n2638 185
R1423 GNDA.n2609 GNDA.n2608 185
R1424 GNDA.n2607 GNDA.n2604 185
R1425 GNDA.n2625 GNDA.n2624 185
R1426 GNDA.n2623 GNDA.n16 185
R1427 GNDA.n2597 GNDA.n2596 185
R1428 GNDA.n2595 GNDA.n2514 185
R1429 GNDA.n2593 GNDA.n2515 185
R1430 GNDA.n2590 GNDA.n2516 185
R1431 GNDA.n2589 GNDA.n2517 185
R1432 GNDA.n2586 GNDA.n2518 185
R1433 GNDA.n2585 GNDA.n2519 185
R1434 GNDA.n2582 GNDA.n2520 185
R1435 GNDA.n2581 GNDA.n2521 185
R1436 GNDA.n2578 GNDA.n2522 185
R1437 GNDA.n2539 GNDA.n2534 185
R1438 GNDA.n2541 GNDA.n2540 185
R1439 GNDA.n2532 GNDA.n2531 185
R1440 GNDA.n2548 GNDA.n2547 185
R1441 GNDA.n2549 GNDA.n2530 185
R1442 GNDA.n2551 GNDA.n2550 185
R1443 GNDA.n2528 GNDA.n2527 185
R1444 GNDA.n2558 GNDA.n2557 185
R1445 GNDA.n2559 GNDA.n2526 185
R1446 GNDA.n2561 GNDA.n2560 185
R1447 GNDA.n2287 GNDA.n2286 185
R1448 GNDA.n2285 GNDA.n2186 185
R1449 GNDA.n2283 GNDA.n2187 185
R1450 GNDA.n2280 GNDA.n2188 185
R1451 GNDA.n2279 GNDA.n2189 185
R1452 GNDA.n2276 GNDA.n2190 185
R1453 GNDA.n2275 GNDA.n2191 185
R1454 GNDA.n2272 GNDA.n2192 185
R1455 GNDA.n2271 GNDA.n2193 185
R1456 GNDA.n2268 GNDA.n2194 185
R1457 GNDA.n2251 GNDA.n2250 185
R1458 GNDA.n2249 GNDA.n2222 185
R1459 GNDA.n2247 GNDA.n2223 185
R1460 GNDA.n2244 GNDA.n2224 185
R1461 GNDA.n2243 GNDA.n2225 185
R1462 GNDA.n2240 GNDA.n2226 185
R1463 GNDA.n2239 GNDA.n2227 185
R1464 GNDA.n2236 GNDA.n2228 185
R1465 GNDA.n2235 GNDA.n2229 185
R1466 GNDA.n2232 GNDA.n2230 185
R1467 GNDA.n1558 GNDA.n1557 185
R1468 GNDA.n1560 GNDA.n1559 185
R1469 GNDA.n1562 GNDA.n1561 185
R1470 GNDA.n1564 GNDA.n1563 185
R1471 GNDA.n1566 GNDA.n1565 185
R1472 GNDA.n1568 GNDA.n1567 185
R1473 GNDA.n1570 GNDA.n1569 185
R1474 GNDA.n1571 GNDA.n467 185
R1475 GNDA.n1575 GNDA.n1574 185
R1476 GNDA.n1540 GNDA.n1539 185
R1477 GNDA.n1542 GNDA.n1541 185
R1478 GNDA.n1544 GNDA.n1543 185
R1479 GNDA.n1546 GNDA.n1545 185
R1480 GNDA.n1548 GNDA.n1547 185
R1481 GNDA.n1550 GNDA.n1549 185
R1482 GNDA.n1552 GNDA.n1551 185
R1483 GNDA.n1554 GNDA.n1553 185
R1484 GNDA.n1556 GNDA.n1555 185
R1485 GNDA.n1522 GNDA.n1521 185
R1486 GNDA.n1524 GNDA.n1523 185
R1487 GNDA.n1526 GNDA.n1525 185
R1488 GNDA.n1528 GNDA.n1527 185
R1489 GNDA.n1530 GNDA.n1529 185
R1490 GNDA.n1532 GNDA.n1531 185
R1491 GNDA.n1534 GNDA.n1533 185
R1492 GNDA.n1536 GNDA.n1535 185
R1493 GNDA.n1538 GNDA.n1537 185
R1494 GNDA.n1520 GNDA.n1519 185
R1495 GNDA.n1514 GNDA.n1513 185
R1496 GNDA.n1512 GNDA.n1511 185
R1497 GNDA.n1507 GNDA.n1506 185
R1498 GNDA.n1505 GNDA.n1504 185
R1499 GNDA.n1499 GNDA.n1498 185
R1500 GNDA.n1495 GNDA.n450 185
R1501 GNDA.n1579 GNDA.n1578 185
R1502 GNDA.n449 GNDA.n447 185
R1503 GNDA.n882 GNDA.n821 185
R1504 GNDA.n896 GNDA.n895 185
R1505 GNDA.n894 GNDA.n822 185
R1506 GNDA.n893 GNDA.n892 185
R1507 GNDA.n891 GNDA.n890 185
R1508 GNDA.n889 GNDA.n888 185
R1509 GNDA.n887 GNDA.n886 185
R1510 GNDA.n885 GNDA.n884 185
R1511 GNDA.n883 GNDA.n798 185
R1512 GNDA.n865 GNDA.n864 185
R1513 GNDA.n867 GNDA.n866 185
R1514 GNDA.n869 GNDA.n868 185
R1515 GNDA.n871 GNDA.n870 185
R1516 GNDA.n873 GNDA.n872 185
R1517 GNDA.n875 GNDA.n874 185
R1518 GNDA.n877 GNDA.n876 185
R1519 GNDA.n879 GNDA.n878 185
R1520 GNDA.n881 GNDA.n880 185
R1521 GNDA.n847 GNDA.n846 185
R1522 GNDA.n849 GNDA.n848 185
R1523 GNDA.n851 GNDA.n850 185
R1524 GNDA.n853 GNDA.n852 185
R1525 GNDA.n855 GNDA.n854 185
R1526 GNDA.n857 GNDA.n856 185
R1527 GNDA.n859 GNDA.n858 185
R1528 GNDA.n861 GNDA.n860 185
R1529 GNDA.n863 GNDA.n862 185
R1530 GNDA.n845 GNDA.n844 185
R1531 GNDA.n839 GNDA.n838 185
R1532 GNDA.n837 GNDA.n836 185
R1533 GNDA.n832 GNDA.n831 185
R1534 GNDA.n827 GNDA.n806 185
R1535 GNDA.n900 GNDA.n899 185
R1536 GNDA.n805 GNDA.n803 185
R1537 GNDA.n906 GNDA.n905 185
R1538 GNDA.n908 GNDA.n907 185
R1539 GNDA.n393 GNDA.n392 185
R1540 GNDA.n394 GNDA.n344 185
R1541 GNDA.n396 GNDA.n395 185
R1542 GNDA.n398 GNDA.n343 185
R1543 GNDA.n401 GNDA.n400 185
R1544 GNDA.n402 GNDA.n342 185
R1545 GNDA.n404 GNDA.n403 185
R1546 GNDA.n406 GNDA.n341 185
R1547 GNDA.n408 GNDA.n407 185
R1548 GNDA.n374 GNDA.n349 185
R1549 GNDA.n377 GNDA.n376 185
R1550 GNDA.n378 GNDA.n348 185
R1551 GNDA.n380 GNDA.n379 185
R1552 GNDA.n382 GNDA.n347 185
R1553 GNDA.n385 GNDA.n384 185
R1554 GNDA.n386 GNDA.n346 185
R1555 GNDA.n388 GNDA.n387 185
R1556 GNDA.n390 GNDA.n345 185
R1557 GNDA.n358 GNDA.n323 185
R1558 GNDA.n360 GNDA.n354 185
R1559 GNDA.n362 GNDA.n361 185
R1560 GNDA.n363 GNDA.n353 185
R1561 GNDA.n365 GNDA.n364 185
R1562 GNDA.n367 GNDA.n351 185
R1563 GNDA.n369 GNDA.n368 185
R1564 GNDA.n370 GNDA.n350 185
R1565 GNDA.n372 GNDA.n371 185
R1566 GNDA.n357 GNDA.n324 185
R1567 GNDA.n332 GNDA.n331 185
R1568 GNDA.n1761 GNDA.n1760 185
R1569 GNDA.n1758 GNDA.n329 185
R1570 GNDA.n1757 GNDA.n334 185
R1571 GNDA.n1755 GNDA.n1754 185
R1572 GNDA.n1746 GNDA.n335 185
R1573 GNDA.n1745 GNDA.n1744 185
R1574 GNDA.n1742 GNDA.n1741 185
R1575 GNDA.n1900 GNDA.n1899 185
R1576 GNDA.n1902 GNDA.n1901 185
R1577 GNDA.n1904 GNDA.n1903 185
R1578 GNDA.n1906 GNDA.n1905 185
R1579 GNDA.n1908 GNDA.n1907 185
R1580 GNDA.n1910 GNDA.n1909 185
R1581 GNDA.n1912 GNDA.n1911 185
R1582 GNDA.n1914 GNDA.n1913 185
R1583 GNDA.n1915 GNDA.n122 185
R1584 GNDA.n1882 GNDA.n1881 185
R1585 GNDA.n1884 GNDA.n1883 185
R1586 GNDA.n1886 GNDA.n1885 185
R1587 GNDA.n1888 GNDA.n1887 185
R1588 GNDA.n1890 GNDA.n1889 185
R1589 GNDA.n1892 GNDA.n1891 185
R1590 GNDA.n1894 GNDA.n1893 185
R1591 GNDA.n1896 GNDA.n1895 185
R1592 GNDA.n1898 GNDA.n1897 185
R1593 GNDA.n1864 GNDA.n1863 185
R1594 GNDA.n1866 GNDA.n1865 185
R1595 GNDA.n1868 GNDA.n1867 185
R1596 GNDA.n1870 GNDA.n1869 185
R1597 GNDA.n1872 GNDA.n1871 185
R1598 GNDA.n1874 GNDA.n1873 185
R1599 GNDA.n1876 GNDA.n1875 185
R1600 GNDA.n1878 GNDA.n1877 185
R1601 GNDA.n1880 GNDA.n1879 185
R1602 GNDA.n1862 GNDA.n1861 185
R1603 GNDA.n1853 GNDA.n1852 185
R1604 GNDA.n1851 GNDA.n105 185
R1605 GNDA.n2158 GNDA.n2157 185
R1606 GNDA.n2141 GNDA.n104 185
R1607 GNDA.n2145 GNDA.n2144 185
R1608 GNDA.n2143 GNDA.n2140 185
R1609 GNDA.n125 GNDA.n123 185
R1610 GNDA.n2154 GNDA.n2153 185
R1611 GNDA.n717 GNDA.n656 185
R1612 GNDA.n732 GNDA.n731 185
R1613 GNDA.n730 GNDA.n657 185
R1614 GNDA.n729 GNDA.n728 185
R1615 GNDA.n727 GNDA.n726 185
R1616 GNDA.n725 GNDA.n724 185
R1617 GNDA.n723 GNDA.n722 185
R1618 GNDA.n721 GNDA.n720 185
R1619 GNDA.n719 GNDA.n718 185
R1620 GNDA.n700 GNDA.n699 185
R1621 GNDA.n702 GNDA.n701 185
R1622 GNDA.n704 GNDA.n703 185
R1623 GNDA.n706 GNDA.n705 185
R1624 GNDA.n708 GNDA.n707 185
R1625 GNDA.n710 GNDA.n709 185
R1626 GNDA.n712 GNDA.n711 185
R1627 GNDA.n714 GNDA.n713 185
R1628 GNDA.n716 GNDA.n715 185
R1629 GNDA.n682 GNDA.n681 185
R1630 GNDA.n684 GNDA.n683 185
R1631 GNDA.n686 GNDA.n685 185
R1632 GNDA.n688 GNDA.n687 185
R1633 GNDA.n690 GNDA.n689 185
R1634 GNDA.n692 GNDA.n691 185
R1635 GNDA.n694 GNDA.n693 185
R1636 GNDA.n696 GNDA.n695 185
R1637 GNDA.n698 GNDA.n697 185
R1638 GNDA.n680 GNDA.n679 185
R1639 GNDA.n674 GNDA.n673 185
R1640 GNDA.n672 GNDA.n671 185
R1641 GNDA.n667 GNDA.n666 185
R1642 GNDA.n662 GNDA.n641 185
R1643 GNDA.n736 GNDA.n735 185
R1644 GNDA.n640 GNDA.n638 185
R1645 GNDA.n742 GNDA.n741 185
R1646 GNDA.n744 GNDA.n743 185
R1647 GNDA.n1459 GNDA.n1458 185
R1648 GNDA.n1461 GNDA.n1460 185
R1649 GNDA.n1463 GNDA.n1462 185
R1650 GNDA.n1465 GNDA.n1464 185
R1651 GNDA.n1467 GNDA.n1466 185
R1652 GNDA.n1469 GNDA.n1468 185
R1653 GNDA.n1471 GNDA.n1470 185
R1654 GNDA.n1473 GNDA.n1472 185
R1655 GNDA.n1474 GNDA.n473 185
R1656 GNDA.n1441 GNDA.n1440 185
R1657 GNDA.n1443 GNDA.n1442 185
R1658 GNDA.n1445 GNDA.n1444 185
R1659 GNDA.n1447 GNDA.n1446 185
R1660 GNDA.n1449 GNDA.n1448 185
R1661 GNDA.n1451 GNDA.n1450 185
R1662 GNDA.n1453 GNDA.n1452 185
R1663 GNDA.n1455 GNDA.n1454 185
R1664 GNDA.n1457 GNDA.n1456 185
R1665 GNDA.n1423 GNDA.n1422 185
R1666 GNDA.n1425 GNDA.n1424 185
R1667 GNDA.n1427 GNDA.n1426 185
R1668 GNDA.n1429 GNDA.n1428 185
R1669 GNDA.n1431 GNDA.n1430 185
R1670 GNDA.n1433 GNDA.n1432 185
R1671 GNDA.n1435 GNDA.n1434 185
R1672 GNDA.n1437 GNDA.n1436 185
R1673 GNDA.n1439 GNDA.n1438 185
R1674 GNDA.n1421 GNDA.n1420 185
R1675 GNDA.n1415 GNDA.n1414 185
R1676 GNDA.n1413 GNDA.n1412 185
R1677 GNDA.n1408 GNDA.n1407 185
R1678 GNDA.n1406 GNDA.n1405 185
R1679 GNDA.n1400 GNDA.n1399 185
R1680 GNDA.n1395 GNDA.n477 185
R1681 GNDA.n1478 GNDA.n1477 185
R1682 GNDA.n476 GNDA.n474 185
R1683 GNDA.n976 GNDA.n975 185
R1684 GNDA.n978 GNDA.n933 185
R1685 GNDA.n981 GNDA.n980 185
R1686 GNDA.n982 GNDA.n932 185
R1687 GNDA.n984 GNDA.n983 185
R1688 GNDA.n986 GNDA.n931 185
R1689 GNDA.n989 GNDA.n988 185
R1690 GNDA.n990 GNDA.n930 185
R1691 GNDA.n995 GNDA.n994 185
R1692 GNDA.n958 GNDA.n938 185
R1693 GNDA.n960 GNDA.n959 185
R1694 GNDA.n962 GNDA.n937 185
R1695 GNDA.n965 GNDA.n964 185
R1696 GNDA.n966 GNDA.n936 185
R1697 GNDA.n968 GNDA.n967 185
R1698 GNDA.n970 GNDA.n935 185
R1699 GNDA.n973 GNDA.n972 185
R1700 GNDA.n974 GNDA.n934 185
R1701 GNDA.n1029 GNDA.n1028 185
R1702 GNDA.n943 GNDA.n917 185
R1703 GNDA.n945 GNDA.n944 185
R1704 GNDA.n947 GNDA.n941 185
R1705 GNDA.n949 GNDA.n948 185
R1706 GNDA.n950 GNDA.n940 185
R1707 GNDA.n952 GNDA.n951 185
R1708 GNDA.n954 GNDA.n939 185
R1709 GNDA.n957 GNDA.n956 185
R1710 GNDA.n1027 GNDA.n916 185
R1711 GNDA.n1025 GNDA.n1024 185
R1712 GNDA.n920 GNDA.n919 185
R1713 GNDA.n1015 GNDA.n1014 185
R1714 GNDA.n1012 GNDA.n923 185
R1715 GNDA.n1010 GNDA.n1009 185
R1716 GNDA.n925 GNDA.n924 185
R1717 GNDA.n1000 GNDA.n999 185
R1718 GNDA.n997 GNDA.n929 185
R1719 GNDA.n2075 GNDA.n2074 185
R1720 GNDA.n2077 GNDA.n2076 185
R1721 GNDA.n2079 GNDA.n2078 185
R1722 GNDA.n2081 GNDA.n2080 185
R1723 GNDA.n2083 GNDA.n2082 185
R1724 GNDA.n2085 GNDA.n2084 185
R1725 GNDA.n2087 GNDA.n2086 185
R1726 GNDA.n2089 GNDA.n2088 185
R1727 GNDA.n2090 GNDA.n161 185
R1728 GNDA.n2057 GNDA.n2056 185
R1729 GNDA.n2059 GNDA.n2058 185
R1730 GNDA.n2061 GNDA.n2060 185
R1731 GNDA.n2063 GNDA.n2062 185
R1732 GNDA.n2065 GNDA.n2064 185
R1733 GNDA.n2067 GNDA.n2066 185
R1734 GNDA.n2069 GNDA.n2068 185
R1735 GNDA.n2071 GNDA.n2070 185
R1736 GNDA.n2073 GNDA.n2072 185
R1737 GNDA.n2039 GNDA.n2038 185
R1738 GNDA.n2041 GNDA.n2040 185
R1739 GNDA.n2043 GNDA.n2042 185
R1740 GNDA.n2045 GNDA.n2044 185
R1741 GNDA.n2047 GNDA.n2046 185
R1742 GNDA.n2049 GNDA.n2048 185
R1743 GNDA.n2051 GNDA.n2050 185
R1744 GNDA.n2053 GNDA.n2052 185
R1745 GNDA.n2055 GNDA.n2054 185
R1746 GNDA.n2037 GNDA.n2036 185
R1747 GNDA.n181 GNDA.n180 185
R1748 GNDA.n179 GNDA.n144 185
R1749 GNDA.n2116 GNDA.n2115 185
R1750 GNDA.n2099 GNDA.n143 185
R1751 GNDA.n2103 GNDA.n2102 185
R1752 GNDA.n2101 GNDA.n2098 185
R1753 GNDA.n164 GNDA.n162 185
R1754 GNDA.n2112 GNDA.n2111 185
R1755 GNDA.n1359 GNDA.n1358 185
R1756 GNDA.n1361 GNDA.n1360 185
R1757 GNDA.n1363 GNDA.n1362 185
R1758 GNDA.n1365 GNDA.n1364 185
R1759 GNDA.n1367 GNDA.n1366 185
R1760 GNDA.n1369 GNDA.n1368 185
R1761 GNDA.n1371 GNDA.n1370 185
R1762 GNDA.n1373 GNDA.n1372 185
R1763 GNDA.n1374 GNDA.n499 185
R1764 GNDA.n1341 GNDA.n1340 185
R1765 GNDA.n1343 GNDA.n1342 185
R1766 GNDA.n1345 GNDA.n1344 185
R1767 GNDA.n1347 GNDA.n1346 185
R1768 GNDA.n1349 GNDA.n1348 185
R1769 GNDA.n1351 GNDA.n1350 185
R1770 GNDA.n1353 GNDA.n1352 185
R1771 GNDA.n1355 GNDA.n1354 185
R1772 GNDA.n1357 GNDA.n1356 185
R1773 GNDA.n1323 GNDA.n1322 185
R1774 GNDA.n1325 GNDA.n1324 185
R1775 GNDA.n1327 GNDA.n1326 185
R1776 GNDA.n1329 GNDA.n1328 185
R1777 GNDA.n1331 GNDA.n1330 185
R1778 GNDA.n1333 GNDA.n1332 185
R1779 GNDA.n1335 GNDA.n1334 185
R1780 GNDA.n1337 GNDA.n1336 185
R1781 GNDA.n1339 GNDA.n1338 185
R1782 GNDA.n1321 GNDA.n1320 185
R1783 GNDA.n1315 GNDA.n1314 185
R1784 GNDA.n1313 GNDA.n1312 185
R1785 GNDA.n1308 GNDA.n1307 185
R1786 GNDA.n1306 GNDA.n1305 185
R1787 GNDA.n1300 GNDA.n1299 185
R1788 GNDA.n1295 GNDA.n503 185
R1789 GNDA.n1378 GNDA.n1377 185
R1790 GNDA.n502 GNDA.n500 185
R1791 GNDA.n211 GNDA.n129 185
R1792 GNDA.n219 GNDA.n211 185
R1793 GNDA.n217 GNDA.n129 185
R1794 GNDA.n217 GNDA.n216 185
R1795 GNDA.n1175 GNDA.n1174 183.948
R1796 GNDA.n1203 GNDA.n1202 183.948
R1797 GNDA.n1176 GNDA.n1175 180.013
R1798 GNDA.n1203 GNDA.n1079 180.013
R1799 GNDA.n425 GNDA.n424 175.546
R1800 GNDA.n1603 GNDA.n424 175.546
R1801 GNDA.n1601 GNDA.n1600 175.546
R1802 GNDA.n1597 GNDA.n1596 175.546
R1803 GNDA.n1593 GNDA.n1592 175.546
R1804 GNDA.n1589 GNDA.n1588 175.546
R1805 GNDA.n1153 GNDA.n426 175.546
R1806 GNDA.n1153 GNDA.n1151 175.546
R1807 GNDA.n1157 GNDA.n1151 175.546
R1808 GNDA.n1157 GNDA.n1149 175.546
R1809 GNDA.n1161 GNDA.n1149 175.546
R1810 GNDA.n1161 GNDA.n1147 175.546
R1811 GNDA.n1165 GNDA.n1147 175.546
R1812 GNDA.n1165 GNDA.n1145 175.546
R1813 GNDA.n1169 GNDA.n1145 175.546
R1814 GNDA.n1169 GNDA.n1106 175.546
R1815 GNDA.n1173 GNDA.n1106 175.546
R1816 GNDA.n1581 GNDA.n429 175.546
R1817 GNDA.n1496 GNDA.n446 175.546
R1818 GNDA.n1502 GNDA.n1501 175.546
R1819 GNDA.n1509 GNDA.n1508 175.546
R1820 GNDA.n1517 GNDA.n1516 175.546
R1821 GNDA.n1143 GNDA.n1107 175.546
R1822 GNDA.n1110 GNDA.n1107 175.546
R1823 GNDA.n1111 GNDA.n1110 175.546
R1824 GNDA.n1114 GNDA.n1111 175.546
R1825 GNDA.n1115 GNDA.n1114 175.546
R1826 GNDA.n1119 GNDA.n1115 175.546
R1827 GNDA.n1120 GNDA.n1119 175.546
R1828 GNDA.n1121 GNDA.n1120 175.546
R1829 GNDA.n1122 GNDA.n1121 175.546
R1830 GNDA.n1122 GNDA.n470 175.546
R1831 GNDA.n1489 GNDA.n470 175.546
R1832 GNDA.n778 GNDA.n777 175.546
R1833 GNDA.n782 GNDA.n781 175.546
R1834 GNDA.n786 GNDA.n785 175.546
R1835 GNDA.n790 GNDA.n789 175.546
R1836 GNDA.n794 GNDA.n793 175.546
R1837 GNDA.n770 GNDA.n769 175.546
R1838 GNDA.n766 GNDA.n765 175.546
R1839 GNDA.n762 GNDA.n761 175.546
R1840 GNDA.n758 GNDA.n757 175.546
R1841 GNDA.n754 GNDA.n257 175.546
R1842 GNDA.n799 GNDA.n753 175.546
R1843 GNDA.n903 GNDA.n902 175.546
R1844 GNDA.n829 GNDA.n828 175.546
R1845 GNDA.n834 GNDA.n833 175.546
R1846 GNDA.n842 GNDA.n841 175.546
R1847 GNDA.n279 GNDA.n270 175.546
R1848 GNDA.n272 GNDA.n271 175.546
R1849 GNDA.n274 GNDA.n273 175.546
R1850 GNDA.n276 GNDA.n275 175.546
R1851 GNDA.n278 GNDA.n277 175.546
R1852 GNDA.n1715 GNDA.n1713 175.546
R1853 GNDA.n1719 GNDA.n1614 175.546
R1854 GNDA.n1723 GNDA.n1721 175.546
R1855 GNDA.n1727 GNDA.n1612 175.546
R1856 GNDA.n1730 GNDA.n1729 175.546
R1857 GNDA.n1707 GNDA.n1706 175.546
R1858 GNDA.n1704 GNDA.n1619 175.546
R1859 GNDA.n1700 GNDA.n1699 175.546
R1860 GNDA.n1697 GNDA.n1622 175.546
R1861 GNDA.n1693 GNDA.n1692 175.546
R1862 GNDA.n1739 GNDA.n1735 175.546
R1863 GNDA.n1739 GNDA.n338 175.546
R1864 GNDA.n1748 GNDA.n338 175.546
R1865 GNDA.n1748 GNDA.n337 175.546
R1866 GNDA.n1752 GNDA.n337 175.546
R1867 GNDA.n1752 GNDA.n328 175.546
R1868 GNDA.n1763 GNDA.n328 175.546
R1869 GNDA.n1763 GNDA.n325 175.546
R1870 GNDA.n1767 GNDA.n325 175.546
R1871 GNDA.n1770 GNDA.n1767 175.546
R1872 GNDA.n1770 GNDA.n317 175.546
R1873 GNDA.n1656 GNDA.n1655 175.546
R1874 GNDA.n1661 GNDA.n1658 175.546
R1875 GNDA.n1664 GNDA.n1663 175.546
R1876 GNDA.n1668 GNDA.n1666 175.546
R1877 GNDA.n1925 GNDA.n320 175.546
R1878 GNDA.n1684 GNDA.n1683 175.546
R1879 GNDA.n1680 GNDA.n1679 175.546
R1880 GNDA.n1677 GNDA.n1660 175.546
R1881 GNDA.n1673 GNDA.n1671 175.546
R1882 GNDA.n1923 GNDA.n322 175.546
R1883 GNDA.n1650 GNDA.n1628 175.546
R1884 GNDA.n1646 GNDA.n1645 175.546
R1885 GNDA.n1643 GNDA.n1631 175.546
R1886 GNDA.n1639 GNDA.n1638 175.546
R1887 GNDA.n1636 GNDA.n1634 175.546
R1888 GNDA.n1919 GNDA.n126 175.546
R1889 GNDA.n2151 GNDA.n126 175.546
R1890 GNDA.n2151 GNDA.n127 175.546
R1891 GNDA.n2147 GNDA.n127 175.546
R1892 GNDA.n2147 GNDA.n101 175.546
R1893 GNDA.n2160 GNDA.n101 175.546
R1894 GNDA.n2160 GNDA.n102 175.546
R1895 GNDA.n1855 GNDA.n102 175.546
R1896 GNDA.n1855 GNDA.n1777 175.546
R1897 GNDA.n1859 GNDA.n1777 175.546
R1898 GNDA.n1859 GNDA.n1849 175.546
R1899 GNDA.n1789 GNDA.n300 175.546
R1900 GNDA.n1825 GNDA.n1824 175.546
R1901 GNDA.n1786 GNDA.n1785 175.546
R1902 GNDA.n1835 GNDA.n1834 175.546
R1903 GNDA.n1781 GNDA.n1780 175.546
R1904 GNDA.n1986 GNDA.n264 175.546
R1905 GNDA.n1982 GNDA.n269 175.546
R1906 GNDA.n1980 GNDA.n1979 175.546
R1907 GNDA.n1976 GNDA.n1975 175.546
R1908 GNDA.n1972 GNDA.n1971 175.546
R1909 GNDA.n528 GNDA.n527 175.546
R1910 GNDA.n532 GNDA.n531 175.546
R1911 GNDA.n536 GNDA.n535 175.546
R1912 GNDA.n540 GNDA.n539 175.546
R1913 GNDA.n544 GNDA.n543 175.546
R1914 GNDA.n746 GNDA.n632 175.546
R1915 GNDA.n739 GNDA.n738 175.546
R1916 GNDA.n664 GNDA.n663 175.546
R1917 GNDA.n669 GNDA.n668 175.546
R1918 GNDA.n677 GNDA.n676 175.546
R1919 GNDA.n553 GNDA.n550 175.546
R1920 GNDA.n556 GNDA.n555 175.546
R1921 GNDA.n561 GNDA.n560 175.546
R1922 GNDA.n564 GNDA.n563 175.546
R1923 GNDA.n568 GNDA.n567 175.546
R1924 GNDA.n1140 GNDA.n1103 175.546
R1925 GNDA.n1140 GNDA.n1109 175.546
R1926 GNDA.n1136 GNDA.n1109 175.546
R1927 GNDA.n1136 GNDA.n1113 175.546
R1928 GNDA.n1132 GNDA.n1113 175.546
R1929 GNDA.n1132 GNDA.n1131 175.546
R1930 GNDA.n1131 GNDA.n1130 175.546
R1931 GNDA.n1130 GNDA.n1117 175.546
R1932 GNDA.n1126 GNDA.n1117 175.546
R1933 GNDA.n1126 GNDA.n472 175.546
R1934 GNDA.n1487 GNDA.n472 175.546
R1935 GNDA.n1177 GNDA.n1101 175.546
R1936 GNDA.n1181 GNDA.n1101 175.546
R1937 GNDA.n1181 GNDA.n1099 175.546
R1938 GNDA.n1186 GNDA.n1099 175.546
R1939 GNDA.n1186 GNDA.n1089 175.546
R1940 GNDA.n1191 GNDA.n1089 175.546
R1941 GNDA.n1191 GNDA.n1088 175.546
R1942 GNDA.n1196 GNDA.n1088 175.546
R1943 GNDA.n1196 GNDA.n1086 175.546
R1944 GNDA.n1200 GNDA.n1086 175.546
R1945 GNDA.n1201 GNDA.n1200 175.546
R1946 GNDA.n1481 GNDA.n1480 175.546
R1947 GNDA.n1397 GNDA.n1396 175.546
R1948 GNDA.n1403 GNDA.n1402 175.546
R1949 GNDA.n1410 GNDA.n1409 175.546
R1950 GNDA.n1418 GNDA.n1417 175.546
R1951 GNDA.n1204 GNDA.n1082 175.546
R1952 GNDA.n1205 GNDA.n1204 175.546
R1953 GNDA.n1208 GNDA.n1205 175.546
R1954 GNDA.n1209 GNDA.n1208 175.546
R1955 GNDA.n1212 GNDA.n1209 175.546
R1956 GNDA.n1213 GNDA.n1212 175.546
R1957 GNDA.n1214 GNDA.n1213 175.546
R1958 GNDA.n1215 GNDA.n1214 175.546
R1959 GNDA.n1219 GNDA.n1215 175.546
R1960 GNDA.n1219 GNDA.n496 175.546
R1961 GNDA.n1389 GNDA.n496 175.546
R1962 GNDA.n589 GNDA.n588 175.546
R1963 GNDA.n588 GNDA.n587 175.546
R1964 GNDA.n584 GNDA.n583 175.546
R1965 GNDA.n581 GNDA.n558 175.546
R1966 GNDA.n577 GNDA.n575 175.546
R1967 GNDA.n573 GNDA.n293 175.546
R1968 GNDA.n597 GNDA.n596 175.546
R1969 GNDA.n601 GNDA.n600 175.546
R1970 GNDA.n605 GNDA.n604 175.546
R1971 GNDA.n609 GNDA.n608 175.546
R1972 GNDA.n613 GNDA.n612 175.546
R1973 GNDA.n1002 GNDA.n928 175.546
R1974 GNDA.n1006 GNDA.n1004 175.546
R1975 GNDA.n1017 GNDA.n922 175.546
R1976 GNDA.n1021 GNDA.n1019 175.546
R1977 GNDA.n1032 GNDA.n915 175.546
R1978 GNDA.n1057 GNDA.n523 175.546
R1979 GNDA.n1053 GNDA.n523 175.546
R1980 GNDA.n1053 GNDA.n617 175.546
R1981 GNDA.n1049 GNDA.n617 175.546
R1982 GNDA.n1049 GNDA.n618 175.546
R1983 GNDA.n1045 GNDA.n618 175.546
R1984 GNDA.n1045 GNDA.n1044 175.546
R1985 GNDA.n1044 GNDA.n620 175.546
R1986 GNDA.n1040 GNDA.n620 175.546
R1987 GNDA.n1040 GNDA.n622 175.546
R1988 GNDA.n626 GNDA.n622 175.546
R1989 GNDA.n1821 GNDA.n1819 175.546
R1990 GNDA.n1827 GNDA.n1787 175.546
R1991 GNDA.n1831 GNDA.n1829 175.546
R1992 GNDA.n1837 GNDA.n1783 175.546
R1993 GNDA.n1840 GNDA.n1839 175.546
R1994 GNDA.n1814 GNDA.n1790 175.546
R1995 GNDA.n1810 GNDA.n1809 175.546
R1996 GNDA.n1807 GNDA.n1793 175.546
R1997 GNDA.n1803 GNDA.n1802 175.546
R1998 GNDA.n1800 GNDA.n1797 175.546
R1999 GNDA.n2093 GNDA.n165 175.546
R2000 GNDA.n2109 GNDA.n165 175.546
R2001 GNDA.n2109 GNDA.n166 175.546
R2002 GNDA.n2105 GNDA.n166 175.546
R2003 GNDA.n2105 GNDA.n140 175.546
R2004 GNDA.n2118 GNDA.n140 175.546
R2005 GNDA.n2118 GNDA.n141 175.546
R2006 GNDA.n183 GNDA.n141 175.546
R2007 GNDA.n183 GNDA.n176 175.546
R2008 GNDA.n2034 GNDA.n176 175.546
R2009 GNDA.n2034 GNDA.n177 175.546
R2010 GNDA.n1998 GNDA.n200 175.546
R2011 GNDA.n2003 GNDA.n200 175.546
R2012 GNDA.n2003 GNDA.n197 175.546
R2013 GNDA.n2007 GNDA.n197 175.546
R2014 GNDA.n2008 GNDA.n2007 175.546
R2015 GNDA.n2009 GNDA.n2008 175.546
R2016 GNDA.n2009 GNDA.n195 175.546
R2017 GNDA.n2014 GNDA.n195 175.546
R2018 GNDA.n2014 GNDA.n192 175.546
R2019 GNDA.n2018 GNDA.n192 175.546
R2020 GNDA.n2019 GNDA.n2018 175.546
R2021 GNDA.n1238 GNDA.n1084 175.546
R2022 GNDA.n1234 GNDA.n1084 175.546
R2023 GNDA.n1234 GNDA.n1207 175.546
R2024 GNDA.n1230 GNDA.n1207 175.546
R2025 GNDA.n1230 GNDA.n1228 175.546
R2026 GNDA.n1228 GNDA.n1227 175.546
R2027 GNDA.n1227 GNDA.n1211 175.546
R2028 GNDA.n1223 GNDA.n1211 175.546
R2029 GNDA.n1223 GNDA.n1217 175.546
R2030 GNDA.n1217 GNDA.n498 175.546
R2031 GNDA.n1387 GNDA.n498 175.546
R2032 GNDA.n1243 GNDA.n1080 175.546
R2033 GNDA.n1243 GNDA.n1078 175.546
R2034 GNDA.n1247 GNDA.n1078 175.546
R2035 GNDA.n1247 GNDA.n1076 175.546
R2036 GNDA.n1251 GNDA.n1076 175.546
R2037 GNDA.n1251 GNDA.n1074 175.546
R2038 GNDA.n1255 GNDA.n1074 175.546
R2039 GNDA.n1255 GNDA.n1072 175.546
R2040 GNDA.n1259 GNDA.n1072 175.546
R2041 GNDA.n1259 GNDA.n1070 175.546
R2042 GNDA.n1263 GNDA.n1070 175.546
R2043 GNDA.n1381 GNDA.n1380 175.546
R2044 GNDA.n1297 GNDA.n1296 175.546
R2045 GNDA.n1303 GNDA.n1302 175.546
R2046 GNDA.n1310 GNDA.n1309 175.546
R2047 GNDA.n1318 GNDA.n1317 175.546
R2048 GNDA.n1267 GNDA.n1068 175.546
R2049 GNDA.n1267 GNDA.n1066 175.546
R2050 GNDA.n1272 GNDA.n1066 175.546
R2051 GNDA.n1272 GNDA.n1064 175.546
R2052 GNDA.n1276 GNDA.n1064 175.546
R2053 GNDA.n1277 GNDA.n1276 175.546
R2054 GNDA.n1279 GNDA.n1277 175.546
R2055 GNDA.n1279 GNDA.n1062 175.546
R2056 GNDA.n1284 GNDA.n1062 175.546
R2057 GNDA.n1284 GNDA.n1060 175.546
R2058 GNDA.n1288 GNDA.n1060 175.546
R2059 GNDA.n285 GNDA.n203 173.881
R2060 GNDA.t191 GNDA.n205 172.876
R2061 GNDA.t191 GNDA.n239 172.615
R2062 GNDA.n1988 GNDA.n203 171.624
R2063 GNDA.n1521 GNDA.n1520 163.333
R2064 GNDA.n846 GNDA.n845 163.333
R2065 GNDA.n358 GNDA.n357 163.333
R2066 GNDA.n1863 GNDA.n1862 163.333
R2067 GNDA.n681 GNDA.n680 163.333
R2068 GNDA.n1422 GNDA.n1421 163.333
R2069 GNDA.n1028 GNDA.n1027 163.333
R2070 GNDA.n2038 GNDA.n2037 163.333
R2071 GNDA.n1322 GNDA.n1321 163.333
R2072 GNDA.t66 GNDA.t300 153.578
R2073 GNDA.n2251 GNDA.n2222 150
R2074 GNDA.n2223 GNDA.n2222 150
R2075 GNDA.n2224 GNDA.n2223 150
R2076 GNDA.n2225 GNDA.n2224 150
R2077 GNDA.n2227 GNDA.n2226 150
R2078 GNDA.n2228 GNDA.n2227 150
R2079 GNDA.n2229 GNDA.n2228 150
R2080 GNDA.n2230 GNDA.n2229 150
R2081 GNDA.n2597 GNDA.n2514 150
R2082 GNDA.n2515 GNDA.n2514 150
R2083 GNDA.n2516 GNDA.n2515 150
R2084 GNDA.n2517 GNDA.n2516 150
R2085 GNDA.n2519 GNDA.n2518 150
R2086 GNDA.n2520 GNDA.n2519 150
R2087 GNDA.n2521 GNDA.n2520 150
R2088 GNDA.n2522 GNDA.n2521 150
R2089 GNDA.n2540 GNDA.n2539 150
R2090 GNDA.n2540 GNDA.n2531 150
R2091 GNDA.n2548 GNDA.n2531 150
R2092 GNDA.n2549 GNDA.n2548 150
R2093 GNDA.n2550 GNDA.n2527 150
R2094 GNDA.n2558 GNDA.n2527 150
R2095 GNDA.n2559 GNDA.n2558 150
R2096 GNDA.n2560 GNDA.n2559 150
R2097 GNDA.n2287 GNDA.n2186 150
R2098 GNDA.n2187 GNDA.n2186 150
R2099 GNDA.n2188 GNDA.n2187 150
R2100 GNDA.n2189 GNDA.n2188 150
R2101 GNDA.n2191 GNDA.n2190 150
R2102 GNDA.n2192 GNDA.n2191 150
R2103 GNDA.n2193 GNDA.n2192 150
R2104 GNDA.n2194 GNDA.n2193 150
R2105 GNDA.n1553 GNDA.n1552 150
R2106 GNDA.n1549 GNDA.n1548 150
R2107 GNDA.n1545 GNDA.n1544 150
R2108 GNDA.n1541 GNDA.n1540 150
R2109 GNDA.n1537 GNDA.n1536 150
R2110 GNDA.n1533 GNDA.n1532 150
R2111 GNDA.n1529 GNDA.n1528 150
R2112 GNDA.n1525 GNDA.n1524 150
R2113 GNDA.n1578 GNDA.n449 150
R2114 GNDA.n1498 GNDA.n450 150
R2115 GNDA.n1506 GNDA.n1505 150
R2116 GNDA.n1513 GNDA.n1512 150
R2117 GNDA.n1561 GNDA.n1560 150
R2118 GNDA.n1565 GNDA.n1564 150
R2119 GNDA.n1569 GNDA.n1568 150
R2120 GNDA.n1575 GNDA.n467 150
R2121 GNDA.n878 GNDA.n877 150
R2122 GNDA.n874 GNDA.n873 150
R2123 GNDA.n870 GNDA.n869 150
R2124 GNDA.n866 GNDA.n865 150
R2125 GNDA.n862 GNDA.n861 150
R2126 GNDA.n858 GNDA.n857 150
R2127 GNDA.n854 GNDA.n853 150
R2128 GNDA.n850 GNDA.n849 150
R2129 GNDA.n907 GNDA.n906 150
R2130 GNDA.n899 GNDA.n805 150
R2131 GNDA.n831 GNDA.n806 150
R2132 GNDA.n838 GNDA.n837 150
R2133 GNDA.n896 GNDA.n822 150
R2134 GNDA.n892 GNDA.n891 150
R2135 GNDA.n888 GNDA.n887 150
R2136 GNDA.n884 GNDA.n883 150
R2137 GNDA.n388 GNDA.n346 150
R2138 GNDA.n384 GNDA.n382 150
R2139 GNDA.n380 GNDA.n348 150
R2140 GNDA.n376 GNDA.n374 150
R2141 GNDA.n372 GNDA.n350 150
R2142 GNDA.n368 GNDA.n367 150
R2143 GNDA.n365 GNDA.n353 150
R2144 GNDA.n361 GNDA.n360 150
R2145 GNDA.n1744 GNDA.n1742 150
R2146 GNDA.n1755 GNDA.n335 150
R2147 GNDA.n1758 GNDA.n1757 150
R2148 GNDA.n1760 GNDA.n332 150
R2149 GNDA.n396 GNDA.n344 150
R2150 GNDA.n400 GNDA.n398 150
R2151 GNDA.n404 GNDA.n342 150
R2152 GNDA.n407 GNDA.n406 150
R2153 GNDA.n1895 GNDA.n1894 150
R2154 GNDA.n1891 GNDA.n1890 150
R2155 GNDA.n1887 GNDA.n1886 150
R2156 GNDA.n1883 GNDA.n1882 150
R2157 GNDA.n1879 GNDA.n1878 150
R2158 GNDA.n1875 GNDA.n1874 150
R2159 GNDA.n1871 GNDA.n1870 150
R2160 GNDA.n1867 GNDA.n1866 150
R2161 GNDA.n2154 GNDA.n123 150
R2162 GNDA.n2144 GNDA.n2143 150
R2163 GNDA.n2157 GNDA.n104 150
R2164 GNDA.n1852 GNDA.n105 150
R2165 GNDA.n1903 GNDA.n1902 150
R2166 GNDA.n1907 GNDA.n1906 150
R2167 GNDA.n1911 GNDA.n1910 150
R2168 GNDA.n1913 GNDA.n122 150
R2169 GNDA.n713 GNDA.n712 150
R2170 GNDA.n709 GNDA.n708 150
R2171 GNDA.n705 GNDA.n704 150
R2172 GNDA.n701 GNDA.n700 150
R2173 GNDA.n697 GNDA.n696 150
R2174 GNDA.n693 GNDA.n692 150
R2175 GNDA.n689 GNDA.n688 150
R2176 GNDA.n685 GNDA.n684 150
R2177 GNDA.n743 GNDA.n742 150
R2178 GNDA.n735 GNDA.n640 150
R2179 GNDA.n666 GNDA.n641 150
R2180 GNDA.n673 GNDA.n672 150
R2181 GNDA.n732 GNDA.n657 150
R2182 GNDA.n728 GNDA.n727 150
R2183 GNDA.n724 GNDA.n723 150
R2184 GNDA.n720 GNDA.n719 150
R2185 GNDA.n1454 GNDA.n1453 150
R2186 GNDA.n1450 GNDA.n1449 150
R2187 GNDA.n1446 GNDA.n1445 150
R2188 GNDA.n1442 GNDA.n1441 150
R2189 GNDA.n1438 GNDA.n1437 150
R2190 GNDA.n1434 GNDA.n1433 150
R2191 GNDA.n1430 GNDA.n1429 150
R2192 GNDA.n1426 GNDA.n1425 150
R2193 GNDA.n1477 GNDA.n476 150
R2194 GNDA.n1399 GNDA.n477 150
R2195 GNDA.n1407 GNDA.n1406 150
R2196 GNDA.n1414 GNDA.n1413 150
R2197 GNDA.n1462 GNDA.n1461 150
R2198 GNDA.n1466 GNDA.n1465 150
R2199 GNDA.n1470 GNDA.n1469 150
R2200 GNDA.n1474 GNDA.n1473 150
R2201 GNDA.n972 GNDA.n970 150
R2202 GNDA.n968 GNDA.n936 150
R2203 GNDA.n964 GNDA.n962 150
R2204 GNDA.n960 GNDA.n938 150
R2205 GNDA.n956 GNDA.n954 150
R2206 GNDA.n952 GNDA.n940 150
R2207 GNDA.n948 GNDA.n947 150
R2208 GNDA.n945 GNDA.n943 150
R2209 GNDA.n999 GNDA.n997 150
R2210 GNDA.n1010 GNDA.n924 150
R2211 GNDA.n1014 GNDA.n1012 150
R2212 GNDA.n1025 GNDA.n919 150
R2213 GNDA.n980 GNDA.n978 150
R2214 GNDA.n984 GNDA.n932 150
R2215 GNDA.n988 GNDA.n986 150
R2216 GNDA.n995 GNDA.n930 150
R2217 GNDA.n2070 GNDA.n2069 150
R2218 GNDA.n2066 GNDA.n2065 150
R2219 GNDA.n2062 GNDA.n2061 150
R2220 GNDA.n2058 GNDA.n2057 150
R2221 GNDA.n2054 GNDA.n2053 150
R2222 GNDA.n2050 GNDA.n2049 150
R2223 GNDA.n2046 GNDA.n2045 150
R2224 GNDA.n2042 GNDA.n2041 150
R2225 GNDA.n2112 GNDA.n162 150
R2226 GNDA.n2102 GNDA.n2101 150
R2227 GNDA.n2115 GNDA.n143 150
R2228 GNDA.n180 GNDA.n144 150
R2229 GNDA.n2078 GNDA.n2077 150
R2230 GNDA.n2082 GNDA.n2081 150
R2231 GNDA.n2086 GNDA.n2085 150
R2232 GNDA.n2088 GNDA.n161 150
R2233 GNDA.n1354 GNDA.n1353 150
R2234 GNDA.n1350 GNDA.n1349 150
R2235 GNDA.n1346 GNDA.n1345 150
R2236 GNDA.n1342 GNDA.n1341 150
R2237 GNDA.n1338 GNDA.n1337 150
R2238 GNDA.n1334 GNDA.n1333 150
R2239 GNDA.n1330 GNDA.n1329 150
R2240 GNDA.n1326 GNDA.n1325 150
R2241 GNDA.n1377 GNDA.n502 150
R2242 GNDA.n1299 GNDA.n503 150
R2243 GNDA.n1307 GNDA.n1306 150
R2244 GNDA.n1314 GNDA.n1313 150
R2245 GNDA.n1362 GNDA.n1361 150
R2246 GNDA.n1366 GNDA.n1365 150
R2247 GNDA.n1370 GNDA.n1369 150
R2248 GNDA.n1374 GNDA.n1373 150
R2249 GNDA.t89 GNDA.t50 147.84
R2250 GNDA.t312 GNDA.t298 144.321
R2251 GNDA.n312 GNDA.n311 139.077
R2252 GNDA.n314 GNDA.n313 139.077
R2253 GNDA.n316 GNDA.n315 139.077
R2254 GNDA.n1953 GNDA.n1952 139.077
R2255 GNDA.n1951 GNDA.n1950 139.077
R2256 GNDA.n1949 GNDA.n1948 139.077
R2257 GNDA.n1947 GNDA.n1946 139.077
R2258 GNDA.n1937 GNDA.n1936 139.077
R2259 GNDA.n1935 GNDA.n1934 139.077
R2260 GNDA.n187 GNDA.n186 139.077
R2261 GNDA.t76 GNDA.t290 139.041
R2262 GNDA.n2025 GNDA.t295 135.69
R2263 GNDA.n211 GNDA.n210 134.268
R2264 GNDA.n217 GNDA.n210 134.268
R2265 GNDA.n796 GNDA.n422 132.721
R2266 GNDA.n1732 GNDA.n1731 132.721
R2267 GNDA.n2030 GNDA.t232 130.001
R2268 GNDA.n1940 GNDA.t249 130.001
R2269 GNDA.n1943 GNDA.t226 130.001
R2270 GNDA.n1956 GNDA.t274 130.001
R2271 GNDA.n1931 GNDA.t252 130.001
R2272 GNDA.n309 GNDA.t246 130.001
R2273 GNDA.n1490 GNDA.n1489 124.832
R2274 GNDA.n291 GNDA.n287 124.832
R2275 GNDA.n1928 GNDA.n1927 124.832
R2276 GNDA.n1921 GNDA.n1920 124.832
R2277 GNDA.n1845 GNDA.n1844 124.832
R2278 GNDA.n1968 GNDA.n1967 124.832
R2279 GNDA.n570 GNDA.n292 124.832
R2280 GNDA.n1487 GNDA.n1486 124.832
R2281 GNDA.n1390 GNDA.n1389 124.832
R2282 GNDA.n1965 GNDA.n293 124.832
R2283 GNDA.n1842 GNDA.n172 124.832
R2284 GNDA.n1387 GNDA.n1386 124.832
R2285 GNDA.n130 GNDA.t291 115.948
R2286 GNDA.n1091 GNDA.t308 115.105
R2287 GNDA.n130 GNDA.t299 114.635
R2288 GNDA.n1092 GNDA.t1 114.635
R2289 GNDA.t210 GNDA.n90 103.665
R2290 GNDA.n2502 GNDA.t194 103.665
R2291 GNDA.t225 GNDA.n1847 101.942
R2292 GNDA.n2120 GNDA.n136 101.718
R2293 GNDA.n52 GNDA.n51 101.718
R2294 GNDA.n2435 GNDA.n68 101.718
R2295 GNDA.n2501 GNDA.n2500 101.718
R2296 GNDA.n2489 GNDA.n2488 101.718
R2297 GNDA.n2461 GNDA.n2460 101.718
R2298 GNDA.n2387 GNDA.n2386 101.718
R2299 GNDA.n2402 GNDA.n2401 101.718
R2300 GNDA.n2364 GNDA.n2363 101.718
R2301 GNDA.n2622 GNDA.n11 101.718
R2302 GNDA.n2606 GNDA.n2504 101.718
R2303 GNDA.n2296 GNDA.n2176 101.718
R2304 GNDA.n2453 GNDA.n2445 101.718
R2305 GNDA.n2376 GNDA.n2372 101.718
R2306 GNDA.n2207 GNDA.n2197 101.718
R2307 GNDA.n2594 GNDA.n2505 101.718
R2308 GNDA.n2591 GNDA.n2506 101.718
R2309 GNDA.n2587 GNDA.n2507 101.718
R2310 GNDA.n2583 GNDA.n2508 101.718
R2311 GNDA.n2579 GNDA.n2509 101.718
R2312 GNDA.n2543 GNDA.n2542 101.718
R2313 GNDA.n2546 GNDA.n2545 101.718
R2314 GNDA.n2553 GNDA.n2552 101.718
R2315 GNDA.n2556 GNDA.n2555 101.718
R2316 GNDA.n2563 GNDA.n2562 101.718
R2317 GNDA.n2284 GNDA.n2177 101.718
R2318 GNDA.n2281 GNDA.n2178 101.718
R2319 GNDA.n2277 GNDA.n2179 101.718
R2320 GNDA.n2273 GNDA.n2180 101.718
R2321 GNDA.n2269 GNDA.n2181 101.718
R2322 GNDA.n2319 GNDA.n2318 101.718
R2323 GNDA.n2353 GNDA.n2352 101.718
R2324 GNDA.n2248 GNDA.n2214 101.718
R2325 GNDA.n2245 GNDA.n2215 101.718
R2326 GNDA.n2241 GNDA.n2216 101.718
R2327 GNDA.n2237 GNDA.n2217 101.718
R2328 GNDA.n2233 GNDA.n2218 101.718
R2329 GNDA.n2253 GNDA.n2220 101.718
R2330 GNDA.n2246 GNDA.n2214 101.718
R2331 GNDA.n2242 GNDA.n2215 101.718
R2332 GNDA.n2238 GNDA.n2216 101.718
R2333 GNDA.n2234 GNDA.n2217 101.718
R2334 GNDA.n2218 GNDA.n2196 101.718
R2335 GNDA.n65 GNDA.n59 101.718
R2336 GNDA.n2641 GNDA.n5 101.718
R2337 GNDA.n2346 GNDA.n2345 101.718
R2338 GNDA.n2312 GNDA.n2311 101.718
R2339 GNDA.n2289 GNDA.n2184 101.718
R2340 GNDA.n2282 GNDA.n2177 101.718
R2341 GNDA.n2278 GNDA.n2178 101.718
R2342 GNDA.n2274 GNDA.n2179 101.718
R2343 GNDA.n2270 GNDA.n2180 101.718
R2344 GNDA.n2266 GNDA.n2181 101.718
R2345 GNDA.n2536 GNDA.n2535 101.718
R2346 GNDA.n2544 GNDA.n2543 101.718
R2347 GNDA.n2545 GNDA.n2529 101.718
R2348 GNDA.n2554 GNDA.n2553 101.718
R2349 GNDA.n2555 GNDA.n2525 101.718
R2350 GNDA.n2564 GNDA.n2563 101.718
R2351 GNDA.n2599 GNDA.n2512 101.718
R2352 GNDA.n2592 GNDA.n2505 101.718
R2353 GNDA.n2588 GNDA.n2506 101.718
R2354 GNDA.n2584 GNDA.n2507 101.718
R2355 GNDA.n2580 GNDA.n2508 101.718
R2356 GNDA.n2576 GNDA.n2509 101.718
R2357 GNDA.n2212 GNDA.n2200 101.718
R2358 GNDA.n2205 GNDA.n2197 101.718
R2359 GNDA.n2381 GNDA.n2373 101.718
R2360 GNDA.n2372 GNDA.n2371 101.718
R2361 GNDA.n2458 GNDA.n2446 101.718
R2362 GNDA.n2451 GNDA.n2445 101.718
R2363 GNDA.n2301 GNDA.n2292 101.718
R2364 GNDA.n2176 GNDA.n2175 101.718
R2365 GNDA.n2611 GNDA.n2602 101.718
R2366 GNDA.n2504 GNDA.n30 101.718
R2367 GNDA.n2627 GNDA.n14 101.718
R2368 GNDA.n2620 GNDA.n11 101.718
R2369 GNDA.n2414 GNDA.n87 101.718
R2370 GNDA.n2425 GNDA.n2424 101.718
R2371 GNDA.n2441 GNDA.n71 101.718
R2372 GNDA.n2482 GNDA.n37 101.718
R2373 GNDA.n2472 GNDA.n2471 101.718
R2374 GNDA.n45 GNDA.n44 101.718
R2375 GNDA.n2131 GNDA.n135 101.718
R2376 GNDA.n221 GNDA.n208 101.718
R2377 GNDA.n213 GNDA.n209 101.718
R2378 GNDA.n212 GNDA.n208 101.718
R2379 GNDA.t191 GNDA.n224 47.6748
R2380 GNDA.n2341 GNDA.n2340 99.0842
R2381 GNDA.n2339 GNDA.n2338 99.0842
R2382 GNDA.n2337 GNDA.n2336 99.0842
R2383 GNDA.n2335 GNDA.n2334 99.0842
R2384 GNDA.n2333 GNDA.n2332 99.0842
R2385 GNDA.n2331 GNDA.n2330 99.0842
R2386 GNDA.n2329 GNDA.n2328 99.0842
R2387 GNDA.n2327 GNDA.n2326 99.0842
R2388 GNDA.n2325 GNDA.n2324 99.0842
R2389 GNDA.n2323 GNDA.n2322 99.0842
R2390 GNDA.n2369 GNDA.n2368 99.0842
R2391 GNDA.n40 GNDA.n39 99.0842
R2392 GNDA.n1997 GNDA.t191 98.9756
R2393 GNDA.n1918 GNDA.n308 98.8538
R2394 GNDA.n2259 GNDA.n2258 94.601
R2395 GNDA.n2572 GNDA.n2571 94.601
R2396 GNDA.n2569 GNDA.n2568 94.601
R2397 GNDA.n2262 GNDA.n2261 94.601
R2398 GNDA.n2095 GNDA.n2094 92.6754
R2399 GNDA.t75 GNDA.t41 92.1471
R2400 GNDA.t122 GNDA.t75 92.1471
R2401 GNDA.t300 GNDA.t122 92.1471
R2402 GNDA.n2127 GNDA.n134 91.069
R2403 GNDA.n2122 GNDA.n134 91.069
R2404 GNDA.n2124 GNDA.n133 91.069
R2405 GNDA.n2125 GNDA.n2124 91.069
R2406 GNDA.n215 GNDA.n211 91.069
R2407 GNDA.n218 GNDA.n217 91.069
R2408 GNDA.t251 GNDA.n1768 90.616
R2409 GNDA.n2360 GNDA.n2359 90.4158
R2410 GNDA.n2349 GNDA.n2348 90.2704
R2411 GNDA.n2348 GNDA.n2342 90.2704
R2412 GNDA.n2315 GNDA.n2314 90.2704
R2413 GNDA.n2314 GNDA.n2308 90.2704
R2414 GNDA.n2399 GNDA.n2398 90.2704
R2415 GNDA.n2378 GNDA.n2374 90.2704
R2416 GNDA.n2374 GNDA.n2370 90.2704
R2417 GNDA.n2455 GNDA.n2447 90.2704
R2418 GNDA.n2450 GNDA.n2447 90.2704
R2419 GNDA.n2485 GNDA.n32 90.2704
R2420 GNDA.n2498 GNDA.n2497 90.2704
R2421 GNDA.n2411 GNDA.n86 90.2704
R2422 GNDA.n2422 GNDA.n2420 90.2704
R2423 GNDA.n2438 GNDA.n72 90.2704
R2424 GNDA.n2434 GNDA.n72 90.2704
R2425 GNDA.n2383 GNDA.n2382 90.2704
R2426 GNDA.n48 GNDA.n47 90.2704
R2427 GNDA.n47 GNDA.n41 90.2704
R2428 GNDA.n57 GNDA.n55 90.2704
R2429 GNDA.n2479 GNDA.n38 90.2704
R2430 GNDA.n2469 GNDA.n2467 90.2704
R2431 GNDA.n62 GNDA.n60 90.2704
R2432 GNDA.n2638 GNDA.n4 90.2704
R2433 GNDA.t0 GNDA.n1058 89.6052
R2434 GNDA.n1152 GNDA.n227 88.5317
R2435 GNDA.n1152 GNDA.n1150 88.5317
R2436 GNDA.n1158 GNDA.n1150 88.5317
R2437 GNDA.n1159 GNDA.n1158 88.5317
R2438 GNDA.n1160 GNDA.n1159 88.5317
R2439 GNDA.n1166 GNDA.n1146 88.5317
R2440 GNDA.n1167 GNDA.n1166 88.5317
R2441 GNDA.n1168 GNDA.n1167 88.5317
R2442 GNDA.n1168 GNDA.n1105 88.5317
R2443 GNDA.n1174 GNDA.n1105 88.5317
R2444 GNDA.n1176 GNDA.n1100 88.5317
R2445 GNDA.n1182 GNDA.n1100 88.5317
R2446 GNDA.n1183 GNDA.n1182 88.5317
R2447 GNDA.n1185 GNDA.n1183 88.5317
R2448 GNDA.n1185 GNDA.n1184 88.5317
R2449 GNDA.n1193 GNDA.n1192 88.5317
R2450 GNDA.n1195 GNDA.n1193 88.5317
R2451 GNDA.n1195 GNDA.n1194 88.5317
R2452 GNDA.n1194 GNDA.n1085 88.5317
R2453 GNDA.n1202 GNDA.n1085 88.5317
R2454 GNDA.n1244 GNDA.n1079 88.5317
R2455 GNDA.n1245 GNDA.n1244 88.5317
R2456 GNDA.n1246 GNDA.n1245 88.5317
R2457 GNDA.n1246 GNDA.n1075 88.5317
R2458 GNDA.n1252 GNDA.n1075 88.5317
R2459 GNDA.n1254 GNDA.n1253 88.5317
R2460 GNDA.n1254 GNDA.n1071 88.5317
R2461 GNDA.n1260 GNDA.n1071 88.5317
R2462 GNDA.n1261 GNDA.n1260 88.5317
R2463 GNDA.n1262 GNDA.n1261 88.5317
R2464 GNDA.t147 GNDA.n167 85.4674
R2465 GNDA.t61 GNDA.t80 84.4682
R2466 GNDA.t297 GNDA.t85 84.4682
R2467 GNDA.t97 GNDA.t292 84.4682
R2468 GNDA.t32 GNDA.t49 84.4682
R2469 GNDA.t121 GNDA.t265 84.4682
R2470 GNDA.t115 GNDA.t131 84.4682
R2471 GNDA.t56 GNDA.t133 84.4682
R2472 GNDA.t282 GNDA.t127 84.4682
R2473 GNDA.t63 GNDA.t301 84.4682
R2474 GNDA.t302 GNDA.t68 84.4682
R2475 GNDA.t119 GNDA.t306 84.4682
R2476 GNDA.t88 GNDA.t293 84.4682
R2477 GNDA.n2148 GNDA.t168 84.4377
R2478 GNDA.n1095 GNDA.n1094 84.306
R2479 GNDA.t34 GNDA.t92 82.3782
R2480 GNDA.t294 GNDA.t47 82.3782
R2481 GNDA.n1237 GNDA.n1203 80.9821
R2482 GNDA.n1175 GNDA.n1104 80.9821
R2483 GNDA.t25 GNDA.t98 80.6288
R2484 GNDA.t67 GNDA.t135 80.6288
R2485 GNDA.n1850 GNDA.t158 80.3188
R2486 GNDA.n2302 GNDA.n2290 76.7893
R2487 GNDA.t218 GNDA.t5 76.7893
R2488 GNDA.t270 GNDA.t110 76.7893
R2489 GNDA.n2612 GNDA.n2503 76.7893
R2490 GNDA.t191 GNDA.n203 76.3879
R2491 GNDA.n1609 GNDA.n1608 76.3222
R2492 GNDA.n1603 GNDA.n412 76.3222
R2493 GNDA.n1600 GNDA.n413 76.3222
R2494 GNDA.n1596 GNDA.n414 76.3222
R2495 GNDA.n1592 GNDA.n415 76.3222
R2496 GNDA.n1585 GNDA.n1584 76.3222
R2497 GNDA.n1582 GNDA.n1581 76.3222
R2498 GNDA.n1496 GNDA.n445 76.3222
R2499 GNDA.n1502 GNDA.n444 76.3222
R2500 GNDA.n1508 GNDA.n443 76.3222
R2501 GNDA.n1517 GNDA.n442 76.3222
R2502 GNDA.n774 GNDA.n417 76.3222
R2503 GNDA.n778 GNDA.n418 76.3222
R2504 GNDA.n782 GNDA.n419 76.3222
R2505 GNDA.n786 GNDA.n420 76.3222
R2506 GNDA.n790 GNDA.n421 76.3222
R2507 GNDA.n794 GNDA.n422 76.3222
R2508 GNDA.n770 GNDA.n252 76.3222
R2509 GNDA.n766 GNDA.n253 76.3222
R2510 GNDA.n762 GNDA.n254 76.3222
R2511 GNDA.n758 GNDA.n255 76.3222
R2512 GNDA.n754 GNDA.n256 76.3222
R2513 GNDA.n1995 GNDA.n1994 76.3222
R2514 GNDA.n913 GNDA.n912 76.3222
R2515 GNDA.n799 GNDA.n752 76.3222
R2516 GNDA.n902 GNDA.n751 76.3222
R2517 GNDA.n829 GNDA.n750 76.3222
R2518 GNDA.n833 GNDA.n749 76.3222
R2519 GNDA.n842 GNDA.n748 76.3222
R2520 GNDA.n280 GNDA.n258 76.3222
R2521 GNDA.n281 GNDA.n270 76.3222
R2522 GNDA.n282 GNDA.n272 76.3222
R2523 GNDA.n283 GNDA.n274 76.3222
R2524 GNDA.n284 GNDA.n276 76.3222
R2525 GNDA.n286 GNDA.n278 76.3222
R2526 GNDA.n1712 GNDA.n1711 76.3222
R2527 GNDA.n1715 GNDA.n1714 76.3222
R2528 GNDA.n1720 GNDA.n1719 76.3222
R2529 GNDA.n1723 GNDA.n1722 76.3222
R2530 GNDA.n1728 GNDA.n1727 76.3222
R2531 GNDA.n1731 GNDA.n1730 76.3222
R2532 GNDA.n1707 GNDA.n1618 76.3222
R2533 GNDA.n1705 GNDA.n1704 76.3222
R2534 GNDA.n1700 GNDA.n1621 76.3222
R2535 GNDA.n1698 GNDA.n1697 76.3222
R2536 GNDA.n1693 GNDA.n1624 76.3222
R2537 GNDA.n1691 GNDA.n1690 76.3222
R2538 GNDA.n1654 GNDA.n1625 76.3222
R2539 GNDA.n1657 GNDA.n1656 76.3222
R2540 GNDA.n1662 GNDA.n1661 76.3222
R2541 GNDA.n1665 GNDA.n1664 76.3222
R2542 GNDA.n1668 GNDA.n1667 76.3222
R2543 GNDA.n1926 GNDA.n1925 76.3222
R2544 GNDA.n1686 GNDA.n1685 76.3222
R2545 GNDA.n1683 GNDA.n1653 76.3222
R2546 GNDA.n1679 GNDA.n1678 76.3222
R2547 GNDA.n1672 GNDA.n1660 76.3222
R2548 GNDA.n1671 GNDA.n1670 76.3222
R2549 GNDA.n1923 GNDA.n1922 76.3222
R2550 GNDA.n1651 GNDA.n1650 76.3222
R2551 GNDA.n1646 GNDA.n1630 76.3222
R2552 GNDA.n1644 GNDA.n1643 76.3222
R2553 GNDA.n1639 GNDA.n1633 76.3222
R2554 GNDA.n1637 GNDA.n1636 76.3222
R2555 GNDA.n1961 GNDA.n299 76.3222
R2556 GNDA.n1960 GNDA.n1959 76.3222
R2557 GNDA.n1789 GNDA.n301 76.3222
R2558 GNDA.n1825 GNDA.n302 76.3222
R2559 GNDA.n1786 GNDA.n303 76.3222
R2560 GNDA.n1835 GNDA.n304 76.3222
R2561 GNDA.n1780 GNDA.n305 76.3222
R2562 GNDA.n1990 GNDA.n1989 76.3222
R2563 GNDA.n1987 GNDA.n1986 76.3222
R2564 GNDA.n1982 GNDA.n268 76.3222
R2565 GNDA.n1979 GNDA.n267 76.3222
R2566 GNDA.n1975 GNDA.n266 76.3222
R2567 GNDA.n1971 GNDA.n265 76.3222
R2568 GNDA.n527 GNDA.n246 76.3222
R2569 GNDA.n531 GNDA.n247 76.3222
R2570 GNDA.n535 GNDA.n248 76.3222
R2571 GNDA.n539 GNDA.n249 76.3222
R2572 GNDA.n543 GNDA.n250 76.3222
R2573 GNDA.n547 GNDA.n251 76.3222
R2574 GNDA.n747 GNDA.n289 76.3222
R2575 GNDA.n632 GNDA.n631 76.3222
R2576 GNDA.n738 GNDA.n630 76.3222
R2577 GNDA.n664 GNDA.n629 76.3222
R2578 GNDA.n668 GNDA.n628 76.3222
R2579 GNDA.n677 GNDA.n627 76.3222
R2580 GNDA.n549 GNDA.n548 76.3222
R2581 GNDA.n554 GNDA.n553 76.3222
R2582 GNDA.n559 GNDA.n556 76.3222
R2583 GNDA.n562 GNDA.n561 76.3222
R2584 GNDA.n566 GNDA.n564 76.3222
R2585 GNDA.n569 GNDA.n568 76.3222
R2586 GNDA.n1485 GNDA.n441 76.3222
R2587 GNDA.n1480 GNDA.n440 76.3222
R2588 GNDA.n1397 GNDA.n439 76.3222
R2589 GNDA.n1403 GNDA.n438 76.3222
R2590 GNDA.n1409 GNDA.n437 76.3222
R2591 GNDA.n1418 GNDA.n436 76.3222
R2592 GNDA.n592 GNDA.n525 76.3222
R2593 GNDA.n587 GNDA.n552 76.3222
R2594 GNDA.n583 GNDA.n582 76.3222
R2595 GNDA.n576 GNDA.n558 76.3222
R2596 GNDA.n575 GNDA.n574 76.3222
R2597 GNDA.n596 GNDA.n240 76.3222
R2598 GNDA.n600 GNDA.n241 76.3222
R2599 GNDA.n604 GNDA.n242 76.3222
R2600 GNDA.n608 GNDA.n243 76.3222
R2601 GNDA.n612 GNDA.n244 76.3222
R2602 GNDA.n522 GNDA.n245 76.3222
R2603 GNDA.n927 GNDA.n294 76.3222
R2604 GNDA.n1003 GNDA.n1002 76.3222
R2605 GNDA.n1006 GNDA.n1005 76.3222
R2606 GNDA.n1018 GNDA.n1017 76.3222
R2607 GNDA.n1021 GNDA.n1020 76.3222
R2608 GNDA.n1033 GNDA.n1032 76.3222
R2609 GNDA.n1818 GNDA.n1817 76.3222
R2610 GNDA.n1821 GNDA.n1820 76.3222
R2611 GNDA.n1828 GNDA.n1827 76.3222
R2612 GNDA.n1831 GNDA.n1830 76.3222
R2613 GNDA.n1838 GNDA.n1837 76.3222
R2614 GNDA.n1841 GNDA.n1840 76.3222
R2615 GNDA.n1815 GNDA.n1814 76.3222
R2616 GNDA.n1810 GNDA.n1792 76.3222
R2617 GNDA.n1808 GNDA.n1807 76.3222
R2618 GNDA.n1803 GNDA.n1795 76.3222
R2619 GNDA.n1801 GNDA.n1800 76.3222
R2620 GNDA.n1796 GNDA.n202 76.3222
R2621 GNDA.n1385 GNDA.n435 76.3222
R2622 GNDA.n1380 GNDA.n434 76.3222
R2623 GNDA.n1297 GNDA.n433 76.3222
R2624 GNDA.n1303 GNDA.n432 76.3222
R2625 GNDA.n1309 GNDA.n431 76.3222
R2626 GNDA.n1318 GNDA.n430 76.3222
R2627 GNDA.n570 GNDA.n569 76.3222
R2628 GNDA.n567 GNDA.n566 76.3222
R2629 GNDA.n563 GNDA.n562 76.3222
R2630 GNDA.n560 GNDA.n559 76.3222
R2631 GNDA.n555 GNDA.n554 76.3222
R2632 GNDA.n550 GNDA.n549 76.3222
R2633 GNDA.n589 GNDA.n525 76.3222
R2634 GNDA.n584 GNDA.n552 76.3222
R2635 GNDA.n582 GNDA.n581 76.3222
R2636 GNDA.n577 GNDA.n576 76.3222
R2637 GNDA.n574 GNDA.n573 76.3222
R2638 GNDA.n1844 GNDA.n305 76.3222
R2639 GNDA.n1781 GNDA.n304 76.3222
R2640 GNDA.n1834 GNDA.n303 76.3222
R2641 GNDA.n1785 GNDA.n302 76.3222
R2642 GNDA.n1824 GNDA.n301 76.3222
R2643 GNDA.n1959 GNDA.n300 76.3222
R2644 GNDA.n1819 GNDA.n1818 76.3222
R2645 GNDA.n1820 GNDA.n1787 76.3222
R2646 GNDA.n1829 GNDA.n1828 76.3222
R2647 GNDA.n1830 GNDA.n1783 76.3222
R2648 GNDA.n1839 GNDA.n1838 76.3222
R2649 GNDA.n1842 GNDA.n1841 76.3222
R2650 GNDA.n1927 GNDA.n1926 76.3222
R2651 GNDA.n1667 GNDA.n320 76.3222
R2652 GNDA.n1666 GNDA.n1665 76.3222
R2653 GNDA.n1663 GNDA.n1662 76.3222
R2654 GNDA.n1658 GNDA.n1657 76.3222
R2655 GNDA.n1655 GNDA.n1654 76.3222
R2656 GNDA.n1685 GNDA.n1684 76.3222
R2657 GNDA.n1680 GNDA.n1653 76.3222
R2658 GNDA.n1678 GNDA.n1677 76.3222
R2659 GNDA.n1673 GNDA.n1672 76.3222
R2660 GNDA.n1670 GNDA.n322 76.3222
R2661 GNDA.n1922 GNDA.n1921 76.3222
R2662 GNDA.n287 GNDA.n286 76.3222
R2663 GNDA.n284 GNDA.n277 76.3222
R2664 GNDA.n283 GNDA.n275 76.3222
R2665 GNDA.n282 GNDA.n273 76.3222
R2666 GNDA.n281 GNDA.n271 76.3222
R2667 GNDA.n280 GNDA.n279 76.3222
R2668 GNDA.n1989 GNDA.n264 76.3222
R2669 GNDA.n1987 GNDA.n269 76.3222
R2670 GNDA.n1980 GNDA.n268 76.3222
R2671 GNDA.n1976 GNDA.n267 76.3222
R2672 GNDA.n1972 GNDA.n266 76.3222
R2673 GNDA.n1968 GNDA.n265 76.3222
R2674 GNDA.n1995 GNDA.n257 76.3222
R2675 GNDA.n757 GNDA.n256 76.3222
R2676 GNDA.n761 GNDA.n255 76.3222
R2677 GNDA.n765 GNDA.n254 76.3222
R2678 GNDA.n769 GNDA.n253 76.3222
R2679 GNDA.n773 GNDA.n252 76.3222
R2680 GNDA.n544 GNDA.n251 76.3222
R2681 GNDA.n540 GNDA.n250 76.3222
R2682 GNDA.n536 GNDA.n249 76.3222
R2683 GNDA.n532 GNDA.n248 76.3222
R2684 GNDA.n528 GNDA.n247 76.3222
R2685 GNDA.n263 GNDA.n246 76.3222
R2686 GNDA.n613 GNDA.n245 76.3222
R2687 GNDA.n609 GNDA.n244 76.3222
R2688 GNDA.n605 GNDA.n243 76.3222
R2689 GNDA.n601 GNDA.n242 76.3222
R2690 GNDA.n597 GNDA.n241 76.3222
R2691 GNDA.n593 GNDA.n240 76.3222
R2692 GNDA.n1584 GNDA.n429 76.3222
R2693 GNDA.n1582 GNDA.n446 76.3222
R2694 GNDA.n1501 GNDA.n445 76.3222
R2695 GNDA.n1509 GNDA.n444 76.3222
R2696 GNDA.n1516 GNDA.n443 76.3222
R2697 GNDA.n1491 GNDA.n442 76.3222
R2698 GNDA.n1481 GNDA.n441 76.3222
R2699 GNDA.n1396 GNDA.n440 76.3222
R2700 GNDA.n1402 GNDA.n439 76.3222
R2701 GNDA.n1410 GNDA.n438 76.3222
R2702 GNDA.n1417 GNDA.n437 76.3222
R2703 GNDA.n1391 GNDA.n436 76.3222
R2704 GNDA.n1381 GNDA.n435 76.3222
R2705 GNDA.n1296 GNDA.n434 76.3222
R2706 GNDA.n1302 GNDA.n433 76.3222
R2707 GNDA.n1310 GNDA.n432 76.3222
R2708 GNDA.n1317 GNDA.n431 76.3222
R2709 GNDA.n1291 GNDA.n430 76.3222
R2710 GNDA.n1692 GNDA.n1691 76.3222
R2711 GNDA.n1624 GNDA.n1622 76.3222
R2712 GNDA.n1699 GNDA.n1698 76.3222
R2713 GNDA.n1621 GNDA.n1619 76.3222
R2714 GNDA.n1706 GNDA.n1705 76.3222
R2715 GNDA.n1618 GNDA.n1616 76.3222
R2716 GNDA.n1634 GNDA.n299 76.3222
R2717 GNDA.n1638 GNDA.n1637 76.3222
R2718 GNDA.n1633 GNDA.n1631 76.3222
R2719 GNDA.n1645 GNDA.n1644 76.3222
R2720 GNDA.n1630 GNDA.n1628 76.3222
R2721 GNDA.n1652 GNDA.n1651 76.3222
R2722 GNDA.n1797 GNDA.n1796 76.3222
R2723 GNDA.n1802 GNDA.n1801 76.3222
R2724 GNDA.n1795 GNDA.n1793 76.3222
R2725 GNDA.n1809 GNDA.n1808 76.3222
R2726 GNDA.n1792 GNDA.n1790 76.3222
R2727 GNDA.n1816 GNDA.n1815 76.3222
R2728 GNDA.n913 GNDA.n753 76.3222
R2729 GNDA.n903 GNDA.n752 76.3222
R2730 GNDA.n828 GNDA.n751 76.3222
R2731 GNDA.n834 GNDA.n750 76.3222
R2732 GNDA.n841 GNDA.n749 76.3222
R2733 GNDA.n823 GNDA.n748 76.3222
R2734 GNDA.n747 GNDA.n746 76.3222
R2735 GNDA.n739 GNDA.n631 76.3222
R2736 GNDA.n663 GNDA.n630 76.3222
R2737 GNDA.n669 GNDA.n629 76.3222
R2738 GNDA.n676 GNDA.n628 76.3222
R2739 GNDA.n658 GNDA.n627 76.3222
R2740 GNDA.n928 GNDA.n927 76.3222
R2741 GNDA.n1004 GNDA.n1003 76.3222
R2742 GNDA.n1005 GNDA.n922 76.3222
R2743 GNDA.n1019 GNDA.n1018 76.3222
R2744 GNDA.n1020 GNDA.n915 76.3222
R2745 GNDA.n1034 GNDA.n1033 76.3222
R2746 GNDA.n1713 GNDA.n1712 76.3222
R2747 GNDA.n1714 GNDA.n1614 76.3222
R2748 GNDA.n1721 GNDA.n1720 76.3222
R2749 GNDA.n1722 GNDA.n1612 76.3222
R2750 GNDA.n1729 GNDA.n1728 76.3222
R2751 GNDA.n777 GNDA.n417 76.3222
R2752 GNDA.n781 GNDA.n418 76.3222
R2753 GNDA.n785 GNDA.n419 76.3222
R2754 GNDA.n789 GNDA.n420 76.3222
R2755 GNDA.n793 GNDA.n421 76.3222
R2756 GNDA.n1609 GNDA.n425 76.3222
R2757 GNDA.n1601 GNDA.n412 76.3222
R2758 GNDA.n1597 GNDA.n413 76.3222
R2759 GNDA.n1593 GNDA.n414 76.3222
R2760 GNDA.n1589 GNDA.n415 76.3222
R2761 GNDA.t261 GNDA.n2225 75.0005
R2762 GNDA.n2226 GNDA.t261 75.0005
R2763 GNDA.n2299 GNDA.t266 75.0005
R2764 GNDA.n2294 GNDA.t266 75.0005
R2765 GNDA.n2210 GNDA.t256 75.0005
R2766 GNDA.n2202 GNDA.t256 75.0005
R2767 GNDA.n2609 GNDA.t283 75.0005
R2768 GNDA.n2604 GNDA.t283 75.0005
R2769 GNDA.n2625 GNDA.t200 75.0005
R2770 GNDA.n16 GNDA.t200 75.0005
R2771 GNDA.t206 GNDA.n2517 75.0005
R2772 GNDA.n2518 GNDA.t206 75.0005
R2773 GNDA.t229 GNDA.n2549 75.0005
R2774 GNDA.n2550 GNDA.t229 75.0005
R2775 GNDA.t243 GNDA.n2189 75.0005
R2776 GNDA.n2190 GNDA.t243 75.0005
R2777 GNDA.n1540 GNDA.n456 74.5978
R2778 GNDA.n1537 GNDA.n456 74.5978
R2779 GNDA.n865 GNDA.n811 74.5978
R2780 GNDA.n862 GNDA.n811 74.5978
R2781 GNDA.n374 GNDA.n373 74.5978
R2782 GNDA.n373 GNDA.n372 74.5978
R2783 GNDA.n1882 GNDA.n111 74.5978
R2784 GNDA.n1879 GNDA.n111 74.5978
R2785 GNDA.n700 GNDA.n646 74.5978
R2786 GNDA.n697 GNDA.n646 74.5978
R2787 GNDA.n1441 GNDA.n483 74.5978
R2788 GNDA.n1438 GNDA.n483 74.5978
R2789 GNDA.n955 GNDA.n938 74.5978
R2790 GNDA.n956 GNDA.n955 74.5978
R2791 GNDA.n2057 GNDA.n150 74.5978
R2792 GNDA.n2054 GNDA.n150 74.5978
R2793 GNDA.n1341 GNDA.n509 74.5978
R2794 GNDA.n1338 GNDA.n509 74.5978
R2795 GNDA.t174 GNDA.n1857 74.1404
R2796 GNDA.t98 GNDA.t105 72.9499
R2797 GNDA.t10 GNDA.t287 72.9499
R2798 GNDA.t142 GNDA.t67 72.9499
R2799 GNDA.n2150 GNDA.t170 70.0216
R2800 GNDA.n1576 GNDA.n449 69.3109
R2801 GNDA.n1576 GNDA.n1575 69.3109
R2802 GNDA.n907 GNDA.n801 69.3109
R2803 GNDA.n883 GNDA.n801 69.3109
R2804 GNDA.n1742 GNDA.n340 69.3109
R2805 GNDA.n407 GNDA.n340 69.3109
R2806 GNDA.n2155 GNDA.n2154 69.3109
R2807 GNDA.n2155 GNDA.n122 69.3109
R2808 GNDA.n743 GNDA.n636 69.3109
R2809 GNDA.n719 GNDA.n636 69.3109
R2810 GNDA.n1475 GNDA.n476 69.3109
R2811 GNDA.n1475 GNDA.n1474 69.3109
R2812 GNDA.n997 GNDA.n996 69.3109
R2813 GNDA.n996 GNDA.n995 69.3109
R2814 GNDA.n2113 GNDA.n2112 69.3109
R2815 GNDA.n2113 GNDA.n161 69.3109
R2816 GNDA.n1375 GNDA.n502 69.3109
R2817 GNDA.n1375 GNDA.n1374 69.3109
R2818 GNDA.t255 GNDA.t307 69.1104
R2819 GNDA.t199 GNDA.t123 69.1104
R2820 GNDA.t207 GNDA.n466 65.8183
R2821 GNDA.t207 GNDA.n465 65.8183
R2822 GNDA.t207 GNDA.n464 65.8183
R2823 GNDA.t207 GNDA.n463 65.8183
R2824 GNDA.t207 GNDA.n454 65.8183
R2825 GNDA.t207 GNDA.n461 65.8183
R2826 GNDA.t207 GNDA.n451 65.8183
R2827 GNDA.t207 GNDA.n462 65.8183
R2828 GNDA.t207 GNDA.n460 65.8183
R2829 GNDA.t207 GNDA.n459 65.8183
R2830 GNDA.t207 GNDA.n458 65.8183
R2831 GNDA.t207 GNDA.n457 65.8183
R2832 GNDA.t207 GNDA.n455 65.8183
R2833 GNDA.t207 GNDA.n453 65.8183
R2834 GNDA.t207 GNDA.n452 65.8183
R2835 GNDA.n1577 GNDA.t207 65.8183
R2836 GNDA.t239 GNDA.n897 65.8183
R2837 GNDA.t239 GNDA.n820 65.8183
R2838 GNDA.t239 GNDA.n819 65.8183
R2839 GNDA.t239 GNDA.n818 65.8183
R2840 GNDA.t239 GNDA.n809 65.8183
R2841 GNDA.t239 GNDA.n816 65.8183
R2842 GNDA.t239 GNDA.n807 65.8183
R2843 GNDA.t239 GNDA.n817 65.8183
R2844 GNDA.t239 GNDA.n815 65.8183
R2845 GNDA.t239 GNDA.n814 65.8183
R2846 GNDA.t239 GNDA.n813 65.8183
R2847 GNDA.t239 GNDA.n812 65.8183
R2848 GNDA.t239 GNDA.n810 65.8183
R2849 GNDA.t239 GNDA.n808 65.8183
R2850 GNDA.n898 GNDA.t239 65.8183
R2851 GNDA.t239 GNDA.n802 65.8183
R2852 GNDA.n391 GNDA.t240 65.8183
R2853 GNDA.n397 GNDA.t240 65.8183
R2854 GNDA.n399 GNDA.t240 65.8183
R2855 GNDA.n405 GNDA.t240 65.8183
R2856 GNDA.n375 GNDA.t240 65.8183
R2857 GNDA.n381 GNDA.t240 65.8183
R2858 GNDA.n383 GNDA.t240 65.8183
R2859 GNDA.n389 GNDA.t240 65.8183
R2860 GNDA.n359 GNDA.t240 65.8183
R2861 GNDA.n355 GNDA.t240 65.8183
R2862 GNDA.n366 GNDA.t240 65.8183
R2863 GNDA.n352 GNDA.t240 65.8183
R2864 GNDA.n356 GNDA.t240 65.8183
R2865 GNDA.n1759 GNDA.t240 65.8183
R2866 GNDA.n1756 GNDA.t240 65.8183
R2867 GNDA.n1743 GNDA.t240 65.8183
R2868 GNDA.t212 GNDA.n121 65.8183
R2869 GNDA.t212 GNDA.n120 65.8183
R2870 GNDA.t212 GNDA.n119 65.8183
R2871 GNDA.t212 GNDA.n118 65.8183
R2872 GNDA.t212 GNDA.n109 65.8183
R2873 GNDA.t212 GNDA.n116 65.8183
R2874 GNDA.t212 GNDA.n107 65.8183
R2875 GNDA.t212 GNDA.n117 65.8183
R2876 GNDA.t212 GNDA.n115 65.8183
R2877 GNDA.t212 GNDA.n114 65.8183
R2878 GNDA.t212 GNDA.n113 65.8183
R2879 GNDA.t212 GNDA.n112 65.8183
R2880 GNDA.t212 GNDA.n110 65.8183
R2881 GNDA.n2156 GNDA.t212 65.8183
R2882 GNDA.t212 GNDA.n108 65.8183
R2883 GNDA.t212 GNDA.n106 65.8183
R2884 GNDA.t208 GNDA.n733 65.8183
R2885 GNDA.t208 GNDA.n655 65.8183
R2886 GNDA.t208 GNDA.n654 65.8183
R2887 GNDA.t208 GNDA.n653 65.8183
R2888 GNDA.t208 GNDA.n644 65.8183
R2889 GNDA.t208 GNDA.n651 65.8183
R2890 GNDA.t208 GNDA.n642 65.8183
R2891 GNDA.t208 GNDA.n652 65.8183
R2892 GNDA.t208 GNDA.n650 65.8183
R2893 GNDA.t208 GNDA.n649 65.8183
R2894 GNDA.t208 GNDA.n648 65.8183
R2895 GNDA.t208 GNDA.n647 65.8183
R2896 GNDA.t208 GNDA.n645 65.8183
R2897 GNDA.t208 GNDA.n643 65.8183
R2898 GNDA.n734 GNDA.t208 65.8183
R2899 GNDA.t208 GNDA.n637 65.8183
R2900 GNDA.t192 GNDA.n493 65.8183
R2901 GNDA.t192 GNDA.n492 65.8183
R2902 GNDA.t192 GNDA.n491 65.8183
R2903 GNDA.t192 GNDA.n490 65.8183
R2904 GNDA.t192 GNDA.n481 65.8183
R2905 GNDA.t192 GNDA.n488 65.8183
R2906 GNDA.t192 GNDA.n478 65.8183
R2907 GNDA.t192 GNDA.n489 65.8183
R2908 GNDA.t192 GNDA.n487 65.8183
R2909 GNDA.t192 GNDA.n486 65.8183
R2910 GNDA.t192 GNDA.n485 65.8183
R2911 GNDA.t192 GNDA.n484 65.8183
R2912 GNDA.t192 GNDA.n482 65.8183
R2913 GNDA.t192 GNDA.n480 65.8183
R2914 GNDA.t192 GNDA.n479 65.8183
R2915 GNDA.n1476 GNDA.t192 65.8183
R2916 GNDA.n977 GNDA.t190 65.8183
R2917 GNDA.n979 GNDA.t190 65.8183
R2918 GNDA.n985 GNDA.t190 65.8183
R2919 GNDA.n987 GNDA.t190 65.8183
R2920 GNDA.n961 GNDA.t190 65.8183
R2921 GNDA.n963 GNDA.t190 65.8183
R2922 GNDA.n969 GNDA.t190 65.8183
R2923 GNDA.n971 GNDA.t190 65.8183
R2924 GNDA.t190 GNDA.n918 65.8183
R2925 GNDA.n946 GNDA.t190 65.8183
R2926 GNDA.n942 GNDA.t190 65.8183
R2927 GNDA.n953 GNDA.t190 65.8183
R2928 GNDA.n1026 GNDA.t190 65.8183
R2929 GNDA.n1013 GNDA.t190 65.8183
R2930 GNDA.n1011 GNDA.t190 65.8183
R2931 GNDA.n998 GNDA.t190 65.8183
R2932 GNDA.t253 GNDA.n160 65.8183
R2933 GNDA.t253 GNDA.n159 65.8183
R2934 GNDA.t253 GNDA.n158 65.8183
R2935 GNDA.t253 GNDA.n157 65.8183
R2936 GNDA.t253 GNDA.n148 65.8183
R2937 GNDA.t253 GNDA.n155 65.8183
R2938 GNDA.t253 GNDA.n146 65.8183
R2939 GNDA.t253 GNDA.n156 65.8183
R2940 GNDA.t253 GNDA.n154 65.8183
R2941 GNDA.t253 GNDA.n153 65.8183
R2942 GNDA.t253 GNDA.n152 65.8183
R2943 GNDA.t253 GNDA.n151 65.8183
R2944 GNDA.t253 GNDA.n149 65.8183
R2945 GNDA.n2114 GNDA.t253 65.8183
R2946 GNDA.t253 GNDA.n147 65.8183
R2947 GNDA.t253 GNDA.n145 65.8183
R2948 GNDA.t216 GNDA.n519 65.8183
R2949 GNDA.t216 GNDA.n518 65.8183
R2950 GNDA.t216 GNDA.n517 65.8183
R2951 GNDA.t216 GNDA.n516 65.8183
R2952 GNDA.t216 GNDA.n507 65.8183
R2953 GNDA.t216 GNDA.n514 65.8183
R2954 GNDA.t216 GNDA.n504 65.8183
R2955 GNDA.t216 GNDA.n515 65.8183
R2956 GNDA.t216 GNDA.n513 65.8183
R2957 GNDA.t216 GNDA.n512 65.8183
R2958 GNDA.t216 GNDA.n511 65.8183
R2959 GNDA.t216 GNDA.n510 65.8183
R2960 GNDA.t216 GNDA.n508 65.8183
R2961 GNDA.t216 GNDA.n506 65.8183
R2962 GNDA.t216 GNDA.n505 65.8183
R2963 GNDA.n1376 GNDA.t216 65.8183
R2964 GNDA.t210 GNDA.t288 65.7614
R2965 GNDA.t2 GNDA.t74 65.7614
R2966 GNDA.t74 GNDA.t31 65.7614
R2967 GNDA.t58 GNDA.t16 65.7614
R2968 GNDA.t133 GNDA.t58 65.7614
R2969 GNDA.t96 GNDA.t40 65.7614
R2970 GNDA.t40 GNDA.t23 65.7614
R2971 GNDA.t23 GNDA.t145 65.7614
R2972 GNDA.t194 GNDA.t83 65.7614
R2973 GNDA.n2254 GNDA.t255 65.271
R2974 GNDA.t138 GNDA.t97 65.271
R2975 GNDA.n2388 GNDA.t54 65.271
R2976 GNDA.n2459 GNDA.t22 65.271
R2977 GNDA.t68 GNDA.t102 65.271
R2978 GNDA.n2600 GNDA.t199 65.271
R2979 GNDA.t191 GNDA.n231 65.0078
R2980 GNDA.n1737 GNDA.t164 63.8432
R2981 GNDA.n2149 GNDA.t186 63.8432
R2982 GNDA.n2106 GNDA.t180 63.8432
R2983 GNDA.n2302 GNDA.t242 61.4316
R2984 GNDA.n2612 GNDA.t228 61.4316
R2985 GNDA.t21 GNDA.n2407 59.7836
R2986 GNDA.t126 GNDA.n2406 59.7836
R2987 GNDA.t73 GNDA.n2405 59.7836
R2988 GNDA.t20 GNDA.n2404 59.7836
R2989 GNDA.n2636 GNDA.t48 59.7836
R2990 GNDA.n2635 GNDA.t29 59.7836
R2991 GNDA.n35 GNDA.t64 59.7836
R2992 GNDA.n2637 GNDA.t24 59.7836
R2993 GNDA.t87 GNDA.n2408 59.7836
R2994 GNDA.n1764 GNDA.t166 59.7243
R2995 GNDA.n1856 GNDA.t188 59.7243
R2996 GNDA.n185 GNDA.t178 59.7243
R2997 GNDA.t39 GNDA.n1736 58.6946
R2998 GNDA.t14 GNDA.n1750 58.6946
R2999 GNDA.t125 GNDA.n1765 58.6946
R3000 GNDA.t207 GNDA.n1576 57.8461
R3001 GNDA.t239 GNDA.n801 57.8461
R3002 GNDA.n340 GNDA.t240 57.8461
R3003 GNDA.t212 GNDA.n2155 57.8461
R3004 GNDA.t208 GNDA.n636 57.8461
R3005 GNDA.t192 GNDA.n1475 57.8461
R3006 GNDA.n996 GNDA.t190 57.8461
R3007 GNDA.t253 GNDA.n2113 57.8461
R3008 GNDA.t216 GNDA.n1375 57.8461
R3009 GNDA.n2213 GNDA.t66 57.5921
R3010 GNDA.t49 GNDA.t94 57.5921
R3011 GNDA.n2403 GNDA.t54 57.5921
R3012 GNDA.t22 GNDA.n33 57.5921
R3013 GNDA.n2642 GNDA.t93 57.5921
R3014 GNDA.t36 GNDA.t63 57.5921
R3015 GNDA.t81 GNDA.n2628 57.5921
R3016 GNDA.t154 GNDA.t4 56.6352
R3017 GNDA.n2136 GNDA.t273 56.6352
R3018 GNDA.t90 GNDA.t150 56.6352
R3019 GNDA.n1588 GNDA.n416 56.3995
R3020 GNDA.n1586 GNDA.n416 56.3995
R3021 GNDA.n1036 GNDA.n626 56.3995
R3022 GNDA.n2020 GNDA.n2019 56.3995
R3023 GNDA.n2021 GNDA.n2020 56.3995
R3024 GNDA.n1036 GNDA.n1035 56.3995
R3025 GNDA.n1289 GNDA.n1288 56.3995
R3026 GNDA.n1290 GNDA.n1289 56.3995
R3027 GNDA.n1732 GNDA.n410 56.3995
R3028 GNDA.n796 GNDA.n423 56.3995
R3029 GNDA.n1930 GNDA.n1929 55.6055
R3030 GNDA.t207 GNDA.n456 55.2026
R3031 GNDA.t239 GNDA.n811 55.2026
R3032 GNDA.n373 GNDA.t240 55.2026
R3033 GNDA.t212 GNDA.n111 55.2026
R3034 GNDA.t208 GNDA.n646 55.2026
R3035 GNDA.t192 GNDA.n483 55.2026
R3036 GNDA.n955 GNDA.t190 55.2026
R3037 GNDA.t253 GNDA.n150 55.2026
R3038 GNDA.t216 GNDA.n509 55.2026
R3039 GNDA.n1848 GNDA.n128 54.5757
R3040 GNDA.n1939 GNDA.n1938 54.5757
R3041 GNDA.t313 GNDA.n2107 54.5757
R3042 GNDA.n178 GNDA.t35 54.5757
R3043 GNDA.t286 GNDA.n2032 54.5757
R3044 GNDA.t172 GNDA.n1856 53.546
R3045 GNDA.n1556 GNDA.n462 53.3664
R3046 GNDA.n1552 GNDA.n451 53.3664
R3047 GNDA.n1548 GNDA.n461 53.3664
R3048 GNDA.n1544 GNDA.n454 53.3664
R3049 GNDA.n1533 GNDA.n457 53.3664
R3050 GNDA.n1529 GNDA.n458 53.3664
R3051 GNDA.n1525 GNDA.n459 53.3664
R3052 GNDA.n1521 GNDA.n460 53.3664
R3053 GNDA.n1578 GNDA.n1577 53.3664
R3054 GNDA.n1498 GNDA.n452 53.3664
R3055 GNDA.n1506 GNDA.n453 53.3664
R3056 GNDA.n1513 GNDA.n455 53.3664
R3057 GNDA.n1560 GNDA.n466 53.3664
R3058 GNDA.n1561 GNDA.n465 53.3664
R3059 GNDA.n1565 GNDA.n464 53.3664
R3060 GNDA.n1569 GNDA.n463 53.3664
R3061 GNDA.n1557 GNDA.n466 53.3664
R3062 GNDA.n1564 GNDA.n465 53.3664
R3063 GNDA.n1568 GNDA.n464 53.3664
R3064 GNDA.n467 GNDA.n463 53.3664
R3065 GNDA.n1541 GNDA.n454 53.3664
R3066 GNDA.n1545 GNDA.n461 53.3664
R3067 GNDA.n1549 GNDA.n451 53.3664
R3068 GNDA.n1553 GNDA.n462 53.3664
R3069 GNDA.n1524 GNDA.n460 53.3664
R3070 GNDA.n1528 GNDA.n459 53.3664
R3071 GNDA.n1532 GNDA.n458 53.3664
R3072 GNDA.n1536 GNDA.n457 53.3664
R3073 GNDA.n1520 GNDA.n455 53.3664
R3074 GNDA.n1512 GNDA.n453 53.3664
R3075 GNDA.n1505 GNDA.n452 53.3664
R3076 GNDA.n1577 GNDA.n450 53.3664
R3077 GNDA.n880 GNDA.n817 53.3664
R3078 GNDA.n877 GNDA.n807 53.3664
R3079 GNDA.n873 GNDA.n816 53.3664
R3080 GNDA.n869 GNDA.n809 53.3664
R3081 GNDA.n858 GNDA.n812 53.3664
R3082 GNDA.n854 GNDA.n813 53.3664
R3083 GNDA.n850 GNDA.n814 53.3664
R3084 GNDA.n846 GNDA.n815 53.3664
R3085 GNDA.n906 GNDA.n802 53.3664
R3086 GNDA.n899 GNDA.n898 53.3664
R3087 GNDA.n831 GNDA.n808 53.3664
R3088 GNDA.n838 GNDA.n810 53.3664
R3089 GNDA.n897 GNDA.n896 53.3664
R3090 GNDA.n822 GNDA.n820 53.3664
R3091 GNDA.n891 GNDA.n819 53.3664
R3092 GNDA.n887 GNDA.n818 53.3664
R3093 GNDA.n897 GNDA.n821 53.3664
R3094 GNDA.n892 GNDA.n820 53.3664
R3095 GNDA.n888 GNDA.n819 53.3664
R3096 GNDA.n884 GNDA.n818 53.3664
R3097 GNDA.n866 GNDA.n809 53.3664
R3098 GNDA.n870 GNDA.n816 53.3664
R3099 GNDA.n874 GNDA.n807 53.3664
R3100 GNDA.n878 GNDA.n817 53.3664
R3101 GNDA.n849 GNDA.n815 53.3664
R3102 GNDA.n853 GNDA.n814 53.3664
R3103 GNDA.n857 GNDA.n813 53.3664
R3104 GNDA.n861 GNDA.n812 53.3664
R3105 GNDA.n845 GNDA.n810 53.3664
R3106 GNDA.n837 GNDA.n808 53.3664
R3107 GNDA.n898 GNDA.n806 53.3664
R3108 GNDA.n805 GNDA.n802 53.3664
R3109 GNDA.n390 GNDA.n389 53.3664
R3110 GNDA.n383 GNDA.n346 53.3664
R3111 GNDA.n382 GNDA.n381 53.3664
R3112 GNDA.n375 GNDA.n348 53.3664
R3113 GNDA.n368 GNDA.n352 53.3664
R3114 GNDA.n366 GNDA.n365 53.3664
R3115 GNDA.n361 GNDA.n355 53.3664
R3116 GNDA.n359 GNDA.n358 53.3664
R3117 GNDA.n1744 GNDA.n1743 53.3664
R3118 GNDA.n1756 GNDA.n1755 53.3664
R3119 GNDA.n1759 GNDA.n1758 53.3664
R3120 GNDA.n356 GNDA.n332 53.3664
R3121 GNDA.n391 GNDA.n344 53.3664
R3122 GNDA.n397 GNDA.n396 53.3664
R3123 GNDA.n400 GNDA.n399 53.3664
R3124 GNDA.n405 GNDA.n404 53.3664
R3125 GNDA.n392 GNDA.n391 53.3664
R3126 GNDA.n398 GNDA.n397 53.3664
R3127 GNDA.n399 GNDA.n342 53.3664
R3128 GNDA.n406 GNDA.n405 53.3664
R3129 GNDA.n376 GNDA.n375 53.3664
R3130 GNDA.n381 GNDA.n380 53.3664
R3131 GNDA.n384 GNDA.n383 53.3664
R3132 GNDA.n389 GNDA.n388 53.3664
R3133 GNDA.n360 GNDA.n359 53.3664
R3134 GNDA.n355 GNDA.n353 53.3664
R3135 GNDA.n367 GNDA.n366 53.3664
R3136 GNDA.n352 GNDA.n350 53.3664
R3137 GNDA.n357 GNDA.n356 53.3664
R3138 GNDA.n1760 GNDA.n1759 53.3664
R3139 GNDA.n1757 GNDA.n1756 53.3664
R3140 GNDA.n1743 GNDA.n335 53.3664
R3141 GNDA.n1898 GNDA.n117 53.3664
R3142 GNDA.n1894 GNDA.n107 53.3664
R3143 GNDA.n1890 GNDA.n116 53.3664
R3144 GNDA.n1886 GNDA.n109 53.3664
R3145 GNDA.n1875 GNDA.n112 53.3664
R3146 GNDA.n1871 GNDA.n113 53.3664
R3147 GNDA.n1867 GNDA.n114 53.3664
R3148 GNDA.n1863 GNDA.n115 53.3664
R3149 GNDA.n123 GNDA.n106 53.3664
R3150 GNDA.n2144 GNDA.n108 53.3664
R3151 GNDA.n2157 GNDA.n2156 53.3664
R3152 GNDA.n1852 GNDA.n110 53.3664
R3153 GNDA.n1902 GNDA.n121 53.3664
R3154 GNDA.n1903 GNDA.n120 53.3664
R3155 GNDA.n1907 GNDA.n119 53.3664
R3156 GNDA.n1911 GNDA.n118 53.3664
R3157 GNDA.n1899 GNDA.n121 53.3664
R3158 GNDA.n1906 GNDA.n120 53.3664
R3159 GNDA.n1910 GNDA.n119 53.3664
R3160 GNDA.n1913 GNDA.n118 53.3664
R3161 GNDA.n1883 GNDA.n109 53.3664
R3162 GNDA.n1887 GNDA.n116 53.3664
R3163 GNDA.n1891 GNDA.n107 53.3664
R3164 GNDA.n1895 GNDA.n117 53.3664
R3165 GNDA.n1866 GNDA.n115 53.3664
R3166 GNDA.n1870 GNDA.n114 53.3664
R3167 GNDA.n1874 GNDA.n113 53.3664
R3168 GNDA.n1878 GNDA.n112 53.3664
R3169 GNDA.n1862 GNDA.n110 53.3664
R3170 GNDA.n2156 GNDA.n105 53.3664
R3171 GNDA.n108 GNDA.n104 53.3664
R3172 GNDA.n2143 GNDA.n106 53.3664
R3173 GNDA.n715 GNDA.n652 53.3664
R3174 GNDA.n712 GNDA.n642 53.3664
R3175 GNDA.n708 GNDA.n651 53.3664
R3176 GNDA.n704 GNDA.n644 53.3664
R3177 GNDA.n693 GNDA.n647 53.3664
R3178 GNDA.n689 GNDA.n648 53.3664
R3179 GNDA.n685 GNDA.n649 53.3664
R3180 GNDA.n681 GNDA.n650 53.3664
R3181 GNDA.n742 GNDA.n637 53.3664
R3182 GNDA.n735 GNDA.n734 53.3664
R3183 GNDA.n666 GNDA.n643 53.3664
R3184 GNDA.n673 GNDA.n645 53.3664
R3185 GNDA.n733 GNDA.n732 53.3664
R3186 GNDA.n657 GNDA.n655 53.3664
R3187 GNDA.n727 GNDA.n654 53.3664
R3188 GNDA.n723 GNDA.n653 53.3664
R3189 GNDA.n733 GNDA.n656 53.3664
R3190 GNDA.n728 GNDA.n655 53.3664
R3191 GNDA.n724 GNDA.n654 53.3664
R3192 GNDA.n720 GNDA.n653 53.3664
R3193 GNDA.n701 GNDA.n644 53.3664
R3194 GNDA.n705 GNDA.n651 53.3664
R3195 GNDA.n709 GNDA.n642 53.3664
R3196 GNDA.n713 GNDA.n652 53.3664
R3197 GNDA.n684 GNDA.n650 53.3664
R3198 GNDA.n688 GNDA.n649 53.3664
R3199 GNDA.n692 GNDA.n648 53.3664
R3200 GNDA.n696 GNDA.n647 53.3664
R3201 GNDA.n680 GNDA.n645 53.3664
R3202 GNDA.n672 GNDA.n643 53.3664
R3203 GNDA.n734 GNDA.n641 53.3664
R3204 GNDA.n640 GNDA.n637 53.3664
R3205 GNDA.n1457 GNDA.n489 53.3664
R3206 GNDA.n1453 GNDA.n478 53.3664
R3207 GNDA.n1449 GNDA.n488 53.3664
R3208 GNDA.n1445 GNDA.n481 53.3664
R3209 GNDA.n1434 GNDA.n484 53.3664
R3210 GNDA.n1430 GNDA.n485 53.3664
R3211 GNDA.n1426 GNDA.n486 53.3664
R3212 GNDA.n1422 GNDA.n487 53.3664
R3213 GNDA.n1477 GNDA.n1476 53.3664
R3214 GNDA.n1399 GNDA.n479 53.3664
R3215 GNDA.n1407 GNDA.n480 53.3664
R3216 GNDA.n1414 GNDA.n482 53.3664
R3217 GNDA.n1461 GNDA.n493 53.3664
R3218 GNDA.n1462 GNDA.n492 53.3664
R3219 GNDA.n1466 GNDA.n491 53.3664
R3220 GNDA.n1470 GNDA.n490 53.3664
R3221 GNDA.n1458 GNDA.n493 53.3664
R3222 GNDA.n1465 GNDA.n492 53.3664
R3223 GNDA.n1469 GNDA.n491 53.3664
R3224 GNDA.n1473 GNDA.n490 53.3664
R3225 GNDA.n1442 GNDA.n481 53.3664
R3226 GNDA.n1446 GNDA.n488 53.3664
R3227 GNDA.n1450 GNDA.n478 53.3664
R3228 GNDA.n1454 GNDA.n489 53.3664
R3229 GNDA.n1425 GNDA.n487 53.3664
R3230 GNDA.n1429 GNDA.n486 53.3664
R3231 GNDA.n1433 GNDA.n485 53.3664
R3232 GNDA.n1437 GNDA.n484 53.3664
R3233 GNDA.n1421 GNDA.n482 53.3664
R3234 GNDA.n1413 GNDA.n480 53.3664
R3235 GNDA.n1406 GNDA.n479 53.3664
R3236 GNDA.n1476 GNDA.n477 53.3664
R3237 GNDA.n971 GNDA.n934 53.3664
R3238 GNDA.n970 GNDA.n969 53.3664
R3239 GNDA.n963 GNDA.n936 53.3664
R3240 GNDA.n962 GNDA.n961 53.3664
R3241 GNDA.n953 GNDA.n952 53.3664
R3242 GNDA.n948 GNDA.n942 53.3664
R3243 GNDA.n946 GNDA.n945 53.3664
R3244 GNDA.n1028 GNDA.n918 53.3664
R3245 GNDA.n999 GNDA.n998 53.3664
R3246 GNDA.n1011 GNDA.n1010 53.3664
R3247 GNDA.n1014 GNDA.n1013 53.3664
R3248 GNDA.n1026 GNDA.n1025 53.3664
R3249 GNDA.n978 GNDA.n977 53.3664
R3250 GNDA.n980 GNDA.n979 53.3664
R3251 GNDA.n985 GNDA.n984 53.3664
R3252 GNDA.n988 GNDA.n987 53.3664
R3253 GNDA.n977 GNDA.n976 53.3664
R3254 GNDA.n979 GNDA.n932 53.3664
R3255 GNDA.n986 GNDA.n985 53.3664
R3256 GNDA.n987 GNDA.n930 53.3664
R3257 GNDA.n961 GNDA.n960 53.3664
R3258 GNDA.n964 GNDA.n963 53.3664
R3259 GNDA.n969 GNDA.n968 53.3664
R3260 GNDA.n972 GNDA.n971 53.3664
R3261 GNDA.n943 GNDA.n918 53.3664
R3262 GNDA.n947 GNDA.n946 53.3664
R3263 GNDA.n942 GNDA.n940 53.3664
R3264 GNDA.n954 GNDA.n953 53.3664
R3265 GNDA.n1027 GNDA.n1026 53.3664
R3266 GNDA.n1013 GNDA.n919 53.3664
R3267 GNDA.n1012 GNDA.n1011 53.3664
R3268 GNDA.n998 GNDA.n924 53.3664
R3269 GNDA.n2073 GNDA.n156 53.3664
R3270 GNDA.n2069 GNDA.n146 53.3664
R3271 GNDA.n2065 GNDA.n155 53.3664
R3272 GNDA.n2061 GNDA.n148 53.3664
R3273 GNDA.n2050 GNDA.n151 53.3664
R3274 GNDA.n2046 GNDA.n152 53.3664
R3275 GNDA.n2042 GNDA.n153 53.3664
R3276 GNDA.n2038 GNDA.n154 53.3664
R3277 GNDA.n162 GNDA.n145 53.3664
R3278 GNDA.n2102 GNDA.n147 53.3664
R3279 GNDA.n2115 GNDA.n2114 53.3664
R3280 GNDA.n180 GNDA.n149 53.3664
R3281 GNDA.n2077 GNDA.n160 53.3664
R3282 GNDA.n2078 GNDA.n159 53.3664
R3283 GNDA.n2082 GNDA.n158 53.3664
R3284 GNDA.n2086 GNDA.n157 53.3664
R3285 GNDA.n2074 GNDA.n160 53.3664
R3286 GNDA.n2081 GNDA.n159 53.3664
R3287 GNDA.n2085 GNDA.n158 53.3664
R3288 GNDA.n2088 GNDA.n157 53.3664
R3289 GNDA.n2058 GNDA.n148 53.3664
R3290 GNDA.n2062 GNDA.n155 53.3664
R3291 GNDA.n2066 GNDA.n146 53.3664
R3292 GNDA.n2070 GNDA.n156 53.3664
R3293 GNDA.n2041 GNDA.n154 53.3664
R3294 GNDA.n2045 GNDA.n153 53.3664
R3295 GNDA.n2049 GNDA.n152 53.3664
R3296 GNDA.n2053 GNDA.n151 53.3664
R3297 GNDA.n2037 GNDA.n149 53.3664
R3298 GNDA.n2114 GNDA.n144 53.3664
R3299 GNDA.n147 GNDA.n143 53.3664
R3300 GNDA.n2101 GNDA.n145 53.3664
R3301 GNDA.n1357 GNDA.n515 53.3664
R3302 GNDA.n1353 GNDA.n504 53.3664
R3303 GNDA.n1349 GNDA.n514 53.3664
R3304 GNDA.n1345 GNDA.n507 53.3664
R3305 GNDA.n1334 GNDA.n510 53.3664
R3306 GNDA.n1330 GNDA.n511 53.3664
R3307 GNDA.n1326 GNDA.n512 53.3664
R3308 GNDA.n1322 GNDA.n513 53.3664
R3309 GNDA.n1377 GNDA.n1376 53.3664
R3310 GNDA.n1299 GNDA.n505 53.3664
R3311 GNDA.n1307 GNDA.n506 53.3664
R3312 GNDA.n1314 GNDA.n508 53.3664
R3313 GNDA.n1361 GNDA.n519 53.3664
R3314 GNDA.n1362 GNDA.n518 53.3664
R3315 GNDA.n1366 GNDA.n517 53.3664
R3316 GNDA.n1370 GNDA.n516 53.3664
R3317 GNDA.n1358 GNDA.n519 53.3664
R3318 GNDA.n1365 GNDA.n518 53.3664
R3319 GNDA.n1369 GNDA.n517 53.3664
R3320 GNDA.n1373 GNDA.n516 53.3664
R3321 GNDA.n1342 GNDA.n507 53.3664
R3322 GNDA.n1346 GNDA.n514 53.3664
R3323 GNDA.n1350 GNDA.n504 53.3664
R3324 GNDA.n1354 GNDA.n515 53.3664
R3325 GNDA.n1325 GNDA.n513 53.3664
R3326 GNDA.n1329 GNDA.n512 53.3664
R3327 GNDA.n1333 GNDA.n511 53.3664
R3328 GNDA.n1337 GNDA.n510 53.3664
R3329 GNDA.n1321 GNDA.n508 53.3664
R3330 GNDA.n1313 GNDA.n506 53.3664
R3331 GNDA.n1306 GNDA.n505 53.3664
R3332 GNDA.n1376 GNDA.n503 53.3664
R3333 GNDA.n1268 GNDA.n1067 52.7091
R3334 GNDA.n1269 GNDA.n1268 52.7091
R3335 GNDA.n1271 GNDA.n1269 52.7091
R3336 GNDA.n1271 GNDA.n1270 52.7091
R3337 GNDA.n1270 GNDA.n235 52.7091
R3338 GNDA.n1278 GNDA.n234 52.7091
R3339 GNDA.n1278 GNDA.n1061 52.7091
R3340 GNDA.n1285 GNDA.n1061 52.7091
R3341 GNDA.n1286 GNDA.n1285 52.7091
R3342 GNDA.n1287 GNDA.n1286 52.7091
R3343 GNDA.n1287 GNDA.n1059 52.7091
R3344 GNDA.n1059 GNDA.t124 52.7091
R3345 GNDA.n1058 GNDA.n521 52.7091
R3346 GNDA.n1052 GNDA.n521 52.7091
R3347 GNDA.n1052 GNDA.n1051 52.7091
R3348 GNDA.n1051 GNDA.n1050 52.7091
R3349 GNDA.n1050 GNDA.n233 52.7091
R3350 GNDA.n1043 GNDA.n232 52.7091
R3351 GNDA.n1043 GNDA.n1042 52.7091
R3352 GNDA.n1042 GNDA.n1041 52.7091
R3353 GNDA.n1041 GNDA.n621 52.7091
R3354 GNDA.n625 GNDA.n621 52.7091
R3355 GNDA.n625 GNDA.n231 52.7091
R3356 GNDA.n1997 GNDA.n199 52.7091
R3357 GNDA.n2004 GNDA.n199 52.7091
R3358 GNDA.n2005 GNDA.n2004 52.7091
R3359 GNDA.n2006 GNDA.n2005 52.7091
R3360 GNDA.n2006 GNDA.n138 52.7091
R3361 GNDA.n194 GNDA.n139 52.7091
R3362 GNDA.n2015 GNDA.n194 52.7091
R3363 GNDA.n2016 GNDA.n2015 52.7091
R3364 GNDA.n2017 GNDA.n2016 52.7091
R3365 GNDA.n2017 GNDA.n189 52.7091
R3366 GNDA.n2022 GNDA.n189 52.7091
R3367 GNDA.t191 GNDA.n1957 51.4866
R3368 GNDA.t191 GNDA.n306 51.4866
R3369 GNDA.n2410 GNDA.t2 50.8162
R3370 GNDA.t145 GNDA.n2633 50.8162
R3371 GNDA.n2443 GNDA.t115 50.8162
R3372 GNDA.t260 GNDA.t297 49.9132
R3373 GNDA.t306 GNDA.t205 49.9132
R3374 GNDA.t160 GNDA.n2149 49.4271
R3375 GNDA.n1938 GNDA.t27 48.3974
R3376 GNDA.t191 GNDA.n1996 47.6748
R3377 GNDA.n1929 GNDA.t3 47.3677
R3378 GNDA.t245 GNDA.t65 46.338
R3379 GNDA.t231 GNDA.t91 46.338
R3380 GNDA.n1160 GNDA.t191 46.2335
R3381 GNDA.n1184 GNDA.t191 46.2335
R3382 GNDA.t191 GNDA.n1252 46.2335
R3383 GNDA.t31 GNDA.n2409 44.838
R3384 GNDA.n2634 GNDA.t96 44.838
R3385 GNDA.n1738 GNDA.t245 43.2488
R3386 GNDA.n2150 GNDA.t160 43.2488
R3387 GNDA.n2107 GNDA.t176 43.2488
R3388 GNDA.t191 GNDA.n1146 42.2987
R3389 GNDA.n1192 GNDA.t191 42.2987
R3390 GNDA.n1253 GNDA.t191 42.2987
R3391 GNDA.t144 GNDA.t89 42.2405
R3392 GNDA.t298 GNDA.t144 42.2405
R3393 GNDA.t13 GNDA.t312 42.2405
R3394 GNDA.t290 GNDA.t13 42.2405
R3395 GNDA.t265 GNDA.t242 42.2344
R3396 GNDA.t228 GNDA.t282 42.2344
R3397 GNDA.n2138 GNDA.t100 42.2191
R3398 GNDA.t191 GNDA.t3 41.1894
R3399 GNDA.t191 GNDA.t27 41.1894
R3400 GNDA.n2410 GNDA.n2171 40.5993
R3401 GNDA.n2633 GNDA.n2632 40.5993
R3402 GNDA.n2134 GNDA.n129 39.3903
R3403 GNDA.n1765 GNDA.t156 39.1299
R3404 GNDA.n2162 GNDA.n2161 39.1299
R3405 GNDA.n1857 GNDA.t172 39.1299
R3406 GNDA.n2033 GNDA.t231 39.1299
R3407 GNDA.n1957 GNDA.n308 38.1002
R3408 GNDA.n1858 GNDA.n128 38.1002
R3409 GNDA.n2119 GNDA.t35 38.1002
R3410 GNDA.n2033 GNDA.t286 38.1002
R3411 GNDA.n1847 GNDA.n306 37.0705
R3412 GNDA.t191 GNDA.t182 36.0408
R3413 GNDA.t191 GNDA.t162 36.0408
R3414 GNDA.t191 GNDA.n235 35.7252
R3415 GNDA.t191 GNDA.n233 35.7252
R3416 GNDA.t191 GNDA.n138 35.7252
R3417 GNDA.n2133 GNDA.n2132 35.3278
R3418 GNDA.t307 GNDA.n2213 34.5555
R3419 GNDA.t80 GNDA.t260 34.5555
R3420 GNDA.t205 GNDA.t88 34.5555
R3421 GNDA.n2628 GNDA.t123 34.5555
R3422 GNDA.n1738 GNDA.t39 33.9813
R3423 GNDA.n1751 GNDA.t14 33.9813
R3424 GNDA.n2137 GNDA.n2136 33.9813
R3425 GNDA.n327 GNDA.t166 32.9516
R3426 GNDA.t188 GNDA.n1850 32.9516
R3427 GNDA.t178 GNDA.n184 32.9516
R3428 GNDA.t191 GNDA.n226 32.9056
R3429 GNDA.t191 GNDA.n225 32.9056
R3430 GNDA.n2026 GNDA.n2025 32.3063
R3431 GNDA.n2649 GNDA.n0 29.8047
R3432 GNDA.t294 GNDA.n171 29.2831
R3433 GNDA.n1749 GNDA.t164 28.8327
R3434 GNDA.t186 GNDA.n2148 28.8327
R3435 GNDA.t180 GNDA.n2096 28.8327
R3436 GNDA.t4 GNDA.n1749 27.803
R3437 GNDA.t289 GNDA.n1764 27.803
R3438 GNDA.n1768 GNDA.t33 27.803
R3439 GNDA.n1558 GNDA.n1555 27.5561
R3440 GNDA.n882 GNDA.n881 27.5561
R3441 GNDA.n393 GNDA.n345 27.5561
R3442 GNDA.n1900 GNDA.n1897 27.5561
R3443 GNDA.n717 GNDA.n716 27.5561
R3444 GNDA.n1459 GNDA.n1456 27.5561
R3445 GNDA.n975 GNDA.n974 27.5561
R3446 GNDA.n2075 GNDA.n2072 27.5561
R3447 GNDA.n1359 GNDA.n1356 27.5561
R3448 GNDA.t94 GNDA.t121 26.8766
R3449 GNDA.t5 GNDA.n2403 26.8766
R3450 GNDA.t110 GNDA.n33 26.8766
R3451 GNDA.t127 GNDA.t36 26.8766
R3452 GNDA.n1539 GNDA.n1538 26.6672
R3453 GNDA.n864 GNDA.n863 26.6672
R3454 GNDA.n371 GNDA.n349 26.6672
R3455 GNDA.n1881 GNDA.n1880 26.6672
R3456 GNDA.n699 GNDA.n698 26.6672
R3457 GNDA.n1440 GNDA.n1439 26.6672
R3458 GNDA.n958 GNDA.n957 26.6672
R3459 GNDA.n2056 GNDA.n2055 26.6672
R3460 GNDA.n1340 GNDA.n1339 26.6672
R3461 GNDA.t156 GNDA.t289 25.7435
R3462 GNDA.t176 GNDA.t28 25.7435
R3463 GNDA.n220 GNDA.n210 25.3679
R3464 GNDA.n2395 GNDA.n2394 24.991
R3465 GNDA.n2491 GNDA.n2490 24.991
R3466 GNDA.n2494 GNDA.n2493 24.991
R3467 GNDA.n2418 GNDA.n2417 24.991
R3468 GNDA.n2428 GNDA.n2427 24.991
R3469 GNDA.n2478 GNDA.n2477 24.991
R3470 GNDA.n2475 GNDA.n2474 24.991
R3471 GNDA.n2366 GNDA.n2365 24.7472
R3472 GNDA.n311 GNDA.t165 24.0005
R3473 GNDA.n311 GNDA.t155 24.0005
R3474 GNDA.n313 GNDA.t183 24.0005
R3475 GNDA.n313 GNDA.t167 24.0005
R3476 GNDA.n315 GNDA.t157 24.0005
R3477 GNDA.n315 GNDA.t185 24.0005
R3478 GNDA.n1952 GNDA.t171 24.0005
R3479 GNDA.n1952 GNDA.t161 24.0005
R3480 GNDA.n1950 GNDA.t187 24.0005
R3481 GNDA.n1950 GNDA.t169 24.0005
R3482 GNDA.n1948 GNDA.t159 24.0005
R3483 GNDA.n1948 GNDA.t189 24.0005
R3484 GNDA.n1946 GNDA.t173 24.0005
R3485 GNDA.n1946 GNDA.t175 24.0005
R3486 GNDA.n1936 GNDA.t153 24.0005
R3487 GNDA.n1936 GNDA.t177 24.0005
R3488 GNDA.n1934 GNDA.t181 24.0005
R3489 GNDA.n1934 GNDA.t163 24.0005
R3490 GNDA.n186 GNDA.t151 24.0005
R3491 GNDA.n186 GNDA.t179 24.0005
R3492 GNDA.n2094 GNDA.t104 23.6841
R3493 GNDA.t28 GNDA.n2106 23.6841
R3494 GNDA.n184 GNDA.t90 23.6841
R3495 GNDA.n2355 GNDA.n2354 22.8576
R3496 GNDA.n2321 GNDA.n2320 22.8576
R3497 GNDA.n2391 GNDA.n2390 22.8576
R3498 GNDA.n2449 GNDA.n2448 22.8576
R3499 GNDA.n2305 GNDA.n2304 22.8576
R3500 GNDA.n2203 GNDA.n2173 22.8576
R3501 GNDA.n2433 GNDA.n2432 22.8576
R3502 GNDA.n2384 GNDA.n73 22.8576
R3503 GNDA.n54 GNDA.n53 22.8576
R3504 GNDA.n2464 GNDA.n2463 22.8576
R3505 GNDA.n2615 GNDA.n2614 22.8576
R3506 GNDA.n2618 GNDA.n2617 22.8576
R3507 GNDA.n2574 GNDA.n2573 22.8576
R3508 GNDA.n2567 GNDA.n2566 22.8576
R3509 GNDA.n2264 GNDA.n2263 22.8576
R3510 GNDA.n2257 GNDA.n2256 22.8576
R3511 GNDA.t170 GNDA.n2137 22.6544
R3512 GNDA.n2108 GNDA.t152 22.6544
R3513 GNDA.n2493 GNDA.n2492 21.6651
R3514 GNDA.t294 GNDA.n167 21.084
R3515 GNDA.n1093 GNDA.n1092 21.0192
R3516 GNDA.n2409 GNDA.t87 20.9249
R3517 GNDA.t29 GNDA.n2634 20.9249
R3518 GNDA.n310 GNDA.n309 20.8233
R3519 GNDA.n1932 GNDA.n1931 20.8233
R3520 GNDA.n1956 GNDA.n1955 20.8233
R3521 GNDA.n1944 GNDA.n1943 20.8233
R3522 GNDA.n1941 GNDA.n1940 20.8233
R3523 GNDA.n2030 GNDA.n2029 20.8233
R3524 GNDA.n61 GNDA.n1 20.7243
R3525 GNDA.n2645 GNDA.n2644 20.7243
R3526 GNDA.t191 GNDA.n223 20.5949
R3527 GNDA.t38 GNDA.n223 20.5949
R3528 GNDA.n1930 GNDA.t33 20.5949
R3529 GNDA.n1939 GNDA.t104 20.5949
R3530 GNDA.n2130 GNDA.t149 20.5949
R3531 GNDA.n2130 GNDA.t191 20.5949
R3532 GNDA.t191 GNDA.n207 19.9378
R3533 GNDA.n83 GNDA.t141 19.7005
R3534 GNDA.n83 GNDA.t60 19.7005
R3535 GNDA.n81 GNDA.t309 19.7005
R3536 GNDA.n81 GNDA.t107 19.7005
R3537 GNDA.n79 GNDA.t310 19.7005
R3538 GNDA.n79 GNDA.t84 19.7005
R3539 GNDA.n77 GNDA.t305 19.7005
R3540 GNDA.n77 GNDA.t140 19.7005
R3541 GNDA.n75 GNDA.t304 19.7005
R3542 GNDA.n75 GNDA.t118 19.7005
R3543 GNDA.n74 GNDA.t9 19.7005
R3544 GNDA.n74 GNDA.t296 19.7005
R3545 GNDA.n26 GNDA.t11 19.7005
R3546 GNDA.n26 GNDA.t82 19.7005
R3547 GNDA.n24 GNDA.t128 19.7005
R3548 GNDA.n24 GNDA.t86 19.7005
R3549 GNDA.n22 GNDA.t101 19.7005
R3550 GNDA.n22 GNDA.t42 19.7005
R3551 GNDA.n20 GNDA.t120 19.7005
R3552 GNDA.n20 GNDA.t62 19.7005
R3553 GNDA.n18 GNDA.t311 19.7005
R3554 GNDA.n18 GNDA.t303 19.7005
R3555 GNDA.n17 GNDA.t51 19.7005
R3556 GNDA.n17 GNDA.t137 19.7005
R3557 GNDA.t191 GNDA.n227 19.6741
R3558 GNDA.n2254 GNDA.t61 19.1977
R3559 GNDA.t85 GNDA.t138 19.1977
R3560 GNDA.n2388 GNDA.t131 19.1977
R3561 GNDA.n2459 GNDA.t56 19.1977
R3562 GNDA.n2642 GNDA.t7 19.1977
R3563 GNDA.t102 GNDA.t119 19.1977
R3564 GNDA.t293 GNDA.n2600 19.1977
R3565 GNDA.n2649 GNDA.n2648 19.008
R3566 GNDA.n1189 GNDA.n1097 18.5605
R3567 GNDA.n1766 GNDA.t184 18.5355
R3568 GNDA.n1858 GNDA.t174 18.5355
R3569 GNDA GNDA.n131 18.1546
R3570 GNDA.n2306 GNDA.n2173 18.1442
R3571 GNDA.n2617 GNDA.n2616 18.1442
R3572 GNDA.n2476 GNDA.n2475 18.0401
R3573 GNDA.n1056 GNDA.n615 17.5843
R3574 GNDA.n1999 GNDA.n201 17.5843
R3575 GNDA.n1265 GNDA.n1264 17.5843
R3576 GNDA.t191 GNDA.n206 17.5058
R3577 GNDA.n2031 GNDA.n167 17.5058
R3578 GNDA.n2367 GNDA.n2366 17.4151
R3579 GNDA.n2394 GNDA.n2393 17.4151
R3580 GNDA.n2492 GNDA.n2491 17.4151
R3581 GNDA.t191 GNDA.n234 16.9844
R3582 GNDA.t191 GNDA.n232 16.9844
R3583 GNDA.t191 GNDA.n139 16.9844
R3584 GNDA.n1607 GNDA.n427 16.9379
R3585 GNDA.n775 GNDA.n772 16.9379
R3586 GNDA.n1710 GNDA.n1709 16.9379
R3587 GNDA.n524 GNDA.n495 16.7709
R3588 GNDA.n1964 GNDA.n1963 16.7709
R3589 GNDA.n1688 GNDA.n290 16.7709
R3590 GNDA.n1992 GNDA.n261 16.7709
R3591 GNDA.n28 GNDA.n27 16.5057
R3592 GNDA.n2360 GNDA.t211 16.0005
R3593 GNDA.n2398 GNDA.t219 16.0005
R3594 GNDA.n2485 GNDA.t271 16.0005
R3595 GNDA.n2497 GNDA.t280 16.0005
R3596 GNDA.n2411 GNDA.t215 16.0005
R3597 GNDA.n2422 GNDA.t234 16.0005
R3598 GNDA.n2383 GNDA.t236 16.0005
R3599 GNDA.n55 GNDA.t278 16.0005
R3600 GNDA.n38 GNDA.t276 16.0005
R3601 GNDA.n2469 GNDA.t195 16.0005
R3602 GNDA.n60 GNDA.t258 16.0005
R3603 GNDA.n2638 GNDA.t268 16.0005
R3604 GNDA.n1559 GNDA.n1558 16.0005
R3605 GNDA.n1562 GNDA.n1559 16.0005
R3606 GNDA.n1563 GNDA.n1562 16.0005
R3607 GNDA.n1566 GNDA.n1563 16.0005
R3608 GNDA.n1567 GNDA.n1566 16.0005
R3609 GNDA.n1570 GNDA.n1567 16.0005
R3610 GNDA.n1571 GNDA.n1570 16.0005
R3611 GNDA.n1574 GNDA.n1571 16.0005
R3612 GNDA.n1555 GNDA.n1554 16.0005
R3613 GNDA.n1554 GNDA.n1551 16.0005
R3614 GNDA.n1551 GNDA.n1550 16.0005
R3615 GNDA.n1550 GNDA.n1547 16.0005
R3616 GNDA.n1547 GNDA.n1546 16.0005
R3617 GNDA.n1546 GNDA.n1543 16.0005
R3618 GNDA.n1543 GNDA.n1542 16.0005
R3619 GNDA.n1542 GNDA.n1539 16.0005
R3620 GNDA.n1538 GNDA.n1535 16.0005
R3621 GNDA.n1535 GNDA.n1534 16.0005
R3622 GNDA.n1534 GNDA.n1531 16.0005
R3623 GNDA.n1531 GNDA.n1530 16.0005
R3624 GNDA.n1530 GNDA.n1527 16.0005
R3625 GNDA.n1527 GNDA.n1526 16.0005
R3626 GNDA.n1526 GNDA.n1523 16.0005
R3627 GNDA.n1523 GNDA.n1522 16.0005
R3628 GNDA.n895 GNDA.n882 16.0005
R3629 GNDA.n895 GNDA.n894 16.0005
R3630 GNDA.n894 GNDA.n893 16.0005
R3631 GNDA.n893 GNDA.n890 16.0005
R3632 GNDA.n890 GNDA.n889 16.0005
R3633 GNDA.n889 GNDA.n886 16.0005
R3634 GNDA.n886 GNDA.n885 16.0005
R3635 GNDA.n885 GNDA.n798 16.0005
R3636 GNDA.n881 GNDA.n879 16.0005
R3637 GNDA.n879 GNDA.n876 16.0005
R3638 GNDA.n876 GNDA.n875 16.0005
R3639 GNDA.n875 GNDA.n872 16.0005
R3640 GNDA.n872 GNDA.n871 16.0005
R3641 GNDA.n871 GNDA.n868 16.0005
R3642 GNDA.n868 GNDA.n867 16.0005
R3643 GNDA.n867 GNDA.n864 16.0005
R3644 GNDA.n863 GNDA.n860 16.0005
R3645 GNDA.n860 GNDA.n859 16.0005
R3646 GNDA.n859 GNDA.n856 16.0005
R3647 GNDA.n856 GNDA.n855 16.0005
R3648 GNDA.n855 GNDA.n852 16.0005
R3649 GNDA.n852 GNDA.n851 16.0005
R3650 GNDA.n851 GNDA.n848 16.0005
R3651 GNDA.n848 GNDA.n847 16.0005
R3652 GNDA.n394 GNDA.n393 16.0005
R3653 GNDA.n395 GNDA.n394 16.0005
R3654 GNDA.n395 GNDA.n343 16.0005
R3655 GNDA.n401 GNDA.n343 16.0005
R3656 GNDA.n402 GNDA.n401 16.0005
R3657 GNDA.n403 GNDA.n402 16.0005
R3658 GNDA.n403 GNDA.n341 16.0005
R3659 GNDA.n408 GNDA.n341 16.0005
R3660 GNDA.n387 GNDA.n345 16.0005
R3661 GNDA.n387 GNDA.n386 16.0005
R3662 GNDA.n386 GNDA.n385 16.0005
R3663 GNDA.n385 GNDA.n347 16.0005
R3664 GNDA.n379 GNDA.n347 16.0005
R3665 GNDA.n379 GNDA.n378 16.0005
R3666 GNDA.n378 GNDA.n377 16.0005
R3667 GNDA.n377 GNDA.n349 16.0005
R3668 GNDA.n371 GNDA.n370 16.0005
R3669 GNDA.n370 GNDA.n369 16.0005
R3670 GNDA.n369 GNDA.n351 16.0005
R3671 GNDA.n364 GNDA.n351 16.0005
R3672 GNDA.n364 GNDA.n363 16.0005
R3673 GNDA.n363 GNDA.n362 16.0005
R3674 GNDA.n362 GNDA.n354 16.0005
R3675 GNDA.n354 GNDA.n323 16.0005
R3676 GNDA.n1901 GNDA.n1900 16.0005
R3677 GNDA.n1904 GNDA.n1901 16.0005
R3678 GNDA.n1905 GNDA.n1904 16.0005
R3679 GNDA.n1908 GNDA.n1905 16.0005
R3680 GNDA.n1909 GNDA.n1908 16.0005
R3681 GNDA.n1912 GNDA.n1909 16.0005
R3682 GNDA.n1914 GNDA.n1912 16.0005
R3683 GNDA.n1915 GNDA.n1914 16.0005
R3684 GNDA.n1897 GNDA.n1896 16.0005
R3685 GNDA.n1896 GNDA.n1893 16.0005
R3686 GNDA.n1893 GNDA.n1892 16.0005
R3687 GNDA.n1892 GNDA.n1889 16.0005
R3688 GNDA.n1889 GNDA.n1888 16.0005
R3689 GNDA.n1888 GNDA.n1885 16.0005
R3690 GNDA.n1885 GNDA.n1884 16.0005
R3691 GNDA.n1884 GNDA.n1881 16.0005
R3692 GNDA.n1880 GNDA.n1877 16.0005
R3693 GNDA.n1877 GNDA.n1876 16.0005
R3694 GNDA.n1876 GNDA.n1873 16.0005
R3695 GNDA.n1873 GNDA.n1872 16.0005
R3696 GNDA.n1872 GNDA.n1869 16.0005
R3697 GNDA.n1869 GNDA.n1868 16.0005
R3698 GNDA.n1868 GNDA.n1865 16.0005
R3699 GNDA.n1865 GNDA.n1864 16.0005
R3700 GNDA.n731 GNDA.n717 16.0005
R3701 GNDA.n731 GNDA.n730 16.0005
R3702 GNDA.n730 GNDA.n729 16.0005
R3703 GNDA.n729 GNDA.n726 16.0005
R3704 GNDA.n726 GNDA.n725 16.0005
R3705 GNDA.n725 GNDA.n722 16.0005
R3706 GNDA.n722 GNDA.n721 16.0005
R3707 GNDA.n721 GNDA.n718 16.0005
R3708 GNDA.n716 GNDA.n714 16.0005
R3709 GNDA.n714 GNDA.n711 16.0005
R3710 GNDA.n711 GNDA.n710 16.0005
R3711 GNDA.n710 GNDA.n707 16.0005
R3712 GNDA.n707 GNDA.n706 16.0005
R3713 GNDA.n706 GNDA.n703 16.0005
R3714 GNDA.n703 GNDA.n702 16.0005
R3715 GNDA.n702 GNDA.n699 16.0005
R3716 GNDA.n698 GNDA.n695 16.0005
R3717 GNDA.n695 GNDA.n694 16.0005
R3718 GNDA.n694 GNDA.n691 16.0005
R3719 GNDA.n691 GNDA.n690 16.0005
R3720 GNDA.n690 GNDA.n687 16.0005
R3721 GNDA.n687 GNDA.n686 16.0005
R3722 GNDA.n686 GNDA.n683 16.0005
R3723 GNDA.n683 GNDA.n682 16.0005
R3724 GNDA.n1460 GNDA.n1459 16.0005
R3725 GNDA.n1463 GNDA.n1460 16.0005
R3726 GNDA.n1464 GNDA.n1463 16.0005
R3727 GNDA.n1467 GNDA.n1464 16.0005
R3728 GNDA.n1468 GNDA.n1467 16.0005
R3729 GNDA.n1471 GNDA.n1468 16.0005
R3730 GNDA.n1472 GNDA.n1471 16.0005
R3731 GNDA.n1472 GNDA.n473 16.0005
R3732 GNDA.n1456 GNDA.n1455 16.0005
R3733 GNDA.n1455 GNDA.n1452 16.0005
R3734 GNDA.n1452 GNDA.n1451 16.0005
R3735 GNDA.n1451 GNDA.n1448 16.0005
R3736 GNDA.n1448 GNDA.n1447 16.0005
R3737 GNDA.n1447 GNDA.n1444 16.0005
R3738 GNDA.n1444 GNDA.n1443 16.0005
R3739 GNDA.n1443 GNDA.n1440 16.0005
R3740 GNDA.n1439 GNDA.n1436 16.0005
R3741 GNDA.n1436 GNDA.n1435 16.0005
R3742 GNDA.n1435 GNDA.n1432 16.0005
R3743 GNDA.n1432 GNDA.n1431 16.0005
R3744 GNDA.n1431 GNDA.n1428 16.0005
R3745 GNDA.n1428 GNDA.n1427 16.0005
R3746 GNDA.n1427 GNDA.n1424 16.0005
R3747 GNDA.n1424 GNDA.n1423 16.0005
R3748 GNDA.n1093 GNDA.n1090 16.0005
R3749 GNDA.n1097 GNDA.n1090 16.0005
R3750 GNDA.n975 GNDA.n933 16.0005
R3751 GNDA.n981 GNDA.n933 16.0005
R3752 GNDA.n982 GNDA.n981 16.0005
R3753 GNDA.n983 GNDA.n982 16.0005
R3754 GNDA.n983 GNDA.n931 16.0005
R3755 GNDA.n989 GNDA.n931 16.0005
R3756 GNDA.n990 GNDA.n989 16.0005
R3757 GNDA.n994 GNDA.n990 16.0005
R3758 GNDA.n974 GNDA.n973 16.0005
R3759 GNDA.n973 GNDA.n935 16.0005
R3760 GNDA.n967 GNDA.n935 16.0005
R3761 GNDA.n967 GNDA.n966 16.0005
R3762 GNDA.n966 GNDA.n965 16.0005
R3763 GNDA.n965 GNDA.n937 16.0005
R3764 GNDA.n959 GNDA.n937 16.0005
R3765 GNDA.n959 GNDA.n958 16.0005
R3766 GNDA.n957 GNDA.n939 16.0005
R3767 GNDA.n951 GNDA.n939 16.0005
R3768 GNDA.n951 GNDA.n950 16.0005
R3769 GNDA.n950 GNDA.n949 16.0005
R3770 GNDA.n949 GNDA.n941 16.0005
R3771 GNDA.n944 GNDA.n941 16.0005
R3772 GNDA.n944 GNDA.n917 16.0005
R3773 GNDA.n1029 GNDA.n917 16.0005
R3774 GNDA.n2076 GNDA.n2075 16.0005
R3775 GNDA.n2079 GNDA.n2076 16.0005
R3776 GNDA.n2080 GNDA.n2079 16.0005
R3777 GNDA.n2083 GNDA.n2080 16.0005
R3778 GNDA.n2084 GNDA.n2083 16.0005
R3779 GNDA.n2087 GNDA.n2084 16.0005
R3780 GNDA.n2089 GNDA.n2087 16.0005
R3781 GNDA.n2090 GNDA.n2089 16.0005
R3782 GNDA.n2072 GNDA.n2071 16.0005
R3783 GNDA.n2071 GNDA.n2068 16.0005
R3784 GNDA.n2068 GNDA.n2067 16.0005
R3785 GNDA.n2067 GNDA.n2064 16.0005
R3786 GNDA.n2064 GNDA.n2063 16.0005
R3787 GNDA.n2063 GNDA.n2060 16.0005
R3788 GNDA.n2060 GNDA.n2059 16.0005
R3789 GNDA.n2059 GNDA.n2056 16.0005
R3790 GNDA.n2055 GNDA.n2052 16.0005
R3791 GNDA.n2052 GNDA.n2051 16.0005
R3792 GNDA.n2051 GNDA.n2048 16.0005
R3793 GNDA.n2048 GNDA.n2047 16.0005
R3794 GNDA.n2047 GNDA.n2044 16.0005
R3795 GNDA.n2044 GNDA.n2043 16.0005
R3796 GNDA.n2043 GNDA.n2040 16.0005
R3797 GNDA.n2040 GNDA.n2039 16.0005
R3798 GNDA.n1360 GNDA.n1359 16.0005
R3799 GNDA.n1363 GNDA.n1360 16.0005
R3800 GNDA.n1364 GNDA.n1363 16.0005
R3801 GNDA.n1367 GNDA.n1364 16.0005
R3802 GNDA.n1368 GNDA.n1367 16.0005
R3803 GNDA.n1371 GNDA.n1368 16.0005
R3804 GNDA.n1372 GNDA.n1371 16.0005
R3805 GNDA.n1372 GNDA.n499 16.0005
R3806 GNDA.n1356 GNDA.n1355 16.0005
R3807 GNDA.n1355 GNDA.n1352 16.0005
R3808 GNDA.n1352 GNDA.n1351 16.0005
R3809 GNDA.n1351 GNDA.n1348 16.0005
R3810 GNDA.n1348 GNDA.n1347 16.0005
R3811 GNDA.n1347 GNDA.n1344 16.0005
R3812 GNDA.n1344 GNDA.n1343 16.0005
R3813 GNDA.n1343 GNDA.n1340 16.0005
R3814 GNDA.n1339 GNDA.n1336 16.0005
R3815 GNDA.n1336 GNDA.n1335 16.0005
R3816 GNDA.n1335 GNDA.n1332 16.0005
R3817 GNDA.n1332 GNDA.n1331 16.0005
R3818 GNDA.n1331 GNDA.n1328 16.0005
R3819 GNDA.n1328 GNDA.n1327 16.0005
R3820 GNDA.n1327 GNDA.n1324 16.0005
R3821 GNDA.n1324 GNDA.n1323 16.0005
R3822 GNDA.t184 GNDA.t125 15.4463
R3823 GNDA.t152 GNDA.t313 15.4463
R3824 GNDA.t288 GNDA.n2410 14.9467
R3825 GNDA.n2633 GNDA.t83 14.9467
R3826 GNDA.t16 GNDA.n2443 14.9467
R3827 GNDA.n2573 GNDA.n2572 14.9255
R3828 GNDA.n2569 GNDA.n2567 14.9255
R3829 GNDA.n2263 GNDA.n2262 14.9255
R3830 GNDA.n2259 GNDA.n2257 14.9255
R3831 GNDA.n1583 GNDA.n226 14.555
R3832 GNDA.n914 GNDA.n225 14.555
R3833 GNDA.n312 GNDA.n310 14.363
R3834 GNDA.n2323 GNDA.n2321 14.0818
R3835 GNDA.n2419 GNDA.n2418 14.0401
R3836 GNDA.n2429 GNDA.n2428 14.0401
R3837 GNDA.n2477 GNDA.n2476 14.0401
R3838 GNDA.n2646 GNDA.n2645 14.0401
R3839 GNDA.n2306 GNDA.n2305 14.0193
R3840 GNDA.n2616 GNDA.n2615 14.0193
R3841 GNDA.n1933 GNDA.n1932 13.8005
R3842 GNDA.n1955 GNDA.n1954 13.8005
R3843 GNDA.n1945 GNDA.n1944 13.8005
R3844 GNDA.n1942 GNDA.n1941 13.8005
R3845 GNDA.n2029 GNDA.n2028 13.8005
R3846 GNDA.n2356 GNDA.n2355 13.8005
R3847 GNDA.n2392 GNDA.n2391 13.8005
R3848 GNDA.n2448 GNDA.n31 13.8005
R3849 GNDA.n2133 GNDA.n132 12.7542
R3850 GNDA.n1751 GNDA.t182 12.3572
R3851 GNDA.n2161 GNDA.t158 12.3572
R3852 GNDA.t150 GNDA.n178 12.3572
R3853 GNDA.n2135 GNDA.n2134 12.2193
R3854 GNDA.n2570 GNDA.n3 12.1567
R3855 GNDA.n2260 GNDA.n2 12.1567
R3856 GNDA.n85 GNDA.n84 11.7557
R3857 GNDA.t124 GNDA.t12 11.7135
R3858 GNDA.n1607 GNDA.n1606 11.6369
R3859 GNDA.n1606 GNDA.n1605 11.6369
R3860 GNDA.n1605 GNDA.n1604 11.6369
R3861 GNDA.n1604 GNDA.n1602 11.6369
R3862 GNDA.n1602 GNDA.n1599 11.6369
R3863 GNDA.n1599 GNDA.n1598 11.6369
R3864 GNDA.n1598 GNDA.n1595 11.6369
R3865 GNDA.n1595 GNDA.n1594 11.6369
R3866 GNDA.n1594 GNDA.n1591 11.6369
R3867 GNDA.n1591 GNDA.n1590 11.6369
R3868 GNDA.n1154 GNDA.n427 11.6369
R3869 GNDA.n1155 GNDA.n1154 11.6369
R3870 GNDA.n1156 GNDA.n1155 11.6369
R3871 GNDA.n1156 GNDA.n1148 11.6369
R3872 GNDA.n1162 GNDA.n1148 11.6369
R3873 GNDA.n1163 GNDA.n1162 11.6369
R3874 GNDA.n1164 GNDA.n1163 11.6369
R3875 GNDA.n1164 GNDA.n1144 11.6369
R3876 GNDA.n1170 GNDA.n1144 11.6369
R3877 GNDA.n1171 GNDA.n1170 11.6369
R3878 GNDA.n1172 GNDA.n1171 11.6369
R3879 GNDA.n776 GNDA.n775 11.6369
R3880 GNDA.n779 GNDA.n776 11.6369
R3881 GNDA.n780 GNDA.n779 11.6369
R3882 GNDA.n783 GNDA.n780 11.6369
R3883 GNDA.n784 GNDA.n783 11.6369
R3884 GNDA.n787 GNDA.n784 11.6369
R3885 GNDA.n788 GNDA.n787 11.6369
R3886 GNDA.n791 GNDA.n788 11.6369
R3887 GNDA.n792 GNDA.n791 11.6369
R3888 GNDA.n795 GNDA.n792 11.6369
R3889 GNDA.n772 GNDA.n771 11.6369
R3890 GNDA.n771 GNDA.n768 11.6369
R3891 GNDA.n768 GNDA.n767 11.6369
R3892 GNDA.n767 GNDA.n764 11.6369
R3893 GNDA.n764 GNDA.n763 11.6369
R3894 GNDA.n763 GNDA.n760 11.6369
R3895 GNDA.n760 GNDA.n759 11.6369
R3896 GNDA.n759 GNDA.n756 11.6369
R3897 GNDA.n756 GNDA.n755 11.6369
R3898 GNDA.n755 GNDA.n259 11.6369
R3899 GNDA.n1993 GNDA.n259 11.6369
R3900 GNDA.n1710 GNDA.n1615 11.6369
R3901 GNDA.n1716 GNDA.n1615 11.6369
R3902 GNDA.n1717 GNDA.n1716 11.6369
R3903 GNDA.n1718 GNDA.n1717 11.6369
R3904 GNDA.n1718 GNDA.n1613 11.6369
R3905 GNDA.n1724 GNDA.n1613 11.6369
R3906 GNDA.n1725 GNDA.n1724 11.6369
R3907 GNDA.n1726 GNDA.n1725 11.6369
R3908 GNDA.n1726 GNDA.n1611 11.6369
R3909 GNDA.n1611 GNDA.n411 11.6369
R3910 GNDA.n526 GNDA.n260 11.6369
R3911 GNDA.n529 GNDA.n526 11.6369
R3912 GNDA.n530 GNDA.n529 11.6369
R3913 GNDA.n533 GNDA.n530 11.6369
R3914 GNDA.n534 GNDA.n533 11.6369
R3915 GNDA.n537 GNDA.n534 11.6369
R3916 GNDA.n538 GNDA.n537 11.6369
R3917 GNDA.n541 GNDA.n538 11.6369
R3918 GNDA.n542 GNDA.n541 11.6369
R3919 GNDA.n545 GNDA.n542 11.6369
R3920 GNDA.n546 GNDA.n545 11.6369
R3921 GNDA.n595 GNDA.n594 11.6369
R3922 GNDA.n598 GNDA.n595 11.6369
R3923 GNDA.n599 GNDA.n598 11.6369
R3924 GNDA.n602 GNDA.n599 11.6369
R3925 GNDA.n603 GNDA.n602 11.6369
R3926 GNDA.n606 GNDA.n603 11.6369
R3927 GNDA.n607 GNDA.n606 11.6369
R3928 GNDA.n610 GNDA.n607 11.6369
R3929 GNDA.n611 GNDA.n610 11.6369
R3930 GNDA.n614 GNDA.n611 11.6369
R3931 GNDA.n615 GNDA.n614 11.6369
R3932 GNDA.n1056 GNDA.n1055 11.6369
R3933 GNDA.n1055 GNDA.n1054 11.6369
R3934 GNDA.n1054 GNDA.n616 11.6369
R3935 GNDA.n1048 GNDA.n616 11.6369
R3936 GNDA.n1048 GNDA.n1047 11.6369
R3937 GNDA.n1047 GNDA.n1046 11.6369
R3938 GNDA.n1046 GNDA.n619 11.6369
R3939 GNDA.n623 GNDA.n619 11.6369
R3940 GNDA.n1039 GNDA.n623 11.6369
R3941 GNDA.n1039 GNDA.n1038 11.6369
R3942 GNDA.n1813 GNDA.n296 11.6369
R3943 GNDA.n1813 GNDA.n1812 11.6369
R3944 GNDA.n1812 GNDA.n1811 11.6369
R3945 GNDA.n1811 GNDA.n1791 11.6369
R3946 GNDA.n1806 GNDA.n1791 11.6369
R3947 GNDA.n1806 GNDA.n1805 11.6369
R3948 GNDA.n1805 GNDA.n1804 11.6369
R3949 GNDA.n1804 GNDA.n1794 11.6369
R3950 GNDA.n1799 GNDA.n1794 11.6369
R3951 GNDA.n1799 GNDA.n1798 11.6369
R3952 GNDA.n1798 GNDA.n201 11.6369
R3953 GNDA.n2000 GNDA.n1999 11.6369
R3954 GNDA.n2002 GNDA.n2000 11.6369
R3955 GNDA.n2002 GNDA.n2001 11.6369
R3956 GNDA.n2001 GNDA.n198 11.6369
R3957 GNDA.n198 GNDA.n196 11.6369
R3958 GNDA.n2010 GNDA.n196 11.6369
R3959 GNDA.n2011 GNDA.n2010 11.6369
R3960 GNDA.n2013 GNDA.n2011 11.6369
R3961 GNDA.n2013 GNDA.n2012 11.6369
R3962 GNDA.n2012 GNDA.n193 11.6369
R3963 GNDA.n1266 GNDA.n1265 11.6369
R3964 GNDA.n1266 GNDA.n1065 11.6369
R3965 GNDA.n1273 GNDA.n1065 11.6369
R3966 GNDA.n1274 GNDA.n1273 11.6369
R3967 GNDA.n1275 GNDA.n1274 11.6369
R3968 GNDA.n1275 GNDA.n1063 11.6369
R3969 GNDA.n1280 GNDA.n1063 11.6369
R3970 GNDA.n1281 GNDA.n1280 11.6369
R3971 GNDA.n1283 GNDA.n1281 11.6369
R3972 GNDA.n1283 GNDA.n1282 11.6369
R3973 GNDA.n1242 GNDA.n1241 11.6369
R3974 GNDA.n1242 GNDA.n1077 11.6369
R3975 GNDA.n1248 GNDA.n1077 11.6369
R3976 GNDA.n1249 GNDA.n1248 11.6369
R3977 GNDA.n1250 GNDA.n1249 11.6369
R3978 GNDA.n1250 GNDA.n1073 11.6369
R3979 GNDA.n1256 GNDA.n1073 11.6369
R3980 GNDA.n1257 GNDA.n1256 11.6369
R3981 GNDA.n1258 GNDA.n1257 11.6369
R3982 GNDA.n1258 GNDA.n1069 11.6369
R3983 GNDA.n1264 GNDA.n1069 11.6369
R3984 GNDA.n1179 GNDA.n1178 11.6369
R3985 GNDA.n1180 GNDA.n1179 11.6369
R3986 GNDA.n1180 GNDA.n1098 11.6369
R3987 GNDA.n1187 GNDA.n1098 11.6369
R3988 GNDA.n1188 GNDA.n1187 11.6369
R3989 GNDA.n1190 GNDA.n1087 11.6369
R3990 GNDA.n1197 GNDA.n1087 11.6369
R3991 GNDA.n1198 GNDA.n1197 11.6369
R3992 GNDA.n1199 GNDA.n1198 11.6369
R3993 GNDA.n1199 GNDA.n1081 11.6369
R3994 GNDA.n1649 GNDA.n1626 11.6369
R3995 GNDA.n1649 GNDA.n1648 11.6369
R3996 GNDA.n1648 GNDA.n1647 11.6369
R3997 GNDA.n1647 GNDA.n1629 11.6369
R3998 GNDA.n1642 GNDA.n1629 11.6369
R3999 GNDA.n1642 GNDA.n1641 11.6369
R4000 GNDA.n1641 GNDA.n1640 11.6369
R4001 GNDA.n1640 GNDA.n1632 11.6369
R4002 GNDA.n1635 GNDA.n1632 11.6369
R4003 GNDA.n1635 GNDA.n298 11.6369
R4004 GNDA.n1962 GNDA.n298 11.6369
R4005 GNDA.n1709 GNDA.n1708 11.6369
R4006 GNDA.n1708 GNDA.n1617 11.6369
R4007 GNDA.n1703 GNDA.n1617 11.6369
R4008 GNDA.n1703 GNDA.n1702 11.6369
R4009 GNDA.n1702 GNDA.n1701 11.6369
R4010 GNDA.n1701 GNDA.n1620 11.6369
R4011 GNDA.n1696 GNDA.n1620 11.6369
R4012 GNDA.n1696 GNDA.n1695 11.6369
R4013 GNDA.n1695 GNDA.n1694 11.6369
R4014 GNDA.n1694 GNDA.n1623 11.6369
R4015 GNDA.n1689 GNDA.n1623 11.6369
R4016 GNDA.t105 GNDA.t32 11.5188
R4017 GNDA.t301 GNDA.t142 11.5188
R4018 GNDA.n2028 GNDA.n2027 11.3792
R4019 GNDA.n28 GNDA.n3 10.8286
R4020 GNDA.t12 GNDA.t0 9.95658
R4021 GNDA.n2431 GNDA.n73 9.8005
R4022 GNDA.n2465 GNDA.n2464 9.8005
R4023 GNDA.n188 GNDA.n0 9.75668
R4024 GNDA.n217 GNDA.t77 9.6005
R4025 GNDA.n211 GNDA.t79 9.6005
R4026 GNDA.n2124 GNDA.t148 9.6005
R4027 GNDA.n134 GNDA.t78 9.6005
R4028 GNDA.n2348 GNDA.t203 9.6005
R4029 GNDA.n2340 GNDA.t109 9.6005
R4030 GNDA.n2340 GNDA.t46 9.6005
R4031 GNDA.n2338 GNDA.t70 9.6005
R4032 GNDA.n2338 GNDA.t44 9.6005
R4033 GNDA.n2336 GNDA.t19 9.6005
R4034 GNDA.n2336 GNDA.t6 9.6005
R4035 GNDA.n2334 GNDA.t55 9.6005
R4036 GNDA.n2334 GNDA.t132 9.6005
R4037 GNDA.n2332 GNDA.t116 9.6005
R4038 GNDA.n2332 GNDA.t129 9.6005
R4039 GNDA.n2330 GNDA.t59 9.6005
R4040 GNDA.n2330 GNDA.t134 9.6005
R4041 GNDA.n2328 GNDA.t57 9.6005
R4042 GNDA.n2328 GNDA.t130 9.6005
R4043 GNDA.n2326 GNDA.t111 9.6005
R4044 GNDA.n2326 GNDA.t53 9.6005
R4045 GNDA.n2324 GNDA.t8 9.6005
R4046 GNDA.n2324 GNDA.t114 9.6005
R4047 GNDA.n2322 GNDA.t72 9.6005
R4048 GNDA.n2322 GNDA.t222 9.6005
R4049 GNDA.n2314 GNDA.t223 9.6005
R4050 GNDA.n2374 GNDA.t197 9.6005
R4051 GNDA.n2368 GNDA.t17 9.6005
R4052 GNDA.n2368 GNDA.t112 9.6005
R4053 GNDA.n2447 GNDA.t263 9.6005
R4054 GNDA.n72 GNDA.t238 9.6005
R4055 GNDA.n39 GNDA.t30 9.6005
R4056 GNDA.n39 GNDA.t117 9.6005
R4057 GNDA.n47 GNDA.t285 9.6005
R4058 GNDA.n2648 GNDA.n1 9.54008
R4059 GNDA.n2432 GNDA.n2431 9.3005
R4060 GNDA.n2465 GNDA.n54 9.3005
R4061 GNDA.n2347 GNDA.n2344 9.14336
R4062 GNDA.n2351 GNDA.n2350 9.14336
R4063 GNDA.n2313 GNDA.n2310 9.14336
R4064 GNDA.n2317 GNDA.n2316 9.14336
R4065 GNDA.n2400 GNDA.n2397 9.14336
R4066 GNDA.n2380 GNDA.n2379 9.14336
R4067 GNDA.n2377 GNDA.n2375 9.14336
R4068 GNDA.n2457 GNDA.n2456 9.14336
R4069 GNDA.n2454 GNDA.n2452 9.14336
R4070 GNDA.n2487 GNDA.n2486 9.14336
R4071 GNDA.n2499 GNDA.n2496 9.14336
R4072 GNDA.n2298 GNDA.n2293 9.14336
R4073 GNDA.n2298 GNDA.n2297 9.14336
R4074 GNDA.n2297 GNDA.n2295 9.14336
R4075 GNDA.n2209 GNDA.n2201 9.14336
R4076 GNDA.n2209 GNDA.n2208 9.14336
R4077 GNDA.n2208 GNDA.n2206 9.14336
R4078 GNDA.n2413 GNDA.n2412 9.14336
R4079 GNDA.n2423 GNDA.n2421 9.14336
R4080 GNDA.n2440 GNDA.n2439 9.14336
R4081 GNDA.n2437 GNDA.n2436 9.14336
R4082 GNDA.n2385 GNDA.n2384 9.14336
R4083 GNDA.n46 GNDA.n43 9.14336
R4084 GNDA.n50 GNDA.n49 9.14336
R4085 GNDA.n2463 GNDA.n56 9.14336
R4086 GNDA.n2481 GNDA.n2480 9.14336
R4087 GNDA.n2470 GNDA.n2468 9.14336
R4088 GNDA.n64 GNDA.n63 9.14336
R4089 GNDA.n2640 GNDA.n2639 9.14336
R4090 GNDA.n2608 GNDA.n2603 9.14336
R4091 GNDA.n2608 GNDA.n2607 9.14336
R4092 GNDA.n2607 GNDA.n2605 9.14336
R4093 GNDA.n2624 GNDA.n15 9.14336
R4094 GNDA.n2624 GNDA.n2623 9.14336
R4095 GNDA.n2623 GNDA.n2621 9.14336
R4096 GNDA.n2596 GNDA.n2513 9.14336
R4097 GNDA.n2596 GNDA.n2595 9.14336
R4098 GNDA.n2595 GNDA.n2593 9.14336
R4099 GNDA.n2593 GNDA.n2590 9.14336
R4100 GNDA.n2590 GNDA.n2589 9.14336
R4101 GNDA.n2589 GNDA.n2586 9.14336
R4102 GNDA.n2586 GNDA.n2585 9.14336
R4103 GNDA.n2585 GNDA.n2582 9.14336
R4104 GNDA.n2582 GNDA.n2581 9.14336
R4105 GNDA.n2581 GNDA.n2578 9.14336
R4106 GNDA.n2578 GNDA.n2577 9.14336
R4107 GNDA.n2537 GNDA.n2534 9.14336
R4108 GNDA.n2541 GNDA.n2534 9.14336
R4109 GNDA.n2541 GNDA.n2532 9.14336
R4110 GNDA.n2547 GNDA.n2532 9.14336
R4111 GNDA.n2547 GNDA.n2530 9.14336
R4112 GNDA.n2551 GNDA.n2530 9.14336
R4113 GNDA.n2551 GNDA.n2528 9.14336
R4114 GNDA.n2557 GNDA.n2528 9.14336
R4115 GNDA.n2557 GNDA.n2526 9.14336
R4116 GNDA.n2561 GNDA.n2526 9.14336
R4117 GNDA.n2561 GNDA.n2524 9.14336
R4118 GNDA.n2286 GNDA.n2185 9.14336
R4119 GNDA.n2286 GNDA.n2285 9.14336
R4120 GNDA.n2285 GNDA.n2283 9.14336
R4121 GNDA.n2283 GNDA.n2280 9.14336
R4122 GNDA.n2280 GNDA.n2279 9.14336
R4123 GNDA.n2279 GNDA.n2276 9.14336
R4124 GNDA.n2276 GNDA.n2275 9.14336
R4125 GNDA.n2275 GNDA.n2272 9.14336
R4126 GNDA.n2272 GNDA.n2271 9.14336
R4127 GNDA.n2271 GNDA.n2268 9.14336
R4128 GNDA.n2268 GNDA.n2267 9.14336
R4129 GNDA.n2250 GNDA.n2221 9.14336
R4130 GNDA.n2250 GNDA.n2249 9.14336
R4131 GNDA.n2249 GNDA.n2247 9.14336
R4132 GNDA.n2247 GNDA.n2244 9.14336
R4133 GNDA.n2244 GNDA.n2243 9.14336
R4134 GNDA.n2243 GNDA.n2240 9.14336
R4135 GNDA.n2240 GNDA.n2239 9.14336
R4136 GNDA.n2239 GNDA.n2236 9.14336
R4137 GNDA.n2236 GNDA.n2235 9.14336
R4138 GNDA.n2235 GNDA.n2232 9.14336
R4139 GNDA.n2232 GNDA.n2231 9.14336
R4140 GNDA.n469 GNDA.n226 8.60107
R4141 GNDA.n1966 GNDA.n225 8.60107
R4142 GNDA.n2362 GNDA.n2361 8.53383
R4143 GNDA.n1750 GNDA.t154 8.23827
R4144 GNDA.t168 GNDA.n2138 8.23827
R4145 GNDA.t162 GNDA.n2119 8.23827
R4146 GNDA.n2023 GNDA.n167 8.19962
R4147 GNDA.t218 GNDA.t18 7.67938
R4148 GNDA.t64 GNDA.t7 7.67938
R4149 GNDA.n131 GNDA.n130 7.56675
R4150 GNDA.n1091 GNDA.n188 7.56675
R4151 GNDA.n2357 GNDA.n2356 7.5005
R4152 GNDA.n1766 GNDA.t92 7.20855
R4153 GNDA.n2096 GNDA.t149 7.20855
R4154 GNDA.t91 GNDA.n185 7.20855
R4155 GNDA.n2032 GNDA.n2031 7.20855
R4156 GNDA.n2647 GNDA.n2 6.78175
R4157 GNDA.n1172 GNDA.n1102 6.72373
R4158 GNDA.n1993 GNDA.n1992 6.72373
R4159 GNDA.n546 GNDA.n524 6.72373
R4160 GNDA.n1240 GNDA.n1081 6.72373
R4161 GNDA.n1963 GNDA.n1962 6.72373
R4162 GNDA.n1689 GNDA.n1688 6.72373
R4163 GNDA.n2357 GNDA.n2 6.688
R4164 GNDA.n1992 GNDA.n260 6.20656
R4165 GNDA.n594 GNDA.n524 6.20656
R4166 GNDA.n1963 GNDA.n296 6.20656
R4167 GNDA.n1241 GNDA.n1240 6.20656
R4168 GNDA.n1178 GNDA.n1102 6.20656
R4169 GNDA.n1688 GNDA.n1626 6.20656
R4170 GNDA.t100 GNDA.t191 6.17883
R4171 GNDA.n1189 GNDA.n1188 6.07727
R4172 GNDA.t24 GNDA.n2636 5.97926
R4173 GNDA.t48 GNDA.n2635 5.97926
R4174 GNDA.n2407 GNDA.t126 5.97926
R4175 GNDA.n2406 GNDA.t73 5.97926
R4176 GNDA.n2405 GNDA.t20 5.97926
R4177 GNDA.n2404 GNDA.t10 5.97926
R4178 GNDA.n2408 GNDA.t21 5.97926
R4179 GNDA.t270 GNDA.n35 5.97926
R4180 GNDA.t93 GNDA.n2637 5.97926
R4181 GNDA.n220 GNDA.n129 5.81868
R4182 GNDA.n220 GNDA.n219 5.81868
R4183 GNDA.n2304 GNDA.n2174 5.78934
R4184 GNDA.n2204 GNDA.n2203 5.78934
R4185 GNDA.n2614 GNDA.n29 5.78934
R4186 GNDA.n2619 GNDA.n2618 5.78934
R4187 GNDA.n2575 GNDA.n2574 5.78934
R4188 GNDA.n2566 GNDA.n2523 5.78934
R4189 GNDA.n2265 GNDA.n2264 5.78934
R4190 GNDA.n2256 GNDA.n2195 5.78934
R4191 GNDA.n131 GNDA.n0 5.737
R4192 GNDA.n2367 GNDA.n2358 5.563
R4193 GNDA.n1190 GNDA.n1189 5.5601
R4194 GNDA.n2307 GNDA.n2306 5.54068
R4195 GNDA.n2616 GNDA.n28 5.54068
R4196 GNDA.n1522 GNDA.n1493 5.51161
R4197 GNDA.n847 GNDA.n825 5.51161
R4198 GNDA.n1772 GNDA.n323 5.51161
R4199 GNDA.n1864 GNDA.n1775 5.51161
R4200 GNDA.n682 GNDA.n660 5.51161
R4201 GNDA.n1423 GNDA.n1393 5.51161
R4202 GNDA.n1030 GNDA.n1029 5.51161
R4203 GNDA.n2039 GNDA.n174 5.51161
R4204 GNDA.n1323 GNDA.n1293 5.51161
R4205 GNDA.n2419 GNDA.n85 5.46925
R4206 GNDA.n1037 GNDA.n624 5.1717
R4207 GNDA.n191 GNDA.n190 5.1717
R4208 GNDA.n1292 GNDA.n520 5.1717
R4209 GNDA.n2162 GNDA.t191 5.14911
R4210 GNDA.t47 GNDA.t248 5.14911
R4211 GNDA.n84 GNDA.n82 5.063
R4212 GNDA.n27 GNDA.n25 5.063
R4213 GNDA.n1587 GNDA.n428 4.9157
R4214 GNDA.n911 GNDA.n797 4.9157
R4215 GNDA.n1734 GNDA.n1733 4.9157
R4216 GNDA.n2646 GNDA.n3 4.71925
R4217 GNDA.n2307 GNDA.n85 4.6255
R4218 GNDA.n2466 GNDA.n2465 4.5005
R4219 GNDA.n2431 GNDA.n2430 4.5005
R4220 GNDA.n2648 GNDA.n2647 4.5005
R4221 GNDA.n2349 GNDA.n2344 4.46219
R4222 GNDA.n2351 GNDA.n2342 4.46219
R4223 GNDA.n2350 GNDA.n2349 4.46219
R4224 GNDA.n2354 GNDA.n2342 4.46219
R4225 GNDA.n2315 GNDA.n2310 4.46219
R4226 GNDA.n2317 GNDA.n2308 4.46219
R4227 GNDA.n2316 GNDA.n2315 4.46219
R4228 GNDA.n2320 GNDA.n2308 4.46219
R4229 GNDA.n2400 GNDA.n2399 4.46219
R4230 GNDA.n2399 GNDA.n2395 4.46219
R4231 GNDA.n2379 GNDA.n2378 4.46219
R4232 GNDA.n2375 GNDA.n2370 4.46219
R4233 GNDA.n2378 GNDA.n2377 4.46219
R4234 GNDA.n2390 GNDA.n2370 4.46219
R4235 GNDA.n2456 GNDA.n2455 4.46219
R4236 GNDA.n2452 GNDA.n2450 4.46219
R4237 GNDA.n2455 GNDA.n2454 4.46219
R4238 GNDA.n2450 GNDA.n2449 4.46219
R4239 GNDA.n2487 GNDA.n32 4.46219
R4240 GNDA.n2490 GNDA.n32 4.46219
R4241 GNDA.n2499 GNDA.n2498 4.46219
R4242 GNDA.n2498 GNDA.n2494 4.46219
R4243 GNDA.n2412 GNDA.n86 4.46219
R4244 GNDA.n2417 GNDA.n86 4.46219
R4245 GNDA.n2421 GNDA.n2420 4.46219
R4246 GNDA.n2427 GNDA.n2420 4.46219
R4247 GNDA.n2439 GNDA.n2438 4.46219
R4248 GNDA.n2436 GNDA.n2434 4.46219
R4249 GNDA.n2438 GNDA.n2437 4.46219
R4250 GNDA.n2434 GNDA.n2433 4.46219
R4251 GNDA.n2385 GNDA.n2382 4.46219
R4252 GNDA.n48 GNDA.n43 4.46219
R4253 GNDA.n50 GNDA.n41 4.46219
R4254 GNDA.n49 GNDA.n48 4.46219
R4255 GNDA.n53 GNDA.n41 4.46219
R4256 GNDA.n57 GNDA.n56 4.46219
R4257 GNDA.n2480 GNDA.n2479 4.46219
R4258 GNDA.n2479 GNDA.n2478 4.46219
R4259 GNDA.n2468 GNDA.n2467 4.46219
R4260 GNDA.n2474 GNDA.n2467 4.46219
R4261 GNDA.n63 GNDA.n62 4.46219
R4262 GNDA.n62 GNDA.n61 4.46219
R4263 GNDA.n2639 GNDA.n4 4.46219
R4264 GNDA.n2644 GNDA.n4 4.46219
R4265 GNDA.n1239 GNDA.n1083 4.26717
R4266 GNDA.n1233 GNDA.n1083 4.26717
R4267 GNDA.n1233 GNDA.n1232 4.26717
R4268 GNDA.n1232 GNDA.n1231 4.26717
R4269 GNDA.n1231 GNDA.n1210 4.26717
R4270 GNDA.n1226 GNDA.n1210 4.26717
R4271 GNDA.n1226 GNDA.n1225 4.26717
R4272 GNDA.n1225 GNDA.n1224 4.26717
R4273 GNDA.n1224 GNDA.n1216 4.26717
R4274 GNDA.n1216 GNDA.n497 4.26717
R4275 GNDA.n1388 GNDA.n497 4.26717
R4276 GNDA.n591 GNDA.n590 4.26717
R4277 GNDA.n590 GNDA.n551 4.26717
R4278 GNDA.n586 GNDA.n551 4.26717
R4279 GNDA.n586 GNDA.n585 4.26717
R4280 GNDA.n585 GNDA.n557 4.26717
R4281 GNDA.n580 GNDA.n557 4.26717
R4282 GNDA.n580 GNDA.n579 4.26717
R4283 GNDA.n579 GNDA.n578 4.26717
R4284 GNDA.n578 GNDA.n565 4.26717
R4285 GNDA.n572 GNDA.n565 4.26717
R4286 GNDA.n572 GNDA.n571 4.26717
R4287 GNDA.n1788 GNDA.n297 4.26717
R4288 GNDA.n1822 GNDA.n1788 4.26717
R4289 GNDA.n1823 GNDA.n1822 4.26717
R4290 GNDA.n1826 GNDA.n1823 4.26717
R4291 GNDA.n1826 GNDA.n1784 4.26717
R4292 GNDA.n1832 GNDA.n1784 4.26717
R4293 GNDA.n1833 GNDA.n1832 4.26717
R4294 GNDA.n1836 GNDA.n1833 4.26717
R4295 GNDA.n1836 GNDA.n1782 4.26717
R4296 GNDA.n1782 GNDA.n1779 4.26717
R4297 GNDA.n1843 GNDA.n1779 4.26717
R4298 GNDA.n1687 GNDA.n1627 4.26717
R4299 GNDA.n1682 GNDA.n1627 4.26717
R4300 GNDA.n1682 GNDA.n1681 4.26717
R4301 GNDA.n1681 GNDA.n1659 4.26717
R4302 GNDA.n1676 GNDA.n1659 4.26717
R4303 GNDA.n1676 GNDA.n1675 4.26717
R4304 GNDA.n1675 GNDA.n1674 4.26717
R4305 GNDA.n1674 GNDA.n1669 4.26717
R4306 GNDA.n1669 GNDA.n321 4.26717
R4307 GNDA.n1924 GNDA.n321 4.26717
R4308 GNDA.n1924 GNDA.n319 4.26717
R4309 GNDA.n1991 GNDA.n262 4.26717
R4310 GNDA.n1985 GNDA.n262 4.26717
R4311 GNDA.n1985 GNDA.n1984 4.26717
R4312 GNDA.n1984 GNDA.n1983 4.26717
R4313 GNDA.n1983 GNDA.n1981 4.26717
R4314 GNDA.n1981 GNDA.n1978 4.26717
R4315 GNDA.n1978 GNDA.n1977 4.26717
R4316 GNDA.n1977 GNDA.n1974 4.26717
R4317 GNDA.n1974 GNDA.n1973 4.26717
R4318 GNDA.n1973 GNDA.n1970 4.26717
R4319 GNDA.n1970 GNDA.n1969 4.26717
R4320 GNDA.n1142 GNDA.n1141 4.26717
R4321 GNDA.n1141 GNDA.n1108 4.26717
R4322 GNDA.n1135 GNDA.n1108 4.26717
R4323 GNDA.n1135 GNDA.n1134 4.26717
R4324 GNDA.n1134 GNDA.n1133 4.26717
R4325 GNDA.n1133 GNDA.n1116 4.26717
R4326 GNDA.n1118 GNDA.n1116 4.26717
R4327 GNDA.n1124 GNDA.n1118 4.26717
R4328 GNDA.n1125 GNDA.n1124 4.26717
R4329 GNDA.n1125 GNDA.n471 4.26717
R4330 GNDA.n1488 GNDA.n471 4.26717
R4331 GNDA GNDA.n2649 4.2117
R4332 GNDA.n2362 GNDA.n2359 4.17148
R4333 GNDA.n2365 GNDA.n2359 4.17148
R4334 GNDA.n2393 GNDA.n2367 4.15675
R4335 GNDA.n2134 GNDA.n2133 4.063
R4336 GNDA.n2409 GNDA.n2172 4.0593
R4337 GNDA.n2634 GNDA.n6 4.0593
R4338 GNDA.n2429 GNDA.n2419 4.0005
R4339 GNDA.n1240 GNDA.n1239 3.93531
R4340 GNDA.n591 GNDA.n524 3.93531
R4341 GNDA.n1963 GNDA.n297 3.93531
R4342 GNDA.n1688 GNDA.n1687 3.93531
R4343 GNDA.n1992 GNDA.n1991 3.93531
R4344 GNDA.n1142 GNDA.n1102 3.93531
R4345 GNDA.t292 GNDA.t25 3.83994
R4346 GNDA.t18 GNDA.t287 3.83994
R4347 GNDA.t135 GNDA.t302 3.83994
R4348 GNDA.n1572 GNDA.n447 3.7893
R4349 GNDA.n1580 GNDA.n1579 3.7893
R4350 GNDA.n1495 GNDA.n448 3.7893
R4351 GNDA.n1499 GNDA.n1497 3.7893
R4352 GNDA.n1504 GNDA.n1500 3.7893
R4353 GNDA.n1511 GNDA.n1510 3.7893
R4354 GNDA.n1514 GNDA.n1494 3.7893
R4355 GNDA.n1519 GNDA.n1515 3.7893
R4356 GNDA.n909 GNDA.n908 3.7893
R4357 GNDA.n905 GNDA.n800 3.7893
R4358 GNDA.n904 GNDA.n803 3.7893
R4359 GNDA.n901 GNDA.n900 3.7893
R4360 GNDA.n827 GNDA.n804 3.7893
R4361 GNDA.n836 GNDA.n835 3.7893
R4362 GNDA.n839 GNDA.n826 3.7893
R4363 GNDA.n844 GNDA.n840 3.7893
R4364 GNDA.n1741 GNDA.n1740 3.7893
R4365 GNDA.n1745 GNDA.n339 3.7893
R4366 GNDA.n1747 GNDA.n1746 3.7893
R4367 GNDA.n1754 GNDA.n336 3.7893
R4368 GNDA.n1753 GNDA.n334 3.7893
R4369 GNDA.n1762 GNDA.n1761 3.7893
R4370 GNDA.n331 GNDA.n330 3.7893
R4371 GNDA.n326 GNDA.n324 3.7893
R4372 GNDA.n2153 GNDA.n124 3.7893
R4373 GNDA.n2152 GNDA.n125 3.7893
R4374 GNDA.n2140 GNDA.n2139 3.7893
R4375 GNDA.n2146 GNDA.n2145 3.7893
R4376 GNDA.n2142 GNDA.n2141 3.7893
R4377 GNDA.n1851 GNDA.n103 3.7893
R4378 GNDA.n1854 GNDA.n1853 3.7893
R4379 GNDA.n1861 GNDA.n1776 3.7893
R4380 GNDA.n745 GNDA.n744 3.7893
R4381 GNDA.n741 GNDA.n635 3.7893
R4382 GNDA.n740 GNDA.n638 3.7893
R4383 GNDA.n737 GNDA.n736 3.7893
R4384 GNDA.n662 GNDA.n639 3.7893
R4385 GNDA.n671 GNDA.n670 3.7893
R4386 GNDA.n674 GNDA.n661 3.7893
R4387 GNDA.n679 GNDA.n675 3.7893
R4388 GNDA.n1482 GNDA.n474 3.7893
R4389 GNDA.n1479 GNDA.n1478 3.7893
R4390 GNDA.n1395 GNDA.n475 3.7893
R4391 GNDA.n1400 GNDA.n1398 3.7893
R4392 GNDA.n1405 GNDA.n1401 3.7893
R4393 GNDA.n1412 GNDA.n1411 3.7893
R4394 GNDA.n1415 GNDA.n1394 3.7893
R4395 GNDA.n1420 GNDA.n1416 3.7893
R4396 GNDA.n992 GNDA.n929 3.7893
R4397 GNDA.n1001 GNDA.n1000 3.7893
R4398 GNDA.n926 GNDA.n925 3.7893
R4399 GNDA.n1009 GNDA.n1007 3.7893
R4400 GNDA.n1008 GNDA.n923 3.7893
R4401 GNDA.n921 GNDA.n920 3.7893
R4402 GNDA.n1024 GNDA.n1022 3.7893
R4403 GNDA.n1023 GNDA.n916 3.7893
R4404 GNDA.n2111 GNDA.n163 3.7893
R4405 GNDA.n2110 GNDA.n164 3.7893
R4406 GNDA.n2098 GNDA.n2097 3.7893
R4407 GNDA.n2104 GNDA.n2103 3.7893
R4408 GNDA.n2100 GNDA.n2099 3.7893
R4409 GNDA.n179 GNDA.n142 3.7893
R4410 GNDA.n182 GNDA.n181 3.7893
R4411 GNDA.n2036 GNDA.n175 3.7893
R4412 GNDA.n1382 GNDA.n500 3.7893
R4413 GNDA.n1379 GNDA.n1378 3.7893
R4414 GNDA.n1295 GNDA.n501 3.7893
R4415 GNDA.n1300 GNDA.n1298 3.7893
R4416 GNDA.n1305 GNDA.n1301 3.7893
R4417 GNDA.n1312 GNDA.n1311 3.7893
R4418 GNDA.n1315 GNDA.n1294 3.7893
R4419 GNDA.n1320 GNDA.n1316 3.7893
R4420 GNDA.n1507 GNDA 3.7381
R4421 GNDA.n832 GNDA 3.7381
R4422 GNDA GNDA.n329 3.7381
R4423 GNDA GNDA.n2158 3.7381
R4424 GNDA.n667 GNDA 3.7381
R4425 GNDA.n1408 GNDA 3.7381
R4426 GNDA GNDA.n1015 3.7381
R4427 GNDA GNDA.n2116 3.7381
R4428 GNDA.n1308 GNDA 3.7381
R4429 GNDA.n2027 GNDA.n188 3.51962
R4430 GNDA.n2258 GNDA.t139 3.42907
R4431 GNDA.n2258 GNDA.t26 3.42907
R4432 GNDA.n2571 GNDA.t136 3.42907
R4433 GNDA.n2571 GNDA.t103 3.42907
R4434 GNDA.n2568 GNDA.t37 3.42907
R4435 GNDA.n2568 GNDA.t143 3.42907
R4436 GNDA.n2261 GNDA.t106 3.42907
R4437 GNDA.n2261 GNDA.t95 3.42907
R4438 GNDA.n2443 GNDA.n66 3.28629
R4439 GNDA.n2300 GNDA.n2293 3.19754
R4440 GNDA.n2295 GNDA.n2174 3.19754
R4441 GNDA.n2211 GNDA.n2201 3.19754
R4442 GNDA.n2206 GNDA.n2204 3.19754
R4443 GNDA.n2610 GNDA.n2603 3.19754
R4444 GNDA.n2605 GNDA.n29 3.19754
R4445 GNDA.n2626 GNDA.n15 3.19754
R4446 GNDA.n2621 GNDA.n2619 3.19754
R4447 GNDA.n2598 GNDA.n2513 3.19754
R4448 GNDA.n2577 GNDA.n2575 3.19754
R4449 GNDA.n2538 GNDA.n2537 3.19754
R4450 GNDA.n2524 GNDA.n2523 3.19754
R4451 GNDA.n2288 GNDA.n2185 3.19754
R4452 GNDA.n2267 GNDA.n2265 3.19754
R4453 GNDA.n2252 GNDA.n2221 3.19754
R4454 GNDA.n2231 GNDA.n2195 3.19754
R4455 GNDA.n1736 GNDA.n206 3.08966
R4456 GNDA.t65 GNDA.n1737 3.08966
R4457 GNDA.n327 GNDA.t38 3.08966
R4458 GNDA.n1769 GNDA.t34 3.08966
R4459 GNDA.n2108 GNDA.t294 3.08966
R4460 GNDA.n2358 GNDA.n2357 2.96925
R4461 GNDA.n2126 GNDA.n133 2.86505
R4462 GNDA.n2127 GNDA.n2126 2.86505
R4463 GNDA.n2125 GNDA.n2121 2.86505
R4464 GNDA.n2122 GNDA.n2121 2.86505
R4465 GNDA.n2128 GNDA.n2127 2.86505
R4466 GNDA.n2123 GNDA.n2122 2.86505
R4467 GNDA.n2132 GNDA.n133 2.86505
R4468 GNDA.n2128 GNDA.n2125 2.86505
R4469 GNDA.n218 GNDA.n214 2.86505
R4470 GNDA.n215 GNDA.n214 2.86505
R4471 GNDA.n216 GNDA.n215 2.86505
R4472 GNDA.n219 GNDA.n218 2.86505
R4473 GNDA.n1573 GNDA.n428 2.6629
R4474 GNDA.n1492 GNDA.n468 2.6629
R4475 GNDA.n911 GNDA.n910 2.6629
R4476 GNDA.n824 GNDA.n288 2.6629
R4477 GNDA.n1734 GNDA.n409 2.6629
R4478 GNDA.n1774 GNDA.n1773 2.6629
R4479 GNDA.n1917 GNDA.n1916 2.6629
R4480 GNDA.n1846 GNDA.n173 2.6629
R4481 GNDA.n634 GNDA.n633 2.6629
R4482 GNDA.n659 GNDA.n295 2.6629
R4483 GNDA.n1484 GNDA.n1483 2.6629
R4484 GNDA.n1392 GNDA.n494 2.6629
R4485 GNDA.n993 GNDA.n991 2.6629
R4486 GNDA.n2092 GNDA.n2091 2.6629
R4487 GNDA.n1384 GNDA.n1383 2.6629
R4488 GNDA.n1493 GNDA.n1492 2.4581
R4489 GNDA.n825 GNDA.n824 2.4581
R4490 GNDA.n1773 GNDA.n1772 2.4581
R4491 GNDA.n1917 GNDA.n1774 2.4581
R4492 GNDA.n1846 GNDA.n1775 2.4581
R4493 GNDA.n633 GNDA.n288 2.4581
R4494 GNDA.n660 GNDA.n659 2.4581
R4495 GNDA.n1484 GNDA.n468 2.4581
R4496 GNDA.n1393 GNDA.n1392 2.4581
R4497 GNDA.n991 GNDA.n295 2.4581
R4498 GNDA.n1030 GNDA.n624 2.4581
R4499 GNDA.n2092 GNDA.n173 2.4581
R4500 GNDA.n190 GNDA.n174 2.4581
R4501 GNDA.n1384 GNDA.n494 2.4581
R4502 GNDA.n1293 GNDA.n1292 2.4581
R4503 GNDA.n1388 GNDA.n494 2.18124
R4504 GNDA.n571 GNDA.n295 2.18124
R4505 GNDA.n1843 GNDA.n173 2.18124
R4506 GNDA.n1774 GNDA.n319 2.18124
R4507 GNDA.n1969 GNDA.n288 2.18124
R4508 GNDA.n1488 GNDA.n468 2.18124
R4509 GNDA.n1518 GNDA.n1493 2.1509
R4510 GNDA.n843 GNDA.n825 2.1509
R4511 GNDA.n1772 GNDA.n1771 2.1509
R4512 GNDA.n1860 GNDA.n1775 2.1509
R4513 GNDA.n678 GNDA.n660 2.1509
R4514 GNDA.n1419 GNDA.n1393 2.1509
R4515 GNDA.n1031 GNDA.n1030 2.1509
R4516 GNDA.n2035 GNDA.n174 2.1509
R4517 GNDA.n1319 GNDA.n1293 2.1509
R4518 GNDA.n1574 GNDA.n1573 2.13383
R4519 GNDA.n910 GNDA.n798 2.13383
R4520 GNDA.n409 GNDA.n408 2.13383
R4521 GNDA.n1916 GNDA.n1915 2.13383
R4522 GNDA.n718 GNDA.n634 2.13383
R4523 GNDA.n1483 GNDA.n473 2.13383
R4524 GNDA.n994 GNDA.n993 2.13383
R4525 GNDA.n2091 GNDA.n2090 2.13383
R4526 GNDA.n1383 GNDA.n499 2.13383
R4527 GNDA.n132 GNDA 2.09787
R4528 GNDA.n495 GNDA.n494 2.08643
R4529 GNDA.n1964 GNDA.n295 2.08643
R4530 GNDA.n1778 GNDA.n173 2.08643
R4531 GNDA.n1774 GNDA.n318 2.08643
R4532 GNDA.n290 GNDA.n288 2.08643
R4533 GNDA.n468 GNDA.n261 2.08643
R4534 GNDA.n1769 GNDA.t251 2.05994
R4535 GNDA.n1918 GNDA.t273 2.05994
R4536 GNDA.n1848 GNDA.t225 2.05994
R4537 GNDA.t248 GNDA.n2095 2.05994
R4538 GNDA.n1573 GNDA.n1572 1.9461
R4539 GNDA.n910 GNDA.n909 1.9461
R4540 GNDA.n1740 GNDA.n409 1.9461
R4541 GNDA.n1916 GNDA.n124 1.9461
R4542 GNDA.n745 GNDA.n634 1.9461
R4543 GNDA.n1483 GNDA.n1482 1.9461
R4544 GNDA.n993 GNDA.n992 1.9461
R4545 GNDA.n2091 GNDA.n163 1.9461
R4546 GNDA.n1383 GNDA.n1382 1.9461
R4547 GNDA.n2647 GNDA.n2646 1.938
R4548 GNDA.n1092 GNDA.n1091 1.90675
R4549 GNDA.n207 GNDA.t76 1.83728
R4550 GNDA.n2407 GNDA.t108 1.54702
R4551 GNDA.n2406 GNDA.t45 1.54702
R4552 GNDA.n2405 GNDA.t69 1.54702
R4553 GNDA.n2404 GNDA.t43 1.54702
R4554 GNDA.n2636 GNDA.t71 1.54702
R4555 GNDA.n2635 GNDA.t221 1.54702
R4556 GNDA.n2408 GNDA.t202 1.54702
R4557 GNDA.n35 GNDA.t52 1.54702
R4558 GNDA.n2637 GNDA.t113 1.54702
R4559 GNDA.n1590 GNDA.n1587 1.47392
R4560 GNDA.n797 GNDA.n795 1.47392
R4561 GNDA.n1733 GNDA.n411 1.47392
R4562 GNDA.n1038 GNDA.n1037 1.47392
R4563 GNDA.n193 GNDA.n191 1.47392
R4564 GNDA.n1282 GNDA.n520 1.47392
R4565 GNDA.n1945 GNDA.n1942 0.96925
R4566 GNDA.n1954 GNDA.n1933 0.96925
R4567 GNDA.n2358 GNDA.n2307 0.922375
R4568 GNDA.n2476 GNDA.n2466 0.8755
R4569 GNDA.n2430 GNDA.n2429 0.8755
R4570 GNDA.n1580 GNDA.n447 0.8197
R4571 GNDA.n1579 GNDA.n448 0.8197
R4572 GNDA.n1497 GNDA.n1495 0.8197
R4573 GNDA.n1500 GNDA.n1499 0.8197
R4574 GNDA.n1510 GNDA.n1507 0.8197
R4575 GNDA.n1511 GNDA.n1494 0.8197
R4576 GNDA.n1515 GNDA.n1514 0.8197
R4577 GNDA.n1519 GNDA.n1518 0.8197
R4578 GNDA.n908 GNDA.n800 0.8197
R4579 GNDA.n905 GNDA.n904 0.8197
R4580 GNDA.n901 GNDA.n803 0.8197
R4581 GNDA.n900 GNDA.n804 0.8197
R4582 GNDA.n835 GNDA.n832 0.8197
R4583 GNDA.n836 GNDA.n826 0.8197
R4584 GNDA.n840 GNDA.n839 0.8197
R4585 GNDA.n844 GNDA.n843 0.8197
R4586 GNDA.n1741 GNDA.n339 0.8197
R4587 GNDA.n1747 GNDA.n1745 0.8197
R4588 GNDA.n1746 GNDA.n336 0.8197
R4589 GNDA.n1754 GNDA.n1753 0.8197
R4590 GNDA.n1762 GNDA.n329 0.8197
R4591 GNDA.n1761 GNDA.n330 0.8197
R4592 GNDA.n331 GNDA.n326 0.8197
R4593 GNDA.n1771 GNDA.n324 0.8197
R4594 GNDA.n2153 GNDA.n2152 0.8197
R4595 GNDA.n2139 GNDA.n125 0.8197
R4596 GNDA.n2146 GNDA.n2140 0.8197
R4597 GNDA.n2145 GNDA.n2142 0.8197
R4598 GNDA.n2158 GNDA.n103 0.8197
R4599 GNDA.n1854 GNDA.n1851 0.8197
R4600 GNDA.n1853 GNDA.n1776 0.8197
R4601 GNDA.n1861 GNDA.n1860 0.8197
R4602 GNDA.n744 GNDA.n635 0.8197
R4603 GNDA.n741 GNDA.n740 0.8197
R4604 GNDA.n737 GNDA.n638 0.8197
R4605 GNDA.n736 GNDA.n639 0.8197
R4606 GNDA.n670 GNDA.n667 0.8197
R4607 GNDA.n671 GNDA.n661 0.8197
R4608 GNDA.n675 GNDA.n674 0.8197
R4609 GNDA.n679 GNDA.n678 0.8197
R4610 GNDA.n1479 GNDA.n474 0.8197
R4611 GNDA.n1478 GNDA.n475 0.8197
R4612 GNDA.n1398 GNDA.n1395 0.8197
R4613 GNDA.n1401 GNDA.n1400 0.8197
R4614 GNDA.n1411 GNDA.n1408 0.8197
R4615 GNDA.n1412 GNDA.n1394 0.8197
R4616 GNDA.n1416 GNDA.n1415 0.8197
R4617 GNDA.n1420 GNDA.n1419 0.8197
R4618 GNDA.n1001 GNDA.n929 0.8197
R4619 GNDA.n1000 GNDA.n926 0.8197
R4620 GNDA.n1007 GNDA.n925 0.8197
R4621 GNDA.n1009 GNDA.n1008 0.8197
R4622 GNDA.n1015 GNDA.n921 0.8197
R4623 GNDA.n1022 GNDA.n920 0.8197
R4624 GNDA.n1024 GNDA.n1023 0.8197
R4625 GNDA.n1031 GNDA.n916 0.8197
R4626 GNDA.n2111 GNDA.n2110 0.8197
R4627 GNDA.n2097 GNDA.n164 0.8197
R4628 GNDA.n2104 GNDA.n2098 0.8197
R4629 GNDA.n2103 GNDA.n2100 0.8197
R4630 GNDA.n2116 GNDA.n142 0.8197
R4631 GNDA.n182 GNDA.n179 0.8197
R4632 GNDA.n181 GNDA.n175 0.8197
R4633 GNDA.n2036 GNDA.n2035 0.8197
R4634 GNDA.n1379 GNDA.n500 0.8197
R4635 GNDA.n1378 GNDA.n501 0.8197
R4636 GNDA.n1298 GNDA.n1295 0.8197
R4637 GNDA.n1301 GNDA.n1300 0.8197
R4638 GNDA.n1311 GNDA.n1308 0.8197
R4639 GNDA.n1312 GNDA.n1294 0.8197
R4640 GNDA.n1316 GNDA.n1315 0.8197
R4641 GNDA.n1320 GNDA.n1319 0.8197
R4642 GNDA.n2393 GNDA.n2392 0.688
R4643 GNDA.n2492 GNDA.n31 0.6255
R4644 GNDA.n1610 GNDA.n207 0.575776
R4645 GNDA.n1504 GNDA 0.5637
R4646 GNDA GNDA.n827 0.5637
R4647 GNDA.n334 GNDA 0.5637
R4648 GNDA.n2141 GNDA 0.5637
R4649 GNDA GNDA.n662 0.5637
R4650 GNDA.n1405 GNDA 0.5637
R4651 GNDA.n923 GNDA 0.5637
R4652 GNDA.n2099 GNDA 0.5637
R4653 GNDA.n1305 GNDA 0.5637
R4654 GNDA.n2028 GNDA.n187 0.563
R4655 GNDA.n1935 GNDA.n187 0.563
R4656 GNDA.n1937 GNDA.n1935 0.563
R4657 GNDA.n1942 GNDA.n1937 0.563
R4658 GNDA.n1947 GNDA.n1945 0.563
R4659 GNDA.n1949 GNDA.n1947 0.563
R4660 GNDA.n1951 GNDA.n1949 0.563
R4661 GNDA.n1953 GNDA.n1951 0.563
R4662 GNDA.n1954 GNDA.n1953 0.563
R4663 GNDA.n1933 GNDA.n316 0.563
R4664 GNDA.n316 GNDA.n314 0.563
R4665 GNDA.n314 GNDA.n312 0.563
R4666 GNDA.n2325 GNDA.n2323 0.563
R4667 GNDA.n2327 GNDA.n2325 0.563
R4668 GNDA.n2329 GNDA.n2327 0.563
R4669 GNDA.n2331 GNDA.n2329 0.563
R4670 GNDA.n2333 GNDA.n2331 0.563
R4671 GNDA.n2335 GNDA.n2333 0.563
R4672 GNDA.n2337 GNDA.n2335 0.563
R4673 GNDA.n2339 GNDA.n2337 0.563
R4674 GNDA.n2341 GNDA.n2339 0.563
R4675 GNDA.n2356 GNDA.n2341 0.563
R4676 GNDA.n2369 GNDA.n31 0.563
R4677 GNDA.n2392 GNDA.n2369 0.563
R4678 GNDA.n2466 GNDA.n40 0.563
R4679 GNDA.n2430 GNDA.n40 0.563
R4680 GNDA.n78 GNDA.n76 0.563
R4681 GNDA.n80 GNDA.n78 0.563
R4682 GNDA.n82 GNDA.n80 0.563
R4683 GNDA.n21 GNDA.n19 0.563
R4684 GNDA.n23 GNDA.n21 0.563
R4685 GNDA.n25 GNDA.n23 0.563
R4686 GNDA.n2572 GNDA.n2570 0.5005
R4687 GNDA.n2570 GNDA.n2569 0.5005
R4688 GNDA.n2262 GNDA.n2260 0.5005
R4689 GNDA.n2260 GNDA.n2259 0.5005
R4690 GNDA.n2026 GNDA.n132 0.276625
R4691 GNDA GNDA.n1503 0.2565
R4692 GNDA.n830 GNDA 0.2565
R4693 GNDA GNDA.n333 0.2565
R4694 GNDA.n2159 GNDA 0.2565
R4695 GNDA.n665 GNDA 0.2565
R4696 GNDA GNDA.n1404 0.2565
R4697 GNDA.n1016 GNDA 0.2565
R4698 GNDA.n2117 GNDA 0.2565
R4699 GNDA GNDA.n1304 0.2565
R4700 GNDA.n2027 GNDA.n2026 0.22375
R4701 GNDA.n1503 GNDA 0.0517
R4702 GNDA GNDA.n830 0.0517
R4703 GNDA.n333 GNDA 0.0517
R4704 GNDA.n2159 GNDA 0.0517
R4705 GNDA GNDA.n665 0.0517
R4706 GNDA.n1404 GNDA 0.0517
R4707 GNDA.n1016 GNDA 0.0517
R4708 GNDA.n2117 GNDA 0.0517
R4709 GNDA.n1304 GNDA 0.0517
R4710 VDDA.n345 VDDA.t213 1212.4
R4711 VDDA.n409 VDDA.t191 1212.4
R4712 VDDA.n105 VDDA.t262 1212.4
R4713 VDDA.n174 VDDA.t274 1212.4
R4714 VDDA.n418 VDDA.t218 905.125
R4715 VDDA.n417 VDDA.t228 905.125
R4716 VDDA.n202 VDDA.t241 794.668
R4717 VDDA.n206 VDDA.t238 794.668
R4718 VDDA.n186 VDDA.t210 794.668
R4719 VDDA.n231 VDDA.t286 794.668
R4720 VDDA.n526 VDDA.t258 708.125
R4721 VDDA.t258 VDDA.n482 708.125
R4722 VDDA.n503 VDDA.t199 708.125
R4723 VDDA.t199 VDDA.n485 708.125
R4724 VDDA.n415 VDDA.n414 682
R4725 VDDA.n548 VDDA.t290 676.966
R4726 VDDA.n418 VDDA.t217 672.274
R4727 VDDA.t226 VDDA.n417 672.274
R4728 VDDA.n505 VDDA.t223 660.001
R4729 VDDA.t257 VDDA.n527 657.76
R4730 VDDA.t198 VDDA.n504 657.76
R4731 VDDA.n430 VDDA.t232 652.076
R4732 VDDA.n464 VDDA.t280 652.076
R4733 VDDA.n246 VDDA.t179 652.076
R4734 VDDA.n279 VDDA.t235 652.076
R4735 VDDA.n11 VDDA.t250 652.076
R4736 VDDA.n44 VDDA.t194 652.076
R4737 VDDA.t254 VDDA.n547 643.038
R4738 VDDA.t201 VDDA.n675 643.037
R4739 VDDA.n676 VDDA.t272 643.037
R4740 VDDA.t266 VDDA.n644 643.037
R4741 VDDA.n645 VDDA.t183 643.037
R4742 VDDA.t245 VDDA.n636 643.037
R4743 VDDA.n637 VDDA.t278 643.037
R4744 VDDA.n309 VDDA.t259 624.725
R4745 VDDA.n72 VDDA.t188 624.725
R4746 VDDA.n595 VDDA.t268 611.909
R4747 VDDA.n319 VDDA.t247 601.867
R4748 VDDA.n84 VDDA.t203 601.867
R4749 VDDA.n653 VDDA.t283 601.867
R4750 VDDA.n669 VDDA.t206 601.867
R4751 VDDA.n380 VDDA.n323 587.407
R4752 VDDA.n388 VDDA.n387 587.407
R4753 VDDA.n374 VDDA.n373 587.407
R4754 VDDA.n354 VDDA.n353 587.407
R4755 VDDA.n134 VDDA.n106 587.407
R4756 VDDA.n119 VDDA.n115 587.407
R4757 VDDA.n145 VDDA.n88 587.407
R4758 VDDA.n153 VDDA.n152 587.407
R4759 VDDA.n573 VDDA.n541 587.407
R4760 VDDA.n569 VDDA.n568 587.407
R4761 VDDA.n586 VDDA.n585 587.407
R4762 VDDA.n580 VDDA.n535 587.407
R4763 VDDA.n463 VDDA.n423 585
R4764 VDDA.n445 VDDA.n444 585
R4765 VDDA.n404 VDDA.n380 585
R4766 VDDA.n403 VDDA.n381 585
R4767 VDDA.n402 VDDA.n382 585
R4768 VDDA.n399 VDDA.n383 585
R4769 VDDA.n398 VDDA.n384 585
R4770 VDDA.n395 VDDA.n385 585
R4771 VDDA.n394 VDDA.n386 585
R4772 VDDA.n391 VDDA.n387 585
R4773 VDDA.n373 VDDA.n372 585
R4774 VDDA.n369 VDDA.n347 585
R4775 VDDA.n368 VDDA.n348 585
R4776 VDDA.n365 VDDA.n349 585
R4777 VDDA.n364 VDDA.n350 585
R4778 VDDA.n361 VDDA.n351 585
R4779 VDDA.n360 VDDA.n352 585
R4780 VDDA.n357 VDDA.n353 585
R4781 VDDA.n278 VDDA.n237 585
R4782 VDDA.n260 VDDA.n259 585
R4783 VDDA.n219 VDDA.n218 585
R4784 VDDA.n216 VDDA.n215 585
R4785 VDDA.n230 VDDA.n179 585
R4786 VDDA.n201 VDDA.n188 585
R4787 VDDA.n169 VDDA.n145 585
R4788 VDDA.n168 VDDA.n146 585
R4789 VDDA.n167 VDDA.n147 585
R4790 VDDA.n164 VDDA.n148 585
R4791 VDDA.n163 VDDA.n149 585
R4792 VDDA.n160 VDDA.n150 585
R4793 VDDA.n159 VDDA.n151 585
R4794 VDDA.n156 VDDA.n152 585
R4795 VDDA.n132 VDDA.n106 585
R4796 VDDA.n131 VDDA.n130 585
R4797 VDDA.n129 VDDA.n109 585
R4798 VDDA.n128 VDDA.n127 585
R4799 VDDA.n126 VDDA.n125 585
R4800 VDDA.n124 VDDA.n114 585
R4801 VDDA.n123 VDDA.n122 585
R4802 VDDA.n121 VDDA.n115 585
R4803 VDDA.n43 VDDA.n2 585
R4804 VDDA.n25 VDDA.n24 585
R4805 VDDA.n585 VDDA.n584 585
R4806 VDDA.n583 VDDA.n580 585
R4807 VDDA.n571 VDDA.n541 585
R4808 VDDA.n570 VDDA.n569 585
R4809 VDDA.n603 VDDA.t185 579.775
R4810 VDDA.n528 VDDA.t230 540.818
R4811 VDDA.n317 VDDA.t249 464.281
R4812 VDDA.n314 VDDA.t249 464.281
R4813 VDDA.n308 VDDA.t261 464.281
R4814 VDDA.t261 VDDA.n307 464.281
R4815 VDDA.n71 VDDA.t190 464.281
R4816 VDDA.t190 VDDA.n70 464.281
R4817 VDDA.t205 VDDA.n63 464.281
R4818 VDDA.n79 VDDA.t205 464.281
R4819 VDDA.t270 VDDA.n594 464.281
R4820 VDDA.t270 VDDA.n616 464.281
R4821 VDDA.n608 VDDA.t187 464.281
R4822 VDDA.t187 VDDA.n607 464.281
R4823 VDDA.n658 VDDA.t285 464.281
R4824 VDDA.n655 VDDA.t285 464.281
R4825 VDDA.n664 VDDA.t209 464.281
R4826 VDDA.t209 VDDA.n625 464.281
R4827 VDDA.n416 VDDA.t225 447.226
R4828 VDDA.n419 VDDA.t216 447.226
R4829 VDDA.n546 VDDA.t253 413.084
R4830 VDDA.n549 VDDA.t289 413.084
R4831 VDDA.n674 VDDA.t200 409.067
R4832 VDDA.n677 VDDA.t271 409.067
R4833 VDDA.n643 VDDA.t265 409.067
R4834 VDDA.n635 VDDA.t244 409.067
R4835 VDDA.n638 VDDA.t277 409.067
R4836 VDDA.t375 VDDA.t257 407.144
R4837 VDDA.t162 VDDA.t375 407.144
R4838 VDDA.t95 VDDA.t162 407.144
R4839 VDDA.t4 VDDA.t95 407.144
R4840 VDDA.t65 VDDA.t4 407.144
R4841 VDDA.t33 VDDA.t65 407.144
R4842 VDDA.t292 VDDA.t33 407.144
R4843 VDDA.t92 VDDA.t292 407.144
R4844 VDDA.t109 VDDA.t92 407.144
R4845 VDDA.t43 VDDA.t109 407.144
R4846 VDDA.t310 VDDA.t43 407.144
R4847 VDDA.t80 VDDA.t310 407.144
R4848 VDDA.t402 VDDA.t80 407.144
R4849 VDDA.t298 VDDA.t402 407.144
R4850 VDDA.t28 VDDA.t298 407.144
R4851 VDDA.t312 VDDA.t28 407.144
R4852 VDDA.t159 VDDA.t312 407.144
R4853 VDDA.t6 VDDA.t159 407.144
R4854 VDDA.t230 VDDA.t6 407.144
R4855 VDDA.t143 VDDA.t198 407.144
R4856 VDDA.t124 VDDA.t143 407.144
R4857 VDDA.t59 VDDA.t124 407.144
R4858 VDDA.t107 VDDA.t59 407.144
R4859 VDDA.t39 VDDA.t107 407.144
R4860 VDDA.t370 VDDA.t39 407.144
R4861 VDDA.t372 VDDA.t370 407.144
R4862 VDDA.t136 VDDA.t372 407.144
R4863 VDDA.t362 VDDA.t136 407.144
R4864 VDDA.t134 VDDA.t362 407.144
R4865 VDDA.t174 VDDA.t134 407.144
R4866 VDDA.t97 VDDA.t174 407.144
R4867 VDDA.t164 VDDA.t97 407.144
R4868 VDDA.t8 VDDA.t164 407.144
R4869 VDDA.t296 VDDA.t8 407.144
R4870 VDDA.t37 VDDA.t296 407.144
R4871 VDDA.t172 VDDA.t37 407.144
R4872 VDDA.t393 VDDA.t172 407.144
R4873 VDDA.t223 VDDA.t393 407.144
R4874 VDDA.n646 VDDA.t182 390.322
R4875 VDDA.n526 VDDA.t256 379.582
R4876 VDDA.n503 VDDA.t197 379.582
R4877 VDDA.t229 VDDA.n529 379.277
R4878 VDDA.t111 VDDA.t254 373.214
R4879 VDDA.t161 VDDA.t111 373.214
R4880 VDDA.t290 VDDA.t161 373.214
R4881 VDDA.t85 VDDA.t201 373.214
R4882 VDDA.t1 VDDA.t85 373.214
R4883 VDDA.t314 VDDA.t1 373.214
R4884 VDDA.t364 VDDA.t314 373.214
R4885 VDDA.t272 VDDA.t364 373.214
R4886 VDDA.t22 VDDA.t266 373.214
R4887 VDDA.t20 VDDA.t22 373.214
R4888 VDDA.t57 VDDA.t20 373.214
R4889 VDDA.t26 VDDA.t57 373.214
R4890 VDDA.t183 VDDA.t26 373.214
R4891 VDDA.t300 VDDA.t245 373.214
R4892 VDDA.t409 VDDA.t300 373.214
R4893 VDDA.t278 VDDA.t409 373.214
R4894 VDDA.n566 VDDA.t219 360.868
R4895 VDDA.n591 VDDA.t176 360.868
R4896 VDDA.n530 VDDA.t229 358.858
R4897 VDDA.t256 VDDA.n525 358.858
R4898 VDDA.n506 VDDA.t222 358.858
R4899 VDDA.t197 VDDA.n502 358.858
R4900 VDDA.n505 VDDA.t224 354.065
R4901 VDDA.n547 VDDA.t255 354.063
R4902 VDDA.n481 VDDA.t231 351.793
R4903 VDDA.n548 VDDA.t291 347.224
R4904 VDDA.n632 VDDA.n631 345.127
R4905 VDDA.n641 VDDA.n640 345.127
R4906 VDDA.n634 VDDA.n633 345.127
R4907 VDDA.n622 VDDA.n621 344.7
R4908 VDDA.n672 VDDA.n671 344.7
R4909 VDDA.n479 VDDA.n478 341.675
R4910 VDDA.n509 VDDA.n508 341.675
R4911 VDDA.n511 VDDA.n510 341.675
R4912 VDDA.n513 VDDA.n512 341.675
R4913 VDDA.n515 VDDA.n514 341.675
R4914 VDDA.n517 VDDA.n516 341.675
R4915 VDDA.n519 VDDA.n518 341.675
R4916 VDDA.n521 VDDA.n520 341.675
R4917 VDDA.n523 VDDA.n522 341.675
R4918 VDDA.n484 VDDA.n483 341.675
R4919 VDDA.n487 VDDA.n486 341.675
R4920 VDDA.n489 VDDA.n488 341.675
R4921 VDDA.n491 VDDA.n490 341.675
R4922 VDDA.n493 VDDA.n492 341.675
R4923 VDDA.n495 VDDA.n494 341.675
R4924 VDDA.n497 VDDA.n496 341.675
R4925 VDDA.n499 VDDA.n498 341.675
R4926 VDDA.n501 VDDA.n500 341.675
R4927 VDDA.n644 VDDA.t267 332.267
R4928 VDDA.n645 VDDA.t184 332.267
R4929 VDDA.n636 VDDA.t246 332.267
R4930 VDDA.n637 VDDA.t279 332.267
R4931 VDDA.n675 VDDA.t202 332.084
R4932 VDDA.n676 VDDA.t273 332.084
R4933 VDDA.n218 VDDA.n210 291.053
R4934 VDDA.n218 VDDA.n217 291.053
R4935 VDDA.n215 VDDA.n208 291.053
R4936 VDDA.n215 VDDA.n214 291.053
R4937 VDDA.n451 VDDA.n423 290.233
R4938 VDDA.n457 VDDA.n423 290.233
R4939 VDDA.n452 VDDA.n423 290.233
R4940 VDDA.n444 VDDA.n432 290.233
R4941 VDDA.n444 VDDA.n437 290.233
R4942 VDDA.n444 VDDA.n442 290.233
R4943 VDDA.n266 VDDA.n237 290.233
R4944 VDDA.n272 VDDA.n237 290.233
R4945 VDDA.n267 VDDA.n237 290.233
R4946 VDDA.n259 VDDA.n248 290.233
R4947 VDDA.n259 VDDA.n253 290.233
R4948 VDDA.n259 VDDA.n258 290.233
R4949 VDDA.n223 VDDA.n179 290.233
R4950 VDDA.n224 VDDA.n179 290.233
R4951 VDDA.n193 VDDA.n188 290.233
R4952 VDDA.n197 VDDA.n188 290.233
R4953 VDDA.n31 VDDA.n2 290.233
R4954 VDDA.n37 VDDA.n2 290.233
R4955 VDDA.n32 VDDA.n2 290.233
R4956 VDDA.n24 VDDA.n13 290.233
R4957 VDDA.n24 VDDA.n18 290.233
R4958 VDDA.n24 VDDA.n23 290.233
R4959 VDDA.n312 VDDA.t248 267.188
R4960 VDDA.t260 VDDA.n311 267.188
R4961 VDDA.t189 VDDA.n74 267.188
R4962 VDDA.n81 VDDA.t204 267.188
R4963 VDDA.n612 VDDA.t269 267.188
R4964 VDDA.t186 VDDA.n610 267.188
R4965 VDDA.t284 VDDA.n660 267.188
R4966 VDDA.n666 VDDA.t207 267.188
R4967 VDDA.t217 VDDA.t145 259.091
R4968 VDDA.t145 VDDA.t226 259.091
R4969 VDDA.t52 VDDA.t220 251.471
R4970 VDDA.t304 VDDA.t52 251.471
R4971 VDDA.t153 VDDA.t304 251.471
R4972 VDDA.t167 VDDA.t153 251.471
R4973 VDDA.t88 VDDA.t167 251.471
R4974 VDDA.t71 VDDA.t88 251.471
R4975 VDDA.t48 VDDA.t71 251.471
R4976 VDDA.t82 VDDA.t48 251.471
R4977 VDDA.t90 VDDA.t82 251.471
R4978 VDDA.t50 VDDA.t90 251.471
R4979 VDDA.t73 VDDA.t50 251.471
R4980 VDDA.t75 VDDA.t73 251.471
R4981 VDDA.t102 VDDA.t75 251.471
R4982 VDDA.t10 VDDA.t102 251.471
R4983 VDDA.t68 VDDA.t10 251.471
R4984 VDDA.t99 VDDA.t68 251.471
R4985 VDDA.t177 VDDA.t99 251.471
R4986 VDDA.n381 VDDA.n380 246.25
R4987 VDDA.n382 VDDA.n381 246.25
R4988 VDDA.n383 VDDA.n382 246.25
R4989 VDDA.n385 VDDA.n384 246.25
R4990 VDDA.n386 VDDA.n385 246.25
R4991 VDDA.n387 VDDA.n386 246.25
R4992 VDDA.n373 VDDA.n347 246.25
R4993 VDDA.n348 VDDA.n347 246.25
R4994 VDDA.n349 VDDA.n348 246.25
R4995 VDDA.n351 VDDA.n350 246.25
R4996 VDDA.n352 VDDA.n351 246.25
R4997 VDDA.n353 VDDA.n352 246.25
R4998 VDDA.n130 VDDA.n106 246.25
R4999 VDDA.n130 VDDA.n129 246.25
R5000 VDDA.n129 VDDA.n128 246.25
R5001 VDDA.n125 VDDA.n124 246.25
R5002 VDDA.n124 VDDA.n123 246.25
R5003 VDDA.n123 VDDA.n115 246.25
R5004 VDDA.n146 VDDA.n145 246.25
R5005 VDDA.n147 VDDA.n146 246.25
R5006 VDDA.n148 VDDA.n147 246.25
R5007 VDDA.n150 VDDA.n149 246.25
R5008 VDDA.n151 VDDA.n150 246.25
R5009 VDDA.n152 VDDA.n151 246.25
R5010 VDDA.n307 VDDA.n302 243.698
R5011 VDDA.n70 VDDA.n65 243.698
R5012 VDDA.n609 VDDA.n608 243.698
R5013 VDDA.n587 VDDA.n586 243.698
R5014 VDDA.n665 VDDA.n664 243.698
R5015 VDDA.n452 VDDA.n449 242.903
R5016 VDDA.n442 VDDA.n428 242.903
R5017 VDDA.n267 VDDA.n264 242.903
R5018 VDDA.n258 VDDA.n242 242.903
R5019 VDDA.n224 VDDA.n182 242.903
R5020 VDDA.n198 VDDA.n197 242.903
R5021 VDDA.n32 VDDA.n29 242.903
R5022 VDDA.n23 VDDA.n7 242.903
R5023 VDDA.n463 VDDA.n462 238.367
R5024 VDDA.n408 VDDA.n407 238.367
R5025 VDDA.n310 VDDA.n309 238.367
R5026 VDDA.n278 VDDA.n277 238.367
R5027 VDDA.n220 VDDA.n219 238.367
R5028 VDDA.n230 VDDA.n229 238.367
R5029 VDDA.n216 VDDA.n183 238.367
R5030 VDDA.n173 VDDA.n172 238.367
R5031 VDDA.n73 VDDA.n72 238.367
R5032 VDDA.n43 VDDA.n42 238.367
R5033 VDDA.n529 VDDA.n528 238.367
R5034 VDDA.n528 VDDA.n480 238.367
R5035 VDDA.n604 VDDA.n600 238.367
R5036 VDDA.n668 VDDA.n667 238.367
R5037 VDDA.t220 VDDA.n575 237.5
R5038 VDDA.n588 VDDA.t177 237.5
R5039 VDDA.n228 VDDA.t287 221.121
R5040 VDDA.t211 VDDA.n221 221.121
R5041 VDDA.n221 VDDA.t239 221.121
R5042 VDDA.n199 VDDA.t242 221.121
R5043 VDDA.t248 VDDA.t115 217.708
R5044 VDDA.t115 VDDA.t171 217.708
R5045 VDDA.t171 VDDA.t120 217.708
R5046 VDDA.t120 VDDA.t130 217.708
R5047 VDDA.t130 VDDA.t56 217.708
R5048 VDDA.t56 VDDA.t140 217.708
R5049 VDDA.t140 VDDA.t79 217.708
R5050 VDDA.t79 VDDA.t406 217.708
R5051 VDDA.t406 VDDA.t392 217.708
R5052 VDDA.t392 VDDA.t64 217.708
R5053 VDDA.t64 VDDA.t260 217.708
R5054 VDDA.t386 VDDA.t189 217.708
R5055 VDDA.t395 VDDA.t386 217.708
R5056 VDDA.t138 VDDA.t395 217.708
R5057 VDDA.t398 VDDA.t138 217.708
R5058 VDDA.t294 VDDA.t398 217.708
R5059 VDDA.t405 VDDA.t294 217.708
R5060 VDDA.t116 VDDA.t405 217.708
R5061 VDDA.t404 VDDA.t116 217.708
R5062 VDDA.t131 VDDA.t404 217.708
R5063 VDDA.t295 VDDA.t131 217.708
R5064 VDDA.t204 VDDA.t295 217.708
R5065 VDDA.t269 VDDA.t41 217.708
R5066 VDDA.t41 VDDA.t186 217.708
R5067 VDDA.t378 VDDA.t284 217.708
R5068 VDDA.t24 VDDA.t378 217.708
R5069 VDDA.t302 VDDA.t24 217.708
R5070 VDDA.t30 VDDA.t302 217.708
R5071 VDDA.t207 VDDA.t30 217.708
R5072 VDDA.n178 VDDA.n177 213.186
R5073 VDDA.n204 VDDA.n203 213.186
R5074 VDDA.n624 VDDA.n623 205.488
R5075 VDDA.n649 VDDA.n648 205.488
R5076 VDDA.n651 VDDA.n650 205.488
R5077 VDDA.n618 VDDA.n617 200.988
R5078 VDDA.n388 VDDA.n329 190.333
R5079 VDDA.n354 VDDA.n335 190.333
R5080 VDDA.n314 VDDA.n313 190.333
R5081 VDDA.n153 VDDA.n142 190.333
R5082 VDDA.n119 VDDA.n95 190.333
R5083 VDDA.n80 VDDA.n79 190.333
R5084 VDDA.n611 VDDA.n594 190.333
R5085 VDDA.n574 VDDA.n573 190.333
R5086 VDDA.n659 VDDA.n658 190.333
R5087 VDDA.n425 VDDA.n424 185
R5088 VDDA.n460 VDDA.n459 185
R5089 VDDA.n461 VDDA.n460 185
R5090 VDDA.n458 VDDA.n450 185
R5091 VDDA.n456 VDDA.n455 185
R5092 VDDA.n454 VDDA.n453 185
R5093 VDDA.n446 VDDA.n445 185
R5094 VDDA.n447 VDDA.n446 185
R5095 VDDA.n431 VDDA.n429 185
R5096 VDDA.n434 VDDA.n433 185
R5097 VDDA.n436 VDDA.n435 185
R5098 VDDA.n439 VDDA.n438 185
R5099 VDDA.n441 VDDA.n440 185
R5100 VDDA.n379 VDDA.n324 185
R5101 VDDA.n405 VDDA.n404 185
R5102 VDDA.n406 VDDA.n405 185
R5103 VDDA.n403 VDDA.n378 185
R5104 VDDA.n402 VDDA.n401 185
R5105 VDDA.n400 VDDA.n399 185
R5106 VDDA.n398 VDDA.n397 185
R5107 VDDA.n396 VDDA.n395 185
R5108 VDDA.n394 VDDA.n393 185
R5109 VDDA.n392 VDDA.n391 185
R5110 VDDA.n390 VDDA.n389 185
R5111 VDDA.n406 VDDA.n329 185
R5112 VDDA.n376 VDDA.n375 185
R5113 VDDA.n377 VDDA.n376 185
R5114 VDDA.n346 VDDA.n336 185
R5115 VDDA.n372 VDDA.n371 185
R5116 VDDA.n370 VDDA.n369 185
R5117 VDDA.n368 VDDA.n367 185
R5118 VDDA.n366 VDDA.n365 185
R5119 VDDA.n364 VDDA.n363 185
R5120 VDDA.n362 VDDA.n361 185
R5121 VDDA.n360 VDDA.n359 185
R5122 VDDA.n358 VDDA.n357 185
R5123 VDDA.n356 VDDA.n355 185
R5124 VDDA.n377 VDDA.n335 185
R5125 VDDA.n304 VDDA.n303 185
R5126 VDDA.n306 VDDA.n305 185
R5127 VDDA.n318 VDDA.n298 185
R5128 VDDA.n312 VDDA.n298 185
R5129 VDDA.n316 VDDA.n299 185
R5130 VDDA.n315 VDDA.n300 185
R5131 VDDA.n313 VDDA.n312 185
R5132 VDDA.n239 VDDA.n238 185
R5133 VDDA.n275 VDDA.n274 185
R5134 VDDA.n276 VDDA.n275 185
R5135 VDDA.n273 VDDA.n265 185
R5136 VDDA.n271 VDDA.n270 185
R5137 VDDA.n269 VDDA.n268 185
R5138 VDDA.n261 VDDA.n260 185
R5139 VDDA.n262 VDDA.n261 185
R5140 VDDA.n247 VDDA.n243 185
R5141 VDDA.n250 VDDA.n249 185
R5142 VDDA.n252 VDDA.n251 185
R5143 VDDA.n255 VDDA.n254 185
R5144 VDDA.n257 VDDA.n256 185
R5145 VDDA.n181 VDDA.n180 185
R5146 VDDA.n227 VDDA.n226 185
R5147 VDDA.n228 VDDA.n227 185
R5148 VDDA.n225 VDDA.n222 185
R5149 VDDA.n209 VDDA.n185 185
R5150 VDDA.n213 VDDA.n184 185
R5151 VDDA.n221 VDDA.n184 185
R5152 VDDA.n212 VDDA.n211 185
R5153 VDDA.n201 VDDA.n200 185
R5154 VDDA.n200 VDDA.n199 185
R5155 VDDA.n190 VDDA.n189 185
R5156 VDDA.n195 VDDA.n194 185
R5157 VDDA.n196 VDDA.n192 185
R5158 VDDA.n144 VDDA.n89 185
R5159 VDDA.n170 VDDA.n169 185
R5160 VDDA.n171 VDDA.n170 185
R5161 VDDA.n168 VDDA.n143 185
R5162 VDDA.n167 VDDA.n166 185
R5163 VDDA.n165 VDDA.n164 185
R5164 VDDA.n163 VDDA.n162 185
R5165 VDDA.n161 VDDA.n160 185
R5166 VDDA.n159 VDDA.n158 185
R5167 VDDA.n157 VDDA.n156 185
R5168 VDDA.n155 VDDA.n154 185
R5169 VDDA.n171 VDDA.n142 185
R5170 VDDA.n136 VDDA.n135 185
R5171 VDDA.n137 VDDA.n136 185
R5172 VDDA.n133 VDDA.n96 185
R5173 VDDA.n132 VDDA.n107 185
R5174 VDDA.n131 VDDA.n108 185
R5175 VDDA.n110 VDDA.n109 185
R5176 VDDA.n127 VDDA.n111 185
R5177 VDDA.n126 VDDA.n112 185
R5178 VDDA.n114 VDDA.n113 185
R5179 VDDA.n122 VDDA.n116 185
R5180 VDDA.n121 VDDA.n117 185
R5181 VDDA.n120 VDDA.n118 185
R5182 VDDA.n137 VDDA.n95 185
R5183 VDDA.n67 VDDA.n66 185
R5184 VDDA.n69 VDDA.n68 185
R5185 VDDA.n83 VDDA.n82 185
R5186 VDDA.n82 VDDA.n81 185
R5187 VDDA.n77 VDDA.n64 185
R5188 VDDA.n78 VDDA.n76 185
R5189 VDDA.n81 VDDA.n80 185
R5190 VDDA.n4 VDDA.n3 185
R5191 VDDA.n40 VDDA.n39 185
R5192 VDDA.n41 VDDA.n40 185
R5193 VDDA.n38 VDDA.n30 185
R5194 VDDA.n36 VDDA.n35 185
R5195 VDDA.n34 VDDA.n33 185
R5196 VDDA.n26 VDDA.n25 185
R5197 VDDA.n27 VDDA.n26 185
R5198 VDDA.n12 VDDA.n8 185
R5199 VDDA.n15 VDDA.n14 185
R5200 VDDA.n17 VDDA.n16 185
R5201 VDDA.n20 VDDA.n19 185
R5202 VDDA.n22 VDDA.n21 185
R5203 VDDA.n602 VDDA.n601 185
R5204 VDDA.n606 VDDA.n605 185
R5205 VDDA.n612 VDDA.n611 185
R5206 VDDA.n599 VDDA.n597 185
R5207 VDDA.n615 VDDA.n614 185
R5208 VDDA.n598 VDDA.n596 185
R5209 VDDA.n612 VDDA.n598 185
R5210 VDDA.n579 VDDA.n578 185
R5211 VDDA.n584 VDDA.n577 185
R5212 VDDA.n588 VDDA.n577 185
R5213 VDDA.n583 VDDA.n582 185
R5214 VDDA.n581 VDDA.n536 185
R5215 VDDA.n590 VDDA.n589 185
R5216 VDDA.n589 VDDA.n588 185
R5217 VDDA.n575 VDDA.n574 185
R5218 VDDA.n572 VDDA.n540 185
R5219 VDDA.n571 VDDA.n542 185
R5220 VDDA.n570 VDDA.n543 185
R5221 VDDA.n545 VDDA.n544 185
R5222 VDDA.n567 VDDA.n539 185
R5223 VDDA.n575 VDDA.n539 185
R5224 VDDA.n663 VDDA.n661 185
R5225 VDDA.n662 VDDA.n626 185
R5226 VDDA.n660 VDDA.n659 185
R5227 VDDA.n657 VDDA.n629 185
R5228 VDDA.n656 VDDA.n630 185
R5229 VDDA.n654 VDDA.n628 185
R5230 VDDA.n660 VDDA.n628 185
R5231 VDDA.t287 VDDA.t67 180.173
R5232 VDDA.t67 VDDA.t380 180.173
R5233 VDDA.t380 VDDA.t157 180.173
R5234 VDDA.t157 VDDA.t3 180.173
R5235 VDDA.t3 VDDA.t211 180.173
R5236 VDDA.t0 VDDA.t239 180.173
R5237 VDDA.t18 VDDA.t0 180.173
R5238 VDDA.t308 VDDA.t18 180.173
R5239 VDDA.t411 VDDA.t308 180.173
R5240 VDDA.t242 VDDA.t411 180.173
R5241 VDDA.t233 VDDA.n447 170.513
R5242 VDDA.n461 VDDA.t281 170.513
R5243 VDDA.t180 VDDA.n262 170.513
R5244 VDDA.n276 VDDA.t236 170.513
R5245 VDDA.t251 VDDA.n27 170.513
R5246 VDDA.n41 VDDA.t195 170.513
R5247 VDDA.n534 VDDA.n533 168.435
R5248 VDDA.n552 VDDA.n551 168.435
R5249 VDDA.n554 VDDA.n553 168.435
R5250 VDDA.n556 VDDA.n555 168.435
R5251 VDDA.n558 VDDA.n557 168.435
R5252 VDDA.n560 VDDA.n559 168.435
R5253 VDDA.n562 VDDA.n561 168.435
R5254 VDDA.n564 VDDA.n563 168.435
R5255 VDDA.n443 VDDA.n422 159.803
R5256 VDDA.n236 VDDA.n235 159.803
R5257 VDDA.n245 VDDA.n244 159.803
R5258 VDDA.n281 VDDA.n280 159.803
R5259 VDDA.n283 VDDA.n282 159.803
R5260 VDDA.n1 VDDA.n0 159.803
R5261 VDDA.n10 VDDA.n9 159.803
R5262 VDDA.n46 VDDA.n45 159.803
R5263 VDDA.n48 VDDA.n47 159.803
R5264 VDDA.n286 VDDA.n285 155.303
R5265 VDDA.n51 VDDA.n50 155.303
R5266 VDDA.n460 VDDA.n425 150
R5267 VDDA.n460 VDDA.n450 150
R5268 VDDA.n455 VDDA.n454 150
R5269 VDDA.n446 VDDA.n429 150
R5270 VDDA.n435 VDDA.n434 150
R5271 VDDA.n440 VDDA.n439 150
R5272 VDDA.n405 VDDA.n324 150
R5273 VDDA.n405 VDDA.n378 150
R5274 VDDA.n401 VDDA.n400 150
R5275 VDDA.n397 VDDA.n396 150
R5276 VDDA.n393 VDDA.n392 150
R5277 VDDA.n389 VDDA.n329 150
R5278 VDDA.n376 VDDA.n336 150
R5279 VDDA.n371 VDDA.n370 150
R5280 VDDA.n367 VDDA.n366 150
R5281 VDDA.n363 VDDA.n362 150
R5282 VDDA.n359 VDDA.n358 150
R5283 VDDA.n355 VDDA.n335 150
R5284 VDDA.n305 VDDA.n303 150
R5285 VDDA.n299 VDDA.n298 150
R5286 VDDA.n313 VDDA.n300 150
R5287 VDDA.n275 VDDA.n239 150
R5288 VDDA.n275 VDDA.n265 150
R5289 VDDA.n270 VDDA.n269 150
R5290 VDDA.n261 VDDA.n243 150
R5291 VDDA.n251 VDDA.n250 150
R5292 VDDA.n256 VDDA.n255 150
R5293 VDDA.n185 VDDA.n184 150
R5294 VDDA.n211 VDDA.n184 150
R5295 VDDA.n227 VDDA.n181 150
R5296 VDDA.n227 VDDA.n222 150
R5297 VDDA.n200 VDDA.n190 150
R5298 VDDA.n194 VDDA.n192 150
R5299 VDDA.n170 VDDA.n89 150
R5300 VDDA.n170 VDDA.n143 150
R5301 VDDA.n166 VDDA.n165 150
R5302 VDDA.n162 VDDA.n161 150
R5303 VDDA.n158 VDDA.n157 150
R5304 VDDA.n154 VDDA.n142 150
R5305 VDDA.n136 VDDA.n96 150
R5306 VDDA.n108 VDDA.n107 150
R5307 VDDA.n111 VDDA.n110 150
R5308 VDDA.n113 VDDA.n112 150
R5309 VDDA.n117 VDDA.n116 150
R5310 VDDA.n118 VDDA.n95 150
R5311 VDDA.n68 VDDA.n66 150
R5312 VDDA.n82 VDDA.n64 150
R5313 VDDA.n80 VDDA.n76 150
R5314 VDDA.n40 VDDA.n4 150
R5315 VDDA.n40 VDDA.n30 150
R5316 VDDA.n35 VDDA.n34 150
R5317 VDDA.n26 VDDA.n8 150
R5318 VDDA.n16 VDDA.n15 150
R5319 VDDA.n21 VDDA.n20 150
R5320 VDDA.n605 VDDA.n601 150
R5321 VDDA.n611 VDDA.n599 150
R5322 VDDA.n614 VDDA.n598 150
R5323 VDDA.n578 VDDA.n577 150
R5324 VDDA.n582 VDDA.n577 150
R5325 VDDA.n589 VDDA.n536 150
R5326 VDDA.n574 VDDA.n540 150
R5327 VDDA.n543 VDDA.n542 150
R5328 VDDA.n544 VDDA.n539 150
R5329 VDDA.n661 VDDA.n626 150
R5330 VDDA.n659 VDDA.n629 150
R5331 VDDA.n630 VDDA.n628 150
R5332 VDDA.t348 VDDA.t233 146.155
R5333 VDDA.t281 VDDA.t348 146.155
R5334 VDDA.t326 VDDA.t180 146.155
R5335 VDDA.t336 VDDA.t326 146.155
R5336 VDDA.t344 VDDA.t336 146.155
R5337 VDDA.t352 VDDA.t344 146.155
R5338 VDDA.t356 VDDA.t352 146.155
R5339 VDDA.t320 VDDA.t356 146.155
R5340 VDDA.t330 VDDA.t320 146.155
R5341 VDDA.t338 VDDA.t330 146.155
R5342 VDDA.t334 VDDA.t338 146.155
R5343 VDDA.t342 VDDA.t334 146.155
R5344 VDDA.t236 VDDA.t342 146.155
R5345 VDDA.t350 VDDA.t251 146.155
R5346 VDDA.t354 VDDA.t350 146.155
R5347 VDDA.t318 VDDA.t354 146.155
R5348 VDDA.t328 VDDA.t318 146.155
R5349 VDDA.t324 VDDA.t328 146.155
R5350 VDDA.t332 VDDA.t324 146.155
R5351 VDDA.t340 VDDA.t332 146.155
R5352 VDDA.t346 VDDA.t340 146.155
R5353 VDDA.t322 VDDA.t346 146.155
R5354 VDDA.t316 VDDA.t322 146.155
R5355 VDDA.t195 VDDA.t316 146.155
R5356 VDDA.n322 VDDA.n321 145.429
R5357 VDDA.n338 VDDA.n337 145.429
R5358 VDDA.n340 VDDA.n339 145.429
R5359 VDDA.n342 VDDA.n341 145.429
R5360 VDDA.n344 VDDA.n343 145.429
R5361 VDDA.n87 VDDA.n86 145.429
R5362 VDDA.n98 VDDA.n97 145.429
R5363 VDDA.n100 VDDA.n99 145.429
R5364 VDDA.n102 VDDA.n101 145.429
R5365 VDDA.n104 VDDA.n103 145.429
R5366 VDDA.t193 VDDA.n383 123.126
R5367 VDDA.n384 VDDA.t193 123.126
R5368 VDDA.t215 VDDA.n349 123.126
R5369 VDDA.n350 VDDA.t215 123.126
R5370 VDDA.n128 VDDA.t264 123.126
R5371 VDDA.n125 VDDA.t264 123.126
R5372 VDDA.t276 VDDA.n148 123.126
R5373 VDDA.n149 VDDA.t276 123.126
R5374 VDDA.t221 VDDA.n541 123.126
R5375 VDDA.n569 VDDA.t221 123.126
R5376 VDDA.n585 VDDA.t178 123.126
R5377 VDDA.n580 VDDA.t178 123.126
R5378 VDDA.n406 VDDA.t192 100.195
R5379 VDDA.t214 VDDA.n377 100.195
R5380 VDDA.t263 VDDA.n137 100.195
R5381 VDDA.n171 VDDA.t275 100.195
R5382 VDDA.n289 VDDA.n287 97.4002
R5383 VDDA.n54 VDDA.n52 97.4002
R5384 VDDA.n297 VDDA.n296 96.8377
R5385 VDDA.n295 VDDA.n294 96.8377
R5386 VDDA.n293 VDDA.n292 96.8377
R5387 VDDA.n291 VDDA.n290 96.8377
R5388 VDDA.n289 VDDA.n288 96.8377
R5389 VDDA.n62 VDDA.n61 96.8377
R5390 VDDA.n60 VDDA.n59 96.8377
R5391 VDDA.n58 VDDA.n57 96.8377
R5392 VDDA.n56 VDDA.n55 96.8377
R5393 VDDA.n54 VDDA.n53 96.8377
R5394 VDDA.t192 VDDA.t16 81.6411
R5395 VDDA.t16 VDDA.t113 81.6411
R5396 VDDA.t113 VDDA.t128 81.6411
R5397 VDDA.t128 VDDA.t399 81.6411
R5398 VDDA.t399 VDDA.t54 81.6411
R5399 VDDA.t54 VDDA.t118 81.6411
R5400 VDDA.t118 VDDA.t141 81.6411
R5401 VDDA.t141 VDDA.t35 81.6411
R5402 VDDA.t35 VDDA.t407 81.6411
R5403 VDDA.t407 VDDA.t122 81.6411
R5404 VDDA.t122 VDDA.t214 81.6411
R5405 VDDA.t61 VDDA.t263 81.6411
R5406 VDDA.t396 VDDA.t61 81.6411
R5407 VDDA.t384 VDDA.t396 81.6411
R5408 VDDA.t387 VDDA.t384 81.6411
R5409 VDDA.t132 VDDA.t387 81.6411
R5410 VDDA.t382 VDDA.t132 81.6411
R5411 VDDA.t368 VDDA.t382 81.6411
R5412 VDDA.t148 VDDA.t368 81.6411
R5413 VDDA.t14 VDDA.t148 81.6411
R5414 VDDA.t366 VDDA.t14 81.6411
R5415 VDDA.t275 VDDA.t366 81.6411
R5416 VDDA.n462 VDDA.n461 65.8183
R5417 VDDA.n461 VDDA.n448 65.8183
R5418 VDDA.n461 VDDA.n449 65.8183
R5419 VDDA.n447 VDDA.n426 65.8183
R5420 VDDA.n447 VDDA.n427 65.8183
R5421 VDDA.n447 VDDA.n428 65.8183
R5422 VDDA.n407 VDDA.n406 65.8183
R5423 VDDA.n406 VDDA.n325 65.8183
R5424 VDDA.n406 VDDA.n326 65.8183
R5425 VDDA.n406 VDDA.n327 65.8183
R5426 VDDA.n406 VDDA.n328 65.8183
R5427 VDDA.n377 VDDA.n330 65.8183
R5428 VDDA.n377 VDDA.n331 65.8183
R5429 VDDA.n377 VDDA.n332 65.8183
R5430 VDDA.n377 VDDA.n333 65.8183
R5431 VDDA.n377 VDDA.n334 65.8183
R5432 VDDA.n311 VDDA.n310 65.8183
R5433 VDDA.n311 VDDA.n302 65.8183
R5434 VDDA.n312 VDDA.n301 65.8183
R5435 VDDA.n277 VDDA.n276 65.8183
R5436 VDDA.n276 VDDA.n263 65.8183
R5437 VDDA.n276 VDDA.n264 65.8183
R5438 VDDA.n262 VDDA.n240 65.8183
R5439 VDDA.n262 VDDA.n241 65.8183
R5440 VDDA.n262 VDDA.n242 65.8183
R5441 VDDA.n229 VDDA.n228 65.8183
R5442 VDDA.n228 VDDA.n182 65.8183
R5443 VDDA.n221 VDDA.n220 65.8183
R5444 VDDA.n221 VDDA.n183 65.8183
R5445 VDDA.n199 VDDA.n191 65.8183
R5446 VDDA.n199 VDDA.n198 65.8183
R5447 VDDA.n172 VDDA.n171 65.8183
R5448 VDDA.n171 VDDA.n138 65.8183
R5449 VDDA.n171 VDDA.n139 65.8183
R5450 VDDA.n171 VDDA.n140 65.8183
R5451 VDDA.n171 VDDA.n141 65.8183
R5452 VDDA.n137 VDDA.n90 65.8183
R5453 VDDA.n137 VDDA.n91 65.8183
R5454 VDDA.n137 VDDA.n92 65.8183
R5455 VDDA.n137 VDDA.n93 65.8183
R5456 VDDA.n137 VDDA.n94 65.8183
R5457 VDDA.n74 VDDA.n73 65.8183
R5458 VDDA.n74 VDDA.n65 65.8183
R5459 VDDA.n81 VDDA.n75 65.8183
R5460 VDDA.n42 VDDA.n41 65.8183
R5461 VDDA.n41 VDDA.n28 65.8183
R5462 VDDA.n41 VDDA.n29 65.8183
R5463 VDDA.n27 VDDA.n5 65.8183
R5464 VDDA.n27 VDDA.n6 65.8183
R5465 VDDA.n27 VDDA.n7 65.8183
R5466 VDDA.n610 VDDA.n609 65.8183
R5467 VDDA.n610 VDDA.n600 65.8183
R5468 VDDA.n613 VDDA.n612 65.8183
R5469 VDDA.n588 VDDA.n587 65.8183
R5470 VDDA.n588 VDDA.n576 65.8183
R5471 VDDA.n575 VDDA.n537 65.8183
R5472 VDDA.n575 VDDA.n538 65.8183
R5473 VDDA.n666 VDDA.n665 65.8183
R5474 VDDA.n667 VDDA.n666 65.8183
R5475 VDDA.n660 VDDA.n627 65.8183
R5476 VDDA.n475 VDDA.t414 59.5681
R5477 VDDA.n474 VDDA.t415 59.5681
R5478 VDDA.n450 VDDA.n448 53.3664
R5479 VDDA.n454 VDDA.n449 53.3664
R5480 VDDA.n462 VDDA.n425 53.3664
R5481 VDDA.n455 VDDA.n448 53.3664
R5482 VDDA.n429 VDDA.n426 53.3664
R5483 VDDA.n435 VDDA.n427 53.3664
R5484 VDDA.n440 VDDA.n428 53.3664
R5485 VDDA.n434 VDDA.n426 53.3664
R5486 VDDA.n439 VDDA.n427 53.3664
R5487 VDDA.n378 VDDA.n325 53.3664
R5488 VDDA.n400 VDDA.n326 53.3664
R5489 VDDA.n396 VDDA.n327 53.3664
R5490 VDDA.n392 VDDA.n328 53.3664
R5491 VDDA.n407 VDDA.n324 53.3664
R5492 VDDA.n401 VDDA.n325 53.3664
R5493 VDDA.n397 VDDA.n326 53.3664
R5494 VDDA.n393 VDDA.n327 53.3664
R5495 VDDA.n389 VDDA.n328 53.3664
R5496 VDDA.n336 VDDA.n330 53.3664
R5497 VDDA.n370 VDDA.n331 53.3664
R5498 VDDA.n366 VDDA.n332 53.3664
R5499 VDDA.n362 VDDA.n333 53.3664
R5500 VDDA.n358 VDDA.n334 53.3664
R5501 VDDA.n371 VDDA.n330 53.3664
R5502 VDDA.n367 VDDA.n331 53.3664
R5503 VDDA.n363 VDDA.n332 53.3664
R5504 VDDA.n359 VDDA.n333 53.3664
R5505 VDDA.n355 VDDA.n334 53.3664
R5506 VDDA.n310 VDDA.n303 53.3664
R5507 VDDA.n305 VDDA.n302 53.3664
R5508 VDDA.n301 VDDA.n299 53.3664
R5509 VDDA.n301 VDDA.n300 53.3664
R5510 VDDA.n265 VDDA.n263 53.3664
R5511 VDDA.n269 VDDA.n264 53.3664
R5512 VDDA.n277 VDDA.n239 53.3664
R5513 VDDA.n270 VDDA.n263 53.3664
R5514 VDDA.n243 VDDA.n240 53.3664
R5515 VDDA.n251 VDDA.n241 53.3664
R5516 VDDA.n256 VDDA.n242 53.3664
R5517 VDDA.n250 VDDA.n240 53.3664
R5518 VDDA.n255 VDDA.n241 53.3664
R5519 VDDA.n211 VDDA.n183 53.3664
R5520 VDDA.n222 VDDA.n182 53.3664
R5521 VDDA.n229 VDDA.n181 53.3664
R5522 VDDA.n220 VDDA.n185 53.3664
R5523 VDDA.n191 VDDA.n190 53.3664
R5524 VDDA.n198 VDDA.n192 53.3664
R5525 VDDA.n194 VDDA.n191 53.3664
R5526 VDDA.n143 VDDA.n138 53.3664
R5527 VDDA.n165 VDDA.n139 53.3664
R5528 VDDA.n161 VDDA.n140 53.3664
R5529 VDDA.n157 VDDA.n141 53.3664
R5530 VDDA.n172 VDDA.n89 53.3664
R5531 VDDA.n166 VDDA.n138 53.3664
R5532 VDDA.n162 VDDA.n139 53.3664
R5533 VDDA.n158 VDDA.n140 53.3664
R5534 VDDA.n154 VDDA.n141 53.3664
R5535 VDDA.n96 VDDA.n90 53.3664
R5536 VDDA.n108 VDDA.n91 53.3664
R5537 VDDA.n111 VDDA.n92 53.3664
R5538 VDDA.n113 VDDA.n93 53.3664
R5539 VDDA.n117 VDDA.n94 53.3664
R5540 VDDA.n107 VDDA.n90 53.3664
R5541 VDDA.n110 VDDA.n91 53.3664
R5542 VDDA.n112 VDDA.n92 53.3664
R5543 VDDA.n116 VDDA.n93 53.3664
R5544 VDDA.n118 VDDA.n94 53.3664
R5545 VDDA.n73 VDDA.n66 53.3664
R5546 VDDA.n68 VDDA.n65 53.3664
R5547 VDDA.n75 VDDA.n64 53.3664
R5548 VDDA.n76 VDDA.n75 53.3664
R5549 VDDA.n30 VDDA.n28 53.3664
R5550 VDDA.n34 VDDA.n29 53.3664
R5551 VDDA.n42 VDDA.n4 53.3664
R5552 VDDA.n35 VDDA.n28 53.3664
R5553 VDDA.n8 VDDA.n5 53.3664
R5554 VDDA.n16 VDDA.n6 53.3664
R5555 VDDA.n21 VDDA.n7 53.3664
R5556 VDDA.n15 VDDA.n5 53.3664
R5557 VDDA.n20 VDDA.n6 53.3664
R5558 VDDA.n609 VDDA.n601 53.3664
R5559 VDDA.n605 VDDA.n600 53.3664
R5560 VDDA.n613 VDDA.n599 53.3664
R5561 VDDA.n614 VDDA.n613 53.3664
R5562 VDDA.n582 VDDA.n576 53.3664
R5563 VDDA.n587 VDDA.n578 53.3664
R5564 VDDA.n576 VDDA.n536 53.3664
R5565 VDDA.n540 VDDA.n537 53.3664
R5566 VDDA.n543 VDDA.n538 53.3664
R5567 VDDA.n542 VDDA.n537 53.3664
R5568 VDDA.n544 VDDA.n538 53.3664
R5569 VDDA.n665 VDDA.n661 53.3664
R5570 VDDA.n667 VDDA.n626 53.3664
R5571 VDDA.n629 VDDA.n627 53.3664
R5572 VDDA.n630 VDDA.n627 53.3664
R5573 VDDA.n474 VDDA.t413 52.3888
R5574 VDDA.n231 VDDA.n230 51.6576
R5575 VDDA.n202 VDDA.n201 51.6576
R5576 VDDA.n476 VDDA.t412 48.9557
R5577 VDDA.n207 VDDA.n206 48.0005
R5578 VDDA.n207 VDDA.n186 48.0005
R5579 VDDA.n419 VDDA.n418 46.6291
R5580 VDDA.n417 VDDA.n416 46.6291
R5581 VDDA.n478 VDDA.t160 39.4005
R5582 VDDA.n478 VDDA.t7 39.4005
R5583 VDDA.n508 VDDA.t29 39.4005
R5584 VDDA.n508 VDDA.t313 39.4005
R5585 VDDA.n510 VDDA.t403 39.4005
R5586 VDDA.n510 VDDA.t299 39.4005
R5587 VDDA.n512 VDDA.t311 39.4005
R5588 VDDA.n512 VDDA.t81 39.4005
R5589 VDDA.n514 VDDA.t110 39.4005
R5590 VDDA.n514 VDDA.t44 39.4005
R5591 VDDA.n516 VDDA.t293 39.4005
R5592 VDDA.n516 VDDA.t93 39.4005
R5593 VDDA.n518 VDDA.t66 39.4005
R5594 VDDA.n518 VDDA.t34 39.4005
R5595 VDDA.n520 VDDA.t96 39.4005
R5596 VDDA.n520 VDDA.t5 39.4005
R5597 VDDA.n522 VDDA.t376 39.4005
R5598 VDDA.n522 VDDA.t163 39.4005
R5599 VDDA.n483 VDDA.t173 39.4005
R5600 VDDA.n483 VDDA.t394 39.4005
R5601 VDDA.n486 VDDA.t297 39.4005
R5602 VDDA.n486 VDDA.t38 39.4005
R5603 VDDA.n488 VDDA.t165 39.4005
R5604 VDDA.n488 VDDA.t9 39.4005
R5605 VDDA.n490 VDDA.t175 39.4005
R5606 VDDA.n490 VDDA.t98 39.4005
R5607 VDDA.n492 VDDA.t363 39.4005
R5608 VDDA.n492 VDDA.t135 39.4005
R5609 VDDA.n494 VDDA.t373 39.4005
R5610 VDDA.n494 VDDA.t137 39.4005
R5611 VDDA.n496 VDDA.t40 39.4005
R5612 VDDA.n496 VDDA.t371 39.4005
R5613 VDDA.n498 VDDA.t60 39.4005
R5614 VDDA.n498 VDDA.t108 39.4005
R5615 VDDA.n500 VDDA.t144 39.4005
R5616 VDDA.n500 VDDA.t125 39.4005
R5617 VDDA.n621 VDDA.t315 39.4005
R5618 VDDA.n621 VDDA.t365 39.4005
R5619 VDDA.n671 VDDA.t86 39.4005
R5620 VDDA.n671 VDDA.t2 39.4005
R5621 VDDA.n631 VDDA.t58 39.4005
R5622 VDDA.n631 VDDA.t27 39.4005
R5623 VDDA.n640 VDDA.t23 39.4005
R5624 VDDA.n640 VDDA.t21 39.4005
R5625 VDDA.n633 VDDA.t301 39.4005
R5626 VDDA.n633 VDDA.t410 39.4005
R5627 VDDA.n473 VDDA.n467 27.9413
R5628 VDDA.n677 VDDA.n676 27.2462
R5629 VDDA.n675 VDDA.n674 27.2462
R5630 VDDA.n646 VDDA.n645 27.2462
R5631 VDDA.n644 VDDA.n643 27.2462
R5632 VDDA.n638 VDDA.n637 27.2462
R5633 VDDA.n636 VDDA.n635 27.2462
R5634 VDDA.n547 VDDA.n546 22.9536
R5635 VDDA.n506 VDDA.n505 22.9536
R5636 VDDA.n464 VDDA.n463 22.8576
R5637 VDDA.n445 VDDA.n430 22.8576
R5638 VDDA.n409 VDDA.n408 22.8576
R5639 VDDA.n375 VDDA.n345 22.8576
R5640 VDDA.n319 VDDA.n318 22.8576
R5641 VDDA.n279 VDDA.n278 22.8576
R5642 VDDA.n260 VDDA.n246 22.8576
R5643 VDDA.n174 VDDA.n173 22.8576
R5644 VDDA.n135 VDDA.n105 22.8576
R5645 VDDA.n84 VDDA.n83 22.8576
R5646 VDDA.n44 VDDA.n43 22.8576
R5647 VDDA.n25 VDDA.n11 22.8576
R5648 VDDA.n604 VDDA.n603 22.8576
R5649 VDDA.n596 VDDA.n595 22.8576
R5650 VDDA.n591 VDDA.n590 22.8576
R5651 VDDA.n567 VDDA.n566 22.8576
R5652 VDDA.n669 VDDA.n668 22.8576
R5653 VDDA.n654 VDDA.n653 22.8576
R5654 VDDA.n414 VDDA.t146 21.8894
R5655 VDDA.n414 VDDA.t227 21.8894
R5656 VDDA.n467 VDDA.n466 20.883
R5657 VDDA.n530 VDDA.n480 20.7243
R5658 VDDA.n525 VDDA.n482 20.7243
R5659 VDDA.n502 VDDA.n485 20.7243
R5660 VDDA.n549 VDDA.n548 20.4312
R5661 VDDA.n473 VDDA.t105 19.9244
R5662 VDDA.n617 VDDA.t270 19.7005
R5663 VDDA.n617 VDDA.t42 19.7005
R5664 VDDA.n623 VDDA.t31 19.7005
R5665 VDDA.n623 VDDA.t208 19.7005
R5666 VDDA.n648 VDDA.t25 19.7005
R5667 VDDA.n648 VDDA.t303 19.7005
R5668 VDDA.n650 VDDA.t285 19.7005
R5669 VDDA.n650 VDDA.t379 19.7005
R5670 VDDA.n320 VDDA.n319 19.613
R5671 VDDA.n85 VDDA.n84 19.613
R5672 VDDA.n177 VDDA.t381 15.7605
R5673 VDDA.n177 VDDA.t158 15.7605
R5674 VDDA.n203 VDDA.t19 15.7605
R5675 VDDA.n203 VDDA.t309 15.7605
R5676 VDDA.n215 VDDA.t240 15.7605
R5677 VDDA.n218 VDDA.t212 15.7605
R5678 VDDA.n179 VDDA.t288 15.7605
R5679 VDDA.n188 VDDA.t243 15.7605
R5680 VDDA.n550 VDDA.n546 15.488
R5681 VDDA.n204 VDDA.n202 14.7224
R5682 VDDA.n502 VDDA.n501 14.6963
R5683 VDDA.n281 VDDA.n279 14.4255
R5684 VDDA.n246 VDDA.n245 14.4255
R5685 VDDA.n46 VDDA.n44 14.4255
R5686 VDDA.n11 VDDA.n10 14.4255
R5687 VDDA.n345 VDDA.n344 14.363
R5688 VDDA.n105 VDDA.n104 14.363
R5689 VDDA.n603 VDDA.n593 14.363
R5690 VDDA.n635 VDDA.n634 14.2693
R5691 VDDA.n550 VDDA.n549 14.238
R5692 VDDA.n595 VDDA.n593 14.0818
R5693 VDDA.n525 VDDA.n524 14.0713
R5694 VDDA.n531 VDDA.n530 14.0713
R5695 VDDA.n507 VDDA.n506 14.0713
R5696 VDDA.n430 VDDA.n422 14.0505
R5697 VDDA.n416 VDDA.n415 14.0505
R5698 VDDA.n465 VDDA.n464 13.8005
R5699 VDDA.n420 VDDA.n419 13.8005
R5700 VDDA.n410 VDDA.n409 13.8005
R5701 VDDA.n206 VDDA.n205 13.8005
R5702 VDDA.n187 VDDA.n186 13.8005
R5703 VDDA.n232 VDDA.n231 13.8005
R5704 VDDA.n175 VDDA.n174 13.8005
R5705 VDDA.n566 VDDA.n565 13.8005
R5706 VDDA.n592 VDDA.n591 13.8005
R5707 VDDA.n674 VDDA.n673 13.8005
R5708 VDDA.n653 VDDA.n652 13.8005
R5709 VDDA.n643 VDDA.n642 13.8005
R5710 VDDA.n639 VDDA.n638 13.8005
R5711 VDDA.n647 VDDA.n646 13.8005
R5712 VDDA.n670 VDDA.n669 13.8005
R5713 VDDA.n678 VDDA.n677 13.8005
R5714 VDDA.n533 VDDA.t69 13.1338
R5715 VDDA.n533 VDDA.t100 13.1338
R5716 VDDA.n551 VDDA.t103 13.1338
R5717 VDDA.n551 VDDA.t11 13.1338
R5718 VDDA.n553 VDDA.t74 13.1338
R5719 VDDA.n553 VDDA.t76 13.1338
R5720 VDDA.n555 VDDA.t91 13.1338
R5721 VDDA.n555 VDDA.t51 13.1338
R5722 VDDA.n557 VDDA.t49 13.1338
R5723 VDDA.n557 VDDA.t83 13.1338
R5724 VDDA.n559 VDDA.t89 13.1338
R5725 VDDA.n559 VDDA.t72 13.1338
R5726 VDDA.n561 VDDA.t154 13.1338
R5727 VDDA.n561 VDDA.t168 13.1338
R5728 VDDA.n563 VDDA.t53 13.1338
R5729 VDDA.n563 VDDA.t305 13.1338
R5730 VDDA.n679 VDDA.n678 11.4105
R5731 VDDA.t234 VDDA.n443 11.2576
R5732 VDDA.n443 VDDA.t349 11.2576
R5733 VDDA.n444 VDDA.t234 11.2576
R5734 VDDA.n423 VDDA.t282 11.2576
R5735 VDDA.n285 VDDA.t357 11.2576
R5736 VDDA.n285 VDDA.t321 11.2576
R5737 VDDA.n235 VDDA.t345 11.2576
R5738 VDDA.n235 VDDA.t353 11.2576
R5739 VDDA.n244 VDDA.t327 11.2576
R5740 VDDA.n244 VDDA.t337 11.2576
R5741 VDDA.n259 VDDA.t181 11.2576
R5742 VDDA.n237 VDDA.t237 11.2576
R5743 VDDA.n280 VDDA.t335 11.2576
R5744 VDDA.n280 VDDA.t343 11.2576
R5745 VDDA.n282 VDDA.t331 11.2576
R5746 VDDA.n282 VDDA.t339 11.2576
R5747 VDDA.n50 VDDA.t325 11.2576
R5748 VDDA.n50 VDDA.t333 11.2576
R5749 VDDA.n0 VDDA.t319 11.2576
R5750 VDDA.n0 VDDA.t329 11.2576
R5751 VDDA.n9 VDDA.t351 11.2576
R5752 VDDA.n9 VDDA.t355 11.2576
R5753 VDDA.n24 VDDA.t252 11.2576
R5754 VDDA.n2 VDDA.t196 11.2576
R5755 VDDA.n45 VDDA.t323 11.2576
R5756 VDDA.n45 VDDA.t317 11.2576
R5757 VDDA.n47 VDDA.t341 11.2576
R5758 VDDA.n47 VDDA.t347 11.2576
R5759 VDDA.n477 VDDA.n476 11.1572
R5760 VDDA.n320 VDDA.n297 10.8443
R5761 VDDA.n85 VDDA.n62 10.8443
R5762 VDDA.n620 VDDA.n619 9.7855
R5763 VDDA.n463 VDDA.n424 9.14336
R5764 VDDA.n459 VDDA.n458 9.14336
R5765 VDDA.n456 VDDA.n453 9.14336
R5766 VDDA.n445 VDDA.n431 9.14336
R5767 VDDA.n436 VDDA.n433 9.14336
R5768 VDDA.n441 VDDA.n438 9.14336
R5769 VDDA.n404 VDDA.n379 9.14336
R5770 VDDA.n404 VDDA.n403 9.14336
R5771 VDDA.n403 VDDA.n402 9.14336
R5772 VDDA.n402 VDDA.n399 9.14336
R5773 VDDA.n399 VDDA.n398 9.14336
R5774 VDDA.n398 VDDA.n395 9.14336
R5775 VDDA.n395 VDDA.n394 9.14336
R5776 VDDA.n394 VDDA.n391 9.14336
R5777 VDDA.n391 VDDA.n390 9.14336
R5778 VDDA.n372 VDDA.n346 9.14336
R5779 VDDA.n372 VDDA.n369 9.14336
R5780 VDDA.n369 VDDA.n368 9.14336
R5781 VDDA.n368 VDDA.n365 9.14336
R5782 VDDA.n365 VDDA.n364 9.14336
R5783 VDDA.n364 VDDA.n361 9.14336
R5784 VDDA.n361 VDDA.n360 9.14336
R5785 VDDA.n360 VDDA.n357 9.14336
R5786 VDDA.n357 VDDA.n356 9.14336
R5787 VDDA.n306 VDDA.n304 9.14336
R5788 VDDA.n316 VDDA.n315 9.14336
R5789 VDDA.n278 VDDA.n238 9.14336
R5790 VDDA.n274 VDDA.n273 9.14336
R5791 VDDA.n271 VDDA.n268 9.14336
R5792 VDDA.n260 VDDA.n247 9.14336
R5793 VDDA.n252 VDDA.n249 9.14336
R5794 VDDA.n257 VDDA.n254 9.14336
R5795 VDDA.n230 VDDA.n180 9.14336
R5796 VDDA.n226 VDDA.n225 9.14336
R5797 VDDA.n201 VDDA.n189 9.14336
R5798 VDDA.n196 VDDA.n195 9.14336
R5799 VDDA.n169 VDDA.n144 9.14336
R5800 VDDA.n169 VDDA.n168 9.14336
R5801 VDDA.n168 VDDA.n167 9.14336
R5802 VDDA.n167 VDDA.n164 9.14336
R5803 VDDA.n164 VDDA.n163 9.14336
R5804 VDDA.n163 VDDA.n160 9.14336
R5805 VDDA.n160 VDDA.n159 9.14336
R5806 VDDA.n159 VDDA.n156 9.14336
R5807 VDDA.n156 VDDA.n155 9.14336
R5808 VDDA.n133 VDDA.n132 9.14336
R5809 VDDA.n132 VDDA.n131 9.14336
R5810 VDDA.n131 VDDA.n109 9.14336
R5811 VDDA.n127 VDDA.n109 9.14336
R5812 VDDA.n127 VDDA.n126 9.14336
R5813 VDDA.n126 VDDA.n114 9.14336
R5814 VDDA.n122 VDDA.n114 9.14336
R5815 VDDA.n122 VDDA.n121 9.14336
R5816 VDDA.n121 VDDA.n120 9.14336
R5817 VDDA.n69 VDDA.n67 9.14336
R5818 VDDA.n78 VDDA.n77 9.14336
R5819 VDDA.n43 VDDA.n3 9.14336
R5820 VDDA.n39 VDDA.n38 9.14336
R5821 VDDA.n36 VDDA.n33 9.14336
R5822 VDDA.n25 VDDA.n12 9.14336
R5823 VDDA.n17 VDDA.n14 9.14336
R5824 VDDA.n22 VDDA.n19 9.14336
R5825 VDDA.n606 VDDA.n602 9.14336
R5826 VDDA.n615 VDDA.n597 9.14336
R5827 VDDA.n584 VDDA.n579 9.14336
R5828 VDDA.n584 VDDA.n583 9.14336
R5829 VDDA.n583 VDDA.n581 9.14336
R5830 VDDA.n572 VDDA.n571 9.14336
R5831 VDDA.n571 VDDA.n570 9.14336
R5832 VDDA.n570 VDDA.n545 9.14336
R5833 VDDA.n663 VDDA.n662 9.14336
R5834 VDDA.n657 VDDA.n656 9.14336
R5835 VDDA.n532 VDDA.n531 8.973
R5836 VDDA.n412 VDDA.n411 8.8755
R5837 VDDA.n233 VDDA.n232 8.688
R5838 VDDA.n234 VDDA.n233 8.28175
R5839 VDDA.n412 VDDA.n286 8.15675
R5840 VDDA.n234 VDDA.n51 8.15675
R5841 VDDA.n296 VDDA.t361 8.0005
R5842 VDDA.n296 VDDA.t170 8.0005
R5843 VDDA.n294 VDDA.t84 8.0005
R5844 VDDA.n294 VDDA.t390 8.0005
R5845 VDDA.n292 VDDA.t94 8.0005
R5846 VDDA.n292 VDDA.t391 8.0005
R5847 VDDA.n290 VDDA.t106 8.0005
R5848 VDDA.n290 VDDA.t139 8.0005
R5849 VDDA.n288 VDDA.t401 8.0005
R5850 VDDA.n288 VDDA.t121 8.0005
R5851 VDDA.n287 VDDA.t377 8.0005
R5852 VDDA.n287 VDDA.t358 8.0005
R5853 VDDA.n61 VDDA.t147 8.0005
R5854 VDDA.n61 VDDA.t360 8.0005
R5855 VDDA.n59 VDDA.t32 8.0005
R5856 VDDA.n59 VDDA.t63 8.0005
R5857 VDDA.n57 VDDA.t374 8.0005
R5858 VDDA.n57 VDDA.t127 8.0005
R5859 VDDA.n55 VDDA.t117 8.0005
R5860 VDDA.n55 VDDA.t126 8.0005
R5861 VDDA.n53 VDDA.t112 8.0005
R5862 VDDA.n53 VDDA.t389 8.0005
R5863 VDDA.n52 VDDA.t359 8.0005
R5864 VDDA.n52 VDDA.t78 8.0005
R5865 VDDA.n321 VDDA.t17 6.56717
R5866 VDDA.n321 VDDA.t114 6.56717
R5867 VDDA.n337 VDDA.t129 6.56717
R5868 VDDA.n337 VDDA.t400 6.56717
R5869 VDDA.n339 VDDA.t55 6.56717
R5870 VDDA.n339 VDDA.t119 6.56717
R5871 VDDA.n341 VDDA.t142 6.56717
R5872 VDDA.n341 VDDA.t36 6.56717
R5873 VDDA.n343 VDDA.t408 6.56717
R5874 VDDA.n343 VDDA.t123 6.56717
R5875 VDDA.n86 VDDA.t15 6.56717
R5876 VDDA.n86 VDDA.t367 6.56717
R5877 VDDA.n97 VDDA.t369 6.56717
R5878 VDDA.n97 VDDA.t149 6.56717
R5879 VDDA.n99 VDDA.t133 6.56717
R5880 VDDA.n99 VDDA.t383 6.56717
R5881 VDDA.n101 VDDA.t385 6.56717
R5882 VDDA.n101 VDDA.t388 6.56717
R5883 VDDA.n103 VDDA.t62 6.56717
R5884 VDDA.n103 VDDA.t397 6.56717
R5885 VDDA.n421 VDDA.n413 6.563
R5886 VDDA.n413 VDDA.n412 6.5005
R5887 VDDA.n413 VDDA.n234 6.5005
R5888 VDDA.n411 VDDA.n410 5.8755
R5889 VDDA.n176 VDDA.n175 5.8755
R5890 VDDA.n408 VDDA.n323 5.33286
R5891 VDDA.n375 VDDA.n374 5.33286
R5892 VDDA.n318 VDDA.n317 5.33286
R5893 VDDA.n309 VDDA.n308 5.33286
R5894 VDDA.n135 VDDA.n134 5.33286
R5895 VDDA.n173 VDDA.n88 5.33286
R5896 VDDA.n72 VDDA.n71 5.33286
R5897 VDDA.n83 VDDA.n63 5.33286
R5898 VDDA.n607 VDDA.n604 5.33286
R5899 VDDA.n616 VDDA.n596 5.33286
R5900 VDDA.n590 VDDA.n535 5.33286
R5901 VDDA.n568 VDDA.n567 5.33286
R5902 VDDA.n668 VDDA.n625 5.33286
R5903 VDDA.n655 VDDA.n654 5.33286
R5904 VDDA.n466 VDDA.n465 5.28175
R5905 VDDA.n421 VDDA.n420 5.28175
R5906 VDDA.n411 VDDA.n320 4.96925
R5907 VDDA.n176 VDDA.n85 4.96925
R5908 VDDA.n619 VDDA.n618 4.7505
R5909 VDDA.n477 VDDA.n473 4.5595
R5910 VDDA.n481 VDDA.n480 4.54311
R5911 VDDA.n529 VDDA.n481 4.54311
R5912 VDDA.n451 VDDA.n424 4.53698
R5913 VDDA.n458 VDDA.n457 4.53698
R5914 VDDA.n453 VDDA.n452 4.53698
R5915 VDDA.n459 VDDA.n451 4.53698
R5916 VDDA.n457 VDDA.n456 4.53698
R5917 VDDA.n432 VDDA.n431 4.53698
R5918 VDDA.n437 VDDA.n436 4.53698
R5919 VDDA.n442 VDDA.n441 4.53698
R5920 VDDA.n433 VDDA.n432 4.53698
R5921 VDDA.n438 VDDA.n437 4.53698
R5922 VDDA.n266 VDDA.n238 4.53698
R5923 VDDA.n273 VDDA.n272 4.53698
R5924 VDDA.n268 VDDA.n267 4.53698
R5925 VDDA.n274 VDDA.n266 4.53698
R5926 VDDA.n272 VDDA.n271 4.53698
R5927 VDDA.n248 VDDA.n247 4.53698
R5928 VDDA.n253 VDDA.n252 4.53698
R5929 VDDA.n258 VDDA.n257 4.53698
R5930 VDDA.n249 VDDA.n248 4.53698
R5931 VDDA.n254 VDDA.n253 4.53698
R5932 VDDA.n223 VDDA.n180 4.53698
R5933 VDDA.n225 VDDA.n224 4.53698
R5934 VDDA.n226 VDDA.n223 4.53698
R5935 VDDA.n193 VDDA.n189 4.53698
R5936 VDDA.n197 VDDA.n196 4.53698
R5937 VDDA.n195 VDDA.n193 4.53698
R5938 VDDA.n31 VDDA.n3 4.53698
R5939 VDDA.n38 VDDA.n37 4.53698
R5940 VDDA.n33 VDDA.n32 4.53698
R5941 VDDA.n39 VDDA.n31 4.53698
R5942 VDDA.n37 VDDA.n36 4.53698
R5943 VDDA.n13 VDDA.n12 4.53698
R5944 VDDA.n18 VDDA.n17 4.53698
R5945 VDDA.n23 VDDA.n22 4.53698
R5946 VDDA.n14 VDDA.n13 4.53698
R5947 VDDA.n19 VDDA.n18 4.53698
R5948 VDDA.n286 VDDA.n284 4.5005
R5949 VDDA.n51 VDDA.n49 4.5005
R5950 VDDA.n618 VDDA.n593 4.5005
R5951 VDDA.n527 VDDA.n482 4.48641
R5952 VDDA.n527 VDDA.n526 4.48641
R5953 VDDA.n504 VDDA.n485 4.48641
R5954 VDDA.n504 VDDA.n503 4.48641
R5955 VDDA.n475 VDDA.n474 4.12334
R5956 VDDA.n379 VDDA.n323 3.75335
R5957 VDDA.n390 VDDA.n388 3.75335
R5958 VDDA.n374 VDDA.n346 3.75335
R5959 VDDA.n356 VDDA.n354 3.75335
R5960 VDDA.n308 VDDA.n304 3.75335
R5961 VDDA.n307 VDDA.n306 3.75335
R5962 VDDA.n317 VDDA.n316 3.75335
R5963 VDDA.n315 VDDA.n314 3.75335
R5964 VDDA.n144 VDDA.n88 3.75335
R5965 VDDA.n155 VDDA.n153 3.75335
R5966 VDDA.n134 VDDA.n133 3.75335
R5967 VDDA.n120 VDDA.n119 3.75335
R5968 VDDA.n71 VDDA.n67 3.75335
R5969 VDDA.n70 VDDA.n69 3.75335
R5970 VDDA.n77 VDDA.n63 3.75335
R5971 VDDA.n79 VDDA.n78 3.75335
R5972 VDDA.n608 VDDA.n602 3.75335
R5973 VDDA.n607 VDDA.n606 3.75335
R5974 VDDA.n597 VDDA.n594 3.75335
R5975 VDDA.n616 VDDA.n615 3.75335
R5976 VDDA.n586 VDDA.n579 3.75335
R5977 VDDA.n581 VDDA.n535 3.75335
R5978 VDDA.n573 VDDA.n572 3.75335
R5979 VDDA.n568 VDDA.n545 3.75335
R5980 VDDA.n664 VDDA.n663 3.75335
R5981 VDDA.n662 VDDA.n625 3.75335
R5982 VDDA.n658 VDDA.n657 3.75335
R5983 VDDA.n656 VDDA.n655 3.75335
R5984 VDDA.n680 VDDA.n679 3.71013
R5985 VDDA.n476 VDDA.n475 3.43377
R5986 VDDA.n209 VDDA.n208 2.8957
R5987 VDDA.n210 VDDA.n209 2.8957
R5988 VDDA.n214 VDDA.n212 2.8957
R5989 VDDA.n217 VDDA.n212 2.8957
R5990 VDDA.n213 VDDA.n210 2.8957
R5991 VDDA.n217 VDDA.n216 2.8957
R5992 VDDA.n219 VDDA.n208 2.8957
R5993 VDDA.n214 VDDA.n213 2.8957
R5994 VDDA.n652 VDDA.n647 2.78175
R5995 VDDA.n673 VDDA.n670 2.78175
R5996 VDDA.n619 VDDA.n592 2.5005
R5997 VDDA.n219 VDDA.n207 2.32777
R5998 VDDA.n680 VDDA.n467 2.1343
R5999 VDDA VDDA.n680 2.0779
R6000 VDDA.n642 VDDA.n639 2.063
R6001 VDDA.n524 VDDA.n507 1.8755
R6002 VDDA.n565 VDDA.n550 1.84425
R6003 VDDA.n565 VDDA.n564 1.0005
R6004 VDDA.n564 VDDA.n562 1.0005
R6005 VDDA.n562 VDDA.n560 1.0005
R6006 VDDA.n560 VDDA.n558 1.0005
R6007 VDDA.n558 VDDA.n556 1.0005
R6008 VDDA.n556 VDDA.n554 1.0005
R6009 VDDA.n554 VDDA.n552 1.0005
R6010 VDDA.n552 VDDA.n534 1.0005
R6011 VDDA.n592 VDDA.n534 1.0005
R6012 VDDA.n466 VDDA.n421 0.938
R6013 VDDA.n205 VDDA.n204 0.922375
R6014 VDDA.n187 VDDA.n178 0.922375
R6015 VDDA.n232 VDDA.n178 0.922375
R6016 VDDA.n532 VDDA.n477 0.840625
R6017 VDDA.n620 VDDA.n532 0.74075
R6018 VDDA.n639 VDDA.n634 0.65675
R6019 VDDA.n465 VDDA.n422 0.6255
R6020 VDDA.n420 VDDA.n415 0.6255
R6021 VDDA.n284 VDDA.n283 0.6255
R6022 VDDA.n283 VDDA.n281 0.6255
R6023 VDDA.n245 VDDA.n236 0.6255
R6024 VDDA.n284 VDDA.n236 0.6255
R6025 VDDA.n49 VDDA.n48 0.6255
R6026 VDDA.n48 VDDA.n46 0.6255
R6027 VDDA.n10 VDDA.n1 0.6255
R6028 VDDA.n49 VDDA.n1 0.6255
R6029 VDDA.n501 VDDA.n499 0.6255
R6030 VDDA.n499 VDDA.n497 0.6255
R6031 VDDA.n497 VDDA.n495 0.6255
R6032 VDDA.n495 VDDA.n493 0.6255
R6033 VDDA.n493 VDDA.n491 0.6255
R6034 VDDA.n491 VDDA.n489 0.6255
R6035 VDDA.n489 VDDA.n487 0.6255
R6036 VDDA.n487 VDDA.n484 0.6255
R6037 VDDA.n507 VDDA.n484 0.6255
R6038 VDDA.n524 VDDA.n523 0.6255
R6039 VDDA.n523 VDDA.n521 0.6255
R6040 VDDA.n521 VDDA.n519 0.6255
R6041 VDDA.n519 VDDA.n517 0.6255
R6042 VDDA.n517 VDDA.n515 0.6255
R6043 VDDA.n515 VDDA.n513 0.6255
R6044 VDDA.n513 VDDA.n511 0.6255
R6045 VDDA.n511 VDDA.n509 0.6255
R6046 VDDA.n509 VDDA.n479 0.6255
R6047 VDDA.n531 VDDA.n479 0.6255
R6048 VDDA.n344 VDDA.n342 0.563
R6049 VDDA.n342 VDDA.n340 0.563
R6050 VDDA.n340 VDDA.n338 0.563
R6051 VDDA.n338 VDDA.n322 0.563
R6052 VDDA.n410 VDDA.n322 0.563
R6053 VDDA.n291 VDDA.n289 0.563
R6054 VDDA.n293 VDDA.n291 0.563
R6055 VDDA.n295 VDDA.n293 0.563
R6056 VDDA.n297 VDDA.n295 0.563
R6057 VDDA.n104 VDDA.n102 0.563
R6058 VDDA.n102 VDDA.n100 0.563
R6059 VDDA.n100 VDDA.n98 0.563
R6060 VDDA.n98 VDDA.n87 0.563
R6061 VDDA.n175 VDDA.n87 0.563
R6062 VDDA.n56 VDDA.n54 0.563
R6063 VDDA.n58 VDDA.n56 0.563
R6064 VDDA.n60 VDDA.n58 0.563
R6065 VDDA.n62 VDDA.n60 0.563
R6066 VDDA.n642 VDDA.n641 0.563
R6067 VDDA.n641 VDDA.n632 0.563
R6068 VDDA.n647 VDDA.n632 0.563
R6069 VDDA.n651 VDDA.n649 0.563
R6070 VDDA.n649 VDDA.n624 0.563
R6071 VDDA.n673 VDDA.n672 0.563
R6072 VDDA.n672 VDDA.n622 0.563
R6073 VDDA.n678 VDDA.n622 0.563
R6074 VDDA.n233 VDDA.n176 0.46925
R6075 VDDA VDDA.n620 0.41175
R6076 VDDA.n205 VDDA.n187 0.3755
R6077 VDDA.n652 VDDA.n651 0.28175
R6078 VDDA.n670 VDDA.n624 0.28175
R6079 VDDA.t169 VDDA.t104 0.1603
R6080 VDDA.t152 VDDA.t77 0.1603
R6081 VDDA.t101 VDDA.t45 0.1603
R6082 VDDA.t70 VDDA.t156 0.1603
R6083 VDDA.t13 VDDA.t306 0.1603
R6084 VDDA.n469 VDDA.t307 0.159278
R6085 VDDA.n470 VDDA.t150 0.159278
R6086 VDDA.n471 VDDA.t47 0.159278
R6087 VDDA.n472 VDDA.t155 0.159278
R6088 VDDA.n472 VDDA.t12 0.1368
R6089 VDDA.n472 VDDA.t169 0.1368
R6090 VDDA.n471 VDDA.t46 0.1368
R6091 VDDA.n471 VDDA.t152 0.1368
R6092 VDDA.n470 VDDA.t87 0.1368
R6093 VDDA.n470 VDDA.t101 0.1368
R6094 VDDA.n469 VDDA.t166 0.1368
R6095 VDDA.n469 VDDA.t70 0.1368
R6096 VDDA.n468 VDDA.t151 0.1368
R6097 VDDA.n468 VDDA.t13 0.1368
R6098 VDDA.n679 VDDA 0.135625
R6099 VDDA.t307 VDDA.n468 0.00152174
R6100 VDDA.t150 VDDA.n469 0.00152174
R6101 VDDA.t47 VDDA.n470 0.00152174
R6102 VDDA.t155 VDDA.n471 0.00152174
R6103 VDDA.t105 VDDA.n472 0.00152174
R6104 bgr_7_0.V_TOP.n0 bgr_7_0.V_TOP.t29 369.534
R6105 bgr_7_0.V_TOP.n23 bgr_7_0.V_TOP.n21 339.961
R6106 bgr_7_0.V_TOP.n23 bgr_7_0.V_TOP.n22 339.272
R6107 bgr_7_0.V_TOP.n19 bgr_7_0.V_TOP.n18 339.272
R6108 bgr_7_0.V_TOP.n27 bgr_7_0.V_TOP.n26 339.272
R6109 bgr_7_0.V_TOP.n29 bgr_7_0.V_TOP.n28 339.272
R6110 bgr_7_0.V_TOP.n24 bgr_7_0.V_TOP.n20 334.772
R6111 bgr_7_0.V_TOP.n39 bgr_7_0.V_TOP.n38 224.934
R6112 bgr_7_0.V_TOP.n38 bgr_7_0.V_TOP.n37 224.934
R6113 bgr_7_0.V_TOP.n37 bgr_7_0.V_TOP.n36 224.934
R6114 bgr_7_0.V_TOP.n36 bgr_7_0.V_TOP.n35 224.934
R6115 bgr_7_0.V_TOP.n35 bgr_7_0.V_TOP.n34 224.934
R6116 bgr_7_0.V_TOP.n34 bgr_7_0.V_TOP.n33 224.934
R6117 bgr_7_0.V_TOP.n33 bgr_7_0.V_TOP.n32 224.934
R6118 bgr_7_0.V_TOP.n1 bgr_7_0.V_TOP.n0 224.934
R6119 bgr_7_0.V_TOP.n2 bgr_7_0.V_TOP.n1 224.934
R6120 bgr_7_0.V_TOP.n3 bgr_7_0.V_TOP.n2 224.934
R6121 bgr_7_0.V_TOP.n4 bgr_7_0.V_TOP.n3 224.934
R6122 bgr_7_0.V_TOP.n5 bgr_7_0.V_TOP.n4 224.934
R6123 bgr_7_0.V_TOP bgr_7_0.V_TOP.t48 214.222
R6124 bgr_7_0.V_TOP.n31 bgr_7_0.V_TOP.n30 163.175
R6125 bgr_7_0.V_TOP.n39 bgr_7_0.V_TOP.t24 144.601
R6126 bgr_7_0.V_TOP.n38 bgr_7_0.V_TOP.t33 144.601
R6127 bgr_7_0.V_TOP.n37 bgr_7_0.V_TOP.t39 144.601
R6128 bgr_7_0.V_TOP.n36 bgr_7_0.V_TOP.t16 144.601
R6129 bgr_7_0.V_TOP.n35 bgr_7_0.V_TOP.t15 144.601
R6130 bgr_7_0.V_TOP.n34 bgr_7_0.V_TOP.t28 144.601
R6131 bgr_7_0.V_TOP.n33 bgr_7_0.V_TOP.t38 144.601
R6132 bgr_7_0.V_TOP.n32 bgr_7_0.V_TOP.t14 144.601
R6133 bgr_7_0.V_TOP.n0 bgr_7_0.V_TOP.t30 144.601
R6134 bgr_7_0.V_TOP.n1 bgr_7_0.V_TOP.t18 144.601
R6135 bgr_7_0.V_TOP.n2 bgr_7_0.V_TOP.t46 144.601
R6136 bgr_7_0.V_TOP.n3 bgr_7_0.V_TOP.t37 144.601
R6137 bgr_7_0.V_TOP.n4 bgr_7_0.V_TOP.t26 144.601
R6138 bgr_7_0.V_TOP.n5 bgr_7_0.V_TOP.t27 144.601
R6139 bgr_7_0.V_TOP.n17 bgr_7_0.V_TOP.t0 108.424
R6140 bgr_7_0.V_TOP.n30 bgr_7_0.V_TOP.t10 95.4467
R6141 bgr_7_0.V_TOP bgr_7_0.V_TOP.n39 69.6227
R6142 bgr_7_0.V_TOP.n32 bgr_7_0.V_TOP.n31 69.6227
R6143 bgr_7_0.V_TOP.n31 bgr_7_0.V_TOP.n5 69.6227
R6144 bgr_7_0.V_TOP.n18 bgr_7_0.V_TOP.t6 39.4005
R6145 bgr_7_0.V_TOP.n18 bgr_7_0.V_TOP.t3 39.4005
R6146 bgr_7_0.V_TOP.n20 bgr_7_0.V_TOP.t11 39.4005
R6147 bgr_7_0.V_TOP.n20 bgr_7_0.V_TOP.t12 39.4005
R6148 bgr_7_0.V_TOP.n22 bgr_7_0.V_TOP.t4 39.4005
R6149 bgr_7_0.V_TOP.n22 bgr_7_0.V_TOP.t9 39.4005
R6150 bgr_7_0.V_TOP.n21 bgr_7_0.V_TOP.t8 39.4005
R6151 bgr_7_0.V_TOP.n21 bgr_7_0.V_TOP.t2 39.4005
R6152 bgr_7_0.V_TOP.n26 bgr_7_0.V_TOP.t1 39.4005
R6153 bgr_7_0.V_TOP.n26 bgr_7_0.V_TOP.t5 39.4005
R6154 bgr_7_0.V_TOP.n28 bgr_7_0.V_TOP.t13 39.4005
R6155 bgr_7_0.V_TOP.n28 bgr_7_0.V_TOP.t7 39.4005
R6156 bgr_7_0.V_TOP.n17 bgr_7_0.V_TOP.n16 37.1479
R6157 bgr_7_0.V_TOP.n19 bgr_7_0.V_TOP.n17 27.8371
R6158 bgr_7_0.V_TOP.n24 bgr_7_0.V_TOP.n23 8.313
R6159 bgr_7_0.V_TOP.n30 bgr_7_0.V_TOP.n29 5.188
R6160 bgr_7_0.V_TOP.n6 bgr_7_0.V_TOP.t31 4.8295
R6161 bgr_7_0.V_TOP.n7 bgr_7_0.V_TOP.t22 4.8295
R6162 bgr_7_0.V_TOP.n8 bgr_7_0.V_TOP.t20 4.8295
R6163 bgr_7_0.V_TOP.n9 bgr_7_0.V_TOP.t45 4.8295
R6164 bgr_7_0.V_TOP.n10 bgr_7_0.V_TOP.t42 4.8295
R6165 bgr_7_0.V_TOP.n11 bgr_7_0.V_TOP.t36 4.8295
R6166 bgr_7_0.V_TOP.n12 bgr_7_0.V_TOP.t17 4.8295
R6167 bgr_7_0.V_TOP.n13 bgr_7_0.V_TOP.t43 4.8295
R6168 bgr_7_0.V_TOP.n14 bgr_7_0.V_TOP.t34 4.8295
R6169 bgr_7_0.V_TOP.n6 bgr_7_0.V_TOP.t35 4.5005
R6170 bgr_7_0.V_TOP.n7 bgr_7_0.V_TOP.t32 4.5005
R6171 bgr_7_0.V_TOP.n8 bgr_7_0.V_TOP.t25 4.5005
R6172 bgr_7_0.V_TOP.n9 bgr_7_0.V_TOP.t21 4.5005
R6173 bgr_7_0.V_TOP.n10 bgr_7_0.V_TOP.t49 4.5005
R6174 bgr_7_0.V_TOP.n11 bgr_7_0.V_TOP.t44 4.5005
R6175 bgr_7_0.V_TOP.n12 bgr_7_0.V_TOP.t23 4.5005
R6176 bgr_7_0.V_TOP.n13 bgr_7_0.V_TOP.t19 4.5005
R6177 bgr_7_0.V_TOP.n16 bgr_7_0.V_TOP.t40 4.5005
R6178 bgr_7_0.V_TOP.n15 bgr_7_0.V_TOP.t47 4.5005
R6179 bgr_7_0.V_TOP.n14 bgr_7_0.V_TOP.t41 4.5005
R6180 bgr_7_0.V_TOP.n25 bgr_7_0.V_TOP.n24 4.5005
R6181 bgr_7_0.V_TOP.n29 bgr_7_0.V_TOP.n27 2.1255
R6182 bgr_7_0.V_TOP.n27 bgr_7_0.V_TOP.n25 2.1255
R6183 bgr_7_0.V_TOP.n25 bgr_7_0.V_TOP.n19 2.1255
R6184 bgr_7_0.V_TOP.n7 bgr_7_0.V_TOP.n6 0.3295
R6185 bgr_7_0.V_TOP.n9 bgr_7_0.V_TOP.n8 0.3295
R6186 bgr_7_0.V_TOP.n11 bgr_7_0.V_TOP.n10 0.3295
R6187 bgr_7_0.V_TOP.n13 bgr_7_0.V_TOP.n12 0.3295
R6188 bgr_7_0.V_TOP.n16 bgr_7_0.V_TOP.n15 0.3295
R6189 bgr_7_0.V_TOP.n15 bgr_7_0.V_TOP.n14 0.3295
R6190 bgr_7_0.V_TOP.n9 bgr_7_0.V_TOP.n7 0.2825
R6191 bgr_7_0.V_TOP.n11 bgr_7_0.V_TOP.n9 0.2825
R6192 bgr_7_0.V_TOP.n13 bgr_7_0.V_TOP.n11 0.2825
R6193 bgr_7_0.V_TOP.n14 bgr_7_0.V_TOP.n13 0.2825
R6194 VOUT-.n8 VOUT-.n0 149.19
R6195 VOUT-.n3 VOUT-.n1 149.19
R6196 VOUT-.n7 VOUT-.n6 148.626
R6197 VOUT-.n5 VOUT-.n4 148.626
R6198 VOUT-.n3 VOUT-.n2 148.626
R6199 VOUT-.n10 VOUT-.n9 144.126
R6200 VOUT-.n91 VOUT-.t18 112.184
R6201 VOUT-.n88 VOUT-.n86 98.9303
R6202 VOUT-.n90 VOUT-.n89 97.8053
R6203 VOUT-.n88 VOUT-.n87 97.8053
R6204 VOUT-.n85 VOUT-.n10 15.0682
R6205 VOUT-.n85 VOUT-.n84 11.5649
R6206 VOUT- VOUT-.n85 9.46925
R6207 VOUT-.n9 VOUT-.t17 6.56717
R6208 VOUT-.n9 VOUT-.t15 6.56717
R6209 VOUT-.n6 VOUT-.t16 6.56717
R6210 VOUT-.n6 VOUT-.t5 6.56717
R6211 VOUT-.n4 VOUT-.t14 6.56717
R6212 VOUT-.n4 VOUT-.t13 6.56717
R6213 VOUT-.n2 VOUT-.t6 6.56717
R6214 VOUT-.n2 VOUT-.t0 6.56717
R6215 VOUT-.n1 VOUT-.t12 6.56717
R6216 VOUT-.n1 VOUT-.t9 6.56717
R6217 VOUT-.n0 VOUT-.t8 6.56717
R6218 VOUT-.n0 VOUT-.t2 6.56717
R6219 VOUT-.n39 VOUT-.t68 4.8295
R6220 VOUT-.n47 VOUT-.t66 4.8295
R6221 VOUT-.n45 VOUT-.t115 4.8295
R6222 VOUT-.n43 VOUT-.t150 4.8295
R6223 VOUT-.n42 VOUT-.t132 4.8295
R6224 VOUT-.n41 VOUT-.t29 4.8295
R6225 VOUT-.n59 VOUT-.t125 4.8295
R6226 VOUT-.n60 VOUT-.t73 4.8295
R6227 VOUT-.n61 VOUT-.t23 4.8295
R6228 VOUT-.n62 VOUT-.t109 4.8295
R6229 VOUT-.n63 VOUT-.t76 4.8295
R6230 VOUT-.n64 VOUT-.t44 4.8295
R6231 VOUT-.n66 VOUT-.t37 4.8295
R6232 VOUT-.n67 VOUT-.t143 4.8295
R6233 VOUT-.n69 VOUT-.t70 4.8295
R6234 VOUT-.n70 VOUT-.t39 4.8295
R6235 VOUT-.n72 VOUT-.t32 4.8295
R6236 VOUT-.n73 VOUT-.t138 4.8295
R6237 VOUT-.n75 VOUT-.t131 4.8295
R6238 VOUT-.n76 VOUT-.t101 4.8295
R6239 VOUT-.n78 VOUT-.t28 4.8295
R6240 VOUT-.n79 VOUT-.t133 4.8295
R6241 VOUT-.n11 VOUT-.t26 4.8295
R6242 VOUT-.n13 VOUT-.t36 4.8295
R6243 VOUT-.n24 VOUT-.t140 4.8295
R6244 VOUT-.n25 VOUT-.t111 4.8295
R6245 VOUT-.n27 VOUT-.t41 4.8295
R6246 VOUT-.n28 VOUT-.t151 4.8295
R6247 VOUT-.n30 VOUT-.t80 4.8295
R6248 VOUT-.n31 VOUT-.t51 4.8295
R6249 VOUT-.n33 VOUT-.t49 4.8295
R6250 VOUT-.n34 VOUT-.t19 4.8295
R6251 VOUT-.n36 VOUT-.t85 4.8295
R6252 VOUT-.n37 VOUT-.t55 4.8295
R6253 VOUT-.n81 VOUT-.t124 4.8295
R6254 VOUT-.n49 VOUT-.t91 4.8154
R6255 VOUT-.n50 VOUT-.t69 4.8154
R6256 VOUT-.n51 VOUT-.t107 4.8154
R6257 VOUT-.n49 VOUT-.t31 4.806
R6258 VOUT-.n50 VOUT-.t149 4.806
R6259 VOUT-.n51 VOUT-.t50 4.806
R6260 VOUT-.n52 VOUT-.t144 4.806
R6261 VOUT-.n52 VOUT-.t83 4.806
R6262 VOUT-.n53 VOUT-.t120 4.806
R6263 VOUT-.n54 VOUT-.t104 4.806
R6264 VOUT-.n55 VOUT-.t137 4.806
R6265 VOUT-.n56 VOUT-.t35 4.806
R6266 VOUT-.n57 VOUT-.t156 4.806
R6267 VOUT-.n14 VOUT-.t71 4.806
R6268 VOUT-.n14 VOUT-.t113 4.806
R6269 VOUT-.n15 VOUT-.t114 4.806
R6270 VOUT-.n15 VOUT-.t24 4.806
R6271 VOUT-.n16 VOUT-.t65 4.806
R6272 VOUT-.n16 VOUT-.t62 4.806
R6273 VOUT-.n17 VOUT-.t154 4.806
R6274 VOUT-.n17 VOUT-.t95 4.806
R6275 VOUT-.n18 VOUT-.t105 4.806
R6276 VOUT-.n18 VOUT-.t126 4.806
R6277 VOUT-.n19 VOUT-.t141 4.806
R6278 VOUT-.n19 VOUT-.t38 4.806
R6279 VOUT-.n20 VOUT-.t92 4.806
R6280 VOUT-.n20 VOUT-.t74 4.806
R6281 VOUT-.n21 VOUT-.t42 4.806
R6282 VOUT-.n22 VOUT-.t82 4.806
R6283 VOUT-.n39 VOUT-.t86 4.5005
R6284 VOUT-.n40 VOUT-.t54 4.5005
R6285 VOUT-.n47 VOUT-.t77 4.5005
R6286 VOUT-.n48 VOUT-.t43 4.5005
R6287 VOUT-.n45 VOUT-.t58 4.5005
R6288 VOUT-.n46 VOUT-.t22 4.5005
R6289 VOUT-.n43 VOUT-.t94 4.5005
R6290 VOUT-.n44 VOUT-.t61 4.5005
R6291 VOUT-.n42 VOUT-.t99 4.5005
R6292 VOUT-.n41 VOUT-.t52 4.5005
R6293 VOUT-.n58 VOUT-.t155 4.5005
R6294 VOUT-.n57 VOUT-.t116 4.5005
R6295 VOUT-.n56 VOUT-.t136 4.5005
R6296 VOUT-.n55 VOUT-.t100 4.5005
R6297 VOUT-.n54 VOUT-.t64 4.5005
R6298 VOUT-.n53 VOUT-.t81 4.5005
R6299 VOUT-.n52 VOUT-.t45 4.5005
R6300 VOUT-.n51 VOUT-.t146 4.5005
R6301 VOUT-.n50 VOUT-.t108 4.5005
R6302 VOUT-.n49 VOUT-.t130 4.5005
R6303 VOUT-.n59 VOUT-.t152 4.5005
R6304 VOUT-.n60 VOUT-.t112 4.5005
R6305 VOUT-.n61 VOUT-.t47 4.5005
R6306 VOUT-.n62 VOUT-.t147 4.5005
R6307 VOUT-.n63 VOUT-.t27 4.5005
R6308 VOUT-.n65 VOUT-.t128 4.5005
R6309 VOUT-.n64 VOUT-.t97 4.5005
R6310 VOUT-.n66 VOUT-.t123 4.5005
R6311 VOUT-.n68 VOUT-.t88 4.5005
R6312 VOUT-.n67 VOUT-.t57 4.5005
R6313 VOUT-.n69 VOUT-.t20 4.5005
R6314 VOUT-.n71 VOUT-.t121 4.5005
R6315 VOUT-.n70 VOUT-.t87 4.5005
R6316 VOUT-.n72 VOUT-.t118 4.5005
R6317 VOUT-.n74 VOUT-.t84 4.5005
R6318 VOUT-.n73 VOUT-.t53 4.5005
R6319 VOUT-.n75 VOUT-.t79 4.5005
R6320 VOUT-.n77 VOUT-.t48 4.5005
R6321 VOUT-.n76 VOUT-.t153 4.5005
R6322 VOUT-.n78 VOUT-.t117 4.5005
R6323 VOUT-.n80 VOUT-.t78 4.5005
R6324 VOUT-.n79 VOUT-.t46 4.5005
R6325 VOUT-.n11 VOUT-.t119 4.5005
R6326 VOUT-.n12 VOUT-.t33 4.5005
R6327 VOUT-.n13 VOUT-.t122 4.5005
R6328 VOUT-.n23 VOUT-.t90 4.5005
R6329 VOUT-.n22 VOUT-.t56 4.5005
R6330 VOUT-.n21 VOUT-.t142 4.5005
R6331 VOUT-.n20 VOUT-.t110 4.5005
R6332 VOUT-.n19 VOUT-.t72 4.5005
R6333 VOUT-.n18 VOUT-.t25 4.5005
R6334 VOUT-.n17 VOUT-.t127 4.5005
R6335 VOUT-.n16 VOUT-.t93 4.5005
R6336 VOUT-.n15 VOUT-.t60 4.5005
R6337 VOUT-.n14 VOUT-.t148 4.5005
R6338 VOUT-.n24 VOUT-.t89 4.5005
R6339 VOUT-.n26 VOUT-.t59 4.5005
R6340 VOUT-.n25 VOUT-.t21 4.5005
R6341 VOUT-.n27 VOUT-.t129 4.5005
R6342 VOUT-.n29 VOUT-.t98 4.5005
R6343 VOUT-.n28 VOUT-.t63 4.5005
R6344 VOUT-.n30 VOUT-.t30 4.5005
R6345 VOUT-.n32 VOUT-.t134 4.5005
R6346 VOUT-.n31 VOUT-.t103 4.5005
R6347 VOUT-.n33 VOUT-.t135 4.5005
R6348 VOUT-.n35 VOUT-.t102 4.5005
R6349 VOUT-.n34 VOUT-.t67 4.5005
R6350 VOUT-.n36 VOUT-.t34 4.5005
R6351 VOUT-.n38 VOUT-.t139 4.5005
R6352 VOUT-.n37 VOUT-.t106 4.5005
R6353 VOUT-.n81 VOUT-.t75 4.5005
R6354 VOUT-.n82 VOUT-.t40 4.5005
R6355 VOUT-.n83 VOUT-.t145 4.5005
R6356 VOUT-.n84 VOUT-.t96 4.5005
R6357 VOUT-.n10 VOUT-.n8 4.5005
R6358 VOUT-.n89 VOUT-.t11 3.42907
R6359 VOUT-.n89 VOUT-.t7 3.42907
R6360 VOUT-.n87 VOUT-.t1 3.42907
R6361 VOUT-.n87 VOUT-.t4 3.42907
R6362 VOUT-.n86 VOUT-.t3 3.42907
R6363 VOUT-.n86 VOUT-.t10 3.42907
R6364 VOUT-.n91 VOUT-.n90 1.30519
R6365 VOUT- VOUT-.n91 1.24269
R6366 VOUT-.n90 VOUT-.n88 1.1255
R6367 VOUT-.n5 VOUT-.n3 0.563
R6368 VOUT-.n7 VOUT-.n5 0.563
R6369 VOUT-.n8 VOUT-.n7 0.563
R6370 VOUT-.n40 VOUT-.n39 0.3295
R6371 VOUT-.n48 VOUT-.n47 0.3295
R6372 VOUT-.n46 VOUT-.n45 0.3295
R6373 VOUT-.n44 VOUT-.n43 0.3295
R6374 VOUT-.n58 VOUT-.n41 0.3295
R6375 VOUT-.n58 VOUT-.n57 0.3295
R6376 VOUT-.n57 VOUT-.n56 0.3295
R6377 VOUT-.n56 VOUT-.n55 0.3295
R6378 VOUT-.n55 VOUT-.n54 0.3295
R6379 VOUT-.n54 VOUT-.n53 0.3295
R6380 VOUT-.n53 VOUT-.n52 0.3295
R6381 VOUT-.n52 VOUT-.n51 0.3295
R6382 VOUT-.n51 VOUT-.n50 0.3295
R6383 VOUT-.n50 VOUT-.n49 0.3295
R6384 VOUT-.n60 VOUT-.n59 0.3295
R6385 VOUT-.n62 VOUT-.n61 0.3295
R6386 VOUT-.n65 VOUT-.n63 0.3295
R6387 VOUT-.n65 VOUT-.n64 0.3295
R6388 VOUT-.n68 VOUT-.n66 0.3295
R6389 VOUT-.n68 VOUT-.n67 0.3295
R6390 VOUT-.n71 VOUT-.n69 0.3295
R6391 VOUT-.n71 VOUT-.n70 0.3295
R6392 VOUT-.n74 VOUT-.n72 0.3295
R6393 VOUT-.n74 VOUT-.n73 0.3295
R6394 VOUT-.n77 VOUT-.n75 0.3295
R6395 VOUT-.n77 VOUT-.n76 0.3295
R6396 VOUT-.n80 VOUT-.n78 0.3295
R6397 VOUT-.n80 VOUT-.n79 0.3295
R6398 VOUT-.n12 VOUT-.n11 0.3295
R6399 VOUT-.n23 VOUT-.n13 0.3295
R6400 VOUT-.n23 VOUT-.n22 0.3295
R6401 VOUT-.n22 VOUT-.n21 0.3295
R6402 VOUT-.n21 VOUT-.n20 0.3295
R6403 VOUT-.n20 VOUT-.n19 0.3295
R6404 VOUT-.n19 VOUT-.n18 0.3295
R6405 VOUT-.n18 VOUT-.n17 0.3295
R6406 VOUT-.n17 VOUT-.n16 0.3295
R6407 VOUT-.n16 VOUT-.n15 0.3295
R6408 VOUT-.n15 VOUT-.n14 0.3295
R6409 VOUT-.n26 VOUT-.n24 0.3295
R6410 VOUT-.n26 VOUT-.n25 0.3295
R6411 VOUT-.n29 VOUT-.n27 0.3295
R6412 VOUT-.n29 VOUT-.n28 0.3295
R6413 VOUT-.n32 VOUT-.n30 0.3295
R6414 VOUT-.n32 VOUT-.n31 0.3295
R6415 VOUT-.n35 VOUT-.n33 0.3295
R6416 VOUT-.n35 VOUT-.n34 0.3295
R6417 VOUT-.n38 VOUT-.n36 0.3295
R6418 VOUT-.n38 VOUT-.n37 0.3295
R6419 VOUT-.n82 VOUT-.n81 0.3295
R6420 VOUT-.n83 VOUT-.n82 0.3295
R6421 VOUT-.n84 VOUT-.n83 0.3295
R6422 VOUT-.n53 VOUT-.n48 0.306
R6423 VOUT-.n54 VOUT-.n46 0.306
R6424 VOUT-.n55 VOUT-.n44 0.306
R6425 VOUT-.n56 VOUT-.n42 0.306
R6426 VOUT-.n58 VOUT-.n40 0.2825
R6427 VOUT-.n60 VOUT-.n58 0.2825
R6428 VOUT-.n62 VOUT-.n60 0.2825
R6429 VOUT-.n65 VOUT-.n62 0.2825
R6430 VOUT-.n68 VOUT-.n65 0.2825
R6431 VOUT-.n71 VOUT-.n68 0.2825
R6432 VOUT-.n74 VOUT-.n71 0.2825
R6433 VOUT-.n77 VOUT-.n74 0.2825
R6434 VOUT-.n80 VOUT-.n77 0.2825
R6435 VOUT-.n23 VOUT-.n12 0.2825
R6436 VOUT-.n26 VOUT-.n23 0.2825
R6437 VOUT-.n29 VOUT-.n26 0.2825
R6438 VOUT-.n32 VOUT-.n29 0.2825
R6439 VOUT-.n35 VOUT-.n32 0.2825
R6440 VOUT-.n38 VOUT-.n35 0.2825
R6441 VOUT-.n82 VOUT-.n38 0.2825
R6442 VOUT-.n82 VOUT-.n80 0.2825
R6443 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 49.197
R6444 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 0.87
R6445 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 0.1603
R6446 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 0.1603
R6447 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 0.1603
R6448 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 0.1603
R6449 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 0.1603
R6450 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 0.1603
R6451 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 0.1603
R6452 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 0.1603
R6453 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 0.1603
R6454 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 0.1603
R6455 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 0.1603
R6456 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 0.1603
R6457 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 0.1603
R6458 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 0.1603
R6459 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 0.1603
R6460 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 0.1603
R6461 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 0.1603
R6462 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 0.1603
R6463 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 0.1603
R6464 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 0.1603
R6465 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 0.1603
R6466 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 0.1603
R6467 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 0.1603
R6468 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 0.1603
R6469 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 0.1603
R6470 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 0.1603
R6471 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 0.1603
R6472 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 0.1603
R6473 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 0.1603
R6474 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 0.1603
R6475 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 0.1603
R6476 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 0.1603
R6477 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 0.1603
R6478 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 0.1603
R6479 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 0.1603
R6480 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 0.1603
R6481 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 0.1603
R6482 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 0.1603
R6483 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 0.1603
R6484 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 0.1603
R6485 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 0.1603
R6486 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 0.1603
R6487 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 0.1603
R6488 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 0.1603
R6489 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 0.1603
R6490 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 0.1603
R6491 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 0.1603
R6492 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 0.1603
R6493 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 0.1603
R6494 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 0.1603
R6495 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 0.1603
R6496 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 0.1603
R6497 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 0.1603
R6498 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 0.1603
R6499 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 0.159278
R6500 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 0.159278
R6501 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 0.159278
R6502 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 0.159278
R6503 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 0.159278
R6504 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 0.159278
R6505 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 0.159278
R6506 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 0.159278
R6507 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 0.159278
R6508 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 0.159278
R6509 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 0.159278
R6510 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 0.159278
R6511 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 0.159278
R6512 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 0.159278
R6513 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 0.159278
R6514 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 0.159278
R6515 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 0.159278
R6516 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 0.159278
R6517 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 0.159278
R6518 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 0.159278
R6519 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 0.159278
R6520 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 0.159278
R6521 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 0.159278
R6522 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 0.159278
R6523 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 0.159278
R6524 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 0.159278
R6525 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 0.159278
R6526 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 0.159278
R6527 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 0.159278
R6528 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 0.159278
R6529 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 0.159278
R6530 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 0.159278
R6531 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 0.159278
R6532 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 0.137822
R6533 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 0.1368
R6534 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 0.1368
R6535 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 0.1368
R6536 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 0.1368
R6537 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 0.1368
R6538 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 0.1368
R6539 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 0.1368
R6540 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 0.1368
R6541 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 0.1368
R6542 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 0.1368
R6543 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 0.1368
R6544 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 0.1368
R6545 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 0.1368
R6546 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 0.1368
R6547 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 0.1368
R6548 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 0.1368
R6549 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 0.1368
R6550 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 0.1368
R6551 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 0.1368
R6552 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 0.1368
R6553 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 0.1368
R6554 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 0.1368
R6555 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 0.1368
R6556 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 0.1368
R6557 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 0.1368
R6558 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 0.1368
R6559 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 0.1368
R6560 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 0.1368
R6561 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 0.1368
R6562 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 0.1368
R6563 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 0.1368
R6564 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 0.1133
R6565 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 0.1133
R6566 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 0.1133
R6567 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 0.1133
R6568 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 0.1133
R6569 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 0.1133
R6570 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 0.1133
R6571 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 0.1133
R6572 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 0.1133
R6573 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 0.1133
R6574 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 0.1133
R6575 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 0.1133
R6576 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 0.1133
R6577 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 0.1133
R6578 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 0.1133
R6579 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 0.1133
R6580 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 0.1133
R6581 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 0.1133
R6582 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 0.00152174
R6583 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 0.00152174
R6584 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 0.00152174
R6585 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 0.00152174
R6586 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 0.00152174
R6587 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 0.00152174
R6588 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 0.00152174
R6589 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 0.00152174
R6590 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 0.00152174
R6591 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 0.00152174
R6592 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 0.00152174
R6593 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 0.00152174
R6594 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 0.00152174
R6595 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 0.00152174
R6596 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 0.00152174
R6597 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 0.00152174
R6598 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 0.00152174
R6599 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 0.00152174
R6600 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 0.00152174
R6601 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 0.00152174
R6602 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 0.00152174
R6603 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 0.00152174
R6604 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 0.00152174
R6605 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 0.00152174
R6606 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 0.00152174
R6607 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 0.00152174
R6608 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 0.00152174
R6609 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 0.00152174
R6610 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 0.00152174
R6611 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 0.00152174
R6612 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 0.00152174
R6613 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 0.00152174
R6614 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 0.00152174
R6615 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 0.00152174
R6616 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 0.00152174
R6617 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t5 554.301
R6618 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t3 442.837
R6619 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 193.869
R6620 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 173.088
R6621 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 86.8857
R6622 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t0 15.7605
R6623 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t1 15.7605
R6624 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t4 9.6005
R6625 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 9.6005
R6626 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 610.534
R6627 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 610.534
R6628 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 488.428
R6629 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 488.428
R6630 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 433.8
R6631 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 433.8
R6632 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 433.8
R6633 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 433.8
R6634 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 433.8
R6635 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 433.8
R6636 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 433.8
R6637 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 433.8
R6638 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 433.8
R6639 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 433.8
R6640 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 433.8
R6641 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 433.8
R6642 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 433.8
R6643 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 433.8
R6644 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 433.8
R6645 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 433.8
R6646 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 277.755
R6647 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 176.733
R6648 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 176.733
R6649 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 176.733
R6650 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 176.733
R6651 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 176.733
R6652 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 176.733
R6653 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 176.733
R6654 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 176.733
R6655 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 176.733
R6656 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 176.733
R6657 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 176.733
R6658 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 176.733
R6659 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 176.733
R6660 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 176.733
R6661 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 175.587
R6662 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 161.3
R6663 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 133.786
R6664 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 121.218
R6665 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 111.778
R6666 bgr_7_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 71.358
R6667 bgr_7_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 63.7817
R6668 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 54.6272
R6669 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 54.6272
R6670 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 19.7005
R6671 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 19.7005
R6672 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 19.7005
R6673 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 19.7005
R6674 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t4 16.0005
R6675 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t3 16.0005
R6676 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t7 16.0005
R6677 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t5 16.0005
R6678 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 0.583833
R6679 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 0.53175
R6680 two_stage_opamp_dummy_magic_14_0.V_source.n26 two_stage_opamp_dummy_magic_14_0.V_source.t34 171.525
R6681 two_stage_opamp_dummy_magic_14_0.V_source.n10 two_stage_opamp_dummy_magic_14_0.V_source.n8 114.469
R6682 two_stage_opamp_dummy_magic_14_0.V_source.n3 two_stage_opamp_dummy_magic_14_0.V_source.n1 114.469
R6683 two_stage_opamp_dummy_magic_14_0.V_source.n18 two_stage_opamp_dummy_magic_14_0.V_source.n17 113.906
R6684 two_stage_opamp_dummy_magic_14_0.V_source.n16 two_stage_opamp_dummy_magic_14_0.V_source.n15 113.906
R6685 two_stage_opamp_dummy_magic_14_0.V_source.n14 two_stage_opamp_dummy_magic_14_0.V_source.n13 113.906
R6686 two_stage_opamp_dummy_magic_14_0.V_source.n12 two_stage_opamp_dummy_magic_14_0.V_source.n11 113.906
R6687 two_stage_opamp_dummy_magic_14_0.V_source.n10 two_stage_opamp_dummy_magic_14_0.V_source.n9 113.906
R6688 two_stage_opamp_dummy_magic_14_0.V_source.n7 two_stage_opamp_dummy_magic_14_0.V_source.n6 113.906
R6689 two_stage_opamp_dummy_magic_14_0.V_source.n5 two_stage_opamp_dummy_magic_14_0.V_source.n4 113.906
R6690 two_stage_opamp_dummy_magic_14_0.V_source.n3 two_stage_opamp_dummy_magic_14_0.V_source.n2 113.906
R6691 two_stage_opamp_dummy_magic_14_0.V_source.n22 two_stage_opamp_dummy_magic_14_0.V_source.n0 102.941
R6692 two_stage_opamp_dummy_magic_14_0.V_source.n38 two_stage_opamp_dummy_magic_14_0.V_source.n37 102.285
R6693 two_stage_opamp_dummy_magic_14_0.V_source.n36 two_stage_opamp_dummy_magic_14_0.V_source.n35 102.284
R6694 two_stage_opamp_dummy_magic_14_0.V_source.n34 two_stage_opamp_dummy_magic_14_0.V_source.n33 102.284
R6695 two_stage_opamp_dummy_magic_14_0.V_source.n32 two_stage_opamp_dummy_magic_14_0.V_source.n31 102.284
R6696 two_stage_opamp_dummy_magic_14_0.V_source.n30 two_stage_opamp_dummy_magic_14_0.V_source.n29 102.284
R6697 two_stage_opamp_dummy_magic_14_0.V_source.n28 two_stage_opamp_dummy_magic_14_0.V_source.n27 102.284
R6698 two_stage_opamp_dummy_magic_14_0.V_source.n26 two_stage_opamp_dummy_magic_14_0.V_source.n25 102.284
R6699 two_stage_opamp_dummy_magic_14_0.V_source.n24 two_stage_opamp_dummy_magic_14_0.V_source.n23 102.284
R6700 two_stage_opamp_dummy_magic_14_0.V_source.n21 two_stage_opamp_dummy_magic_14_0.V_source.n20 97.7845
R6701 two_stage_opamp_dummy_magic_14_0.V_source.n17 two_stage_opamp_dummy_magic_14_0.V_source.t1 16.0005
R6702 two_stage_opamp_dummy_magic_14_0.V_source.n17 two_stage_opamp_dummy_magic_14_0.V_source.t6 16.0005
R6703 two_stage_opamp_dummy_magic_14_0.V_source.n15 two_stage_opamp_dummy_magic_14_0.V_source.t7 16.0005
R6704 two_stage_opamp_dummy_magic_14_0.V_source.n15 two_stage_opamp_dummy_magic_14_0.V_source.t40 16.0005
R6705 two_stage_opamp_dummy_magic_14_0.V_source.n13 two_stage_opamp_dummy_magic_14_0.V_source.t36 16.0005
R6706 two_stage_opamp_dummy_magic_14_0.V_source.n13 two_stage_opamp_dummy_magic_14_0.V_source.t35 16.0005
R6707 two_stage_opamp_dummy_magic_14_0.V_source.n11 two_stage_opamp_dummy_magic_14_0.V_source.t4 16.0005
R6708 two_stage_opamp_dummy_magic_14_0.V_source.n11 two_stage_opamp_dummy_magic_14_0.V_source.t38 16.0005
R6709 two_stage_opamp_dummy_magic_14_0.V_source.n9 two_stage_opamp_dummy_magic_14_0.V_source.t5 16.0005
R6710 two_stage_opamp_dummy_magic_14_0.V_source.n9 two_stage_opamp_dummy_magic_14_0.V_source.t3 16.0005
R6711 two_stage_opamp_dummy_magic_14_0.V_source.n8 two_stage_opamp_dummy_magic_14_0.V_source.t32 16.0005
R6712 two_stage_opamp_dummy_magic_14_0.V_source.n8 two_stage_opamp_dummy_magic_14_0.V_source.t10 16.0005
R6713 two_stage_opamp_dummy_magic_14_0.V_source.n6 two_stage_opamp_dummy_magic_14_0.V_source.t30 16.0005
R6714 two_stage_opamp_dummy_magic_14_0.V_source.n6 two_stage_opamp_dummy_magic_14_0.V_source.t8 16.0005
R6715 two_stage_opamp_dummy_magic_14_0.V_source.n4 two_stage_opamp_dummy_magic_14_0.V_source.t39 16.0005
R6716 two_stage_opamp_dummy_magic_14_0.V_source.n4 two_stage_opamp_dummy_magic_14_0.V_source.t2 16.0005
R6717 two_stage_opamp_dummy_magic_14_0.V_source.n2 two_stage_opamp_dummy_magic_14_0.V_source.t9 16.0005
R6718 two_stage_opamp_dummy_magic_14_0.V_source.n2 two_stage_opamp_dummy_magic_14_0.V_source.t31 16.0005
R6719 two_stage_opamp_dummy_magic_14_0.V_source.n1 two_stage_opamp_dummy_magic_14_0.V_source.t37 16.0005
R6720 two_stage_opamp_dummy_magic_14_0.V_source.n1 two_stage_opamp_dummy_magic_14_0.V_source.t0 16.0005
R6721 two_stage_opamp_dummy_magic_14_0.V_source.n35 two_stage_opamp_dummy_magic_14_0.V_source.t27 9.6005
R6722 two_stage_opamp_dummy_magic_14_0.V_source.n35 two_stage_opamp_dummy_magic_14_0.V_source.t17 9.6005
R6723 two_stage_opamp_dummy_magic_14_0.V_source.n33 two_stage_opamp_dummy_magic_14_0.V_source.t23 9.6005
R6724 two_stage_opamp_dummy_magic_14_0.V_source.n33 two_stage_opamp_dummy_magic_14_0.V_source.t15 9.6005
R6725 two_stage_opamp_dummy_magic_14_0.V_source.n31 two_stage_opamp_dummy_magic_14_0.V_source.t26 9.6005
R6726 two_stage_opamp_dummy_magic_14_0.V_source.n31 two_stage_opamp_dummy_magic_14_0.V_source.t16 9.6005
R6727 two_stage_opamp_dummy_magic_14_0.V_source.n29 two_stage_opamp_dummy_magic_14_0.V_source.t22 9.6005
R6728 two_stage_opamp_dummy_magic_14_0.V_source.n29 two_stage_opamp_dummy_magic_14_0.V_source.t12 9.6005
R6729 two_stage_opamp_dummy_magic_14_0.V_source.n27 two_stage_opamp_dummy_magic_14_0.V_source.t20 9.6005
R6730 two_stage_opamp_dummy_magic_14_0.V_source.n27 two_stage_opamp_dummy_magic_14_0.V_source.t28 9.6005
R6731 two_stage_opamp_dummy_magic_14_0.V_source.n25 two_stage_opamp_dummy_magic_14_0.V_source.t18 9.6005
R6732 two_stage_opamp_dummy_magic_14_0.V_source.n25 two_stage_opamp_dummy_magic_14_0.V_source.t24 9.6005
R6733 two_stage_opamp_dummy_magic_14_0.V_source.n23 two_stage_opamp_dummy_magic_14_0.V_source.t14 9.6005
R6734 two_stage_opamp_dummy_magic_14_0.V_source.n23 two_stage_opamp_dummy_magic_14_0.V_source.t21 9.6005
R6735 two_stage_opamp_dummy_magic_14_0.V_source.n20 two_stage_opamp_dummy_magic_14_0.V_source.t13 9.6005
R6736 two_stage_opamp_dummy_magic_14_0.V_source.n20 two_stage_opamp_dummy_magic_14_0.V_source.t25 9.6005
R6737 two_stage_opamp_dummy_magic_14_0.V_source.n0 two_stage_opamp_dummy_magic_14_0.V_source.t33 9.6005
R6738 two_stage_opamp_dummy_magic_14_0.V_source.n0 two_stage_opamp_dummy_magic_14_0.V_source.t11 9.6005
R6739 two_stage_opamp_dummy_magic_14_0.V_source.t29 two_stage_opamp_dummy_magic_14_0.V_source.n38 9.6005
R6740 two_stage_opamp_dummy_magic_14_0.V_source.n38 two_stage_opamp_dummy_magic_14_0.V_source.t19 9.6005
R6741 two_stage_opamp_dummy_magic_14_0.V_source.n21 two_stage_opamp_dummy_magic_14_0.V_source.n19 9.17758
R6742 two_stage_opamp_dummy_magic_14_0.V_source.n18 two_stage_opamp_dummy_magic_14_0.V_source.n16 4.6255
R6743 two_stage_opamp_dummy_magic_14_0.V_source.n22 two_stage_opamp_dummy_magic_14_0.V_source.n21 4.5005
R6744 two_stage_opamp_dummy_magic_14_0.V_source.n28 two_stage_opamp_dummy_magic_14_0.V_source.n26 0.563
R6745 two_stage_opamp_dummy_magic_14_0.V_source.n30 two_stage_opamp_dummy_magic_14_0.V_source.n28 0.563
R6746 two_stage_opamp_dummy_magic_14_0.V_source.n32 two_stage_opamp_dummy_magic_14_0.V_source.n30 0.563
R6747 two_stage_opamp_dummy_magic_14_0.V_source.n34 two_stage_opamp_dummy_magic_14_0.V_source.n32 0.563
R6748 two_stage_opamp_dummy_magic_14_0.V_source.n36 two_stage_opamp_dummy_magic_14_0.V_source.n34 0.563
R6749 two_stage_opamp_dummy_magic_14_0.V_source.n37 two_stage_opamp_dummy_magic_14_0.V_source.n36 0.563
R6750 two_stage_opamp_dummy_magic_14_0.V_source.n12 two_stage_opamp_dummy_magic_14_0.V_source.n10 0.563
R6751 two_stage_opamp_dummy_magic_14_0.V_source.n14 two_stage_opamp_dummy_magic_14_0.V_source.n12 0.563
R6752 two_stage_opamp_dummy_magic_14_0.V_source.n16 two_stage_opamp_dummy_magic_14_0.V_source.n14 0.563
R6753 two_stage_opamp_dummy_magic_14_0.V_source.n5 two_stage_opamp_dummy_magic_14_0.V_source.n3 0.563
R6754 two_stage_opamp_dummy_magic_14_0.V_source.n7 two_stage_opamp_dummy_magic_14_0.V_source.n5 0.563
R6755 two_stage_opamp_dummy_magic_14_0.V_source.n24 two_stage_opamp_dummy_magic_14_0.V_source.n22 0.563
R6756 two_stage_opamp_dummy_magic_14_0.V_source.n37 two_stage_opamp_dummy_magic_14_0.V_source.n24 0.563
R6757 two_stage_opamp_dummy_magic_14_0.V_source.n19 two_stage_opamp_dummy_magic_14_0.V_source.n18 0.234875
R6758 two_stage_opamp_dummy_magic_14_0.V_source.n19 two_stage_opamp_dummy_magic_14_0.V_source.n7 0.234875
R6759 VOUT+.n8 VOUT+.n6 149.19
R6760 VOUT+.n14 VOUT+.n13 149.19
R6761 VOUT+.n12 VOUT+.n11 148.626
R6762 VOUT+.n10 VOUT+.n9 148.626
R6763 VOUT+.n8 VOUT+.n7 148.626
R6764 VOUT+.n16 VOUT+.n15 144.126
R6765 VOUT+.n5 VOUT+.t10 112.184
R6766 VOUT+.n2 VOUT+.n0 98.9303
R6767 VOUT+.n4 VOUT+.n3 97.8053
R6768 VOUT+.n2 VOUT+.n1 97.8053
R6769 VOUT+.n91 VOUT+.n16 15.0682
R6770 VOUT+.n91 VOUT+.n90 11.5649
R6771 VOUT+ VOUT+.n91 9.2505
R6772 VOUT+.n15 VOUT+.t1 6.56717
R6773 VOUT+.n15 VOUT+.t18 6.56717
R6774 VOUT+.n13 VOUT+.t6 6.56717
R6775 VOUT+.n13 VOUT+.t13 6.56717
R6776 VOUT+.n11 VOUT+.t5 6.56717
R6777 VOUT+.n11 VOUT+.t9 6.56717
R6778 VOUT+.n9 VOUT+.t17 6.56717
R6779 VOUT+.n9 VOUT+.t3 6.56717
R6780 VOUT+.n7 VOUT+.t4 6.56717
R6781 VOUT+.n7 VOUT+.t7 6.56717
R6782 VOUT+.n6 VOUT+.t12 6.56717
R6783 VOUT+.n6 VOUT+.t0 6.56717
R6784 VOUT+.n45 VOUT+.t56 4.8295
R6785 VOUT+.n47 VOUT+.t105 4.8295
R6786 VOUT+.n48 VOUT+.t29 4.8295
R6787 VOUT+.n50 VOUT+.t60 4.8295
R6788 VOUT+.n52 VOUT+.t115 4.8295
R6789 VOUT+.n63 VOUT+.t20 4.8295
R6790 VOUT+.n66 VOUT+.t31 4.8295
R6791 VOUT+.n65 VOUT+.t121 4.8295
R6792 VOUT+.n68 VOUT+.t67 4.8295
R6793 VOUT+.n67 VOUT+.t152 4.8295
R6794 VOUT+.n69 VOUT+.t131 4.8295
R6795 VOUT+.n70 VOUT+.t118 4.8295
R6796 VOUT+.n72 VOUT+.t89 4.8295
R6797 VOUT+.n73 VOUT+.t76 4.8295
R6798 VOUT+.n75 VOUT+.t127 4.8295
R6799 VOUT+.n76 VOUT+.t110 4.8295
R6800 VOUT+.n78 VOUT+.t84 4.8295
R6801 VOUT+.n79 VOUT+.t68 4.8295
R6802 VOUT+.n81 VOUT+.t42 4.8295
R6803 VOUT+.n82 VOUT+.t30 4.8295
R6804 VOUT+.n84 VOUT+.t81 4.8295
R6805 VOUT+.n85 VOUT+.t64 4.8295
R6806 VOUT+.n17 VOUT+.t150 4.8295
R6807 VOUT+.n28 VOUT+.t75 4.8295
R6808 VOUT+.n30 VOUT+.t54 4.8295
R6809 VOUT+.n31 VOUT+.t34 4.8295
R6810 VOUT+.n33 VOUT+.t95 4.8295
R6811 VOUT+.n34 VOUT+.t79 4.8295
R6812 VOUT+.n36 VOUT+.t134 4.8295
R6813 VOUT+.n37 VOUT+.t122 4.8295
R6814 VOUT+.n39 VOUT+.t102 4.8295
R6815 VOUT+.n40 VOUT+.t82 4.8295
R6816 VOUT+.n42 VOUT+.t137 4.8295
R6817 VOUT+.n43 VOUT+.t126 4.8295
R6818 VOUT+.n87 VOUT+.t28 4.8295
R6819 VOUT+.n56 VOUT+.t57 4.8154
R6820 VOUT+.n55 VOUT+.t33 4.8154
R6821 VOUT+.n54 VOUT+.t77 4.8154
R6822 VOUT+.n62 VOUT+.t116 4.806
R6823 VOUT+.n61 VOUT+.t147 4.806
R6824 VOUT+.n60 VOUT+.t43 4.806
R6825 VOUT+.n59 VOUT+.t83 4.806
R6826 VOUT+.n58 VOUT+.t63 4.806
R6827 VOUT+.n57 VOUT+.t26 4.806
R6828 VOUT+.n57 VOUT+.t103 4.806
R6829 VOUT+.n56 VOUT+.t135 4.806
R6830 VOUT+.n55 VOUT+.t120 4.806
R6831 VOUT+.n54 VOUT+.t155 4.806
R6832 VOUT+.n27 VOUT+.t91 4.806
R6833 VOUT+.n26 VOUT+.t38 4.806
R6834 VOUT+.n25 VOUT+.t130 4.806
R6835 VOUT+.n25 VOUT+.t90 4.806
R6836 VOUT+.n24 VOUT+.t80 4.806
R6837 VOUT+.n24 VOUT+.t128 4.806
R6838 VOUT+.n23 VOUT+.t124 4.806
R6839 VOUT+.n23 VOUT+.t32 4.806
R6840 VOUT+.n22 VOUT+.t70 4.806
R6841 VOUT+.n22 VOUT+.t73 4.806
R6842 VOUT+.n21 VOUT+.t23 4.806
R6843 VOUT+.n21 VOUT+.t108 4.806
R6844 VOUT+.n20 VOUT+.t62 4.806
R6845 VOUT+.n20 VOUT+.t19 4.806
R6846 VOUT+.n19 VOUT+.t151 4.806
R6847 VOUT+.n19 VOUT+.t49 4.806
R6848 VOUT+.n46 VOUT+.t132 4.5005
R6849 VOUT+.n45 VOUT+.t96 4.5005
R6850 VOUT+.n47 VOUT+.t69 4.5005
R6851 VOUT+.n48 VOUT+.t139 4.5005
R6852 VOUT+.n49 VOUT+.t109 4.5005
R6853 VOUT+.n50 VOUT+.t37 4.5005
R6854 VOUT+.n51 VOUT+.t144 4.5005
R6855 VOUT+.n52 VOUT+.t21 4.5005
R6856 VOUT+.n53 VOUT+.t125 4.5005
R6857 VOUT+.n54 VOUT+.t119 4.5005
R6858 VOUT+.n55 VOUT+.t78 4.5005
R6859 VOUT+.n56 VOUT+.t97 4.5005
R6860 VOUT+.n57 VOUT+.t61 4.5005
R6861 VOUT+.n58 VOUT+.t27 4.5005
R6862 VOUT+.n59 VOUT+.t41 4.5005
R6863 VOUT+.n60 VOUT+.t145 4.5005
R6864 VOUT+.n61 VOUT+.t113 4.5005
R6865 VOUT+.n62 VOUT+.t72 4.5005
R6866 VOUT+.n64 VOUT+.t92 4.5005
R6867 VOUT+.n63 VOUT+.t55 4.5005
R6868 VOUT+.n66 VOUT+.t50 4.5005
R6869 VOUT+.n65 VOUT+.t156 4.5005
R6870 VOUT+.n68 VOUT+.t86 4.5005
R6871 VOUT+.n67 VOUT+.t47 4.5005
R6872 VOUT+.n69 VOUT+.t94 4.5005
R6873 VOUT+.n71 VOUT+.t39 4.5005
R6874 VOUT+.n70 VOUT+.t146 4.5005
R6875 VOUT+.n72 VOUT+.t53 4.5005
R6876 VOUT+.n74 VOUT+.t142 4.5005
R6877 VOUT+.n73 VOUT+.t112 4.5005
R6878 VOUT+.n75 VOUT+.t88 4.5005
R6879 VOUT+.n77 VOUT+.t35 4.5005
R6880 VOUT+.n76 VOUT+.t140 4.5005
R6881 VOUT+.n78 VOUT+.t46 4.5005
R6882 VOUT+.n80 VOUT+.t136 4.5005
R6883 VOUT+.n79 VOUT+.t104 4.5005
R6884 VOUT+.n81 VOUT+.t149 4.5005
R6885 VOUT+.n83 VOUT+.t99 4.5005
R6886 VOUT+.n82 VOUT+.t65 4.5005
R6887 VOUT+.n84 VOUT+.t40 4.5005
R6888 VOUT+.n86 VOUT+.t133 4.5005
R6889 VOUT+.n85 VOUT+.t98 4.5005
R6890 VOUT+.n18 VOUT+.t45 4.5005
R6891 VOUT+.n17 VOUT+.t101 4.5005
R6892 VOUT+.n19 VOUT+.t85 4.5005
R6893 VOUT+.n20 VOUT+.t48 4.5005
R6894 VOUT+.n21 VOUT+.t138 4.5005
R6895 VOUT+.n22 VOUT+.t107 4.5005
R6896 VOUT+.n23 VOUT+.t71 4.5005
R6897 VOUT+.n24 VOUT+.t25 4.5005
R6898 VOUT+.n25 VOUT+.t129 4.5005
R6899 VOUT+.n26 VOUT+.t87 4.5005
R6900 VOUT+.n27 VOUT+.t52 4.5005
R6901 VOUT+.n29 VOUT+.t141 4.5005
R6902 VOUT+.n28 VOUT+.t111 4.5005
R6903 VOUT+.n30 VOUT+.t24 4.5005
R6904 VOUT+.n32 VOUT+.t114 4.5005
R6905 VOUT+.n31 VOUT+.t74 4.5005
R6906 VOUT+.n33 VOUT+.t59 4.5005
R6907 VOUT+.n35 VOUT+.t148 4.5005
R6908 VOUT+.n34 VOUT+.t117 4.5005
R6909 VOUT+.n36 VOUT+.t100 4.5005
R6910 VOUT+.n38 VOUT+.t44 4.5005
R6911 VOUT+.n37 VOUT+.t153 4.5005
R6912 VOUT+.n39 VOUT+.t66 4.5005
R6913 VOUT+.n41 VOUT+.t154 4.5005
R6914 VOUT+.n40 VOUT+.t123 4.5005
R6915 VOUT+.n42 VOUT+.t106 4.5005
R6916 VOUT+.n44 VOUT+.t51 4.5005
R6917 VOUT+.n43 VOUT+.t22 4.5005
R6918 VOUT+.n90 VOUT+.t36 4.5005
R6919 VOUT+.n89 VOUT+.t143 4.5005
R6920 VOUT+.n88 VOUT+.t93 4.5005
R6921 VOUT+.n87 VOUT+.t58 4.5005
R6922 VOUT+.n16 VOUT+.n14 4.5005
R6923 VOUT+.n3 VOUT+.t8 3.42907
R6924 VOUT+.n3 VOUT+.t15 3.42907
R6925 VOUT+.n1 VOUT+.t14 3.42907
R6926 VOUT+.n1 VOUT+.t11 3.42907
R6927 VOUT+.n0 VOUT+.t16 3.42907
R6928 VOUT+.n0 VOUT+.t2 3.42907
R6929 VOUT+ VOUT+.n5 1.46144
R6930 VOUT+.n5 VOUT+.n4 1.30519
R6931 VOUT+.n4 VOUT+.n2 1.1255
R6932 VOUT+.n10 VOUT+.n8 0.563
R6933 VOUT+.n12 VOUT+.n10 0.563
R6934 VOUT+.n14 VOUT+.n12 0.563
R6935 VOUT+.n46 VOUT+.n45 0.3295
R6936 VOUT+.n49 VOUT+.n48 0.3295
R6937 VOUT+.n51 VOUT+.n50 0.3295
R6938 VOUT+.n53 VOUT+.n52 0.3295
R6939 VOUT+.n55 VOUT+.n54 0.3295
R6940 VOUT+.n56 VOUT+.n55 0.3295
R6941 VOUT+.n57 VOUT+.n56 0.3295
R6942 VOUT+.n58 VOUT+.n57 0.3295
R6943 VOUT+.n59 VOUT+.n58 0.3295
R6944 VOUT+.n60 VOUT+.n59 0.3295
R6945 VOUT+.n61 VOUT+.n60 0.3295
R6946 VOUT+.n62 VOUT+.n61 0.3295
R6947 VOUT+.n64 VOUT+.n62 0.3295
R6948 VOUT+.n64 VOUT+.n63 0.3295
R6949 VOUT+.n66 VOUT+.n65 0.3295
R6950 VOUT+.n68 VOUT+.n67 0.3295
R6951 VOUT+.n71 VOUT+.n69 0.3295
R6952 VOUT+.n71 VOUT+.n70 0.3295
R6953 VOUT+.n74 VOUT+.n72 0.3295
R6954 VOUT+.n74 VOUT+.n73 0.3295
R6955 VOUT+.n77 VOUT+.n75 0.3295
R6956 VOUT+.n77 VOUT+.n76 0.3295
R6957 VOUT+.n80 VOUT+.n78 0.3295
R6958 VOUT+.n80 VOUT+.n79 0.3295
R6959 VOUT+.n83 VOUT+.n81 0.3295
R6960 VOUT+.n83 VOUT+.n82 0.3295
R6961 VOUT+.n86 VOUT+.n84 0.3295
R6962 VOUT+.n86 VOUT+.n85 0.3295
R6963 VOUT+.n18 VOUT+.n17 0.3295
R6964 VOUT+.n20 VOUT+.n19 0.3295
R6965 VOUT+.n21 VOUT+.n20 0.3295
R6966 VOUT+.n22 VOUT+.n21 0.3295
R6967 VOUT+.n23 VOUT+.n22 0.3295
R6968 VOUT+.n24 VOUT+.n23 0.3295
R6969 VOUT+.n25 VOUT+.n24 0.3295
R6970 VOUT+.n26 VOUT+.n25 0.3295
R6971 VOUT+.n27 VOUT+.n26 0.3295
R6972 VOUT+.n29 VOUT+.n27 0.3295
R6973 VOUT+.n29 VOUT+.n28 0.3295
R6974 VOUT+.n32 VOUT+.n30 0.3295
R6975 VOUT+.n32 VOUT+.n31 0.3295
R6976 VOUT+.n35 VOUT+.n33 0.3295
R6977 VOUT+.n35 VOUT+.n34 0.3295
R6978 VOUT+.n38 VOUT+.n36 0.3295
R6979 VOUT+.n38 VOUT+.n37 0.3295
R6980 VOUT+.n41 VOUT+.n39 0.3295
R6981 VOUT+.n41 VOUT+.n40 0.3295
R6982 VOUT+.n44 VOUT+.n42 0.3295
R6983 VOUT+.n44 VOUT+.n43 0.3295
R6984 VOUT+.n90 VOUT+.n89 0.3295
R6985 VOUT+.n89 VOUT+.n88 0.3295
R6986 VOUT+.n88 VOUT+.n87 0.3295
R6987 VOUT+.n61 VOUT+.n47 0.306
R6988 VOUT+.n60 VOUT+.n49 0.306
R6989 VOUT+.n59 VOUT+.n51 0.306
R6990 VOUT+.n58 VOUT+.n53 0.306
R6991 VOUT+.n64 VOUT+.n46 0.2825
R6992 VOUT+.n66 VOUT+.n64 0.2825
R6993 VOUT+.n68 VOUT+.n66 0.2825
R6994 VOUT+.n71 VOUT+.n68 0.2825
R6995 VOUT+.n74 VOUT+.n71 0.2825
R6996 VOUT+.n77 VOUT+.n74 0.2825
R6997 VOUT+.n80 VOUT+.n77 0.2825
R6998 VOUT+.n83 VOUT+.n80 0.2825
R6999 VOUT+.n86 VOUT+.n83 0.2825
R7000 VOUT+.n29 VOUT+.n18 0.2825
R7001 VOUT+.n32 VOUT+.n29 0.2825
R7002 VOUT+.n35 VOUT+.n32 0.2825
R7003 VOUT+.n38 VOUT+.n35 0.2825
R7004 VOUT+.n41 VOUT+.n38 0.2825
R7005 VOUT+.n44 VOUT+.n41 0.2825
R7006 VOUT+.n88 VOUT+.n44 0.2825
R7007 VOUT+.n88 VOUT+.n86 0.2825
R7008 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 50.3211
R7009 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 0.1603
R7010 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 0.1603
R7011 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 0.1603
R7012 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 0.1603
R7013 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 0.1603
R7014 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 0.1603
R7015 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 0.1603
R7016 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 0.1603
R7017 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 0.1603
R7018 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 0.1603
R7019 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 0.1603
R7020 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 0.1603
R7021 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 0.1603
R7022 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 0.1603
R7023 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 0.1603
R7024 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 0.1603
R7025 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 0.1603
R7026 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 0.1603
R7027 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 0.1603
R7028 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 0.1603
R7029 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 0.1603
R7030 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 0.1603
R7031 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 0.1603
R7032 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 0.1603
R7033 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 0.1603
R7034 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 0.1603
R7035 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 0.1603
R7036 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 0.1603
R7037 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 0.1603
R7038 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 0.1603
R7039 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 0.1603
R7040 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 0.1603
R7041 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 0.1603
R7042 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 0.1603
R7043 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 0.1603
R7044 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 0.1603
R7045 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 0.1603
R7046 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 0.1603
R7047 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 0.1603
R7048 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 0.1603
R7049 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 0.1603
R7050 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 0.1603
R7051 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 0.1603
R7052 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 0.1603
R7053 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 0.1603
R7054 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 0.1603
R7055 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 0.1603
R7056 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 0.1603
R7057 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 0.1603
R7058 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 0.1603
R7059 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 0.1603
R7060 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 0.1603
R7061 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 0.1603
R7062 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 0.1603
R7063 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 0.159278
R7064 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 0.159278
R7065 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 0.159278
R7066 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 0.159278
R7067 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 0.159278
R7068 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 0.159278
R7069 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 0.159278
R7070 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 0.159278
R7071 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 0.159278
R7072 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 0.159278
R7073 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 0.159278
R7074 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 0.159278
R7075 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 0.159278
R7076 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 0.159278
R7077 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 0.159278
R7078 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 0.159278
R7079 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 0.159278
R7080 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 0.159278
R7081 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 0.159278
R7082 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 0.159278
R7083 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 0.159278
R7084 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 0.159278
R7085 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 0.159278
R7086 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 0.159278
R7087 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 0.159278
R7088 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 0.159278
R7089 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 0.159278
R7090 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 0.159278
R7091 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 0.159278
R7092 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 0.159278
R7093 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 0.159278
R7094 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 0.159278
R7095 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 0.159278
R7096 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 0.137822
R7097 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 0.1368
R7098 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 0.1368
R7099 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 0.1368
R7100 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 0.1368
R7101 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 0.1368
R7102 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 0.1368
R7103 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 0.1368
R7104 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 0.1368
R7105 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 0.1368
R7106 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 0.1368
R7107 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 0.1368
R7108 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 0.1368
R7109 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 0.1368
R7110 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 0.1368
R7111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 0.1368
R7112 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 0.1368
R7113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 0.1368
R7114 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 0.1368
R7115 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 0.1368
R7116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 0.1368
R7117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 0.1368
R7118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 0.1368
R7119 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 0.1368
R7120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 0.1368
R7121 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 0.1368
R7122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 0.1368
R7123 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 0.1368
R7124 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 0.1368
R7125 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 0.1368
R7126 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 0.1368
R7127 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 0.1368
R7128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 0.1133
R7129 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 0.1133
R7130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 0.1133
R7131 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 0.1133
R7132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 0.1133
R7133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 0.1133
R7134 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 0.1133
R7135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 0.1133
R7136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 0.1133
R7137 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 0.1133
R7138 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 0.1133
R7139 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 0.1133
R7140 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 0.1133
R7141 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 0.1133
R7142 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 0.1133
R7143 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 0.1133
R7144 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 0.1133
R7145 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 0.1133
R7146 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 0.00152174
R7147 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 0.00152174
R7148 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 0.00152174
R7149 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 0.00152174
R7150 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 0.00152174
R7151 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 0.00152174
R7152 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 0.00152174
R7153 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 0.00152174
R7154 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 0.00152174
R7155 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 0.00152174
R7156 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 0.00152174
R7157 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 0.00152174
R7158 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 0.00152174
R7159 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 0.00152174
R7160 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 0.00152174
R7161 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 0.00152174
R7162 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 0.00152174
R7163 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 0.00152174
R7164 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 0.00152174
R7165 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 0.00152174
R7166 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 0.00152174
R7167 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 0.00152174
R7168 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 0.00152174
R7169 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 0.00152174
R7170 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 0.00152174
R7171 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 0.00152174
R7172 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 0.00152174
R7173 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 0.00152174
R7174 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 0.00152174
R7175 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 0.00152174
R7176 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 0.00152174
R7177 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 0.00152174
R7178 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 0.00152174
R7179 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 0.00152174
R7180 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 0.00152174
R7181 two_stage_opamp_dummy_magic_14_0.X.n47 two_stage_opamp_dummy_magic_14_0.X.t43 1172.87
R7182 two_stage_opamp_dummy_magic_14_0.X.n43 two_stage_opamp_dummy_magic_14_0.X.t48 1172.87
R7183 two_stage_opamp_dummy_magic_14_0.X.n50 two_stage_opamp_dummy_magic_14_0.X.t46 996.134
R7184 two_stage_opamp_dummy_magic_14_0.X.n49 two_stage_opamp_dummy_magic_14_0.X.t33 996.134
R7185 two_stage_opamp_dummy_magic_14_0.X.n48 two_stage_opamp_dummy_magic_14_0.X.t50 996.134
R7186 two_stage_opamp_dummy_magic_14_0.X.n47 two_stage_opamp_dummy_magic_14_0.X.t28 996.134
R7187 two_stage_opamp_dummy_magic_14_0.X.n43 two_stage_opamp_dummy_magic_14_0.X.t35 996.134
R7188 two_stage_opamp_dummy_magic_14_0.X.n44 two_stage_opamp_dummy_magic_14_0.X.t51 996.134
R7189 two_stage_opamp_dummy_magic_14_0.X.n45 two_stage_opamp_dummy_magic_14_0.X.t39 996.134
R7190 two_stage_opamp_dummy_magic_14_0.X.n46 two_stage_opamp_dummy_magic_14_0.X.t31 996.134
R7191 two_stage_opamp_dummy_magic_14_0.X.n37 two_stage_opamp_dummy_magic_14_0.X.t47 690.867
R7192 two_stage_opamp_dummy_magic_14_0.X.n32 two_stage_opamp_dummy_magic_14_0.X.t25 690.867
R7193 two_stage_opamp_dummy_magic_14_0.X.n28 two_stage_opamp_dummy_magic_14_0.X.t30 530.201
R7194 two_stage_opamp_dummy_magic_14_0.X.n23 two_stage_opamp_dummy_magic_14_0.X.t36 530.201
R7195 two_stage_opamp_dummy_magic_14_0.X.n37 two_stage_opamp_dummy_magic_14_0.X.t32 514.134
R7196 two_stage_opamp_dummy_magic_14_0.X.n38 two_stage_opamp_dummy_magic_14_0.X.t27 514.134
R7197 two_stage_opamp_dummy_magic_14_0.X.n39 two_stage_opamp_dummy_magic_14_0.X.t41 514.134
R7198 two_stage_opamp_dummy_magic_14_0.X.n36 two_stage_opamp_dummy_magic_14_0.X.t54 514.134
R7199 two_stage_opamp_dummy_magic_14_0.X.n35 two_stage_opamp_dummy_magic_14_0.X.t37 514.134
R7200 two_stage_opamp_dummy_magic_14_0.X.n34 two_stage_opamp_dummy_magic_14_0.X.t44 514.134
R7201 two_stage_opamp_dummy_magic_14_0.X.n33 two_stage_opamp_dummy_magic_14_0.X.t29 514.134
R7202 two_stage_opamp_dummy_magic_14_0.X.n32 two_stage_opamp_dummy_magic_14_0.X.t42 514.134
R7203 two_stage_opamp_dummy_magic_14_0.X.n30 two_stage_opamp_dummy_magic_14_0.X.t52 353.467
R7204 two_stage_opamp_dummy_magic_14_0.X.n29 two_stage_opamp_dummy_magic_14_0.X.t38 353.467
R7205 two_stage_opamp_dummy_magic_14_0.X.n28 two_stage_opamp_dummy_magic_14_0.X.t45 353.467
R7206 two_stage_opamp_dummy_magic_14_0.X.n23 two_stage_opamp_dummy_magic_14_0.X.t53 353.467
R7207 two_stage_opamp_dummy_magic_14_0.X.n24 two_stage_opamp_dummy_magic_14_0.X.t40 353.467
R7208 two_stage_opamp_dummy_magic_14_0.X.n25 two_stage_opamp_dummy_magic_14_0.X.t26 353.467
R7209 two_stage_opamp_dummy_magic_14_0.X.n26 two_stage_opamp_dummy_magic_14_0.X.t49 353.467
R7210 two_stage_opamp_dummy_magic_14_0.X.n27 two_stage_opamp_dummy_magic_14_0.X.t34 353.467
R7211 two_stage_opamp_dummy_magic_14_0.X.n50 two_stage_opamp_dummy_magic_14_0.X.n49 176.733
R7212 two_stage_opamp_dummy_magic_14_0.X.n49 two_stage_opamp_dummy_magic_14_0.X.n48 176.733
R7213 two_stage_opamp_dummy_magic_14_0.X.n48 two_stage_opamp_dummy_magic_14_0.X.n47 176.733
R7214 two_stage_opamp_dummy_magic_14_0.X.n44 two_stage_opamp_dummy_magic_14_0.X.n43 176.733
R7215 two_stage_opamp_dummy_magic_14_0.X.n45 two_stage_opamp_dummy_magic_14_0.X.n44 176.733
R7216 two_stage_opamp_dummy_magic_14_0.X.n46 two_stage_opamp_dummy_magic_14_0.X.n45 176.733
R7217 two_stage_opamp_dummy_magic_14_0.X.n30 two_stage_opamp_dummy_magic_14_0.X.n29 176.733
R7218 two_stage_opamp_dummy_magic_14_0.X.n29 two_stage_opamp_dummy_magic_14_0.X.n28 176.733
R7219 two_stage_opamp_dummy_magic_14_0.X.n24 two_stage_opamp_dummy_magic_14_0.X.n23 176.733
R7220 two_stage_opamp_dummy_magic_14_0.X.n25 two_stage_opamp_dummy_magic_14_0.X.n24 176.733
R7221 two_stage_opamp_dummy_magic_14_0.X.n26 two_stage_opamp_dummy_magic_14_0.X.n25 176.733
R7222 two_stage_opamp_dummy_magic_14_0.X.n27 two_stage_opamp_dummy_magic_14_0.X.n26 176.733
R7223 two_stage_opamp_dummy_magic_14_0.X.n39 two_stage_opamp_dummy_magic_14_0.X.n38 176.733
R7224 two_stage_opamp_dummy_magic_14_0.X.n38 two_stage_opamp_dummy_magic_14_0.X.n37 176.733
R7225 two_stage_opamp_dummy_magic_14_0.X.n33 two_stage_opamp_dummy_magic_14_0.X.n32 176.733
R7226 two_stage_opamp_dummy_magic_14_0.X.n34 two_stage_opamp_dummy_magic_14_0.X.n33 176.733
R7227 two_stage_opamp_dummy_magic_14_0.X.n35 two_stage_opamp_dummy_magic_14_0.X.n34 176.733
R7228 two_stage_opamp_dummy_magic_14_0.X.n36 two_stage_opamp_dummy_magic_14_0.X.n35 176.733
R7229 two_stage_opamp_dummy_magic_14_0.X.n52 two_stage_opamp_dummy_magic_14_0.X.n51 166.258
R7230 two_stage_opamp_dummy_magic_14_0.X.n2 two_stage_opamp_dummy_magic_14_0.X.n0 163.626
R7231 two_stage_opamp_dummy_magic_14_0.X.n8 two_stage_opamp_dummy_magic_14_0.X.n7 163.001
R7232 two_stage_opamp_dummy_magic_14_0.X.n6 two_stage_opamp_dummy_magic_14_0.X.n5 163.001
R7233 two_stage_opamp_dummy_magic_14_0.X.n4 two_stage_opamp_dummy_magic_14_0.X.n3 163.001
R7234 two_stage_opamp_dummy_magic_14_0.X.n2 two_stage_opamp_dummy_magic_14_0.X.n1 163.001
R7235 two_stage_opamp_dummy_magic_14_0.X.n41 two_stage_opamp_dummy_magic_14_0.X.n31 161.541
R7236 two_stage_opamp_dummy_magic_14_0.X.n41 two_stage_opamp_dummy_magic_14_0.X.n40 161.541
R7237 two_stage_opamp_dummy_magic_14_0.X.n10 two_stage_opamp_dummy_magic_14_0.X.n9 158.501
R7238 two_stage_opamp_dummy_magic_14_0.X.n13 two_stage_opamp_dummy_magic_14_0.X.n11 117.888
R7239 two_stage_opamp_dummy_magic_14_0.X.n21 two_stage_opamp_dummy_magic_14_0.X.n20 117.326
R7240 two_stage_opamp_dummy_magic_14_0.X.n19 two_stage_opamp_dummy_magic_14_0.X.n18 117.326
R7241 two_stage_opamp_dummy_magic_14_0.X.n17 two_stage_opamp_dummy_magic_14_0.X.n16 117.326
R7242 two_stage_opamp_dummy_magic_14_0.X.n15 two_stage_opamp_dummy_magic_14_0.X.n14 117.326
R7243 two_stage_opamp_dummy_magic_14_0.X.n13 two_stage_opamp_dummy_magic_14_0.X.n12 117.326
R7244 two_stage_opamp_dummy_magic_14_0.X.n31 two_stage_opamp_dummy_magic_14_0.X.n30 54.6272
R7245 two_stage_opamp_dummy_magic_14_0.X.n31 two_stage_opamp_dummy_magic_14_0.X.n27 54.6272
R7246 two_stage_opamp_dummy_magic_14_0.X.n40 two_stage_opamp_dummy_magic_14_0.X.n39 54.6272
R7247 two_stage_opamp_dummy_magic_14_0.X.n40 two_stage_opamp_dummy_magic_14_0.X.n36 54.6272
R7248 two_stage_opamp_dummy_magic_14_0.X.n51 two_stage_opamp_dummy_magic_14_0.X.n50 53.3126
R7249 two_stage_opamp_dummy_magic_14_0.X.n51 two_stage_opamp_dummy_magic_14_0.X.n46 53.3126
R7250 two_stage_opamp_dummy_magic_14_0.X.t15 two_stage_opamp_dummy_magic_14_0.X.n52 49.8023
R7251 two_stage_opamp_dummy_magic_14_0.X.n20 two_stage_opamp_dummy_magic_14_0.X.t16 16.0005
R7252 two_stage_opamp_dummy_magic_14_0.X.n20 two_stage_opamp_dummy_magic_14_0.X.t24 16.0005
R7253 two_stage_opamp_dummy_magic_14_0.X.n18 two_stage_opamp_dummy_magic_14_0.X.t2 16.0005
R7254 two_stage_opamp_dummy_magic_14_0.X.n18 two_stage_opamp_dummy_magic_14_0.X.t19 16.0005
R7255 two_stage_opamp_dummy_magic_14_0.X.n16 two_stage_opamp_dummy_magic_14_0.X.t3 16.0005
R7256 two_stage_opamp_dummy_magic_14_0.X.n16 two_stage_opamp_dummy_magic_14_0.X.t9 16.0005
R7257 two_stage_opamp_dummy_magic_14_0.X.n14 two_stage_opamp_dummy_magic_14_0.X.t8 16.0005
R7258 two_stage_opamp_dummy_magic_14_0.X.n14 two_stage_opamp_dummy_magic_14_0.X.t13 16.0005
R7259 two_stage_opamp_dummy_magic_14_0.X.n12 two_stage_opamp_dummy_magic_14_0.X.t18 16.0005
R7260 two_stage_opamp_dummy_magic_14_0.X.n12 two_stage_opamp_dummy_magic_14_0.X.t10 16.0005
R7261 two_stage_opamp_dummy_magic_14_0.X.n11 two_stage_opamp_dummy_magic_14_0.X.t1 16.0005
R7262 two_stage_opamp_dummy_magic_14_0.X.n11 two_stage_opamp_dummy_magic_14_0.X.t17 16.0005
R7263 two_stage_opamp_dummy_magic_14_0.X.n22 two_stage_opamp_dummy_magic_14_0.X.n10 15.8443
R7264 two_stage_opamp_dummy_magic_14_0.X.n42 two_stage_opamp_dummy_magic_14_0.X.n41 13.4693
R7265 two_stage_opamp_dummy_magic_14_0.X.n9 two_stage_opamp_dummy_magic_14_0.X.t11 11.2576
R7266 two_stage_opamp_dummy_magic_14_0.X.n9 two_stage_opamp_dummy_magic_14_0.X.t14 11.2576
R7267 two_stage_opamp_dummy_magic_14_0.X.n7 two_stage_opamp_dummy_magic_14_0.X.t21 11.2576
R7268 two_stage_opamp_dummy_magic_14_0.X.n7 two_stage_opamp_dummy_magic_14_0.X.t6 11.2576
R7269 two_stage_opamp_dummy_magic_14_0.X.n5 two_stage_opamp_dummy_magic_14_0.X.t0 11.2576
R7270 two_stage_opamp_dummy_magic_14_0.X.n5 two_stage_opamp_dummy_magic_14_0.X.t22 11.2576
R7271 two_stage_opamp_dummy_magic_14_0.X.n3 two_stage_opamp_dummy_magic_14_0.X.t20 11.2576
R7272 two_stage_opamp_dummy_magic_14_0.X.n3 two_stage_opamp_dummy_magic_14_0.X.t4 11.2576
R7273 two_stage_opamp_dummy_magic_14_0.X.n1 two_stage_opamp_dummy_magic_14_0.X.t23 11.2576
R7274 two_stage_opamp_dummy_magic_14_0.X.n1 two_stage_opamp_dummy_magic_14_0.X.t7 11.2576
R7275 two_stage_opamp_dummy_magic_14_0.X.n0 two_stage_opamp_dummy_magic_14_0.X.t5 11.2576
R7276 two_stage_opamp_dummy_magic_14_0.X.n0 two_stage_opamp_dummy_magic_14_0.X.t12 11.2576
R7277 two_stage_opamp_dummy_magic_14_0.X.n52 two_stage_opamp_dummy_magic_14_0.X.n42 7.09425
R7278 two_stage_opamp_dummy_magic_14_0.X.n22 two_stage_opamp_dummy_magic_14_0.X.n21 6.3755
R7279 two_stage_opamp_dummy_magic_14_0.X.n10 two_stage_opamp_dummy_magic_14_0.X.n8 5.1255
R7280 two_stage_opamp_dummy_magic_14_0.X.n42 two_stage_opamp_dummy_magic_14_0.X.n22 1.40675
R7281 two_stage_opamp_dummy_magic_14_0.X.n4 two_stage_opamp_dummy_magic_14_0.X.n2 0.6255
R7282 two_stage_opamp_dummy_magic_14_0.X.n6 two_stage_opamp_dummy_magic_14_0.X.n4 0.6255
R7283 two_stage_opamp_dummy_magic_14_0.X.n8 two_stage_opamp_dummy_magic_14_0.X.n6 0.6255
R7284 two_stage_opamp_dummy_magic_14_0.X.n15 two_stage_opamp_dummy_magic_14_0.X.n13 0.563
R7285 two_stage_opamp_dummy_magic_14_0.X.n17 two_stage_opamp_dummy_magic_14_0.X.n15 0.563
R7286 two_stage_opamp_dummy_magic_14_0.X.n19 two_stage_opamp_dummy_magic_14_0.X.n17 0.563
R7287 two_stage_opamp_dummy_magic_14_0.X.n21 two_stage_opamp_dummy_magic_14_0.X.n19 0.563
R7288 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 144.827
R7289 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 134.577
R7290 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 118.986
R7291 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 100.6
R7292 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 100.038
R7293 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 100.038
R7294 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 100.038
R7295 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 100.038
R7296 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 37.4067
R7297 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 33.705
R7298 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 24.0005
R7299 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 24.0005
R7300 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 24.0005
R7301 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 24.0005
R7302 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 8.0005
R7303 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 8.0005
R7304 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 8.0005
R7305 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 8.0005
R7306 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 8.0005
R7307 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 8.0005
R7308 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 8.0005
R7309 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 8.0005
R7310 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 8.0005
R7311 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 8.0005
R7312 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 5.6255
R7313 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 0.563
R7314 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 0.563
R7315 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 0.563
R7316 bgr_7_0.V_CMFB_S2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 0.047375
R7317 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 525.38
R7318 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 525.38
R7319 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 358.288
R7320 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 358.288
R7321 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 281.168
R7322 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 281.168
R7323 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 281.168
R7324 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 281.168
R7325 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 244.214
R7326 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 244.214
R7327 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 166.019
R7328 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 166.019
R7329 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 116.013
R7330 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 116.013
R7331 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 77.1205
R7332 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 77.1205
R7333 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 36.8755
R7334 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 688.859
R7335 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 651.343
R7336 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 647.968
R7337 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 514.134
R7338 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 214.056
R7339 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 174.726
R7340 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 174.726
R7341 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 174.726
R7342 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 174.726
R7343 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 173.591
R7344 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 169.216
R7345 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 169.216
R7346 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 128.534
R7347 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 128.534
R7348 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 125.736
R7349 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 46.6411
R7350 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 13.1338
R7351 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 13.1338
R7352 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 13.1338
R7353 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 13.1338
R7354 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 13.1338
R7355 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 13.1338
R7356 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 10.0317
R7357 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 4.3755
R7358 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 3.03175
R7359 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 1.53175
R7360 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 two_stage_opamp_dummy_magic_14_0.err_amp_out.t4 686.271
R7361 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 179.195
R7362 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 101.055
R7363 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 two_stage_opamp_dummy_magic_14_0.err_amp_out.t0 15.7605
R7364 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 two_stage_opamp_dummy_magic_14_0.err_amp_out.t3 15.7605
R7365 two_stage_opamp_dummy_magic_14_0.err_amp_out.t1 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 9.6005
R7366 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 two_stage_opamp_dummy_magic_14_0.err_amp_out.t2 9.6005
R7367 bgr_7_0.Vin+.n3 bgr_7_0.Vin+.n2 526.183
R7368 bgr_7_0.Vin+.n1 bgr_7_0.Vin+.n0 514.134
R7369 bgr_7_0.Vin+.n0 bgr_7_0.Vin+.t8 303.259
R7370 bgr_7_0.Vin+.n5 bgr_7_0.Vin+.n3 227.169
R7371 bgr_7_0.Vin+.n0 bgr_7_0.Vin+.t9 174.726
R7372 bgr_7_0.Vin+.n1 bgr_7_0.Vin+.t6 174.726
R7373 bgr_7_0.Vin+.n2 bgr_7_0.Vin+.t10 174.726
R7374 bgr_7_0.Vin+.n7 bgr_7_0.Vin+.n6 168.435
R7375 bgr_7_0.Vin+.n5 bgr_7_0.Vin+.n4 168.435
R7376 bgr_7_0.Vin+.n8 bgr_7_0.Vin+.t1 158.989
R7377 bgr_7_0.Vin+.n2 bgr_7_0.Vin+.n1 128.534
R7378 bgr_7_0.Vin+.t0 bgr_7_0.Vin+.n8 119.067
R7379 bgr_7_0.Vin+.n3 bgr_7_0.Vin+.t7 96.4005
R7380 bgr_7_0.Vin+.n8 bgr_7_0.Vin+.n7 35.0317
R7381 bgr_7_0.Vin+.n6 bgr_7_0.Vin+.t2 13.1338
R7382 bgr_7_0.Vin+.n6 bgr_7_0.Vin+.t5 13.1338
R7383 bgr_7_0.Vin+.n4 bgr_7_0.Vin+.t4 13.1338
R7384 bgr_7_0.Vin+.n4 bgr_7_0.Vin+.t3 13.1338
R7385 bgr_7_0.Vin+.n7 bgr_7_0.Vin+.n5 2.1255
R7386 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 344.837
R7387 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 344.274
R7388 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 292.5
R7389 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 209.251
R7390 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 208.689
R7391 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 208.689
R7392 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 208.689
R7393 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 208.689
R7394 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 120.305
R7395 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 52.3363
R7396 bgr_7_0.V_CMFB_S1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 52.1563
R7397 bgr_7_0.V_CMFB_S1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 41.2477
R7398 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 39.4005
R7399 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 39.4005
R7400 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 39.4005
R7401 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 39.4005
R7402 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 39.4005
R7403 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 39.4005
R7404 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 19.7005
R7405 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 19.7005
R7406 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 19.7005
R7407 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 19.7005
R7408 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 19.7005
R7409 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 19.7005
R7410 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 19.7005
R7411 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 19.7005
R7412 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 19.7005
R7413 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 19.7005
R7414 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 5.90675
R7415 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 0.563
R7416 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 0.563
R7417 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 0.563
R7418 bgr_7_0.V_mir1.n20 bgr_7_0.V_mir1.n19 325.473
R7419 bgr_7_0.V_mir1.n13 bgr_7_0.V_mir1.n12 325.473
R7420 bgr_7_0.V_mir1.n4 bgr_7_0.V_mir1.n3 325.473
R7421 bgr_7_0.V_mir1.n16 bgr_7_0.V_mir1.t19 310.488
R7422 bgr_7_0.V_mir1.n9 bgr_7_0.V_mir1.t21 310.488
R7423 bgr_7_0.V_mir1.n0 bgr_7_0.V_mir1.t20 310.488
R7424 bgr_7_0.V_mir1.n7 bgr_7_0.V_mir1.t0 278.312
R7425 bgr_7_0.V_mir1.n7 bgr_7_0.V_mir1.n6 228.939
R7426 bgr_7_0.V_mir1.n8 bgr_7_0.V_mir1.n5 224.439
R7427 bgr_7_0.V_mir1.n18 bgr_7_0.V_mir1.t11 184.097
R7428 bgr_7_0.V_mir1.n11 bgr_7_0.V_mir1.t7 184.097
R7429 bgr_7_0.V_mir1.n2 bgr_7_0.V_mir1.t5 184.097
R7430 bgr_7_0.V_mir1.n17 bgr_7_0.V_mir1.n16 167.094
R7431 bgr_7_0.V_mir1.n10 bgr_7_0.V_mir1.n9 167.094
R7432 bgr_7_0.V_mir1.n1 bgr_7_0.V_mir1.n0 167.094
R7433 bgr_7_0.V_mir1.n13 bgr_7_0.V_mir1.n11 152
R7434 bgr_7_0.V_mir1.n4 bgr_7_0.V_mir1.n2 152
R7435 bgr_7_0.V_mir1.n19 bgr_7_0.V_mir1.n18 152
R7436 bgr_7_0.V_mir1.n16 bgr_7_0.V_mir1.t22 120.501
R7437 bgr_7_0.V_mir1.n17 bgr_7_0.V_mir1.t15 120.501
R7438 bgr_7_0.V_mir1.n9 bgr_7_0.V_mir1.t17 120.501
R7439 bgr_7_0.V_mir1.n10 bgr_7_0.V_mir1.t13 120.501
R7440 bgr_7_0.V_mir1.n0 bgr_7_0.V_mir1.t18 120.501
R7441 bgr_7_0.V_mir1.n1 bgr_7_0.V_mir1.t9 120.501
R7442 bgr_7_0.V_mir1.n6 bgr_7_0.V_mir1.t4 48.0005
R7443 bgr_7_0.V_mir1.n6 bgr_7_0.V_mir1.t3 48.0005
R7444 bgr_7_0.V_mir1.n5 bgr_7_0.V_mir1.t2 48.0005
R7445 bgr_7_0.V_mir1.n5 bgr_7_0.V_mir1.t1 48.0005
R7446 bgr_7_0.V_mir1.n18 bgr_7_0.V_mir1.n17 40.7027
R7447 bgr_7_0.V_mir1.n11 bgr_7_0.V_mir1.n10 40.7027
R7448 bgr_7_0.V_mir1.n2 bgr_7_0.V_mir1.n1 40.7027
R7449 bgr_7_0.V_mir1.n12 bgr_7_0.V_mir1.t8 39.4005
R7450 bgr_7_0.V_mir1.n12 bgr_7_0.V_mir1.t14 39.4005
R7451 bgr_7_0.V_mir1.n3 bgr_7_0.V_mir1.t6 39.4005
R7452 bgr_7_0.V_mir1.n3 bgr_7_0.V_mir1.t10 39.4005
R7453 bgr_7_0.V_mir1.n20 bgr_7_0.V_mir1.t12 39.4005
R7454 bgr_7_0.V_mir1.t16 bgr_7_0.V_mir1.n20 39.4005
R7455 bgr_7_0.V_mir1.n15 bgr_7_0.V_mir1.n4 15.8005
R7456 bgr_7_0.V_mir1.n19 bgr_7_0.V_mir1.n15 15.8005
R7457 bgr_7_0.V_mir1.n14 bgr_7_0.V_mir1.n13 9.3005
R7458 bgr_7_0.V_mir1.n8 bgr_7_0.V_mir1.n7 5.8755
R7459 bgr_7_0.V_mir1.n15 bgr_7_0.V_mir1.n14 4.5005
R7460 bgr_7_0.V_mir1.n14 bgr_7_0.V_mir1.n8 0.78175
R7461 bgr_7_0.1st_Vout_1 bgr_7_0.1st_Vout_1.t13 354.854
R7462 bgr_7_0.1st_Vout_1.n5 bgr_7_0.1st_Vout_1.t21 346.8
R7463 bgr_7_0.1st_Vout_1.n20 bgr_7_0.1st_Vout_1.n19 339.522
R7464 bgr_7_0.1st_Vout_1.n7 bgr_7_0.1st_Vout_1.n6 339.522
R7465 bgr_7_0.1st_Vout_1.n15 bgr_7_0.1st_Vout_1.n14 335.022
R7466 bgr_7_0.1st_Vout_1.n11 bgr_7_0.1st_Vout_1.t10 275.909
R7467 bgr_7_0.1st_Vout_1.n11 bgr_7_0.1st_Vout_1.n10 227.909
R7468 bgr_7_0.1st_Vout_1.n13 bgr_7_0.1st_Vout_1.n12 222.034
R7469 bgr_7_0.1st_Vout_1.n17 bgr_7_0.1st_Vout_1.t22 184.097
R7470 bgr_7_0.1st_Vout_1.n17 bgr_7_0.1st_Vout_1.t32 184.097
R7471 bgr_7_0.1st_Vout_1.n8 bgr_7_0.1st_Vout_1.t16 184.097
R7472 bgr_7_0.1st_Vout_1.n8 bgr_7_0.1st_Vout_1.t36 184.097
R7473 bgr_7_0.1st_Vout_1.n18 bgr_7_0.1st_Vout_1.n17 166.05
R7474 bgr_7_0.1st_Vout_1.n9 bgr_7_0.1st_Vout_1.n8 166.05
R7475 bgr_7_0.1st_Vout_1.n5 bgr_7_0.1st_Vout_1.n4 54.2759
R7476 bgr_7_0.1st_Vout_1.n12 bgr_7_0.1st_Vout_1.t6 48.0005
R7477 bgr_7_0.1st_Vout_1.n12 bgr_7_0.1st_Vout_1.t8 48.0005
R7478 bgr_7_0.1st_Vout_1.n10 bgr_7_0.1st_Vout_1.t7 48.0005
R7479 bgr_7_0.1st_Vout_1.n10 bgr_7_0.1st_Vout_1.t9 48.0005
R7480 bgr_7_0.1st_Vout_1.n19 bgr_7_0.1st_Vout_1.t4 39.4005
R7481 bgr_7_0.1st_Vout_1.n19 bgr_7_0.1st_Vout_1.t2 39.4005
R7482 bgr_7_0.1st_Vout_1.n6 bgr_7_0.1st_Vout_1.t0 39.4005
R7483 bgr_7_0.1st_Vout_1.n6 bgr_7_0.1st_Vout_1.t3 39.4005
R7484 bgr_7_0.1st_Vout_1.n14 bgr_7_0.1st_Vout_1.t5 39.4005
R7485 bgr_7_0.1st_Vout_1.n14 bgr_7_0.1st_Vout_1.t1 39.4005
R7486 bgr_7_0.1st_Vout_1.n0 bgr_7_0.1st_Vout_1.t11 4.8295
R7487 bgr_7_0.1st_Vout_1.n0 bgr_7_0.1st_Vout_1.t29 4.8295
R7488 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t31 4.8295
R7489 bgr_7_0.1st_Vout_1.n1 bgr_7_0.1st_Vout_1.t20 4.8295
R7490 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t24 4.8295
R7491 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t14 4.8295
R7492 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t30 4.8295
R7493 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t18 4.8295
R7494 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t23 4.8295
R7495 bgr_7_0.1st_Vout_1.n0 bgr_7_0.1st_Vout_1.t15 4.5005
R7496 bgr_7_0.1st_Vout_1.n0 bgr_7_0.1st_Vout_1.t35 4.5005
R7497 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t34 4.5005
R7498 bgr_7_0.1st_Vout_1.n1 bgr_7_0.1st_Vout_1.t28 4.5005
R7499 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t27 4.5005
R7500 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.t19 4.5005
R7501 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t33 4.5005
R7502 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t26 4.5005
R7503 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.t25 4.5005
R7504 bgr_7_0.1st_Vout_1.n4 bgr_7_0.1st_Vout_1.t17 4.5005
R7505 bgr_7_0.1st_Vout_1.n4 bgr_7_0.1st_Vout_1.t12 4.5005
R7506 bgr_7_0.1st_Vout_1.n13 bgr_7_0.1st_Vout_1.n11 4.5005
R7507 bgr_7_0.1st_Vout_1.n16 bgr_7_0.1st_Vout_1.n15 4.5005
R7508 bgr_7_0.1st_Vout_1.n20 bgr_7_0.1st_Vout_1.n18 1.3755
R7509 bgr_7_0.1st_Vout_1.n16 bgr_7_0.1st_Vout_1.n9 1.3755
R7510 bgr_7_0.1st_Vout_1.n7 bgr_7_0.1st_Vout_1.n5 1.188
R7511 bgr_7_0.1st_Vout_1.n3 bgr_7_0.1st_Vout_1.n2 0.8935
R7512 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.n0 0.8935
R7513 bgr_7_0.1st_Vout_1.n15 bgr_7_0.1st_Vout_1.n13 0.78175
R7514 bgr_7_0.1st_Vout_1.n4 bgr_7_0.1st_Vout_1.n3 0.6585
R7515 bgr_7_0.1st_Vout_1.n2 bgr_7_0.1st_Vout_1.n1 0.6585
R7516 bgr_7_0.1st_Vout_1.n18 bgr_7_0.1st_Vout_1.n16 0.6255
R7517 bgr_7_0.1st_Vout_1.n9 bgr_7_0.1st_Vout_1.n7 0.6255
R7518 bgr_7_0.1st_Vout_1 bgr_7_0.1st_Vout_1.n20 0.438
R7519 bgr_7_0.1st_Vout_2.n0 bgr_7_0.1st_Vout_2.t33 355.293
R7520 bgr_7_0.1st_Vout_2.n1 bgr_7_0.1st_Vout_2.t34 346.8
R7521 bgr_7_0.1st_Vout_2.n12 bgr_7_0.1st_Vout_2.n1 339.522
R7522 bgr_7_0.1st_Vout_2.n0 bgr_7_0.1st_Vout_2.n5 339.522
R7523 bgr_7_0.1st_Vout_2.n3 bgr_7_0.1st_Vout_2.n10 335.022
R7524 bgr_7_0.1st_Vout_2.n8 bgr_7_0.1st_Vout_2.t10 275.909
R7525 bgr_7_0.1st_Vout_2.n8 bgr_7_0.1st_Vout_2.n7 227.909
R7526 bgr_7_0.1st_Vout_2.n3 bgr_7_0.1st_Vout_2.n9 222.034
R7527 bgr_7_0.1st_Vout_2.n11 bgr_7_0.1st_Vout_2.t16 184.097
R7528 bgr_7_0.1st_Vout_2.n11 bgr_7_0.1st_Vout_2.t27 184.097
R7529 bgr_7_0.1st_Vout_2.n6 bgr_7_0.1st_Vout_2.t13 184.097
R7530 bgr_7_0.1st_Vout_2.n6 bgr_7_0.1st_Vout_2.t24 184.097
R7531 bgr_7_0.1st_Vout_2.n1 bgr_7_0.1st_Vout_2.n11 166.05
R7532 bgr_7_0.1st_Vout_2.n0 bgr_7_0.1st_Vout_2.n6 166.05
R7533 bgr_7_0.1st_Vout_2.n1 bgr_7_0.1st_Vout_2.n4 52.9634
R7534 bgr_7_0.1st_Vout_2.n9 bgr_7_0.1st_Vout_2.t9 48.0005
R7535 bgr_7_0.1st_Vout_2.n9 bgr_7_0.1st_Vout_2.t1 48.0005
R7536 bgr_7_0.1st_Vout_2.n7 bgr_7_0.1st_Vout_2.t6 48.0005
R7537 bgr_7_0.1st_Vout_2.n7 bgr_7_0.1st_Vout_2.t2 48.0005
R7538 bgr_7_0.1st_Vout_2.n10 bgr_7_0.1st_Vout_2.t3 39.4005
R7539 bgr_7_0.1st_Vout_2.n10 bgr_7_0.1st_Vout_2.t5 39.4005
R7540 bgr_7_0.1st_Vout_2.n5 bgr_7_0.1st_Vout_2.t7 39.4005
R7541 bgr_7_0.1st_Vout_2.n5 bgr_7_0.1st_Vout_2.t4 39.4005
R7542 bgr_7_0.1st_Vout_2.n12 bgr_7_0.1st_Vout_2.t8 39.4005
R7543 bgr_7_0.1st_Vout_2.t0 bgr_7_0.1st_Vout_2.n12 39.4005
R7544 bgr_7_0.1st_Vout_2.n0 bgr_7_0.1st_Vout_2.n3 5.28175
R7545 bgr_7_0.1st_Vout_2.n1 bgr_7_0.1st_Vout_2.n0 5.188
R7546 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t17 4.8295
R7547 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t35 4.8295
R7548 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t11 4.8295
R7549 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t26 4.8295
R7550 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t30 4.8295
R7551 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t19 4.8295
R7552 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t36 4.8295
R7553 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t25 4.8295
R7554 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t18 4.8295
R7555 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t12 4.5005
R7556 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t32 4.5005
R7557 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t31 4.5005
R7558 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t23 4.5005
R7559 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t22 4.5005
R7560 bgr_7_0.1st_Vout_2.n2 bgr_7_0.1st_Vout_2.t15 4.5005
R7561 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t29 4.5005
R7562 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t21 4.5005
R7563 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t28 4.5005
R7564 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t20 4.5005
R7565 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.t14 4.5005
R7566 bgr_7_0.1st_Vout_2.n3 bgr_7_0.1st_Vout_2.n8 4.5005
R7567 bgr_7_0.1st_Vout_2.n4 bgr_7_0.1st_Vout_2.n2 3.1025
R7568 bgr_7_0.cap_res2.t20 bgr_7_0.cap_res2.t17 121.245
R7569 bgr_7_0.cap_res2.t12 bgr_7_0.cap_res2.t6 0.1603
R7570 bgr_7_0.cap_res2.t5 bgr_7_0.cap_res2.t0 0.1603
R7571 bgr_7_0.cap_res2.t10 bgr_7_0.cap_res2.t4 0.1603
R7572 bgr_7_0.cap_res2.t3 bgr_7_0.cap_res2.t19 0.1603
R7573 bgr_7_0.cap_res2.t18 bgr_7_0.cap_res2.t15 0.1603
R7574 bgr_7_0.cap_res2.n1 bgr_7_0.cap_res2.t2 0.159278
R7575 bgr_7_0.cap_res2.n2 bgr_7_0.cap_res2.t9 0.159278
R7576 bgr_7_0.cap_res2.n3 bgr_7_0.cap_res2.t16 0.159278
R7577 bgr_7_0.cap_res2.n4 bgr_7_0.cap_res2.t11 0.159278
R7578 bgr_7_0.cap_res2.n4 bgr_7_0.cap_res2.t14 0.1368
R7579 bgr_7_0.cap_res2.n4 bgr_7_0.cap_res2.t12 0.1368
R7580 bgr_7_0.cap_res2.n3 bgr_7_0.cap_res2.t8 0.1368
R7581 bgr_7_0.cap_res2.n3 bgr_7_0.cap_res2.t5 0.1368
R7582 bgr_7_0.cap_res2.n2 bgr_7_0.cap_res2.t13 0.1368
R7583 bgr_7_0.cap_res2.n2 bgr_7_0.cap_res2.t10 0.1368
R7584 bgr_7_0.cap_res2.n1 bgr_7_0.cap_res2.t7 0.1368
R7585 bgr_7_0.cap_res2.n1 bgr_7_0.cap_res2.t3 0.1368
R7586 bgr_7_0.cap_res2.n0 bgr_7_0.cap_res2.t1 0.1368
R7587 bgr_7_0.cap_res2.n0 bgr_7_0.cap_res2.t18 0.1368
R7588 bgr_7_0.cap_res2.t2 bgr_7_0.cap_res2.n0 0.00152174
R7589 bgr_7_0.cap_res2.t9 bgr_7_0.cap_res2.n1 0.00152174
R7590 bgr_7_0.cap_res2.t16 bgr_7_0.cap_res2.n2 0.00152174
R7591 bgr_7_0.cap_res2.t11 bgr_7_0.cap_res2.n3 0.00152174
R7592 bgr_7_0.cap_res2.t17 bgr_7_0.cap_res2.n4 0.00152174
R7593 two_stage_opamp_dummy_magic_14_0.Vb2.n25 two_stage_opamp_dummy_magic_14_0.Vb2.t31 650.273
R7594 two_stage_opamp_dummy_magic_14_0.Vb2.n27 two_stage_opamp_dummy_magic_14_0.Vb2.t0 650.273
R7595 two_stage_opamp_dummy_magic_14_0.Vb2.n4 two_stage_opamp_dummy_magic_14_0.Vb2.t12 611.739
R7596 two_stage_opamp_dummy_magic_14_0.Vb2.n0 two_stage_opamp_dummy_magic_14_0.Vb2.t22 611.739
R7597 two_stage_opamp_dummy_magic_14_0.Vb2.n13 two_stage_opamp_dummy_magic_14_0.Vb2.t13 611.739
R7598 two_stage_opamp_dummy_magic_14_0.Vb2.n9 two_stage_opamp_dummy_magic_14_0.Vb2.t23 611.739
R7599 two_stage_opamp_dummy_magic_14_0.Vb2.n28 two_stage_opamp_dummy_magic_14_0.Vb2.t27 445.423
R7600 two_stage_opamp_dummy_magic_14_0.Vb2.n4 two_stage_opamp_dummy_magic_14_0.Vb2.t17 421.75
R7601 two_stage_opamp_dummy_magic_14_0.Vb2.n5 two_stage_opamp_dummy_magic_14_0.Vb2.t24 421.75
R7602 two_stage_opamp_dummy_magic_14_0.Vb2.n6 two_stage_opamp_dummy_magic_14_0.Vb2.t28 421.75
R7603 two_stage_opamp_dummy_magic_14_0.Vb2.n7 two_stage_opamp_dummy_magic_14_0.Vb2.t29 421.75
R7604 two_stage_opamp_dummy_magic_14_0.Vb2.n0 two_stage_opamp_dummy_magic_14_0.Vb2.t26 421.75
R7605 two_stage_opamp_dummy_magic_14_0.Vb2.n1 two_stage_opamp_dummy_magic_14_0.Vb2.t19 421.75
R7606 two_stage_opamp_dummy_magic_14_0.Vb2.n2 two_stage_opamp_dummy_magic_14_0.Vb2.t14 421.75
R7607 two_stage_opamp_dummy_magic_14_0.Vb2.n3 two_stage_opamp_dummy_magic_14_0.Vb2.t32 421.75
R7608 two_stage_opamp_dummy_magic_14_0.Vb2.n13 two_stage_opamp_dummy_magic_14_0.Vb2.t18 421.75
R7609 two_stage_opamp_dummy_magic_14_0.Vb2.n14 two_stage_opamp_dummy_magic_14_0.Vb2.t25 421.75
R7610 two_stage_opamp_dummy_magic_14_0.Vb2.n15 two_stage_opamp_dummy_magic_14_0.Vb2.t21 421.75
R7611 two_stage_opamp_dummy_magic_14_0.Vb2.n16 two_stage_opamp_dummy_magic_14_0.Vb2.t30 421.75
R7612 two_stage_opamp_dummy_magic_14_0.Vb2.n9 two_stage_opamp_dummy_magic_14_0.Vb2.t16 421.75
R7613 two_stage_opamp_dummy_magic_14_0.Vb2.n10 two_stage_opamp_dummy_magic_14_0.Vb2.t20 421.75
R7614 two_stage_opamp_dummy_magic_14_0.Vb2.n11 two_stage_opamp_dummy_magic_14_0.Vb2.t15 421.75
R7615 two_stage_opamp_dummy_magic_14_0.Vb2.n12 two_stage_opamp_dummy_magic_14_0.Vb2.t11 421.75
R7616 two_stage_opamp_dummy_magic_14_0.Vb2.n30 two_stage_opamp_dummy_magic_14_0.Vb2.n17 169.352
R7617 two_stage_opamp_dummy_magic_14_0.Vb2.n5 two_stage_opamp_dummy_magic_14_0.Vb2.n4 167.094
R7618 two_stage_opamp_dummy_magic_14_0.Vb2.n6 two_stage_opamp_dummy_magic_14_0.Vb2.n5 167.094
R7619 two_stage_opamp_dummy_magic_14_0.Vb2.n7 two_stage_opamp_dummy_magic_14_0.Vb2.n6 167.094
R7620 two_stage_opamp_dummy_magic_14_0.Vb2.n1 two_stage_opamp_dummy_magic_14_0.Vb2.n0 167.094
R7621 two_stage_opamp_dummy_magic_14_0.Vb2.n2 two_stage_opamp_dummy_magic_14_0.Vb2.n1 167.094
R7622 two_stage_opamp_dummy_magic_14_0.Vb2.n3 two_stage_opamp_dummy_magic_14_0.Vb2.n2 167.094
R7623 two_stage_opamp_dummy_magic_14_0.Vb2.n14 two_stage_opamp_dummy_magic_14_0.Vb2.n13 167.094
R7624 two_stage_opamp_dummy_magic_14_0.Vb2.n15 two_stage_opamp_dummy_magic_14_0.Vb2.n14 167.094
R7625 two_stage_opamp_dummy_magic_14_0.Vb2.n16 two_stage_opamp_dummy_magic_14_0.Vb2.n15 167.094
R7626 two_stage_opamp_dummy_magic_14_0.Vb2.n10 two_stage_opamp_dummy_magic_14_0.Vb2.n9 167.094
R7627 two_stage_opamp_dummy_magic_14_0.Vb2.n11 two_stage_opamp_dummy_magic_14_0.Vb2.n10 167.094
R7628 two_stage_opamp_dummy_magic_14_0.Vb2.n12 two_stage_opamp_dummy_magic_14_0.Vb2.n11 167.094
R7629 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.Vb2.n8 161.477
R7630 two_stage_opamp_dummy_magic_14_0.Vb2.n27 two_stage_opamp_dummy_magic_14_0.Vb2.n26 160.06
R7631 two_stage_opamp_dummy_magic_14_0.Vb2.n20 two_stage_opamp_dummy_magic_14_0.Vb2.n18 140.857
R7632 two_stage_opamp_dummy_magic_14_0.Vb2.n22 two_stage_opamp_dummy_magic_14_0.Vb2.n21 139.608
R7633 two_stage_opamp_dummy_magic_14_0.Vb2.n24 two_stage_opamp_dummy_magic_14_0.Vb2.n23 139.608
R7634 two_stage_opamp_dummy_magic_14_0.Vb2.n20 two_stage_opamp_dummy_magic_14_0.Vb2.n19 139.608
R7635 two_stage_opamp_dummy_magic_14_0.Vb2.n25 two_stage_opamp_dummy_magic_14_0.Vb2.n24 61.3349
R7636 two_stage_opamp_dummy_magic_14_0.Vb2.n8 two_stage_opamp_dummy_magic_14_0.Vb2.n7 49.8072
R7637 two_stage_opamp_dummy_magic_14_0.Vb2.n8 two_stage_opamp_dummy_magic_14_0.Vb2.n3 49.8072
R7638 two_stage_opamp_dummy_magic_14_0.Vb2.n17 two_stage_opamp_dummy_magic_14_0.Vb2.n16 49.8072
R7639 two_stage_opamp_dummy_magic_14_0.Vb2.n17 two_stage_opamp_dummy_magic_14_0.Vb2.n12 49.8072
R7640 two_stage_opamp_dummy_magic_14_0.Vb2.n18 two_stage_opamp_dummy_magic_14_0.Vb2.t6 24.0005
R7641 two_stage_opamp_dummy_magic_14_0.Vb2.n18 two_stage_opamp_dummy_magic_14_0.Vb2.t8 24.0005
R7642 two_stage_opamp_dummy_magic_14_0.Vb2.n21 two_stage_opamp_dummy_magic_14_0.Vb2.t4 24.0005
R7643 two_stage_opamp_dummy_magic_14_0.Vb2.n21 two_stage_opamp_dummy_magic_14_0.Vb2.t2 24.0005
R7644 two_stage_opamp_dummy_magic_14_0.Vb2.n23 two_stage_opamp_dummy_magic_14_0.Vb2.t9 24.0005
R7645 two_stage_opamp_dummy_magic_14_0.Vb2.n23 two_stage_opamp_dummy_magic_14_0.Vb2.t3 24.0005
R7646 two_stage_opamp_dummy_magic_14_0.Vb2.n19 two_stage_opamp_dummy_magic_14_0.Vb2.t5 24.0005
R7647 two_stage_opamp_dummy_magic_14_0.Vb2.n19 two_stage_opamp_dummy_magic_14_0.Vb2.t7 24.0005
R7648 two_stage_opamp_dummy_magic_14_0.Vb2.n30 two_stage_opamp_dummy_magic_14_0.Vb2.n29 12.8443
R7649 two_stage_opamp_dummy_magic_14_0.Vb2.n26 two_stage_opamp_dummy_magic_14_0.Vb2.t1 11.2576
R7650 two_stage_opamp_dummy_magic_14_0.Vb2.n26 two_stage_opamp_dummy_magic_14_0.Vb2.t10 11.2576
R7651 two_stage_opamp_dummy_magic_14_0.Vb2.n22 two_stage_opamp_dummy_magic_14_0.Vb2.n20 7.563
R7652 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.Vb2.n30 7.2505
R7653 two_stage_opamp_dummy_magic_14_0.Vb2.n29 two_stage_opamp_dummy_magic_14_0.Vb2.n25 4.54113
R7654 two_stage_opamp_dummy_magic_14_0.Vb2.n28 two_stage_opamp_dummy_magic_14_0.Vb2.n27 2.84425
R7655 two_stage_opamp_dummy_magic_14_0.Vb2.n24 two_stage_opamp_dummy_magic_14_0.Vb2.n22 1.2505
R7656 two_stage_opamp_dummy_magic_14_0.Vb2.n29 two_stage_opamp_dummy_magic_14_0.Vb2.n28 0.928625
R7657 two_stage_opamp_dummy_magic_14_0.VD3.n23 two_stage_opamp_dummy_magic_14_0.VD3.t25 652.076
R7658 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.t22 652.076
R7659 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n2 585
R7660 two_stage_opamp_dummy_magic_14_0.VD3.n37 two_stage_opamp_dummy_magic_14_0.VD3.n36 585
R7661 two_stage_opamp_dummy_magic_14_0.VD3.n43 two_stage_opamp_dummy_magic_14_0.VD3.n2 290.233
R7662 two_stage_opamp_dummy_magic_14_0.VD3.n49 two_stage_opamp_dummy_magic_14_0.VD3.n2 290.233
R7663 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n2 290.233
R7664 two_stage_opamp_dummy_magic_14_0.VD3.n36 two_stage_opamp_dummy_magic_14_0.VD3.n25 290.233
R7665 two_stage_opamp_dummy_magic_14_0.VD3.n36 two_stage_opamp_dummy_magic_14_0.VD3.n30 290.233
R7666 two_stage_opamp_dummy_magic_14_0.VD3.n36 two_stage_opamp_dummy_magic_14_0.VD3.n35 290.233
R7667 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n41 242.903
R7668 two_stage_opamp_dummy_magic_14_0.VD3.n35 two_stage_opamp_dummy_magic_14_0.VD3.n7 242.903
R7669 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n54 238.367
R7670 two_stage_opamp_dummy_magic_14_0.VD3.n4 two_stage_opamp_dummy_magic_14_0.VD3.n3 185
R7671 two_stage_opamp_dummy_magic_14_0.VD3.n52 two_stage_opamp_dummy_magic_14_0.VD3.n51 185
R7672 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.n52 185
R7673 two_stage_opamp_dummy_magic_14_0.VD3.n50 two_stage_opamp_dummy_magic_14_0.VD3.n42 185
R7674 two_stage_opamp_dummy_magic_14_0.VD3.n48 two_stage_opamp_dummy_magic_14_0.VD3.n47 185
R7675 two_stage_opamp_dummy_magic_14_0.VD3.n46 two_stage_opamp_dummy_magic_14_0.VD3.n45 185
R7676 two_stage_opamp_dummy_magic_14_0.VD3.n38 two_stage_opamp_dummy_magic_14_0.VD3.n37 185
R7677 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n38 185
R7678 two_stage_opamp_dummy_magic_14_0.VD3.n24 two_stage_opamp_dummy_magic_14_0.VD3.n8 185
R7679 two_stage_opamp_dummy_magic_14_0.VD3.n27 two_stage_opamp_dummy_magic_14_0.VD3.n26 185
R7680 two_stage_opamp_dummy_magic_14_0.VD3.n29 two_stage_opamp_dummy_magic_14_0.VD3.n28 185
R7681 two_stage_opamp_dummy_magic_14_0.VD3.n32 two_stage_opamp_dummy_magic_14_0.VD3.n31 185
R7682 two_stage_opamp_dummy_magic_14_0.VD3.n34 two_stage_opamp_dummy_magic_14_0.VD3.n33 185
R7683 two_stage_opamp_dummy_magic_14_0.VD3.t26 two_stage_opamp_dummy_magic_14_0.VD3.n39 170.513
R7684 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.t23 170.513
R7685 two_stage_opamp_dummy_magic_14_0.VD3.n11 two_stage_opamp_dummy_magic_14_0.VD3.n9 163.626
R7686 two_stage_opamp_dummy_magic_14_0.VD3.n19 two_stage_opamp_dummy_magic_14_0.VD3.n18 163.001
R7687 two_stage_opamp_dummy_magic_14_0.VD3.n17 two_stage_opamp_dummy_magic_14_0.VD3.n16 163.001
R7688 two_stage_opamp_dummy_magic_14_0.VD3.n15 two_stage_opamp_dummy_magic_14_0.VD3.n14 163.001
R7689 two_stage_opamp_dummy_magic_14_0.VD3.n13 two_stage_opamp_dummy_magic_14_0.VD3.n12 163.001
R7690 two_stage_opamp_dummy_magic_14_0.VD3.n11 two_stage_opamp_dummy_magic_14_0.VD3.n10 163.001
R7691 two_stage_opamp_dummy_magic_14_0.VD3.n62 two_stage_opamp_dummy_magic_14_0.VD3.n61 159.804
R7692 two_stage_opamp_dummy_magic_14_0.VD3.n1 two_stage_opamp_dummy_magic_14_0.VD3.n0 159.803
R7693 two_stage_opamp_dummy_magic_14_0.VD3.n21 two_stage_opamp_dummy_magic_14_0.VD3.n20 159.803
R7694 two_stage_opamp_dummy_magic_14_0.VD3.n58 two_stage_opamp_dummy_magic_14_0.VD3.n57 159.803
R7695 two_stage_opamp_dummy_magic_14_0.VD3.n60 two_stage_opamp_dummy_magic_14_0.VD3.n59 159.803
R7696 two_stage_opamp_dummy_magic_14_0.VD3.n52 two_stage_opamp_dummy_magic_14_0.VD3.n4 150
R7697 two_stage_opamp_dummy_magic_14_0.VD3.n52 two_stage_opamp_dummy_magic_14_0.VD3.n42 150
R7698 two_stage_opamp_dummy_magic_14_0.VD3.n47 two_stage_opamp_dummy_magic_14_0.VD3.n46 150
R7699 two_stage_opamp_dummy_magic_14_0.VD3.n38 two_stage_opamp_dummy_magic_14_0.VD3.n8 150
R7700 two_stage_opamp_dummy_magic_14_0.VD3.n28 two_stage_opamp_dummy_magic_14_0.VD3.n27 150
R7701 two_stage_opamp_dummy_magic_14_0.VD3.n33 two_stage_opamp_dummy_magic_14_0.VD3.n32 150
R7702 two_stage_opamp_dummy_magic_14_0.VD3.t4 two_stage_opamp_dummy_magic_14_0.VD3.t26 146.155
R7703 two_stage_opamp_dummy_magic_14_0.VD3.t12 two_stage_opamp_dummy_magic_14_0.VD3.t4 146.155
R7704 two_stage_opamp_dummy_magic_14_0.VD3.t8 two_stage_opamp_dummy_magic_14_0.VD3.t12 146.155
R7705 two_stage_opamp_dummy_magic_14_0.VD3.t14 two_stage_opamp_dummy_magic_14_0.VD3.t8 146.155
R7706 two_stage_opamp_dummy_magic_14_0.VD3.t18 two_stage_opamp_dummy_magic_14_0.VD3.t14 146.155
R7707 two_stage_opamp_dummy_magic_14_0.VD3.t0 two_stage_opamp_dummy_magic_14_0.VD3.t18 146.155
R7708 two_stage_opamp_dummy_magic_14_0.VD3.t6 two_stage_opamp_dummy_magic_14_0.VD3.t0 146.155
R7709 two_stage_opamp_dummy_magic_14_0.VD3.t2 two_stage_opamp_dummy_magic_14_0.VD3.t6 146.155
R7710 two_stage_opamp_dummy_magic_14_0.VD3.t10 two_stage_opamp_dummy_magic_14_0.VD3.t2 146.155
R7711 two_stage_opamp_dummy_magic_14_0.VD3.t16 two_stage_opamp_dummy_magic_14_0.VD3.t10 146.155
R7712 two_stage_opamp_dummy_magic_14_0.VD3.t23 two_stage_opamp_dummy_magic_14_0.VD3.t16 146.155
R7713 two_stage_opamp_dummy_magic_14_0.VD3.n54 two_stage_opamp_dummy_magic_14_0.VD3.n53 65.8183
R7714 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.n40 65.8183
R7715 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.n41 65.8183
R7716 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n5 65.8183
R7717 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n6 65.8183
R7718 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n7 65.8183
R7719 two_stage_opamp_dummy_magic_14_0.VD3.n42 two_stage_opamp_dummy_magic_14_0.VD3.n40 53.3664
R7720 two_stage_opamp_dummy_magic_14_0.VD3.n46 two_stage_opamp_dummy_magic_14_0.VD3.n41 53.3664
R7721 two_stage_opamp_dummy_magic_14_0.VD3.n54 two_stage_opamp_dummy_magic_14_0.VD3.n4 53.3664
R7722 two_stage_opamp_dummy_magic_14_0.VD3.n47 two_stage_opamp_dummy_magic_14_0.VD3.n40 53.3664
R7723 two_stage_opamp_dummy_magic_14_0.VD3.n8 two_stage_opamp_dummy_magic_14_0.VD3.n5 53.3664
R7724 two_stage_opamp_dummy_magic_14_0.VD3.n28 two_stage_opamp_dummy_magic_14_0.VD3.n6 53.3664
R7725 two_stage_opamp_dummy_magic_14_0.VD3.n33 two_stage_opamp_dummy_magic_14_0.VD3.n7 53.3664
R7726 two_stage_opamp_dummy_magic_14_0.VD3.n27 two_stage_opamp_dummy_magic_14_0.VD3.n5 53.3664
R7727 two_stage_opamp_dummy_magic_14_0.VD3.n32 two_stage_opamp_dummy_magic_14_0.VD3.n6 53.3664
R7728 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.n55 22.8576
R7729 two_stage_opamp_dummy_magic_14_0.VD3.n37 two_stage_opamp_dummy_magic_14_0.VD3.n23 22.8576
R7730 two_stage_opamp_dummy_magic_14_0.VD3.n58 two_stage_opamp_dummy_magic_14_0.VD3.n56 14.4255
R7731 two_stage_opamp_dummy_magic_14_0.VD3.n22 two_stage_opamp_dummy_magic_14_0.VD3.n19 14.188
R7732 two_stage_opamp_dummy_magic_14_0.VD3.n23 two_stage_opamp_dummy_magic_14_0.VD3.n22 13.8005
R7733 two_stage_opamp_dummy_magic_14_0.VD3.n0 two_stage_opamp_dummy_magic_14_0.VD3.t9 11.2576
R7734 two_stage_opamp_dummy_magic_14_0.VD3.n0 two_stage_opamp_dummy_magic_14_0.VD3.t15 11.2576
R7735 two_stage_opamp_dummy_magic_14_0.VD3.n20 two_stage_opamp_dummy_magic_14_0.VD3.t5 11.2576
R7736 two_stage_opamp_dummy_magic_14_0.VD3.n20 two_stage_opamp_dummy_magic_14_0.VD3.t13 11.2576
R7737 two_stage_opamp_dummy_magic_14_0.VD3.n36 two_stage_opamp_dummy_magic_14_0.VD3.t27 11.2576
R7738 two_stage_opamp_dummy_magic_14_0.VD3.n2 two_stage_opamp_dummy_magic_14_0.VD3.t24 11.2576
R7739 two_stage_opamp_dummy_magic_14_0.VD3.n57 two_stage_opamp_dummy_magic_14_0.VD3.t11 11.2576
R7740 two_stage_opamp_dummy_magic_14_0.VD3.n57 two_stage_opamp_dummy_magic_14_0.VD3.t17 11.2576
R7741 two_stage_opamp_dummy_magic_14_0.VD3.n59 two_stage_opamp_dummy_magic_14_0.VD3.t7 11.2576
R7742 two_stage_opamp_dummy_magic_14_0.VD3.n59 two_stage_opamp_dummy_magic_14_0.VD3.t3 11.2576
R7743 two_stage_opamp_dummy_magic_14_0.VD3.n18 two_stage_opamp_dummy_magic_14_0.VD3.t28 11.2576
R7744 two_stage_opamp_dummy_magic_14_0.VD3.n18 two_stage_opamp_dummy_magic_14_0.VD3.t20 11.2576
R7745 two_stage_opamp_dummy_magic_14_0.VD3.n16 two_stage_opamp_dummy_magic_14_0.VD3.t35 11.2576
R7746 two_stage_opamp_dummy_magic_14_0.VD3.n16 two_stage_opamp_dummy_magic_14_0.VD3.t30 11.2576
R7747 two_stage_opamp_dummy_magic_14_0.VD3.n14 two_stage_opamp_dummy_magic_14_0.VD3.t33 11.2576
R7748 two_stage_opamp_dummy_magic_14_0.VD3.n14 two_stage_opamp_dummy_magic_14_0.VD3.t34 11.2576
R7749 two_stage_opamp_dummy_magic_14_0.VD3.n12 two_stage_opamp_dummy_magic_14_0.VD3.t32 11.2576
R7750 two_stage_opamp_dummy_magic_14_0.VD3.n12 two_stage_opamp_dummy_magic_14_0.VD3.t31 11.2576
R7751 two_stage_opamp_dummy_magic_14_0.VD3.n10 two_stage_opamp_dummy_magic_14_0.VD3.t37 11.2576
R7752 two_stage_opamp_dummy_magic_14_0.VD3.n10 two_stage_opamp_dummy_magic_14_0.VD3.t29 11.2576
R7753 two_stage_opamp_dummy_magic_14_0.VD3.n9 two_stage_opamp_dummy_magic_14_0.VD3.t21 11.2576
R7754 two_stage_opamp_dummy_magic_14_0.VD3.n9 two_stage_opamp_dummy_magic_14_0.VD3.t36 11.2576
R7755 two_stage_opamp_dummy_magic_14_0.VD3.t19 two_stage_opamp_dummy_magic_14_0.VD3.n62 11.2576
R7756 two_stage_opamp_dummy_magic_14_0.VD3.n62 two_stage_opamp_dummy_magic_14_0.VD3.t1 11.2576
R7757 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n3 9.14336
R7758 two_stage_opamp_dummy_magic_14_0.VD3.n51 two_stage_opamp_dummy_magic_14_0.VD3.n50 9.14336
R7759 two_stage_opamp_dummy_magic_14_0.VD3.n48 two_stage_opamp_dummy_magic_14_0.VD3.n45 9.14336
R7760 two_stage_opamp_dummy_magic_14_0.VD3.n37 two_stage_opamp_dummy_magic_14_0.VD3.n24 9.14336
R7761 two_stage_opamp_dummy_magic_14_0.VD3.n29 two_stage_opamp_dummy_magic_14_0.VD3.n26 9.14336
R7762 two_stage_opamp_dummy_magic_14_0.VD3.n34 two_stage_opamp_dummy_magic_14_0.VD3.n31 9.14336
R7763 two_stage_opamp_dummy_magic_14_0.VD3.n43 two_stage_opamp_dummy_magic_14_0.VD3.n3 4.53698
R7764 two_stage_opamp_dummy_magic_14_0.VD3.n50 two_stage_opamp_dummy_magic_14_0.VD3.n49 4.53698
R7765 two_stage_opamp_dummy_magic_14_0.VD3.n45 two_stage_opamp_dummy_magic_14_0.VD3.n44 4.53698
R7766 two_stage_opamp_dummy_magic_14_0.VD3.n51 two_stage_opamp_dummy_magic_14_0.VD3.n43 4.53698
R7767 two_stage_opamp_dummy_magic_14_0.VD3.n49 two_stage_opamp_dummy_magic_14_0.VD3.n48 4.53698
R7768 two_stage_opamp_dummy_magic_14_0.VD3.n25 two_stage_opamp_dummy_magic_14_0.VD3.n24 4.53698
R7769 two_stage_opamp_dummy_magic_14_0.VD3.n30 two_stage_opamp_dummy_magic_14_0.VD3.n29 4.53698
R7770 two_stage_opamp_dummy_magic_14_0.VD3.n35 two_stage_opamp_dummy_magic_14_0.VD3.n34 4.53698
R7771 two_stage_opamp_dummy_magic_14_0.VD3.n26 two_stage_opamp_dummy_magic_14_0.VD3.n25 4.53698
R7772 two_stage_opamp_dummy_magic_14_0.VD3.n31 two_stage_opamp_dummy_magic_14_0.VD3.n30 4.53698
R7773 two_stage_opamp_dummy_magic_14_0.VD3.n61 two_stage_opamp_dummy_magic_14_0.VD3.n60 0.6255
R7774 two_stage_opamp_dummy_magic_14_0.VD3.n60 two_stage_opamp_dummy_magic_14_0.VD3.n58 0.6255
R7775 two_stage_opamp_dummy_magic_14_0.VD3.n13 two_stage_opamp_dummy_magic_14_0.VD3.n11 0.6255
R7776 two_stage_opamp_dummy_magic_14_0.VD3.n15 two_stage_opamp_dummy_magic_14_0.VD3.n13 0.6255
R7777 two_stage_opamp_dummy_magic_14_0.VD3.n17 two_stage_opamp_dummy_magic_14_0.VD3.n15 0.6255
R7778 two_stage_opamp_dummy_magic_14_0.VD3.n19 two_stage_opamp_dummy_magic_14_0.VD3.n17 0.6255
R7779 two_stage_opamp_dummy_magic_14_0.VD3.n22 two_stage_opamp_dummy_magic_14_0.VD3.n21 0.6255
R7780 two_stage_opamp_dummy_magic_14_0.VD3.n21 two_stage_opamp_dummy_magic_14_0.VD3.n1 0.6255
R7781 two_stage_opamp_dummy_magic_14_0.VD3.n61 two_stage_opamp_dummy_magic_14_0.VD3.n1 0.6255
R7782 two_stage_opamp_dummy_magic_14_0.Y.n47 two_stage_opamp_dummy_magic_14_0.Y.t30 1172.87
R7783 two_stage_opamp_dummy_magic_14_0.Y.n43 two_stage_opamp_dummy_magic_14_0.Y.t36 1172.87
R7784 two_stage_opamp_dummy_magic_14_0.Y.n50 two_stage_opamp_dummy_magic_14_0.Y.t54 996.134
R7785 two_stage_opamp_dummy_magic_14_0.Y.n49 two_stage_opamp_dummy_magic_14_0.Y.t40 996.134
R7786 two_stage_opamp_dummy_magic_14_0.Y.n48 two_stage_opamp_dummy_magic_14_0.Y.t26 996.134
R7787 two_stage_opamp_dummy_magic_14_0.Y.n47 two_stage_opamp_dummy_magic_14_0.Y.t43 996.134
R7788 two_stage_opamp_dummy_magic_14_0.Y.n43 two_stage_opamp_dummy_magic_14_0.Y.t52 996.134
R7789 two_stage_opamp_dummy_magic_14_0.Y.n44 two_stage_opamp_dummy_magic_14_0.Y.t46 996.134
R7790 two_stage_opamp_dummy_magic_14_0.Y.n45 two_stage_opamp_dummy_magic_14_0.Y.t51 996.134
R7791 two_stage_opamp_dummy_magic_14_0.Y.n46 two_stage_opamp_dummy_magic_14_0.Y.t37 996.134
R7792 two_stage_opamp_dummy_magic_14_0.Y.n35 two_stage_opamp_dummy_magic_14_0.Y.t35 690.867
R7793 two_stage_opamp_dummy_magic_14_0.Y.n32 two_stage_opamp_dummy_magic_14_0.Y.t41 690.867
R7794 two_stage_opamp_dummy_magic_14_0.Y.n26 two_stage_opamp_dummy_magic_14_0.Y.t48 530.201
R7795 two_stage_opamp_dummy_magic_14_0.Y.n23 two_stage_opamp_dummy_magic_14_0.Y.t53 530.201
R7796 two_stage_opamp_dummy_magic_14_0.Y.n35 two_stage_opamp_dummy_magic_14_0.Y.t49 514.134
R7797 two_stage_opamp_dummy_magic_14_0.Y.n36 two_stage_opamp_dummy_magic_14_0.Y.t33 514.134
R7798 two_stage_opamp_dummy_magic_14_0.Y.n37 two_stage_opamp_dummy_magic_14_0.Y.t47 514.134
R7799 two_stage_opamp_dummy_magic_14_0.Y.n38 two_stage_opamp_dummy_magic_14_0.Y.t31 514.134
R7800 two_stage_opamp_dummy_magic_14_0.Y.n39 two_stage_opamp_dummy_magic_14_0.Y.t44 514.134
R7801 two_stage_opamp_dummy_magic_14_0.Y.n34 two_stage_opamp_dummy_magic_14_0.Y.t27 514.134
R7802 two_stage_opamp_dummy_magic_14_0.Y.n33 two_stage_opamp_dummy_magic_14_0.Y.t50 514.134
R7803 two_stage_opamp_dummy_magic_14_0.Y.n32 two_stage_opamp_dummy_magic_14_0.Y.t28 514.134
R7804 two_stage_opamp_dummy_magic_14_0.Y.n30 two_stage_opamp_dummy_magic_14_0.Y.t25 353.467
R7805 two_stage_opamp_dummy_magic_14_0.Y.n29 two_stage_opamp_dummy_magic_14_0.Y.t42 353.467
R7806 two_stage_opamp_dummy_magic_14_0.Y.n28 two_stage_opamp_dummy_magic_14_0.Y.t29 353.467
R7807 two_stage_opamp_dummy_magic_14_0.Y.n27 two_stage_opamp_dummy_magic_14_0.Y.t45 353.467
R7808 two_stage_opamp_dummy_magic_14_0.Y.n26 two_stage_opamp_dummy_magic_14_0.Y.t32 353.467
R7809 two_stage_opamp_dummy_magic_14_0.Y.n23 two_stage_opamp_dummy_magic_14_0.Y.t39 353.467
R7810 two_stage_opamp_dummy_magic_14_0.Y.n24 two_stage_opamp_dummy_magic_14_0.Y.t34 353.467
R7811 two_stage_opamp_dummy_magic_14_0.Y.n25 two_stage_opamp_dummy_magic_14_0.Y.t38 353.467
R7812 two_stage_opamp_dummy_magic_14_0.Y.n50 two_stage_opamp_dummy_magic_14_0.Y.n49 176.733
R7813 two_stage_opamp_dummy_magic_14_0.Y.n49 two_stage_opamp_dummy_magic_14_0.Y.n48 176.733
R7814 two_stage_opamp_dummy_magic_14_0.Y.n48 two_stage_opamp_dummy_magic_14_0.Y.n47 176.733
R7815 two_stage_opamp_dummy_magic_14_0.Y.n44 two_stage_opamp_dummy_magic_14_0.Y.n43 176.733
R7816 two_stage_opamp_dummy_magic_14_0.Y.n45 two_stage_opamp_dummy_magic_14_0.Y.n44 176.733
R7817 two_stage_opamp_dummy_magic_14_0.Y.n46 two_stage_opamp_dummy_magic_14_0.Y.n45 176.733
R7818 two_stage_opamp_dummy_magic_14_0.Y.n30 two_stage_opamp_dummy_magic_14_0.Y.n29 176.733
R7819 two_stage_opamp_dummy_magic_14_0.Y.n29 two_stage_opamp_dummy_magic_14_0.Y.n28 176.733
R7820 two_stage_opamp_dummy_magic_14_0.Y.n28 two_stage_opamp_dummy_magic_14_0.Y.n27 176.733
R7821 two_stage_opamp_dummy_magic_14_0.Y.n27 two_stage_opamp_dummy_magic_14_0.Y.n26 176.733
R7822 two_stage_opamp_dummy_magic_14_0.Y.n24 two_stage_opamp_dummy_magic_14_0.Y.n23 176.733
R7823 two_stage_opamp_dummy_magic_14_0.Y.n25 two_stage_opamp_dummy_magic_14_0.Y.n24 176.733
R7824 two_stage_opamp_dummy_magic_14_0.Y.n39 two_stage_opamp_dummy_magic_14_0.Y.n38 176.733
R7825 two_stage_opamp_dummy_magic_14_0.Y.n38 two_stage_opamp_dummy_magic_14_0.Y.n37 176.733
R7826 two_stage_opamp_dummy_magic_14_0.Y.n37 two_stage_opamp_dummy_magic_14_0.Y.n36 176.733
R7827 two_stage_opamp_dummy_magic_14_0.Y.n36 two_stage_opamp_dummy_magic_14_0.Y.n35 176.733
R7828 two_stage_opamp_dummy_magic_14_0.Y.n33 two_stage_opamp_dummy_magic_14_0.Y.n32 176.733
R7829 two_stage_opamp_dummy_magic_14_0.Y.n34 two_stage_opamp_dummy_magic_14_0.Y.n33 176.733
R7830 two_stage_opamp_dummy_magic_14_0.Y.n52 two_stage_opamp_dummy_magic_14_0.Y.n51 166.258
R7831 two_stage_opamp_dummy_magic_14_0.Y.n2 two_stage_opamp_dummy_magic_14_0.Y.n0 163.626
R7832 two_stage_opamp_dummy_magic_14_0.Y.n8 two_stage_opamp_dummy_magic_14_0.Y.n7 163.001
R7833 two_stage_opamp_dummy_magic_14_0.Y.n6 two_stage_opamp_dummy_magic_14_0.Y.n5 163.001
R7834 two_stage_opamp_dummy_magic_14_0.Y.n4 two_stage_opamp_dummy_magic_14_0.Y.n3 163.001
R7835 two_stage_opamp_dummy_magic_14_0.Y.n2 two_stage_opamp_dummy_magic_14_0.Y.n1 163.001
R7836 two_stage_opamp_dummy_magic_14_0.Y.n41 two_stage_opamp_dummy_magic_14_0.Y.n31 161.541
R7837 two_stage_opamp_dummy_magic_14_0.Y.n41 two_stage_opamp_dummy_magic_14_0.Y.n40 161.541
R7838 two_stage_opamp_dummy_magic_14_0.Y.n10 two_stage_opamp_dummy_magic_14_0.Y.n9 158.501
R7839 two_stage_opamp_dummy_magic_14_0.Y.n13 two_stage_opamp_dummy_magic_14_0.Y.n11 117.888
R7840 two_stage_opamp_dummy_magic_14_0.Y.n21 two_stage_opamp_dummy_magic_14_0.Y.n20 117.326
R7841 two_stage_opamp_dummy_magic_14_0.Y.n19 two_stage_opamp_dummy_magic_14_0.Y.n18 117.326
R7842 two_stage_opamp_dummy_magic_14_0.Y.n17 two_stage_opamp_dummy_magic_14_0.Y.n16 117.326
R7843 two_stage_opamp_dummy_magic_14_0.Y.n15 two_stage_opamp_dummy_magic_14_0.Y.n14 117.326
R7844 two_stage_opamp_dummy_magic_14_0.Y.n13 two_stage_opamp_dummy_magic_14_0.Y.n12 117.326
R7845 two_stage_opamp_dummy_magic_14_0.Y.n31 two_stage_opamp_dummy_magic_14_0.Y.n30 54.6272
R7846 two_stage_opamp_dummy_magic_14_0.Y.n31 two_stage_opamp_dummy_magic_14_0.Y.n25 54.6272
R7847 two_stage_opamp_dummy_magic_14_0.Y.n40 two_stage_opamp_dummy_magic_14_0.Y.n39 54.6272
R7848 two_stage_opamp_dummy_magic_14_0.Y.n40 two_stage_opamp_dummy_magic_14_0.Y.n34 54.6272
R7849 two_stage_opamp_dummy_magic_14_0.Y.n51 two_stage_opamp_dummy_magic_14_0.Y.n50 53.3126
R7850 two_stage_opamp_dummy_magic_14_0.Y.n51 two_stage_opamp_dummy_magic_14_0.Y.n46 53.3126
R7851 two_stage_opamp_dummy_magic_14_0.Y.t16 two_stage_opamp_dummy_magic_14_0.Y.n52 49.8031
R7852 two_stage_opamp_dummy_magic_14_0.Y.n20 two_stage_opamp_dummy_magic_14_0.Y.t17 16.0005
R7853 two_stage_opamp_dummy_magic_14_0.Y.n20 two_stage_opamp_dummy_magic_14_0.Y.t22 16.0005
R7854 two_stage_opamp_dummy_magic_14_0.Y.n18 two_stage_opamp_dummy_magic_14_0.Y.t13 16.0005
R7855 two_stage_opamp_dummy_magic_14_0.Y.n18 two_stage_opamp_dummy_magic_14_0.Y.t21 16.0005
R7856 two_stage_opamp_dummy_magic_14_0.Y.n16 two_stage_opamp_dummy_magic_14_0.Y.t15 16.0005
R7857 two_stage_opamp_dummy_magic_14_0.Y.n16 two_stage_opamp_dummy_magic_14_0.Y.t18 16.0005
R7858 two_stage_opamp_dummy_magic_14_0.Y.n14 two_stage_opamp_dummy_magic_14_0.Y.t12 16.0005
R7859 two_stage_opamp_dummy_magic_14_0.Y.n14 two_stage_opamp_dummy_magic_14_0.Y.t19 16.0005
R7860 two_stage_opamp_dummy_magic_14_0.Y.n12 two_stage_opamp_dummy_magic_14_0.Y.t14 16.0005
R7861 two_stage_opamp_dummy_magic_14_0.Y.n12 two_stage_opamp_dummy_magic_14_0.Y.t11 16.0005
R7862 two_stage_opamp_dummy_magic_14_0.Y.n11 two_stage_opamp_dummy_magic_14_0.Y.t23 16.0005
R7863 two_stage_opamp_dummy_magic_14_0.Y.n11 two_stage_opamp_dummy_magic_14_0.Y.t24 16.0005
R7864 two_stage_opamp_dummy_magic_14_0.Y.n22 two_stage_opamp_dummy_magic_14_0.Y.n10 15.8443
R7865 two_stage_opamp_dummy_magic_14_0.Y.n42 two_stage_opamp_dummy_magic_14_0.Y.n41 13.4693
R7866 two_stage_opamp_dummy_magic_14_0.Y.n9 two_stage_opamp_dummy_magic_14_0.Y.t2 11.2576
R7867 two_stage_opamp_dummy_magic_14_0.Y.n9 two_stage_opamp_dummy_magic_14_0.Y.t20 11.2576
R7868 two_stage_opamp_dummy_magic_14_0.Y.n7 two_stage_opamp_dummy_magic_14_0.Y.t0 11.2576
R7869 two_stage_opamp_dummy_magic_14_0.Y.n7 two_stage_opamp_dummy_magic_14_0.Y.t5 11.2576
R7870 two_stage_opamp_dummy_magic_14_0.Y.n5 two_stage_opamp_dummy_magic_14_0.Y.t9 11.2576
R7871 two_stage_opamp_dummy_magic_14_0.Y.n5 two_stage_opamp_dummy_magic_14_0.Y.t3 11.2576
R7872 two_stage_opamp_dummy_magic_14_0.Y.n3 two_stage_opamp_dummy_magic_14_0.Y.t1 11.2576
R7873 two_stage_opamp_dummy_magic_14_0.Y.n3 two_stage_opamp_dummy_magic_14_0.Y.t4 11.2576
R7874 two_stage_opamp_dummy_magic_14_0.Y.n1 two_stage_opamp_dummy_magic_14_0.Y.t8 11.2576
R7875 two_stage_opamp_dummy_magic_14_0.Y.n1 two_stage_opamp_dummy_magic_14_0.Y.t6 11.2576
R7876 two_stage_opamp_dummy_magic_14_0.Y.n0 two_stage_opamp_dummy_magic_14_0.Y.t10 11.2576
R7877 two_stage_opamp_dummy_magic_14_0.Y.n0 two_stage_opamp_dummy_magic_14_0.Y.t7 11.2576
R7878 two_stage_opamp_dummy_magic_14_0.Y.n52 two_stage_opamp_dummy_magic_14_0.Y.n42 7.09425
R7879 two_stage_opamp_dummy_magic_14_0.Y.n22 two_stage_opamp_dummy_magic_14_0.Y.n21 6.3755
R7880 two_stage_opamp_dummy_magic_14_0.Y.n10 two_stage_opamp_dummy_magic_14_0.Y.n8 5.1255
R7881 two_stage_opamp_dummy_magic_14_0.Y.n42 two_stage_opamp_dummy_magic_14_0.Y.n22 1.40675
R7882 two_stage_opamp_dummy_magic_14_0.Y.n4 two_stage_opamp_dummy_magic_14_0.Y.n2 0.6255
R7883 two_stage_opamp_dummy_magic_14_0.Y.n6 two_stage_opamp_dummy_magic_14_0.Y.n4 0.6255
R7884 two_stage_opamp_dummy_magic_14_0.Y.n8 two_stage_opamp_dummy_magic_14_0.Y.n6 0.6255
R7885 two_stage_opamp_dummy_magic_14_0.Y.n15 two_stage_opamp_dummy_magic_14_0.Y.n13 0.563
R7886 two_stage_opamp_dummy_magic_14_0.Y.n17 two_stage_opamp_dummy_magic_14_0.Y.n15 0.563
R7887 two_stage_opamp_dummy_magic_14_0.Y.n19 two_stage_opamp_dummy_magic_14_0.Y.n17 0.563
R7888 two_stage_opamp_dummy_magic_14_0.Y.n21 two_stage_opamp_dummy_magic_14_0.Y.n19 0.563
R7889 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 345.264
R7890 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 344.7
R7891 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 292.5
R7892 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 209.251
R7893 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 208.689
R7894 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 208.689
R7895 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 208.689
R7896 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 208.689
R7897 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 120.305
R7898 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 52.763
R7899 bgr_7_0.V_CMFB_S3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 51.7297
R7900 bgr_7_0.V_CMFB_S3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 41.2477
R7901 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 39.4005
R7902 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 39.4005
R7903 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 39.4005
R7904 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 39.4005
R7905 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 39.4005
R7906 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 39.4005
R7907 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 19.7005
R7908 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 19.7005
R7909 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 19.7005
R7910 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 19.7005
R7911 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 19.7005
R7912 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 19.7005
R7913 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 19.7005
R7914 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 19.7005
R7915 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 19.7005
R7916 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 19.7005
R7917 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 5.90675
R7918 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 0.563
R7919 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 0.563
R7920 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 0.563
R7921 bgr_7_0.V_CUR_REF_REG.n4 bgr_7_0.V_CUR_REF_REG.n3 526.183
R7922 bgr_7_0.V_CUR_REF_REG.n2 bgr_7_0.V_CUR_REF_REG.n1 514.134
R7923 bgr_7_0.V_CUR_REF_REG.n5 bgr_7_0.V_CUR_REF_REG.n0 378.053
R7924 bgr_7_0.V_CUR_REF_REG.n1 bgr_7_0.V_CUR_REF_REG.t5 303.259
R7925 bgr_7_0.V_CUR_REF_REG.n5 bgr_7_0.V_CUR_REF_REG.n4 210.169
R7926 bgr_7_0.V_CUR_REF_REG.n1 bgr_7_0.V_CUR_REF_REG.t3 174.726
R7927 bgr_7_0.V_CUR_REF_REG.n2 bgr_7_0.V_CUR_REF_REG.t7 174.726
R7928 bgr_7_0.V_CUR_REF_REG.n3 bgr_7_0.V_CUR_REF_REG.t4 174.726
R7929 bgr_7_0.V_CUR_REF_REG.t0 bgr_7_0.V_CUR_REF_REG.n5 153.474
R7930 bgr_7_0.V_CUR_REF_REG.n3 bgr_7_0.V_CUR_REF_REG.n2 128.534
R7931 bgr_7_0.V_CUR_REF_REG.n4 bgr_7_0.V_CUR_REF_REG.t6 96.4005
R7932 bgr_7_0.V_CUR_REF_REG.n0 bgr_7_0.V_CUR_REF_REG.t2 39.4005
R7933 bgr_7_0.V_CUR_REF_REG.n0 bgr_7_0.V_CUR_REF_REG.t1 39.4005
R7934 bgr_7_0.V_p_2.n1 bgr_7_0.V_p_2.n2 229.562
R7935 bgr_7_0.V_p_2.n1 bgr_7_0.V_p_2.n5 228.939
R7936 bgr_7_0.V_p_2.n0 bgr_7_0.V_p_2.n4 228.939
R7937 bgr_7_0.V_p_2.n0 bgr_7_0.V_p_2.n3 228.939
R7938 bgr_7_0.V_p_2.n6 bgr_7_0.V_p_2.n1 228.938
R7939 bgr_7_0.V_p_2.n0 bgr_7_0.V_p_2.t5 98.7279
R7940 bgr_7_0.V_p_2.n5 bgr_7_0.V_p_2.t8 48.0005
R7941 bgr_7_0.V_p_2.n5 bgr_7_0.V_p_2.t0 48.0005
R7942 bgr_7_0.V_p_2.n4 bgr_7_0.V_p_2.t3 48.0005
R7943 bgr_7_0.V_p_2.n4 bgr_7_0.V_p_2.t10 48.0005
R7944 bgr_7_0.V_p_2.n3 bgr_7_0.V_p_2.t6 48.0005
R7945 bgr_7_0.V_p_2.n3 bgr_7_0.V_p_2.t1 48.0005
R7946 bgr_7_0.V_p_2.n2 bgr_7_0.V_p_2.t9 48.0005
R7947 bgr_7_0.V_p_2.n2 bgr_7_0.V_p_2.t2 48.0005
R7948 bgr_7_0.V_p_2.t4 bgr_7_0.V_p_2.n6 48.0005
R7949 bgr_7_0.V_p_2.n6 bgr_7_0.V_p_2.t7 48.0005
R7950 bgr_7_0.V_p_2.n1 bgr_7_0.V_p_2.n0 1.8755
R7951 a_7460_23988.t0 a_7460_23988.t1 178.133
R7952 two_stage_opamp_dummy_magic_14_0.VD2.n13 two_stage_opamp_dummy_magic_14_0.VD2.n11 146.47
R7953 two_stage_opamp_dummy_magic_14_0.VD2.n17 two_stage_opamp_dummy_magic_14_0.VD2.n15 146.469
R7954 two_stage_opamp_dummy_magic_14_0.VD2.n17 two_stage_opamp_dummy_magic_14_0.VD2.n16 145.906
R7955 two_stage_opamp_dummy_magic_14_0.VD2.n1 two_stage_opamp_dummy_magic_14_0.VD2.n18 145.906
R7956 two_stage_opamp_dummy_magic_14_0.VD2.n0 two_stage_opamp_dummy_magic_14_0.VD2.n14 145.906
R7957 two_stage_opamp_dummy_magic_14_0.VD2.n13 two_stage_opamp_dummy_magic_14_0.VD2.n12 145.906
R7958 two_stage_opamp_dummy_magic_14_0.VD2.n7 two_stage_opamp_dummy_magic_14_0.VD2.n5 114.469
R7959 two_stage_opamp_dummy_magic_14_0.VD2.n4 two_stage_opamp_dummy_magic_14_0.VD2.n2 114.469
R7960 two_stage_opamp_dummy_magic_14_0.VD2.n7 two_stage_opamp_dummy_magic_14_0.VD2.n6 113.906
R7961 two_stage_opamp_dummy_magic_14_0.VD2.n4 two_stage_opamp_dummy_magic_14_0.VD2.n3 113.906
R7962 two_stage_opamp_dummy_magic_14_0.VD2.n10 two_stage_opamp_dummy_magic_14_0.VD2.n9 109.406
R7963 two_stage_opamp_dummy_magic_14_0.VD2.n16 two_stage_opamp_dummy_magic_14_0.VD2.t0 16.0005
R7964 two_stage_opamp_dummy_magic_14_0.VD2.n16 two_stage_opamp_dummy_magic_14_0.VD2.t12 16.0005
R7965 two_stage_opamp_dummy_magic_14_0.VD2.n18 two_stage_opamp_dummy_magic_14_0.VD2.t20 16.0005
R7966 two_stage_opamp_dummy_magic_14_0.VD2.n18 two_stage_opamp_dummy_magic_14_0.VD2.t3 16.0005
R7967 two_stage_opamp_dummy_magic_14_0.VD2.n9 two_stage_opamp_dummy_magic_14_0.VD2.t13 16.0005
R7968 two_stage_opamp_dummy_magic_14_0.VD2.n9 two_stage_opamp_dummy_magic_14_0.VD2.t9 16.0005
R7969 two_stage_opamp_dummy_magic_14_0.VD2.n6 two_stage_opamp_dummy_magic_14_0.VD2.t11 16.0005
R7970 two_stage_opamp_dummy_magic_14_0.VD2.n6 two_stage_opamp_dummy_magic_14_0.VD2.t5 16.0005
R7971 two_stage_opamp_dummy_magic_14_0.VD2.n5 two_stage_opamp_dummy_magic_14_0.VD2.t14 16.0005
R7972 two_stage_opamp_dummy_magic_14_0.VD2.n5 two_stage_opamp_dummy_magic_14_0.VD2.t10 16.0005
R7973 two_stage_opamp_dummy_magic_14_0.VD2.n3 two_stage_opamp_dummy_magic_14_0.VD2.t1 16.0005
R7974 two_stage_opamp_dummy_magic_14_0.VD2.n3 two_stage_opamp_dummy_magic_14_0.VD2.t4 16.0005
R7975 two_stage_opamp_dummy_magic_14_0.VD2.n2 two_stage_opamp_dummy_magic_14_0.VD2.t17 16.0005
R7976 two_stage_opamp_dummy_magic_14_0.VD2.n2 two_stage_opamp_dummy_magic_14_0.VD2.t8 16.0005
R7977 two_stage_opamp_dummy_magic_14_0.VD2.n14 two_stage_opamp_dummy_magic_14_0.VD2.t18 16.0005
R7978 two_stage_opamp_dummy_magic_14_0.VD2.n14 two_stage_opamp_dummy_magic_14_0.VD2.t2 16.0005
R7979 two_stage_opamp_dummy_magic_14_0.VD2.n12 two_stage_opamp_dummy_magic_14_0.VD2.t21 16.0005
R7980 two_stage_opamp_dummy_magic_14_0.VD2.n12 two_stage_opamp_dummy_magic_14_0.VD2.t19 16.0005
R7981 two_stage_opamp_dummy_magic_14_0.VD2.n11 two_stage_opamp_dummy_magic_14_0.VD2.t15 16.0005
R7982 two_stage_opamp_dummy_magic_14_0.VD2.n11 two_stage_opamp_dummy_magic_14_0.VD2.t6 16.0005
R7983 two_stage_opamp_dummy_magic_14_0.VD2.n15 two_stage_opamp_dummy_magic_14_0.VD2.t7 16.0005
R7984 two_stage_opamp_dummy_magic_14_0.VD2.n15 two_stage_opamp_dummy_magic_14_0.VD2.t16 16.0005
R7985 two_stage_opamp_dummy_magic_14_0.VD2 two_stage_opamp_dummy_magic_14_0.VD2.n1 4.64633
R7986 two_stage_opamp_dummy_magic_14_0.VD2.n10 two_stage_opamp_dummy_magic_14_0.VD2.n8 4.5005
R7987 two_stage_opamp_dummy_magic_14_0.VD2.n8 two_stage_opamp_dummy_magic_14_0.VD2.n7 0.563
R7988 two_stage_opamp_dummy_magic_14_0.VD2.n8 two_stage_opamp_dummy_magic_14_0.VD2.n4 0.563
R7989 two_stage_opamp_dummy_magic_14_0.VD2.n0 two_stage_opamp_dummy_magic_14_0.VD2.n13 0.563
R7990 two_stage_opamp_dummy_magic_14_0.VD2.n1 two_stage_opamp_dummy_magic_14_0.VD2.n17 0.563
R7991 two_stage_opamp_dummy_magic_14_0.VD2 two_stage_opamp_dummy_magic_14_0.VD2.n10 0.46925
R7992 two_stage_opamp_dummy_magic_14_0.VD2.n1 two_stage_opamp_dummy_magic_14_0.VD2.n0 0.46925
R7993 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 479.322
R7994 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 479.322
R7995 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 479.322
R7996 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 479.322
R7997 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 178.625
R7998 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 177.987
R7999 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 175.013
R8000 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 165.8
R8001 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 165.8
R8002 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 24.0005
R8003 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 24.0005
R8004 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 15.7605
R8005 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 15.7605
R8006 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 15.7605
R8007 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 15.7605
R8008 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 1.76612
R8009 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 0.641125
R8010 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 187.315
R8011 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 177.755
R8012 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t0 15.7605
R8013 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t1 15.7605
R8014 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t2 15.7605
R8015 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t3 15.7605
R8016 two_stage_opamp_dummy_magic_14_0.Vb1.n14 two_stage_opamp_dummy_magic_14_0.Vb1.t20 449.868
R8017 two_stage_opamp_dummy_magic_14_0.Vb1.n10 two_stage_opamp_dummy_magic_14_0.Vb1.t26 449.868
R8018 two_stage_opamp_dummy_magic_14_0.Vb1.n5 two_stage_opamp_dummy_magic_14_0.Vb1.t12 449.868
R8019 two_stage_opamp_dummy_magic_14_0.Vb1.n1 two_stage_opamp_dummy_magic_14_0.Vb1.t18 449.868
R8020 two_stage_opamp_dummy_magic_14_0.Vb1.n23 two_stage_opamp_dummy_magic_14_0.Vb1.t7 449.868
R8021 two_stage_opamp_dummy_magic_14_0.Vb1.n22 two_stage_opamp_dummy_magic_14_0.Vb1.t5 449.868
R8022 two_stage_opamp_dummy_magic_14_0.Vb1.n14 two_stage_opamp_dummy_magic_14_0.Vb1.t29 273.134
R8023 two_stage_opamp_dummy_magic_14_0.Vb1.n15 two_stage_opamp_dummy_magic_14_0.Vb1.t14 273.134
R8024 two_stage_opamp_dummy_magic_14_0.Vb1.n16 two_stage_opamp_dummy_magic_14_0.Vb1.t25 273.134
R8025 two_stage_opamp_dummy_magic_14_0.Vb1.n17 two_stage_opamp_dummy_magic_14_0.Vb1.t32 273.134
R8026 two_stage_opamp_dummy_magic_14_0.Vb1.n13 two_stage_opamp_dummy_magic_14_0.Vb1.t22 273.134
R8027 two_stage_opamp_dummy_magic_14_0.Vb1.n12 two_stage_opamp_dummy_magic_14_0.Vb1.t17 273.134
R8028 two_stage_opamp_dummy_magic_14_0.Vb1.n11 two_stage_opamp_dummy_magic_14_0.Vb1.t27 273.134
R8029 two_stage_opamp_dummy_magic_14_0.Vb1.n10 two_stage_opamp_dummy_magic_14_0.Vb1.t16 273.134
R8030 two_stage_opamp_dummy_magic_14_0.Vb1.n5 two_stage_opamp_dummy_magic_14_0.Vb1.t23 273.134
R8031 two_stage_opamp_dummy_magic_14_0.Vb1.n6 two_stage_opamp_dummy_magic_14_0.Vb1.t13 273.134
R8032 two_stage_opamp_dummy_magic_14_0.Vb1.n7 two_stage_opamp_dummy_magic_14_0.Vb1.t24 273.134
R8033 two_stage_opamp_dummy_magic_14_0.Vb1.n8 two_stage_opamp_dummy_magic_14_0.Vb1.t31 273.134
R8034 two_stage_opamp_dummy_magic_14_0.Vb1.n4 two_stage_opamp_dummy_magic_14_0.Vb1.t21 273.134
R8035 two_stage_opamp_dummy_magic_14_0.Vb1.n3 two_stage_opamp_dummy_magic_14_0.Vb1.t30 273.134
R8036 two_stage_opamp_dummy_magic_14_0.Vb1.n2 two_stage_opamp_dummy_magic_14_0.Vb1.t19 273.134
R8037 two_stage_opamp_dummy_magic_14_0.Vb1.n1 two_stage_opamp_dummy_magic_14_0.Vb1.t28 273.134
R8038 two_stage_opamp_dummy_magic_14_0.Vb1.n23 two_stage_opamp_dummy_magic_14_0.Vb1.t3 273.134
R8039 two_stage_opamp_dummy_magic_14_0.Vb1.n22 two_stage_opamp_dummy_magic_14_0.Vb1.t1 273.134
R8040 bgr_7_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb1.n0 217.895
R8041 two_stage_opamp_dummy_magic_14_0.Vb1.n17 two_stage_opamp_dummy_magic_14_0.Vb1.n16 176.733
R8042 two_stage_opamp_dummy_magic_14_0.Vb1.n16 two_stage_opamp_dummy_magic_14_0.Vb1.n15 176.733
R8043 two_stage_opamp_dummy_magic_14_0.Vb1.n15 two_stage_opamp_dummy_magic_14_0.Vb1.n14 176.733
R8044 two_stage_opamp_dummy_magic_14_0.Vb1.n11 two_stage_opamp_dummy_magic_14_0.Vb1.n10 176.733
R8045 two_stage_opamp_dummy_magic_14_0.Vb1.n12 two_stage_opamp_dummy_magic_14_0.Vb1.n11 176.733
R8046 two_stage_opamp_dummy_magic_14_0.Vb1.n13 two_stage_opamp_dummy_magic_14_0.Vb1.n12 176.733
R8047 two_stage_opamp_dummy_magic_14_0.Vb1.n8 two_stage_opamp_dummy_magic_14_0.Vb1.n7 176.733
R8048 two_stage_opamp_dummy_magic_14_0.Vb1.n7 two_stage_opamp_dummy_magic_14_0.Vb1.n6 176.733
R8049 two_stage_opamp_dummy_magic_14_0.Vb1.n6 two_stage_opamp_dummy_magic_14_0.Vb1.n5 176.733
R8050 two_stage_opamp_dummy_magic_14_0.Vb1.n2 two_stage_opamp_dummy_magic_14_0.Vb1.n1 176.733
R8051 two_stage_opamp_dummy_magic_14_0.Vb1.n3 two_stage_opamp_dummy_magic_14_0.Vb1.n2 176.733
R8052 two_stage_opamp_dummy_magic_14_0.Vb1.n4 two_stage_opamp_dummy_magic_14_0.Vb1.n3 176.733
R8053 two_stage_opamp_dummy_magic_14_0.Vb1.n19 two_stage_opamp_dummy_magic_14_0.Vb1.n9 173.207
R8054 two_stage_opamp_dummy_magic_14_0.Vb1.n19 two_stage_opamp_dummy_magic_14_0.Vb1.n18 165.8
R8055 two_stage_opamp_dummy_magic_14_0.Vb1.n26 two_stage_opamp_dummy_magic_14_0.Vb1.n24 152
R8056 two_stage_opamp_dummy_magic_14_0.Vb1.n21 two_stage_opamp_dummy_magic_14_0.Vb1.n20 113.906
R8057 two_stage_opamp_dummy_magic_14_0.Vb1.n29 two_stage_opamp_dummy_magic_14_0.Vb1.n28 113.906
R8058 two_stage_opamp_dummy_magic_14_0.Vb1.n26 two_stage_opamp_dummy_magic_14_0.Vb1.n25 100.106
R8059 two_stage_opamp_dummy_magic_14_0.Vb1.n21 two_stage_opamp_dummy_magic_14_0.Vb1.t15 65.0512
R8060 two_stage_opamp_dummy_magic_14_0.Vb1.n18 two_stage_opamp_dummy_magic_14_0.Vb1.n17 54.6272
R8061 two_stage_opamp_dummy_magic_14_0.Vb1.n18 two_stage_opamp_dummy_magic_14_0.Vb1.n13 54.6272
R8062 two_stage_opamp_dummy_magic_14_0.Vb1.n9 two_stage_opamp_dummy_magic_14_0.Vb1.n8 54.6272
R8063 two_stage_opamp_dummy_magic_14_0.Vb1.n9 two_stage_opamp_dummy_magic_14_0.Vb1.n4 54.6272
R8064 bgr_7_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb1.n30 45.8755
R8065 two_stage_opamp_dummy_magic_14_0.Vb1.n24 two_stage_opamp_dummy_magic_14_0.Vb1.n23 45.5227
R8066 two_stage_opamp_dummy_magic_14_0.Vb1.n24 two_stage_opamp_dummy_magic_14_0.Vb1.n22 45.5227
R8067 two_stage_opamp_dummy_magic_14_0.Vb1.n30 two_stage_opamp_dummy_magic_14_0.Vb1.n29 24.8755
R8068 two_stage_opamp_dummy_magic_14_0.Vb1.n0 two_stage_opamp_dummy_magic_14_0.Vb1.t0 19.7005
R8069 two_stage_opamp_dummy_magic_14_0.Vb1.n0 two_stage_opamp_dummy_magic_14_0.Vb1.t9 19.7005
R8070 two_stage_opamp_dummy_magic_14_0.Vb1.n25 two_stage_opamp_dummy_magic_14_0.Vb1.t2 16.0005
R8071 two_stage_opamp_dummy_magic_14_0.Vb1.n25 two_stage_opamp_dummy_magic_14_0.Vb1.t4 16.0005
R8072 two_stage_opamp_dummy_magic_14_0.Vb1.n20 two_stage_opamp_dummy_magic_14_0.Vb1.t10 16.0005
R8073 two_stage_opamp_dummy_magic_14_0.Vb1.n20 two_stage_opamp_dummy_magic_14_0.Vb1.t6 16.0005
R8074 two_stage_opamp_dummy_magic_14_0.Vb1.n28 two_stage_opamp_dummy_magic_14_0.Vb1.t8 16.0005
R8075 two_stage_opamp_dummy_magic_14_0.Vb1.n28 two_stage_opamp_dummy_magic_14_0.Vb1.t11 16.0005
R8076 two_stage_opamp_dummy_magic_14_0.Vb1.n27 two_stage_opamp_dummy_magic_14_0.Vb1.n26 13.8005
R8077 two_stage_opamp_dummy_magic_14_0.Vb1.n30 two_stage_opamp_dummy_magic_14_0.Vb1.n19 2.07862
R8078 two_stage_opamp_dummy_magic_14_0.Vb1.n27 two_stage_opamp_dummy_magic_14_0.Vb1.n21 0.563
R8079 two_stage_opamp_dummy_magic_14_0.Vb1.n29 two_stage_opamp_dummy_magic_14_0.Vb1.n27 0.563
R8080 two_stage_opamp_dummy_magic_14_0.VD1.n11 two_stage_opamp_dummy_magic_14_0.VD1.n9 146.47
R8081 two_stage_opamp_dummy_magic_14_0.VD1.n6 two_stage_opamp_dummy_magic_14_0.VD1.n4 146.47
R8082 two_stage_opamp_dummy_magic_14_0.VD1.n13 two_stage_opamp_dummy_magic_14_0.VD1.n12 145.906
R8083 two_stage_opamp_dummy_magic_14_0.VD1.n11 two_stage_opamp_dummy_magic_14_0.VD1.n10 145.906
R8084 two_stage_opamp_dummy_magic_14_0.VD1.n8 two_stage_opamp_dummy_magic_14_0.VD1.n7 145.906
R8085 two_stage_opamp_dummy_magic_14_0.VD1.n6 two_stage_opamp_dummy_magic_14_0.VD1.n5 145.906
R8086 two_stage_opamp_dummy_magic_14_0.VD1.n19 two_stage_opamp_dummy_magic_14_0.VD1.n18 114.469
R8087 two_stage_opamp_dummy_magic_14_0.VD1.n2 two_stage_opamp_dummy_magic_14_0.VD1.n0 114.469
R8088 two_stage_opamp_dummy_magic_14_0.VD1.n18 two_stage_opamp_dummy_magic_14_0.VD1.n17 113.906
R8089 two_stage_opamp_dummy_magic_14_0.VD1.n2 two_stage_opamp_dummy_magic_14_0.VD1.n1 113.906
R8090 two_stage_opamp_dummy_magic_14_0.VD1.n15 two_stage_opamp_dummy_magic_14_0.VD1.n3 109.406
R8091 two_stage_opamp_dummy_magic_14_0.VD1.n17 two_stage_opamp_dummy_magic_14_0.VD1.t7 16.0005
R8092 two_stage_opamp_dummy_magic_14_0.VD1.n17 two_stage_opamp_dummy_magic_14_0.VD1.t12 16.0005
R8093 two_stage_opamp_dummy_magic_14_0.VD1.n3 two_stage_opamp_dummy_magic_14_0.VD1.t9 16.0005
R8094 two_stage_opamp_dummy_magic_14_0.VD1.n3 two_stage_opamp_dummy_magic_14_0.VD1.t4 16.0005
R8095 two_stage_opamp_dummy_magic_14_0.VD1.n12 two_stage_opamp_dummy_magic_14_0.VD1.t2 16.0005
R8096 two_stage_opamp_dummy_magic_14_0.VD1.n12 two_stage_opamp_dummy_magic_14_0.VD1.t16 16.0005
R8097 two_stage_opamp_dummy_magic_14_0.VD1.n10 two_stage_opamp_dummy_magic_14_0.VD1.t14 16.0005
R8098 two_stage_opamp_dummy_magic_14_0.VD1.n10 two_stage_opamp_dummy_magic_14_0.VD1.t1 16.0005
R8099 two_stage_opamp_dummy_magic_14_0.VD1.n9 two_stage_opamp_dummy_magic_14_0.VD1.t3 16.0005
R8100 two_stage_opamp_dummy_magic_14_0.VD1.n9 two_stage_opamp_dummy_magic_14_0.VD1.t19 16.0005
R8101 two_stage_opamp_dummy_magic_14_0.VD1.n7 two_stage_opamp_dummy_magic_14_0.VD1.t17 16.0005
R8102 two_stage_opamp_dummy_magic_14_0.VD1.n7 two_stage_opamp_dummy_magic_14_0.VD1.t21 16.0005
R8103 two_stage_opamp_dummy_magic_14_0.VD1.n5 two_stage_opamp_dummy_magic_14_0.VD1.t0 16.0005
R8104 two_stage_opamp_dummy_magic_14_0.VD1.n5 two_stage_opamp_dummy_magic_14_0.VD1.t15 16.0005
R8105 two_stage_opamp_dummy_magic_14_0.VD1.n4 two_stage_opamp_dummy_magic_14_0.VD1.t18 16.0005
R8106 two_stage_opamp_dummy_magic_14_0.VD1.n4 two_stage_opamp_dummy_magic_14_0.VD1.t20 16.0005
R8107 two_stage_opamp_dummy_magic_14_0.VD1.n1 two_stage_opamp_dummy_magic_14_0.VD1.t10 16.0005
R8108 two_stage_opamp_dummy_magic_14_0.VD1.n1 two_stage_opamp_dummy_magic_14_0.VD1.t5 16.0005
R8109 two_stage_opamp_dummy_magic_14_0.VD1.n0 two_stage_opamp_dummy_magic_14_0.VD1.t11 16.0005
R8110 two_stage_opamp_dummy_magic_14_0.VD1.n0 two_stage_opamp_dummy_magic_14_0.VD1.t6 16.0005
R8111 two_stage_opamp_dummy_magic_14_0.VD1.n19 two_stage_opamp_dummy_magic_14_0.VD1.t8 16.0005
R8112 two_stage_opamp_dummy_magic_14_0.VD1.t13 two_stage_opamp_dummy_magic_14_0.VD1.n19 16.0005
R8113 two_stage_opamp_dummy_magic_14_0.VD1.n15 two_stage_opamp_dummy_magic_14_0.VD1.n14 5.11508
R8114 two_stage_opamp_dummy_magic_14_0.VD1.n16 two_stage_opamp_dummy_magic_14_0.VD1.n15 4.5005
R8115 two_stage_opamp_dummy_magic_14_0.VD1.n13 two_stage_opamp_dummy_magic_14_0.VD1.n11 0.563
R8116 two_stage_opamp_dummy_magic_14_0.VD1.n8 two_stage_opamp_dummy_magic_14_0.VD1.n6 0.563
R8117 two_stage_opamp_dummy_magic_14_0.VD1.n16 two_stage_opamp_dummy_magic_14_0.VD1.n2 0.563
R8118 two_stage_opamp_dummy_magic_14_0.VD1.n18 two_stage_opamp_dummy_magic_14_0.VD1.n16 0.563
R8119 two_stage_opamp_dummy_magic_14_0.VD1.n14 two_stage_opamp_dummy_magic_14_0.VD1.n13 0.234875
R8120 two_stage_opamp_dummy_magic_14_0.VD1.n14 two_stage_opamp_dummy_magic_14_0.VD1.n8 0.234875
R8121 a_6930_22564.t0 a_6930_22564.t1 178.133
R8122 bgr_7_0.PFET_GATE_10uA.n16 bgr_7_0.PFET_GATE_10uA.t18 565.114
R8123 bgr_7_0.PFET_GATE_10uA.n19 bgr_7_0.PFET_GATE_10uA.t15 530.201
R8124 bgr_7_0.PFET_GATE_10uA.n21 bgr_7_0.PFET_GATE_10uA.t14 409.7
R8125 bgr_7_0.PFET_GATE_10uA.n6 bgr_7_0.PFET_GATE_10uA.t12 369.534
R8126 bgr_7_0.PFET_GATE_10uA.n5 bgr_7_0.PFET_GATE_10uA.t11 369.534
R8127 bgr_7_0.PFET_GATE_10uA.n2 bgr_7_0.PFET_GATE_10uA.t20 369.534
R8128 bgr_7_0.PFET_GATE_10uA.n1 bgr_7_0.PFET_GATE_10uA.t19 369.534
R8129 bgr_7_0.PFET_GATE_10uA.n19 bgr_7_0.PFET_GATE_10uA.t21 353.467
R8130 bgr_7_0.PFET_GATE_10uA.n20 bgr_7_0.PFET_GATE_10uA.t10 353.467
R8131 bgr_7_0.PFET_GATE_10uA.n10 bgr_7_0.PFET_GATE_10uA.n8 341.397
R8132 bgr_7_0.PFET_GATE_10uA.n12 bgr_7_0.PFET_GATE_10uA.n11 339.272
R8133 bgr_7_0.PFET_GATE_10uA.n10 bgr_7_0.PFET_GATE_10uA.n9 339.272
R8134 bgr_7_0.PFET_GATE_10uA.n15 bgr_7_0.PFET_GATE_10uA.n14 334.772
R8135 bgr_7_0.PFET_GATE_10uA.n0 bgr_7_0.PFET_GATE_10uA.t17 325.351
R8136 bgr_7_0.PFET_GATE_10uA.n4 bgr_7_0.PFET_GATE_10uA.n0 202.364
R8137 bgr_7_0.PFET_GATE_10uA.n6 bgr_7_0.PFET_GATE_10uA.t22 192.8
R8138 bgr_7_0.PFET_GATE_10uA.n5 bgr_7_0.PFET_GATE_10uA.t16 192.8
R8139 bgr_7_0.PFET_GATE_10uA.n2 bgr_7_0.PFET_GATE_10uA.t13 192.8
R8140 bgr_7_0.PFET_GATE_10uA.n1 bgr_7_0.PFET_GATE_10uA.t24 192.8
R8141 bgr_7_0.PFET_GATE_10uA.n0 bgr_7_0.PFET_GATE_10uA.t23 192.8
R8142 bgr_7_0.PFET_GATE_10uA.n20 bgr_7_0.PFET_GATE_10uA.n19 176.733
R8143 bgr_7_0.PFET_GATE_10uA.n18 bgr_7_0.PFET_GATE_10uA.n7 168.166
R8144 bgr_7_0.PFET_GATE_10uA bgr_7_0.PFET_GATE_10uA.n21 166.071
R8145 bgr_7_0.PFET_GATE_10uA.n4 bgr_7_0.PFET_GATE_10uA.n3 166.071
R8146 bgr_7_0.PFET_GATE_10uA.n16 bgr_7_0.PFET_GATE_10uA.t6 137.386
R8147 bgr_7_0.PFET_GATE_10uA.n13 bgr_7_0.PFET_GATE_10uA.t9 100.635
R8148 bgr_7_0.PFET_GATE_10uA.n7 bgr_7_0.PFET_GATE_10uA.n6 56.2338
R8149 bgr_7_0.PFET_GATE_10uA.n7 bgr_7_0.PFET_GATE_10uA.n5 56.2338
R8150 bgr_7_0.PFET_GATE_10uA.n21 bgr_7_0.PFET_GATE_10uA.n20 56.2338
R8151 bgr_7_0.PFET_GATE_10uA.n3 bgr_7_0.PFET_GATE_10uA.n2 56.2338
R8152 bgr_7_0.PFET_GATE_10uA.n3 bgr_7_0.PFET_GATE_10uA.n1 56.2338
R8153 bgr_7_0.PFET_GATE_10uA.n14 bgr_7_0.PFET_GATE_10uA.t8 39.4005
R8154 bgr_7_0.PFET_GATE_10uA.n14 bgr_7_0.PFET_GATE_10uA.t1 39.4005
R8155 bgr_7_0.PFET_GATE_10uA.n11 bgr_7_0.PFET_GATE_10uA.t3 39.4005
R8156 bgr_7_0.PFET_GATE_10uA.n11 bgr_7_0.PFET_GATE_10uA.t5 39.4005
R8157 bgr_7_0.PFET_GATE_10uA.n9 bgr_7_0.PFET_GATE_10uA.t2 39.4005
R8158 bgr_7_0.PFET_GATE_10uA.n9 bgr_7_0.PFET_GATE_10uA.t4 39.4005
R8159 bgr_7_0.PFET_GATE_10uA.n8 bgr_7_0.PFET_GATE_10uA.t0 39.4005
R8160 bgr_7_0.PFET_GATE_10uA.n8 bgr_7_0.PFET_GATE_10uA.t7 39.4005
R8161 bgr_7_0.PFET_GATE_10uA.n18 bgr_7_0.PFET_GATE_10uA.n17 27.5005
R8162 bgr_7_0.PFET_GATE_10uA.n17 bgr_7_0.PFET_GATE_10uA.n15 9.53175
R8163 bgr_7_0.PFET_GATE_10uA bgr_7_0.PFET_GATE_10uA.n4 5.2505
R8164 bgr_7_0.PFET_GATE_10uA.n15 bgr_7_0.PFET_GATE_10uA.n13 4.5005
R8165 bgr_7_0.PFET_GATE_10uA bgr_7_0.PFET_GATE_10uA.n18 2.34425
R8166 bgr_7_0.PFET_GATE_10uA.n12 bgr_7_0.PFET_GATE_10uA.n10 2.1255
R8167 bgr_7_0.PFET_GATE_10uA.n13 bgr_7_0.PFET_GATE_10uA.n12 2.1255
R8168 bgr_7_0.PFET_GATE_10uA.n17 bgr_7_0.PFET_GATE_10uA.n16 1.78175
R8169 bgr_7_0.cap_res1.t0 bgr_7_0.cap_res1.t10 121.245
R8170 bgr_7_0.cap_res1.t16 bgr_7_0.cap_res1.t19 0.1603
R8171 bgr_7_0.cap_res1.t9 bgr_7_0.cap_res1.t15 0.1603
R8172 bgr_7_0.cap_res1.t14 bgr_7_0.cap_res1.t18 0.1603
R8173 bgr_7_0.cap_res1.t7 bgr_7_0.cap_res1.t13 0.1603
R8174 bgr_7_0.cap_res1.t1 bgr_7_0.cap_res1.t6 0.1603
R8175 bgr_7_0.cap_res1.n1 bgr_7_0.cap_res1.t17 0.159278
R8176 bgr_7_0.cap_res1.n2 bgr_7_0.cap_res1.t2 0.159278
R8177 bgr_7_0.cap_res1.n3 bgr_7_0.cap_res1.t8 0.159278
R8178 bgr_7_0.cap_res1.n4 bgr_7_0.cap_res1.t3 0.159278
R8179 bgr_7_0.cap_res1.n4 bgr_7_0.cap_res1.t16 0.1368
R8180 bgr_7_0.cap_res1.n4 bgr_7_0.cap_res1.t12 0.1368
R8181 bgr_7_0.cap_res1.n3 bgr_7_0.cap_res1.t9 0.1368
R8182 bgr_7_0.cap_res1.n3 bgr_7_0.cap_res1.t5 0.1368
R8183 bgr_7_0.cap_res1.n2 bgr_7_0.cap_res1.t14 0.1368
R8184 bgr_7_0.cap_res1.n2 bgr_7_0.cap_res1.t11 0.1368
R8185 bgr_7_0.cap_res1.n1 bgr_7_0.cap_res1.t7 0.1368
R8186 bgr_7_0.cap_res1.n1 bgr_7_0.cap_res1.t4 0.1368
R8187 bgr_7_0.cap_res1.n0 bgr_7_0.cap_res1.t1 0.1368
R8188 bgr_7_0.cap_res1.n0 bgr_7_0.cap_res1.t20 0.1368
R8189 bgr_7_0.cap_res1.t17 bgr_7_0.cap_res1.n0 0.00152174
R8190 bgr_7_0.cap_res1.t2 bgr_7_0.cap_res1.n1 0.00152174
R8191 bgr_7_0.cap_res1.t8 bgr_7_0.cap_res1.n2 0.00152174
R8192 bgr_7_0.cap_res1.t3 bgr_7_0.cap_res1.n3 0.00152174
R8193 bgr_7_0.cap_res1.t10 bgr_7_0.cap_res1.n4 0.00152174
R8194 bgr_7_0.V_mir2.n20 bgr_7_0.V_mir2.n19 325.473
R8195 bgr_7_0.V_mir2.n13 bgr_7_0.V_mir2.n12 325.473
R8196 bgr_7_0.V_mir2.n8 bgr_7_0.V_mir2.n7 325.473
R8197 bgr_7_0.V_mir2.n16 bgr_7_0.V_mir2.t21 310.488
R8198 bgr_7_0.V_mir2.n9 bgr_7_0.V_mir2.t22 310.488
R8199 bgr_7_0.V_mir2.n4 bgr_7_0.V_mir2.t20 310.488
R8200 bgr_7_0.V_mir2.n2 bgr_7_0.V_mir2.t14 278.312
R8201 bgr_7_0.V_mir2.n2 bgr_7_0.V_mir2.n1 228.939
R8202 bgr_7_0.V_mir2.n3 bgr_7_0.V_mir2.n0 224.439
R8203 bgr_7_0.V_mir2.n18 bgr_7_0.V_mir2.t10 184.097
R8204 bgr_7_0.V_mir2.n11 bgr_7_0.V_mir2.t8 184.097
R8205 bgr_7_0.V_mir2.n6 bgr_7_0.V_mir2.t0 184.097
R8206 bgr_7_0.V_mir2.n17 bgr_7_0.V_mir2.n16 167.094
R8207 bgr_7_0.V_mir2.n10 bgr_7_0.V_mir2.n9 167.094
R8208 bgr_7_0.V_mir2.n5 bgr_7_0.V_mir2.n4 167.094
R8209 bgr_7_0.V_mir2.n13 bgr_7_0.V_mir2.n11 152
R8210 bgr_7_0.V_mir2.n8 bgr_7_0.V_mir2.n6 152
R8211 bgr_7_0.V_mir2.n19 bgr_7_0.V_mir2.n18 152
R8212 bgr_7_0.V_mir2.n16 bgr_7_0.V_mir2.t19 120.501
R8213 bgr_7_0.V_mir2.n17 bgr_7_0.V_mir2.t6 120.501
R8214 bgr_7_0.V_mir2.n9 bgr_7_0.V_mir2.t18 120.501
R8215 bgr_7_0.V_mir2.n10 bgr_7_0.V_mir2.t2 120.501
R8216 bgr_7_0.V_mir2.n4 bgr_7_0.V_mir2.t17 120.501
R8217 bgr_7_0.V_mir2.n5 bgr_7_0.V_mir2.t4 120.501
R8218 bgr_7_0.V_mir2.n1 bgr_7_0.V_mir2.t16 48.0005
R8219 bgr_7_0.V_mir2.n1 bgr_7_0.V_mir2.t12 48.0005
R8220 bgr_7_0.V_mir2.n0 bgr_7_0.V_mir2.t15 48.0005
R8221 bgr_7_0.V_mir2.n0 bgr_7_0.V_mir2.t13 48.0005
R8222 bgr_7_0.V_mir2.n18 bgr_7_0.V_mir2.n17 40.7027
R8223 bgr_7_0.V_mir2.n11 bgr_7_0.V_mir2.n10 40.7027
R8224 bgr_7_0.V_mir2.n6 bgr_7_0.V_mir2.n5 40.7027
R8225 bgr_7_0.V_mir2.n12 bgr_7_0.V_mir2.t3 39.4005
R8226 bgr_7_0.V_mir2.n12 bgr_7_0.V_mir2.t9 39.4005
R8227 bgr_7_0.V_mir2.n7 bgr_7_0.V_mir2.t5 39.4005
R8228 bgr_7_0.V_mir2.n7 bgr_7_0.V_mir2.t1 39.4005
R8229 bgr_7_0.V_mir2.n20 bgr_7_0.V_mir2.t7 39.4005
R8230 bgr_7_0.V_mir2.t11 bgr_7_0.V_mir2.n20 39.4005
R8231 bgr_7_0.V_mir2.n14 bgr_7_0.V_mir2.n13 15.8005
R8232 bgr_7_0.V_mir2.n14 bgr_7_0.V_mir2.n8 15.8005
R8233 bgr_7_0.V_mir2.n19 bgr_7_0.V_mir2.n15 9.3005
R8234 bgr_7_0.V_mir2.n3 bgr_7_0.V_mir2.n2 5.8755
R8235 bgr_7_0.V_mir2.n15 bgr_7_0.V_mir2.n14 4.5005
R8236 bgr_7_0.V_mir2.n15 bgr_7_0.V_mir2.n3 0.78175
R8237 bgr_7_0.Vin-.n8 bgr_7_0.Vin-.t12 688.859
R8238 bgr_7_0.Vin-.n10 bgr_7_0.Vin-.n9 514.134
R8239 bgr_7_0.Vin-.n7 bgr_7_0.Vin-.n6 351.522
R8240 bgr_7_0.Vin-.n12 bgr_7_0.Vin-.n11 213.4
R8241 bgr_7_0.Vin-.n8 bgr_7_0.Vin-.t8 174.726
R8242 bgr_7_0.Vin-.n9 bgr_7_0.Vin-.t10 174.726
R8243 bgr_7_0.Vin-.n10 bgr_7_0.Vin-.t9 174.726
R8244 bgr_7_0.Vin-.n11 bgr_7_0.Vin-.t11 174.726
R8245 bgr_7_0.Vin-.n5 bgr_7_0.Vin-.n3 173.029
R8246 bgr_7_0.Vin-.n5 bgr_7_0.Vin-.n4 168.654
R8247 bgr_7_0.Vin-.n22 bgr_7_0.Vin-.n21 141.667
R8248 bgr_7_0.Vin-.n9 bgr_7_0.Vin-.n8 128.534
R8249 bgr_7_0.Vin-.n11 bgr_7_0.Vin-.n10 128.534
R8250 bgr_7_0.Vin-.n13 bgr_7_0.Vin-.t7 119.099
R8251 bgr_7_0.Vin-.n23 bgr_7_0.Vin-.n22 84.0884
R8252 bgr_7_0.Vin-.n18 bgr_7_0.Vin-.n17 83.5719
R8253 bgr_7_0.Vin-.n19 bgr_7_0.Vin-.n0 83.5719
R8254 bgr_7_0.Vin-.n20 bgr_7_0.Vin-.n1 83.5719
R8255 bgr_7_0.Vin-.n15 bgr_7_0.Vin-.t2 65.0299
R8256 bgr_7_0.Vin-.n6 bgr_7_0.Vin-.t0 39.4005
R8257 bgr_7_0.Vin-.n6 bgr_7_0.Vin-.t1 39.4005
R8258 bgr_7_0.Vin-.n14 bgr_7_0.Vin-.n13 28.813
R8259 bgr_7_0.Vin-.n19 bgr_7_0.Vin-.n18 26.074
R8260 bgr_7_0.Vin-.n20 bgr_7_0.Vin-.n19 26.074
R8261 bgr_7_0.Vin-.n22 bgr_7_0.Vin-.n20 26.074
R8262 bgr_7_0.Vin-.n13 bgr_7_0.Vin-.n12 16.188
R8263 bgr_7_0.Vin-.n4 bgr_7_0.Vin-.t3 13.1338
R8264 bgr_7_0.Vin-.n4 bgr_7_0.Vin-.t5 13.1338
R8265 bgr_7_0.Vin-.n3 bgr_7_0.Vin-.t6 13.1338
R8266 bgr_7_0.Vin-.n3 bgr_7_0.Vin-.t4 13.1338
R8267 bgr_7_0.Vin-.n12 bgr_7_0.Vin-.n7 11.2193
R8268 bgr_7_0.Vin-.n7 bgr_7_0.Vin-.n5 3.8755
R8269 bgr_7_0.Vin-.n24 bgr_7_0.Vin-.n23 1.56836
R8270 bgr_7_0.Vin-.n17 bgr_7_0.Vin-.n15 1.56363
R8271 bgr_7_0.Vin-.n25 bgr_7_0.Vin-.n24 1.5505
R8272 bgr_7_0.Vin-.n16 bgr_7_0.Vin-.n2 1.5505
R8273 bgr_7_0.Vin-.n23 bgr_7_0.Vin-.n1 1.14402
R8274 bgr_7_0.Vin-.n16 bgr_7_0.Vin-.n0 0.885803
R8275 bgr_7_0.Vin-.n17 bgr_7_0.Vin-.n16 0.77514
R8276 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_7_0.Vin-.n0 0.756696
R8277 bgr_7_0.Vin-.n25 bgr_7_0.Vin-.n1 0.701365
R8278 bgr_7_0.Vin-.n15 bgr_7_0.Vin-.n14 0.530034
R8279 bgr_7_0.Vin-.n18 bgr_7_0.Vin-.t2 0.290206
R8280 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_7_0.Vin-.n25 0.203382
R8281 bgr_7_0.Vin-.n24 bgr_7_0.Vin-.n2 0.0183571
R8282 bgr_7_0.Vin-.n14 bgr_7_0.Vin-.n2 0.00817857
R8283 bgr_7_0.V_p_1.n1 bgr_7_0.V_p_1.n5 229.562
R8284 bgr_7_0.V_p_1.n1 bgr_7_0.V_p_1.n4 228.939
R8285 bgr_7_0.V_p_1.n0 bgr_7_0.V_p_1.n3 228.939
R8286 bgr_7_0.V_p_1.n0 bgr_7_0.V_p_1.n2 228.939
R8287 bgr_7_0.V_p_1.n6 bgr_7_0.V_p_1.n1 228.938
R8288 bgr_7_0.V_p_1.n0 bgr_7_0.V_p_1.t5 98.7279
R8289 bgr_7_0.V_p_1.n5 bgr_7_0.V_p_1.t8 48.0005
R8290 bgr_7_0.V_p_1.n5 bgr_7_0.V_p_1.t0 48.0005
R8291 bgr_7_0.V_p_1.n4 bgr_7_0.V_p_1.t10 48.0005
R8292 bgr_7_0.V_p_1.n4 bgr_7_0.V_p_1.t2 48.0005
R8293 bgr_7_0.V_p_1.n3 bgr_7_0.V_p_1.t3 48.0005
R8294 bgr_7_0.V_p_1.n3 bgr_7_0.V_p_1.t6 48.0005
R8295 bgr_7_0.V_p_1.n2 bgr_7_0.V_p_1.t9 48.0005
R8296 bgr_7_0.V_p_1.n2 bgr_7_0.V_p_1.t1 48.0005
R8297 bgr_7_0.V_p_1.t4 bgr_7_0.V_p_1.n6 48.0005
R8298 bgr_7_0.V_p_1.n6 bgr_7_0.V_p_1.t7 48.0005
R8299 bgr_7_0.V_p_1.n1 bgr_7_0.V_p_1.n0 1.8755
R8300 VIN-.n9 VIN-.t1 490.572
R8301 VIN-.n4 VIN-.t2 449.868
R8302 VIN-.n0 VIN-.t4 449.868
R8303 VIN-.n4 VIN-.t7 273.134
R8304 VIN-.n5 VIN-.t3 273.134
R8305 VIN-.n6 VIN-.t8 273.134
R8306 VIN-.n7 VIN-.t0 273.134
R8307 VIN-.n3 VIN-.t6 273.134
R8308 VIN-.n2 VIN-.t10 273.134
R8309 VIN-.n1 VIN-.t5 273.134
R8310 VIN-.n0 VIN-.t9 273.134
R8311 VIN-.n7 VIN-.n6 176.733
R8312 VIN-.n6 VIN-.n5 176.733
R8313 VIN-.n5 VIN-.n4 176.733
R8314 VIN-.n1 VIN-.n0 176.733
R8315 VIN-.n2 VIN-.n1 176.733
R8316 VIN-.n3 VIN-.n2 176.733
R8317 VIN-.n9 VIN-.n8 165.8
R8318 VIN-.n8 VIN-.n7 56.2338
R8319 VIN-.n8 VIN-.n3 56.2338
R8320 VIN- VIN-.n9 2.14112
R8321 two_stage_opamp_dummy_magic_14_0.Vb1_2.n2 two_stage_opamp_dummy_magic_14_0.Vb1_2.n1 114.469
R8322 two_stage_opamp_dummy_magic_14_0.Vb1_2.n1 two_stage_opamp_dummy_magic_14_0.Vb1_2.n0 113.906
R8323 two_stage_opamp_dummy_magic_14_0.Vb1_2.n1 two_stage_opamp_dummy_magic_14_0.Vb1_2.t4 96.77
R8324 two_stage_opamp_dummy_magic_14_0.Vb1_2.n0 two_stage_opamp_dummy_magic_14_0.Vb1_2.t0 16.0005
R8325 two_stage_opamp_dummy_magic_14_0.Vb1_2.n0 two_stage_opamp_dummy_magic_14_0.Vb1_2.t2 16.0005
R8326 two_stage_opamp_dummy_magic_14_0.Vb1_2.t3 two_stage_opamp_dummy_magic_14_0.Vb1_2.n2 16.0005
R8327 two_stage_opamp_dummy_magic_14_0.Vb1_2.n2 two_stage_opamp_dummy_magic_14_0.Vb1_2.t1 16.0005
R8328 two_stage_opamp_dummy_magic_14_0.VD4.n28 two_stage_opamp_dummy_magic_14_0.VD4.t23 652.076
R8329 two_stage_opamp_dummy_magic_14_0.VD4.n61 two_stage_opamp_dummy_magic_14_0.VD4.t20 652.076
R8330 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n13 585
R8331 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n41 585
R8332 two_stage_opamp_dummy_magic_14_0.VD4.n48 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8333 two_stage_opamp_dummy_magic_14_0.VD4.n54 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8334 two_stage_opamp_dummy_magic_14_0.VD4.n49 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8335 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n30 290.233
R8336 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n35 290.233
R8337 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n40 290.233
R8338 two_stage_opamp_dummy_magic_14_0.VD4.n49 two_stage_opamp_dummy_magic_14_0.VD4.n46 242.903
R8339 two_stage_opamp_dummy_magic_14_0.VD4.n40 two_stage_opamp_dummy_magic_14_0.VD4.n18 242.903
R8340 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n59 238.367
R8341 two_stage_opamp_dummy_magic_14_0.VD4.n15 two_stage_opamp_dummy_magic_14_0.VD4.n14 185
R8342 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n56 185
R8343 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n57 185
R8344 two_stage_opamp_dummy_magic_14_0.VD4.n55 two_stage_opamp_dummy_magic_14_0.VD4.n47 185
R8345 two_stage_opamp_dummy_magic_14_0.VD4.n53 two_stage_opamp_dummy_magic_14_0.VD4.n52 185
R8346 two_stage_opamp_dummy_magic_14_0.VD4.n51 two_stage_opamp_dummy_magic_14_0.VD4.n50 185
R8347 two_stage_opamp_dummy_magic_14_0.VD4.n43 two_stage_opamp_dummy_magic_14_0.VD4.n42 185
R8348 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n43 185
R8349 two_stage_opamp_dummy_magic_14_0.VD4.n29 two_stage_opamp_dummy_magic_14_0.VD4.n19 185
R8350 two_stage_opamp_dummy_magic_14_0.VD4.n32 two_stage_opamp_dummy_magic_14_0.VD4.n31 185
R8351 two_stage_opamp_dummy_magic_14_0.VD4.n34 two_stage_opamp_dummy_magic_14_0.VD4.n33 185
R8352 two_stage_opamp_dummy_magic_14_0.VD4.n37 two_stage_opamp_dummy_magic_14_0.VD4.n36 185
R8353 two_stage_opamp_dummy_magic_14_0.VD4.n39 two_stage_opamp_dummy_magic_14_0.VD4.n38 185
R8354 two_stage_opamp_dummy_magic_14_0.VD4.t24 two_stage_opamp_dummy_magic_14_0.VD4.n44 170.513
R8355 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.t21 170.513
R8356 two_stage_opamp_dummy_magic_14_0.VD4.n2 two_stage_opamp_dummy_magic_14_0.VD4.n0 163.626
R8357 two_stage_opamp_dummy_magic_14_0.VD4.n10 two_stage_opamp_dummy_magic_14_0.VD4.n9 163.001
R8358 two_stage_opamp_dummy_magic_14_0.VD4.n8 two_stage_opamp_dummy_magic_14_0.VD4.n7 163.001
R8359 two_stage_opamp_dummy_magic_14_0.VD4.n6 two_stage_opamp_dummy_magic_14_0.VD4.n5 163.001
R8360 two_stage_opamp_dummy_magic_14_0.VD4.n4 two_stage_opamp_dummy_magic_14_0.VD4.n3 163.001
R8361 two_stage_opamp_dummy_magic_14_0.VD4.n2 two_stage_opamp_dummy_magic_14_0.VD4.n1 163.001
R8362 two_stage_opamp_dummy_magic_14_0.VD4.n12 two_stage_opamp_dummy_magic_14_0.VD4.n11 159.804
R8363 two_stage_opamp_dummy_magic_14_0.VD4.n21 two_stage_opamp_dummy_magic_14_0.VD4.n20 159.803
R8364 two_stage_opamp_dummy_magic_14_0.VD4.n23 two_stage_opamp_dummy_magic_14_0.VD4.n22 159.803
R8365 two_stage_opamp_dummy_magic_14_0.VD4.n25 two_stage_opamp_dummy_magic_14_0.VD4.n24 159.803
R8366 two_stage_opamp_dummy_magic_14_0.VD4.n27 two_stage_opamp_dummy_magic_14_0.VD4.n26 159.803
R8367 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n15 150
R8368 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n47 150
R8369 two_stage_opamp_dummy_magic_14_0.VD4.n52 two_stage_opamp_dummy_magic_14_0.VD4.n51 150
R8370 two_stage_opamp_dummy_magic_14_0.VD4.n43 two_stage_opamp_dummy_magic_14_0.VD4.n19 150
R8371 two_stage_opamp_dummy_magic_14_0.VD4.n33 two_stage_opamp_dummy_magic_14_0.VD4.n32 150
R8372 two_stage_opamp_dummy_magic_14_0.VD4.n38 two_stage_opamp_dummy_magic_14_0.VD4.n37 150
R8373 two_stage_opamp_dummy_magic_14_0.VD4.t10 two_stage_opamp_dummy_magic_14_0.VD4.t24 146.155
R8374 two_stage_opamp_dummy_magic_14_0.VD4.t6 two_stage_opamp_dummy_magic_14_0.VD4.t10 146.155
R8375 two_stage_opamp_dummy_magic_14_0.VD4.t12 two_stage_opamp_dummy_magic_14_0.VD4.t6 146.155
R8376 two_stage_opamp_dummy_magic_14_0.VD4.t16 two_stage_opamp_dummy_magic_14_0.VD4.t12 146.155
R8377 two_stage_opamp_dummy_magic_14_0.VD4.t0 two_stage_opamp_dummy_magic_14_0.VD4.t16 146.155
R8378 two_stage_opamp_dummy_magic_14_0.VD4.t2 two_stage_opamp_dummy_magic_14_0.VD4.t0 146.155
R8379 two_stage_opamp_dummy_magic_14_0.VD4.t4 two_stage_opamp_dummy_magic_14_0.VD4.t2 146.155
R8380 two_stage_opamp_dummy_magic_14_0.VD4.t8 two_stage_opamp_dummy_magic_14_0.VD4.t4 146.155
R8381 two_stage_opamp_dummy_magic_14_0.VD4.t14 two_stage_opamp_dummy_magic_14_0.VD4.t8 146.155
R8382 two_stage_opamp_dummy_magic_14_0.VD4.t18 two_stage_opamp_dummy_magic_14_0.VD4.t14 146.155
R8383 two_stage_opamp_dummy_magic_14_0.VD4.t21 two_stage_opamp_dummy_magic_14_0.VD4.t18 146.155
R8384 two_stage_opamp_dummy_magic_14_0.VD4.n59 two_stage_opamp_dummy_magic_14_0.VD4.n58 65.8183
R8385 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n45 65.8183
R8386 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n46 65.8183
R8387 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n16 65.8183
R8388 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n17 65.8183
R8389 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n18 65.8183
R8390 two_stage_opamp_dummy_magic_14_0.VD4.n47 two_stage_opamp_dummy_magic_14_0.VD4.n45 53.3664
R8391 two_stage_opamp_dummy_magic_14_0.VD4.n51 two_stage_opamp_dummy_magic_14_0.VD4.n46 53.3664
R8392 two_stage_opamp_dummy_magic_14_0.VD4.n59 two_stage_opamp_dummy_magic_14_0.VD4.n15 53.3664
R8393 two_stage_opamp_dummy_magic_14_0.VD4.n52 two_stage_opamp_dummy_magic_14_0.VD4.n45 53.3664
R8394 two_stage_opamp_dummy_magic_14_0.VD4.n19 two_stage_opamp_dummy_magic_14_0.VD4.n16 53.3664
R8395 two_stage_opamp_dummy_magic_14_0.VD4.n33 two_stage_opamp_dummy_magic_14_0.VD4.n17 53.3664
R8396 two_stage_opamp_dummy_magic_14_0.VD4.n38 two_stage_opamp_dummy_magic_14_0.VD4.n18 53.3664
R8397 two_stage_opamp_dummy_magic_14_0.VD4.n32 two_stage_opamp_dummy_magic_14_0.VD4.n16 53.3664
R8398 two_stage_opamp_dummy_magic_14_0.VD4.n37 two_stage_opamp_dummy_magic_14_0.VD4.n17 53.3664
R8399 two_stage_opamp_dummy_magic_14_0.VD4.n61 two_stage_opamp_dummy_magic_14_0.VD4.n60 22.8576
R8400 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n28 22.8576
R8401 two_stage_opamp_dummy_magic_14_0.VD4.n28 two_stage_opamp_dummy_magic_14_0.VD4.n27 14.4255
R8402 two_stage_opamp_dummy_magic_14_0.VD4.n62 two_stage_opamp_dummy_magic_14_0.VD4.n61 13.8005
R8403 two_stage_opamp_dummy_magic_14_0.VD4.n20 two_stage_opamp_dummy_magic_14_0.VD4.t5 11.2576
R8404 two_stage_opamp_dummy_magic_14_0.VD4.n20 two_stage_opamp_dummy_magic_14_0.VD4.t9 11.2576
R8405 two_stage_opamp_dummy_magic_14_0.VD4.n22 two_stage_opamp_dummy_magic_14_0.VD4.t1 11.2576
R8406 two_stage_opamp_dummy_magic_14_0.VD4.n22 two_stage_opamp_dummy_magic_14_0.VD4.t3 11.2576
R8407 two_stage_opamp_dummy_magic_14_0.VD4.n24 two_stage_opamp_dummy_magic_14_0.VD4.t13 11.2576
R8408 two_stage_opamp_dummy_magic_14_0.VD4.n24 two_stage_opamp_dummy_magic_14_0.VD4.t17 11.2576
R8409 two_stage_opamp_dummy_magic_14_0.VD4.n26 two_stage_opamp_dummy_magic_14_0.VD4.t11 11.2576
R8410 two_stage_opamp_dummy_magic_14_0.VD4.n26 two_stage_opamp_dummy_magic_14_0.VD4.t7 11.2576
R8411 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.t25 11.2576
R8412 two_stage_opamp_dummy_magic_14_0.VD4.n13 two_stage_opamp_dummy_magic_14_0.VD4.t22 11.2576
R8413 two_stage_opamp_dummy_magic_14_0.VD4.n9 two_stage_opamp_dummy_magic_14_0.VD4.t26 11.2576
R8414 two_stage_opamp_dummy_magic_14_0.VD4.n9 two_stage_opamp_dummy_magic_14_0.VD4.t29 11.2576
R8415 two_stage_opamp_dummy_magic_14_0.VD4.n7 two_stage_opamp_dummy_magic_14_0.VD4.t32 11.2576
R8416 two_stage_opamp_dummy_magic_14_0.VD4.n7 two_stage_opamp_dummy_magic_14_0.VD4.t35 11.2576
R8417 two_stage_opamp_dummy_magic_14_0.VD4.n5 two_stage_opamp_dummy_magic_14_0.VD4.t36 11.2576
R8418 two_stage_opamp_dummy_magic_14_0.VD4.n5 two_stage_opamp_dummy_magic_14_0.VD4.t37 11.2576
R8419 two_stage_opamp_dummy_magic_14_0.VD4.n3 two_stage_opamp_dummy_magic_14_0.VD4.t28 11.2576
R8420 two_stage_opamp_dummy_magic_14_0.VD4.n3 two_stage_opamp_dummy_magic_14_0.VD4.t30 11.2576
R8421 two_stage_opamp_dummy_magic_14_0.VD4.n1 two_stage_opamp_dummy_magic_14_0.VD4.t33 11.2576
R8422 two_stage_opamp_dummy_magic_14_0.VD4.n1 two_stage_opamp_dummy_magic_14_0.VD4.t31 11.2576
R8423 two_stage_opamp_dummy_magic_14_0.VD4.n0 two_stage_opamp_dummy_magic_14_0.VD4.t34 11.2576
R8424 two_stage_opamp_dummy_magic_14_0.VD4.n0 two_stage_opamp_dummy_magic_14_0.VD4.t27 11.2576
R8425 two_stage_opamp_dummy_magic_14_0.VD4.n11 two_stage_opamp_dummy_magic_14_0.VD4.t15 11.2576
R8426 two_stage_opamp_dummy_magic_14_0.VD4.n11 two_stage_opamp_dummy_magic_14_0.VD4.t19 11.2576
R8427 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n14 9.14336
R8428 two_stage_opamp_dummy_magic_14_0.VD4.n56 two_stage_opamp_dummy_magic_14_0.VD4.n55 9.14336
R8429 two_stage_opamp_dummy_magic_14_0.VD4.n53 two_stage_opamp_dummy_magic_14_0.VD4.n50 9.14336
R8430 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n29 9.14336
R8431 two_stage_opamp_dummy_magic_14_0.VD4.n34 two_stage_opamp_dummy_magic_14_0.VD4.n31 9.14336
R8432 two_stage_opamp_dummy_magic_14_0.VD4.n39 two_stage_opamp_dummy_magic_14_0.VD4.n36 9.14336
R8433 two_stage_opamp_dummy_magic_14_0.VD4.n63 two_stage_opamp_dummy_magic_14_0.VD4.n10 8.2505
R8434 two_stage_opamp_dummy_magic_14_0.VD4.n63 two_stage_opamp_dummy_magic_14_0.VD4.n62 5.8755
R8435 two_stage_opamp_dummy_magic_14_0.VD4.n48 two_stage_opamp_dummy_magic_14_0.VD4.n14 4.53698
R8436 two_stage_opamp_dummy_magic_14_0.VD4.n55 two_stage_opamp_dummy_magic_14_0.VD4.n54 4.53698
R8437 two_stage_opamp_dummy_magic_14_0.VD4.n50 two_stage_opamp_dummy_magic_14_0.VD4.n49 4.53698
R8438 two_stage_opamp_dummy_magic_14_0.VD4.n56 two_stage_opamp_dummy_magic_14_0.VD4.n48 4.53698
R8439 two_stage_opamp_dummy_magic_14_0.VD4.n54 two_stage_opamp_dummy_magic_14_0.VD4.n53 4.53698
R8440 two_stage_opamp_dummy_magic_14_0.VD4.n30 two_stage_opamp_dummy_magic_14_0.VD4.n29 4.53698
R8441 two_stage_opamp_dummy_magic_14_0.VD4.n35 two_stage_opamp_dummy_magic_14_0.VD4.n34 4.53698
R8442 two_stage_opamp_dummy_magic_14_0.VD4.n40 two_stage_opamp_dummy_magic_14_0.VD4.n39 4.53698
R8443 two_stage_opamp_dummy_magic_14_0.VD4.n31 two_stage_opamp_dummy_magic_14_0.VD4.n30 4.53698
R8444 two_stage_opamp_dummy_magic_14_0.VD4.n36 two_stage_opamp_dummy_magic_14_0.VD4.n35 4.53698
R8445 two_stage_opamp_dummy_magic_14_0.VD4.n4 two_stage_opamp_dummy_magic_14_0.VD4.n2 0.6255
R8446 two_stage_opamp_dummy_magic_14_0.VD4.n6 two_stage_opamp_dummy_magic_14_0.VD4.n4 0.6255
R8447 two_stage_opamp_dummy_magic_14_0.VD4.n8 two_stage_opamp_dummy_magic_14_0.VD4.n6 0.6255
R8448 two_stage_opamp_dummy_magic_14_0.VD4.n10 two_stage_opamp_dummy_magic_14_0.VD4.n8 0.6255
R8449 two_stage_opamp_dummy_magic_14_0.VD4.n62 two_stage_opamp_dummy_magic_14_0.VD4.n12 0.6255
R8450 two_stage_opamp_dummy_magic_14_0.VD4.n27 two_stage_opamp_dummy_magic_14_0.VD4.n25 0.6255
R8451 two_stage_opamp_dummy_magic_14_0.VD4.n25 two_stage_opamp_dummy_magic_14_0.VD4.n23 0.6255
R8452 two_stage_opamp_dummy_magic_14_0.VD4.n23 two_stage_opamp_dummy_magic_14_0.VD4.n21 0.6255
R8453 two_stage_opamp_dummy_magic_14_0.VD4.n21 two_stage_opamp_dummy_magic_14_0.VD4.n12 0.6255
R8454 two_stage_opamp_dummy_magic_14_0.VD4 two_stage_opamp_dummy_magic_14_0.VD4.n63 0.063
R8455 VIN+.n9 VIN+.t7 490.572
R8456 VIN+.n4 VIN+.t4 449.868
R8457 VIN+.n0 VIN+.t8 449.868
R8458 VIN+.n4 VIN+.t10 273.134
R8459 VIN+.n5 VIN+.t1 273.134
R8460 VIN+.n6 VIN+.t6 273.134
R8461 VIN+.n7 VIN+.t0 273.134
R8462 VIN+.n3 VIN+.t5 273.134
R8463 VIN+.n2 VIN+.t3 273.134
R8464 VIN+.n1 VIN+.t9 273.134
R8465 VIN+.n0 VIN+.t2 273.134
R8466 VIN+.n7 VIN+.n6 176.733
R8467 VIN+.n6 VIN+.n5 176.733
R8468 VIN+.n5 VIN+.n4 176.733
R8469 VIN+.n1 VIN+.n0 176.733
R8470 VIN+.n2 VIN+.n1 176.733
R8471 VIN+.n3 VIN+.n2 176.733
R8472 VIN+.n9 VIN+.n8 165.8
R8473 VIN+.n8 VIN+.n7 56.2338
R8474 VIN+.n8 VIN+.n3 56.2338
R8475 VIN+ VIN+.n9 2.14112
R8476 bgr_7_0.START_UP.n4 bgr_7_0.START_UP.t6 238.322
R8477 bgr_7_0.START_UP.n4 bgr_7_0.START_UP.t7 238.322
R8478 bgr_7_0.START_UP.n3 bgr_7_0.START_UP.n1 175.56
R8479 bgr_7_0.START_UP.n3 bgr_7_0.START_UP.n2 168.936
R8480 bgr_7_0.START_UP.n5 bgr_7_0.START_UP.n4 166.925
R8481 bgr_7_0.START_UP.n0 bgr_7_0.START_UP.t1 130.001
R8482 bgr_7_0.START_UP.n0 bgr_7_0.START_UP.t0 81.7074
R8483 bgr_7_0.START_UP bgr_7_0.START_UP.n0 36.9489
R8484 bgr_7_0.START_UP bgr_7_0.START_UP.n5 13.4693
R8485 bgr_7_0.START_UP.n1 bgr_7_0.START_UP.t2 13.1338
R8486 bgr_7_0.START_UP.n1 bgr_7_0.START_UP.t4 13.1338
R8487 bgr_7_0.START_UP.n2 bgr_7_0.START_UP.t3 13.1338
R8488 bgr_7_0.START_UP.n2 bgr_7_0.START_UP.t5 13.1338
R8489 bgr_7_0.START_UP.n5 bgr_7_0.START_UP.n3 4.21925
R8490 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 144.827
R8491 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 134.577
R8492 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 118.986
R8493 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 100.6
R8494 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 100.038
R8495 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 100.038
R8496 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 100.038
R8497 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 100.038
R8498 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 37.4067
R8499 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 33.705
R8500 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 24.0005
R8501 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 24.0005
R8502 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 24.0005
R8503 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 24.0005
R8504 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 8.0005
R8505 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 8.0005
R8506 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 8.0005
R8507 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 8.0005
R8508 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 8.0005
R8509 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 8.0005
R8510 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 8.0005
R8511 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 8.0005
R8512 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 8.0005
R8513 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 8.0005
R8514 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 5.6255
R8515 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 0.563
R8516 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 0.563
R8517 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 0.563
R8518 bgr_7_0.V_CMFB_S4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 0.047375
R8519 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 365.07
R8520 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_p.t1 15.7605
R8521 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_p.t0 15.7605
R8522 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_p.t3 15.7605
R8523 two_stage_opamp_dummy_magic_14_0.V_err_p.t2 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 15.7605
R8524 two_stage_opamp_dummy_magic_14_0.V_p_mir.n2 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 112.686
R8525 two_stage_opamp_dummy_magic_14_0.V_p_mir.n2 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 106.394
R8526 two_stage_opamp_dummy_magic_14_0.V_p_mir.n3 two_stage_opamp_dummy_magic_14_0.V_p_mir.n2 96.9586
R8527 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 two_stage_opamp_dummy_magic_14_0.V_p_mir.t0 16.0005
R8528 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 two_stage_opamp_dummy_magic_14_0.V_p_mir.t1 16.0005
R8529 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 two_stage_opamp_dummy_magic_14_0.V_p_mir.t2 9.6005
R8530 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 two_stage_opamp_dummy_magic_14_0.V_p_mir.t5 9.6005
R8531 two_stage_opamp_dummy_magic_14_0.V_p_mir.n3 two_stage_opamp_dummy_magic_14_0.V_p_mir.t4 9.6005
R8532 two_stage_opamp_dummy_magic_14_0.V_p_mir.t3 two_stage_opamp_dummy_magic_14_0.V_p_mir.n3 9.6005
R8533 a_5980_2720.t0 a_5980_2720.t1 169.905
R8534 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t2 652.076
R8535 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t6 652.076
R8536 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 585
R8537 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 585
R8538 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 290.233
R8539 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 290.233
R8540 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 290.233
R8541 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 290.233
R8542 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 290.233
R8543 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 290.233
R8544 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 242.903
R8545 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 242.903
R8546 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 238.367
R8547 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 185
R8548 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 185
R8549 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 185
R8550 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 185
R8551 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 185
R8552 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 185
R8553 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 185
R8554 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 185
R8555 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 185
R8556 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 185
R8557 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 185
R8558 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 185
R8559 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 185
R8560 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 170.513
R8561 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 170.513
R8562 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 169.694
R8563 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 155.303
R8564 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 150
R8565 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 150
R8566 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 150
R8567 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 150
R8568 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 150
R8569 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 150
R8570 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 146.155
R8571 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 146.155
R8572 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 65.8183
R8573 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 65.8183
R8574 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 65.8183
R8575 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 65.8183
R8576 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 65.8183
R8577 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 65.8183
R8578 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 53.3664
R8579 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 53.3664
R8580 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 53.3664
R8581 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 53.3664
R8582 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 53.3664
R8583 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 53.3664
R8584 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 53.3664
R8585 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 53.3664
R8586 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 53.3664
R8587 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 22.8576
R8588 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 22.8576
R8589 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 14.4255
R8590 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 14.0505
R8591 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t1 11.2576
R8592 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t4 11.2576
R8593 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t10 11.2576
R8594 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t9 11.2576
R8595 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t8 11.2576
R8596 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 11.2576
R8597 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 9.14336
R8598 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 9.14336
R8599 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 9.14336
R8600 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 9.14336
R8601 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 9.14336
R8602 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 9.14336
R8603 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 4.53698
R8604 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 4.53698
R8605 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 4.53698
R8606 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 4.53698
R8607 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 4.53698
R8608 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 4.53698
R8609 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 4.53698
R8610 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 4.53698
R8611 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 4.53698
R8612 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 4.53698
R8613 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 4.5005
R8614 a_14010_2720.t0 a_14010_2720.t1 169.905
R8615 bgr_7_0.START_UP_NFET1 bgr_7_0.START_UP_NFET1.t0 141.653
R8616 a_12530_23988.t0 a_12530_23988.t1 178.133
R8617 two_stage_opamp_dummy_magic_14_0.V_tot.n2 two_stage_opamp_dummy_magic_14_0.V_tot.t5 648.28
R8618 two_stage_opamp_dummy_magic_14_0.V_tot.n1 two_stage_opamp_dummy_magic_14_0.V_tot.t4 648.28
R8619 two_stage_opamp_dummy_magic_14_0.V_tot.n0 two_stage_opamp_dummy_magic_14_0.V_tot.t2 116.546
R8620 two_stage_opamp_dummy_magic_14_0.V_tot.n3 two_stage_opamp_dummy_magic_14_0.V_tot.t3 116.546
R8621 two_stage_opamp_dummy_magic_14_0.V_tot.n0 two_stage_opamp_dummy_magic_14_0.V_tot.t1 107.328
R8622 two_stage_opamp_dummy_magic_14_0.V_tot.t0 two_stage_opamp_dummy_magic_14_0.V_tot.n3 107.328
R8623 two_stage_opamp_dummy_magic_14_0.V_tot.n3 two_stage_opamp_dummy_magic_14_0.V_tot.n2 35.3494
R8624 two_stage_opamp_dummy_magic_14_0.V_tot.n1 two_stage_opamp_dummy_magic_14_0.V_tot.n0 35.3494
R8625 two_stage_opamp_dummy_magic_14_0.V_tot.n2 two_stage_opamp_dummy_magic_14_0.V_tot.n1 1.563
R8626 a_7580_22380.t0 a_7580_22380.t1 178.133
R8627 a_14330_5524.t0 a_14330_5524.t1 262.248
R8628 a_6810_23838.t0 a_6810_23838.t1 178.133
R8629 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R8630 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R8631 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R8632 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R8633 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R8634 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R8635 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R8636 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R8637 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8638 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R8639 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R8640 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R8641 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R8642 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R8643 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R8644 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R8645 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R8646 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R8647 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R8648 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R8649 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R8650 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8651 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R8652 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R8653 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R8654 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8655 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R8656 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R8657 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R8658 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R8659 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R8660 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R8661 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8662 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R8663 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R8664 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R8665 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R8666 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R8667 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R8668 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R8669 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R8670 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R8671 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R8672 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R8673 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R8674 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R8675 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R8676 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R8677 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R8678 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R8679 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R8680 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R8681 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R8682 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8683 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8684 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8685 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8686 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8687 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8688 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8689 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R8690 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8691 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8692 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8693 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8694 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R8695 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R8696 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8697 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8698 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8699 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8700 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8701 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8702 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8703 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8704 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8705 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8706 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8707 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R8708 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R8709 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R8710 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8711 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8712 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8713 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R8714 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8715 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8716 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8717 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R8718 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8719 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8720 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8721 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8722 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8723 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8724 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8725 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8726 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8727 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8728 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8729 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8730 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R8731 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R8732 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8733 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8734 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8735 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8736 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R8737 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R8738 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R8739 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R8740 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R8741 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R8742 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R8743 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R8744 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R8745 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R8746 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R8747 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R8748 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R8749 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R8750 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R8751 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R8752 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R8753 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R8754 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R8755 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R8756 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8757 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R8758 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R8759 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R8760 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R8761 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R8762 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R8763 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R8764 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R8765 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R8766 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R8767 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R8768 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R8769 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R8770 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8771 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R8772 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R8773 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R8774 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R8775 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R8776 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R8777 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R8778 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R8779 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R8780 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R8781 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R8782 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R8783 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R8784 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R8785 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R8786 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R8787 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R8788 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8789 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R8790 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R8791 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R8792 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R8793 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R8794 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R8795 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R8796 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R8797 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R8798 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R8799 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R8800 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R8801 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R8802 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R8803 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R8804 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8805 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R8806 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R8807 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8808 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R8809 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R8810 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R8811 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R8812 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R8813 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R8814 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R8815 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R8816 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8817 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R8818 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R8819 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8820 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R8821 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8822 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8823 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R8824 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R8825 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R8826 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R8827 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R8828 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R8829 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R8830 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R8831 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R8832 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R8833 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R8834 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R8835 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R8836 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R8837 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8838 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R8839 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R8840 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R8841 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8842 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R8843 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8844 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R8845 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8846 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8847 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8848 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R8849 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8850 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R8851 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R8852 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R8853 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R8854 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R8855 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R8856 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R8857 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R8858 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R8859 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8860 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R8861 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8862 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8863 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R8864 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8865 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8866 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R8867 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R8868 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8869 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8870 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8871 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8872 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R8873 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8874 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8875 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R8876 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R8877 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R8878 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R8879 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R8880 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R8881 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R8882 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8883 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R8884 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8885 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8886 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8887 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R8888 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R8889 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R8890 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8891 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R8892 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8893 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8894 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8895 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8896 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R8897 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8898 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8899 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R8900 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R8901 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R8902 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R8903 a_12410_22380.t0 a_12410_22380.t1 178.133
R8904 a_13060_22630.t0 a_13060_22630.t1 178.133
R8905 a_5420_5524.t0 a_5420_5524.t1 262.248
R8906 a_14450_5524.t0 a_14450_5524.t1 169.905
R8907 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 692.967
R8908 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 two_stage_opamp_dummy_magic_14_0.Vb2_2.t3 652.076
R8909 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 652.076
R8910 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 587.407
R8911 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 587.407
R8912 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 585
R8913 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 585
R8914 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 585
R8915 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 585
R8916 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8917 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8918 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8919 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 246.25
R8920 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 246.25
R8921 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 243.698
R8922 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 242.903
R8923 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 238.367
R8924 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 185
R8925 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 185
R8926 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 185
R8927 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 185
R8928 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 185
R8929 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 185
R8930 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 185
R8931 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 185
R8932 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 185
R8933 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 185
R8934 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 185
R8935 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 185
R8936 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 185
R8937 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.t4 170.513
R8938 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.t7 170.513
R8939 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 155.304
R8940 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 150
R8941 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 150
R8942 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 150
R8943 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 150
R8944 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 150
R8945 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 150
R8946 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 two_stage_opamp_dummy_magic_14_0.Vb2_2.t4 146.155
R8947 two_stage_opamp_dummy_magic_14_0.Vb2_2.t7 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 146.155
R8948 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 65.8183
R8949 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 65.8183
R8950 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 65.8183
R8951 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 65.8183
R8952 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 65.8183
R8953 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 65.8183
R8954 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 53.3664
R8955 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 53.3664
R8956 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 53.3664
R8957 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 53.3664
R8958 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 53.3664
R8959 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 53.3664
R8960 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 53.3664
R8961 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 53.3664
R8962 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 53.3664
R8963 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 22.8576
R8964 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 22.8576
R8965 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 two_stage_opamp_dummy_magic_14_0.Vb2_2.t9 21.8894
R8966 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 two_stage_opamp_dummy_magic_14_0.Vb2_2.t2 21.8894
R8967 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 14.4255
R8968 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 14.0505
R8969 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 two_stage_opamp_dummy_magic_14_0.Vb2_2.t8 11.2576
R8970 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 11.2576
R8971 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 two_stage_opamp_dummy_magic_14_0.Vb2_2.t1 11.2576
R8972 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 9.14336
R8973 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 9.14336
R8974 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 9.14336
R8975 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 9.14336
R8976 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 9.14336
R8977 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 9.14336
R8978 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 9.14336
R8979 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 5.33286
R8980 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 4.53698
R8981 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 4.53698
R8982 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 4.53698
R8983 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 4.53698
R8984 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 4.53698
R8985 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 4.5005
R8986 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 3.75335
R8987 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 3.75335
R8988 a_5540_5524.t0 a_5540_5524.t1 169.905
R8989 a_13180_23838.t0 a_13180_23838.t1 178.133
C0 bgr_7_0.NFET_GATE_10uA bgr_7_0.START_UP_NFET1 0.351171f
C1 bgr_7_0.V_TOP bgr_7_0.PFET_GATE_10uA 0.211901f
C2 bgr_7_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.Vb2 0.538734f
C3 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.V_err_gate 2.05055f
C4 bgr_7_0.1st_Vout_1 m2_10730_16580# 0.075543f
C5 two_stage_opamp_dummy_magic_14_0.V_err_gate VOUT- 0.038574f
C6 bgr_7_0.START_UP_NFET1 bgr_7_0.START_UP 0.145663f
C7 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_7_0.START_UP 0.08188f
C8 bgr_7_0.NFET_GATE_10uA bgr_7_0.PFET_GATE_10uA 0.011067f
C9 li_11260_5990# VIN- 0.024834f
C10 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter m1_10050_19490# 0.013969f
C11 two_stage_opamp_dummy_magic_14_0.V_err_gate bgr_7_0.PFET_GATE_10uA 0.091127f
C12 two_stage_opamp_dummy_magic_14_0.cap_res_X VOUT+ 0.037134f
C13 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.Vb2 0.615806f
C14 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref VOUT+ 0.039491f
C15 two_stage_opamp_dummy_magic_14_0.cap_res_X VOUT- 51.0191f
C16 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01158f
C17 m1_4880_3600# m2_4880_3600# 0.016063f
C18 two_stage_opamp_dummy_magic_14_0.VD4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.044674f
C19 bgr_7_0.V_TOP VDDA 13.2423f
C20 two_stage_opamp_dummy_magic_14_0.V_err_mir_p VDDA 0.671453f
C21 bgr_7_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 1.67069f
C22 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_7_0.1st_Vout_1 0.042752f
C23 two_stage_opamp_dummy_magic_14_0.VD2 VIN+ 1.00068f
C24 bgr_7_0.NFET_GATE_10uA VDDA 0.214521f
C25 two_stage_opamp_dummy_magic_14_0.V_err_gate VDDA 2.16767f
C26 bgr_7_0.START_UP VDDA 1.09224f
C27 bgr_7_0.V_TOP bgr_7_0.NFET_GATE_10uA 0.049214f
C28 two_stage_opamp_dummy_magic_14_0.Vb2 m1_10050_19490# 0.08176f
C29 bgr_7_0.V_TOP two_stage_opamp_dummy_magic_14_0.V_err_gate 0.08195f
C30 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_gate 0.429395f
C31 li_8860_5990# VIN+ 0.024834f
C32 two_stage_opamp_dummy_magic_14_0.cap_res_X VDDA 0.455327f
C33 bgr_7_0.V_TOP bgr_7_0.START_UP 0.792764f
C34 bgr_7_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_err_gate 3.51904f
C35 two_stage_opamp_dummy_magic_14_0.VD2 VDDA 0.020765f
C36 VOUT+ VOUT- 0.397591f
C37 two_stage_opamp_dummy_magic_14_0.VD4 VOUT+ 0.030624f
C38 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref VDDA 2.78293f
C39 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C40 bgr_7_0.NFET_GATE_10uA bgr_7_0.START_UP 1.64125f
C41 bgr_7_0.PFET_GATE_10uA m2_9370_16580# 0.012f
C42 two_stage_opamp_dummy_magic_14_0.Vb2 VOUT- 0.058721f
C43 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.VD4 1.23588f
C44 bgr_7_0.1st_Vout_1 VDDA 0.896465f
C45 bgr_7_0.START_UP_NFET1 bgr_7_0.PFET_GATE_10uA 0.0108f
C46 bgr_7_0.V_TOP two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.583702f
C47 bgr_7_0.V_TOP bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C48 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.047306f
C49 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.V_err_gate 0.33348f
C50 bgr_7_0.V_TOP bgr_7_0.1st_Vout_1 2.47405f
C51 bgr_7_0.V_TOP m2_10730_16580# 0.012f
C52 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.804289f
C53 bgr_7_0.START_UP two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 1.36583f
C54 bgr_7_0.NFET_GATE_10uA bgr_7_0.1st_Vout_1 0.03875f
C55 two_stage_opamp_dummy_magic_14_0.V_err_gate bgr_7_0.1st_Vout_1 0.041119f
C56 VDDA VOUT+ 5.85678f
C57 bgr_7_0.START_UP bgr_7_0.1st_Vout_1 0.04354f
C58 bgr_7_0.START_UP_NFET1 VDDA 0.167059f
C59 two_stage_opamp_dummy_magic_14_0.Vb2 VDDA 1.45884f
C60 VIN+ VIN- 0.102537f
C61 VDDA VOUT- 5.85978f
C62 two_stage_opamp_dummy_magic_14_0.VD4 VDDA 4.49131f
C63 two_stage_opamp_dummy_magic_14_0.V_err_gate m1_10050_19490# 0.091711f
C64 bgr_7_0.PFET_GATE_10uA VDDA 8.31389f
C65 bgr_7_0.V_TOP two_stage_opamp_dummy_magic_14_0.Vb2 0.936691f
C66 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.VD4 0.0195f
C67 two_stage_opamp_dummy_magic_14_0.VD2 li_8860_5990# 0.07273f
C68 VIN- GNDA 1.63494f
C69 VIN+ GNDA 1.64352f
C70 VOUT- GNDA 15.731145f
C71 VOUT+ GNDA 15.764891f
C72 VDDA GNDA 0.122563p
C73 m2_4880_3600# GNDA 0.05269f $ **FLOATING
C74 m2_10730_16580# GNDA 0.0105f $ **FLOATING
C75 m2_9370_16580# GNDA 0.010002f $ **FLOATING
C76 m1_4880_3600# GNDA 0.059696f $ **FLOATING
C77 m1_10050_19490# GNDA 0.259273f $ **FLOATING
C78 li_11260_5990# GNDA 0.01959f $ **FLOATING
C79 li_8860_5990# GNDA 0.01959f $ **FLOATING
C80 two_stage_opamp_dummy_magic_14_0.cap_res_X GNDA 32.97403f
C81 two_stage_opamp_dummy_magic_14_0.VD2 GNDA 2.16451f
C82 two_stage_opamp_dummy_magic_14_0.V_err_mir_p GNDA 0.098428f
C83 bgr_7_0.1st_Vout_1 GNDA 7.823503f
C84 bgr_7_0.START_UP GNDA 5.877477f
C85 bgr_7_0.START_UP_NFET1 GNDA 4.29564f
C86 two_stage_opamp_dummy_magic_14_0.V_err_gate GNDA 9.02901f
C87 two_stage_opamp_dummy_magic_14_0.Vb2 GNDA 7.399733f
C88 bgr_7_0.NFET_GATE_10uA GNDA 7.21715f
C89 bgr_7_0.V_TOP GNDA 9.961141f
C90 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8955f
C91 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref GNDA 7.1992f
C92 bgr_7_0.PFET_GATE_10uA GNDA 6.316023f
C93 two_stage_opamp_dummy_magic_14_0.VD4 GNDA 4.986378f
C94 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 GNDA 0.020756f
C95 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 GNDA 0.020756f
C96 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 GNDA 0.075443f
C97 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 GNDA 0.020756f
C98 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 GNDA 0.020756f
C99 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 GNDA 0.062693f
C100 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 GNDA 1.2228f
C101 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 GNDA 0.255002f
C102 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 GNDA 0.062269f
C103 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 GNDA 0.062269f
C104 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 GNDA 0.259745f
C105 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 GNDA 0.062269f
C106 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 GNDA 0.062269f
C107 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 GNDA 0.258789f
C108 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 GNDA 0.3553f
C109 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 GNDA 0.062269f
C110 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 GNDA 0.062269f
C111 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 GNDA 0.258789f
C112 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 GNDA 0.185392f
C113 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 GNDA 0.062269f
C114 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 GNDA 0.062269f
C115 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 GNDA 0.258789f
C116 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 GNDA 0.185392f
C117 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 GNDA 0.062269f
C118 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 GNDA 0.062269f
C119 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 GNDA 0.258789f
C120 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 GNDA 0.257209f
C121 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 GNDA 1.47144f
C122 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 GNDA 1.81834f
C123 bgr_7_0.V_CMFB_S4 GNDA 0.010378f
C124 bgr_7_0.START_UP.t0 GNDA 1.06745f
C125 bgr_7_0.START_UP.t1 GNDA 0.02806f
C126 bgr_7_0.START_UP.n0 GNDA 0.714928f
C127 bgr_7_0.START_UP.t2 GNDA 0.026778f
C128 bgr_7_0.START_UP.t4 GNDA 0.026778f
C129 bgr_7_0.START_UP.n1 GNDA 0.097147f
C130 bgr_7_0.START_UP.t3 GNDA 0.026778f
C131 bgr_7_0.START_UP.t5 GNDA 0.026778f
C132 bgr_7_0.START_UP.n2 GNDA 0.08937f
C133 bgr_7_0.START_UP.n3 GNDA 0.462855f
C134 bgr_7_0.START_UP.t7 GNDA 0.010062f
C135 bgr_7_0.START_UP.t6 GNDA 0.010062f
C136 bgr_7_0.START_UP.n4 GNDA 0.028407f
C137 bgr_7_0.START_UP.n5 GNDA 0.260836f
C138 two_stage_opamp_dummy_magic_14_0.VD4.t34 GNDA 0.03131f
C139 two_stage_opamp_dummy_magic_14_0.VD4.t27 GNDA 0.03131f
C140 two_stage_opamp_dummy_magic_14_0.VD4.n0 GNDA 0.109961f
C141 two_stage_opamp_dummy_magic_14_0.VD4.t33 GNDA 0.03131f
C142 two_stage_opamp_dummy_magic_14_0.VD4.t31 GNDA 0.03131f
C143 two_stage_opamp_dummy_magic_14_0.VD4.n1 GNDA 0.109583f
C144 two_stage_opamp_dummy_magic_14_0.VD4.n2 GNDA 0.204478f
C145 two_stage_opamp_dummy_magic_14_0.VD4.t28 GNDA 0.03131f
C146 two_stage_opamp_dummy_magic_14_0.VD4.t30 GNDA 0.03131f
C147 two_stage_opamp_dummy_magic_14_0.VD4.n3 GNDA 0.109583f
C148 two_stage_opamp_dummy_magic_14_0.VD4.n4 GNDA 0.106006f
C149 two_stage_opamp_dummy_magic_14_0.VD4.t36 GNDA 0.03131f
C150 two_stage_opamp_dummy_magic_14_0.VD4.t37 GNDA 0.03131f
C151 two_stage_opamp_dummy_magic_14_0.VD4.n5 GNDA 0.109583f
C152 two_stage_opamp_dummy_magic_14_0.VD4.n6 GNDA 0.106006f
C153 two_stage_opamp_dummy_magic_14_0.VD4.t32 GNDA 0.03131f
C154 two_stage_opamp_dummy_magic_14_0.VD4.t35 GNDA 0.03131f
C155 two_stage_opamp_dummy_magic_14_0.VD4.n7 GNDA 0.109583f
C156 two_stage_opamp_dummy_magic_14_0.VD4.n8 GNDA 0.106006f
C157 two_stage_opamp_dummy_magic_14_0.VD4.t26 GNDA 0.03131f
C158 two_stage_opamp_dummy_magic_14_0.VD4.t29 GNDA 0.03131f
C159 two_stage_opamp_dummy_magic_14_0.VD4.n9 GNDA 0.109583f
C160 two_stage_opamp_dummy_magic_14_0.VD4.n10 GNDA 0.15577f
C161 two_stage_opamp_dummy_magic_14_0.VD4.t15 GNDA 0.03131f
C162 two_stage_opamp_dummy_magic_14_0.VD4.t19 GNDA 0.03131f
C163 two_stage_opamp_dummy_magic_14_0.VD4.n11 GNDA 0.108502f
C164 two_stage_opamp_dummy_magic_14_0.VD4.n12 GNDA 0.106192f
C165 two_stage_opamp_dummy_magic_14_0.VD4.t22 GNDA 0.03131f
C166 two_stage_opamp_dummy_magic_14_0.VD4.n13 GNDA 0.093929f
C167 two_stage_opamp_dummy_magic_14_0.VD4.n14 GNDA 0.03131f
C168 two_stage_opamp_dummy_magic_14_0.VD4.n15 GNDA 0.017891f
C169 two_stage_opamp_dummy_magic_14_0.VD4.n18 GNDA 0.014487f
C170 two_stage_opamp_dummy_magic_14_0.VD4.n19 GNDA 0.017891f
C171 two_stage_opamp_dummy_magic_14_0.VD4.t23 GNDA 0.054896f
C172 two_stage_opamp_dummy_magic_14_0.VD4.t5 GNDA 0.03131f
C173 two_stage_opamp_dummy_magic_14_0.VD4.t9 GNDA 0.03131f
C174 two_stage_opamp_dummy_magic_14_0.VD4.n20 GNDA 0.108502f
C175 two_stage_opamp_dummy_magic_14_0.VD4.n21 GNDA 0.106192f
C176 two_stage_opamp_dummy_magic_14_0.VD4.t1 GNDA 0.03131f
C177 two_stage_opamp_dummy_magic_14_0.VD4.t3 GNDA 0.03131f
C178 two_stage_opamp_dummy_magic_14_0.VD4.n22 GNDA 0.108502f
C179 two_stage_opamp_dummy_magic_14_0.VD4.n23 GNDA 0.106192f
C180 two_stage_opamp_dummy_magic_14_0.VD4.t13 GNDA 0.03131f
C181 two_stage_opamp_dummy_magic_14_0.VD4.t17 GNDA 0.03131f
C182 two_stage_opamp_dummy_magic_14_0.VD4.n24 GNDA 0.108502f
C183 two_stage_opamp_dummy_magic_14_0.VD4.n25 GNDA 0.106192f
C184 two_stage_opamp_dummy_magic_14_0.VD4.t11 GNDA 0.03131f
C185 two_stage_opamp_dummy_magic_14_0.VD4.t7 GNDA 0.03131f
C186 two_stage_opamp_dummy_magic_14_0.VD4.n26 GNDA 0.108502f
C187 two_stage_opamp_dummy_magic_14_0.VD4.n27 GNDA 0.135959f
C188 two_stage_opamp_dummy_magic_14_0.VD4.n28 GNDA 0.046623f
C189 two_stage_opamp_dummy_magic_14_0.VD4.n29 GNDA 0.03131f
C190 two_stage_opamp_dummy_magic_14_0.VD4.n31 GNDA 0.03131f
C191 two_stage_opamp_dummy_magic_14_0.VD4.n32 GNDA 0.017891f
C192 two_stage_opamp_dummy_magic_14_0.VD4.n33 GNDA 0.017891f
C193 two_stage_opamp_dummy_magic_14_0.VD4.n34 GNDA 0.03131f
C194 two_stage_opamp_dummy_magic_14_0.VD4.n36 GNDA 0.03131f
C195 two_stage_opamp_dummy_magic_14_0.VD4.n37 GNDA 0.017891f
C196 two_stage_opamp_dummy_magic_14_0.VD4.n38 GNDA 0.017891f
C197 two_stage_opamp_dummy_magic_14_0.VD4.n39 GNDA 0.03131f
C198 two_stage_opamp_dummy_magic_14_0.VD4.n40 GNDA 0.031583f
C199 two_stage_opamp_dummy_magic_14_0.VD4.t25 GNDA 0.03131f
C200 two_stage_opamp_dummy_magic_14_0.VD4.n41 GNDA 0.093929f
C201 two_stage_opamp_dummy_magic_14_0.VD4.n42 GNDA 0.030183f
C202 two_stage_opamp_dummy_magic_14_0.VD4.n43 GNDA 0.017891f
C203 two_stage_opamp_dummy_magic_14_0.VD4.n44 GNDA 0.261659f
C204 two_stage_opamp_dummy_magic_14_0.VD4.t24 GNDA 0.226771f
C205 two_stage_opamp_dummy_magic_14_0.VD4.t10 GNDA 0.209327f
C206 two_stage_opamp_dummy_magic_14_0.VD4.t6 GNDA 0.209327f
C207 two_stage_opamp_dummy_magic_14_0.VD4.t12 GNDA 0.209327f
C208 two_stage_opamp_dummy_magic_14_0.VD4.t16 GNDA 0.209327f
C209 two_stage_opamp_dummy_magic_14_0.VD4.t0 GNDA 0.209327f
C210 two_stage_opamp_dummy_magic_14_0.VD4.t2 GNDA 0.209327f
C211 two_stage_opamp_dummy_magic_14_0.VD4.t4 GNDA 0.209327f
C212 two_stage_opamp_dummy_magic_14_0.VD4.t8 GNDA 0.209327f
C213 two_stage_opamp_dummy_magic_14_0.VD4.t14 GNDA 0.209327f
C214 two_stage_opamp_dummy_magic_14_0.VD4.t18 GNDA 0.209327f
C215 two_stage_opamp_dummy_magic_14_0.VD4.t21 GNDA 0.226771f
C216 two_stage_opamp_dummy_magic_14_0.VD4.n46 GNDA 0.014487f
C217 two_stage_opamp_dummy_magic_14_0.VD4.n47 GNDA 0.017891f
C218 two_stage_opamp_dummy_magic_14_0.VD4.n49 GNDA 0.031583f
C219 two_stage_opamp_dummy_magic_14_0.VD4.n50 GNDA 0.03131f
C220 two_stage_opamp_dummy_magic_14_0.VD4.n51 GNDA 0.017891f
C221 two_stage_opamp_dummy_magic_14_0.VD4.n52 GNDA 0.017891f
C222 two_stage_opamp_dummy_magic_14_0.VD4.n53 GNDA 0.03131f
C223 two_stage_opamp_dummy_magic_14_0.VD4.n55 GNDA 0.03131f
C224 two_stage_opamp_dummy_magic_14_0.VD4.n56 GNDA 0.03131f
C225 two_stage_opamp_dummy_magic_14_0.VD4.n57 GNDA 0.017891f
C226 two_stage_opamp_dummy_magic_14_0.VD4.n58 GNDA 0.261659f
C227 two_stage_opamp_dummy_magic_14_0.VD4.n59 GNDA 0.013886f
C228 two_stage_opamp_dummy_magic_14_0.VD4.n60 GNDA 0.034188f
C229 two_stage_opamp_dummy_magic_14_0.VD4.t20 GNDA 0.054896f
C230 two_stage_opamp_dummy_magic_14_0.VD4.n61 GNDA 0.045275f
C231 two_stage_opamp_dummy_magic_14_0.VD4.n62 GNDA 0.073673f
C232 two_stage_opamp_dummy_magic_14_0.VD4.n63 GNDA 0.091958f
C233 bgr_7_0.Vin-.n0 GNDA 0.069747f
C234 bgr_7_0.Vin-.n1 GNDA 0.078367f
C235 bgr_7_0.Vin-.n2 GNDA 0.113033f
C236 bgr_7_0.Vin-.t2 GNDA 0.261601f
C237 bgr_7_0.Vin-.t6 GNDA 0.027101f
C238 bgr_7_0.Vin-.t4 GNDA 0.027101f
C239 bgr_7_0.Vin-.n3 GNDA 0.094346f
C240 bgr_7_0.Vin-.t3 GNDA 0.027101f
C241 bgr_7_0.Vin-.t5 GNDA 0.027101f
C242 bgr_7_0.Vin-.n4 GNDA 0.090091f
C243 bgr_7_0.Vin-.n5 GNDA 0.386489f
C244 bgr_7_0.Vin-.n6 GNDA 0.027681f
C245 bgr_7_0.Vin-.n7 GNDA 0.366254f
C246 bgr_7_0.Vin-.t12 GNDA 0.022346f
C247 bgr_7_0.Vin-.n8 GNDA 0.026209f
C248 bgr_7_0.Vin-.n9 GNDA 0.021455f
C249 bgr_7_0.Vin-.n10 GNDA 0.021455f
C250 bgr_7_0.Vin-.n11 GNDA 0.036491f
C251 bgr_7_0.Vin-.n12 GNDA 0.497932f
C252 bgr_7_0.Vin-.t7 GNDA 0.117924f
C253 bgr_7_0.Vin-.n13 GNDA 0.65583f
C254 bgr_7_0.Vin-.n14 GNDA 1.073f
C255 bgr_7_0.Vin-.n15 GNDA 0.471409f
C256 bgr_7_0.Vin-.n16 GNDA 0.07053f
C257 bgr_7_0.Vin-.n17 GNDA 0.119504f
C258 bgr_7_0.Vin-.n18 GNDA 0.069875f
C259 bgr_7_0.Vin-.n19 GNDA 0.138215f
C260 bgr_7_0.Vin-.n20 GNDA 0.138215f
C261 bgr_7_0.Vin-.n21 GNDA -0.269519f
C262 bgr_7_0.Vin-.n22 GNDA 0.445457f
C263 bgr_7_0.Vin-.n23 GNDA 0.213551f
C264 bgr_7_0.Vin-.n24 GNDA 0.403461f
C265 bgr_7_0.Vin-.n25 GNDA 0.0384f
C266 bgr_7_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.040751f
C267 bgr_7_0.V_mir2.t7 GNDA 0.019293f
C268 bgr_7_0.V_mir2.n0 GNDA 0.025223f
C269 bgr_7_0.V_mir2.t14 GNDA 0.041163f
C270 bgr_7_0.V_mir2.n1 GNDA 0.027381f
C271 bgr_7_0.V_mir2.n2 GNDA 0.451535f
C272 bgr_7_0.V_mir2.n3 GNDA 0.146338f
C273 bgr_7_0.V_mir2.t4 GNDA 0.023151f
C274 bgr_7_0.V_mir2.t17 GNDA 0.023151f
C275 bgr_7_0.V_mir2.t20 GNDA 0.037369f
C276 bgr_7_0.V_mir2.n4 GNDA 0.041731f
C277 bgr_7_0.V_mir2.n5 GNDA 0.028507f
C278 bgr_7_0.V_mir2.t0 GNDA 0.02939f
C279 bgr_7_0.V_mir2.n6 GNDA 0.044354f
C280 bgr_7_0.V_mir2.t5 GNDA 0.019293f
C281 bgr_7_0.V_mir2.t1 GNDA 0.019293f
C282 bgr_7_0.V_mir2.n7 GNDA 0.044166f
C283 bgr_7_0.V_mir2.n8 GNDA 0.109943f
C284 bgr_7_0.V_mir2.t2 GNDA 0.023151f
C285 bgr_7_0.V_mir2.t18 GNDA 0.023151f
C286 bgr_7_0.V_mir2.t22 GNDA 0.037369f
C287 bgr_7_0.V_mir2.n9 GNDA 0.041731f
C288 bgr_7_0.V_mir2.n10 GNDA 0.028507f
C289 bgr_7_0.V_mir2.t8 GNDA 0.02939f
C290 bgr_7_0.V_mir2.n11 GNDA 0.044354f
C291 bgr_7_0.V_mir2.t3 GNDA 0.019293f
C292 bgr_7_0.V_mir2.t9 GNDA 0.019293f
C293 bgr_7_0.V_mir2.n12 GNDA 0.044166f
C294 bgr_7_0.V_mir2.n13 GNDA 0.111042f
C295 bgr_7_0.V_mir2.n14 GNDA 0.381359f
C296 bgr_7_0.V_mir2.n15 GNDA 0.051125f
C297 bgr_7_0.V_mir2.t6 GNDA 0.023151f
C298 bgr_7_0.V_mir2.t19 GNDA 0.023151f
C299 bgr_7_0.V_mir2.t21 GNDA 0.037369f
C300 bgr_7_0.V_mir2.n16 GNDA 0.041731f
C301 bgr_7_0.V_mir2.n17 GNDA 0.028507f
C302 bgr_7_0.V_mir2.t10 GNDA 0.02939f
C303 bgr_7_0.V_mir2.n18 GNDA 0.044354f
C304 bgr_7_0.V_mir2.n19 GNDA 0.085095f
C305 bgr_7_0.V_mir2.n20 GNDA 0.044166f
C306 bgr_7_0.V_mir2.t11 GNDA 0.019293f
C307 bgr_7_0.cap_res1.t12 GNDA 0.331712f
C308 bgr_7_0.cap_res1.t19 GNDA 0.349187f
C309 bgr_7_0.cap_res1.t16 GNDA 0.350452f
C310 bgr_7_0.cap_res1.t5 GNDA 0.331712f
C311 bgr_7_0.cap_res1.t15 GNDA 0.349187f
C312 bgr_7_0.cap_res1.t9 GNDA 0.350452f
C313 bgr_7_0.cap_res1.t11 GNDA 0.331712f
C314 bgr_7_0.cap_res1.t18 GNDA 0.349187f
C315 bgr_7_0.cap_res1.t14 GNDA 0.350452f
C316 bgr_7_0.cap_res1.t4 GNDA 0.331712f
C317 bgr_7_0.cap_res1.t13 GNDA 0.349187f
C318 bgr_7_0.cap_res1.t7 GNDA 0.350452f
C319 bgr_7_0.cap_res1.t20 GNDA 0.331712f
C320 bgr_7_0.cap_res1.t6 GNDA 0.349187f
C321 bgr_7_0.cap_res1.t1 GNDA 0.350452f
C322 bgr_7_0.cap_res1.n0 GNDA 0.23406f
C323 bgr_7_0.cap_res1.t17 GNDA 0.186395f
C324 bgr_7_0.cap_res1.n1 GNDA 0.253961f
C325 bgr_7_0.cap_res1.t2 GNDA 0.186395f
C326 bgr_7_0.cap_res1.n2 GNDA 0.253961f
C327 bgr_7_0.cap_res1.t8 GNDA 0.186395f
C328 bgr_7_0.cap_res1.n3 GNDA 0.253961f
C329 bgr_7_0.cap_res1.t3 GNDA 0.186395f
C330 bgr_7_0.cap_res1.n4 GNDA 0.253961f
C331 bgr_7_0.cap_res1.t10 GNDA 0.363549f
C332 bgr_7_0.cap_res1.t0 GNDA 0.08421f
C333 bgr_7_0.PFET_GATE_10uA.t23 GNDA 0.020962f
C334 bgr_7_0.PFET_GATE_10uA.t17 GNDA 0.031035f
C335 bgr_7_0.PFET_GATE_10uA.n0 GNDA 0.066714f
C336 bgr_7_0.PFET_GATE_10uA.t24 GNDA 0.020962f
C337 bgr_7_0.PFET_GATE_10uA.t19 GNDA 0.030987f
C338 bgr_7_0.PFET_GATE_10uA.n1 GNDA 0.034144f
C339 bgr_7_0.PFET_GATE_10uA.t13 GNDA 0.020962f
C340 bgr_7_0.PFET_GATE_10uA.t20 GNDA 0.030987f
C341 bgr_7_0.PFET_GATE_10uA.n2 GNDA 0.034144f
C342 bgr_7_0.PFET_GATE_10uA.n3 GNDA 0.031856f
C343 bgr_7_0.PFET_GATE_10uA.n4 GNDA 0.659441f
C344 bgr_7_0.PFET_GATE_10uA.t16 GNDA 0.020962f
C345 bgr_7_0.PFET_GATE_10uA.t11 GNDA 0.030987f
C346 bgr_7_0.PFET_GATE_10uA.n5 GNDA 0.034144f
C347 bgr_7_0.PFET_GATE_10uA.t22 GNDA 0.020962f
C348 bgr_7_0.PFET_GATE_10uA.t12 GNDA 0.030987f
C349 bgr_7_0.PFET_GATE_10uA.n6 GNDA 0.034144f
C350 bgr_7_0.PFET_GATE_10uA.n7 GNDA 0.034254f
C351 bgr_7_0.PFET_GATE_10uA.t9 GNDA 0.314052f
C352 bgr_7_0.PFET_GATE_10uA.t0 GNDA 0.021499f
C353 bgr_7_0.PFET_GATE_10uA.t7 GNDA 0.021499f
C354 bgr_7_0.PFET_GATE_10uA.n8 GNDA 0.05495f
C355 bgr_7_0.PFET_GATE_10uA.t2 GNDA 0.021499f
C356 bgr_7_0.PFET_GATE_10uA.t4 GNDA 0.021499f
C357 bgr_7_0.PFET_GATE_10uA.n9 GNDA 0.05353f
C358 bgr_7_0.PFET_GATE_10uA.n10 GNDA 0.523597f
C359 bgr_7_0.PFET_GATE_10uA.t3 GNDA 0.021499f
C360 bgr_7_0.PFET_GATE_10uA.t5 GNDA 0.021499f
C361 bgr_7_0.PFET_GATE_10uA.n11 GNDA 0.05353f
C362 bgr_7_0.PFET_GATE_10uA.n12 GNDA 0.296907f
C363 bgr_7_0.PFET_GATE_10uA.n13 GNDA 0.606116f
C364 bgr_7_0.PFET_GATE_10uA.t8 GNDA 0.021499f
C365 bgr_7_0.PFET_GATE_10uA.t1 GNDA 0.021499f
C366 bgr_7_0.PFET_GATE_10uA.n14 GNDA 0.051852f
C367 bgr_7_0.PFET_GATE_10uA.n15 GNDA 0.276809f
C368 bgr_7_0.PFET_GATE_10uA.t6 GNDA 0.466209f
C369 bgr_7_0.PFET_GATE_10uA.t18 GNDA 0.062934f
C370 bgr_7_0.PFET_GATE_10uA.n16 GNDA 1.92661f
C371 bgr_7_0.PFET_GATE_10uA.n17 GNDA 0.778649f
C372 bgr_7_0.PFET_GATE_10uA.n18 GNDA 0.763078f
C373 bgr_7_0.PFET_GATE_10uA.t10 GNDA 0.045148f
C374 bgr_7_0.PFET_GATE_10uA.t21 GNDA 0.045148f
C375 bgr_7_0.PFET_GATE_10uA.t15 GNDA 0.054823f
C376 bgr_7_0.PFET_GATE_10uA.n19 GNDA 0.054823f
C377 bgr_7_0.PFET_GATE_10uA.n20 GNDA 0.03127f
C378 bgr_7_0.PFET_GATE_10uA.t14 GNDA 0.048555f
C379 bgr_7_0.PFET_GATE_10uA.n21 GNDA 0.053269f
C380 two_stage_opamp_dummy_magic_14_0.Vb1.t0 GNDA 0.011829f
C381 two_stage_opamp_dummy_magic_14_0.Vb1.t9 GNDA 0.011829f
C382 two_stage_opamp_dummy_magic_14_0.Vb1.n0 GNDA 0.041331f
C383 two_stage_opamp_dummy_magic_14_0.Vb1.t18 GNDA 0.011794f
C384 two_stage_opamp_dummy_magic_14_0.Vb1.n1 GNDA 0.012824f
C385 two_stage_opamp_dummy_magic_14_0.Vb1.t12 GNDA 0.011794f
C386 two_stage_opamp_dummy_magic_14_0.Vb1.n5 GNDA 0.012824f
C387 two_stage_opamp_dummy_magic_14_0.Vb1.n9 GNDA 0.013132f
C388 two_stage_opamp_dummy_magic_14_0.Vb1.t26 GNDA 0.011794f
C389 two_stage_opamp_dummy_magic_14_0.Vb1.n10 GNDA 0.012824f
C390 two_stage_opamp_dummy_magic_14_0.Vb1.t20 GNDA 0.011794f
C391 two_stage_opamp_dummy_magic_14_0.Vb1.n14 GNDA 0.012824f
C392 two_stage_opamp_dummy_magic_14_0.Vb1.n19 GNDA 0.194378f
C393 two_stage_opamp_dummy_magic_14_0.Vb1.t15 GNDA 0.265569f
C394 two_stage_opamp_dummy_magic_14_0.Vb1.n20 GNDA 0.031226f
C395 two_stage_opamp_dummy_magic_14_0.Vb1.n21 GNDA 0.20356f
C396 two_stage_opamp_dummy_magic_14_0.Vb1.t5 GNDA 0.011794f
C397 two_stage_opamp_dummy_magic_14_0.Vb1.n22 GNDA 0.012126f
C398 two_stage_opamp_dummy_magic_14_0.Vb1.t7 GNDA 0.011794f
C399 two_stage_opamp_dummy_magic_14_0.Vb1.n23 GNDA 0.012126f
C400 two_stage_opamp_dummy_magic_14_0.Vb1.n25 GNDA 0.027604f
C401 two_stage_opamp_dummy_magic_14_0.Vb1.n26 GNDA 0.029894f
C402 two_stage_opamp_dummy_magic_14_0.Vb1.n27 GNDA 0.02412f
C403 two_stage_opamp_dummy_magic_14_0.Vb1.n28 GNDA 0.031226f
C404 two_stage_opamp_dummy_magic_14_0.Vb1.n29 GNDA 0.223662f
C405 two_stage_opamp_dummy_magic_14_0.Vb1.n30 GNDA 0.449117f
C406 bgr_7_0.VB1_CUR_BIAS GNDA 0.461318f
C407 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 GNDA 0.026703f
C408 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 GNDA 0.026703f
C409 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 GNDA 0.406043f
C410 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 GNDA 0.066758f
C411 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 GNDA 0.066758f
C412 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 GNDA 0.204527f
C413 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 GNDA 0.074546f
C414 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 GNDA 0.074546f
C415 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 GNDA 0.111974f
C416 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 GNDA 0.413267f
C417 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 GNDA 0.066758f
C418 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 GNDA 0.066758f
C419 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 GNDA 0.203641f
C420 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 GNDA 0.316207f
C421 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 GNDA 0.074546f
C422 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 GNDA 0.074546f
C423 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 GNDA 0.111974f
C424 bgr_7_0.V_CUR_REF_REG.n0 GNDA 0.05674f
C425 bgr_7_0.V_CUR_REF_REG.t5 GNDA 0.011381f
C426 bgr_7_0.V_CUR_REF_REG.n1 GNDA 0.024409f
C427 bgr_7_0.V_CUR_REF_REG.n2 GNDA 0.018995f
C428 bgr_7_0.V_CUR_REF_REG.n3 GNDA 0.019251f
C429 bgr_7_0.V_CUR_REF_REG.n4 GNDA 0.035481f
C430 bgr_7_0.V_CUR_REF_REG.n5 GNDA 1.74641f
C431 bgr_7_0.V_CUR_REF_REG.t0 GNDA 0.244345f
C432 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 GNDA 0.016424f
C433 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 GNDA 0.016424f
C434 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 GNDA 0.041188f
C435 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 GNDA 0.016424f
C436 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 GNDA 0.016424f
C437 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 GNDA 0.040971f
C438 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 GNDA 0.364219f
C439 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 GNDA 0.016424f
C440 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 GNDA 0.016424f
C441 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 GNDA 0.032849f
C442 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 GNDA 0.061063f
C443 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 GNDA 0.206842f
C444 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 GNDA 0.032849f
C445 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 GNDA 0.032849f
C446 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 GNDA 0.097616f
C447 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 GNDA 0.032849f
C448 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 GNDA 0.032849f
C449 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 GNDA 0.097184f
C450 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 GNDA 0.332426f
C451 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 GNDA 0.032849f
C452 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 GNDA 0.032849f
C453 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 GNDA 0.097184f
C454 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 GNDA 0.172178f
C455 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 GNDA 0.032849f
C456 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 GNDA 0.032849f
C457 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 GNDA 0.097184f
C458 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 GNDA 0.172178f
C459 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 GNDA 0.032849f
C460 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 GNDA 0.032849f
C461 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 GNDA 0.097184f
C462 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 GNDA 0.240026f
C463 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 GNDA 1.40468f
C464 bgr_7_0.V_CMFB_S3 GNDA 0.917995f
C465 two_stage_opamp_dummy_magic_14_0.Y.t10 GNDA 0.031899f
C466 two_stage_opamp_dummy_magic_14_0.Y.t7 GNDA 0.031899f
C467 two_stage_opamp_dummy_magic_14_0.Y.n0 GNDA 0.112032f
C468 two_stage_opamp_dummy_magic_14_0.Y.t8 GNDA 0.031899f
C469 two_stage_opamp_dummy_magic_14_0.Y.t6 GNDA 0.031899f
C470 two_stage_opamp_dummy_magic_14_0.Y.n1 GNDA 0.111647f
C471 two_stage_opamp_dummy_magic_14_0.Y.n2 GNDA 0.20833f
C472 two_stage_opamp_dummy_magic_14_0.Y.t1 GNDA 0.031899f
C473 two_stage_opamp_dummy_magic_14_0.Y.t4 GNDA 0.031899f
C474 two_stage_opamp_dummy_magic_14_0.Y.n3 GNDA 0.111647f
C475 two_stage_opamp_dummy_magic_14_0.Y.n4 GNDA 0.108003f
C476 two_stage_opamp_dummy_magic_14_0.Y.t9 GNDA 0.031899f
C477 two_stage_opamp_dummy_magic_14_0.Y.t3 GNDA 0.031899f
C478 two_stage_opamp_dummy_magic_14_0.Y.n5 GNDA 0.111647f
C479 two_stage_opamp_dummy_magic_14_0.Y.n6 GNDA 0.108003f
C480 two_stage_opamp_dummy_magic_14_0.Y.t0 GNDA 0.031899f
C481 two_stage_opamp_dummy_magic_14_0.Y.t5 GNDA 0.031899f
C482 two_stage_opamp_dummy_magic_14_0.Y.n7 GNDA 0.111647f
C483 two_stage_opamp_dummy_magic_14_0.Y.n8 GNDA 0.127209f
C484 two_stage_opamp_dummy_magic_14_0.Y.t2 GNDA 0.031899f
C485 two_stage_opamp_dummy_magic_14_0.Y.t20 GNDA 0.031899f
C486 two_stage_opamp_dummy_magic_14_0.Y.n9 GNDA 0.109409f
C487 two_stage_opamp_dummy_magic_14_0.Y.n10 GNDA 0.179923f
C488 two_stage_opamp_dummy_magic_14_0.Y.t23 GNDA 0.013671f
C489 two_stage_opamp_dummy_magic_14_0.Y.t24 GNDA 0.013671f
C490 two_stage_opamp_dummy_magic_14_0.Y.n11 GNDA 0.050047f
C491 two_stage_opamp_dummy_magic_14_0.Y.t14 GNDA 0.013671f
C492 two_stage_opamp_dummy_magic_14_0.Y.t11 GNDA 0.013671f
C493 two_stage_opamp_dummy_magic_14_0.Y.n12 GNDA 0.049628f
C494 two_stage_opamp_dummy_magic_14_0.Y.n13 GNDA 0.181951f
C495 two_stage_opamp_dummy_magic_14_0.Y.t12 GNDA 0.013671f
C496 two_stage_opamp_dummy_magic_14_0.Y.t19 GNDA 0.013671f
C497 two_stage_opamp_dummy_magic_14_0.Y.n14 GNDA 0.049628f
C498 two_stage_opamp_dummy_magic_14_0.Y.n15 GNDA 0.094375f
C499 two_stage_opamp_dummy_magic_14_0.Y.t15 GNDA 0.013671f
C500 two_stage_opamp_dummy_magic_14_0.Y.t18 GNDA 0.013671f
C501 two_stage_opamp_dummy_magic_14_0.Y.n16 GNDA 0.049628f
C502 two_stage_opamp_dummy_magic_14_0.Y.n17 GNDA 0.094375f
C503 two_stage_opamp_dummy_magic_14_0.Y.t13 GNDA 0.013671f
C504 two_stage_opamp_dummy_magic_14_0.Y.t21 GNDA 0.013671f
C505 two_stage_opamp_dummy_magic_14_0.Y.n18 GNDA 0.049628f
C506 two_stage_opamp_dummy_magic_14_0.Y.n19 GNDA 0.094375f
C507 two_stage_opamp_dummy_magic_14_0.Y.t17 GNDA 0.013671f
C508 two_stage_opamp_dummy_magic_14_0.Y.t22 GNDA 0.013671f
C509 two_stage_opamp_dummy_magic_14_0.Y.n20 GNDA 0.049628f
C510 two_stage_opamp_dummy_magic_14_0.Y.n21 GNDA 0.141822f
C511 two_stage_opamp_dummy_magic_14_0.Y.n22 GNDA 0.195875f
C512 two_stage_opamp_dummy_magic_14_0.Y.t38 GNDA 0.01914f
C513 two_stage_opamp_dummy_magic_14_0.Y.t34 GNDA 0.01914f
C514 two_stage_opamp_dummy_magic_14_0.Y.t39 GNDA 0.01914f
C515 two_stage_opamp_dummy_magic_14_0.Y.t53 GNDA 0.023241f
C516 two_stage_opamp_dummy_magic_14_0.Y.n23 GNDA 0.023241f
C517 two_stage_opamp_dummy_magic_14_0.Y.n24 GNDA 0.015038f
C518 two_stage_opamp_dummy_magic_14_0.Y.n25 GNDA 0.013264f
C519 two_stage_opamp_dummy_magic_14_0.Y.t25 GNDA 0.01914f
C520 two_stage_opamp_dummy_magic_14_0.Y.t42 GNDA 0.01914f
C521 two_stage_opamp_dummy_magic_14_0.Y.t29 GNDA 0.01914f
C522 two_stage_opamp_dummy_magic_14_0.Y.t45 GNDA 0.01914f
C523 two_stage_opamp_dummy_magic_14_0.Y.t32 GNDA 0.01914f
C524 two_stage_opamp_dummy_magic_14_0.Y.t48 GNDA 0.023241f
C525 two_stage_opamp_dummy_magic_14_0.Y.n26 GNDA 0.023241f
C526 two_stage_opamp_dummy_magic_14_0.Y.n27 GNDA 0.015038f
C527 two_stage_opamp_dummy_magic_14_0.Y.n28 GNDA 0.015038f
C528 two_stage_opamp_dummy_magic_14_0.Y.n29 GNDA 0.015038f
C529 two_stage_opamp_dummy_magic_14_0.Y.n30 GNDA 0.013264f
C530 two_stage_opamp_dummy_magic_14_0.Y.n31 GNDA 0.013782f
C531 two_stage_opamp_dummy_magic_14_0.Y.t27 GNDA 0.029393f
C532 two_stage_opamp_dummy_magic_14_0.Y.t50 GNDA 0.029393f
C533 two_stage_opamp_dummy_magic_14_0.Y.t28 GNDA 0.029393f
C534 two_stage_opamp_dummy_magic_14_0.Y.t41 GNDA 0.033415f
C535 two_stage_opamp_dummy_magic_14_0.Y.n32 GNDA 0.030156f
C536 two_stage_opamp_dummy_magic_14_0.Y.n33 GNDA 0.018456f
C537 two_stage_opamp_dummy_magic_14_0.Y.n34 GNDA 0.016682f
C538 two_stage_opamp_dummy_magic_14_0.Y.t44 GNDA 0.029393f
C539 two_stage_opamp_dummy_magic_14_0.Y.t31 GNDA 0.029393f
C540 two_stage_opamp_dummy_magic_14_0.Y.t47 GNDA 0.029393f
C541 two_stage_opamp_dummy_magic_14_0.Y.t33 GNDA 0.029393f
C542 two_stage_opamp_dummy_magic_14_0.Y.t49 GNDA 0.029393f
C543 two_stage_opamp_dummy_magic_14_0.Y.t35 GNDA 0.033415f
C544 two_stage_opamp_dummy_magic_14_0.Y.n35 GNDA 0.030156f
C545 two_stage_opamp_dummy_magic_14_0.Y.n36 GNDA 0.018456f
C546 two_stage_opamp_dummy_magic_14_0.Y.n37 GNDA 0.018456f
C547 two_stage_opamp_dummy_magic_14_0.Y.n38 GNDA 0.018456f
C548 two_stage_opamp_dummy_magic_14_0.Y.n39 GNDA 0.016682f
C549 two_stage_opamp_dummy_magic_14_0.Y.n40 GNDA 0.013782f
C550 two_stage_opamp_dummy_magic_14_0.Y.n41 GNDA 0.12298f
C551 two_stage_opamp_dummy_magic_14_0.Y.n42 GNDA 0.15804f
C552 two_stage_opamp_dummy_magic_14_0.Y.t37 GNDA 0.060153f
C553 two_stage_opamp_dummy_magic_14_0.Y.t51 GNDA 0.060153f
C554 two_stage_opamp_dummy_magic_14_0.Y.t46 GNDA 0.060153f
C555 two_stage_opamp_dummy_magic_14_0.Y.t52 GNDA 0.060153f
C556 two_stage_opamp_dummy_magic_14_0.Y.t36 GNDA 0.064067f
C557 two_stage_opamp_dummy_magic_14_0.Y.n43 GNDA 0.050771f
C558 two_stage_opamp_dummy_magic_14_0.Y.n44 GNDA 0.028709f
C559 two_stage_opamp_dummy_magic_14_0.Y.n45 GNDA 0.028709f
C560 two_stage_opamp_dummy_magic_14_0.Y.n46 GNDA 0.026942f
C561 two_stage_opamp_dummy_magic_14_0.Y.t54 GNDA 0.060153f
C562 two_stage_opamp_dummy_magic_14_0.Y.t40 GNDA 0.060153f
C563 two_stage_opamp_dummy_magic_14_0.Y.t26 GNDA 0.060153f
C564 two_stage_opamp_dummy_magic_14_0.Y.t43 GNDA 0.060153f
C565 two_stage_opamp_dummy_magic_14_0.Y.t30 GNDA 0.064067f
C566 two_stage_opamp_dummy_magic_14_0.Y.n47 GNDA 0.050771f
C567 two_stage_opamp_dummy_magic_14_0.Y.n48 GNDA 0.028709f
C568 two_stage_opamp_dummy_magic_14_0.Y.n49 GNDA 0.028709f
C569 two_stage_opamp_dummy_magic_14_0.Y.n50 GNDA 0.026942f
C570 two_stage_opamp_dummy_magic_14_0.Y.n51 GNDA 0.016389f
C571 two_stage_opamp_dummy_magic_14_0.Y.n52 GNDA 0.506605f
C572 two_stage_opamp_dummy_magic_14_0.Y.t16 GNDA 0.43926f
C573 two_stage_opamp_dummy_magic_14_0.VD3.t1 GNDA 0.03131f
C574 two_stage_opamp_dummy_magic_14_0.VD3.t9 GNDA 0.03131f
C575 two_stage_opamp_dummy_magic_14_0.VD3.t15 GNDA 0.03131f
C576 two_stage_opamp_dummy_magic_14_0.VD3.n0 GNDA 0.108502f
C577 two_stage_opamp_dummy_magic_14_0.VD3.n1 GNDA 0.106192f
C578 two_stage_opamp_dummy_magic_14_0.VD3.t24 GNDA 0.03131f
C579 two_stage_opamp_dummy_magic_14_0.VD3.n2 GNDA 0.093929f
C580 two_stage_opamp_dummy_magic_14_0.VD3.n3 GNDA 0.03131f
C581 two_stage_opamp_dummy_magic_14_0.VD3.n4 GNDA 0.017891f
C582 two_stage_opamp_dummy_magic_14_0.VD3.n7 GNDA 0.014487f
C583 two_stage_opamp_dummy_magic_14_0.VD3.n8 GNDA 0.017891f
C584 two_stage_opamp_dummy_magic_14_0.VD3.t25 GNDA 0.054896f
C585 two_stage_opamp_dummy_magic_14_0.VD3.t21 GNDA 0.03131f
C586 two_stage_opamp_dummy_magic_14_0.VD3.t36 GNDA 0.03131f
C587 two_stage_opamp_dummy_magic_14_0.VD3.n9 GNDA 0.109961f
C588 two_stage_opamp_dummy_magic_14_0.VD3.t37 GNDA 0.03131f
C589 two_stage_opamp_dummy_magic_14_0.VD3.t29 GNDA 0.03131f
C590 two_stage_opamp_dummy_magic_14_0.VD3.n10 GNDA 0.109583f
C591 two_stage_opamp_dummy_magic_14_0.VD3.n11 GNDA 0.204478f
C592 two_stage_opamp_dummy_magic_14_0.VD3.t32 GNDA 0.03131f
C593 two_stage_opamp_dummy_magic_14_0.VD3.t31 GNDA 0.03131f
C594 two_stage_opamp_dummy_magic_14_0.VD3.n12 GNDA 0.109583f
C595 two_stage_opamp_dummy_magic_14_0.VD3.n13 GNDA 0.106006f
C596 two_stage_opamp_dummy_magic_14_0.VD3.t33 GNDA 0.03131f
C597 two_stage_opamp_dummy_magic_14_0.VD3.t34 GNDA 0.03131f
C598 two_stage_opamp_dummy_magic_14_0.VD3.n14 GNDA 0.109583f
C599 two_stage_opamp_dummy_magic_14_0.VD3.n15 GNDA 0.106006f
C600 two_stage_opamp_dummy_magic_14_0.VD3.t35 GNDA 0.03131f
C601 two_stage_opamp_dummy_magic_14_0.VD3.t30 GNDA 0.03131f
C602 two_stage_opamp_dummy_magic_14_0.VD3.n16 GNDA 0.109583f
C603 two_stage_opamp_dummy_magic_14_0.VD3.n17 GNDA 0.106006f
C604 two_stage_opamp_dummy_magic_14_0.VD3.t28 GNDA 0.03131f
C605 two_stage_opamp_dummy_magic_14_0.VD3.t20 GNDA 0.03131f
C606 two_stage_opamp_dummy_magic_14_0.VD3.n18 GNDA 0.109583f
C607 two_stage_opamp_dummy_magic_14_0.VD3.n19 GNDA 0.195671f
C608 two_stage_opamp_dummy_magic_14_0.VD3.t5 GNDA 0.03131f
C609 two_stage_opamp_dummy_magic_14_0.VD3.t13 GNDA 0.03131f
C610 two_stage_opamp_dummy_magic_14_0.VD3.n20 GNDA 0.108502f
C611 two_stage_opamp_dummy_magic_14_0.VD3.n21 GNDA 0.106192f
C612 two_stage_opamp_dummy_magic_14_0.VD3.n22 GNDA 0.129308f
C613 two_stage_opamp_dummy_magic_14_0.VD3.n23 GNDA 0.045275f
C614 two_stage_opamp_dummy_magic_14_0.VD3.n24 GNDA 0.03131f
C615 two_stage_opamp_dummy_magic_14_0.VD3.n26 GNDA 0.03131f
C616 two_stage_opamp_dummy_magic_14_0.VD3.n27 GNDA 0.017891f
C617 two_stage_opamp_dummy_magic_14_0.VD3.n28 GNDA 0.017891f
C618 two_stage_opamp_dummy_magic_14_0.VD3.n29 GNDA 0.03131f
C619 two_stage_opamp_dummy_magic_14_0.VD3.n31 GNDA 0.03131f
C620 two_stage_opamp_dummy_magic_14_0.VD3.n32 GNDA 0.017891f
C621 two_stage_opamp_dummy_magic_14_0.VD3.n33 GNDA 0.017891f
C622 two_stage_opamp_dummy_magic_14_0.VD3.n34 GNDA 0.03131f
C623 two_stage_opamp_dummy_magic_14_0.VD3.n35 GNDA 0.031583f
C624 two_stage_opamp_dummy_magic_14_0.VD3.t27 GNDA 0.03131f
C625 two_stage_opamp_dummy_magic_14_0.VD3.n36 GNDA 0.093929f
C626 two_stage_opamp_dummy_magic_14_0.VD3.n37 GNDA 0.030183f
C627 two_stage_opamp_dummy_magic_14_0.VD3.n38 GNDA 0.017891f
C628 two_stage_opamp_dummy_magic_14_0.VD3.n39 GNDA 0.261659f
C629 two_stage_opamp_dummy_magic_14_0.VD3.t26 GNDA 0.226771f
C630 two_stage_opamp_dummy_magic_14_0.VD3.t4 GNDA 0.209327f
C631 two_stage_opamp_dummy_magic_14_0.VD3.t12 GNDA 0.209327f
C632 two_stage_opamp_dummy_magic_14_0.VD3.t8 GNDA 0.209327f
C633 two_stage_opamp_dummy_magic_14_0.VD3.t14 GNDA 0.209327f
C634 two_stage_opamp_dummy_magic_14_0.VD3.t18 GNDA 0.209327f
C635 two_stage_opamp_dummy_magic_14_0.VD3.t0 GNDA 0.209327f
C636 two_stage_opamp_dummy_magic_14_0.VD3.t6 GNDA 0.209327f
C637 two_stage_opamp_dummy_magic_14_0.VD3.t2 GNDA 0.209327f
C638 two_stage_opamp_dummy_magic_14_0.VD3.t10 GNDA 0.209327f
C639 two_stage_opamp_dummy_magic_14_0.VD3.t16 GNDA 0.209327f
C640 two_stage_opamp_dummy_magic_14_0.VD3.t23 GNDA 0.226771f
C641 two_stage_opamp_dummy_magic_14_0.VD3.n41 GNDA 0.014487f
C642 two_stage_opamp_dummy_magic_14_0.VD3.n42 GNDA 0.017891f
C643 two_stage_opamp_dummy_magic_14_0.VD3.n44 GNDA 0.031583f
C644 two_stage_opamp_dummy_magic_14_0.VD3.n45 GNDA 0.03131f
C645 two_stage_opamp_dummy_magic_14_0.VD3.n46 GNDA 0.017891f
C646 two_stage_opamp_dummy_magic_14_0.VD3.n47 GNDA 0.017891f
C647 two_stage_opamp_dummy_magic_14_0.VD3.n48 GNDA 0.03131f
C648 two_stage_opamp_dummy_magic_14_0.VD3.n50 GNDA 0.03131f
C649 two_stage_opamp_dummy_magic_14_0.VD3.n51 GNDA 0.03131f
C650 two_stage_opamp_dummy_magic_14_0.VD3.n52 GNDA 0.017891f
C651 two_stage_opamp_dummy_magic_14_0.VD3.n53 GNDA 0.261659f
C652 two_stage_opamp_dummy_magic_14_0.VD3.n54 GNDA 0.013886f
C653 two_stage_opamp_dummy_magic_14_0.VD3.n55 GNDA 0.034188f
C654 two_stage_opamp_dummy_magic_14_0.VD3.t22 GNDA 0.054896f
C655 two_stage_opamp_dummy_magic_14_0.VD3.n56 GNDA 0.046623f
C656 two_stage_opamp_dummy_magic_14_0.VD3.t11 GNDA 0.03131f
C657 two_stage_opamp_dummy_magic_14_0.VD3.t17 GNDA 0.03131f
C658 two_stage_opamp_dummy_magic_14_0.VD3.n57 GNDA 0.108502f
C659 two_stage_opamp_dummy_magic_14_0.VD3.n58 GNDA 0.135959f
C660 two_stage_opamp_dummy_magic_14_0.VD3.t7 GNDA 0.03131f
C661 two_stage_opamp_dummy_magic_14_0.VD3.t3 GNDA 0.03131f
C662 two_stage_opamp_dummy_magic_14_0.VD3.n59 GNDA 0.108502f
C663 two_stage_opamp_dummy_magic_14_0.VD3.n60 GNDA 0.106192f
C664 two_stage_opamp_dummy_magic_14_0.VD3.n61 GNDA 0.106192f
C665 two_stage_opamp_dummy_magic_14_0.VD3.n62 GNDA 0.108502f
C666 two_stage_opamp_dummy_magic_14_0.VD3.t19 GNDA 0.03131f
C667 two_stage_opamp_dummy_magic_14_0.Vb2.t32 GNDA 0.043632f
C668 two_stage_opamp_dummy_magic_14_0.Vb2.t14 GNDA 0.043632f
C669 two_stage_opamp_dummy_magic_14_0.Vb2.t19 GNDA 0.043632f
C670 two_stage_opamp_dummy_magic_14_0.Vb2.t26 GNDA 0.043632f
C671 two_stage_opamp_dummy_magic_14_0.Vb2.t22 GNDA 0.050351f
C672 two_stage_opamp_dummy_magic_14_0.Vb2.n0 GNDA 0.04088f
C673 two_stage_opamp_dummy_magic_14_0.Vb2.n1 GNDA 0.025122f
C674 two_stage_opamp_dummy_magic_14_0.Vb2.n2 GNDA 0.025122f
C675 two_stage_opamp_dummy_magic_14_0.Vb2.n3 GNDA 0.023309f
C676 two_stage_opamp_dummy_magic_14_0.Vb2.t29 GNDA 0.043632f
C677 two_stage_opamp_dummy_magic_14_0.Vb2.t28 GNDA 0.043632f
C678 two_stage_opamp_dummy_magic_14_0.Vb2.t24 GNDA 0.043632f
C679 two_stage_opamp_dummy_magic_14_0.Vb2.t17 GNDA 0.043632f
C680 two_stage_opamp_dummy_magic_14_0.Vb2.t12 GNDA 0.050351f
C681 two_stage_opamp_dummy_magic_14_0.Vb2.n4 GNDA 0.04088f
C682 two_stage_opamp_dummy_magic_14_0.Vb2.n5 GNDA 0.025122f
C683 two_stage_opamp_dummy_magic_14_0.Vb2.n6 GNDA 0.025122f
C684 two_stage_opamp_dummy_magic_14_0.Vb2.n7 GNDA 0.023309f
C685 two_stage_opamp_dummy_magic_14_0.Vb2.n8 GNDA 0.013512f
C686 two_stage_opamp_dummy_magic_14_0.Vb2.t11 GNDA 0.043632f
C687 two_stage_opamp_dummy_magic_14_0.Vb2.t15 GNDA 0.043632f
C688 two_stage_opamp_dummy_magic_14_0.Vb2.t20 GNDA 0.043632f
C689 two_stage_opamp_dummy_magic_14_0.Vb2.t16 GNDA 0.043632f
C690 two_stage_opamp_dummy_magic_14_0.Vb2.t23 GNDA 0.050351f
C691 two_stage_opamp_dummy_magic_14_0.Vb2.n9 GNDA 0.04088f
C692 two_stage_opamp_dummy_magic_14_0.Vb2.n10 GNDA 0.025122f
C693 two_stage_opamp_dummy_magic_14_0.Vb2.n11 GNDA 0.025122f
C694 two_stage_opamp_dummy_magic_14_0.Vb2.n12 GNDA 0.023309f
C695 two_stage_opamp_dummy_magic_14_0.Vb2.t30 GNDA 0.043632f
C696 two_stage_opamp_dummy_magic_14_0.Vb2.t21 GNDA 0.043632f
C697 two_stage_opamp_dummy_magic_14_0.Vb2.t25 GNDA 0.043632f
C698 two_stage_opamp_dummy_magic_14_0.Vb2.t18 GNDA 0.043632f
C699 two_stage_opamp_dummy_magic_14_0.Vb2.t13 GNDA 0.050351f
C700 two_stage_opamp_dummy_magic_14_0.Vb2.n13 GNDA 0.04088f
C701 two_stage_opamp_dummy_magic_14_0.Vb2.n14 GNDA 0.025122f
C702 two_stage_opamp_dummy_magic_14_0.Vb2.n15 GNDA 0.025122f
C703 two_stage_opamp_dummy_magic_14_0.Vb2.n16 GNDA 0.023309f
C704 two_stage_opamp_dummy_magic_14_0.Vb2.n17 GNDA 0.016397f
C705 two_stage_opamp_dummy_magic_14_0.Vb2.n18 GNDA 0.03003f
C706 two_stage_opamp_dummy_magic_14_0.Vb2.n19 GNDA 0.029147f
C707 two_stage_opamp_dummy_magic_14_0.Vb2.n20 GNDA 0.303104f
C708 two_stage_opamp_dummy_magic_14_0.Vb2.n21 GNDA 0.029147f
C709 two_stage_opamp_dummy_magic_14_0.Vb2.n22 GNDA 0.204441f
C710 two_stage_opamp_dummy_magic_14_0.Vb2.n23 GNDA 0.029147f
C711 two_stage_opamp_dummy_magic_14_0.Vb2.n24 GNDA 0.808923f
C712 two_stage_opamp_dummy_magic_14_0.Vb2.t31 GNDA 0.053353f
C713 two_stage_opamp_dummy_magic_14_0.Vb2.n25 GNDA 0.723168f
C714 two_stage_opamp_dummy_magic_14_0.Vb2.t1 GNDA 0.030851f
C715 two_stage_opamp_dummy_magic_14_0.Vb2.t10 GNDA 0.030851f
C716 two_stage_opamp_dummy_magic_14_0.Vb2.n26 GNDA 0.107063f
C717 two_stage_opamp_dummy_magic_14_0.Vb2.t0 GNDA 0.053353f
C718 two_stage_opamp_dummy_magic_14_0.Vb2.n27 GNDA 0.18525f
C719 two_stage_opamp_dummy_magic_14_0.Vb2.t27 GNDA 0.031502f
C720 two_stage_opamp_dummy_magic_14_0.Vb2.n28 GNDA 0.094361f
C721 two_stage_opamp_dummy_magic_14_0.Vb2.n29 GNDA 0.154162f
C722 two_stage_opamp_dummy_magic_14_0.Vb2.n30 GNDA 0.287807f
C723 bgr_7_0.cap_res2.t6 GNDA 0.358376f
C724 bgr_7_0.cap_res2.t12 GNDA 0.359675f
C725 bgr_7_0.cap_res2.t14 GNDA 0.340442f
C726 bgr_7_0.cap_res2.t0 GNDA 0.358376f
C727 bgr_7_0.cap_res2.t5 GNDA 0.359675f
C728 bgr_7_0.cap_res2.t8 GNDA 0.340442f
C729 bgr_7_0.cap_res2.t4 GNDA 0.358376f
C730 bgr_7_0.cap_res2.t10 GNDA 0.359675f
C731 bgr_7_0.cap_res2.t13 GNDA 0.340442f
C732 bgr_7_0.cap_res2.t19 GNDA 0.358376f
C733 bgr_7_0.cap_res2.t3 GNDA 0.359675f
C734 bgr_7_0.cap_res2.t7 GNDA 0.340442f
C735 bgr_7_0.cap_res2.t15 GNDA 0.358376f
C736 bgr_7_0.cap_res2.t18 GNDA 0.359675f
C737 bgr_7_0.cap_res2.t1 GNDA 0.340442f
C738 bgr_7_0.cap_res2.n0 GNDA 0.24022f
C739 bgr_7_0.cap_res2.t2 GNDA 0.1913f
C740 bgr_7_0.cap_res2.n1 GNDA 0.260644f
C741 bgr_7_0.cap_res2.t9 GNDA 0.1913f
C742 bgr_7_0.cap_res2.n2 GNDA 0.260644f
C743 bgr_7_0.cap_res2.t16 GNDA 0.1913f
C744 bgr_7_0.cap_res2.n3 GNDA 0.260644f
C745 bgr_7_0.cap_res2.t11 GNDA 0.1913f
C746 bgr_7_0.cap_res2.n4 GNDA 0.260644f
C747 bgr_7_0.cap_res2.t17 GNDA 0.373116f
C748 bgr_7_0.cap_res2.t20 GNDA 0.086426f
C749 bgr_7_0.1st_Vout_2.n0 GNDA 0.237573f
C750 bgr_7_0.1st_Vout_2.n1 GNDA 0.723004f
C751 bgr_7_0.1st_Vout_2.n2 GNDA 1.43086f
C752 bgr_7_0.1st_Vout_2.n3 GNDA 0.104399f
C753 bgr_7_0.1st_Vout_2.n4 GNDA 1.45767f
C754 bgr_7_0.1st_Vout_2.t33 GNDA 0.017308f
C755 bgr_7_0.1st_Vout_2.n5 GNDA 0.018179f
C756 bgr_7_0.1st_Vout_2.t24 GNDA 0.010986f
C757 bgr_7_0.1st_Vout_2.t13 GNDA 0.010986f
C758 bgr_7_0.1st_Vout_2.n6 GNDA 0.024439f
C759 bgr_7_0.1st_Vout_2.n7 GNDA 0.010417f
C760 bgr_7_0.1st_Vout_2.t10 GNDA 0.015189f
C761 bgr_7_0.1st_Vout_2.n8 GNDA 0.157567f
C762 bgr_7_0.1st_Vout_2.n10 GNDA 0.017425f
C763 bgr_7_0.1st_Vout_2.t27 GNDA 0.010986f
C764 bgr_7_0.1st_Vout_2.t16 GNDA 0.010986f
C765 bgr_7_0.1st_Vout_2.n11 GNDA 0.024439f
C766 bgr_7_0.1st_Vout_2.t28 GNDA 0.288462f
C767 bgr_7_0.1st_Vout_2.t17 GNDA 0.293375f
C768 bgr_7_0.1st_Vout_2.t12 GNDA 0.288462f
C769 bgr_7_0.1st_Vout_2.t32 GNDA 0.288462f
C770 bgr_7_0.1st_Vout_2.t35 GNDA 0.293375f
C771 bgr_7_0.1st_Vout_2.t11 GNDA 0.293375f
C772 bgr_7_0.1st_Vout_2.t31 GNDA 0.288462f
C773 bgr_7_0.1st_Vout_2.t23 GNDA 0.288462f
C774 bgr_7_0.1st_Vout_2.t26 GNDA 0.293375f
C775 bgr_7_0.1st_Vout_2.t30 GNDA 0.293375f
C776 bgr_7_0.1st_Vout_2.t22 GNDA 0.288462f
C777 bgr_7_0.1st_Vout_2.t15 GNDA 0.288462f
C778 bgr_7_0.1st_Vout_2.t19 GNDA 0.293375f
C779 bgr_7_0.1st_Vout_2.t36 GNDA 0.293375f
C780 bgr_7_0.1st_Vout_2.t29 GNDA 0.288462f
C781 bgr_7_0.1st_Vout_2.t21 GNDA 0.288462f
C782 bgr_7_0.1st_Vout_2.t25 GNDA 0.293375f
C783 bgr_7_0.1st_Vout_2.t18 GNDA 0.293375f
C784 bgr_7_0.1st_Vout_2.t14 GNDA 0.288462f
C785 bgr_7_0.1st_Vout_2.t20 GNDA 0.288462f
C786 bgr_7_0.1st_Vout_2.t34 GNDA 0.018845f
C787 bgr_7_0.1st_Vout_2.n12 GNDA 0.018179f
C788 bgr_7_0.1st_Vout_1.n0 GNDA 0.538712f
C789 bgr_7_0.1st_Vout_1.n1 GNDA 0.236313f
C790 bgr_7_0.1st_Vout_1.n2 GNDA 0.973284f
C791 bgr_7_0.1st_Vout_1.n3 GNDA 0.907198f
C792 bgr_7_0.1st_Vout_1.n4 GNDA 0.891647f
C793 bgr_7_0.1st_Vout_1.t11 GNDA 0.358463f
C794 bgr_7_0.1st_Vout_1.t15 GNDA 0.35246f
C795 bgr_7_0.1st_Vout_1.t29 GNDA 0.358463f
C796 bgr_7_0.1st_Vout_1.t35 GNDA 0.35246f
C797 bgr_7_0.1st_Vout_1.t31 GNDA 0.358463f
C798 bgr_7_0.1st_Vout_1.t34 GNDA 0.35246f
C799 bgr_7_0.1st_Vout_1.t20 GNDA 0.358463f
C800 bgr_7_0.1st_Vout_1.t28 GNDA 0.35246f
C801 bgr_7_0.1st_Vout_1.t24 GNDA 0.358463f
C802 bgr_7_0.1st_Vout_1.t27 GNDA 0.35246f
C803 bgr_7_0.1st_Vout_1.t14 GNDA 0.358463f
C804 bgr_7_0.1st_Vout_1.t19 GNDA 0.35246f
C805 bgr_7_0.1st_Vout_1.t30 GNDA 0.358463f
C806 bgr_7_0.1st_Vout_1.t33 GNDA 0.35246f
C807 bgr_7_0.1st_Vout_1.t18 GNDA 0.358463f
C808 bgr_7_0.1st_Vout_1.t26 GNDA 0.35246f
C809 bgr_7_0.1st_Vout_1.t23 GNDA 0.358463f
C810 bgr_7_0.1st_Vout_1.t25 GNDA 0.35246f
C811 bgr_7_0.1st_Vout_1.t17 GNDA 0.35246f
C812 bgr_7_0.1st_Vout_1.t12 GNDA 0.35246f
C813 bgr_7_0.1st_Vout_1.t21 GNDA 0.023025f
C814 bgr_7_0.1st_Vout_1.n5 GNDA 0.715456f
C815 bgr_7_0.1st_Vout_1.n6 GNDA 0.022212f
C816 bgr_7_0.1st_Vout_1.n7 GNDA 0.104674f
C817 bgr_7_0.1st_Vout_1.t36 GNDA 0.013423f
C818 bgr_7_0.1st_Vout_1.t16 GNDA 0.013423f
C819 bgr_7_0.1st_Vout_1.n8 GNDA 0.029862f
C820 bgr_7_0.1st_Vout_1.n9 GNDA 0.082514f
C821 bgr_7_0.1st_Vout_1.t10 GNDA 0.018559f
C822 bgr_7_0.1st_Vout_1.n10 GNDA 0.012728f
C823 bgr_7_0.1st_Vout_1.n11 GNDA 0.192525f
C824 bgr_7_0.1st_Vout_1.n12 GNDA 0.011517f
C825 bgr_7_0.1st_Vout_1.n13 GNDA 0.048842f
C826 bgr_7_0.1st_Vout_1.n14 GNDA 0.021291f
C827 bgr_7_0.1st_Vout_1.n15 GNDA 0.078719f
C828 bgr_7_0.1st_Vout_1.n16 GNDA 0.038771f
C829 bgr_7_0.1st_Vout_1.t32 GNDA 0.013423f
C830 bgr_7_0.1st_Vout_1.t22 GNDA 0.013423f
C831 bgr_7_0.1st_Vout_1.n17 GNDA 0.029862f
C832 bgr_7_0.1st_Vout_1.n18 GNDA 0.082514f
C833 bgr_7_0.1st_Vout_1.n19 GNDA 0.022212f
C834 bgr_7_0.1st_Vout_1.n20 GNDA 0.104674f
C835 bgr_7_0.1st_Vout_1.t13 GNDA 0.021069f
C836 bgr_7_0.V_mir1.t12 GNDA 0.019293f
C837 bgr_7_0.V_mir1.t5 GNDA 0.02939f
C838 bgr_7_0.V_mir1.t9 GNDA 0.023151f
C839 bgr_7_0.V_mir1.t18 GNDA 0.023151f
C840 bgr_7_0.V_mir1.t20 GNDA 0.037369f
C841 bgr_7_0.V_mir1.n0 GNDA 0.041731f
C842 bgr_7_0.V_mir1.n1 GNDA 0.028507f
C843 bgr_7_0.V_mir1.n2 GNDA 0.044354f
C844 bgr_7_0.V_mir1.t6 GNDA 0.019293f
C845 bgr_7_0.V_mir1.t10 GNDA 0.019293f
C846 bgr_7_0.V_mir1.n3 GNDA 0.044166f
C847 bgr_7_0.V_mir1.n4 GNDA 0.109943f
C848 bgr_7_0.V_mir1.n5 GNDA 0.025223f
C849 bgr_7_0.V_mir1.t0 GNDA 0.041163f
C850 bgr_7_0.V_mir1.n6 GNDA 0.027381f
C851 bgr_7_0.V_mir1.n7 GNDA 0.451535f
C852 bgr_7_0.V_mir1.n8 GNDA 0.146338f
C853 bgr_7_0.V_mir1.t7 GNDA 0.02939f
C854 bgr_7_0.V_mir1.t13 GNDA 0.023151f
C855 bgr_7_0.V_mir1.t17 GNDA 0.023151f
C856 bgr_7_0.V_mir1.t21 GNDA 0.037369f
C857 bgr_7_0.V_mir1.n9 GNDA 0.041731f
C858 bgr_7_0.V_mir1.n10 GNDA 0.028507f
C859 bgr_7_0.V_mir1.n11 GNDA 0.044354f
C860 bgr_7_0.V_mir1.t8 GNDA 0.019293f
C861 bgr_7_0.V_mir1.t14 GNDA 0.019293f
C862 bgr_7_0.V_mir1.n12 GNDA 0.044166f
C863 bgr_7_0.V_mir1.n13 GNDA 0.085095f
C864 bgr_7_0.V_mir1.n14 GNDA 0.051125f
C865 bgr_7_0.V_mir1.n15 GNDA 0.381359f
C866 bgr_7_0.V_mir1.t11 GNDA 0.02939f
C867 bgr_7_0.V_mir1.t15 GNDA 0.023151f
C868 bgr_7_0.V_mir1.t22 GNDA 0.023151f
C869 bgr_7_0.V_mir1.t19 GNDA 0.037369f
C870 bgr_7_0.V_mir1.n16 GNDA 0.041731f
C871 bgr_7_0.V_mir1.n17 GNDA 0.028507f
C872 bgr_7_0.V_mir1.n18 GNDA 0.044354f
C873 bgr_7_0.V_mir1.n19 GNDA 0.111042f
C874 bgr_7_0.V_mir1.n20 GNDA 0.044166f
C875 bgr_7_0.V_mir1.t16 GNDA 0.019293f
C876 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 GNDA 0.016424f
C877 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 GNDA 0.016424f
C878 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 GNDA 0.041171f
C879 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 GNDA 0.016424f
C880 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 GNDA 0.016424f
C881 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 GNDA 0.040954f
C882 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 GNDA 0.363992f
C883 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 GNDA 0.016424f
C884 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 GNDA 0.016424f
C885 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 GNDA 0.032849f
C886 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 GNDA 0.061089f
C887 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 GNDA 0.206842f
C888 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 GNDA 0.032849f
C889 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 GNDA 0.032849f
C890 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 GNDA 0.097616f
C891 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 GNDA 0.032849f
C892 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 GNDA 0.032849f
C893 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 GNDA 0.097184f
C894 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 GNDA 0.332426f
C895 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 GNDA 0.032849f
C896 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 GNDA 0.032849f
C897 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 GNDA 0.097184f
C898 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 GNDA 0.172178f
C899 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 GNDA 0.032849f
C900 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 GNDA 0.032849f
C901 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 GNDA 0.097184f
C902 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 GNDA 0.172178f
C903 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 GNDA 0.032849f
C904 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 GNDA 0.032849f
C905 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 GNDA 0.097184f
C906 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 GNDA 0.240026f
C907 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 GNDA 1.40468f
C908 bgr_7_0.V_CMFB_S1 GNDA 0.918231f
C909 bgr_7_0.Vin+.t1 GNDA 0.173951f
C910 bgr_7_0.Vin+.t7 GNDA 0.010696f
C911 bgr_7_0.Vin+.t8 GNDA 0.025367f
C912 bgr_7_0.Vin+.t9 GNDA 0.01649f
C913 bgr_7_0.Vin+.n0 GNDA 0.054406f
C914 bgr_7_0.Vin+.t6 GNDA 0.01649f
C915 bgr_7_0.Vin+.n1 GNDA 0.042338f
C916 bgr_7_0.Vin+.t10 GNDA 0.01649f
C917 bgr_7_0.Vin+.n2 GNDA 0.042909f
C918 bgr_7_0.Vin+.n3 GNDA 0.130793f
C919 bgr_7_0.Vin+.t4 GNDA 0.05348f
C920 bgr_7_0.Vin+.t3 GNDA 0.05348f
C921 bgr_7_0.Vin+.n4 GNDA 0.176679f
C922 bgr_7_0.Vin+.n5 GNDA 1.27851f
C923 bgr_7_0.Vin+.t2 GNDA 0.05348f
C924 bgr_7_0.Vin+.t5 GNDA 0.05348f
C925 bgr_7_0.Vin+.n6 GNDA 0.176679f
C926 bgr_7_0.Vin+.n7 GNDA 1.06525f
C927 bgr_7_0.Vin+.n8 GNDA 1.7265f
C928 bgr_7_0.Vin+.t0 GNDA 0.232527f
C929 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 GNDA 0.067008f
C930 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 GNDA 0.065881f
C931 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 GNDA 0.477431f
C932 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 GNDA 0.307683f
C933 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 GNDA 0.048115f
C934 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 GNDA 0.017992f
C935 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 GNDA 0.056432f
C936 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 GNDA 0.017992f
C937 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 GNDA 0.046195f
C938 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 GNDA 0.017992f
C939 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 GNDA 0.046195f
C940 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 GNDA 0.017992f
C941 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 GNDA 0.080073f
C942 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 GNDA 1.60088f
C943 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 GNDA 0.058352f
C944 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 GNDA 0.058352f
C945 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 GNDA 0.205513f
C946 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 GNDA 0.058352f
C947 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 GNDA 0.058352f
C948 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 GNDA 0.195539f
C949 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 GNDA 0.913816f
C950 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 GNDA 0.058352f
C951 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 GNDA 0.058352f
C952 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 GNDA 0.195539f
C953 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 GNDA 0.653448f
C954 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 GNDA 1.34823f
C955 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 GNDA 0.102986f
C956 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 GNDA 0.279533f
C957 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 GNDA 0.258036f
C958 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 GNDA 0.258036f
C959 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 GNDA 0.306249f
C960 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 GNDA 0.161758f
C961 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 GNDA 0.102403f
C962 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 GNDA 0.099835f
C963 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 GNDA 0.531165f
C964 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 GNDA 0.258036f
C965 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 GNDA 0.258036f
C966 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 GNDA 0.306249f
C967 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 GNDA 0.161758f
C968 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 GNDA 0.102403f
C969 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 GNDA 0.279533f
C970 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 GNDA 0.099835f
C971 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 GNDA 0.531165f
C972 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 GNDA 0.102986f
C973 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 GNDA 0.020231f
C974 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 GNDA 0.020231f
C975 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 GNDA 0.073533f
C976 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 GNDA 0.020231f
C977 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 GNDA 0.020231f
C978 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 GNDA 0.061105f
C979 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 GNDA 1.19184f
C980 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 GNDA 0.248547f
C981 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 GNDA 0.060692f
C982 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 GNDA 0.060692f
C983 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 GNDA 0.253169f
C984 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 GNDA 0.060692f
C985 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 GNDA 0.060692f
C986 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 GNDA 0.252238f
C987 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 GNDA 0.346305f
C988 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 GNDA 0.060692f
C989 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 GNDA 0.060692f
C990 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 GNDA 0.252238f
C991 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 GNDA 0.180699f
C992 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 GNDA 0.060692f
C993 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 GNDA 0.060692f
C994 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 GNDA 0.252238f
C995 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 GNDA 0.180699f
C996 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 GNDA 0.060692f
C997 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 GNDA 0.060692f
C998 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 GNDA 0.252238f
C999 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 GNDA 0.250697f
C1000 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 GNDA 1.43419f
C1001 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 GNDA 1.77231f
C1002 bgr_7_0.V_CMFB_S2 GNDA 0.010115f
C1003 two_stage_opamp_dummy_magic_14_0.X.t5 GNDA 0.031899f
C1004 two_stage_opamp_dummy_magic_14_0.X.t12 GNDA 0.031899f
C1005 two_stage_opamp_dummy_magic_14_0.X.n0 GNDA 0.112032f
C1006 two_stage_opamp_dummy_magic_14_0.X.t23 GNDA 0.031899f
C1007 two_stage_opamp_dummy_magic_14_0.X.t7 GNDA 0.031899f
C1008 two_stage_opamp_dummy_magic_14_0.X.n1 GNDA 0.111647f
C1009 two_stage_opamp_dummy_magic_14_0.X.n2 GNDA 0.20833f
C1010 two_stage_opamp_dummy_magic_14_0.X.t20 GNDA 0.031899f
C1011 two_stage_opamp_dummy_magic_14_0.X.t4 GNDA 0.031899f
C1012 two_stage_opamp_dummy_magic_14_0.X.n3 GNDA 0.111647f
C1013 two_stage_opamp_dummy_magic_14_0.X.n4 GNDA 0.108003f
C1014 two_stage_opamp_dummy_magic_14_0.X.t0 GNDA 0.031899f
C1015 two_stage_opamp_dummy_magic_14_0.X.t22 GNDA 0.031899f
C1016 two_stage_opamp_dummy_magic_14_0.X.n5 GNDA 0.111647f
C1017 two_stage_opamp_dummy_magic_14_0.X.n6 GNDA 0.108003f
C1018 two_stage_opamp_dummy_magic_14_0.X.t21 GNDA 0.031899f
C1019 two_stage_opamp_dummy_magic_14_0.X.t6 GNDA 0.031899f
C1020 two_stage_opamp_dummy_magic_14_0.X.n7 GNDA 0.111647f
C1021 two_stage_opamp_dummy_magic_14_0.X.n8 GNDA 0.127209f
C1022 two_stage_opamp_dummy_magic_14_0.X.t11 GNDA 0.031899f
C1023 two_stage_opamp_dummy_magic_14_0.X.t14 GNDA 0.031899f
C1024 two_stage_opamp_dummy_magic_14_0.X.n9 GNDA 0.109409f
C1025 two_stage_opamp_dummy_magic_14_0.X.n10 GNDA 0.179923f
C1026 two_stage_opamp_dummy_magic_14_0.X.t1 GNDA 0.013671f
C1027 two_stage_opamp_dummy_magic_14_0.X.t17 GNDA 0.013671f
C1028 two_stage_opamp_dummy_magic_14_0.X.n11 GNDA 0.050047f
C1029 two_stage_opamp_dummy_magic_14_0.X.t18 GNDA 0.013671f
C1030 two_stage_opamp_dummy_magic_14_0.X.t10 GNDA 0.013671f
C1031 two_stage_opamp_dummy_magic_14_0.X.n12 GNDA 0.049628f
C1032 two_stage_opamp_dummy_magic_14_0.X.n13 GNDA 0.181951f
C1033 two_stage_opamp_dummy_magic_14_0.X.t8 GNDA 0.013671f
C1034 two_stage_opamp_dummy_magic_14_0.X.t13 GNDA 0.013671f
C1035 two_stage_opamp_dummy_magic_14_0.X.n14 GNDA 0.049628f
C1036 two_stage_opamp_dummy_magic_14_0.X.n15 GNDA 0.094375f
C1037 two_stage_opamp_dummy_magic_14_0.X.t3 GNDA 0.013671f
C1038 two_stage_opamp_dummy_magic_14_0.X.t9 GNDA 0.013671f
C1039 two_stage_opamp_dummy_magic_14_0.X.n16 GNDA 0.049628f
C1040 two_stage_opamp_dummy_magic_14_0.X.n17 GNDA 0.094375f
C1041 two_stage_opamp_dummy_magic_14_0.X.t2 GNDA 0.013671f
C1042 two_stage_opamp_dummy_magic_14_0.X.t19 GNDA 0.013671f
C1043 two_stage_opamp_dummy_magic_14_0.X.n18 GNDA 0.049628f
C1044 two_stage_opamp_dummy_magic_14_0.X.n19 GNDA 0.094375f
C1045 two_stage_opamp_dummy_magic_14_0.X.t16 GNDA 0.013671f
C1046 two_stage_opamp_dummy_magic_14_0.X.t24 GNDA 0.013671f
C1047 two_stage_opamp_dummy_magic_14_0.X.n20 GNDA 0.049628f
C1048 two_stage_opamp_dummy_magic_14_0.X.n21 GNDA 0.141822f
C1049 two_stage_opamp_dummy_magic_14_0.X.n22 GNDA 0.195875f
C1050 two_stage_opamp_dummy_magic_14_0.X.t34 GNDA 0.01914f
C1051 two_stage_opamp_dummy_magic_14_0.X.t49 GNDA 0.01914f
C1052 two_stage_opamp_dummy_magic_14_0.X.t26 GNDA 0.01914f
C1053 two_stage_opamp_dummy_magic_14_0.X.t40 GNDA 0.01914f
C1054 two_stage_opamp_dummy_magic_14_0.X.t53 GNDA 0.01914f
C1055 two_stage_opamp_dummy_magic_14_0.X.t36 GNDA 0.023241f
C1056 two_stage_opamp_dummy_magic_14_0.X.n23 GNDA 0.023241f
C1057 two_stage_opamp_dummy_magic_14_0.X.n24 GNDA 0.015038f
C1058 two_stage_opamp_dummy_magic_14_0.X.n25 GNDA 0.015038f
C1059 two_stage_opamp_dummy_magic_14_0.X.n26 GNDA 0.015038f
C1060 two_stage_opamp_dummy_magic_14_0.X.n27 GNDA 0.013264f
C1061 two_stage_opamp_dummy_magic_14_0.X.t52 GNDA 0.01914f
C1062 two_stage_opamp_dummy_magic_14_0.X.t38 GNDA 0.01914f
C1063 two_stage_opamp_dummy_magic_14_0.X.t45 GNDA 0.01914f
C1064 two_stage_opamp_dummy_magic_14_0.X.t30 GNDA 0.023241f
C1065 two_stage_opamp_dummy_magic_14_0.X.n28 GNDA 0.023241f
C1066 two_stage_opamp_dummy_magic_14_0.X.n29 GNDA 0.015038f
C1067 two_stage_opamp_dummy_magic_14_0.X.n30 GNDA 0.013264f
C1068 two_stage_opamp_dummy_magic_14_0.X.n31 GNDA 0.013782f
C1069 two_stage_opamp_dummy_magic_14_0.X.t54 GNDA 0.029393f
C1070 two_stage_opamp_dummy_magic_14_0.X.t37 GNDA 0.029393f
C1071 two_stage_opamp_dummy_magic_14_0.X.t44 GNDA 0.029393f
C1072 two_stage_opamp_dummy_magic_14_0.X.t29 GNDA 0.029393f
C1073 two_stage_opamp_dummy_magic_14_0.X.t42 GNDA 0.029393f
C1074 two_stage_opamp_dummy_magic_14_0.X.t25 GNDA 0.033415f
C1075 two_stage_opamp_dummy_magic_14_0.X.n32 GNDA 0.030156f
C1076 two_stage_opamp_dummy_magic_14_0.X.n33 GNDA 0.018456f
C1077 two_stage_opamp_dummy_magic_14_0.X.n34 GNDA 0.018456f
C1078 two_stage_opamp_dummy_magic_14_0.X.n35 GNDA 0.018456f
C1079 two_stage_opamp_dummy_magic_14_0.X.n36 GNDA 0.016682f
C1080 two_stage_opamp_dummy_magic_14_0.X.t41 GNDA 0.029393f
C1081 two_stage_opamp_dummy_magic_14_0.X.t27 GNDA 0.029393f
C1082 two_stage_opamp_dummy_magic_14_0.X.t32 GNDA 0.029393f
C1083 two_stage_opamp_dummy_magic_14_0.X.t47 GNDA 0.033415f
C1084 two_stage_opamp_dummy_magic_14_0.X.n37 GNDA 0.030156f
C1085 two_stage_opamp_dummy_magic_14_0.X.n38 GNDA 0.018456f
C1086 two_stage_opamp_dummy_magic_14_0.X.n39 GNDA 0.016682f
C1087 two_stage_opamp_dummy_magic_14_0.X.n40 GNDA 0.013782f
C1088 two_stage_opamp_dummy_magic_14_0.X.n41 GNDA 0.12298f
C1089 two_stage_opamp_dummy_magic_14_0.X.n42 GNDA 0.15804f
C1090 two_stage_opamp_dummy_magic_14_0.X.t31 GNDA 0.060153f
C1091 two_stage_opamp_dummy_magic_14_0.X.t39 GNDA 0.060153f
C1092 two_stage_opamp_dummy_magic_14_0.X.t51 GNDA 0.060153f
C1093 two_stage_opamp_dummy_magic_14_0.X.t35 GNDA 0.060153f
C1094 two_stage_opamp_dummy_magic_14_0.X.t48 GNDA 0.064067f
C1095 two_stage_opamp_dummy_magic_14_0.X.n43 GNDA 0.050771f
C1096 two_stage_opamp_dummy_magic_14_0.X.n44 GNDA 0.028709f
C1097 two_stage_opamp_dummy_magic_14_0.X.n45 GNDA 0.028709f
C1098 two_stage_opamp_dummy_magic_14_0.X.n46 GNDA 0.026942f
C1099 two_stage_opamp_dummy_magic_14_0.X.t46 GNDA 0.060153f
C1100 two_stage_opamp_dummy_magic_14_0.X.t33 GNDA 0.060153f
C1101 two_stage_opamp_dummy_magic_14_0.X.t50 GNDA 0.060153f
C1102 two_stage_opamp_dummy_magic_14_0.X.t28 GNDA 0.060153f
C1103 two_stage_opamp_dummy_magic_14_0.X.t43 GNDA 0.064067f
C1104 two_stage_opamp_dummy_magic_14_0.X.n47 GNDA 0.050771f
C1105 two_stage_opamp_dummy_magic_14_0.X.n48 GNDA 0.028709f
C1106 two_stage_opamp_dummy_magic_14_0.X.n49 GNDA 0.028709f
C1107 two_stage_opamp_dummy_magic_14_0.X.n50 GNDA 0.026942f
C1108 two_stage_opamp_dummy_magic_14_0.X.n51 GNDA 0.016389f
C1109 two_stage_opamp_dummy_magic_14_0.X.n52 GNDA 0.506608f
C1110 two_stage_opamp_dummy_magic_14_0.X.t15 GNDA 0.439257f
C1111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 GNDA 0.345142f
C1112 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 GNDA 0.346293f
C1113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 GNDA 0.186001f
C1114 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 GNDA 0.198613f
C1115 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 GNDA 0.345142f
C1116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 GNDA 0.346293f
C1117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 GNDA 0.186001f
C1118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 GNDA 0.217197f
C1119 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 GNDA 0.345142f
C1120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 GNDA 0.346293f
C1121 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 GNDA 0.186001f
C1122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 GNDA 0.217197f
C1123 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 GNDA 0.345142f
C1124 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 GNDA 0.346293f
C1125 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 GNDA 0.186001f
C1126 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 GNDA 0.217197f
C1127 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 GNDA 0.345142f
C1128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 GNDA 0.346293f
C1129 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 GNDA 0.364878f
C1130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 GNDA 0.364878f
C1131 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 GNDA 0.186001f
C1132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 GNDA 0.217197f
C1133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 GNDA 0.345142f
C1134 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 GNDA 0.346293f
C1135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 GNDA 0.364878f
C1136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 GNDA 0.364878f
C1137 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 GNDA 0.186001f
C1138 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 GNDA 0.217197f
C1139 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 GNDA 0.346293f
C1140 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 GNDA 0.347548f
C1141 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 GNDA 0.346293f
C1142 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 GNDA 0.349008f
C1143 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 GNDA 0.379597f
C1144 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 GNDA 0.328964f
C1145 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 GNDA 0.346293f
C1146 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 GNDA 0.347548f
C1147 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 GNDA 0.328964f
C1148 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 GNDA 0.346293f
C1149 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 GNDA 0.347548f
C1150 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 GNDA 0.346293f
C1151 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 GNDA 0.347548f
C1152 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 GNDA 0.346293f
C1153 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 GNDA 0.347548f
C1154 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 GNDA 0.346293f
C1155 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 GNDA 0.347548f
C1156 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 GNDA 0.346293f
C1157 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 GNDA 0.347548f
C1158 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 GNDA 0.346293f
C1159 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 GNDA 0.347548f
C1160 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 GNDA 0.346293f
C1161 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 GNDA 0.347548f
C1162 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 GNDA 0.346293f
C1163 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 GNDA 0.347548f
C1164 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 GNDA 0.346293f
C1165 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 GNDA 0.347548f
C1166 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 GNDA 0.346293f
C1167 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 GNDA 0.347548f
C1168 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 GNDA 0.346293f
C1169 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 GNDA 0.347548f
C1170 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 GNDA 0.346293f
C1171 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 GNDA 0.347548f
C1172 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 GNDA 0.346293f
C1173 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 GNDA 0.347548f
C1174 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 GNDA 0.346293f
C1175 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 GNDA 0.347548f
C1176 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 GNDA 0.346293f
C1177 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 GNDA 0.347548f
C1178 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 GNDA 0.346293f
C1179 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 GNDA 0.347548f
C1180 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 GNDA 0.346293f
C1181 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 GNDA 0.347548f
C1182 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 GNDA 0.346293f
C1183 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 GNDA 0.347548f
C1184 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 GNDA 0.346293f
C1185 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 GNDA 0.347548f
C1186 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 GNDA 0.346293f
C1187 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 GNDA 0.347548f
C1188 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 GNDA 0.346293f
C1189 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 GNDA 0.347548f
C1190 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 GNDA 0.346293f
C1191 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 GNDA 0.347548f
C1192 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 GNDA 0.346293f
C1193 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 GNDA 0.347548f
C1194 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 GNDA 0.346293f
C1195 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 GNDA 0.347548f
C1196 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 GNDA 0.346293f
C1197 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 GNDA 0.347548f
C1198 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 GNDA 0.345142f
C1199 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 GNDA 0.346293f
C1200 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 GNDA 0.186001f
C1201 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 GNDA 0.198613f
C1202 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 GNDA 0.345142f
C1203 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 GNDA 0.346293f
C1204 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 GNDA 0.186001f
C1205 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 GNDA 0.217197f
C1206 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 GNDA 0.345142f
C1207 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 GNDA 0.346293f
C1208 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 GNDA 0.186001f
C1209 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 GNDA 0.217197f
C1210 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 GNDA 0.345142f
C1211 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 GNDA 0.346293f
C1212 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 GNDA 0.186001f
C1213 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 GNDA 0.217197f
C1214 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 GNDA 0.345142f
C1215 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 GNDA 0.346293f
C1216 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 GNDA 0.186001f
C1217 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 GNDA 0.217197f
C1218 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 GNDA 0.345142f
C1219 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 GNDA 0.346293f
C1220 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 GNDA 0.186001f
C1221 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 GNDA 0.217197f
C1222 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 GNDA 0.345142f
C1223 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 GNDA 0.346293f
C1224 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 GNDA 0.186001f
C1225 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 GNDA 0.217197f
C1226 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 GNDA 0.346293f
C1227 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 GNDA 0.186001f
C1228 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 GNDA 0.197462f
C1229 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 GNDA 0.346293f
C1230 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 GNDA 0.186001f
C1231 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 GNDA 0.197462f
C1232 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 GNDA 0.346293f
C1233 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 GNDA 0.347548f
C1234 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 GNDA 0.346293f
C1235 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 GNDA 0.347548f
C1236 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 GNDA 0.167416f
C1237 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 GNDA 0.215942f
C1238 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 GNDA 0.18485f
C1239 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 GNDA 0.234527f
C1240 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 GNDA 0.18485f
C1241 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 GNDA 0.251856f
C1242 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 GNDA 0.18485f
C1243 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 GNDA 0.251856f
C1244 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 GNDA 0.18485f
C1245 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 GNDA 0.251856f
C1246 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 GNDA 0.18485f
C1247 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 GNDA 0.251856f
C1248 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 GNDA 0.18485f
C1249 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 GNDA 0.251856f
C1250 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 GNDA 0.18485f
C1251 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 GNDA 0.251856f
C1252 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 GNDA 0.18485f
C1253 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 GNDA 0.251856f
C1254 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 GNDA 0.18485f
C1255 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 GNDA 0.251856f
C1256 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 GNDA 0.18485f
C1257 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 GNDA 0.251856f
C1258 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 GNDA 0.18485f
C1259 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 GNDA 0.251856f
C1260 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 GNDA 0.18485f
C1261 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 GNDA 0.251856f
C1262 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 GNDA 0.18485f
C1263 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 GNDA 0.251856f
C1264 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 GNDA 0.18485f
C1265 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 GNDA 0.251856f
C1266 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 GNDA 0.18485f
C1267 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 GNDA 0.251856f
C1268 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 GNDA 0.18485f
C1269 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 GNDA 0.234527f
C1270 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 GNDA 0.345142f
C1271 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 GNDA 0.167416f
C1272 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 GNDA 0.217197f
C1273 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 GNDA 0.345142f
C1274 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 GNDA 0.346293f
C1275 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 GNDA 0.364878f
C1276 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 GNDA 0.186001f
C1277 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 GNDA 0.217197f
C1278 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 GNDA 0.345142f
C1279 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 GNDA 0.217197f
C1280 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 GNDA 0.186001f
C1281 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 GNDA 0.364878f
C1282 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 GNDA 0.364878f
C1283 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 GNDA 0.730561f
C1284 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 GNDA 0.29977f
C1285 VOUT+.t16 GNDA 0.04876f
C1286 VOUT+.t2 GNDA 0.04876f
C1287 VOUT+.n0 GNDA 0.22634f
C1288 VOUT+.t14 GNDA 0.04876f
C1289 VOUT+.t11 GNDA 0.04876f
C1290 VOUT+.n1 GNDA 0.22561f
C1291 VOUT+.n2 GNDA 0.138742f
C1292 VOUT+.t8 GNDA 0.04876f
C1293 VOUT+.t15 GNDA 0.04876f
C1294 VOUT+.n3 GNDA 0.22561f
C1295 VOUT+.n4 GNDA 0.077288f
C1296 VOUT+.t10 GNDA 0.081164f
C1297 VOUT+.n5 GNDA 0.091784f
C1298 VOUT+.t12 GNDA 0.041794f
C1299 VOUT+.t0 GNDA 0.041794f
C1300 VOUT+.n6 GNDA 0.168982f
C1301 VOUT+.t4 GNDA 0.041794f
C1302 VOUT+.t7 GNDA 0.041794f
C1303 VOUT+.n7 GNDA 0.16868f
C1304 VOUT+.n8 GNDA 0.164566f
C1305 VOUT+.t17 GNDA 0.041794f
C1306 VOUT+.t3 GNDA 0.041794f
C1307 VOUT+.n9 GNDA 0.16868f
C1308 VOUT+.n10 GNDA 0.084872f
C1309 VOUT+.t5 GNDA 0.041794f
C1310 VOUT+.t9 GNDA 0.041794f
C1311 VOUT+.n11 GNDA 0.16868f
C1312 VOUT+.n12 GNDA 0.084872f
C1313 VOUT+.t6 GNDA 0.041794f
C1314 VOUT+.t13 GNDA 0.041794f
C1315 VOUT+.n13 GNDA 0.168981f
C1316 VOUT+.n14 GNDA 0.100592f
C1317 VOUT+.t1 GNDA 0.041794f
C1318 VOUT+.t18 GNDA 0.041794f
C1319 VOUT+.n15 GNDA 0.166683f
C1320 VOUT+.n16 GNDA 0.135258f
C1321 VOUT+.t45 GNDA 0.278629f
C1322 VOUT+.t150 GNDA 0.283374f
C1323 VOUT+.t101 GNDA 0.278629f
C1324 VOUT+.n17 GNDA 0.186811f
C1325 VOUT+.n18 GNDA 0.1219f
C1326 VOUT+.t91 GNDA 0.28278f
C1327 VOUT+.t38 GNDA 0.28278f
C1328 VOUT+.t130 GNDA 0.28278f
C1329 VOUT+.t90 GNDA 0.28278f
C1330 VOUT+.t80 GNDA 0.28278f
C1331 VOUT+.t128 GNDA 0.28278f
C1332 VOUT+.t124 GNDA 0.28278f
C1333 VOUT+.t32 GNDA 0.28278f
C1334 VOUT+.t70 GNDA 0.28278f
C1335 VOUT+.t73 GNDA 0.28278f
C1336 VOUT+.t23 GNDA 0.28278f
C1337 VOUT+.t108 GNDA 0.28278f
C1338 VOUT+.t62 GNDA 0.28278f
C1339 VOUT+.t19 GNDA 0.28278f
C1340 VOUT+.t151 GNDA 0.28278f
C1341 VOUT+.t49 GNDA 0.28278f
C1342 VOUT+.t85 GNDA 0.278629f
C1343 VOUT+.n19 GNDA 0.305154f
C1344 VOUT+.t48 GNDA 0.278629f
C1345 VOUT+.n20 GNDA 0.357397f
C1346 VOUT+.t138 GNDA 0.278629f
C1347 VOUT+.n21 GNDA 0.357397f
C1348 VOUT+.t107 GNDA 0.278629f
C1349 VOUT+.n22 GNDA 0.357397f
C1350 VOUT+.t71 GNDA 0.278629f
C1351 VOUT+.n23 GNDA 0.357397f
C1352 VOUT+.t25 GNDA 0.278629f
C1353 VOUT+.n24 GNDA 0.357397f
C1354 VOUT+.t129 GNDA 0.278629f
C1355 VOUT+.n25 GNDA 0.357397f
C1356 VOUT+.t87 GNDA 0.278629f
C1357 VOUT+.n26 GNDA 0.239648f
C1358 VOUT+.t52 GNDA 0.278629f
C1359 VOUT+.n27 GNDA 0.239648f
C1360 VOUT+.t141 GNDA 0.278629f
C1361 VOUT+.t75 GNDA 0.283374f
C1362 VOUT+.t111 GNDA 0.278629f
C1363 VOUT+.n28 GNDA 0.186811f
C1364 VOUT+.n29 GNDA 0.226386f
C1365 VOUT+.t54 GNDA 0.283374f
C1366 VOUT+.t24 GNDA 0.278629f
C1367 VOUT+.n30 GNDA 0.186811f
C1368 VOUT+.t114 GNDA 0.278629f
C1369 VOUT+.t34 GNDA 0.283374f
C1370 VOUT+.t74 GNDA 0.278629f
C1371 VOUT+.n31 GNDA 0.186811f
C1372 VOUT+.n32 GNDA 0.226386f
C1373 VOUT+.t95 GNDA 0.283374f
C1374 VOUT+.t59 GNDA 0.278629f
C1375 VOUT+.n33 GNDA 0.186811f
C1376 VOUT+.t148 GNDA 0.278629f
C1377 VOUT+.t79 GNDA 0.283374f
C1378 VOUT+.t117 GNDA 0.278629f
C1379 VOUT+.n34 GNDA 0.186811f
C1380 VOUT+.n35 GNDA 0.226386f
C1381 VOUT+.t134 GNDA 0.283374f
C1382 VOUT+.t100 GNDA 0.278629f
C1383 VOUT+.n36 GNDA 0.186811f
C1384 VOUT+.t44 GNDA 0.278629f
C1385 VOUT+.t122 GNDA 0.283374f
C1386 VOUT+.t153 GNDA 0.278629f
C1387 VOUT+.n37 GNDA 0.186811f
C1388 VOUT+.n38 GNDA 0.226386f
C1389 VOUT+.t102 GNDA 0.283374f
C1390 VOUT+.t66 GNDA 0.278629f
C1391 VOUT+.n39 GNDA 0.186811f
C1392 VOUT+.t154 GNDA 0.278629f
C1393 VOUT+.t82 GNDA 0.283374f
C1394 VOUT+.t123 GNDA 0.278629f
C1395 VOUT+.n40 GNDA 0.186811f
C1396 VOUT+.n41 GNDA 0.226386f
C1397 VOUT+.t137 GNDA 0.283374f
C1398 VOUT+.t106 GNDA 0.278629f
C1399 VOUT+.n42 GNDA 0.186811f
C1400 VOUT+.t51 GNDA 0.278629f
C1401 VOUT+.t126 GNDA 0.283374f
C1402 VOUT+.t22 GNDA 0.278629f
C1403 VOUT+.n43 GNDA 0.186811f
C1404 VOUT+.n44 GNDA 0.226386f
C1405 VOUT+.t132 GNDA 0.278629f
C1406 VOUT+.t56 GNDA 0.283374f
C1407 VOUT+.t96 GNDA 0.278629f
C1408 VOUT+.n45 GNDA 0.186811f
C1409 VOUT+.n46 GNDA 0.1219f
C1410 VOUT+.t116 GNDA 0.28278f
C1411 VOUT+.t105 GNDA 0.283374f
C1412 VOUT+.t69 GNDA 0.278629f
C1413 VOUT+.n47 GNDA 0.182458f
C1414 VOUT+.t147 GNDA 0.28278f
C1415 VOUT+.t29 GNDA 0.283374f
C1416 VOUT+.t139 GNDA 0.278629f
C1417 VOUT+.n48 GNDA 0.186811f
C1418 VOUT+.t109 GNDA 0.278629f
C1419 VOUT+.n49 GNDA 0.117546f
C1420 VOUT+.t43 GNDA 0.28278f
C1421 VOUT+.t60 GNDA 0.283374f
C1422 VOUT+.t37 GNDA 0.278629f
C1423 VOUT+.n50 GNDA 0.186811f
C1424 VOUT+.t144 GNDA 0.278629f
C1425 VOUT+.n51 GNDA 0.117546f
C1426 VOUT+.t83 GNDA 0.28278f
C1427 VOUT+.t115 GNDA 0.283374f
C1428 VOUT+.t21 GNDA 0.278629f
C1429 VOUT+.n52 GNDA 0.186811f
C1430 VOUT+.t125 GNDA 0.278629f
C1431 VOUT+.n53 GNDA 0.117546f
C1432 VOUT+.t63 GNDA 0.28278f
C1433 VOUT+.t26 GNDA 0.28278f
C1434 VOUT+.t103 GNDA 0.28278f
C1435 VOUT+.t57 GNDA 0.283013f
C1436 VOUT+.t135 GNDA 0.28278f
C1437 VOUT+.t33 GNDA 0.283013f
C1438 VOUT+.t120 GNDA 0.28278f
C1439 VOUT+.t77 GNDA 0.283013f
C1440 VOUT+.t155 GNDA 0.28278f
C1441 VOUT+.t119 GNDA 0.278629f
C1442 VOUT+.n54 GNDA 0.308404f
C1443 VOUT+.t78 GNDA 0.278629f
C1444 VOUT+.n55 GNDA 0.360646f
C1445 VOUT+.t97 GNDA 0.278629f
C1446 VOUT+.n56 GNDA 0.360646f
C1447 VOUT+.t61 GNDA 0.278629f
C1448 VOUT+.n57 GNDA 0.357397f
C1449 VOUT+.t27 GNDA 0.278629f
C1450 VOUT+.n58 GNDA 0.296245f
C1451 VOUT+.t41 GNDA 0.278629f
C1452 VOUT+.n59 GNDA 0.296245f
C1453 VOUT+.t145 GNDA 0.278629f
C1454 VOUT+.n60 GNDA 0.296245f
C1455 VOUT+.t113 GNDA 0.278629f
C1456 VOUT+.n61 GNDA 0.296245f
C1457 VOUT+.t72 GNDA 0.278629f
C1458 VOUT+.n62 GNDA 0.239648f
C1459 VOUT+.t92 GNDA 0.278629f
C1460 VOUT+.t20 GNDA 0.283374f
C1461 VOUT+.t55 GNDA 0.278629f
C1462 VOUT+.n63 GNDA 0.186811f
C1463 VOUT+.n64 GNDA 0.226386f
C1464 VOUT+.t31 GNDA 0.283374f
C1465 VOUT+.t50 GNDA 0.278629f
C1466 VOUT+.t121 GNDA 0.283374f
C1467 VOUT+.t156 GNDA 0.278629f
C1468 VOUT+.n65 GNDA 0.186811f
C1469 VOUT+.n66 GNDA 0.291297f
C1470 VOUT+.t67 GNDA 0.283374f
C1471 VOUT+.t86 GNDA 0.278629f
C1472 VOUT+.t152 GNDA 0.283374f
C1473 VOUT+.t47 GNDA 0.278629f
C1474 VOUT+.n67 GNDA 0.186811f
C1475 VOUT+.n68 GNDA 0.291297f
C1476 VOUT+.t131 GNDA 0.283374f
C1477 VOUT+.t94 GNDA 0.278629f
C1478 VOUT+.n69 GNDA 0.186811f
C1479 VOUT+.t39 GNDA 0.278629f
C1480 VOUT+.t118 GNDA 0.283374f
C1481 VOUT+.t146 GNDA 0.278629f
C1482 VOUT+.n70 GNDA 0.186811f
C1483 VOUT+.n71 GNDA 0.226386f
C1484 VOUT+.t89 GNDA 0.283374f
C1485 VOUT+.t53 GNDA 0.278629f
C1486 VOUT+.n72 GNDA 0.186811f
C1487 VOUT+.t142 GNDA 0.278629f
C1488 VOUT+.t76 GNDA 0.283374f
C1489 VOUT+.t112 GNDA 0.278629f
C1490 VOUT+.n73 GNDA 0.186811f
C1491 VOUT+.n74 GNDA 0.226386f
C1492 VOUT+.t127 GNDA 0.283374f
C1493 VOUT+.t88 GNDA 0.278629f
C1494 VOUT+.n75 GNDA 0.186811f
C1495 VOUT+.t35 GNDA 0.278629f
C1496 VOUT+.t110 GNDA 0.283374f
C1497 VOUT+.t140 GNDA 0.278629f
C1498 VOUT+.n76 GNDA 0.186811f
C1499 VOUT+.n77 GNDA 0.226386f
C1500 VOUT+.t84 GNDA 0.283374f
C1501 VOUT+.t46 GNDA 0.278629f
C1502 VOUT+.n78 GNDA 0.186811f
C1503 VOUT+.t136 GNDA 0.278629f
C1504 VOUT+.t68 GNDA 0.283374f
C1505 VOUT+.t104 GNDA 0.278629f
C1506 VOUT+.n79 GNDA 0.186811f
C1507 VOUT+.n80 GNDA 0.226386f
C1508 VOUT+.t42 GNDA 0.283374f
C1509 VOUT+.t149 GNDA 0.278629f
C1510 VOUT+.n81 GNDA 0.186811f
C1511 VOUT+.t99 GNDA 0.278629f
C1512 VOUT+.t30 GNDA 0.283374f
C1513 VOUT+.t65 GNDA 0.278629f
C1514 VOUT+.n82 GNDA 0.186811f
C1515 VOUT+.n83 GNDA 0.226386f
C1516 VOUT+.t81 GNDA 0.283374f
C1517 VOUT+.t40 GNDA 0.278629f
C1518 VOUT+.n84 GNDA 0.186811f
C1519 VOUT+.t133 GNDA 0.278629f
C1520 VOUT+.t64 GNDA 0.283374f
C1521 VOUT+.t98 GNDA 0.278629f
C1522 VOUT+.n85 GNDA 0.186811f
C1523 VOUT+.n86 GNDA 0.226386f
C1524 VOUT+.t28 GNDA 0.283374f
C1525 VOUT+.t58 GNDA 0.278629f
C1526 VOUT+.n87 GNDA 0.186811f
C1527 VOUT+.t93 GNDA 0.278629f
C1528 VOUT+.n88 GNDA 0.226386f
C1529 VOUT+.t143 GNDA 0.278629f
C1530 VOUT+.n89 GNDA 0.1219f
C1531 VOUT+.t36 GNDA 0.278629f
C1532 VOUT+.n90 GNDA 0.177758f
C1533 VOUT+.n91 GNDA 0.205844f
C1534 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 GNDA 0.013072f
C1535 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 GNDA 0.013072f
C1536 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 GNDA 0.026144f
C1537 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 GNDA 0.013072f
C1538 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 GNDA 0.013072f
C1539 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 GNDA 0.065442f
C1540 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 GNDA 0.108875f
C1541 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 GNDA 0.017402f
C1542 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 GNDA 0.017402f
C1543 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 GNDA 0.017402f
C1544 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 GNDA 0.017402f
C1545 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 GNDA 0.017402f
C1546 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 GNDA 0.017402f
C1547 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 GNDA 0.017402f
C1548 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 GNDA 0.017402f
C1549 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 GNDA 0.017402f
C1550 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 GNDA 0.017402f
C1551 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 GNDA 0.017402f
C1552 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 GNDA 0.017402f
C1553 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 GNDA 0.017402f
C1554 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 GNDA 0.017402f
C1555 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 GNDA 0.017402f
C1556 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 GNDA 0.020311f
C1557 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 GNDA 0.01915f
C1558 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 GNDA 0.01201f
C1559 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 GNDA 0.01201f
C1560 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 GNDA 0.01201f
C1561 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 GNDA 0.01201f
C1562 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 GNDA 0.01201f
C1563 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 GNDA 0.01201f
C1564 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 GNDA 0.01201f
C1565 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 GNDA 0.01201f
C1566 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 GNDA 0.01201f
C1567 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 GNDA 0.01201f
C1568 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 GNDA 0.01201f
C1569 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 GNDA 0.01201f
C1570 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 GNDA 0.01201f
C1571 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 GNDA 0.010738f
C1572 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 GNDA 0.017402f
C1573 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 GNDA 0.020311f
C1574 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 GNDA 0.017878f
C1575 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 GNDA 0.018177f
C1576 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 GNDA 0.018384f
C1577 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 GNDA 0.018384f
C1578 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 GNDA 0.02545f
C1579 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 GNDA 0.161233f
C1580 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 GNDA 0.033195f
C1581 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 GNDA 0.037735f
C1582 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 GNDA 0.116306f
C1583 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 GNDA 0.407855f
C1584 bgr_7_0.TAIL_CUR_MIR_BIAS GNDA 0.548373f
C1585 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 GNDA 0.346251f
C1586 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 GNDA 0.347506f
C1587 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 GNDA 0.346251f
C1588 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 GNDA 0.348966f
C1589 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 GNDA 0.379551f
C1590 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 GNDA 0.346251f
C1591 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 GNDA 0.347506f
C1592 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 GNDA 0.328924f
C1593 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 GNDA 0.346251f
C1594 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 GNDA 0.347506f
C1595 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 GNDA 0.328924f
C1596 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 GNDA 0.346251f
C1597 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 GNDA 0.347506f
C1598 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 GNDA 0.346251f
C1599 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 GNDA 0.347506f
C1600 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 GNDA 0.346251f
C1601 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 GNDA 0.347506f
C1602 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 GNDA 0.346251f
C1603 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 GNDA 0.347506f
C1604 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 GNDA 0.346251f
C1605 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 GNDA 0.347506f
C1606 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 GNDA 0.346251f
C1607 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 GNDA 0.347506f
C1608 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 GNDA 0.346251f
C1609 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 GNDA 0.347506f
C1610 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 GNDA 0.346251f
C1611 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 GNDA 0.347506f
C1612 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 GNDA 0.346251f
C1613 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 GNDA 0.347506f
C1614 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 GNDA 0.346251f
C1615 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 GNDA 0.347506f
C1616 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 GNDA 0.346251f
C1617 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 GNDA 0.347506f
C1618 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 GNDA 0.346251f
C1619 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 GNDA 0.347506f
C1620 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 GNDA 0.346251f
C1621 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 GNDA 0.347506f
C1622 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 GNDA 0.346251f
C1623 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 GNDA 0.347506f
C1624 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 GNDA 0.346251f
C1625 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 GNDA 0.347506f
C1626 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 GNDA 0.346251f
C1627 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 GNDA 0.347506f
C1628 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 GNDA 0.346251f
C1629 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 GNDA 0.347506f
C1630 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 GNDA 0.346251f
C1631 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 GNDA 0.347506f
C1632 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 GNDA 0.346251f
C1633 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 GNDA 0.347506f
C1634 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 GNDA 0.346251f
C1635 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 GNDA 0.347506f
C1636 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 GNDA 0.346251f
C1637 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 GNDA 0.347506f
C1638 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 GNDA 0.346251f
C1639 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 GNDA 0.347506f
C1640 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 GNDA 0.346251f
C1641 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 GNDA 0.347506f
C1642 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 GNDA 0.346251f
C1643 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 GNDA 0.347506f
C1644 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 GNDA 0.346251f
C1645 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 GNDA 0.347506f
C1646 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 GNDA 0.3451f
C1647 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 GNDA 0.346251f
C1648 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 GNDA 0.185978f
C1649 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 GNDA 0.198589f
C1650 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 GNDA 0.3451f
C1651 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 GNDA 0.346251f
C1652 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 GNDA 0.185978f
C1653 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 GNDA 0.217171f
C1654 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 GNDA 0.3451f
C1655 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 GNDA 0.346251f
C1656 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 GNDA 0.185978f
C1657 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 GNDA 0.217171f
C1658 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 GNDA 0.3451f
C1659 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 GNDA 0.346251f
C1660 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 GNDA 0.185978f
C1661 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 GNDA 0.217171f
C1662 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 GNDA 0.3451f
C1663 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 GNDA 0.346251f
C1664 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 GNDA 0.185978f
C1665 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 GNDA 0.217171f
C1666 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 GNDA 0.3451f
C1667 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 GNDA 0.346251f
C1668 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 GNDA 0.185978f
C1669 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 GNDA 0.217171f
C1670 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 GNDA 0.3451f
C1671 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 GNDA 0.346251f
C1672 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 GNDA 0.185978f
C1673 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 GNDA 0.217171f
C1674 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 GNDA 0.346251f
C1675 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 GNDA 0.185978f
C1676 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 GNDA 0.197438f
C1677 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 GNDA 0.346251f
C1678 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 GNDA 0.185978f
C1679 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 GNDA 0.197438f
C1680 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 GNDA 0.346251f
C1681 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 GNDA 0.347506f
C1682 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 GNDA 0.167396f
C1683 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 GNDA 0.215916f
C1684 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 GNDA 0.184828f
C1685 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 GNDA 0.234498f
C1686 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 GNDA 0.184828f
C1687 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 GNDA 0.251826f
C1688 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 GNDA 0.184828f
C1689 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 GNDA 0.251826f
C1690 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 GNDA 0.184828f
C1691 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 GNDA 0.251826f
C1692 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 GNDA 0.184828f
C1693 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 GNDA 0.251826f
C1694 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 GNDA 0.184828f
C1695 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 GNDA 0.251826f
C1696 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 GNDA 0.184828f
C1697 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 GNDA 0.251826f
C1698 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 GNDA 0.184828f
C1699 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 GNDA 0.251826f
C1700 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 GNDA 0.184828f
C1701 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 GNDA 0.251826f
C1702 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 GNDA 0.184828f
C1703 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 GNDA 0.251826f
C1704 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 GNDA 0.184828f
C1705 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 GNDA 0.251826f
C1706 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 GNDA 0.184828f
C1707 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 GNDA 0.251826f
C1708 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 GNDA 0.184828f
C1709 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 GNDA 0.251826f
C1710 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 GNDA 0.184828f
C1711 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 GNDA 0.251826f
C1712 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 GNDA 0.184828f
C1713 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 GNDA 0.251826f
C1714 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 GNDA 0.184828f
C1715 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 GNDA 0.234498f
C1716 two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 GNDA 0.3451f
C1717 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 GNDA 0.167396f
C1718 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 GNDA 0.217171f
C1719 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 GNDA 0.3451f
C1720 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 GNDA 0.346251f
C1721 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 GNDA 0.364834f
C1722 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 GNDA 0.185978f
C1723 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 GNDA 0.217171f
C1724 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 GNDA 0.3451f
C1725 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 GNDA 0.346251f
C1726 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 GNDA 0.185978f
C1727 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 GNDA 0.198589f
C1728 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 GNDA 0.3451f
C1729 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 GNDA 0.346251f
C1730 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 GNDA 0.185978f
C1731 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 GNDA 0.217171f
C1732 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 GNDA 0.3451f
C1733 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 GNDA 0.346251f
C1734 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 GNDA 0.185978f
C1735 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 GNDA 0.217171f
C1736 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 GNDA 0.3451f
C1737 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 GNDA 0.346251f
C1738 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 GNDA 0.185978f
C1739 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 GNDA 0.217171f
C1740 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 GNDA 0.3451f
C1741 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 GNDA 0.346251f
C1742 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 GNDA 0.364834f
C1743 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 GNDA 0.364834f
C1744 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 GNDA 0.185978f
C1745 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 GNDA 0.217171f
C1746 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 GNDA 0.3451f
C1747 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 GNDA 0.346251f
C1748 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 GNDA 0.364834f
C1749 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 GNDA 0.364834f
C1750 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 GNDA 0.185978f
C1751 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 GNDA 0.217171f
C1752 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 GNDA 0.3451f
C1753 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 GNDA 0.217171f
C1754 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 GNDA 0.185978f
C1755 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 GNDA 0.364834f
C1756 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 GNDA 0.364834f
C1757 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 GNDA 0.430822f
C1758 two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 GNDA 0.292647f
C1759 VOUT-.t8 GNDA 0.041794f
C1760 VOUT-.t2 GNDA 0.041794f
C1761 VOUT-.n0 GNDA 0.168982f
C1762 VOUT-.t12 GNDA 0.041794f
C1763 VOUT-.t9 GNDA 0.041794f
C1764 VOUT-.n1 GNDA 0.168981f
C1765 VOUT-.t6 GNDA 0.041794f
C1766 VOUT-.t0 GNDA 0.041794f
C1767 VOUT-.n2 GNDA 0.16868f
C1768 VOUT-.n3 GNDA 0.164567f
C1769 VOUT-.t14 GNDA 0.041794f
C1770 VOUT-.t13 GNDA 0.041794f
C1771 VOUT-.n4 GNDA 0.16868f
C1772 VOUT-.n5 GNDA 0.084872f
C1773 VOUT-.t16 GNDA 0.041794f
C1774 VOUT-.t5 GNDA 0.041794f
C1775 VOUT-.n6 GNDA 0.16868f
C1776 VOUT-.n7 GNDA 0.084872f
C1777 VOUT-.n8 GNDA 0.100591f
C1778 VOUT-.t17 GNDA 0.041794f
C1779 VOUT-.t15 GNDA 0.041794f
C1780 VOUT-.n9 GNDA 0.166683f
C1781 VOUT-.n10 GNDA 0.135258f
C1782 VOUT-.t26 GNDA 0.283374f
C1783 VOUT-.t119 GNDA 0.278628f
C1784 VOUT-.n11 GNDA 0.186811f
C1785 VOUT-.t33 GNDA 0.278628f
C1786 VOUT-.n12 GNDA 0.1219f
C1787 VOUT-.t36 GNDA 0.283374f
C1788 VOUT-.t122 GNDA 0.278628f
C1789 VOUT-.n13 GNDA 0.186811f
C1790 VOUT-.t90 GNDA 0.278628f
C1791 VOUT-.t82 GNDA 0.28278f
C1792 VOUT-.t42 GNDA 0.28278f
C1793 VOUT-.t92 GNDA 0.28278f
C1794 VOUT-.t74 GNDA 0.28278f
C1795 VOUT-.t141 GNDA 0.28278f
C1796 VOUT-.t38 GNDA 0.28278f
C1797 VOUT-.t105 GNDA 0.28278f
C1798 VOUT-.t126 GNDA 0.28278f
C1799 VOUT-.t154 GNDA 0.28278f
C1800 VOUT-.t95 GNDA 0.28278f
C1801 VOUT-.t65 GNDA 0.28278f
C1802 VOUT-.t62 GNDA 0.28278f
C1803 VOUT-.t114 GNDA 0.28278f
C1804 VOUT-.t24 GNDA 0.28278f
C1805 VOUT-.t71 GNDA 0.28278f
C1806 VOUT-.t113 GNDA 0.28278f
C1807 VOUT-.t148 GNDA 0.278628f
C1808 VOUT-.n14 GNDA 0.305154f
C1809 VOUT-.t60 GNDA 0.278628f
C1810 VOUT-.n15 GNDA 0.357397f
C1811 VOUT-.t93 GNDA 0.278628f
C1812 VOUT-.n16 GNDA 0.357397f
C1813 VOUT-.t127 GNDA 0.278628f
C1814 VOUT-.n17 GNDA 0.357397f
C1815 VOUT-.t25 GNDA 0.278628f
C1816 VOUT-.n18 GNDA 0.357397f
C1817 VOUT-.t72 GNDA 0.278628f
C1818 VOUT-.n19 GNDA 0.357397f
C1819 VOUT-.t110 GNDA 0.278628f
C1820 VOUT-.n20 GNDA 0.357397f
C1821 VOUT-.t142 GNDA 0.278628f
C1822 VOUT-.n21 GNDA 0.239648f
C1823 VOUT-.t56 GNDA 0.278628f
C1824 VOUT-.n22 GNDA 0.239648f
C1825 VOUT-.n23 GNDA 0.226386f
C1826 VOUT-.t140 GNDA 0.283374f
C1827 VOUT-.t89 GNDA 0.278628f
C1828 VOUT-.n24 GNDA 0.186811f
C1829 VOUT-.t59 GNDA 0.278628f
C1830 VOUT-.t111 GNDA 0.283374f
C1831 VOUT-.t21 GNDA 0.278628f
C1832 VOUT-.n25 GNDA 0.186811f
C1833 VOUT-.n26 GNDA 0.226386f
C1834 VOUT-.t41 GNDA 0.283374f
C1835 VOUT-.t129 GNDA 0.278628f
C1836 VOUT-.n27 GNDA 0.186811f
C1837 VOUT-.t98 GNDA 0.278628f
C1838 VOUT-.t151 GNDA 0.283374f
C1839 VOUT-.t63 GNDA 0.278628f
C1840 VOUT-.n28 GNDA 0.186811f
C1841 VOUT-.n29 GNDA 0.226386f
C1842 VOUT-.t80 GNDA 0.283374f
C1843 VOUT-.t30 GNDA 0.278628f
C1844 VOUT-.n30 GNDA 0.186811f
C1845 VOUT-.t134 GNDA 0.278628f
C1846 VOUT-.t51 GNDA 0.283374f
C1847 VOUT-.t103 GNDA 0.278628f
C1848 VOUT-.n31 GNDA 0.186811f
C1849 VOUT-.n32 GNDA 0.226386f
C1850 VOUT-.t49 GNDA 0.283374f
C1851 VOUT-.t135 GNDA 0.278628f
C1852 VOUT-.n33 GNDA 0.186811f
C1853 VOUT-.t102 GNDA 0.278628f
C1854 VOUT-.t19 GNDA 0.283374f
C1855 VOUT-.t67 GNDA 0.278628f
C1856 VOUT-.n34 GNDA 0.186811f
C1857 VOUT-.n35 GNDA 0.226386f
C1858 VOUT-.t85 GNDA 0.283374f
C1859 VOUT-.t34 GNDA 0.278628f
C1860 VOUT-.n36 GNDA 0.186811f
C1861 VOUT-.t139 GNDA 0.278628f
C1862 VOUT-.t55 GNDA 0.283374f
C1863 VOUT-.t106 GNDA 0.278628f
C1864 VOUT-.n37 GNDA 0.186811f
C1865 VOUT-.n38 GNDA 0.226386f
C1866 VOUT-.t68 GNDA 0.283374f
C1867 VOUT-.t86 GNDA 0.278628f
C1868 VOUT-.n39 GNDA 0.186811f
C1869 VOUT-.t54 GNDA 0.278628f
C1870 VOUT-.n40 GNDA 0.1219f
C1871 VOUT-.t29 GNDA 0.283374f
C1872 VOUT-.t52 GNDA 0.278628f
C1873 VOUT-.n41 GNDA 0.186811f
C1874 VOUT-.t155 GNDA 0.278628f
C1875 VOUT-.t156 GNDA 0.28278f
C1876 VOUT-.t132 GNDA 0.283374f
C1877 VOUT-.t99 GNDA 0.278628f
C1878 VOUT-.n42 GNDA 0.182458f
C1879 VOUT-.t35 GNDA 0.28278f
C1880 VOUT-.t150 GNDA 0.283374f
C1881 VOUT-.t94 GNDA 0.278628f
C1882 VOUT-.n43 GNDA 0.186811f
C1883 VOUT-.t61 GNDA 0.278628f
C1884 VOUT-.n44 GNDA 0.117546f
C1885 VOUT-.t137 GNDA 0.28278f
C1886 VOUT-.t115 GNDA 0.283374f
C1887 VOUT-.t58 GNDA 0.278628f
C1888 VOUT-.n45 GNDA 0.186811f
C1889 VOUT-.t22 GNDA 0.278628f
C1890 VOUT-.n46 GNDA 0.117546f
C1891 VOUT-.t104 GNDA 0.28278f
C1892 VOUT-.t66 GNDA 0.283374f
C1893 VOUT-.t77 GNDA 0.278628f
C1894 VOUT-.n47 GNDA 0.186811f
C1895 VOUT-.t43 GNDA 0.278628f
C1896 VOUT-.n48 GNDA 0.117546f
C1897 VOUT-.t120 GNDA 0.28278f
C1898 VOUT-.t144 GNDA 0.28278f
C1899 VOUT-.t83 GNDA 0.28278f
C1900 VOUT-.t107 GNDA 0.283013f
C1901 VOUT-.t50 GNDA 0.28278f
C1902 VOUT-.t69 GNDA 0.283013f
C1903 VOUT-.t149 GNDA 0.28278f
C1904 VOUT-.t91 GNDA 0.283013f
C1905 VOUT-.t31 GNDA 0.28278f
C1906 VOUT-.t130 GNDA 0.278628f
C1907 VOUT-.n49 GNDA 0.308404f
C1908 VOUT-.t108 GNDA 0.278628f
C1909 VOUT-.n50 GNDA 0.360646f
C1910 VOUT-.t146 GNDA 0.278628f
C1911 VOUT-.n51 GNDA 0.360646f
C1912 VOUT-.t45 GNDA 0.278628f
C1913 VOUT-.n52 GNDA 0.357397f
C1914 VOUT-.t81 GNDA 0.278628f
C1915 VOUT-.n53 GNDA 0.296245f
C1916 VOUT-.t64 GNDA 0.278628f
C1917 VOUT-.n54 GNDA 0.296245f
C1918 VOUT-.t100 GNDA 0.278628f
C1919 VOUT-.n55 GNDA 0.296245f
C1920 VOUT-.t136 GNDA 0.278628f
C1921 VOUT-.n56 GNDA 0.296245f
C1922 VOUT-.t116 GNDA 0.278628f
C1923 VOUT-.n57 GNDA 0.239648f
C1924 VOUT-.n58 GNDA 0.226386f
C1925 VOUT-.t125 GNDA 0.283374f
C1926 VOUT-.t152 GNDA 0.278628f
C1927 VOUT-.n59 GNDA 0.186811f
C1928 VOUT-.t112 GNDA 0.278628f
C1929 VOUT-.t73 GNDA 0.283374f
C1930 VOUT-.n60 GNDA 0.291297f
C1931 VOUT-.t23 GNDA 0.283374f
C1932 VOUT-.t47 GNDA 0.278628f
C1933 VOUT-.n61 GNDA 0.186811f
C1934 VOUT-.t147 GNDA 0.278628f
C1935 VOUT-.t109 GNDA 0.283374f
C1936 VOUT-.n62 GNDA 0.291297f
C1937 VOUT-.t76 GNDA 0.283374f
C1938 VOUT-.t27 GNDA 0.278628f
C1939 VOUT-.n63 GNDA 0.186811f
C1940 VOUT-.t128 GNDA 0.278628f
C1941 VOUT-.t44 GNDA 0.283374f
C1942 VOUT-.t97 GNDA 0.278628f
C1943 VOUT-.n64 GNDA 0.186811f
C1944 VOUT-.n65 GNDA 0.226386f
C1945 VOUT-.t37 GNDA 0.283374f
C1946 VOUT-.t123 GNDA 0.278628f
C1947 VOUT-.n66 GNDA 0.186811f
C1948 VOUT-.t88 GNDA 0.278628f
C1949 VOUT-.t143 GNDA 0.283374f
C1950 VOUT-.t57 GNDA 0.278628f
C1951 VOUT-.n67 GNDA 0.186811f
C1952 VOUT-.n68 GNDA 0.226386f
C1953 VOUT-.t70 GNDA 0.283374f
C1954 VOUT-.t20 GNDA 0.278628f
C1955 VOUT-.n69 GNDA 0.186811f
C1956 VOUT-.t121 GNDA 0.278628f
C1957 VOUT-.t39 GNDA 0.283374f
C1958 VOUT-.t87 GNDA 0.278628f
C1959 VOUT-.n70 GNDA 0.186811f
C1960 VOUT-.n71 GNDA 0.226386f
C1961 VOUT-.t32 GNDA 0.283374f
C1962 VOUT-.t118 GNDA 0.278628f
C1963 VOUT-.n72 GNDA 0.186811f
C1964 VOUT-.t84 GNDA 0.278628f
C1965 VOUT-.t138 GNDA 0.283374f
C1966 VOUT-.t53 GNDA 0.278628f
C1967 VOUT-.n73 GNDA 0.186811f
C1968 VOUT-.n74 GNDA 0.226386f
C1969 VOUT-.t131 GNDA 0.283374f
C1970 VOUT-.t79 GNDA 0.278628f
C1971 VOUT-.n75 GNDA 0.186811f
C1972 VOUT-.t48 GNDA 0.278628f
C1973 VOUT-.t101 GNDA 0.283374f
C1974 VOUT-.t153 GNDA 0.278628f
C1975 VOUT-.n76 GNDA 0.186811f
C1976 VOUT-.n77 GNDA 0.226386f
C1977 VOUT-.t28 GNDA 0.283374f
C1978 VOUT-.t117 GNDA 0.278628f
C1979 VOUT-.n78 GNDA 0.186811f
C1980 VOUT-.t78 GNDA 0.278628f
C1981 VOUT-.t133 GNDA 0.283374f
C1982 VOUT-.t46 GNDA 0.278628f
C1983 VOUT-.n79 GNDA 0.186811f
C1984 VOUT-.n80 GNDA 0.226386f
C1985 VOUT-.t124 GNDA 0.283374f
C1986 VOUT-.t75 GNDA 0.278628f
C1987 VOUT-.n81 GNDA 0.186811f
C1988 VOUT-.t40 GNDA 0.278628f
C1989 VOUT-.n82 GNDA 0.226386f
C1990 VOUT-.t145 GNDA 0.278628f
C1991 VOUT-.n83 GNDA 0.1219f
C1992 VOUT-.t96 GNDA 0.278628f
C1993 VOUT-.n84 GNDA 0.177758f
C1994 VOUT-.n85 GNDA 0.20704f
C1995 VOUT-.t3 GNDA 0.04876f
C1996 VOUT-.t10 GNDA 0.04876f
C1997 VOUT-.n86 GNDA 0.22634f
C1998 VOUT-.t1 GNDA 0.04876f
C1999 VOUT-.t4 GNDA 0.04876f
C2000 VOUT-.n87 GNDA 0.22561f
C2001 VOUT-.n88 GNDA 0.138742f
C2002 VOUT-.t11 GNDA 0.04876f
C2003 VOUT-.t7 GNDA 0.04876f
C2004 VOUT-.n89 GNDA 0.22561f
C2005 VOUT-.n90 GNDA 0.077288f
C2006 VOUT-.t18 GNDA 0.081164f
C2007 VOUT-.n91 GNDA 0.089334f
C2008 bgr_7_0.V_TOP.t24 GNDA 0.095448f
C2009 bgr_7_0.V_TOP.t33 GNDA 0.095448f
C2010 bgr_7_0.V_TOP.t39 GNDA 0.095448f
C2011 bgr_7_0.V_TOP.t16 GNDA 0.095448f
C2012 bgr_7_0.V_TOP.t15 GNDA 0.095448f
C2013 bgr_7_0.V_TOP.t28 GNDA 0.095448f
C2014 bgr_7_0.V_TOP.t38 GNDA 0.095448f
C2015 bgr_7_0.V_TOP.t14 GNDA 0.095448f
C2016 bgr_7_0.V_TOP.t27 GNDA 0.095448f
C2017 bgr_7_0.V_TOP.t26 GNDA 0.095448f
C2018 bgr_7_0.V_TOP.t37 GNDA 0.095448f
C2019 bgr_7_0.V_TOP.t46 GNDA 0.095448f
C2020 bgr_7_0.V_TOP.t18 GNDA 0.095448f
C2021 bgr_7_0.V_TOP.t30 GNDA 0.095448f
C2022 bgr_7_0.V_TOP.t29 GNDA 0.124774f
C2023 bgr_7_0.V_TOP.n0 GNDA 0.069758f
C2024 bgr_7_0.V_TOP.n1 GNDA 0.050905f
C2025 bgr_7_0.V_TOP.n2 GNDA 0.050905f
C2026 bgr_7_0.V_TOP.n3 GNDA 0.050905f
C2027 bgr_7_0.V_TOP.n4 GNDA 0.050905f
C2028 bgr_7_0.V_TOP.n5 GNDA 0.04747f
C2029 bgr_7_0.V_TOP.t10 GNDA 0.122745f
C2030 bgr_7_0.V_TOP.t40 GNDA 0.36361f
C2031 bgr_7_0.V_TOP.t31 GNDA 0.369803f
C2032 bgr_7_0.V_TOP.t35 GNDA 0.36361f
C2033 bgr_7_0.V_TOP.n6 GNDA 0.243789f
C2034 bgr_7_0.V_TOP.t32 GNDA 0.36361f
C2035 bgr_7_0.V_TOP.t22 GNDA 0.369803f
C2036 bgr_7_0.V_TOP.n7 GNDA 0.311966f
C2037 bgr_7_0.V_TOP.t20 GNDA 0.369803f
C2038 bgr_7_0.V_TOP.t25 GNDA 0.36361f
C2039 bgr_7_0.V_TOP.n8 GNDA 0.243789f
C2040 bgr_7_0.V_TOP.t21 GNDA 0.36361f
C2041 bgr_7_0.V_TOP.t45 GNDA 0.369803f
C2042 bgr_7_0.V_TOP.n9 GNDA 0.380142f
C2043 bgr_7_0.V_TOP.t42 GNDA 0.369803f
C2044 bgr_7_0.V_TOP.t49 GNDA 0.36361f
C2045 bgr_7_0.V_TOP.n10 GNDA 0.243789f
C2046 bgr_7_0.V_TOP.t44 GNDA 0.36361f
C2047 bgr_7_0.V_TOP.t36 GNDA 0.369803f
C2048 bgr_7_0.V_TOP.n11 GNDA 0.380142f
C2049 bgr_7_0.V_TOP.t17 GNDA 0.369803f
C2050 bgr_7_0.V_TOP.t23 GNDA 0.36361f
C2051 bgr_7_0.V_TOP.n12 GNDA 0.243789f
C2052 bgr_7_0.V_TOP.t19 GNDA 0.36361f
C2053 bgr_7_0.V_TOP.t43 GNDA 0.369803f
C2054 bgr_7_0.V_TOP.n13 GNDA 0.380142f
C2055 bgr_7_0.V_TOP.t34 GNDA 0.369803f
C2056 bgr_7_0.V_TOP.t41 GNDA 0.36361f
C2057 bgr_7_0.V_TOP.n14 GNDA 0.311966f
C2058 bgr_7_0.V_TOP.t47 GNDA 0.36361f
C2059 bgr_7_0.V_TOP.n15 GNDA 0.159079f
C2060 bgr_7_0.V_TOP.n16 GNDA 0.544408f
C2061 bgr_7_0.V_TOP.t0 GNDA 0.102288f
C2062 bgr_7_0.V_TOP.n17 GNDA 0.724299f
C2063 bgr_7_0.V_TOP.n18 GNDA 0.022634f
C2064 bgr_7_0.V_TOP.n19 GNDA 0.414649f
C2065 bgr_7_0.V_TOP.n20 GNDA 0.021924f
C2066 bgr_7_0.V_TOP.n21 GNDA 0.022786f
C2067 bgr_7_0.V_TOP.n22 GNDA 0.022634f
C2068 bgr_7_0.V_TOP.n23 GNDA 0.209756f
C2069 bgr_7_0.V_TOP.n24 GNDA 0.127416f
C2070 bgr_7_0.V_TOP.n25 GNDA 0.072722f
C2071 bgr_7_0.V_TOP.n26 GNDA 0.022634f
C2072 bgr_7_0.V_TOP.n27 GNDA 0.125537f
C2073 bgr_7_0.V_TOP.n28 GNDA 0.022634f
C2074 bgr_7_0.V_TOP.n29 GNDA 0.124344f
C2075 bgr_7_0.V_TOP.n30 GNDA 0.273328f
C2076 bgr_7_0.V_TOP.n31 GNDA 0.019234f
C2077 bgr_7_0.V_TOP.n32 GNDA 0.04747f
C2078 bgr_7_0.V_TOP.n33 GNDA 0.050905f
C2079 bgr_7_0.V_TOP.n34 GNDA 0.050905f
C2080 bgr_7_0.V_TOP.n35 GNDA 0.050905f
C2081 bgr_7_0.V_TOP.n36 GNDA 0.050905f
C2082 bgr_7_0.V_TOP.n37 GNDA 0.050905f
C2083 bgr_7_0.V_TOP.n38 GNDA 0.050905f
C2084 bgr_7_0.V_TOP.n39 GNDA 0.04747f
C2085 bgr_7_0.V_TOP.t48 GNDA 0.109989f
C2086 VDDA.t319 GNDA 0.02154f
C2087 VDDA.t329 GNDA 0.02154f
C2088 VDDA.n0 GNDA 0.074646f
C2089 VDDA.n1 GNDA 0.073056f
C2090 VDDA.t196 GNDA 0.02154f
C2091 VDDA.n2 GNDA 0.06462f
C2092 VDDA.n3 GNDA 0.02154f
C2093 VDDA.n4 GNDA 0.012309f
C2094 VDDA.n8 GNDA 0.012309f
C2095 VDDA.t250 GNDA 0.037766f
C2096 VDDA.t351 GNDA 0.02154f
C2097 VDDA.t355 GNDA 0.02154f
C2098 VDDA.n9 GNDA 0.074646f
C2099 VDDA.n10 GNDA 0.093535f
C2100 VDDA.n11 GNDA 0.032075f
C2101 VDDA.n12 GNDA 0.02154f
C2102 VDDA.n14 GNDA 0.02154f
C2103 VDDA.n15 GNDA 0.012309f
C2104 VDDA.n16 GNDA 0.012309f
C2105 VDDA.n17 GNDA 0.02154f
C2106 VDDA.n19 GNDA 0.02154f
C2107 VDDA.n20 GNDA 0.012309f
C2108 VDDA.n21 GNDA 0.012309f
C2109 VDDA.n22 GNDA 0.02154f
C2110 VDDA.n23 GNDA 0.021728f
C2111 VDDA.t252 GNDA 0.02154f
C2112 VDDA.n24 GNDA 0.06462f
C2113 VDDA.n25 GNDA 0.020764f
C2114 VDDA.n26 GNDA 0.012309f
C2115 VDDA.n27 GNDA 0.180012f
C2116 VDDA.t251 GNDA 0.15601f
C2117 VDDA.t350 GNDA 0.144009f
C2118 VDDA.t354 GNDA 0.144009f
C2119 VDDA.t318 GNDA 0.144009f
C2120 VDDA.t328 GNDA 0.144009f
C2121 VDDA.t324 GNDA 0.144009f
C2122 VDDA.t332 GNDA 0.144009f
C2123 VDDA.t340 GNDA 0.144009f
C2124 VDDA.t346 GNDA 0.144009f
C2125 VDDA.t322 GNDA 0.144009f
C2126 VDDA.t316 GNDA 0.144009f
C2127 VDDA.t195 GNDA 0.15601f
C2128 VDDA.n30 GNDA 0.012309f
C2129 VDDA.n32 GNDA 0.021728f
C2130 VDDA.n33 GNDA 0.02154f
C2131 VDDA.n34 GNDA 0.012309f
C2132 VDDA.n35 GNDA 0.012309f
C2133 VDDA.n36 GNDA 0.02154f
C2134 VDDA.n38 GNDA 0.02154f
C2135 VDDA.n39 GNDA 0.02154f
C2136 VDDA.n40 GNDA 0.012309f
C2137 VDDA.n41 GNDA 0.180012f
C2138 VDDA.n43 GNDA 0.02352f
C2139 VDDA.t194 GNDA 0.037766f
C2140 VDDA.n44 GNDA 0.032075f
C2141 VDDA.t323 GNDA 0.02154f
C2142 VDDA.t317 GNDA 0.02154f
C2143 VDDA.n45 GNDA 0.074646f
C2144 VDDA.n46 GNDA 0.093535f
C2145 VDDA.t341 GNDA 0.02154f
C2146 VDDA.t347 GNDA 0.02154f
C2147 VDDA.n47 GNDA 0.074646f
C2148 VDDA.n48 GNDA 0.073056f
C2149 VDDA.n49 GNDA 0.019694f
C2150 VDDA.t325 GNDA 0.02154f
C2151 VDDA.t333 GNDA 0.02154f
C2152 VDDA.n50 GNDA 0.073099f
C2153 VDDA.n51 GNDA 0.08421f
C2154 VDDA.t359 GNDA 0.018463f
C2155 VDDA.t78 GNDA 0.018463f
C2156 VDDA.n52 GNDA 0.076351f
C2157 VDDA.t112 GNDA 0.018463f
C2158 VDDA.t389 GNDA 0.018463f
C2159 VDDA.n53 GNDA 0.076058f
C2160 VDDA.n54 GNDA 0.105454f
C2161 VDDA.t117 GNDA 0.018463f
C2162 VDDA.t126 GNDA 0.018463f
C2163 VDDA.n55 GNDA 0.076058f
C2164 VDDA.n56 GNDA 0.055027f
C2165 VDDA.t374 GNDA 0.018463f
C2166 VDDA.t127 GNDA 0.018463f
C2167 VDDA.n57 GNDA 0.076058f
C2168 VDDA.n58 GNDA 0.055027f
C2169 VDDA.t32 GNDA 0.018463f
C2170 VDDA.t63 GNDA 0.018463f
C2171 VDDA.n59 GNDA 0.076058f
C2172 VDDA.n60 GNDA 0.055027f
C2173 VDDA.t147 GNDA 0.018463f
C2174 VDDA.t360 GNDA 0.018463f
C2175 VDDA.n61 GNDA 0.076058f
C2176 VDDA.n62 GNDA 0.111004f
C2177 VDDA.t203 GNDA 0.018605f
C2178 VDDA.n64 GNDA 0.012309f
C2179 VDDA.n65 GNDA 0.010117f
C2180 VDDA.n66 GNDA 0.012309f
C2181 VDDA.t188 GNDA 0.019444f
C2182 VDDA.n67 GNDA 0.02154f
C2183 VDDA.n68 GNDA 0.012309f
C2184 VDDA.n69 GNDA 0.02154f
C2185 VDDA.n70 GNDA 0.029969f
C2186 VDDA.t190 GNDA 0.032451f
C2187 VDDA.n72 GNDA 0.04927f
C2188 VDDA.n74 GNDA 0.10893f
C2189 VDDA.t189 GNDA 0.090467f
C2190 VDDA.t386 GNDA 0.081236f
C2191 VDDA.t395 GNDA 0.081236f
C2192 VDDA.t138 GNDA 0.081236f
C2193 VDDA.t398 GNDA 0.081236f
C2194 VDDA.t294 GNDA 0.081236f
C2195 VDDA.t405 GNDA 0.081236f
C2196 VDDA.t116 GNDA 0.081236f
C2197 VDDA.t404 GNDA 0.081236f
C2198 VDDA.t131 GNDA 0.081236f
C2199 VDDA.t295 GNDA 0.081236f
C2200 VDDA.t204 GNDA 0.090467f
C2201 VDDA.n76 GNDA 0.012309f
C2202 VDDA.n77 GNDA 0.02154f
C2203 VDDA.n78 GNDA 0.02154f
C2204 VDDA.t205 GNDA 0.032451f
C2205 VDDA.n79 GNDA 0.027132f
C2206 VDDA.n80 GNDA 0.012954f
C2207 VDDA.n81 GNDA 0.10893f
C2208 VDDA.n82 GNDA 0.012309f
C2209 VDDA.n83 GNDA 0.024411f
C2210 VDDA.n84 GNDA 0.039446f
C2211 VDDA.n85 GNDA 0.173383f
C2212 VDDA.t15 GNDA 0.036925f
C2213 VDDA.t367 GNDA 0.036925f
C2214 VDDA.n86 GNDA 0.14814f
C2215 VDDA.n87 GNDA 0.075259f
C2216 VDDA.n89 GNDA 0.012309f
C2217 VDDA.n95 GNDA 0.012954f
C2218 VDDA.n96 GNDA 0.012309f
C2219 VDDA.t262 GNDA 0.044741f
C2220 VDDA.t369 GNDA 0.036925f
C2221 VDDA.t149 GNDA 0.036925f
C2222 VDDA.n97 GNDA 0.14814f
C2223 VDDA.n98 GNDA 0.075259f
C2224 VDDA.t133 GNDA 0.036925f
C2225 VDDA.t383 GNDA 0.036925f
C2226 VDDA.n99 GNDA 0.14814f
C2227 VDDA.n100 GNDA 0.075259f
C2228 VDDA.t385 GNDA 0.036925f
C2229 VDDA.t388 GNDA 0.036925f
C2230 VDDA.n101 GNDA 0.14814f
C2231 VDDA.n102 GNDA 0.075259f
C2232 VDDA.t62 GNDA 0.036925f
C2233 VDDA.t397 GNDA 0.036925f
C2234 VDDA.n103 GNDA 0.14814f
C2235 VDDA.n104 GNDA 0.095235f
C2236 VDDA.n105 GNDA 0.036834f
C2237 VDDA.n106 GNDA 0.024488f
C2238 VDDA.n107 GNDA 0.012309f
C2239 VDDA.n108 GNDA 0.012309f
C2240 VDDA.n109 GNDA 0.02154f
C2241 VDDA.n110 GNDA 0.012309f
C2242 VDDA.n111 GNDA 0.012309f
C2243 VDDA.n112 GNDA 0.012309f
C2244 VDDA.n113 GNDA 0.012309f
C2245 VDDA.n114 GNDA 0.02154f
C2246 VDDA.n115 GNDA 0.024488f
C2247 VDDA.n116 GNDA 0.012309f
C2248 VDDA.n117 GNDA 0.012309f
C2249 VDDA.n118 GNDA 0.012309f
C2250 VDDA.n119 GNDA 0.031178f
C2251 VDDA.n120 GNDA 0.02154f
C2252 VDDA.n121 GNDA 0.02154f
C2253 VDDA.n122 GNDA 0.02154f
C2254 VDDA.n123 GNDA 0.012309f
C2255 VDDA.n124 GNDA 0.012309f
C2256 VDDA.n126 GNDA 0.02154f
C2257 VDDA.n127 GNDA 0.02154f
C2258 VDDA.n129 GNDA 0.012309f
C2259 VDDA.n130 GNDA 0.012309f
C2260 VDDA.n131 GNDA 0.02154f
C2261 VDDA.n132 GNDA 0.02154f
C2262 VDDA.n133 GNDA 0.02154f
C2263 VDDA.n135 GNDA 0.024411f
C2264 VDDA.n136 GNDA 0.012309f
C2265 VDDA.n137 GNDA 0.290481f
C2266 VDDA.t263 GNDA 0.241247f
C2267 VDDA.t61 GNDA 0.21663f
C2268 VDDA.t396 GNDA 0.21663f
C2269 VDDA.t384 GNDA 0.21663f
C2270 VDDA.t387 GNDA 0.21663f
C2271 VDDA.t132 GNDA 0.21663f
C2272 VDDA.t382 GNDA 0.21663f
C2273 VDDA.t368 GNDA 0.21663f
C2274 VDDA.t148 GNDA 0.21663f
C2275 VDDA.t14 GNDA 0.21663f
C2276 VDDA.t366 GNDA 0.21663f
C2277 VDDA.t275 GNDA 0.241247f
C2278 VDDA.n142 GNDA 0.012954f
C2279 VDDA.n143 GNDA 0.012309f
C2280 VDDA.n144 GNDA 0.02154f
C2281 VDDA.n145 GNDA 0.024488f
C2282 VDDA.n146 GNDA 0.012309f
C2283 VDDA.n147 GNDA 0.012309f
C2284 VDDA.n150 GNDA 0.012309f
C2285 VDDA.n151 GNDA 0.012309f
C2286 VDDA.n152 GNDA 0.024488f
C2287 VDDA.n153 GNDA 0.031178f
C2288 VDDA.n154 GNDA 0.012309f
C2289 VDDA.n155 GNDA 0.02154f
C2290 VDDA.n156 GNDA 0.02154f
C2291 VDDA.n157 GNDA 0.012309f
C2292 VDDA.n158 GNDA 0.012309f
C2293 VDDA.n159 GNDA 0.02154f
C2294 VDDA.n160 GNDA 0.02154f
C2295 VDDA.n161 GNDA 0.012309f
C2296 VDDA.n162 GNDA 0.012309f
C2297 VDDA.n163 GNDA 0.02154f
C2298 VDDA.n164 GNDA 0.02154f
C2299 VDDA.n165 GNDA 0.012309f
C2300 VDDA.n166 GNDA 0.012309f
C2301 VDDA.n167 GNDA 0.02154f
C2302 VDDA.n168 GNDA 0.02154f
C2303 VDDA.n169 GNDA 0.02154f
C2304 VDDA.n170 GNDA 0.012309f
C2305 VDDA.n171 GNDA 0.290481f
C2306 VDDA.n173 GNDA 0.027166f
C2307 VDDA.t274 GNDA 0.044741f
C2308 VDDA.n174 GNDA 0.03602f
C2309 VDDA.n175 GNDA 0.050069f
C2310 VDDA.n176 GNDA 0.066112f
C2311 VDDA.t381 GNDA 0.015386f
C2312 VDDA.t158 GNDA 0.015386f
C2313 VDDA.n177 GNDA 0.053052f
C2314 VDDA.n178 GNDA 0.068604f
C2315 VDDA.t288 GNDA 0.015386f
C2316 VDDA.n179 GNDA 0.046157f
C2317 VDDA.n180 GNDA 0.02154f
C2318 VDDA.n181 GNDA 0.012309f
C2319 VDDA.t239 GNDA 0.109315f
C2320 VDDA.n184 GNDA 0.012309f
C2321 VDDA.n185 GNDA 0.012309f
C2322 VDDA.t210 GNDA 0.02312f
C2323 VDDA.n186 GNDA 0.03154f
C2324 VDDA.n187 GNDA 0.026736f
C2325 VDDA.t241 GNDA 0.02312f
C2326 VDDA.t243 GNDA 0.015386f
C2327 VDDA.n188 GNDA 0.046157f
C2328 VDDA.n189 GNDA 0.02154f
C2329 VDDA.n190 GNDA 0.012309f
C2330 VDDA.t0 GNDA 0.09816f
C2331 VDDA.t18 GNDA 0.09816f
C2332 VDDA.t308 GNDA 0.09816f
C2333 VDDA.t411 GNDA 0.09816f
C2334 VDDA.t242 GNDA 0.109315f
C2335 VDDA.n192 GNDA 0.012309f
C2336 VDDA.n194 GNDA 0.012309f
C2337 VDDA.n195 GNDA 0.02154f
C2338 VDDA.n196 GNDA 0.02154f
C2339 VDDA.n197 GNDA 0.021728f
C2340 VDDA.n199 GNDA 0.131624f
C2341 VDDA.n200 GNDA 0.012309f
C2342 VDDA.n201 GNDA 0.023599f
C2343 VDDA.n202 GNDA 0.033709f
C2344 VDDA.t19 GNDA 0.015386f
C2345 VDDA.t309 GNDA 0.015386f
C2346 VDDA.n203 GNDA 0.053052f
C2347 VDDA.n204 GNDA 0.091359f
C2348 VDDA.n205 GNDA 0.026736f
C2349 VDDA.t238 GNDA 0.02312f
C2350 VDDA.n206 GNDA 0.03154f
C2351 VDDA.n207 GNDA 0.016493f
C2352 VDDA.t212 GNDA 0.015386f
C2353 VDDA.n209 GNDA 0.033848f
C2354 VDDA.n211 GNDA 0.012309f
C2355 VDDA.n212 GNDA 0.033848f
C2356 VDDA.n213 GNDA 0.033848f
C2357 VDDA.t240 GNDA 0.015386f
C2358 VDDA.n215 GNDA 0.046157f
C2359 VDDA.n216 GNDA 0.033219f
C2360 VDDA.n218 GNDA 0.046157f
C2361 VDDA.n219 GNDA 0.026449f
C2362 VDDA.n221 GNDA 0.120469f
C2363 VDDA.t211 GNDA 0.109315f
C2364 VDDA.t3 GNDA 0.09816f
C2365 VDDA.t157 GNDA 0.09816f
C2366 VDDA.t380 GNDA 0.09816f
C2367 VDDA.t67 GNDA 0.09816f
C2368 VDDA.t287 GNDA 0.109315f
C2369 VDDA.n222 GNDA 0.012309f
C2370 VDDA.n224 GNDA 0.021728f
C2371 VDDA.n225 GNDA 0.02154f
C2372 VDDA.n226 GNDA 0.02154f
C2373 VDDA.n227 GNDA 0.012309f
C2374 VDDA.n228 GNDA 0.131624f
C2375 VDDA.n230 GNDA 0.026354f
C2376 VDDA.t286 GNDA 0.02312f
C2377 VDDA.n231 GNDA 0.032189f
C2378 VDDA.n232 GNDA 0.090099f
C2379 VDDA.n233 GNDA 0.098176f
C2380 VDDA.n234 GNDA 0.151029f
C2381 VDDA.t345 GNDA 0.02154f
C2382 VDDA.t353 GNDA 0.02154f
C2383 VDDA.n235 GNDA 0.074646f
C2384 VDDA.n236 GNDA 0.073056f
C2385 VDDA.t237 GNDA 0.02154f
C2386 VDDA.n237 GNDA 0.06462f
C2387 VDDA.n238 GNDA 0.02154f
C2388 VDDA.n239 GNDA 0.012309f
C2389 VDDA.n243 GNDA 0.012309f
C2390 VDDA.t179 GNDA 0.037766f
C2391 VDDA.t327 GNDA 0.02154f
C2392 VDDA.t337 GNDA 0.02154f
C2393 VDDA.n244 GNDA 0.074646f
C2394 VDDA.n245 GNDA 0.093535f
C2395 VDDA.n246 GNDA 0.032075f
C2396 VDDA.n247 GNDA 0.02154f
C2397 VDDA.n249 GNDA 0.02154f
C2398 VDDA.n250 GNDA 0.012309f
C2399 VDDA.n251 GNDA 0.012309f
C2400 VDDA.n252 GNDA 0.02154f
C2401 VDDA.n254 GNDA 0.02154f
C2402 VDDA.n255 GNDA 0.012309f
C2403 VDDA.n256 GNDA 0.012309f
C2404 VDDA.n257 GNDA 0.02154f
C2405 VDDA.n258 GNDA 0.021728f
C2406 VDDA.t181 GNDA 0.02154f
C2407 VDDA.n259 GNDA 0.06462f
C2408 VDDA.n260 GNDA 0.020764f
C2409 VDDA.n261 GNDA 0.012309f
C2410 VDDA.n262 GNDA 0.180012f
C2411 VDDA.t180 GNDA 0.15601f
C2412 VDDA.t326 GNDA 0.144009f
C2413 VDDA.t336 GNDA 0.144009f
C2414 VDDA.t344 GNDA 0.144009f
C2415 VDDA.t352 GNDA 0.144009f
C2416 VDDA.t356 GNDA 0.144009f
C2417 VDDA.t320 GNDA 0.144009f
C2418 VDDA.t330 GNDA 0.144009f
C2419 VDDA.t338 GNDA 0.144009f
C2420 VDDA.t334 GNDA 0.144009f
C2421 VDDA.t342 GNDA 0.144009f
C2422 VDDA.t236 GNDA 0.15601f
C2423 VDDA.n265 GNDA 0.012309f
C2424 VDDA.n267 GNDA 0.021728f
C2425 VDDA.n268 GNDA 0.02154f
C2426 VDDA.n269 GNDA 0.012309f
C2427 VDDA.n270 GNDA 0.012309f
C2428 VDDA.n271 GNDA 0.02154f
C2429 VDDA.n273 GNDA 0.02154f
C2430 VDDA.n274 GNDA 0.02154f
C2431 VDDA.n275 GNDA 0.012309f
C2432 VDDA.n276 GNDA 0.180012f
C2433 VDDA.n278 GNDA 0.02352f
C2434 VDDA.t235 GNDA 0.037766f
C2435 VDDA.n279 GNDA 0.032075f
C2436 VDDA.t335 GNDA 0.02154f
C2437 VDDA.t343 GNDA 0.02154f
C2438 VDDA.n280 GNDA 0.074646f
C2439 VDDA.n281 GNDA 0.093535f
C2440 VDDA.t331 GNDA 0.02154f
C2441 VDDA.t339 GNDA 0.02154f
C2442 VDDA.n282 GNDA 0.074646f
C2443 VDDA.n283 GNDA 0.073056f
C2444 VDDA.n284 GNDA 0.019694f
C2445 VDDA.t357 GNDA 0.02154f
C2446 VDDA.t321 GNDA 0.02154f
C2447 VDDA.n285 GNDA 0.073099f
C2448 VDDA.n286 GNDA 0.08421f
C2449 VDDA.t377 GNDA 0.018463f
C2450 VDDA.t358 GNDA 0.018463f
C2451 VDDA.n287 GNDA 0.076351f
C2452 VDDA.t401 GNDA 0.018463f
C2453 VDDA.t121 GNDA 0.018463f
C2454 VDDA.n288 GNDA 0.076058f
C2455 VDDA.n289 GNDA 0.105454f
C2456 VDDA.t106 GNDA 0.018463f
C2457 VDDA.t139 GNDA 0.018463f
C2458 VDDA.n290 GNDA 0.076058f
C2459 VDDA.n291 GNDA 0.055027f
C2460 VDDA.t94 GNDA 0.018463f
C2461 VDDA.t391 GNDA 0.018463f
C2462 VDDA.n292 GNDA 0.076058f
C2463 VDDA.n293 GNDA 0.055027f
C2464 VDDA.t84 GNDA 0.018463f
C2465 VDDA.t390 GNDA 0.018463f
C2466 VDDA.n294 GNDA 0.076058f
C2467 VDDA.n295 GNDA 0.055027f
C2468 VDDA.t361 GNDA 0.018463f
C2469 VDDA.t170 GNDA 0.018463f
C2470 VDDA.n296 GNDA 0.076058f
C2471 VDDA.n297 GNDA 0.111004f
C2472 VDDA.t247 GNDA 0.018605f
C2473 VDDA.n298 GNDA 0.012309f
C2474 VDDA.t249 GNDA 0.032451f
C2475 VDDA.n299 GNDA 0.012309f
C2476 VDDA.n300 GNDA 0.012309f
C2477 VDDA.n302 GNDA 0.010117f
C2478 VDDA.n303 GNDA 0.012309f
C2479 VDDA.t259 GNDA 0.019444f
C2480 VDDA.n304 GNDA 0.02154f
C2481 VDDA.n305 GNDA 0.012309f
C2482 VDDA.n306 GNDA 0.02154f
C2483 VDDA.n307 GNDA 0.029969f
C2484 VDDA.t261 GNDA 0.032451f
C2485 VDDA.n309 GNDA 0.04927f
C2486 VDDA.n311 GNDA 0.10893f
C2487 VDDA.t260 GNDA 0.090467f
C2488 VDDA.t64 GNDA 0.081236f
C2489 VDDA.t392 GNDA 0.081236f
C2490 VDDA.t406 GNDA 0.081236f
C2491 VDDA.t79 GNDA 0.081236f
C2492 VDDA.t140 GNDA 0.081236f
C2493 VDDA.t56 GNDA 0.081236f
C2494 VDDA.t130 GNDA 0.081236f
C2495 VDDA.t120 GNDA 0.081236f
C2496 VDDA.t171 GNDA 0.081236f
C2497 VDDA.t115 GNDA 0.081236f
C2498 VDDA.t248 GNDA 0.090467f
C2499 VDDA.n312 GNDA 0.10893f
C2500 VDDA.n313 GNDA 0.012954f
C2501 VDDA.n314 GNDA 0.027132f
C2502 VDDA.n315 GNDA 0.02154f
C2503 VDDA.n316 GNDA 0.02154f
C2504 VDDA.n318 GNDA 0.024411f
C2505 VDDA.n319 GNDA 0.039446f
C2506 VDDA.n320 GNDA 0.173383f
C2507 VDDA.t17 GNDA 0.036925f
C2508 VDDA.t114 GNDA 0.036925f
C2509 VDDA.n321 GNDA 0.14814f
C2510 VDDA.n322 GNDA 0.075259f
C2511 VDDA.n324 GNDA 0.012309f
C2512 VDDA.n329 GNDA 0.012954f
C2513 VDDA.n335 GNDA 0.012954f
C2514 VDDA.n336 GNDA 0.012309f
C2515 VDDA.t213 GNDA 0.044741f
C2516 VDDA.t129 GNDA 0.036925f
C2517 VDDA.t400 GNDA 0.036925f
C2518 VDDA.n337 GNDA 0.14814f
C2519 VDDA.n338 GNDA 0.075259f
C2520 VDDA.t55 GNDA 0.036925f
C2521 VDDA.t119 GNDA 0.036925f
C2522 VDDA.n339 GNDA 0.14814f
C2523 VDDA.n340 GNDA 0.075259f
C2524 VDDA.t142 GNDA 0.036925f
C2525 VDDA.t36 GNDA 0.036925f
C2526 VDDA.n341 GNDA 0.14814f
C2527 VDDA.n342 GNDA 0.075259f
C2528 VDDA.t408 GNDA 0.036925f
C2529 VDDA.t123 GNDA 0.036925f
C2530 VDDA.n343 GNDA 0.14814f
C2531 VDDA.n344 GNDA 0.095235f
C2532 VDDA.n345 GNDA 0.036834f
C2533 VDDA.n346 GNDA 0.02154f
C2534 VDDA.n347 GNDA 0.012309f
C2535 VDDA.n348 GNDA 0.012309f
C2536 VDDA.n351 GNDA 0.012309f
C2537 VDDA.n352 GNDA 0.012309f
C2538 VDDA.n353 GNDA 0.024488f
C2539 VDDA.n354 GNDA 0.031178f
C2540 VDDA.n355 GNDA 0.012309f
C2541 VDDA.n356 GNDA 0.02154f
C2542 VDDA.n357 GNDA 0.02154f
C2543 VDDA.n358 GNDA 0.012309f
C2544 VDDA.n359 GNDA 0.012309f
C2545 VDDA.n360 GNDA 0.02154f
C2546 VDDA.n361 GNDA 0.02154f
C2547 VDDA.n362 GNDA 0.012309f
C2548 VDDA.n363 GNDA 0.012309f
C2549 VDDA.n364 GNDA 0.02154f
C2550 VDDA.n365 GNDA 0.02154f
C2551 VDDA.n366 GNDA 0.012309f
C2552 VDDA.n367 GNDA 0.012309f
C2553 VDDA.n368 GNDA 0.02154f
C2554 VDDA.n369 GNDA 0.02154f
C2555 VDDA.n370 GNDA 0.012309f
C2556 VDDA.n371 GNDA 0.012309f
C2557 VDDA.n372 GNDA 0.02154f
C2558 VDDA.n373 GNDA 0.024488f
C2559 VDDA.n375 GNDA 0.024411f
C2560 VDDA.n376 GNDA 0.012309f
C2561 VDDA.n377 GNDA 0.290481f
C2562 VDDA.t214 GNDA 0.241247f
C2563 VDDA.t122 GNDA 0.21663f
C2564 VDDA.t407 GNDA 0.21663f
C2565 VDDA.t35 GNDA 0.21663f
C2566 VDDA.t141 GNDA 0.21663f
C2567 VDDA.t118 GNDA 0.21663f
C2568 VDDA.t54 GNDA 0.21663f
C2569 VDDA.t399 GNDA 0.21663f
C2570 VDDA.t128 GNDA 0.21663f
C2571 VDDA.t113 GNDA 0.21663f
C2572 VDDA.t16 GNDA 0.21663f
C2573 VDDA.t192 GNDA 0.241247f
C2574 VDDA.n378 GNDA 0.012309f
C2575 VDDA.n379 GNDA 0.02154f
C2576 VDDA.n380 GNDA 0.024488f
C2577 VDDA.n381 GNDA 0.012309f
C2578 VDDA.n382 GNDA 0.012309f
C2579 VDDA.n385 GNDA 0.012309f
C2580 VDDA.n386 GNDA 0.012309f
C2581 VDDA.n387 GNDA 0.024488f
C2582 VDDA.n388 GNDA 0.031178f
C2583 VDDA.n389 GNDA 0.012309f
C2584 VDDA.n390 GNDA 0.02154f
C2585 VDDA.n391 GNDA 0.02154f
C2586 VDDA.n392 GNDA 0.012309f
C2587 VDDA.n393 GNDA 0.012309f
C2588 VDDA.n394 GNDA 0.02154f
C2589 VDDA.n395 GNDA 0.02154f
C2590 VDDA.n396 GNDA 0.012309f
C2591 VDDA.n397 GNDA 0.012309f
C2592 VDDA.n398 GNDA 0.02154f
C2593 VDDA.n399 GNDA 0.02154f
C2594 VDDA.n400 GNDA 0.012309f
C2595 VDDA.n401 GNDA 0.012309f
C2596 VDDA.n402 GNDA 0.02154f
C2597 VDDA.n403 GNDA 0.02154f
C2598 VDDA.n404 GNDA 0.02154f
C2599 VDDA.n405 GNDA 0.012309f
C2600 VDDA.n406 GNDA 0.290481f
C2601 VDDA.n408 GNDA 0.027166f
C2602 VDDA.t191 GNDA 0.044741f
C2603 VDDA.n409 GNDA 0.03602f
C2604 VDDA.n410 GNDA 0.050069f
C2605 VDDA.n411 GNDA 0.130788f
C2606 VDDA.n412 GNDA 0.155578f
C2607 VDDA.n413 GNDA 0.144484f
C2608 VDDA.t146 GNDA 0.011078f
C2609 VDDA.t227 GNDA 0.011078f
C2610 VDDA.n414 GNDA 0.025703f
C2611 VDDA.n415 GNDA 0.083393f
C2612 VDDA.t218 GNDA 0.039304f
C2613 VDDA.t225 GNDA 0.022724f
C2614 VDDA.n416 GNDA 0.044951f
C2615 VDDA.t228 GNDA 0.039304f
C2616 VDDA.n417 GNDA 0.07379f
C2617 VDDA.t226 GNDA 0.1317f
C2618 VDDA.t145 GNDA 0.081236f
C2619 VDDA.t217 GNDA 0.1317f
C2620 VDDA.n418 GNDA 0.07379f
C2621 VDDA.t216 GNDA 0.022724f
C2622 VDDA.n419 GNDA 0.044636f
C2623 VDDA.n420 GNDA 0.041764f
C2624 VDDA.n421 GNDA 0.059172f
C2625 VDDA.n422 GNDA 0.086762f
C2626 VDDA.t282 GNDA 0.02154f
C2627 VDDA.n423 GNDA 0.06462f
C2628 VDDA.n424 GNDA 0.02154f
C2629 VDDA.n425 GNDA 0.012309f
C2630 VDDA.n429 GNDA 0.012309f
C2631 VDDA.t232 GNDA 0.037766f
C2632 VDDA.n430 GNDA 0.031462f
C2633 VDDA.n431 GNDA 0.02154f
C2634 VDDA.n433 GNDA 0.02154f
C2635 VDDA.n434 GNDA 0.012309f
C2636 VDDA.n435 GNDA 0.012309f
C2637 VDDA.n436 GNDA 0.02154f
C2638 VDDA.n438 GNDA 0.02154f
C2639 VDDA.n439 GNDA 0.012309f
C2640 VDDA.n440 GNDA 0.012309f
C2641 VDDA.n441 GNDA 0.02154f
C2642 VDDA.n442 GNDA 0.021728f
C2643 VDDA.t349 GNDA 0.02154f
C2644 VDDA.n443 GNDA 0.074646f
C2645 VDDA.t234 GNDA 0.04308f
C2646 VDDA.n444 GNDA 0.06462f
C2647 VDDA.n445 GNDA 0.020764f
C2648 VDDA.n446 GNDA 0.012309f
C2649 VDDA.n447 GNDA 0.180012f
C2650 VDDA.t233 GNDA 0.15601f
C2651 VDDA.t348 GNDA 0.144009f
C2652 VDDA.t281 GNDA 0.15601f
C2653 VDDA.n450 GNDA 0.012309f
C2654 VDDA.n452 GNDA 0.021728f
C2655 VDDA.n453 GNDA 0.02154f
C2656 VDDA.n454 GNDA 0.012309f
C2657 VDDA.n455 GNDA 0.012309f
C2658 VDDA.n456 GNDA 0.02154f
C2659 VDDA.n458 GNDA 0.02154f
C2660 VDDA.n459 GNDA 0.02154f
C2661 VDDA.n460 GNDA 0.012309f
C2662 VDDA.n461 GNDA 0.180012f
C2663 VDDA.n463 GNDA 0.02352f
C2664 VDDA.t280 GNDA 0.037766f
C2665 VDDA.n464 GNDA 0.031147f
C2666 VDDA.n465 GNDA 0.041764f
C2667 VDDA.n466 GNDA 0.17463f
C2668 VDDA.n467 GNDA 3.30688f
C2669 VDDA.t104 GNDA 0.344023f
C2670 VDDA.t169 GNDA 0.345269f
C2671 VDDA.t12 GNDA 0.326807f
C2672 VDDA.t77 GNDA 0.344023f
C2673 VDDA.t152 GNDA 0.345269f
C2674 VDDA.t46 GNDA 0.326807f
C2675 VDDA.t45 GNDA 0.344023f
C2676 VDDA.t101 GNDA 0.345269f
C2677 VDDA.t87 GNDA 0.326807f
C2678 VDDA.t156 GNDA 0.344023f
C2679 VDDA.t70 GNDA 0.345269f
C2680 VDDA.t166 GNDA 0.326807f
C2681 VDDA.t306 GNDA 0.344023f
C2682 VDDA.t13 GNDA 0.345269f
C2683 VDDA.t151 GNDA 0.326807f
C2684 VDDA.n468 GNDA 0.230599f
C2685 VDDA.t307 GNDA 0.183638f
C2686 VDDA.n469 GNDA 0.250205f
C2687 VDDA.t150 GNDA 0.183638f
C2688 VDDA.n470 GNDA 0.250205f
C2689 VDDA.t47 GNDA 0.183638f
C2690 VDDA.n471 GNDA 0.250205f
C2691 VDDA.t155 GNDA 0.183638f
C2692 VDDA.n472 GNDA 0.250205f
C2693 VDDA.t105 GNDA 0.321703f
C2694 VDDA.n473 GNDA 2.85702f
C2695 VDDA.t412 GNDA 0.680378f
C2696 VDDA.t414 GNDA 0.725153f
C2697 VDDA.t415 GNDA 0.724869f
C2698 VDDA.t413 GNDA 0.697582f
C2699 VDDA.n474 GNDA 0.485588f
C2700 VDDA.n475 GNDA 0.238462f
C2701 VDDA.n476 GNDA 0.346623f
C2702 VDDA.n477 GNDA 0.632719f
C2703 VDDA.n478 GNDA 0.015479f
C2704 VDDA.n479 GNDA 0.06268f
C2705 VDDA.n480 GNDA 0.026027f
C2706 VDDA.t231 GNDA 0.021407f
C2707 VDDA.n482 GNDA 0.026027f
C2708 VDDA.n483 GNDA 0.015479f
C2709 VDDA.n484 GNDA 0.06268f
C2710 VDDA.t224 GNDA 0.021556f
C2711 VDDA.n485 GNDA 0.026027f
C2712 VDDA.n486 GNDA 0.015479f
C2713 VDDA.n487 GNDA 0.06268f
C2714 VDDA.n488 GNDA 0.015479f
C2715 VDDA.n489 GNDA 0.06268f
C2716 VDDA.n490 GNDA 0.015479f
C2717 VDDA.n491 GNDA 0.06268f
C2718 VDDA.n492 GNDA 0.015479f
C2719 VDDA.n493 GNDA 0.06268f
C2720 VDDA.n494 GNDA 0.015479f
C2721 VDDA.n495 GNDA 0.06268f
C2722 VDDA.n496 GNDA 0.015479f
C2723 VDDA.n497 GNDA 0.06268f
C2724 VDDA.n498 GNDA 0.015479f
C2725 VDDA.n499 GNDA 0.06268f
C2726 VDDA.n500 GNDA 0.015479f
C2727 VDDA.n501 GNDA 0.090075f
C2728 VDDA.n502 GNDA 0.023864f
C2729 VDDA.t197 GNDA 0.022718f
C2730 VDDA.t199 GNDA 0.021407f
C2731 VDDA.n503 GNDA 0.041033f
C2732 VDDA.n504 GNDA 0.062374f
C2733 VDDA.t198 GNDA 0.077355f
C2734 VDDA.t143 GNDA 0.051696f
C2735 VDDA.t124 GNDA 0.051696f
C2736 VDDA.t59 GNDA 0.051696f
C2737 VDDA.t107 GNDA 0.051696f
C2738 VDDA.t39 GNDA 0.051696f
C2739 VDDA.t370 GNDA 0.051696f
C2740 VDDA.t372 GNDA 0.051696f
C2741 VDDA.t136 GNDA 0.051696f
C2742 VDDA.t362 GNDA 0.051696f
C2743 VDDA.t134 GNDA 0.051696f
C2744 VDDA.t174 GNDA 0.051696f
C2745 VDDA.t97 GNDA 0.051696f
C2746 VDDA.t164 GNDA 0.051696f
C2747 VDDA.t8 GNDA 0.051696f
C2748 VDDA.t296 GNDA 0.051696f
C2749 VDDA.t37 GNDA 0.051696f
C2750 VDDA.t172 GNDA 0.051696f
C2751 VDDA.t393 GNDA 0.051696f
C2752 VDDA.t223 GNDA 0.078855f
C2753 VDDA.n505 GNDA 0.112279f
C2754 VDDA.t222 GNDA 0.015234f
C2755 VDDA.n506 GNDA 0.025175f
C2756 VDDA.n507 GNDA 0.045844f
C2757 VDDA.n508 GNDA 0.015479f
C2758 VDDA.n509 GNDA 0.06268f
C2759 VDDA.n510 GNDA 0.015479f
C2760 VDDA.n511 GNDA 0.06268f
C2761 VDDA.n512 GNDA 0.015479f
C2762 VDDA.n513 GNDA 0.06268f
C2763 VDDA.n514 GNDA 0.015479f
C2764 VDDA.n515 GNDA 0.06268f
C2765 VDDA.n516 GNDA 0.015479f
C2766 VDDA.n517 GNDA 0.06268f
C2767 VDDA.n518 GNDA 0.015479f
C2768 VDDA.n519 GNDA 0.06268f
C2769 VDDA.n520 GNDA 0.015479f
C2770 VDDA.n521 GNDA 0.06268f
C2771 VDDA.n522 GNDA 0.015479f
C2772 VDDA.n523 GNDA 0.06268f
C2773 VDDA.n524 GNDA 0.045844f
C2774 VDDA.n525 GNDA 0.022647f
C2775 VDDA.t256 GNDA 0.022718f
C2776 VDDA.t258 GNDA 0.021407f
C2777 VDDA.n526 GNDA 0.041033f
C2778 VDDA.n527 GNDA 0.062374f
C2779 VDDA.t257 GNDA 0.077355f
C2780 VDDA.t375 GNDA 0.051696f
C2781 VDDA.t162 GNDA 0.051696f
C2782 VDDA.t95 GNDA 0.051696f
C2783 VDDA.t4 GNDA 0.051696f
C2784 VDDA.t65 GNDA 0.051696f
C2785 VDDA.t33 GNDA 0.051696f
C2786 VDDA.t292 GNDA 0.051696f
C2787 VDDA.t92 GNDA 0.051696f
C2788 VDDA.t109 GNDA 0.051696f
C2789 VDDA.t43 GNDA 0.051696f
C2790 VDDA.t310 GNDA 0.051696f
C2791 VDDA.t80 GNDA 0.051696f
C2792 VDDA.t402 GNDA 0.051696f
C2793 VDDA.t298 GNDA 0.051696f
C2794 VDDA.t28 GNDA 0.051696f
C2795 VDDA.t312 GNDA 0.051696f
C2796 VDDA.t159 GNDA 0.051696f
C2797 VDDA.t6 GNDA 0.051696f
C2798 VDDA.t230 GNDA 0.063868f
C2799 VDDA.n528 GNDA 0.075861f
C2800 VDDA.n529 GNDA 0.041198f
C2801 VDDA.t229 GNDA 0.022707f
C2802 VDDA.n530 GNDA 0.022647f
C2803 VDDA.n531 GNDA 0.106245f
C2804 VDDA.n532 GNDA 0.204847f
C2805 VDDA.t69 GNDA 0.018463f
C2806 VDDA.t100 GNDA 0.018463f
C2807 VDDA.n533 GNDA 0.060995f
C2808 VDDA.n534 GNDA 0.078706f
C2809 VDDA.n536 GNDA 0.012309f
C2810 VDDA.n539 GNDA 0.012309f
C2811 VDDA.n540 GNDA 0.012309f
C2812 VDDA.n541 GNDA 0.021411f
C2813 VDDA.n542 GNDA 0.012309f
C2814 VDDA.n543 GNDA 0.012309f
C2815 VDDA.n544 GNDA 0.012309f
C2816 VDDA.n545 GNDA 0.02154f
C2817 VDDA.t219 GNDA 0.088038f
C2818 VDDA.t253 GNDA 0.011667f
C2819 VDDA.n546 GNDA 0.030232f
C2820 VDDA.t291 GNDA 0.024572f
C2821 VDDA.t255 GNDA 0.021556f
C2822 VDDA.n547 GNDA 0.10784f
C2823 VDDA.t254 GNDA 0.074677f
C2824 VDDA.t111 GNDA 0.047388f
C2825 VDDA.t161 GNDA 0.047388f
C2826 VDDA.t290 GNDA 0.076321f
C2827 VDDA.n548 GNDA 0.112944f
C2828 VDDA.t289 GNDA 0.011667f
C2829 VDDA.n549 GNDA 0.030002f
C2830 VDDA.n550 GNDA 0.090252f
C2831 VDDA.t103 GNDA 0.018463f
C2832 VDDA.t11 GNDA 0.018463f
C2833 VDDA.n551 GNDA 0.060995f
C2834 VDDA.n552 GNDA 0.078706f
C2835 VDDA.t74 GNDA 0.018463f
C2836 VDDA.t76 GNDA 0.018463f
C2837 VDDA.n553 GNDA 0.060995f
C2838 VDDA.n554 GNDA 0.078706f
C2839 VDDA.t91 GNDA 0.018463f
C2840 VDDA.t51 GNDA 0.018463f
C2841 VDDA.n555 GNDA 0.060995f
C2842 VDDA.n556 GNDA 0.078706f
C2843 VDDA.t49 GNDA 0.018463f
C2844 VDDA.t83 GNDA 0.018463f
C2845 VDDA.n557 GNDA 0.060995f
C2846 VDDA.n558 GNDA 0.078706f
C2847 VDDA.t89 GNDA 0.018463f
C2848 VDDA.t72 GNDA 0.018463f
C2849 VDDA.n559 GNDA 0.060995f
C2850 VDDA.n560 GNDA 0.078706f
C2851 VDDA.t154 GNDA 0.018463f
C2852 VDDA.t168 GNDA 0.018463f
C2853 VDDA.n561 GNDA 0.060995f
C2854 VDDA.n562 GNDA 0.078706f
C2855 VDDA.t53 GNDA 0.018463f
C2856 VDDA.t305 GNDA 0.018463f
C2857 VDDA.n563 GNDA 0.060995f
C2858 VDDA.n564 GNDA 0.078706f
C2859 VDDA.n565 GNDA 0.042023f
C2860 VDDA.n566 GNDA 0.032879f
C2861 VDDA.n567 GNDA 0.024411f
C2862 VDDA.n569 GNDA 0.021411f
C2863 VDDA.n570 GNDA 0.02154f
C2864 VDDA.n571 GNDA 0.02154f
C2865 VDDA.n572 GNDA 0.02154f
C2866 VDDA.n573 GNDA 0.031178f
C2867 VDDA.n574 GNDA 0.012954f
C2868 VDDA.n575 GNDA 0.172627f
C2869 VDDA.t220 GNDA 0.183089f
C2870 VDDA.t52 GNDA 0.18832f
C2871 VDDA.t304 GNDA 0.18832f
C2872 VDDA.t153 GNDA 0.18832f
C2873 VDDA.t167 GNDA 0.18832f
C2874 VDDA.t88 GNDA 0.18832f
C2875 VDDA.t71 GNDA 0.18832f
C2876 VDDA.t48 GNDA 0.18832f
C2877 VDDA.t82 GNDA 0.18832f
C2878 VDDA.t90 GNDA 0.18832f
C2879 VDDA.t50 GNDA 0.18832f
C2880 VDDA.t73 GNDA 0.18832f
C2881 VDDA.t75 GNDA 0.18832f
C2882 VDDA.t102 GNDA 0.18832f
C2883 VDDA.t10 GNDA 0.18832f
C2884 VDDA.t68 GNDA 0.18832f
C2885 VDDA.t99 GNDA 0.18832f
C2886 VDDA.t177 GNDA 0.183089f
C2887 VDDA.n577 GNDA 0.012309f
C2888 VDDA.n578 GNDA 0.012309f
C2889 VDDA.n579 GNDA 0.02154f
C2890 VDDA.n580 GNDA 0.021411f
C2891 VDDA.n581 GNDA 0.02154f
C2892 VDDA.n582 GNDA 0.012309f
C2893 VDDA.n583 GNDA 0.02154f
C2894 VDDA.n584 GNDA 0.02154f
C2895 VDDA.n585 GNDA 0.021411f
C2896 VDDA.n586 GNDA 0.034015f
C2897 VDDA.n587 GNDA 0.010117f
C2898 VDDA.n588 GNDA 0.172627f
C2899 VDDA.n589 GNDA 0.012309f
C2900 VDDA.n590 GNDA 0.024411f
C2901 VDDA.t176 GNDA 0.088038f
C2902 VDDA.n591 GNDA 0.032879f
C2903 VDDA.n592 GNDA 0.048485f
C2904 VDDA.n593 GNDA 0.053331f
C2905 VDDA.n594 GNDA 0.027132f
C2906 VDDA.t268 GNDA 0.01812f
C2907 VDDA.n595 GNDA 0.024998f
C2908 VDDA.n596 GNDA 0.024411f
C2909 VDDA.n597 GNDA 0.02154f
C2910 VDDA.n598 GNDA 0.012309f
C2911 VDDA.n599 GNDA 0.012309f
C2912 VDDA.n601 GNDA 0.012309f
C2913 VDDA.n602 GNDA 0.02154f
C2914 VDDA.t185 GNDA 0.017703f
C2915 VDDA.n603 GNDA 0.024946f
C2916 VDDA.n604 GNDA 0.027166f
C2917 VDDA.n605 GNDA 0.012309f
C2918 VDDA.n606 GNDA 0.02154f
C2919 VDDA.t187 GNDA 0.032451f
C2920 VDDA.n608 GNDA 0.029969f
C2921 VDDA.n609 GNDA 0.010117f
C2922 VDDA.n610 GNDA 0.10893f
C2923 VDDA.t186 GNDA 0.090467f
C2924 VDDA.t41 GNDA 0.081236f
C2925 VDDA.t269 GNDA 0.090467f
C2926 VDDA.n611 GNDA 0.012954f
C2927 VDDA.n612 GNDA 0.10893f
C2928 VDDA.n614 GNDA 0.012309f
C2929 VDDA.n615 GNDA 0.02154f
C2930 VDDA.t270 GNDA 0.044759f
C2931 VDDA.t42 GNDA 0.012309f
C2932 VDDA.n617 GNDA 0.034921f
C2933 VDDA.n618 GNDA 0.058656f
C2934 VDDA.n619 GNDA 0.120237f
C2935 VDDA.n620 GNDA 0.167134f
C2936 VDDA.n621 GNDA 0.015352f
C2937 VDDA.n622 GNDA 0.054191f
C2938 VDDA.t273 GNDA 0.022437f
C2939 VDDA.t202 GNDA 0.022437f
C2940 VDDA.t200 GNDA 0.01212f
C2941 VDDA.t31 GNDA 0.012309f
C2942 VDDA.t208 GNDA 0.012309f
C2943 VDDA.n623 GNDA 0.035949f
C2944 VDDA.n624 GNDA 0.061596f
C2945 VDDA.n626 GNDA 0.012309f
C2946 VDDA.n628 GNDA 0.012309f
C2947 VDDA.n629 GNDA 0.012309f
C2948 VDDA.t285 GNDA 0.044759f
C2949 VDDA.n630 GNDA 0.012309f
C2950 VDDA.t283 GNDA 0.018605f
C2951 VDDA.n631 GNDA 0.015358f
C2952 VDDA.n632 GNDA 0.054185f
C2953 VDDA.t184 GNDA 0.022449f
C2954 VDDA.t267 GNDA 0.022449f
C2955 VDDA.t265 GNDA 0.01212f
C2956 VDDA.n633 GNDA 0.015358f
C2957 VDDA.n634 GNDA 0.0734f
C2958 VDDA.t279 GNDA 0.022449f
C2959 VDDA.t246 GNDA 0.022449f
C2960 VDDA.t244 GNDA 0.01212f
C2961 VDDA.n635 GNDA 0.025579f
C2962 VDDA.n636 GNDA 0.064062f
C2963 VDDA.t245 GNDA 0.067513f
C2964 VDDA.t300 GNDA 0.047388f
C2965 VDDA.t409 GNDA 0.047388f
C2966 VDDA.t278 GNDA 0.067513f
C2967 VDDA.n637 GNDA 0.064061f
C2968 VDDA.t277 GNDA 0.01212f
C2969 VDDA.n638 GNDA 0.024926f
C2970 VDDA.n639 GNDA 0.040792f
C2971 VDDA.n640 GNDA 0.015358f
C2972 VDDA.n641 GNDA 0.054185f
C2973 VDDA.n642 GNDA 0.039869f
C2974 VDDA.n643 GNDA 0.024926f
C2975 VDDA.n644 GNDA 0.064062f
C2976 VDDA.t266 GNDA 0.067513f
C2977 VDDA.t22 GNDA 0.047388f
C2978 VDDA.t20 GNDA 0.047388f
C2979 VDDA.t57 GNDA 0.047388f
C2980 VDDA.t26 GNDA 0.047388f
C2981 VDDA.t183 GNDA 0.067513f
C2982 VDDA.n645 GNDA 0.064061f
C2983 VDDA.t182 GNDA 0.012504f
C2984 VDDA.n646 GNDA 0.025311f
C2985 VDDA.n647 GNDA 0.046946f
C2986 VDDA.t25 GNDA 0.012309f
C2987 VDDA.t303 GNDA 0.012309f
C2988 VDDA.n648 GNDA 0.035949f
C2989 VDDA.n649 GNDA 0.064366f
C2990 VDDA.t379 GNDA 0.012309f
C2991 VDDA.n650 GNDA 0.035949f
C2992 VDDA.n651 GNDA 0.061596f
C2993 VDDA.n652 GNDA 0.044177f
C2994 VDDA.n653 GNDA 0.026154f
C2995 VDDA.n654 GNDA 0.024411f
C2996 VDDA.n656 GNDA 0.02154f
C2997 VDDA.n657 GNDA 0.02154f
C2998 VDDA.n658 GNDA 0.027132f
C2999 VDDA.n659 GNDA 0.012954f
C3000 VDDA.n660 GNDA 0.10893f
C3001 VDDA.t284 GNDA 0.090467f
C3002 VDDA.t378 GNDA 0.081236f
C3003 VDDA.t24 GNDA 0.081236f
C3004 VDDA.t302 GNDA 0.081236f
C3005 VDDA.t30 GNDA 0.081236f
C3006 VDDA.t207 GNDA 0.090467f
C3007 VDDA.n661 GNDA 0.012309f
C3008 VDDA.n662 GNDA 0.02154f
C3009 VDDA.n663 GNDA 0.02154f
C3010 VDDA.t209 GNDA 0.032451f
C3011 VDDA.n664 GNDA 0.029969f
C3012 VDDA.n665 GNDA 0.010117f
C3013 VDDA.n666 GNDA 0.10893f
C3014 VDDA.n668 GNDA 0.027166f
C3015 VDDA.t206 GNDA 0.018605f
C3016 VDDA.n669 GNDA 0.026154f
C3017 VDDA.n670 GNDA 0.044177f
C3018 VDDA.n671 GNDA 0.015352f
C3019 VDDA.n672 GNDA 0.054191f
C3020 VDDA.n673 GNDA 0.046946f
C3021 VDDA.n674 GNDA 0.024926f
C3022 VDDA.n675 GNDA 0.064073f
C3023 VDDA.t201 GNDA 0.067513f
C3024 VDDA.t85 GNDA 0.047388f
C3025 VDDA.t1 GNDA 0.047388f
C3026 VDDA.t314 GNDA 0.047388f
C3027 VDDA.t364 GNDA 0.047388f
C3028 VDDA.t272 GNDA 0.067513f
C3029 VDDA.n676 GNDA 0.064073f
C3030 VDDA.t271 GNDA 0.01212f
C3031 VDDA.n677 GNDA 0.024926f
C3032 VDDA.n678 GNDA 0.124452f
C3033 VDDA.n679 GNDA 0.145292f
C3034 VDDA.n680 GNDA 0.692647f
C3035 two_stage_opamp_dummy_magic_14_0.Vb3.t2 GNDA 0.014695f
C3036 two_stage_opamp_dummy_magic_14_0.Vb3.t4 GNDA 0.014695f
C3037 two_stage_opamp_dummy_magic_14_0.Vb3.n0 GNDA 0.047335f
C3038 two_stage_opamp_dummy_magic_14_0.Vb3.t5 GNDA 0.014695f
C3039 two_stage_opamp_dummy_magic_14_0.Vb3.t0 GNDA 0.014695f
C3040 two_stage_opamp_dummy_magic_14_0.Vb3.n1 GNDA 0.047335f
C3041 two_stage_opamp_dummy_magic_14_0.Vb3.n2 GNDA 0.260957f
C3042 two_stage_opamp_dummy_magic_14_0.Vb3.t1 GNDA 0.014695f
C3043 two_stage_opamp_dummy_magic_14_0.Vb3.t3 GNDA 0.014695f
C3044 two_stage_opamp_dummy_magic_14_0.Vb3.n3 GNDA 0.044386f
C3045 two_stage_opamp_dummy_magic_14_0.Vb3.n4 GNDA 0.790392f
C3046 two_stage_opamp_dummy_magic_14_0.Vb3.t6 GNDA 0.051434f
C3047 two_stage_opamp_dummy_magic_14_0.Vb3.t7 GNDA 0.051434f
C3048 two_stage_opamp_dummy_magic_14_0.Vb3.n5 GNDA 0.181328f
C3049 two_stage_opamp_dummy_magic_14_0.Vb3.t24 GNDA 0.072742f
C3050 two_stage_opamp_dummy_magic_14_0.Vb3.t22 GNDA 0.072742f
C3051 two_stage_opamp_dummy_magic_14_0.Vb3.t27 GNDA 0.072742f
C3052 two_stage_opamp_dummy_magic_14_0.Vb3.t9 GNDA 0.072742f
C3053 two_stage_opamp_dummy_magic_14_0.Vb3.t11 GNDA 0.083944f
C3054 two_stage_opamp_dummy_magic_14_0.Vb3.n6 GNDA 0.068153f
C3055 two_stage_opamp_dummy_magic_14_0.Vb3.n7 GNDA 0.041882f
C3056 two_stage_opamp_dummy_magic_14_0.Vb3.n8 GNDA 0.041882f
C3057 two_stage_opamp_dummy_magic_14_0.Vb3.n9 GNDA 0.03886f
C3058 two_stage_opamp_dummy_magic_14_0.Vb3.t20 GNDA 0.072742f
C3059 two_stage_opamp_dummy_magic_14_0.Vb3.t16 GNDA 0.072742f
C3060 two_stage_opamp_dummy_magic_14_0.Vb3.t13 GNDA 0.072742f
C3061 two_stage_opamp_dummy_magic_14_0.Vb3.t25 GNDA 0.072742f
C3062 two_stage_opamp_dummy_magic_14_0.Vb3.t28 GNDA 0.083944f
C3063 two_stage_opamp_dummy_magic_14_0.Vb3.n10 GNDA 0.068153f
C3064 two_stage_opamp_dummy_magic_14_0.Vb3.n11 GNDA 0.041882f
C3065 two_stage_opamp_dummy_magic_14_0.Vb3.n12 GNDA 0.041882f
C3066 two_stage_opamp_dummy_magic_14_0.Vb3.n13 GNDA 0.03886f
C3067 two_stage_opamp_dummy_magic_14_0.Vb3.n14 GNDA 0.042711f
C3068 two_stage_opamp_dummy_magic_14_0.Vb3.t8 GNDA 0.072742f
C3069 two_stage_opamp_dummy_magic_14_0.Vb3.t10 GNDA 0.072742f
C3070 two_stage_opamp_dummy_magic_14_0.Vb3.t14 GNDA 0.072742f
C3071 two_stage_opamp_dummy_magic_14_0.Vb3.t18 GNDA 0.072742f
C3072 two_stage_opamp_dummy_magic_14_0.Vb3.t23 GNDA 0.083944f
C3073 two_stage_opamp_dummy_magic_14_0.Vb3.n15 GNDA 0.068153f
C3074 two_stage_opamp_dummy_magic_14_0.Vb3.n16 GNDA 0.041882f
C3075 two_stage_opamp_dummy_magic_14_0.Vb3.n17 GNDA 0.041882f
C3076 two_stage_opamp_dummy_magic_14_0.Vb3.n18 GNDA 0.03886f
C3077 two_stage_opamp_dummy_magic_14_0.Vb3.t26 GNDA 0.072742f
C3078 two_stage_opamp_dummy_magic_14_0.Vb3.t21 GNDA 0.072742f
C3079 two_stage_opamp_dummy_magic_14_0.Vb3.t17 GNDA 0.072742f
C3080 two_stage_opamp_dummy_magic_14_0.Vb3.t19 GNDA 0.072742f
C3081 two_stage_opamp_dummy_magic_14_0.Vb3.t15 GNDA 0.083944f
C3082 two_stage_opamp_dummy_magic_14_0.Vb3.n19 GNDA 0.068153f
C3083 two_stage_opamp_dummy_magic_14_0.Vb3.n20 GNDA 0.041882f
C3084 two_stage_opamp_dummy_magic_14_0.Vb3.n21 GNDA 0.041882f
C3085 two_stage_opamp_dummy_magic_14_0.Vb3.n22 GNDA 0.03886f
C3086 two_stage_opamp_dummy_magic_14_0.Vb3.n23 GNDA 0.044462f
C3087 two_stage_opamp_dummy_magic_14_0.Vb3.n24 GNDA 1.22508f
C3088 two_stage_opamp_dummy_magic_14_0.Vb3.t12 GNDA 0.089166f
C3089 two_stage_opamp_dummy_magic_14_0.Vb3.n25 GNDA 0.309961f
C3090 two_stage_opamp_dummy_magic_14_0.Vb3.n26 GNDA 0.918527f
C3091 bgr_7_0.VB3_CUR_BIAS GNDA 1.64457f
C3092 bgr_7_0.NFET_GATE_10uA.t0 GNDA 0.01675f
C3093 bgr_7_0.NFET_GATE_10uA.t4 GNDA 0.01675f
C3094 bgr_7_0.NFET_GATE_10uA.n0 GNDA 0.047127f
C3095 bgr_7_0.NFET_GATE_10uA.t18 GNDA 0.016332f
C3096 bgr_7_0.NFET_GATE_10uA.t6 GNDA 0.016332f
C3097 bgr_7_0.NFET_GATE_10uA.t14 GNDA 0.016332f
C3098 bgr_7_0.NFET_GATE_10uA.t19 GNDA 0.016332f
C3099 bgr_7_0.NFET_GATE_10uA.t5 GNDA 0.016332f
C3100 bgr_7_0.NFET_GATE_10uA.t13 GNDA 0.016332f
C3101 bgr_7_0.NFET_GATE_10uA.t12 GNDA 0.024143f
C3102 bgr_7_0.NFET_GATE_10uA.n1 GNDA 0.029878f
C3103 bgr_7_0.NFET_GATE_10uA.n2 GNDA 0.021357f
C3104 bgr_7_0.NFET_GATE_10uA.n3 GNDA 0.018081f
C3105 bgr_7_0.NFET_GATE_10uA.t15 GNDA 0.016332f
C3106 bgr_7_0.NFET_GATE_10uA.t8 GNDA 0.016332f
C3107 bgr_7_0.NFET_GATE_10uA.t21 GNDA 0.016332f
C3108 bgr_7_0.NFET_GATE_10uA.t16 GNDA 0.024143f
C3109 bgr_7_0.NFET_GATE_10uA.n4 GNDA 0.029878f
C3110 bgr_7_0.NFET_GATE_10uA.n5 GNDA 0.021357f
C3111 bgr_7_0.NFET_GATE_10uA.n6 GNDA 0.018081f
C3112 bgr_7_0.NFET_GATE_10uA.t20 GNDA 0.016332f
C3113 bgr_7_0.NFET_GATE_10uA.t7 GNDA 0.024143f
C3114 bgr_7_0.NFET_GATE_10uA.n7 GNDA 0.026602f
C3115 bgr_7_0.NFET_GATE_10uA.n8 GNDA 0.029239f
C3116 bgr_7_0.NFET_GATE_10uA.t11 GNDA 0.016332f
C3117 bgr_7_0.NFET_GATE_10uA.t22 GNDA 0.024143f
C3118 bgr_7_0.NFET_GATE_10uA.n9 GNDA 0.026602f
C3119 bgr_7_0.NFET_GATE_10uA.t9 GNDA 0.016332f
C3120 bgr_7_0.NFET_GATE_10uA.t17 GNDA 0.016332f
C3121 bgr_7_0.NFET_GATE_10uA.t23 GNDA 0.016332f
C3122 bgr_7_0.NFET_GATE_10uA.t10 GNDA 0.024143f
C3123 bgr_7_0.NFET_GATE_10uA.n10 GNDA 0.029878f
C3124 bgr_7_0.NFET_GATE_10uA.n11 GNDA 0.021357f
C3125 bgr_7_0.NFET_GATE_10uA.n12 GNDA 0.018081f
C3126 bgr_7_0.NFET_GATE_10uA.n13 GNDA 0.029239f
C3127 bgr_7_0.NFET_GATE_10uA.n14 GNDA 0.67829f
C3128 bgr_7_0.NFET_GATE_10uA.n15 GNDA 0.024928f
C3129 bgr_7_0.NFET_GATE_10uA.n16 GNDA 0.018081f
C3130 bgr_7_0.NFET_GATE_10uA.n17 GNDA 0.021357f
C3131 bgr_7_0.NFET_GATE_10uA.n18 GNDA 0.029878f
C3132 bgr_7_0.NFET_GATE_10uA.t3 GNDA 0.038251f
C3133 bgr_7_0.NFET_GATE_10uA.n19 GNDA 0.366469f
C3134 bgr_7_0.NFET_GATE_10uA.t1 GNDA 0.01675f
C3135 bgr_7_0.NFET_GATE_10uA.t2 GNDA 0.01675f
C3136 bgr_7_0.NFET_GATE_10uA.n20 GNDA 0.069531f
.ends

